-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
v+TOCidNyF9wWiYjrVwGF6wNP2yzfW+j4BqfV9eXqPOIExt4nt+HKRKTxG+iNSz/yJEKp8bE7ak3
PAP8l/b7QkAy9yc+kDvVAL6iXzdJXUhKXsMieKClt6rBxC71vDoJxo0TXNlVkA81opD0nnb2ZWPY
YuBry/BiWFY8AhYpu5INX3pZNzEuCT22pxCWPQopkGqm6cp26BD55ikDQG+J4U9FGyP7czqAaN5y
n/FwnZErfWvqUWQd8IABDbWa0HkT6x/1Sr7zQ3JzHUhbNYKd+W1xoGutbQvz/i4D1SP2y9b3t/1g
Fnl9m4Pr8bzF41jmt8lRTiu+g8kckVre5jfKeA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3360)
`protect data_block
/O1J3/GOyfo1otPmYL7IJNEaop5jtqa1Ofu56CwFrXBewjQNsDABJuZeAQMxB7TcYwUS8zsF/us5
0w4MkH3Z5YmST3KjhqhkQUK9TLkZJ8T03JWg5k8nCmIJts+jq/Cj2txRpqjDTS1jQWXV+XnB4xlc
QXjmCHMnMX0hiJbYgYmAgVQ/j8vcjvBVfAayLQXjXXlIJnfxRzqnVant8JS2CMRfCR9CSwxWfrav
rLM/H9i3aIzOMiQsH82d1X7P0pwBtf/ICxg3MFfOA9U6CGeBQlRSG/jn4OnMexdLJ9oX5xqQFQsV
L7fw8E7HCvMQ7O6N1PmCw8fu7yaQOwBbk0lWPgP/E9rwR6tYhA6Sq419dtQq9JqUz/OppyPDgLEG
32awN/0v7YuzJwHK/t1x5iN9hlWyQ1jSDL1NVDHZvFlf+Qi8I7Fgmoxc3R8Jd0L3dtbXnTX9VO28
pAu2F7VJInKItJrzsY+zQfSauwURZfPNoDZX4vSJ1Cea1ORVu9Kj8+nuPQnJibu5bhJ4H8zB8NxW
Hj1jQgDyvgpRF+50J8wtlIbNQLmXh5mOoVD0qfncfzaGwguJ+CnD3ty34A9zPd7gSQB3AD6JPyg9
mimUIKfDX0H8nDEB3ae+E6NKmtn3FuYWcFlQA14kR3Rm7QctWaEnqyY5GaCBJlDmNz+2Trva/hJn
oIISTjBd8ZBGj5ODg2/3o0hM6MxruyCI0DdDxSJwQ8kzwXK1eSbrLEmTY/BZzBvzAVkbR1tZEUIW
sAnqdDoAnGOtBlst2A2rJ5KlOohdM7h2c3sav02VGpWTUNgPyDk7I3Iirl2LnuJ9QI30M9zKnqWk
8NcQVQmETtQ+mAhosQJ8b39rJjqnS/Bjr2WgBs8nzWsN3j5WGK5uTWn26GIu8GiZn2aEKENMHV9n
S4R59EJrHHxFdmjiSfS75/BFkN2APBuNMbxf+0LL4t8yigACdHbXrDCVaYbFe7MsKzyaaqOV8meF
fES1DkXJJT0FwN0YY4qoNj2luVR0VIDuiGUw9Cv/0eoiuayCv9woyFOBZ+0TrDl8xq2tRwFDMflK
Cjsj4AAbuyUL5hQTx4Rhl1UiE5cUDPHhDcUajDP8+yTfn/BZs6c4XUD6D2B5WuvMDooDTHGDE8W4
68KiT/p374eOiosGt7bNWUVJOTmZc+nkCgoH0Dy+dJGD8WbfWJdKtzhNu+8FXbyQK8VrFxM7EAIx
7wsDNwKZdpaJWqW7rfygI+Bak3z1coZyxG2CCMOjyKKAzdNUnYeg74rc2ydwRzUuZgHbtGbdXkSA
FvGyMdiJHUJ/ZQjN2XdK74LYlzU8wfmFsztGVBk6giV2xvlv3uoHUIaPXWSn3L1z3x/9v2JmYlZm
qMmF0xzYuJEyRcwCQQWMM+V/6Lz7Uvb6/6IWEhEtq16+C9V7MgMd/asnAfX6/yc3Ojp4C2vwnJh1
KMOxE4qDqr1N8nbEHvjLYeH+bTxfQqKMVqczGTrWN2I5IwT0x+pbPJ4IB+K1geCv0xa8rhvbfcdx
NVKO0OoLh52ywLVXHftgS+p+FRMU2moPKrGWYHXVjH8uHmHDMxfzTfZM/EMKxsH8CB2ymzZEPwf7
W5UB3jLJ7mUSsLbAbNn5bgeHZaYbiIQf+yQvd5kpzSzz7zSUtd24QyeBzbPyZNP9LICGxWA6po9m
QxPEUhVH2LNoaVBtK+RPeEmLNgh4JQG1hUYVjzVm5kmiRtpRpbJXVTvgQjNdoHlM6/UQ0TutL/3e
KzDtj9oz7TkTGoHFxlgqj0cKJHxaU6F4H7CDndcFyDWVxFjCcoKs6hmAzPQMiAahctWlm52SMV2H
3FOHwKghG+Ntykf7PUfN9NQbIOTIhY8lvakL1ZmfuIdXfAUdK59LGH4kyARuOjyQAwx7wstqefif
bQr7FyVmNKPpLtQdU93ob+DM/PmGToN3nT7mRVQriXFE4XPEtNb7fZKMOjbU/BnapQUzdOnLiPm1
bHpsHOa2Uk/NNp4wQHpxtbVUQnDRg9kwH0rsuf91suUMXbPDEPrEW5H5v9KyzG/mgwDPurvjXN0b
9Ra6v7FMG+i8kuBVVBBCjl38s4g67wDDleu7zEAWbsEmASt7GLPJIGEIJz2yLIU+gKOmZiSbzR0N
QzPMOIR8PT+0D5INrzDbYprOTtB5z4cppM8Gw5ZoImqpKQFZGArzT+EFYzC1ZUrNhOZILzkwXMOZ
iVkXSu5VPM8oPrGqV5NuNW7hEP1vSS7J5dT5wrfSov641pZe07IsertwbNxiuko4NNruiI8smCY6
qCx8XWrnru6ssFCIa+APG/8ZOapohkCCJSSZ3DcAyFLDQVxyCr2fuGaCFDF3KGAKRiAmhsybbQZp
z9IkD4IfQLbIdJystNH/nNo5zdVkTuY0Fp9ilOVxfk4hNxawMhYQx4xxzqHpooesIxb3Bs05boVy
LA1iVsvXSufW49UGKfdFseA2QNqKgsErbx5SeXX7vJlCjz/KH671O0I5Frd03n3KrOkd4jscYfdW
F3CXTqIEuEziK2PGQQ4kCbyGOGh1ZNW8/1nHcRmTi+fLRa6cl9Qq4XN6WKcGyuKjvbuS46X6Cpl2
SrIUxL4SgppyO/+Y5FQPc2NDY9UNWbd+5p6wpLw2fzfImwWZNKN6bVpOKHYhLe8s9yB2jlTuMeNh
IozdJddCnNHLr+Au3SaLbK6lxLkeu/DBhzl4pntHF1mYcKE61pPvh+5j1cp1qwobix823+3Jtack
OgijWvTFi+UQSTyBwZaYigtJHmBZpmx0DlWm9x8NSAbKGEXQtjqpaut1E/uY1dpRIzvQINI6S4GM
/l5v/kPDkShWiMXDJw9QcyKxyc7TFuWNNLOqmsjF4qQeZdTzeB8XU7NCetHv3Ll2pEsDp5NES5b2
bFO1eATDF4mPvlXkd+/OHCOObEPHvnTyWMZ6+eivN1n5S7Ma10dhlHOx1XgACb0j4cJiVLi6h9wi
hqGFWFJliA2V/6AfVV/q3JxVU9pVsE+JazS7B0ENszoYYT8jwAdY/ZLe5gNfjl5xlu0MF0FFvfAf
qasQcq7P66q7rm1imr3p9EU6/ZNEULm5s2KdaQGU6PCXsrp8vCCx+obx9QJG29nvAl98mSzJeyag
gn+FodDeoZveQ8vjdhxPGXqvNxINtW7cv7d/SI66YpJwbUs2skSi1ic42BtHGdvlO8bGF+90IshC
KGqoG+voqSVlvjNR8rORnnQ3zJUB/qUH5bXuYsb0b8I7TTsx/hyyxTCaioMR0xAKkRfxZiCBTHut
voBaFIpMol/fJHW7sZvOlnD7uQmCeh7EIE0wV315WUOXApJxRkWooTWutlu+BArCTMjQkyQJd76T
VWxnzupLySV6K250sTwR/Oq1riga1XODdf0h5CECqlthVllCZaHHE83a4465+F8V8FFCEf89b8rU
wVdiULJIoE7Y5h1GpkgPkWTUx/wQmBr82yRffDwVuVXOyKewOFS9ozWoTFmIUZw/tmHrWNITjpTc
St7PWyNxauGzgMPeS4mQEawCq55qal0KGSlL+yZrCsNSwB4ZoqWzMFgR3YSJk40L34wb3BochNGr
wRvk/NGqxW2UOtB7yXRE4azj30FJQ2Ji6YAb9uSYpCU7I83VZdN3QfsrNm9T0jt0dbpVfVZ5jIHF
RvvRqoiufmH24JUwNbjOXc0zVyZkcCn8+3qvwHyY6vJY1D3tGwwnCiByXuhdubNCCnzcrA78A986
6kCioxexMG1499sy+we0MGZD+SAu1PaElBHkk+wH3Gf6nVqGsfNUoST+2qJL5YBBPn2I7rSUM1Nh
6n2jU5huoFrGKZhPmX+UZPO1ak2AK0eKfy9AtoGILey/VJTi0+GymX1AIiH+ZVTd3YQOnStVCbd+
Gk2ByHLTfmsAoY5h7N2GEw5ZBJwZ0yFEsTsOpy3fsoFSLrIyifvaMI+EIrPG/FCwC7/8eRuaUpYY
Q8JdlVnOTqzMrl3EyXx5YmV6lz1QHt6phHdsCO61zQw8TZLXWe2slQNjyfjpIXKk1wwJffft6UEo
0JKjp317igcHsw4J0WO//NdOiOdPY/QfMRrAYJqB3plCehLSDZSa2uBDyiQl33R2g6uR6Ow0u8f2
us/thGGUtLNBV8HumCTcQ1vJH6+zVH9dtcqpBL+blR3sBLoKRsYyOkJWJfnqiApz14f/UdEBGVZM
j73ENPQ/xbaCBL6mufTqYCH12iTvMEUedSFc82yVXESRneq5aPZBZeY/NA4ZtOssdj6ZWkFUWXsG
e2yXc9NHYTeQUunf/pWGiJlpEMwzvuZBKn9EWd+Xe42pgebj8px6sdTbbg2O9XH8DaBjrZWVOUMP
Nc6aRHPgXrY5RX4pBuduCKPvHbm+w/0OtESARONxa7Po6hmjcBRBD2leqDX9Sx+PsVDeVwTY3pHU
FlR5C8Q+9sV9WKFjpW2BsAaBykUO2zGIiQHz1q/sJYvYB2Sb+vA7qm2TA0TBGGZxEggSNt2h
`protect end_protected
