-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Sl2YmNJM1YhrN/VKaoVwaHC3oSre76RRjqV8TIBrfOeFJu/XhuRo68bt0/NKIL/giGSQ2uDfD5s7
0LrrLnz+gSKb31rWbSXHzJpPONtBoNnBpTWoCL9IGwZ3jljuk11Fb/G81kZQGVuxmU7OAEMno6nf
zxfmB415iaVh19xvD4XLyQ40MQBEHTc0RjLb5mt8QkcmRndrlTTG2WQ4t7AR1iCVrJtgKUlbcVCX
iVlmByMKOHyIL+GqV1BbndXveTz2meIQTmtWOqlKnceXW52cZHGkmb0t0GPy8wRgvdcqaSCHdkU1
ioXjDbZxBSxex1QD3n8MqfNK1CsAAlCjx1qz2A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
M70SKUxuzafh1Ogce3ytB4YC5tRKMLxu0CeL5gWKZSVsVs9jxT4TZCeXSJsXNKMVbiP7rM4gTP7s
7XW5HTwRNUtOTb+TtfhOyfpjHOJShC7AnE5bJyj7X/Si1CY39F97TgD/o99i/1EIS7Hc3v83om+b
Mumnos11q1vzPCwzHtzBcSRpSwSwdqr7kfNCXArJ8DQiLpYdqh8hW4BcR6nDa+8why0FLKvL0OKe
su2qcrXvkvUMpnKGfm8gUCazrXVFj8+5sCmTAMO+BCPFh8eUJggTxT1xNwG9FsaPRuelWgvfO2sw
b9+dXfMGOAHI0bqeNuCyBVZ8xH6+btSW9u259labcQci3BfmPxQED6pldK+dGGyDWDbrdIXZZgaa
8TxsOd5WwTacV3My1fL/RlDd4jHD6mW7pDaCePEYwWxHFkD7VWvDQkYwOpSxSC/UNhYJYr8vmJ+p
giVRPeCMPOd63A1cCcFAPHmoG+Pdq9ZL5AjskBGTSs/nDOKiAubHoiJW+m98RiSIe24qmQUwqnDF
6frs+YpGu/a0YwCfGWvt1L8tNIL58BDgoXa0m+oCa3n6V7r2f2F7juRCyWTvp8FHZirxuLAop8ws
ci711OHsqXiv7YnAtSNcqzXrveLqO6wMP/cOktnxSoQi5sepkKIlTRV+/GZH6kHy0p+M/WNT5XHK
gd0XNOYLuYB3prTWZrRsI8kAq0/K3fhfFhe5UbueSSjKn722DEUfYCJ+9Q4IK7FsaJbanSkXLVur
yM/2tfg6y0vSpvB/BCJuPTHuCgQQjlY/HZYbK0qAuR8B3F4yU+zIRQJHLBPTXD5HVgx+vSeiDUAe
VUzuPXROuvnvekSodNh3+leW+7V0cpEDybBHz9r1IoVRWmJI/eA/qWYjCQVZXjd4PcIEbICKjoSF
7wOqEiT0QQfqpqpoWE/bFuKkyQ2HFy5wzPILIGFe4D2yVMUgzlGuc5ZsQJNIPcQXr0yL0d9tX78t
oaTQpr9oRA5VJYn1bnYhkEmGPFEbSJoiwK2RcQe/4qydbh0mxwtINiTW77vJvWAiNQ7+LSpOq4oX
spAecFWRoy6MQ+n1jWJGXyp5WSYAsbNW+Ep9WAuWC2OJMxJrH8THNa4JHW78hivCVUEulcSTlJfi
wXhBsc/hW1mZBS4F2xUeabwHbQ4xGAmz4GfgWntCMi8K0LRYyu2wMHUjZmxHDqtl/e1xDPeLfK1h
cXiM2EyFD+p3eMPMrHOwpg2OaiHeezdBTXiBv2r6EpqqTMTVZQ9xGyh2XE0V+pzBtN6T1Adb2voi
FUTdqaXr5y9fN7cZaftC55MT9TeLUyUACHMSDYEgX41BIBYkQ3LPsVnI4Q1Is7sav5ZrlOtihfgv
4C6Umb05kVyB/LiggmUbshhb9kK7eDUt1J1LAJ7AL3sGSU2qjDUVdvC/8uF0QfJ3hIGWYOg8B/lo
6ikwdiqkJO1L1fNT+C0OMCgngEjAfACJb3Edi14O/xsJvzjlMAhYUgaJcCq3U480TGT1/Q1x8da9
zZJBTADPTsOcMWNHR/cUd70GxW7N9CqdCc2/G+8O8kGlMaUGIBOYNMzhw90HrU/SYwGt6ui1cndK
unYoLsH2v7LT4L6rk0LeFwPWOzgk/sahIgIasAXSPj7t09sjrVvKb7F0WPoY8bupQ5ZyW/W1NwmZ
lftJxbTviFKOhmik+bvZZYIz/EliCfqFeEq/wAN5MjpFrC4Hh+SxG3OVOHzKkhPz4X08BNsKbjwX
790I1O+iBKPz6Dl2GNi00x3rwB+r60Qh6U0zWLDeJnVbeI/D1zr9ToCVTVxCAgB14nzlksXCgOhL
Edzzig8/t6ks2brNd7MOUcSiLKEhZQRnaal+A9xLGS+u5b/UwDWPxWAkXYQWDUKyoDgQ9R655LA/
foZqjeasxG5Ejy8Vd96wrdQRMERQC0aN0zvEA2Vrld4KZZFGq1YmWl/yn3tmjnJCjk6mhDHuOKET
8pfiRt/JWpJtmlaP+EDb9vWxt7NRNy2ACPQzsvxO40dc4K7BrIyo4PK4uegPC+bJiPuHw6Oas2Rb
ngfyFSos04lyDwUHF8+FkmfOSu7oK7aMtrZ7SIlFWkVMQ1wkuuNTbq5UJIIkM0I/u+q626y/N3vr
XBLSYGlW/G+8dGAnY5YiGxTfqUXFriad1cmRmDoHt0ntwC8l7gJbFaq4hYMtmhSkMoFJtyJKrP+n
olxl9ctAZ7yz4cob9rf8g4m0DERQSn+E/UIlb5BKu16Dr8NuF3pRlCptBRRgA8fCwSWcLh42SDCV
Zdyii7fKgVaIE7r0kpifEF8NDObMZ/hg/+1MdumaKueUHahF+pe2lJ6XhET7p9xBzy02oIE/X7i9
VyBAOlihrutVwfhy88oXKtMt3A0GOjSkzngMMN26UapxvxG1/KADNakMMRjGVHDnsDgVfvpNjcAt
b37jxtmS8VnEbNybtvnqOiGpw2hB15blEfgScPsXZVk39Y1eKmoLH3o4s0YQQ+/7eA4tjYjEzh9g
9aNhLxuRPJx9Z4P8BZoMpBJEmTkkcxkC5X9HOeiQLvAu6/32n85xmfEFD67TVcRs0vMAvnGQcSX3
nj6qhH3aZNCEaAS0VjAFurCg7vzo8KLZM1Qrx+fJROweM4gcSd7e+Agsbf6HJHBwKBTUmFA7aWkF
5yx0SQhrdXlJMwz9nb4J4rgFs4UCJgB+3N+uX5TpIiaS3jMAiYAiBy1ViMgU+LRQdLI7JcxSijYV
FopncLY/yxi1FGO0ZJz0I4zOgPX1NROSGRZjHctB6F43FxU5amVOOxKSCOB7TPBDMU2MbSKUJHia
mO1GFp1EWOIGybBaqsEBHCvpKLHCT5KRO44T0fFEPOAEbEDD6E1z6Fd3k9lxfo+UxItXZ9e5kWzR
nZuhLcc4uP2ORP/AdDXu85KQIZSYT6Q36uyPVwcFpDDiifFzlQ9MCYRpsBTR+KVDyXFBH9cOQGB/
XB6sDdCkzmTnMkKZTzsSq6yNm/7sYoGTxM2Ks2J6CFm5o5KBZP0zkneRNpSYXgvjxc67CPzjBqzX
zF9jxE3hMTnHzIioZyV9h9JZQF3sHWv4xoQE9QNIDVUqAj8Ym1wUrt2y09Gnp+eouNnQty3Al1Zb
IjiT8jbB/4tq10FLcFc4pMujkxN7Bba9vGnFlLbSJG/TZqFxylllZtue0s19fusWmSqYpK1jBFG8
/0sTQZi1fHM/U/DCLcIxrG8djMF4R6mn8gecpypzDdo9p/NeJeiuEoxntAkMjUlxqbS2kdTUZbpa
WLoQCzm42Ak0DmBruv+OQdInPWj01hmohX1opaj+hvzEGWXY8L2MraFlsHPY3iXxFUhlarWT32+v
BXzKIrSTSVO4ky90Tk368lzww/Uz8FFRGl8xBP9mbcxR9UgACVuz+JgSnR0aWkTDsnuPVSBHtjLJ
sXBXxB3YpHErMzp1PptqVrYASTiTkSgIghUFnP/FK4srrLlswCpUOatxd0gROPgX0D8kz8cKOu5d
rFg1RlBCosvkQGRH4W7QsECQMHOtd1B00iktujmLkI6h7RPB8VKb0tB2Of6f5Zw+Ve19piZF9W3p
3wUzb2MiokEuhsXhxnBbfCTxiBxEGHxh8tt2He1KhVFFKFAta5YES/+Q2MJbJ/3rMyqke9B+tmAT
orrQVpWJ83ZxHHbkPqo4Kcm/lk2THLPaB2uBwI03vpJbB9mf/xTMxg78JIzRmmYupSWP+CfkJNse
z5AeuT1iZB3u54aAUBGh2h+JW86yciYVZ7/jXQAjn5nZ82yEtRIayap3Xq/dWQZdZbCV6hzxcD0Y
eGQS3oGZN9Wze7nsKh5yn683m5jpmWPTNvXAxTMPO6SdlUtICwRKIkqijjsthgkvMjnO0HNbrKEY
zEAp+daSs06mkz1t77v9e7hsx0RNsb5gwWsk6CySQXNB4/QNUndFa7eVCkCGiS/dNbNq3W7yoRgB
2KsQCJxgKynICIYElMlWeS09RbGXV35KjXBRWDRnMEfU5X7TBCXvI7KqvaarFeJ2pBGgIh06yAxq
oVG8WZmxdPOHoj4b2Y6/Cnh3ThuKzZZcgooUonhAZ2/74rdGmoJ+fw87UTFUMCI3XSOXdMubKDWt
PZV2xpkWLX9RL0slt0m/xNlYK7aAUb7CDL+5hMGq9KoClAY9Jqut0YoDV+NGFlBZeWnQZ+RxNA0F
PJ0etTMMygSsasMsJHNPAZQsGvRhV1qavedCkGDDd3V2r7y7tkk5Z1oUko93+WAYrfVaqKedOQ8n
zue55OKiPuWnjyc1dGF3aJGBWPlnlyitxYbW/umL8T4JHYJ38ikPJqJDZvmYlA5us5pb2NSHKdjL
OmXgZLvBkSuum7rGW4UlXGoMEm6yzXOCq33SAjLmBImvoBTZIUQHWVeDENq/Fd53tnLXcT5MgAmm
21P1HWYAjdwRUrknUZ41QSGhwOXrvr+o9lHkAOxiIOixpoAY4xuZMcO5gImboiHvGE47DCvt6BlW
qTHhVV3dOKRMd3ZOILrWe5f1xR4sE3Ndna8CpFrPU4Gu1kdwj6rkVkUmr/7ANK7ri0V54UDL2rhs
iq0UA5FRX2YwX8tKiK5uYBhlncLeWYtm53aHXmoBCyRow53Wx8G/QCd7L7A7IHmBPVKNyKtNXgd6
EvNw9cvv/H3/4Ow2HIMCHjzCf5PebzXyJdcwczUlpdimLGj/Zkj5em+oBmt4GlQjGDSHdw0az8Za
cVCVlhWOMKEMNuOIaF+lmK0gPlsrdIb6R+Fi6aPCgBnNt/4GNb40cWkqrx+MUD6pmQIHi9iJSzsZ
0svye+L2yIwc37+eKc97aY7tNVWq9dyaPyVnuyiF9UhAmqNMkG1CCfz/M7zo1vxBPzbIieQEpjah
rpA21gf8b8xVGI4vGfldFxbGZ6ouASVu1Fb77FZcrq6ExdXUgDzHi1fOauSv4WNVYf3KOw987QDQ
tVw6MtKKvQGTyszkJePBcn8qykGfwBht3slSlYltr/9HaOxIe3bi2U+VNHobwPsSSjnr5VSKy/gW
ZK30BRc5LBjt9uY9/4MpEY/TD8OHZSc/4J0zIC9uNDNRU8u+4LyaespnugWXaFbk8GTbZsefmIc0
PBnHAe7rtAUBA0OlF2yk30E6b9pnyKhkfeBXkjgl0WhQX0RNNLzujbpr+o3NiwNONqQNuJgKAXwb
A7G1PhOlE1zt8iMxwvryDjBHyq1v//EAR95Juc/iltuto4U74X9IRPwv0wju9tEBI9aif/uNMLiI
DphCtgm3OgF7diX5WUYSlTyzz+3Zvpjj3EY47s7sPoWRPMNt8S/I9cN2sBFzU8SceVSb5HsQXQ2r
kZ5n/4CiLdfDXV1h5qZhPZdnPPB7bEqVYF8gk3GaFt39MNsb3I1MRjGyCrbl8TYQmmuaxp8hyEk8
bGwV3a0uJgRO60pVWkePcgvrvkCDhi7UdUxOgDpiGB+EIruuCcShI1xt4vbMZDLrFjnRzh7hcNOw
fokGevM8YT1SFvjIvka5hzatffY780EAKbNXl0Kf3zpiuos+9QJXeY4NmIBstqXi5ecLZuStGHdJ
RoCfZhKAh57dEsdRHulDxEvwRLkosowPAAbkZf6ccu2c+qeZUQDslU1X7hnX7yzd+cBOfjPYG3In
QVT7oPgCNQ+n+xd4c1Duq0m6NabOcxsHNUD/gQNUqOKXFKuIIHogRJ9QRoGkHnMCCsw1nuZKCkmH
Olk3qr4TmE73yXmGfLHf4Ef3kR5HuTjLEQ6bTNGQNgXVBFRCZXmgFb515dASxRYjaxt+utBX4QCn
ssTpjU+PEzYm1B3CN2pR6Bg2sTUHuiQqWAo3zIKLHHUvCCSacrevnw8q2N4nRFoF0n8Gj7GC8Faf
u8LA4tS6iAP63Daqq3Vpj7MTgzsl0MwV1jeVrK2mAq225OuMyTn1X/sPo9kZ+5bhnUx3Evu4sZmN
cvGOiP+0/RoJPC531Ce2tpRLFVaButqeQ/KK23n9E+Go3v+3/wei5VCRAI3UTZ2dE0cuDos3TL6n
NXLr2ghOO+dSjirYhmeBq539kyRAMBnDCuuxGvDO3Fr1rhuqayhIRq6xSq/mkm1naPQn0WhnslFR
Rr/uxcZS9rqm4dGWzVxgphrnZ+Z5trkGEDcv8TixCSuF7U6xroCzMm0+5f7kXwZXCyz8pfzXpyah
H+jSkPbkTstIOLWJyzwzDY2Dk9I1uIX/Ivhu78bNPuFb2Al+m0l0Rh0zB44nEoZ0RqjleFTt0OlT
Q2V7Ifpuq1uoPtGAuBVpaSCOPkZJtbLhmkcz0jvDQMZPm7KP3bfPP/AkkhaECrhdniEazH6XhNbF
yDLPgINuqaPCzLOgg5wyOi/60wkiSNU30fs/lHB9x/xonHyxUEftWzYSjC6WVW/2VDLiQ/qbvmEu
WXUOYjFbGJwZsnf6BMDyhytuvYD2N00RQAJqut7CbYH4Akb+pzK0t4lGrfFKyV1BewAjx/7ElouO
x/zkR7HOu8X15uYTQOfmp2TbOY98MCAyfzMrlKZKsWrZyAsbdS9HcoQXruRQouo93/X5MjZ8Va4Q
m/9q+9cs6avOrhu3ZF/ScQDHMKtWisZqQNUVbq0enmuEu7qxOy+0xHeOAGXGYvsjhcdjZNkMhk1n
LVHYD2B/uIFPhqY1Y8mDMt0G4pKeCtqGPhKi16Y5oK5U16QVi0O6BOSIcg9d0bvpL9z/ngbOzOTs
BoZk1r5jPiOIs2XnA+/72/EhMF6OhGt3wZ2LjUhpbKQjk+mXKq/Qhqlsy/l56y3rJaL87zyUEGVK
i54jo15aY3Aue7NBp3t6esI6YQuwf+2csJfvC71oQAai+RYHnHkl2QnC6XyGgETleXMuUnbgMpwl
qqBjDqVac3shAQofV+lFLJIVWkYybmGbhQAL5hvqU0s7sLTt7QC3GGy/rA/84J7aR34FIW1LXpF3
se+GYopPVe3/HF20kmoqnC903cbVALhkhhs21SD2nbyTnubqL70MoM0999ZKHE3jhGerA3BzlLLv
O89d7q04vD6pLQFnTVAwyZ7/AKZs1pYZwZBmFYTnL0Ev3z+c3NVAkA9wfHo3OVNKILc39xnqrrFG
TQHVCPZ+SoOGMFaAh8K1KkmSm9sINcJlpRwY+PhmPg9KLqK2Kj0FOE8k7GMDmsFqIrPoHPyN1wsU
Gq1kQCYc4JW6qiA7n1QZgm5Pl5rh93+Xf4r0NZ8M8F8t8bLscTNr9vXm3kOK5j9zLQP1jeL+8lgB
NpOFjCE3NZ7UFx5KtK4W4qh3Dnp5dvET6mUUiKJmjzXcmqTzl5nvVAxnMd70+SPa8rI6Sua7+gui
OrCKpEIKne/uho+CXU16YtAYdy/M8HALs38Vq5n554D4KXi6EdBZLCCS7V9W84mRMn49cZEJ6Cgh
bmA//gu8uc9GZVGhSB+h0mtm8XcXdWnKZF/1ffXWigogKs6Zgt2AZanbQOMaMZ1T6ipKhC8OcwX7
MQJGq5j73koIgfpOIXHCLPjQSIUYTmpvgJeiXwaeYG6jp+ggWyC+sppyc+1iw9obMY1mt0yvkJgK
GgxUSd8c7zsxpO07F+GHCb3Mx6z2H4ZyVmEk1k66eFhEbFSHsuFYzAHB1e9BNmkeLL3FkUMIOIQ6
qqkaS0ed+Sjm0hT+IjkqabD0Q4/Ov4vh07pUqpcgTNuDCBQmdcy3F9CT56t/ZHC8jswFDge4MjiO
jmlm2eNzME0503khvu8rWhCEUmHBSk64hrP1F+pJTekJ8CWN+d0FPJPv6gMFwe/nhy/Sc0Ups6Tk
Ix+NNo9tcHvf1etRaOVglxJxoSCAcP9qnM00HXrVQQFr56zCpu2HUp/JDVf6yjMyvTwWxr5fBFod
6vOdNoaJODz9iiYqwljnP1vCYcSIubL0pytuWqsjOam29BZWZ6FvrwW7s/ArgJFjrJLCIav4AcUA
XQ1CeAIeJ7I0aHUI1nlah7g51Vm98EyHz11HyaPtQMkU5mLbJZsjeoKWfGUpDpVnJcfluXPp/JTF
LVTi2Rhu4naem3Nw5V0YrZPYzKg4bpzgBy/5ncS1HCjRnRlbEOe+cDU6iYoK9yxbaGfE3u/bdoWv
oUYQT+MMhroAWYHcKjXgIeOLWz8JJL3Gs/DgF/x8BDhuOVtyKRVYD0D2f+XoPkDqXVXs99MP0mMr
13pyz/YyD9MqpTpegaiD0SM9FYiajSAFmDwL65QpPfn459OW99WROV7gKFYDG4K7SVqiWpEGSpH3
9k5y+RAcvIx52X0c38AvTLbvbO5WiLxTqDv5X4kamcwXDOf7aAxyDzd9ulkQgF9sDD3U77MYmG2+
42SOikhVz4lg7r9EpVKQoiHxqPTffZoa1kqAO4dbfkX8rjRDhlQPB2StX4sEl+zas/Ep3ggkpRi2
GMac1Ph7mrU+8C3bpwCna1JFLDVgxz1OLKtzbf7v2uFAyfsIEZZ2TQs6JsPd6MtEWfb7L6qYrJVk
nRzCQEyKmjG8Untk3y1mlO61cq7FvVt+am4Flc9BHn75XoPdD+OospOENolTUFtZLCS4CMk9jsQb
lhOCo5LsSn0KxwW34fcG118j9/lf0nlI+BWtGooiOImqot6g5WiTODaBQLU4gAG59/LVZ0TqxfDV
YgT7X37FqIAQ0hdfR8/WNLcnxtMy7jI14vXDzZFkXGeZFIbjb8ocvdVF0T/rX7pXfs1Fdq1EEUQi
l0cCw8ISk6gBYCfBzToB3vhsGziPbPsSplx3/d2EfkAM8YLX5MltrLy13SbswAkNBSr0SJe/hSce
WKMPSGTdiDGFHOJETy+GWKX76f2MbIXbbMsZ3XGd8fuv1HbMmwArwUZq7D1jMSWHBjI6sJzAF9iH
4g4hmdTutoWAv5opP+z7T8xsrP+jF/FDNPaZNKzyhwBB+J4A/2r9OHTbEBM+a7K1RwT9Fekrgsfg
eJADCDSBqz3CdTsenGtlUtIKv44Uycv40oy+6O0t8eJkgGRpGiuvwmoJxOhx/zmjF36l9vk7TM0J
DXl7Oi6KM7NzpwNbYN1U7ToVvvMnNV4gnmRYDXoXxOzL/ohhxqw1RYBce+pBzr03LPizw7j7Mj+H
boITqCIlDK/Gi897vNJxOIiNiFaRH67h2EcDVAnFV/7enmvzdQr1w+roEact4jTq/wDZMhE1PWIH
4AOI5kDwyCBb93i0crdWCxJ0vhZn/Vut32qMV31DtV/LgwOfd80Y2c0KfkcWBru0HUCSnJU8vvvT
0soaGgJ/g4TmwNdDYacCuYOl7w367U+0kHDpV38ZS7W3T2hfFanlmEOphWI3lIvGyTtUWpErNyif
0G5yl5+Ck8vsrP9qrt47xFcQYtADKUu8NA8dA8r9LI4k5pSOcdJuQcAhvoaDGhzE0ODMsRQjIcQp
n1bEbH3K4xdU8akW6OynNxU8SmXluXRqvigYiOAcpF/73xX7sEiXvDfIf0gXD0iNUld4CIc2FmRp
NKkrQE3Ga5uSI10nT2iNMIxv6uevXZ4ZTF9ocMYn7fIin3c3tRODfTGL0QvQ57w+F5nxIOM8dPJj
J30VWao1lZbwZ+HWOh7zxfVLaUwhomcXfXUpjPGW/trQ3uj3Xrj2SWMPxA9JVaLXE5dTx6OWFsz/
QRDW6pG0saiED2x5+mBRsHdWRF4+Nn2SwoO+eZVF/Qh9EGjTStui2I6oxefyrrqi35LeGwAl0aVk
uTqMsKLZNuRD0GnjPeJ90stlkIMouL2OtzWPaO/+Sn6QakFsTPfc3v+PYGHU7BzkzxqBMtiHmzMH
aXwbR8fN1kI3oD325olu3SX2u0BQ5V2YRdmLhRJik5kfrrQEBpUQ0604FyLa7NowJEloX2Hk3VS8
cmpZReLk/VARjSopn8I1UZhv8s6bNyhJWv80CH90Nwtw9BSXJDin5OWFILzc/POhmBX14FtCSapo
FpbrHxNPMDHOlYtitIWP2RG1HhDjwS+x5TvLrzIpR0xMIULCjzA6icjEeinWeihXKp6fXaARvFSS
q2GgeUpCQYPHG2DreC8TBeY/8HTjIcIstJt7rcNPfhoW12yHyNB5h/fbP3dfMleod4B59bydpi4+
3gHSkxBrCKiSIyGbvd5L3xheWlxAxzVO1e+KajL9z8xm2z+QGPqL5OGdIAdG78eAxDo6OMmsV/+P
P3FDTc4VTY3vvwle23QmdTM7OD88f8CJ5zH7/CGy7qa7Xp2gKR0Bry/8x6fMFKy4+xDHYP89pPZ1
0KICbZ/b2JmQHub8U8R7WmrnC4HoIKdKnA5J0EH3n13v0uDjGaqLNbUV5FTE6sPilfcwRuLKXgdb
PFZsKyPrH1LvLmxALqXevs7b6brzje8Ni4YZ+aWE8jb4Msh08l3Ek5579RBwzdYwQO55ka2WSvfa
nRYP7IuhYPVKoFAMQLTpy3VtcK6S0dhyFvUe3liv8XOYSqs8uK9Npmk6VBLWQdtgqISWicHeDzcb
am4RxIP/P7TbyFs0FUVec5mER2tyarymhmcME8ZwWNcEx3DN38iyZ1R8B4LQ+aosxuRL89gw5WII
akkyeGmadtI1arubNlq5pL/Bgv9SWH8X6vpIW4qzkotVqoJ4UFJifXo7KFfwj1k0Wt345GlLTxd2
XNaHoy4MofbWY//FvJNi135Klm8URKxqbJAt9l7KAC1nuYIO6Bbb/yx1gG5iXzSBdPcabOWafmw4
QOjils72urvA4G7xUGtuKMohu+YW+3ncwVKE3ufOXygdOYxz9se/W4UVv2MxCnzJo/3rC+leHu+U
YIlr1QeGvHoyga4sW9ajQZdNFn6BQ9/QRur7orFyBEfJ9nCweFVhDRukSAXeusLKnt9ncVOauUMk
OvYkpuoac+ZBRmoGAinkYwU/qCGRxamwyjKMNE0wsBhvDngcJZBEI9NO6i4K0eVkjgKjS714POmC
fX1OdgivSvfmjh3QtPibqt6LuvqjuUAIRvmI9bpxuG6LxYI02Jqh+mJoYO0JEyMzvool3c0keA4E
zIATyAuMZmUVklaSP839x992jjdPMDH6vqkeVB7YBDvMZKhfdnuxxDE4RLRDjbiESxzGUH8rddBk
hSowPvX8otS+XzZg24PJ5mDXl9Ud4kLEnKC3bwBKeu9dKnnua/ZrWBY2xdnHQ6fWOyrsdpn6RiYk
76DhWnSMZYVsfuy4xoRuN3UeAKdH4BX2LPyZ2fiKdGYeWNnjM5INFymv58Q30V7TMB+UcrgqyTeR
HdmQajOBKJRatMRIy+39e+COo9QO1eQenuoxnTVLI/UG8Jl2nIXG8m6GuaW5UsKK2Nh4t4e0l4Cu
Nop8qEtfStlrdPbOveuYtedBSNw5jhF5y0V8lHOWyu07rzGvi3saECBKRbAWlV0tlja3I181UA4g
7eEQDGpNi0Dw5Fa2rRWqcF8diK4/qelhbSjUDxakFo8EdHxcvXPvFSwe+RFVbyEOm6Ie7U2CJasp
pFzSnRTi0S3nzI9Cjo0QQ/SMyxd3u3cp+LDKDTFp91FjfiW5LK4YMQt7h4f1+TnYTydow3hQP2mt
Gq4mX0leb6L/7V5JNnNUod38fXPaI+BE8Nj3+csfBvkLxuJxtOz3+KX36d5qmRnW+HrNHaYbKFTn
4BfTCDEsHd/l5PPMxKmXNvPAXI28CaoYP6L8hXm3P5c0wczQ/jCM9uLiYJHJb9n2mApyWHSejmwd
85Co9S2k+qhJsEq91pq4vkikfEGNs+zVRtx7wUqR1+13uYoJVBdBbO72QMLymud7ZOnx/To9S6LF
ntVwbyGUumsVvlYDgF03pMf9rIyuFTHiHWkHq8uqW8DjaJFn1uQQHNUactzZ/FSCBsZxF1TdkGMu
00CDm2Z4QnC4TWzg6kgnCbjvTTmUDRLkGZ7289NXQaNoX0nPUliiGfLsunLhdAx2QPIQFhiNIWPL
y/ipGIJhZ6yPq++oD/YkR/LO32z7tibNSvVTUuKi3kHpYKllpvozVQxW2Ax0o6ck0t5/b/5GX4+g
h9yjLIXOA7+rIF31s8uvBu1kJwBiY+IgLf2COyevu7goGE0WZnUt088W0CIZpgjGbunL1oIEjbXD
fh/FmmGAv3J/dTa7wZiluIS2r991FHw/2/J1zq6Kvae7lC4vcKk2CssUXQ6v1XkPSc+0IQnd8+zD
kIHIZqas7utBN5TjT/pNJwnbXdR8IJdsXVpfH+m9urbFcwhBxRv7j817bPipzL9S+4ACpxbL3j2u
aBW5I/T06rihakVYgVpkerZDKi5nMSogtoY7idzUUp3vwah7gUKubUjP18xk8YZnrHKNww+yR/am
ziUl0jJ7HG+NhkQrR3sqq/AtdgntxG+7/4j8cYCxyJAfEqVRbhkgDjbRi8QEad+Pua4ZqydmuL40
f7E4UCVd7LRtlzrRYMoNkyvgq+u1ezFJLfp/TW/peUICiV7wiJAU3Ha/1/5E0xcseob1m4HHHLUc
VgNwL8VASzwvStuAg4OoTTgUvOS4FUCyzQgZlTPRvmBhWOGogWeOqhCvYPvWYqaD1l5phEZ8owZh
OSLYTeeIvBM3HKUvzo+BjwUAy2KFIChDNmWcIqP6IwtfvcQWZ/0W4tKY94nCAuimNF504NVoVzNz
142NZ0anKvI1Rl2kLZ3EAv+QANxHyjwEXMabUgfrTKTironz6SDEHJUNjaPmVD3kqZmNuLbs+Iag
wc0nTfxJ4Z1QS2JoGyF2XrYLSep98a58EHBWo4gdwiCWYjWp1p1/zg1mHwvApl+/T/tCwAnmy5hJ
790QeVAno/Lofqj/Ihrs44UXUgD2zeaGxcu6tkPqH7bMSFjRJXvoepk9pLmpUu2JsKRnc1Talu3i
HWPrGi0vVXoLdItwfbuXMTw3D8us1KL8KTlCeItkUkKnLeRRVlegV3A7ntpM41HZMBfiuVFedwJQ
01/o/0jpUehi7Z18ChVyklTNs/nD2zYr1C3BBoxTC3cqR41vRkKmal/w9TdkoO0A66ciUyLMRRN6
fQPUxKvvYQNb1N8HhqQMB6RqNRIprDCdqkhDqbeJb0ke0fWh04ohQE/fTjlh3sUC6gohbcmyigjz
oNkr+oei6EUQhOKDmkko/F1TxHRFz3Ssn5Z6nJ0j2Pzmqd4ibaLvHBQ+I40Tci70nnkjuYiOdo+9
CvE9EVXmMNIdghySqpO6ENH9i2wQRCpax2sMa3qouWHXNjptFV1FczotX11ygySzAp05oWCe0WyL
KUMGOzf/W9bKTcGWHeGDo4kon5uw3EodZYUG2EfQfc2WlZ3hEb4nDO5ilfzyd1buOJRg8I0DwWK8
Rg2F4DQj3wBuFm9foM2X2Di6Ju9DcVz46bJPay43Ju42lrtI6v75j9D9CTQIlpE/rONoy8NpJl2A
odY0oo9bmgawz9NS6jF6/dK1UpMf8T/4AfPRNMM2qEtgoxn2/ysRUBqNl4mJ/A7hhmCC65BDUihq
Sdo4VwKQK6zoam++mvd30w5WAx4FOSXg2j9+KTRxuKXZC+AVjQiV1gTp8qO4/8f4sIazSIYNg50X
tOrY9dgWvvZHxjCnTmiDBlyT6h82xK2hEL6LjRPNdWRDuOa+4+k0o2m1csai2ZOPJVmAwY1QtZ6K
YO2UGtBYNRuLR8ulLsVZ7YWbIDoZyV7SixpHznb8LOgcdO8cYAXz15TnIPaoF5Z2GVRj9luWadXZ
A8AJBEcSdiJWA3Tli+KaDnakYQy64/Rx3K/MBrDhTYa+lXxzNkVlefAtCa3AQlDMBcmdcGMlyvz7
W15Ml6z8lwXqTqAzTf+Ux9VZQSHXTuj0nw3byBDHsOSA72f0Y0sYhTqxnOtTchdBVUEMxX7/zVYX
1CXrBfXuhnyIJIAJJeJQJXbe+XaD2A9h0n80c2IOwu7uNdTTl1Lh3RCH49Pa7gGM8J415uA0BqAx
aY6HjVAP43dOUNR1BGL60QVLD5CXzzKU5II5nctjX1W+d7DOLq7p5fBB+FlMu0ek6/06FD1lK/oB
iGpIapHFdyR59zOpFJzTIZIoY1Sx05MeGTIQcYOJL8NG44CrmvI4Vd4gZQ10f2SmBCJBL6CLJn8A
JoPqT/TAYVZJ8BBjuoLP+qXhjglrAj2WbrhKQ5S3SPwEh3MgxYOYQBUQdt4CkNcZK31bs5uWLQfq
weIjk4bGvS+GP3fRFksFG9lYtOnu6pSYX8XDr1h5fx4OqYmn5eTS+LGmYFnDKvP6yBE1ga+3Xt26
/IRP3cJq7DTDeunnX+7oPdpqxWRKld24ja9dbDy6bf3XUECDQitghk/jFBxRuqfGOhiF173l/O3R
07WFd+4fWumoLsF0A2BSbXTaaQuwlKPGuPOvTKD0BBnQVpV0vLVru8Irm5fg24J4V6dGimKgwaUu
6uLwPH/7TqDZ8syPMtusjlryE+8ryr7blHZiSavp2cdpohNoZXmqHIXtHi2W3fVCjqfHqQcCHgaW
4kRDzWjlEOdMlVIvQ9hvhL3/e303P/lwaK6hF+oPyI1qnnSDz3D72yXped2NdR0wF1Lij7Ym3TBH
FHkUeGA/B3MhOoWQ8HhmR9bf/Qh6RKK7jBrGJGFjmhT2v5phQuX0HrrCvRT7crJn+sWzq6UJuBkN
M5bfjxdQe+EMRWC7f/mutNYwyEk0PfskhumEHk4GRLzZeh24ebwmujW9PvAnOHB9OnWMiHC55I5h
lfNmhEekM+nq3WGONfEUT1aGTS1Axma8FwCZHI3v42cyLBxZCSr1p+3YIxyus8Ha5kGBkzJemQfO
PnBjFPismVsaoCir25v+Sl9LUjaNOI3Gh8+NBgZQKjM49AkL6ouQpMSaumeHHnLnpvZsxPfZiPRA
z4u4rJP78BkgAG2B5CvhtIVt7/s/BooDedouS303dFadWOrdpN5REzuV5hO6UXnCdVziZWOHyYT4
Lt+9D8WmRh7CelZ05RujelFYGuw4TEpXdcZzVE2cM6EWwQK06vc+GNG50MNxZaCq00HRxq+H+2rY
K4AjtAm2mm69cubheqhybQTuxNz5AuiujvTtMNbq+stkcz4g5QJ9vtsf/7Qhlvgm+Vg3zBVyMw/b
QgnJAJUDsWrDAskrre1BQiPldGcEnWC1SPlcqR0lTN/HNIUAr8NDIXQ67kotjmuVBt5t5XfQHWj/
2DjybDWg7hbAiuIh0uuGxr/XKqS3wNVkROqw1hIuL8glmapTdmAoZt070ePqzgpeXTTJLLTAhUws
X5N/r+Qulp3uXtDPk42E5zj++pWOshtsRQK7vYP9aSTVIHFUOYQb9LsIULEiG+KNEbBm7PxuwGMb
77yrw/Ih3Us6LZZ4SrU7svj62J+zrOKlYJfllSbcNFTASeMXBdRHKPAZC/tHM+5Qy3KJjCftx634
6fVOfdnsCKo771zI60sTF+PDf25UEPYTLfPnPLp1TG6Iq/msMw3KuTU5np+Vo+FKX7oAin0ty8la
HISVmC6LShYbKqfudbyeUxiYejogX7AUHw91GQx6kypc27lIHX0WBfJcaaBFpfwUgu6euez12UM/
NSVp5rAiqzifdSTjyzH0KfQNcqH50gpORlnS+lxuyvSF0kVVlmFtM2VicuY67m70Ei8/Vcj6D9zQ
IUKB+3BHvY5O30RSPUfSHPpXp7cka1imZNKRSVIEvGXehISmqDw1C/Y7tUrO2A5gdodyLR+5esNT
PUkReT5mueFXE3HUkgfYQmn6kWhXrejbLieAkXN3KaYZ4uYhdO1QTIk3JBx/o1u8mj9iMAexjeAd
HBbFV/czhqFFG4XEw4hZKYbR4w9Tl8NKL3z0Hwepje8+Db35hCnsTmbNWMGOZnx4PxDkTgmm4BB6
eZaLRxyh5DH2nJxYi2Z1PPnD662fFEALj8w6Tmp/RykFQIC0xGnZiz67+0QYvP3bEWNKxdbEJDN8
qr2WVDXPM9fy+EJUuAzWWsg7Wg0gTIC9BtZkEvFZKQi21/y9Inz3dLER+3NuWDIiCrM5iPZiklbm
DhIrYhM+OPnDm5AmSja55ksyx9yz7JWtr7GwSpmTNubWdTRRR5JBl83NjNod9bMHquwq5vCfX/rF
cWyRZXWzyub9k/jYn4HY/sBvV++fXNMp74zNLCq29KCKWDjAMWhKbtObHghKGJxu01FIPvhbxbs0
OSewhy6VxIGL8u9/LPCz3uz7KihZHBrZ0b01ORmDiIEsEL+pRUHXvCBo9eJrJtzHIe42A7AqXEHu
E6HYs2IgFG9A99wjvOd259vux0mQ8gHePSw0cSqa9tzVb0vOG3g/uSx8X/Cr+nWilwhoygrr0lNA
uj6PFJqrOz51hlDvdszmz8KDnRbQy+FhV7VMDMYzAXwv09ltI6ZvcSyrp2Q3MUbsFt/QPsQ3+DlB
Z2+IigYlqGUZakzC8nnmc3Q+oakCZAZwDYSNlODQLdxVCmtWRAfkxB8wF2K6E+XDfAYBMyjkkEG8
iOVx13x+jMxIFVvgSCSX/zN73hiKfVRpUhM++tDfXKfv082vE2spCSNpMIaIm3hsJB1RM0qxHEQ5
L5JmsYEr3tsoM19rnCslvjJQbPpXjOQt86ZTqGEWl3HY3WHicVW2mUd8qaH8Wfr1a8fyuH8hsYMF
nVfvzTptaGjfrSEF3Fae6NCJDl13xKN8F34X55HL4kMEOYONVdhbcmDOV2mQThdX3tt5IaCO6j1I
uV+EsWvEBbEvnqebamuzxCSsK6sD4H2VYUOlL6mDSyYcHXTUoF03w+X7nNEiL3b7EC8ehDSb3nDZ
57IE/V7Vv4jOK8JSJQHdys3vMaeOpzzY/sjPN9lJTGxwK1d6m/xRAC5mmUBXfW+PDiINti3bwmF8
uARc0l1V/CPiWaKljEA2OfqgvA5QVvgNAtJgqHEzlK2GIHcAI42tZFlVjCSXb1hSzYh7ZaYaQAzs
OLxC5Brt33ehmfDpXGN9sJ2O11AM7FYKdCleeUYyLeLVbHZXbB6cMlk88/U39QYhOM6d+U8HCyns
uskHkyhHwjpCHhrKlwBi6+EUUfPBAV6WDFLyO/Qde1nKV0YpuXUKzvP6exho1oFmlYj6lC79+Gbh
fDxpfZDwlA/uLrIgc9U4oe77EAKQ/Pxb+AFVw8HiPxQ9JyC9UPY+LUU71gn6F/BQhEJ+Dh1fYDPs
E6L2joEzgXJKJ7Hc+FXhoRmpgk4UTbSfFpY5X6oDEJMM5k4YuZ9sFCehJnihn0c8Q2nEPAULUg6L
fzevpYOIFLG5DdQxpIpdUQf3wCw7zjLDxmxJ+xVEcJeGvWR+8a4YVGialKJ+nGkHJrAaf7kADIKj
ThPriwTUsC5IwJcjgHN4C2Q1syKdjmACcN8FQ9BqepskuqrVJYqI7i35Zmd/J7rz1Qd+IFVGbHYI
4Ytg05fita7ZwUStfl8qv/h0eXIdfmelB1HUgQ1zK439P/zZv4l/3vkm2fUjYU6KlMFTQhBktkb6
KM+BzdgO23WQJRc4amzgjLw/1d1WF39ulKCUfo41PIyonnPwhtWRCaTb8yoXc1o0mjAVKgNo1Y5I
FmXn+XgwP/9Gt1/hTHTF8sdnXG7y0vs36CM4Tdz2XVbCCLOR25DfvQ8U8czJ/HExTOmgdlohoN3t
UE/itr1EQwnOURUHem4OonKq/Y9wZpsRBvSdhcBFI6yztJCekwrjrRfR/hCtP4uHbcUWS/SjGFEB
eajhZfdz/Yx6MtA3Qbbhe7Cq4J4v8pKwwikfEU0xKcwm9qTatxkwr2f8wKJl+5RnfPThJzALF9FG
/MITNjGROXpeCS4rfyJYLhh5fLf8efZo8fJh4UjNO41/gQRGogBOdc4Mcwajr9GcEJMr0gvociIF
Lhz2I41tyhEj15gfEWm+/ivrOtWj5B4jp2b049FV9pIedsc/qq3Od5+0FosNZS3vAT+3Co0YtRlc
r/S8JxTV/y3WlkZ5ZMSyLqSj6/IJQW721OCnupzJfwg4BhyfQTyQEVx3DjOMlQixcLgoo7Tt1SMf
dqkoX693z/IU4fEY746j0wDm/3NTI7/0bu49EkWj0ds169V672ku1rx3FvzeTQdB67l8ERIC7uJE
QP/jkl6+MoVLikN5N+DlX8BJHHpYdx/zMmMgfh2RUXbTW+Unc8MdH8KKk2VLSQrYUAoK1V2R/DRv
zTzs7ei22JY0UOrsUg2Et/jOpPxzXlR8KnJy5qCFgU4/74JMiSg/CymI1ybmIo0tgKXpzhqJ5fVh
1U70HJU7iVEMllqwINbolEexm1V1Q8bQ9ZMg6flWuf05g6z+ghxEGyq+qKm4b3CvvIQ92JzLAFhq
G18QGU97u9Js8O/DJ2AHJh2qDTTpmOr5dM/7z0+QZYW578+ML5YsuEyN7AziYKB3Qyi+LVKPX9SW
6epm7DYZw0T59HgJBQ5V228Lf0yWdAjHboCHdu35FPE5km0Ini6yrhIzg4yssnrizxdZ/rW403OT
EDvYI5o1e/E7WF8eL6PtEA6W8ffweJ4p4EsuXjw2vU3UtXMejg+p2NubBdKZOu2niR5AWJ8o/nr8
kJlG42AOCgTJORoyisXE2SkybSkk4USSNYkS3uC2ERYhE83X1arXRQycw+dUr9o/HUiwb/KMBzBR
MrPGm9u7zdEPwMKQjRvXRiqb4ZiA9d/TOa4u9mgttGLdYUxBJ90UOqK7vGT42XFbvw8XsoIiZTmW
rhl8rCB7Hxu+hK8HW56p+MjxHDK1AfOgRyqiZqgV2CVfOfaGu3YpG/KHeETOFNoBJTqmZMSoLLef
8W1IcerUfKTIf7w94SL4CtQklctrEABPt0KBH4cuRKajRTY2KY62HsFiUuhvqpzYdstLZjzArjLc
B6Gan0aRvC1iGwY3oPtU0ZfDJl2/via6iuUO5I9eZie962Y8O4K7Xhx+V7CXZqlW73GYt0UySbj2
yaguMB4jYsT3vzmhNJ0rnSYZ9ZYlWcEzngHuz9h7Zr1sNXM+xCk3el+P8hKAGr8LMqjc+r/WM46d
xw6kP5Wx9Wz7vWac8WihaqhjHanZriSREnZmR0JGU7Czh6BPvtcSMx+VBXT63ovZ0EaEv8pOoCay
oY23F+EtPAgBYA9OrdJCK1slbxSApxCo5W4TnQEM6S3WRmhH8lznIlI1L9tl3Tn8YtWSfDIoW0K6
WjKt6P75Y9vwLQLxftbnKogm7EmBFflwFitJ9cwNowyPegYZZ/SOcbeZxO23pmW7U9V8aYQpsi+3
vR1jhIcTsZ/g6v7uIoQg8XpquS5RQcu6CC8GFcvTyTI48Ieq6iI6DRMcPYQ0RZqzrxjd+pLf+xVV
4aU3Tvy9itFostmE77qxZWY+Sd+9yICAB6SzT/xqM/m6pyYM6unk0dLrLVaWLBfnmZmy5RIrQXQA
DYz1/f5WkAUlqOZvYrlFyuahguNtVL43lUosN29DN/bOWPX0TfIHVdFJhsMIYNomcog1KQ6dC/FG
gm8Ux5O/RGVZgAIrKQ/+4c8qYwrmsD6pjnaT91ZfpysSfp0zM3S/k3kLO5y/EpRisQ+OIwC+dbWt
QIjyt+mWtJWML9oi7oyb2mZTgW3eACsNgBsfP+fnEnavqbH9fYevFHFUmyuqk7PbHOcGWKbaXMeD
PZEMoBJz9fEB+nhWLMqncEf1wD1q/MME1ogX2XID0Ib0czsMBDe0GVK/cyzVmNUvC5K6T9/S1eWV
JolGkmRdHAULjO7fIykaAXhD+gn2lVpYqPQt0rPcuLCZZZy0+RqJ72R9QD5h2XQ2I/ZSLGYhp2hD
hvoervrHG3K96nif611sEqGsNxYswQ9VqQAn0kTLJdceqdnMLF5w5GBpR+EwS6QL94/N/NHbO4iZ
bijr/AdYjHBuGNrf3Rml5d8wN+GxY3+cJrpqPnVzleY+k7zhYfVP4NPLPX9XycgqzuWkbB1Y0ENY
+W503AsbD3vxpkYzN/nZK/iHGHfMnYAvgmqCwfelkCS6wSQ5+OC8LYfnLCOYo5whw4IcKozKRFkC
oilv+bzwmp2U5khY7RH9T6tkL8GpxuAtRSo7eTm5RdZ1mTZ6hPBzpK6LxcfigG4XA0ooaoYDARSC
OzBw/qzfV/FmPxaAz2znV9Leafi6+mfa36SUsSUV7tjEhgQSnpujzg8zo0ls4Yxx4WRUz6Z8PJ0Z
Hc4ILc3xgf/UtgtID8LvxrqQ03jsWRDfKYRN5TwG6iXiguSb1nK3uWUvFZTc+ONAX8rGy/jVT7B2
J36qxSUVkQjvUVJMw5K90HsSB38JBU6Otmcsdei00pmAlui09Y/G+dXSHHs1xO92xJ/oO3BaZlX6
DvRHknXL5INXDSv//5UPDoGBgQtbJM+u8VR9jzsLvb8c2IEuggNNbndzqUfIgIicoWUDUKaqvqtG
8xpe/7nV0hU4PZYVUM8VfuENEwk2QRaC0F7HEcY8a38SA3xG0iDMA8CwNaNul6abmRvU918p/I6P
nXTFaLuFWRK/RIP6z1fdhlQvUGFOO5nHiOJw3eNq6VlAe0Pn5KdqcfTZJ2C58iTju25U42JT67S3
JONNskY2nMefHWLw2h5xcd+j3xClAyl6UWqj/WU/ocivx2uFj8Dm+RiQwtwwD/zk4miN5wIzoiBN
nfDKDyABCtLgKImRiNFeHXog/TCxzMLDkR4HTjdYFcc4++UxBJIYGFuqkzi5Be4JxpYQ3Xs/Z9U4
tA+51XXvM/1lH9/2toyigShtISzEAIpXeQOv6b7ETohSaU8NiorOb2yy0zZQaRT9WrQBImm4fTGK
ZZyX4/KGliDfJdNWPuXz75fzFhO7+dHljm5qr/UgpNxO2A9vMP3XlwAqJDYWpKwn46sIAB+MgH+J
zqLmONAIyKTkeugUNXpH+n3mHJR4xFfsVvIqJeRrhLVizWSUf9zuBUC7k83K3R69s+GlZWkfspdo
9/EMi/NnK+CCIKBxZr9Hrr9x0D/o35GHuejKZF1LQTAgTJYfSVSkAtaSM51ItMsgCKMHs6hIta88
x1qQP3PvE0YgjvS6pVuEZI+ICV8UI7MBcnhukq6TiaSy2/E5J/FLdSe1wy9NGn8phT7wj/neVq0L
BnYYxqV9SWfCIgguebFT91ocnVxfTIOcnyplg6MXGFSn7Ur7yTr5/ZmNgKZISw+vQye83GDzKWAc
CfhV1Rd4UlfMsMd2cvbl4+nIHhC6K82+er4vUPOn9sIq7zOdOKs3MZcZa8IcB7njK6B1DGEnJbvK
qJOvBQCozi16igdGL80fn6aRoEjOcpE8EmsyTA8E5gx5n1Y+8ezCfohXt0+nPOKRRFXISbfk3h/L
KkK9t8Eq/fvSC37th2tUDVzFlvP9rIn1CaxY314EAEn4+nFo7UbjXNnynC2RydouvBQcpwNz+2wm
31hlZKdBju8+Uum5Uw9/hwrCMEfdPA7LyCwtRqiEpjZaC7BowC1pnx6vWX+PRETZGIQj0kEdSnIc
E5NUucbt0XuXLJlccjLUSo6nN7sOjZaE2ktBbcqbZsllW7xrJ9NHFrZJ5NKeTe4vKefMnf0lgfJJ
lj6siXUEDVzXJKSskiTDwk0C2WgDqVHRVUlzlDZNO2NRVsDWT4OS2jz6aOTdKUUqsEagyzZZRO3B
Ayw6OsFfMOP0C4JCYK8EDcN9FZJG7dzkqtXrwHcu8XiSblrxYEbwEc50pMCucLZf+0OcuIb+rJFM
kG8qrHMqFSPlBmsqin9mFj9NvT+MriCS6LiTtlVQ9Ec1h3gqGEyvenKm4yL7qme0Wmm5xGmHulyZ
dUM7phoJgSpdVpgb97/XwN3sv2sw+P6Yg6EcUprN9EygyxmDTEXcH++oepXkXJtokEtwegOvmyno
vIHWg/Sg3607aWGwkFyRqgjp8wTJOT0mwn4ruK5AwCPcnAL7/h8UK8ISUaaLaebgzr2ZxP5h8LgP
ag3f/DuHYanqDOsYBEBerauCe4e13xaalF4C1274mrvjv+t7Eh5t0zIpbYr0q0HZdKZvKu/3Uxag
bIuxkPf7sJSBvPHYOUOm5Prg+KEnsXN4EmJq04km/7KlAI9bdEalRfDKmZhAaVlG2sF050a7NNcV
+5kocR8iYjHdw1IwKuy2jeeqgruLZ2T+s5K6clKC+xJrTjqCPFLqvckFWVDHq5YuZs2AWeWi/5r8
Hh3L4W3mMFe92/NzFx+/4f/q6/ERAyedJFeS1VbwnJJ9aRuO3EGFXTQ9/GCa4PjJMccBbm9Cb6/3
h84AMpDkptTM7f1PbBLwfaRYXQE30rTKX2u5fgPjWI4Jc/aQPc0/wn7EHXePZ/Fq3pMc2PJxaeXs
WWAzTgvZ3Xt/TfRNGFJTmm6Zs8tZY/SZAcZ2u0dd1YS9JNwTYggSJa+4YfXD/CligMtV0CCIbonr
V1wzNxv9w1grgKMqDFavEmdsPLARpRQyJIOxogTGcGRj50Xpoo7u6sxPoxA5NmTYf9gcztfcuQm4
YkZGkOXVorfkeUy7eJQIPu9E8bcFNsycSgje/uI+JrUeT6uKtAMB15BVtR4ORSn0CHGZIo+Q9gKy
gkFpjq6DUDuPurnBg9oOlzCqHLjj8XvZmUh8OVNgRhap6MkybBZzQCT2aQVnapN3GtZf46qpBCsu
4E62FSWHXWH26eXPTt/sUjs/aT7WHRRTLMARpAS21jnmYTx15Qk2XCPqe42vzpU6f0Pe7sSGoRdq
akIHDrCEHY3H06OvSh+cCE2UeQCwxsaoCKaCgY83x3ni/fCoUnZm781aVg5cnz9LIcwE2ecDXsx/
HEmgNIfz0Thi1Aohsg/xMhYrvBjxXWwzJTaav/JWRL0eUKvohIiYefLqUPRQAGu1FhCWQyA7QYtQ
/XMsM7TET/kjgW2kI9PMA5CvZzW5VGpKYY4eP+PwtwaTayaA+P9h5lIUu2lgi8jXShkthIXxcgwr
Yirguu/xnhUFBFQPDdY5Sw1WfLYANXACro0wZ9gVAcwkB5ete/4LyWoKW7C4yrd/o5OVlK2hT6Mf
tVmE7HrsiTjmaaXPElwceaTLmsWZbZoh31HaDnBqBwDgW/nzz7BE+kwUIcA+aW6s/ARKZHrGLDp/
Pee15tclP2I41kJXW5UG+lMsedUhZBkNsdzsztv0ujpRD6+ClT+0s+D7y+Im8AUqobJT8vfWPTFb
IsKPuQE0AOp9dA45rd9VeBwPGQ3kV+sSxnJbJ0JU2F5JOWzx5X/whCeSgvuXbBmfQBCbzYU6h7G2
nOZu2w8PjDIfv0W4WR2qhxpTbSnCZv4BCweyVRh6TL/tMTMCvI8Q0rijBODGyplTzHIJ5Sh7uRfs
bQZjZ1vv5ikUbyO+0W07z6ewhjV9R5qil0ZlHZEdRtwkCmHoZeuimnYAUpGl12frhQRmMpJaGGKL
Q7DO+ufzrGhGEc132zj5POUtf8MKz8Xol+C4qnPlWS9y+2/4IlpiDokV/YLz1uwr2KhA6Mu3Xwrg
S3a9C9N8Me0IH1NJZtMPTBH+S8tmYMAiMAlL/djR+m6v++1KuCKH+HI7yeFGK/uDy8sXkPuKHogl
HxqI5i3+UNVqt9ob3BP6bSmMNym7Eez7yn+YcHA7XYpMVEXXky6ceZlZnr9EGVsvjbHAphL+ZCvl
WJIEV0G4f6hZlQVhRAZgeMLYK9MfTUI5Hc4Al00+VseujPQzUlBjK+zW7IECD/mOMq6ntbikNtmm
UIlfncoG07/KvftGFmVAGnaRxxK+GI4Far6LL1mtCb1iXI93pr7tMh7Zaq4n9+HPhjl/Xj6HhSvB
5pLf9ExkFA24J2NOmWS4T1hPQ2+o/74HIxi8F0J2Qr6xtuHLmwx4SpBLxgPZlIBH5AqV4NvVWqkB
M6JTiXLwjXBKogo8rx8Wv9M/A13N60jIkYB/HJOn2EtbUNr0MQ1N9e+0JIZAIG4TrfLKgre1dEkK
atM3oij6iFbY/Ib7dCEUx9t7m6ASX9lsBHSRQLtq683eGp7aSu3WAAlDGwePGHPeUwK4iBzJOqRR
HZj4GzXiGg/QRhV++96tig6TktEtQRq5vtwVJzAZ+seh2DVk9dt9PH5MC6q5AeeQv9FR8O8pSg/z
b63sQwD4F/zZhDYd2WK+btBbAUq0zKk4dG3qZW3+niVWAYxPgHYLaDLgYo4/4KBzjdljjGI+OWY0
m34m6qOJudsHG6yjZgNnrMTlQ1MlZiD5D0wndHdNRF6KuTo22ruYyU0Ze/rU6j0oJpsATz+hxYDH
/nkUxxeWBsMO1SyjVNEG8+u5r56YXZxmvlwzQvg39sHp8OwuFa9V7jmpipdKDGWdH/N3Dv3FdiAl
WVAugT8IlRdgFV671zUEZGYkCmAAs/xqj3Dr5kkToG2NUDi/Y1o9Gxc+nd3yAvHflFS44OE+b3L7
ltPI//hkVddI1H8+0CPZ8o5YGyNhHykMEZXZTG+FOARSETfjpuVE0TSCaxtqH29PXbwVETAFpmAb
XzZ4yiXCKWV4tqDdk5ZFeN6gDlbQZbe4DsSkCX6TOTsJ4oPRP2cD7Q10uBfrp8YnbTURvR5+EuNF
VXFNBB08uEHT46j/0HqzpQ+BR2R23dXfLOZ+GYJ2GIaOF2DzdGkZA/auFu41pkK1P8wqn0F2xIN/
QpCCPJyTs9qtApaRVLkMBs8eB5brxYHXaNixaKoW1iZdMW0Nu+NyFEGlE/TUPi1p9Uumwg/D9Wdc
xpFkSqFdxnx4YdEVrOF5Mqt/eCKqAHYxBnU56a2LfRR5+o8Ve8UlUbuaJYOEUxiOHk2IlJg1Y2fg
yVU9roJOvbhyHLinahgy3HrG7uX4J7W3mAxvxSYgjKYp3T3xe9/H7Y8efbDYr0A9Ge5qEiiw4pZS
oFGhoAcDQlgtq0llXv1hxWOu2wrIEijgYor8lQPNOKyTfkjOmgT/7XdUru0UyYGiCD2uz2WKF6BR
StXQ7KFl0iWO21p2X/B17afw+FRcrrR+2vRc+FI7jSPwsh561ibT8pyZ8s+FUeId/Zfdd91KXurb
k/5bNo4xuyrteQf42yd//tNf2cfskG70C+j+m9yRkkvBXdHDOiH/tpjgns23sjbVAkdv+XHUmmQm
IJ8mKu7OzJf37JkCKgwc9wWn+1TSCSkcfniTzRfKqFmTLANU+mH8AKhck0ivRspUMQyB5APasA+J
2Vx9urKfjwJwTKtpB8dSIsSTVtXBT4A3sVEQvX2dC7R+ig+mkNOqm4EgKTaR593VSUJAqJ+FWqjr
9stfwQ/40Mp2WGeQwahrnfpLlG1R/pVOXOxIIYFndv/lD/B5xEh1JJPWlGgNsemawM4i++Qbl6+u
xeB5Uc4Dre9jhkp7wXQuELfpUMz1huRZ4I2q3BAEtTuT+MASvWykWW5LyWQ1EkPbqrrlBJKsl8gO
rm4/zCtJShwuVwlnmYi7u755VIWI73VsnZB66ul7RYcQKMEKcbOUCyJLa0NaZ6sICctpfSHTxw3Z
jjOgOdkwWB1tlm5NCcYensOtf66mAXUSl5cpglrzsh4JdE5pBJq9GmtXA/nbw96e/FPJKwwskuhv
PZDQUxs6wysF+OV7uW2wjFU/c7P+wo/XsnqmAitexY1CO4xmkgN5QHDquzMXX7LoZjj4D6ahnqeN
gLzAxUjHTyoJ9dM6ux4B56VbTp+xtEX1zOtU2bfWXgP25QoIfEENMXB/X75ypQpNosi3td2NX8E2
Q17VQvKWttJAc6AFdHT9raHrfA+tsrI1BP6opczpFFtjoTNYOr18UOdesmspUhw3u9ser5koKdbY
e+kH/9tEQbmKrDx33p/OALl1x9pNCwnE9KmIOD6goA/BmlD2IIBcvoe1M8pFO7BGdsxU3lmepP5/
d8qSN9OriWahGQc398E18Oxl8WgUYSmtIimscm9fR/G2lcXXkODoCogJBLYsRTgHpN6+vUQk68yS
YQSCZBunQMf3ke91l9ovQFaTPzcjqbATx+9Ok+INwURv5X7sdVJe70QuvJb3ysTcN9JYYi+jsX0C
PUjoivJIayHYYOoqsxnCUxF4YTvzAaWOl1E83gaBgEIZ7Q071N1kg9C2QgRTybJo199XFLpLFKBM
hVErGw/TsSo9ich81GkdR2964Hvyr6DsD3a0YT6YDrVmJ5hHhgaM+VgUPlQjCySmY9lU23GtQVvC
LGVPNGMLAxQtD9/9Xq0I92zLsPb58QcSkQNoUjJzO4EsjTPLLmuYgHVyeCihd3JNK6nj/ucK9Jls
MO9k+TzEmTDhMiQpwDg6CCqx0FVp5tUg7jBv6GTSwfMzW/gzP2wPvExatDqKE9QC1Z2yJueYcxrE
cb1ugTRVXBNKN5Md/mB66HEQ4gte6BatZhseS/YW/Ud7c2r4NJ1+hbh2YQ6lvylbNggOFnt6CFfo
n6xnLupVzJrULBXcIKUepvRflIHiShfJP+ZyLAZdthrQlXnwQGD37vmlu68SAjc2lfKldx6hkvks
5ZPWlO9XYehn4CBOx+YQPLsNBgP0xoq/IoDtN5LReJ18V4XODueKLN91nTx01ODlJoJqP7++P+8B
/3O1lQ4qkFyAJmwq0jl4wOxtSRCCKysz5CODBq9byGvsQTnh34aqIimMxMhUgLn+L7Q3jrmigjez
T3lphNKtWQtbFIpJWURcNnSYdREb0lZspgndjhmVbCb1nY36AvhIldgOamO1OPrVIuoXl1smJorY
kWlRiaCll0tzlkmzsaEwnb8zV5v7CAZW1bBdJ0QT1Zk62bmpExz0FRV8KYNe3qxz4iKUhFB0jkPa
GRz4Ox1PHOy8dd7Bk5/W9Lattu//OTV755E0kMfV6V8q3ybCSfjNWD7RNfQ99Pch5V1oCMDNnloq
JcRRFb1MSYMb0OEG5rZmban/zGmjsw2fn2nu5ZHr2Nlqw+aOdUaZ/kNeB6ChytHQHsZ7fuWG/pF1
kPG1lkLjknYi3vY5nJW1aiyy95fZDN6bQF8dx/HNRNqkQ7m9ZXdVYQzmU4ses8b5yMHhLHvo3JCz
gJ2COU+K7nm9BsM2DVkZw6J8xiwJr76xYlEs12zyQAFzwyQXBWNkQuDR6IWny0nUqbKx2GjcoGer
poaQc1GMC+Kjxo/IAf+9Bj/0gj078hDb/45yQ+cV5YvGNq4RvdmDP2Y+YlsHN6b7Qy6s/ECA/CWR
zSE1wC/8mHUU1a1NtHjNOP9QG9oY+OzmF8xSk9rD4WzlZrNqua5RavfZ96MxD8GJ+GnmiwtZPzjx
5gcinwaSmEyF4alVUU/Su5SFtSDbWqF9EKRRzw5DOhbkbl4b7VGU+bhdogvCNaKCarTJ9gg6+cWV
vkZuM3hRqD+oaDHrIzhVvi3KUuweU7FGT1j5Y7zxaPz38KQYTdX9OCj7xY3ePlT+fJ9ob03AKXk3
iSluYsViY0hh3FpMpZKpey8xMoCXItw8gn6azPjQNolyqIrbZFRn8MU+07AD4XXHUXplAPv8uxdK
vczdnJYvT0ajlmTfO28XZUtUREiLVlW61q4Ydd5vRKnWIctsESpSUPc6y6A2v55FMWTlFav0Onig
rGUD5fp+P3x5UuKMxHk6FlCtOb2yFD2h9tUayrDY1lR9PFxHpEAtYjcZt0YPB5AXzGIV6rFO1epX
rH2OdWeFfTditSu4xJ16YKpElTQGZO51Lu3sqLAfdYzEW43CUvObniUIxB8ykKvnXvaNCS9tuztE
zdPX1gn4XAva3tn2W0/CJae4lmAxNBOsz4LiSeODOTPks24fTLKe8MsVHU6IztIut1Y/t3qJjpOi
CtinDir7jvw7KxNbS6q0gTo478G1NrfY0aPbEajQj7/PGDWBCod+cI6/oDn+1jITLoMyb4k6GDQV
HQwk06yV0Cs8octnS3i4dSimgQXj6idgOGEXcL+V55/6c9NNsOZ8zXRc9dCvuZLygICll3QDUUDp
MyR4NHKJgzB7yfLlXKwOvM0uTL7dkPjfgQnp5nznyYjC+JthKOPto07guRSdTyYF41mdJvj6NZqB
I7ocEpxDsLN1jG501ebTChkpK2kPPZU9YuA9Hn64iXxBVVIRrBYelCA+Ay7DdoWSVJoumfAqLy7w
AeCvaHqtadJ2showR7Qft1M85A+E5xHUiogimBQv8sE0pvXQPrU2yBwCf58OOp2EpkEsjgGQSO8o
t5u2l+2zCImiEkZe0SKwd6RWMG2nO2l1c/U2ZKIqkqzXWXwWkAR61XDasRXWs1TPuzeM3R3l1s38
ST7M3fJ//5QMjtAL/1qESaB27Qa9nuAqrDN4tmnknq19TKocJt/e4SO9HOipwqmJilWBhHlexNaZ
2eTy4/H5kIkpKaTBdPHS/5+yGI+3hmkzOFpMbkYYxyJPM2t+zqXC2ik2GhQ5fcMVZXAgsKPPQFX5
dnjgXZ4EPAn1xi0qXQtvxLSlA9jFMRXjXg2iu7s/f0ker+BEj8H4rP5/ujBRDvZpQ//2MJeB86DT
hChFMi1rUhGOJ296dZJv7XT/VlLFYxRTnFp6qQg+sx2u4z8IUep6BA0GCcxdfJFTB/yhrWEMxj8r
gCbEVMip+HfUwm/4ud11YdFotS7gwTY0L4ssmU3qMvgGRfjrg/1Gi3cWtS9aZMPv5CPd/TvE2N+O
sH4VtW+KfWkWUK7iVv305j9cCFxrL82kBjZzxd25N8FKeBUGXBxIxa6UerKawnBnht+/L13hERC9
CFsmc5dO7k3+O16I83Wt/f5aTZeyG3xh8p+sGxZciALvMx3RUPU/atmgbfSaLexYvaEePCUeBw0W
uDvzQ1UqoBpmLDuAjIzgSwBIVyBIUECy9uTgVo2LgIZeAZKiz2bRFvo7W3fziO4cbfwOtzbumjJI
H1RLppKSXTPXbRHvhN1zM5IaMi1dGZCKDHQd1EWElTgupu6XPypvNu5GbWJNeqoRZmKHGaPRzqov
vnOPYMy/n1keR4BWRfeFl0BXIqoqiLzcmKF/Cqiz959o3XxU7jtbkPyhyOP37M1LUWPNdYf2BTQv
FxtcDrAaUc3eEalAQrqgN72LKvk3o8QpuJK0FseIoM8tj1o3uO9xoBqbkszlZiI/q/lNGFkhR2YX
1ZGvp0wUZoA46pX4LMH4Rj/kJEGv/PGdekkxLPPIOe6cB+HoQbSD59spe9+7Bbu/P1GSs2ot0kmp
VxTkcWZlIQAD99QOOdBkSjzRm7EP8teXpFo9ytDDuJ+F1fH8RCLKiKNEygiobdRI0qMbnPXDK0OM
zdPbjIyvXJhpw82bL8OSEenottGRuNTPGIkCJiZrnYfYy/xJK5Gh0aZKRkFklO7XIOuctZTqc4YF
NvZ/zZSAuX7fVV8+MzxL1pRqboREyFovmpYdrfIR7MnLxzEgi9KHE0XZMc5/lvv7y0uwlY1ndN35
p7riqGjkLPUJvx0BWWlTrbEP0UBhDVdDuWNeAyk3+C3zuxV/dPzFlVcqzxE1vz4JMSyozdIWjK0p
NBkvvQyd3YR9wmGAUeOFvDIHnvNS5hEiy1ZrqDSnRwpUy5GQAn33O4T3jTDLn20NThZ77NoG5HLP
MzIKRzN+jPQU62DU5qE2Z/j4C2Mx8DsBNq3aQ3i4C6ZauJLgvNhAKESFSxZ06iblaCXyKL4pxfHA
Hg7s2HNoXkCkDlbOVkoa5S2CbNCclE+UurfDQRlsPOAutpTMhR6IMueP8Gu5BaN2hQELVOFefE+G
hM+MJ/DVSjQPyd0yIXG7rQW5+tUbkyZxKsSwjHWyTMoTbPsPyIJjq2vBGeekL8HKbFP9rvognLpj
I/hISieXfwVWJMuD/AzBu2ZKIqfFcVR5sumjTgYWA5YEUE3GIsVWUZIoyGyvDJDhLcB4U2O/AyQL
RZYP9MRYWpe3E68kqdRKetCpMjqr30108BP17/B/B4e+EkN+jGvnh5wWpQYSskYOfzmRRpE8Uo8N
nWRlMw56IAfJ2z73i0+yutLFCH1PrlfaLVBnP/8CNKWSocItGBRyJjjjN6S2UTaCtxZFxynVUoEU
/SKBOlXYObIok/l7YNUzfyyEONFeYOAcnKJ0aLA2C+dxBgMNOp8q9mpTSRmEskYMu/ChOXyGYo0D
prAbBqrAiimWgd9CZwRA/KrfMye18qeGcHHoMti9ZLn0TR9h/Bpp4Q6ikuT+AwVAAZkldRhN+TR8
XVB8FIOUlPsU3b7svjkpwpfya2QDGSB+1SESmXQCrTxl5Ji8QmzFxQsf53wHdNaWNyUzJWi3Poa9
NiaPEgJYJo8YarCrwG6Pq3uZzkGmbH+8G4c1IbmziQZrZjNdy2+6Xcw2mM+1NTICkGyzLxJmt/GU
jwlQZ6bd69R/xcP1tISMvQAH+7jqdCL28HC3jfKV1IPVKumtGfLmjrvJcI4P6e4t5LOEHyjqXFGk
53WK7WRBzzkUUK3QjB/gVuG/Vbg4DjfjRiYTur8RF/+QFrMzsOqsCHblxXcb2TIzOIXlsQKL2aac
wYgncrHYA+rygYEIv2oQiDk/B6cs7YN1wPnY69ychILLJKd7dgk/2nfAHjJj60DU0H14P4kpgL51
h2so15/YWVL9d9ih7O9BGzoKkiLDdWuy4AHv2WegIhVaB4Vhu+LChHxJpvRJdDoyFPRecdv2jRou
3a6P5KUTIvU7ViVt5wa70emfQyfO4ZVpOkw+SMU2BMle39nhh7/OBCMfsx9VXmiAdhZd5bAavrWH
Ioqm0DoUxzapY5ebjTqsizU0P2PzVKKZ8aSHvPuTV776gNKc03mi57a/RJl8ycrptWVFwzyS2W8Z
3P0CXN3oWko/4BesogP8TIKekqDXeM744oQsjYGyM3ox/sxSPrCSNq56S6HHxw+mFErcnWJQh+kV
7pEuz311J7uMs0Wzwjt6G7W5iTSzNTTiAWQQXVaQtZaQ76GPpcTyKCbJfvxf+L+RmVutAjV9vIYD
qYyCTxuc/L7GxEW3PX5DcKT1jt3b1f2hz1WDz3OOndfE0ircYgrDqeXvk2t/vVF3oyszq/8nPudd
VjiVl2xOyL7UaJzafxQBIY6Bgb5XzUhmNicE+JwJWerPl9Qe5pTjWvFSxWZl+8OJl33QUHZuU9rF
fZ4jNkZ96r+FowZKNkTeuhdfDhgYk/VZt8JsghUXMs6qmSNMzD46CPji2TSjohmFCLgDq1m6OLtG
kHVSURuNqtzIItvGfYFOB31q5tImXmeHlt/MHa3wzAhOAGTBjkvN5uTb0GCm9YIGk2jCesGnqhMt
4Y2i/LUbzQae9Prj+B05pPirDPmsCO2k+xxBXxjW4iE4XdxbVL9k2vbfz83TCNROJ1ebAEQEynE+
ilFyMrbKNPnjKovTk+WKoRBFgdDBwj0TAdcnhld2gvyx/obtgVr1dDBX3vHVWeqFGv/t1u4iCIzG
90a+gRQKj84vKiuwSeYOFE9l05g3dUXaZKnhJCvtJLuyLAXA4E2cH0tFjdycju/qMjGB+PIBnL9Y
xwuHCy0Ay3eAzO4EEEKKaAmJPWv5+o+BwnaQDTeEGtj1HdJjcc9bg7fjjO+ylqmNZkQ2/S+Re7fr
lX8VjbjTNr9k4/on3EOwbmpB8vrHL/Bv5jshZs9FlCJdMAZDqn6KuF1DKbi0sp7jkZJOuzb9VDIF
p311Ku8WCNgj8bog9K8Dhintli0XNY2ZtMDsTHqPSTHlKXCl3scBZKO1chdS6iBV4eF9fo+o978l
Cy8pzV/lmGJzk4gY5p0hNZe/ND+zdBFMfrc0/t4p+aUEUW8cJE9UbJ4bd7+Ga0c40EbN7Q1U773V
GT7mcY5b+zSsJrsd9KYRZ1MVUXXjJFj+uGSeF41zcuQz10hcYHmqaJEba2FDh8Xvzy2DVpl5HPDw
FASx7NiVlGnJvggoKH9ibgXrVzHHVZCS/CA5fSYVISJ+kzbSX9rGwltsB4mHMY71sdXeLVnXrx1z
mfKht369akKcGMQcTdoyPqelFHwDHEK8Ox5fao55ZuzQmE2eIXMFbApoHIRSh9MiJWDMzoOhMW7c
peEjHo3gtkJLQAMnma6bjpyBsR78ENpk9f+Kf6spU8niaiHEE9ysL9DhS01sj4ya54edRjGWJyHU
jBwEiDK4lEZdE6ZmoGUY59iDVRM0RnNjW1UkCmoevNwAve/NDed48Ia8/rv6kO+7uN/ydTDTGdw9
WBqavx1KaU6iF9Cgy6dSDK6ixxWVHCKItFzexhvVs8WSPbHX9Y/k/XHu7uV3+7Ze5o0dVl/27EVH
sZ8dk+P+1Loe4xTww5FZinhHZuYVue/6nbwcQNtgFw6u6QmX8md2VsvtcTIfiOhS9PicqFkPtcWO
dIaHccSlhODaZp7WgWyzEgKb9WYGJ40RprO2P5/20UZCfYy203AQ8fF6pnrP+ZiI7DQSGOwGXZ3G
6uvp/ztDhVDeSiBgOYTTF+WQj6QSv2XdFYnAmOH8yXe2P8JZ4AsPCCfZ8kJzrWQ9OEsie6eGpe57
99e0GgIaPPhAzF5ivC35RslucmgYc1kH4Ms5EgCI+anyShw/F59DV9Ww86xyB7GlSi8sOu0Ef5KA
tjIVwI0hWiSQcBJYxriow2Rv2g5z7EbghbCOoAd0jVuuR1UeWvrLctkjnO6bHeQtlUl+PcTR3RhS
PUCYZFSBCyLNxepc3CCQwWFpKRaIFwTA4aNciONvdAChv4K5nuKWUg8eDq8Vcr/nBf26QkJaC592
WwxPuAEowtGA9glfKxWjcLujI+Dw9yDsbZ/IOVEqnNjd300I8Mp956n2KDKtdpcJ+YyOKFZeGr3+
4WkVbeVQBXoZvUSOhX2Qx/Fl3FNFebSkgqoHW1BbirPr7ruasCo7K5XYya2ekGJq9kJcX2VfuTNB
VswcqpebGUuKkbqq9uQe+EQ1saCNvW8IegJ/CqsD2Qn2/0Kh9QBDJK0lIqpWh5cxf87xC+Cb9I+Q
jAALeYnwfikWm7B7xkfRn/KIxG7ecwQi9/9le5yYcYXc9xVrad5Sek5KOYGPpK4h+LwmPvq8us8V
ilJVPZyjIKT2WHa8DLX1ht2VnCqzxbXQ1uS+1FulFgbZ+EGkTEK0yPEFycSg4FboVNmqYh6RKrwr
CzLc2c4+4XGy3nlAp5VYXMvr5h+EnoSS+qF+G3VJENZv6qEIbLUEms5Fj81eCRmq5udJlBL0g2bF
HQpLrM2UUaL+A9kHxVOanMmY5TCnaFd6gMV2jccc00WRs8tZp4wxO9WP+tjAlzFwbPLCJs93FqHr
aIVYVhn6n4sDNrP+1CKdz7YQOrreb1fITTJ85eFDfs9WevJLkSZ7TFpLszahX0lecrPDhVttHhVE
FqyhfS9nf2zNzepreNAIioNKGyRjV4lEwAJcH815+gbmI0u8z53XYImcsqTKT38s7uY6mZiRfJDU
GfLTuCUsgSojr5hH3KES/MHs8D08V/VyW1x5G8ZfA4idf+aD4VoV7B4O1WfZGUHlEaZboY4IT4pg
fLLBMsEfRTR1wfJ0KICwdeH+VW/WF5H0PKWruSK1iN/cwHeag2Ay+j5iDnumA3XN1f2Nd5vLjwNu
AibALHiTNP+YEVdbOyqAqjxZK8zrkVFcNVoL6pkglgG8iKzkW3HHvfVXbSsYBACJA5ZTN2SQ/oS1
7joaPP/U5yHomGq1ZeHPPBXfFzheQ7pyz+jthlPw98Su45TBlUjBw4bNtalvhkcf5KmjerdmcsUF
nJtxJLYUNJwGQ0IrSTREMOODlX1qguJ+GD4iuhwtQpKQ1/qP+AHxwQ0ALxJW7pU+zjP/vDOPSQDq
KSg3/tfC+VkLGz9ht8gibzFUW+i3u32xUxnRwxJ3NxYu8F/B72hlpkkt/h3JNh1lanBTXNRfsBV/
JilxNI23UoTtxBOPky7LTSml3BzhwQh7E8GAuJDwQZBBVxjy49aTe1NxkAvMQPItMEFwYYg5l5Cd
pv6tg+MENebg2Lzake//Jn7DMx/vcDVpBL7eCxXkFzLbLnNMaSxylY611FIETPLfO3dWS6ZfwHHF
8moBorRahoWXDAakHMaT9sPW/+hhpvGafu8rgSpn4R33sqcGWKb7/8RY51mWb9b7wb1OD+hbgvrz
bGyJdf0dfI2nGSDWJYEJhO5s7y1IRvZ3DMw0U3Lsyqr2CeyJzULOmzBHxlJK31syH0WiJe0HiMnR
1XZiXEPtWSt2F18slf7xs8G0KoRHI1aWju9w2U2usOkaMaWxkPRGCup0WRduiP/6TI9fxhlOOkj3
JtfofekNMReq13lO98kSYm8b2pkhgAEb/zLKt+i/bQYRcNhp+UKmEoCAaJkg5NVb/U8SycB4D1Lk
RoWDC22QuUMLzQjVSEFu+DLGw4gMt7GFNtkq3DrtZhQ8Jar+CO1SxhopbQjwtnwvCdnOMjcMyjdS
19Ni5Z+wZ3XYArzfu9zqHeskFoUoFmyA46TqmDECJOfDschybk3p0OStoeOlK7NBxqavlcEOzj8U
0/BSw6nW5ATZrBOHx3xDbBxUmfE+U+smr29Vtn4uqJoTgZOeu4WED/d9dWv8Y/UoCbJqlo9j7TcB
rxNL7ii3DoQMazOGN8LZZVjh2arwC36l1YkiP/tHhYIx6eqqpGEBPx9MsVMBreZnTtQZ2DKHIdwW
EYAYis0P7sxtMKEIJOfVcjQdg/xb2OVpYWOX9XMvA6/oPUnCO9yeoROTt6FD31ob2SONVSbnB5ZQ
1wwTpzsmAbilAGmsx49qtd+/BicMjVBd87rlq7el1DPZasX9QJnhD60QR5oQdtfT/orxbo9MRGT8
U6iY3mfpOQuQLV5J1u3ypp5FozatAA/JWmu1FaDN0mIgSXDY6tHSGxvzFoa4gA6/10GxUiosoX9c
jja2dInOFldBvetmwctIT/Ekrrb9eSgq3IEmVW/bpz9N33QvVa5txfKQrf4FOlqKgSaDoUhDGI+2
HsHznhtTzZBWR0jSjoLWInyA5z3Fg/XCiaQhYbyB8nSrMI3oGCZ4I4MKsX7PM8KhhD/UpuHoma9z
yzL0hhZgR4Merz9KeyQNDcZ+FXiOS1PIXLUiNqD/BxFuSLo/h83rIrQAMVEz7bB7s77d9dzKPkHo
gGqPcjT/MgnHOxrgDoGQamk2CwOuDcRm2lhcYixQvKqeFdQPa6tP1AxAZqfZcK5Atw7dhsrIIZao
RYtnfxZLJrs6LXkquVvT+ULHBB5owL3OQV5VJMmcPi+iyZ4nbwlnZGWQW6J6+MX9zN+DPXUVL3l9
DJAbAy0N3rDSdIb4bEom43JN6NmhtHZCJtaKaV+ORvTykZKpWT6/j5Haah1lABk5OCg25AInoNCk
vcoxOEq9piborzZU0n40BFZYr6wvRLln20pP/WzHcyBCxitEesM0Ih5krrW3ULE6dPupLfXfbAXq
tAxbMChnSKxxxzcvrf+nwBeae9w3GtXaZc39ZP0aNLR/R/dC6JuM4IlMAiJ7h+s0CM+lycGDAQUW
GyLIo9lw/lbwKa+7komQg2rvQSBF0lMvI652VewqoLhfVYm9dj2bo3hyLSC223mC6ekcrZyOzh1M
WGbgkHWn6/MBVA0as2umwozWVKMkyJuT0ySmb1aRsY11+r7/NJSZ8VwquYf21fFpYwgFb8yGk+aS
jj+QKpgSGr+P01I9XgFSs0ZJTLo5ceVRwe26fkWS4CIGCfVEFfNByxRbSHf5Wmdz1PW9pt7/isX/
0Jcr24X+4nyi7vF2/Mu4uOkMXPWx3UuvEshqqKUaKdKjoGvR2atwcCMHYGk97inBvSH5yCW7QZM6
oRcjiqmnJQw3SFoH0wp8y7L+fib/RRH+fzhtl9UcQRp854iSVexTDElQA3LnJfjrTP8vbiuu6jW3
LEMuEPKmaeVfBuus9pMzJ1rlAtD2l7mp4DBJXIH+l9OSfrF6QbluLGsnJ/HDpw0i7dd2qqWHr3Jp
0Z05uB2oBib037JO11xdEUgH+J1PVRPHSS+2/LvlySPWWgaEDbtUuIgsErzcTP4jklmjCFcwazUI
sjamSWuFnYKg9R6zgrc5o4Y71/3hqfdsjousPtYPvA1xTmpIBluOcH1Kdcc9M0kJLfBjDfiXft8o
ODevXeBlm1wSacCNkqFUfpt0y7qstFmi8AC/A5+XZFZyNMAf7Rh02sLqc6PGoSXY2jo8CkbyDhfM
SAKNcR1mPPDj4iRHYKVwdhDZQg9nnh+WpelLzjGeZogSNCzx8P+MCb5/XlrasQKrCUpjw9nmkY2Y
a2E4hJP/hL1WLt5VsR+lxF2DYbbHhHIfsj9Xyb3Tmvu1ZvRhY/Rw3bycmm6WH3RmanxzjkbEa9V3
EGV0EiVAKJn/2B2jWj4mk5d/r+H42su4UcTLFD8MtfD4hRu6Vsijs7l+PHZSLdjlp3soWVefzrLU
5T5pNtvo/U1rsi75rnr9Okfpzyv8lIUUTgxB/thRBpzFME6DT1eLoOfZBFD0gd9CpzAON4CdqvPh
CscQy7Rxu2XstOiOMWyGInGLWl6hYVUPVNrY56J62QcUr5wfThWKlU3ADEyqwmfObQzA/3U29pvE
bP4YiowWDyw9EXfx2OXRlfTtWfVGmCvf0ngaV1HsigPiQILhQ9qBjK/n2AVIHISVMDdzOro+nMui
JfF2ughFSMDUXv0po1gLk3fjVQSM8/3NzAgsO30SAOt+7ZIDWbL00CDjuC1OeigNOftAI7PcefKW
N37MmJoziw0lKstG4QER8nWluz3K83FbkyqDMwLALuXXlaNPb1bnH59tq325uLvPm1OF6U/Gi71M
JQnafAdk91k1hLhBQt/xbACgEdNWZ2davcEFgfquj3NnUcOKY6uSPgzBEfeL7NsLozMBTPkCCOLk
dSd4+RR3AdGKl6vTD79MSYNoEN38GoYh26/k6dupd7Nx+3fpoDlTYgsFTJtNFs+DaFby5/Uuwj+X
Ba29EE+k7eAVmZk5rhVBBqOdpcQ0Z6qYoOkDB0P7chEhM3eEUvWXZYSas0OUqY+5EFs4lX03yCxw
OT+Ddc9Ajthn799FAHJHAyyWPXu3d2k5Jcsm4+JYVeU89qBKqxesypgPn+JNVpsQV2FsZ9K0bQZz
td5aqVF8VVT1uzGJvDX4lFzgtbiHQ5qqsDYKPz5YxPprvOlOkv6oTFsfk3xRbYfk2gveJPN5Uu0y
o04RnuSRJkHq3uzJh4T3JcvSxKryeQkn+9DySd9Qe79iMLbO2toyWQBNLgwOZ4gBG+WoqKMdN0bu
NSy5/pq9yV/EfVPKYh8tktT9pjouk65gLQ//x4mtDjFD1AY4b0JwMcQzJ6Halgo8KTmqml/nJdzO
9kEvLA6RgwhTLhddRrOugIMcDlzCd9RkNxg+aiiVlbnRWBFZfDg8y8/2P1x+sgwwcDHB0mQAs+UR
gIrAgkwzCAxp3RCAO81qErxHaoF3YgvJZ+dFXwelhBiLLFkUHsZIVLdBAH+w39sR+FeFQxpEjcUp
OXrKqChvVkUCHccRKiTdbL35ATVB3WryTJevO599mhqoXRsqLg+GCNhX1jt2rgtGiX7f9c9DWShB
Vs+cql+/UQnVayYhEJxFJuhRfzBco24sQP4hY/32YpSHeZKmFFLRascA89YdIE1Bdkp2tKfbXjjX
m1sidzNBCQ6ZNgDrebVsHfz5R8aL8ma/9QfcDgIPyK3mLbCD+vE2vLOgdz3xsthEiXvxAPsMxXmr
+YWJXZlbUdDxguka2xQxZ5CpaLJ3f8vW1oNFQIbXIRfbp2LbfiiUMw13AWtYPD70dEgFzHGFZOC8
6F2Zc41IDyWSKFL31yE5XxtCAwUdHXcw7HsZuLlQyrsvP6yMBvhfARe9nImbMkWLS1iZ8ksSt5uK
fxBOqMqI1Mngvr1prByxKhj8EFbcvNsNVQLv8S/UAR9JJD7gc+OCMGVOYiyJ/BdzrnwMEMHdUSE1
6SQ+vgkr0DL4TyMKhCOiPXiew3fFeElzEYv3eM+/uVzXSOr7ETr2jrq2liymLBCWo3ySyIwzF5Y3
cp4Ozf3NCKFKzIwgdxlFJwmeIGe/fGz+plb+g36+KG76u7MjBVP8AM/VwQpDJB60VNPsvrokAkvn
1p6QLvfMz4sYWCiu5+IOlr4us9DFfnQCH+ExSOfSaurHgH4tLn+PrjhhoVLmdZflR4rU2D9LZIYS
6+lqClvirXC6V8+qz8yopaYBwXAXK23KYbRFr6a0kYgVbLXC2wUCn5RtzcFliZN8iOcRq1qXKJdt
tDCvlc5gqBCbq4YsuLmHjEdxMbUZqi7tXfYkzIdvsUSRvehIDTm3XiQEU/Nf/ySSPveS3P29QDcX
BXIvlIKRtLEmkOih/yTwWXgChhWH9bCzXOupC+TrfFK8fhZCZgIIyxlTny0bZ/FpQ0JtHCARNL2t
DzwcSowai3hFvi11tdhbdH8zodmlQLeu4sNeXVriz4yTpwQsS8lsCFiZvnBMJNlRSoN2bUpEOAr5
YS4hPrX0HWSvxB3Ud3T2LfOh+6r/3I/tIJonTY8ej1wICkNnH57CPFmDq4VnLJ0XFaA+HqkgeiFi
tNljssLZSMPBUQ2adij+GY9UheqhEs5El4f2W/IgNGYer4TAkMKGTt72plB8bCRW90aklWvvJ+yT
IuOu+CnG/b6pE+yr4CRzA8pHQJTFWCLjF3pNepqeFTzhurNKLCs+5op7VvfPzyC/40MtXBUeMlEw
FNBB9lbcZfuhW8JTfPN53BZRbgdJDwQ1mkcq5cnnvwmU+3AmOaL8wD3bdvZz7fNhTnJlFD0qxJk3
Yxwl48VTp0ay/IRP+SC9tXNc5gFmwvBNhjBX5LvKrt+LVNrVTc0GQALmF4S0kylKbCXG2tn3J9/I
3tDiPTD5BlPLZHejm67+3WUzzhvQJKmJZIQeti+JiL54r1yxJwJZWeABrTxIip2gJPwKxpChI9Ag
mqMD3JAQtWojfiV7nkrNN9cVSVogjxuEyPhAB0Un8Rp3vG2xhUZeQZIuhEsxJbC0cIqCz0fLthLS
FT7h0O4nmyfxboeMoO6HYOk1ADyysNrvH9eYodBU2wTYu8xsCxViT8R+xHvHBqIxkAkGJ9rBCbtn
NPtpyYCdYx9tRZfVSTo+2hhp/ITI4zdBq5X/3DEmHAveTK3OkRBAj9xkwKtQTeWYZMHHycP8Sxaw
4iME5bDE6BIDf6tEwtvm1EOHW0Xwmaa1FrTg9m9Yp7L/YFfj4WMhNAg3iDDOc15R9tP4mf5wILAC
jbBG1i0sKpmXf1RIjM07wm+9ocU38TBF46b30NFxyPGOcIvNRMa2Pwn5qb0nqWhpKGaiIZv4lzEJ
ZV/uIDH18aDcLnXw/fG0MikyHXXkAqdnl74jrHlUjc0Zz8niqeLij0XTZLQ1kOf6fsMwdekMn8tG
Xpt7iTJxGlpu+rWx1SUWuhQTNR+Y7ed/ZJVllYgUJF/6vnQXs0aAsZ/216hzzwoM/Zf0Z9mDYcPm
jTUTEAfUt85K+IKOQHcyPcrI/RwvLJ5k4OugYewO4ViWEfCf9InIrMLyBdyuIWscJQjsVigHyM27
HlkTsg0FefEqQjBw/Fa5CxvwIJlnGJ6cJLoiD0pAgihGRHc7rFPgrCQIz5bNLNCHpJWOMAlNmjBm
0+H1HZJDSFJhrOjJYHXOpqsjuziJe1r0skrMfPPQA93BsKFVTWeNcDz6ddkvMjWYYqTYlvAPnocT
dpH6IUckBkKCS8/jpZaqbtksUiZ4XzmaeUEQ6pMIp+OkRTDfmjQCVIpnxajVFNAmRSGtrYEUwHSo
yQs/CZVy6phP9vOmwtFEW2KBzTd6Rojavm+ScidYFmv8RmCaxXMRaBz5686+T2n++1M+4/vwUq8p
Rd8XPWjBRtj8L+4MB0m17BViGpIynL1fPDZFHxcFqYt1KTghsS1URCUbVME+0SrEdJT+lc54bVTJ
NzZlNDfaLwbD2ixr+K0lQI48rCDaPrTJKeLJcUnvXgGbQyPtb5g9GirykfBV5qIvFtbemInd8qMT
s3D6Yty3/Sa0B6aiC9emhnHArmoSmxjaq3VthZ5ZM5FTNBxvsy9U8P7rFLFk9fXSLPVbEWcABqct
PMSdj8eiUcARq4ufjV0IV6lAkrpq36Ty4JSBQQ10hz1OfpOmPI65zZrbvclinIPG2TQmBrvMh+1W
cIl+8tzu1O0OFY/7MSihJeFjce3kew+DWrMD0hgV7hrToTBtT9D/Y28TqAzJM/5rpf5DIUl7kOm1
fa5chWtsW5iuJcnYJq1Hd2HUqGve6gidyW6bdrjeice6GlrrX07b/l3K+WhcB6vZcXFlxyFKMDSb
sB95cL8Q2hiBl35yo17KfqC0FjeHUFo1xDHSF5aCu63DrY3N6THTbf5V/M6Hqr2XNjP+0xtfvLDV
jFADR+zuRiVV9bwCWmSVjL2YgKU+Gt2oG34SroQZtMxZjCifYYigFMQmaQyXk1oeH/8s3DoiJuot
wVFtF2+lY1Prh6oECq2faxynxvVyzYLsuodINbeA4EBzjG4IA0/bD3kiKy6L0p+/WFLRLvyoxVN9
vvqg/CYiWX6ldxm101avOO3JbPkM+qWwt3HtrbgaPM2lCHceD/DqupXGoUNUX2HGIAss8lTwBgvx
WzbJVWAO13lPY/rehm5qjn3fdkxHdagPE4TIRxLcKxi3nxOxaK3tLnGu/EqAOPvVGuKWHZKXVMZ2
1oz8wGH5jAihQzc4poDNtMDfcB4wFNdW+FxbIvc93JEqBEeDv4j8Hr16PgTJt5SgDRYJOkgU+lUL
axtemdkPcQjgjNa+8Nd24iNeQzheWQvYH8zLv2Rvy5tdaKqu4rZG/qeOPilAXNekiuoLM3nIyVGZ
iarOSQSme+LEIfLkspRSSrmSOzhHjjo35J60l7CpXf82C4B0XydOy4lyFYJ0YlUmlhcaBSY/+vi1
5aClySKY7YJJ73lYp1uARA3kwaaMmbvAw/UojoMb0KyNWgHZb1LTlOwdLzo5zoktpRbBYSpoBNSr
HTmyJp0fnn+pdO0JOiFD2b1pAgxaFsadJE54KPpEEfkD0u4feTFwpAgkhzAGYEqITYCCnXfgFX8y
cRpBZK+M5cnE7zBWjKy3doPvQXj3HGIYWkVQoH9LPuH1Cmrs7GrOB0QWOIxaPzP/lblSfc7s8b03
DQmSTtnLs0njKGFZLYOZ6fV9/ZcBqpLlV5VlyuuLL75YqxIjKzoJNoOSzdGNipQ0HZjFr2Kozzcc
AxixGw0+VF6xUZpz1ntR4KhN6a2AfVQsC71LkU+YD1aBIujqUUCHGxxOn7UhsfifH7CyQHDwTzWv
6JXEgUA+mV3QjUpj+3nPiYBfrf6j9JPxfo6k673/T+g8h4v0OEYRvqZ9We1VXNtChp6SdYuPGN3n
ajGvKrgJnQB/oSCdjzxQ8jsn+rd0o7YE5CPVUVEgTWb+ereAvNigQlNiH1CLY0SE4q7qOxUFbZiM
9AHANZ5s6dKqLJVvmdrQx9iWgp/VHGqwqX6H143pg3g/0ANNgzPp0nTnIIOKQkcSzTA56FDwxzWS
F6wRMt3+wu4CndMRpS8nclBkfgM12rNJBv8sV7yeEVRiSmQLaysMd3zzfuEMEmZdpPm9qWV2Duxa
ESjUiyXlDGmXraqAOdrwP2mSeTzj/YoyLYPmFgFkU2bd7uLKJKjlMQPomc5lJJwA8FnDVzKfsHTz
ua9Ks9fJsMaVGqGVczDfS4p5FfVx4vQ004PGpY6zWQpfNBEnfjkJmVE44bcKTVmiPuktHcIZtF2X
2fbnW/zHOiSjlXjbvLEfkPetGCYqTbrozlMecAj+AWDprrxMEvUPeD8Qm2FEzJo0+DGxFJ5y/koE
YCzLLYEr9haBFPInxKTQmIV45kXzOKv4Owr1Nv9FrS/NJtNHav9k/6PzCBnWYqwgxMk6aVJZSgsH
SiH8bvTfWSNJRZIk4gkWCjfHryllhNLgpyX65gAFK0Zw94/5LCd314LaFgjRxk81/MgBL/jRUM2r
M9/aVjyMxmWDq6DVUfOFE0lQlmr/REvKSV7Nbdz7ZB7P8fx/nlYgsB4KYYmghqrA6k/nHERx7J+/
AOprgzQ1tchag82Lwbj1G7UmmATpM7kFvaOJeH8CnuOpsWP0z/oU7RI7mB+Spj3whoBJNplLDAZr
RXhDseAnPwsEP6FyMl3LD67ERIZmUSLah4ii0RMEt2ZLcAz+11K4wYj2vw/sHQ/0B+SPo8v4HlAw
AgAT/OKGrosPfJknLw7y66EnMMemnwsRPecsx1eloCjz3YFXqgI3KEDrXLt55Jn4QiKglSPKtUlD
5EW+/GqrN5M8I64eVeSpMeqfFx3JkAEcqNeFHWXCbmWo3WiXrufAYN3I47TSmQpP/HhDMtsYt0ZN
V+cq/Ceotaicb1VckDrfangfw+hmeuvTlPW4pt+Z48Vxn/50x56gK6F0O+84uVkG+orR5s6B4GM6
NIkul47u6PwZfOh6bBzUXlCzC8FSSXuNc64PnE+ufha5fHA/y/67mIow1AVOfYyTmmH5iJAqa1gC
zlBY86zFvg+pUI02lC0mUJlYsaKy7qO7tZCZGdxLlIHwek/2vI0vam+Z+4G5XqrYAhi4f1gd9JdP
/ghkSG2L+DRf84jt1MlAMmjjDMdI9K83k+qiWCm1lk3LIGcKRH8AFpTuppvARFP3NUQ5iSRoZ/0X
EFS3kD/t0kVTiAaItR2ZmI/3/Nktr3pccqysCyuMqZ5b+Cfi9LtYOd0QrMXLk9B9O1BGgCz6uPkh
xzkttqZD9olDDtMtD0zhJxObZdyWLqQcTFcCEokTJo5cYp3+HCATiJv208c95IeSAczGIetasAvl
bnfOrzGu4x92X19yPvlVZ988frdXQ97CHNT7g2Ldoe4gTW/SR7w4p3qcPLH6tBuiVVJibZTe+VoN
5DirTXjTFhYOlkbenxJAI4aYW6YMuQmghuJh5qCQV9kiTbOP42vJceBxmy3WRizdXK5ZhInmw9FI
92mP4QMEqReSTLhd16Rjt6/OlMyGx0eFE7SKuV0LOKXdNtnBko8pmsUaXyCmaBng4Y2E4QXQWV95
zcNhC/4IUfQiuafiI7G0uLgVKxMj+uqwYUPNdOu5PDX69LfgTXhguKATJ42YdA1FfZnAqPDSyQmA
y+6DkkIFvX9EervYYQ6uMgVxFerkSzR0WBO8+FhQciZK3Mc76RlgjhCZtYj3nBVtuRL6yAZ4uBRs
6OF5mIVXQ+jCVmbkENhSgNiqOZA6P1fcUS6sINMyWThjCEfNsaX1bhYIHkE8Wxj1hPD40sRtN8oS
2dp5T1iqWVOKI7r9cXVSgt7OGoOqD2mHmiopgzUAHXL6AME2u6JWtu72CZB+kee/nRiuRHSY37l4
E7yJ7MHFMvcJXHRmlPCZkzy6hVy9SETcKjV+UOxVSahndi72Ro/cByuytCdg6cb3TmVpea9JRbDa
rDuRlYI30sEn4+mE8ZgBtrdPIAHzB5VVC9mW/PjcFeMBQKQUr7CCN6FDPifFATFEXk8UzhAGLph7
c8xz5NM43+kKh9VZNNPA84Ho8z4qQDPNXWna93tYumUoUeI8eGCGAbgOIvjQJUBdrcxcGoSWpv8B
zlTsPz2McuI0AMyuZqH1NhwUVvwsM1OV6JBRgQ4I2bSLMdRjSaOXFs5bgBbcNEcN2rCi7COnxhyO
5qbrl36BF3cRf7igqFHXQDOzmtWjRzwiN3P1EuDSZggd6AY6wy/DlFz6bCFrS9aKBw7jBKsaLzje
aKaJ34pHPwcithPv0pbhDgYpQSMtIxe2szMRYpoLVc7yuBa0avoYKEikbUaCdFyrTujw8NiujUy1
MJftm0AIiMsO1I5ReM65LI3Fnd7XbTBk8TnBtiI1FHoFiBtWzPCiMInlcMW1kDed59O4IkIhihvY
gY3vLN2qHOoDBcmXcuUj4nHBd9ZdFDnoc5LJ/oS/N7nLu875awXNNjjZtRlVLYmB3ARxKi+HdU0N
3wn3+DHJ9kUO3DBylmKaaM8bqjHgsaJSR8vZ9Wg5pPdK44ZNGkHF4vB36pmFkbf8iXwlfqb/GbWG
gaCE4Y3b6YEDLreh/Xs9vUl+1ES9cAIWdvV6GDFviF64o1YUTyjU520Xdrlv94IgRJ7QVy8RInO4
+OigQ4XagE+ganD7LbNNVfwkyqB4cVbxSjO5H0fp2/94R1Z2bgsRdKPAaZI5U/KG7LcQOdmwdZM2
orxrWJw4XrfZi2lZEd1lURODYsXeehTkZwwtHQ/irxMfJ1TzymkuPPRCXUpaxlVI/8YPFTI0YpX6
PfGZ8i81BDnmBy+Fm6LBTkbjMJm8C0fzpRFG4L00BXw+0uVSg8DA3bfhoplSRG1n3cgCYuxZA7gN
eH2wSrdrM92ffqmhbRuxqGDoFowdvfdFJMOwtcp2kLIZGKvvuMiNdCG+ylICzqG3sGdFEJzUKTZH
VpbSKpyPqtDCIUqd320FAJdRr7Mo7m+O0Qt5r6jnLtT6XyZB8JknZYSfnZyL9iAE/Dfh4i+tsT/d
R54qGf+B4nqcNIXJCL2wUfvGODAgdZRGIkFFiftW3JZQlSgJe4CnMqoFIkSVj1iW5wVWnEEYP7yB
CIefFZZY7ADDCo2ZNpk1fsaYVR8f47vmwsP5GFO3G32RwAEkuK1PO6BXO+hM2BOYyuOJi69fnTD4
OFJm/C2OLZI6Fnpb1/d2XLfTyzyT/qoD6TWz2hrFSR3stjNfGh7gLHZ+3GUGaTNifSSQFWQueib3
NbQyNL7Q7X3Col+PcY0ptqMSW1+cBaNmZ2U2zrY6+awO9drrqvycgj5Cq2PB5oYpzuOL610FgAqR
sxCE0pC92nJy/WVGSWf12eFW+kNMfz4PIa1bJ7sVll91g1EhnCJD5RnS+kkWyvgtvve9+Ope0SoN
/Jy+2xNZoTIBE5MyzsgGJI8Q4J1d0sO+tNMoOcrnl5ZN774TizmR9xD1Q7Bwzig6Rjd4HMPriBRu
/KgihXgkoilZxS5Tv1wMezU2MWzM1WxfCZ7OSw+h7zvPC81gc5XJr5DaOud7RwfOhZa7J1CtWSbE
c+r/jWT+8JRULSZkzA8ivlt8JczlH11N9/KsfjBU4rhFipABVYIfH9Fm5IAthbLa8UJLU/jrngpt
ibNEIicWbFXfUFkXLoOFTJY+6V9Yy38R3xuedfXDJ507M5CA+oOxhes+lMYXypUi5/GyJU2vuMmJ
fr/jpK4Ta6ka5JbkJyTBMlou3Dwg9zRe9MgyI8Lq5vX0L5KlBTXfQkGvspENyd6kqhsCFS+D5ltE
db+HnoRZqK5edoyHp+hVCGYJpjjukUML/P5sNBkbAKwrCA6KK7FMzQjujvRHCuErnRphKWVxklL1
u3AZCJEa+8lmVcFhMjAJuJ/hMAUDlkyETFnLiUc80ApGUoHuD9rGDulcmEf5KyhMdeAkGL9sSvFX
NsjXz6shHCRYKSfJQhCb9B78/cG9P/FZnwI5lTIuJzymXgYPglsJxWpQ8GEbqOPUbMLISuiluBO4
FRTmqm+Kp4Ac1rfULAlor8Qi/fLP/0A7tVrVDtQvHfqhCBdf3dUHzWorYS7r5NBIlS/z1Skqrxt1
mGOBPPTJl/WtP31hFRdg4+QQJ7eYOIoaOdAAhtrjln/uhc1lT7DGG6Q4+DUH+Ns9yy4fIFIeXBWn
RbTNDf0ouJ7YSu5UhPNcokHmaHjinMGcTAlaS7whQet4fAh0vlwDOdJAlsVMFqsFCyzdizGGtqyn
sNcBKwv5PB7z3P/oExiroWk11X39RkWepWePnRPCuTupzMx+BbGz4rnGVxMhCm6ddGp2Vz4/QczX
EIfHELOegswDuY5XQPEGk7ZtTQjXk5ezPM/KYby44iHE5SDvtDXxg4LWyJIotEZ5TdHO0+YELwtP
yWrtgI3h0Jn6Nq1esu1azbb/GgtqxfuNvoCedmoNBPcdItd8YzbGTUNV4caIoNtG/bSlLwcJNasQ
bMOkEVRe9rsTyJESy9y0A88ddG2rHMo9go+5oEuPbdGS/ail3rGCJhgcarew8IR9xwsfBDcKpTsd
1Dr37aP9N0DpDaLcoaWCJTUH0UqrOUaEcelVPqO+SvYP8AI4fL8dzVL5CtTAGQZEnZHd3WMNw9n1
XIsCWSmL1FUtp7FW3neMJTgqfQy1+/ff4NaFJ5x3g7+T31CSZQEeSnm756HSxvqkKfUEpc1Jf/Fr
RG5tDNheZ6XKB1DpWJT555UiDw2cHXnTVhFeiOosvCQUudpoOZXrLYVjGjZb+0CT0D7BSCOPa2xJ
S2V009saRyAaR5//AapXTaThshRDZzhEnIfNE+OHLE81cf4fA9wudP9aejpVe9ZmeWaqwrcpVHgc
naeTBjCJs8G0lyxIQgSMmzr5ITDjzxsvtDDIKpYT7Wul4xCdX1wlWFe80dxzAIptYCW5DqT2MwLJ
timcfIm1+XFPb5flYjmCDgv0PV32DGXZBjbfYxUXlUPQnTkHu5wVxkLTEpVFI3uPoeO8/0PF4W/a
wQ9R24pkg9k17cIYeFL/u+kHM+jxJ0X5xxdhn47Jg0sKgljyy8nAhpDlgnk1vcI3IrazrNTaYHZ9
0bP8WczP5dVRf0Qq+1W5Ab6+aQsCZfkSaeHBAaHtu19sPztInTBMQ7mtOlAwZjiToNvdPQJMzqHQ
ufPP1pAVnWrTMoFLYNTfILX77UQ5Taq3sxDkjxAmWCaiwTehfVFxtmwcXT85HwhBBv2tZJY/osau
SRNo/IOBeTCmIuwM4FX/m/xx7CphtxIdpUgMX+Mcy4iRpF5XlSSSn/J0ZNeoY/8CGUjaHEOCe1Ek
qgaQW37zZQYLBa0Sq1xfha5NRucCN2OMeCHeqFvmILtt+J6emDFANWWtXfqmTb+k7GGh5dDsGdk6
dYvCNz0MivGcYwsGK1St5ofmknmT3+QBvf5xWgB3ZZ6cP8ZdEklMy+ZGguvm6d6xdNvHLpC79l28
C09689rVWJfb4OEioLUY52nM4RTrm0ALFaq/LigPbvpceRT70fmr7Vtq64Im1eGQpGuL5sfOxfOA
ad27QH/7gNOM4+Jupas/hygmW1bg9oF9xBJ9A9uaJGa5qnfdAZFcKawb2CpIo4SN6dYOPd6GoqZi
B2v+maMcRoxmBRY4LoXvCBXkFi1/3yEMit5EqqStSQajsqrv3OP5yQxq3nygKePk1ORMXxQ+VboO
fA3rBKDHNucmBE4Sd/bx+T4B5wvhDb3b6E0+wlG9uyacH1+KUm29scW8CxqJoODgBTt+8u2FxW32
pSfVqs43viux3J1C6jBQaE71LSyWNm9M/XzwkAtGb2B8KiyKD9asdKwWry8f/Q12l+gghK7TNdlv
MI1d3uULmv2uLE6tAwEuK8OWqITweIbia5sKCOOGBoiNzUqKwsgAP7NwsvzvHOZS3N+iD9Fot+g+
27LIInU+frqenySaq/G/yG8BFerbLuY9TBfVTBVLxafMafqlSvwQtmHZwMMEfKkBt/ioK5mJeW0i
CoKEGFuU+DiUrXELkfQeU1TwC9F4ULMRrnnxG+ayv9jh8lSLtrAhtD07mE8KK6tOQjY7HgLWiMna
T4yJ357Dkxy8l9LjfKKOrlMIWKbPRU6/Y3cWZpFCap/A/Ej9bOJ+8Opq1yaMISJdUbKw7ZjltqoH
z+gDIJJD4uBMJGjpVu4T/ucMwdr1JhOeQC/5pNj+YxJD3dFqXmfaY+l3jqhMTsFtzOODrDlVuAzv
6yNJaGpcsyoSZTxiPhkAcShRBfvYUB91kf0b/fIf9XP3UNvfPAMtYEDFmL57LQ9Bl0av9/kICAp6
zz5YwqT5S+0y4fIHZRfEaizuvcmXLjUve+hiUlGifBMR2CpgLIhbl6yHbtqJTsqXZujRV/StbjG+
dkxIUcIulCSqFP5O6hqlbR6ODDuI/yNmPaUEVsUJ7hsbcpdf4ndCAiL5t8DyAPswBq5Ob1opMLVu
CKhGOW8e4DRp9Q4TC7gNCbeZFkeYeCqRtELaNPCyUb0ORF8YT9n1psvgSobrcauTvYgojrjoyFaR
WogOOdxzaFVTl1cSS+QXz46+QPsmi9V2/ySEgtmK0kE2MSBjQJsQ9CE9/IPOVan/eeRJecRg5oig
SS5NVTt3IqK27vZgIu/wXvkZeAcr8jAlvkwBXrIuelw0pm6nPKyRBjeeeUBYudsqBdM6Y0wPYBTw
U4fd193LCmwQzh0lu9lbHRppYeh84IKRkdGhGwe9bbHhjtbmOIeQuFjP/9ma7UkUCjcRodRzgoqA
hUfk8bhzh77Ntgq+hQ1TOkCNEkRXjATJ5k5mjIifQ4JR7DWaa/oM1wHudW/YkkevuEMWShGm2hxb
WH7ktnOXyXygZW4KWDSBq1gL8z3UPkGLZT7VBtvv7E5FcllhFcF3tF6BuH5q5t77xlWqdhgYUgnE
zneS0NJ8hTtE/TI//HqEriJXAXmUhsoRnR4wz/X28oadKLIUuUjd9OBcQMw4s3CFa5nQlEeBuncF
55t+I/cEV5jXBGpfoDbnsJDha3iRUIsrT//V6N/rdJQFJPu8y9oxxCCK3M2Lbf9gRzSwgmF01GMQ
ajnObq5WD8NdOvPfIbLaq7WTn1N8jd5vsTv6wLHvPxX96r5dvXb+ELacXwy7707ekSNVaDvmTMZ5
oylKLAcmsMPXf4e11cUzdAQiMlFBSiZbC1xXi2NkcRa+CMZ2l2araUL/tY/nxDwftDFGBD7B25w0
tW0Vnp7zmJKg5pZfgX5IuHEtCsKDzBOQvM+7f8u5JyE8tPnIr+nZ/qjBT6m6WOrYfwSihZS4vYYw
6T5BVQ3vOFHeE/N8Ie+yoYIL0jIAH7QEf39h4VPYdwvCH/ZHw/CVwRxpehSh6ea4oT4BbR7m5eWE
0tfecGO5YNrMC8827/da1wy3phDq8i/aaeLdP1FHfXw12vJWMDbFrOCSMAYFYQIJ8mb3HN41oql/
APOOM+1sGVqUcJcfTNuJEvFgsFRXBbEFpSfQeYsjw6f7OUWdHJMmW0NDpJ4PST8nRq3RHyob2EvM
qZj3XE4oqgDEfLyIdVXWq2V9PwH0jrxKJ6IxSf8cAcZSterBFw6TD9Pns/eU3ZCAp9ToNKAeQaGU
Edc0aYv+k6lFRm147dbg/+gRpHCiHKDsng4SOC4D8M2H/jOhpLirZHJH0vuyxcEwYkb4PjRJ4A07
0I10PzDRiVPK4mjrc0jGfh3AG6FbwIv2dHzFpINvlUhJNABttwzHaD84+6qmcTGLwW/f/lyi/zoT
/PikTliLJbD/2g/oW/ITycvAnFg4ntqeiV/dWgdbftk1wljG70nPTNqUi2oTGAZvV60B+V1yEABX
qzbdGfIXL+M261T0+je2YhWxuwZ/25BxFFlYnDeA/IsaJmIMhK87pU88K0zX4lKHCP4z/SYv1SPx
FvDapackW3GPTqHoZfSzMzAt9YA6LDKlAnUxR45vUbtpqgfkdjsz+NMcW1B7narS+BpXSt1r3Dmb
+Vo6u8oJ0Utm0vv1S+xMVjI3LG58sL017ef6pxZKpD0csVe9ZHcx4zDV+i6s5QfzUsgxSt6sT8sU
XIA+f7O9SkA9TVOXG/yQvnGC/6Jx2liiElavH0WhYncOV54PFRBFC/eA6XAAVQFZneTUGH/zHQA+
tBXn5zyydF0DQfcDB2qvF9YJkpUJz/EemFDofJxxi8y2LbKK2jM1mBLgCFMM/rmEf46Dadb0Q25Q
ugvVl0B3aio9fQzZrlDnkw7qApv8A7ljrqKTLEYSqqQ080B/1Z62Hu/E9kVeV392aCKTpHu3xEU3
SdUzXXGdWE3jS/9ugcmwSxbbrLq4f06YxeNMOsB4MsyilRorjD9mE/SZt2bd4q/Ntrss9ShiG0c0
RWCK1yi9RRv/xlH/lwyFrYfOOZ46aB/aQ5FgfwdPPaZCdPMjDwP2xUvldmPb9BPzhjUDmZubUEZ9
YwUwf1eu0j2NWQxD/LbqlnhjKw2COvuIr9f2hwElv1J+55mn6OdddOvLWzMNei9OCVq81/PCXyhe
wiVd581VtZ5yX+S31G3BBIP0L7Ss7TDp3JqgmOUDglC6Bg5fUTYEdjAKf5N1Oni2B8AQdU5eaSwN
JaFSSqnCt0tKcrBxI0oNXvW0S6MCHMNWySGSfDCOHrchKYTwO8CZzH+MKW/8HjlF4pM3hiYEsDJZ
TO129Txd2J9pwS9MXgmK94/tH1FC0R3byoJrAoUwgnn1tNtKtgD/q8wOgQ44tAdd29P8frx32jyJ
WqScLM7vB4jgwpZH52lIoaujWDloCjs+Fd1WANXe5kCA+zJef1dEmZE7fkvwrH+7jkSgJf6FgYn0
L71vRwl1iGShbVFVtEEORj/XhXAHBzpP238xH2u9tFM88Wanzqr30QPQIr7xdwytzHb7Cgs2apQh
wv3kPLF7AgoMfOTVxzWPzRa3eFLrIljBpOJEAKc+R9ZJQc7YaKw+j1ZyZr2JqGcUSVyKuAwNmg6J
cBDZKVvOyLMIdfBc5ylX7BdGP9TDpdDbX2DOnIpk/bBzYMPWFROM/+23PR9S+UjWY2ETdU1CZFl5
0WFv8mheWW0dPNMhxBUrM/d7Yxxh4Qm03V4xpEnwXGSoeJsgqZWoksy+jWik6ng5xxaS1x6yij69
F2rq9uE9wcUB7bWAPxaF4c8CAWi7RQWCRO7wjtdFOR4ScZrw1AOWiMr3Ig+CQiW/Rd5gttADPNs9
qKfly4+XXq7iSjoCRD1SSFgVYx/tWBY2B2rxAo0yKFuCIq03L78+WCsxGWRKGGOe8atIt6mjHU5R
/DrxQoW/8scBG09pEYTsBdcSWOfxGOM3vD3VP1ReBs1bCClH9Ma110o242YlxTOKfetI4JPN/Qdw
fbGcPLJuQU0PXuUZM0uGKzjApC4zCloNuQ2xblK0Wc7ADTczssI44vzvvD8Unn0kXuXC5rfxV7mh
nNmwNTlgC+S7qFFDizSJzgt0QpxvltX1NRa+7dNtl/DHxaIWZ0y4Hbee02W+5yfQsahaL4dInusC
r6UuJnj2XcXmlveIRbnE+i6dtNehEIv5wp5uFp1Us+5Aedx0kyjDGxX7xlUzJjrxRCex+DkAwQcU
qAYapogjrVreWnvNqU5kk+X5JU7+XLujpR3I9EWOtF7+tzCLW13d5Ht8pi1gOK13TAkj9DWqxvon
tko102NXV/pcPUtO6ptXSynO+bvAIbZIoTg0dXGPBr3oG0ra6PqhK+qcvnoUJDnhbNsPDmeKw5Yv
nThvfAFBdJ7mE3HOhB3sBPXvvpIrbCT0Ev68g8faqovSRgUtAuQRWAu+96Lmu+0MBYLFwJNUj1gg
yuqGEa0lNSrRfGS7GaxRBGWxFn1W3jD1q81w0KTHbzU5tItBfSAQl+eMbSYr0BPXf1qjeXp+LDeA
TBIENkxinqV7wLzzhdgJC9+643az5RJulG8QRJY8gwWXWZFsWzbGqUHIG1bHZuyeMigTWi31H4gv
WDlrjJFbnvHlu4zQKTwx8zZRWMCiHFq1C5G0pmXqpWnt5OaDkktPpUM0hcw5FAHKvLXTYpgkCIW3
UHPZ3q+tdaRd6fIliQrxgyucffvwgH6K0MrxCOV4P73vfYAPAnvQkD4IiIzpHdtN8QTkBygWWd8V
IRpkPzYLgPedgzOIR6bx/fDFxyB+VZUdoAR4BfMsLsdu+nmHfhygAlQ1cp9ntdKiCO+J0mcg5G6U
YYpD7nENwY3zwEU7TEc3OROQy+7g7m2nvluezLegxgnfgUWnj+PC4uPH/rPJrygvrObpd3czKRic
8rLapIndcpBLhAkKAEl3Q552z8MtvmiAiRareWoBngfO09XLBwL5TDg57j36+lDIwTEugb9oEblP
7LE1zSPx1/n3iOxfLaxdqfNDmSnBezx/Jjgv7SUdyr75q+Oe99+mOr4H92+DFtvCAGK/2NGbmIuh
xDu6JxPqm8pGQIwyhjw5OBUyi2pXg8auhqXkGmRPmfdAEp4FDT0wUvso06/sJgcUpfGUGshEu54+
c3PhSSd7So5SMZP37tRsF3VyjCFsZfj7+a+L3gzEY0DsKtQ7XnwFjuWSozrqpDhVx+lPsjooiRen
s553+PP1+U4R8ei/u1hG4d1Fh08r3uTDyjxMIjONB3ooCTCCDq79YcdceywOEiNIyv66/G4pWfPz
zXI3ehSAG3ntGl2TZ4FlHSaQPNp0Cf7qjO0e4/7ZH/X5U5gXixjC2S9N4Bl2yD+7ITbu2hV64j3p
QDIPgFZdqZtV+ZcVluWNE06ZU1p1M2sAvcPx3zeBpGIiaJxHVu8xlxwhnEfNQ5cUmca7IxdeYK2N
QRb0CRuGAsFtYYTaCjtP4ZexFkZvL+pA1IR+BBPmIk8WuwfltYysmpyXI6ySXIGzGabjP6BAGDJP
N2IfO50xAFxv4wNpxL+QeWI2/X9RffBARbCXiEzwgGUYUf6jEI7fL5xRyseuRdUP3jEJ3rZ29lxj
Asmu1MA/7OLZ9TW2B6BUWxPCeJyCTxhc4meeFqvah4vdZLkuAgLCldW2vnrzXBQVhba3D1JuGftb
ENas7xOIKn2ZuyyzqXY3zxToAY/5qSegF2D8T8EdYJteQplKOeAuVuHre6mgmLGFlik4ab5ks4tX
RDm41Hc4zikneRqz5I35LLyhKyseCV3H8qpplmexqs5VdnmcfA5UhYsPgAagG+1ZKF0zIaHWAeJi
UPc/8bpAyuGXfZnpVvFrndidbnZU0PHOr5rEWJO97yMuEtzsC6mvmatO+9fNluUHsjHi1lOI5yg0
HjxKI4NoAhVYgD9NkkH9CS9DD50oh5AuG64Qpwtd+b+oArSs4AwVUDsv2WLuevw1LEWnHTM9RuvD
VHFGXNitLhy50DVL6mMlMw4Evpt4UzDCd4Lx3yCm4j9lOlI5gvydTKg3M/mHp720RDdxGMfsVIhi
x9RavrKr/stjg/pLSHoTle+DFVeUO+V377DqcJta7gd5VCAyE4/hhN+IpX//PhGto8IzCzivtYK1
WwP2pT8C6mO5Xjaodk7dgT7JXbe9tf60eidjah3GDqjee/XTkGJkXKIeWjW/o4NT0e2CaZmFjp3O
SkHAfab2BNdje1DQeRVfhY2gm3PExqU3+zNCLeIgGTSK9fDulQxY/NiT19hhNACtEx/+SyzR+VTO
No0VzKeRnKo1KmNTPCLnODQCwv+/kKsNwV5RlaY32qusxSCGZ3B4Uoik9YG4dUYSe6rgRyRg9C7c
MrO1qS5Lq0DpURDGkkxO11x4tZwi+6HQTcxa5VmfXmbzf//SlCjWyz72bIEGJRZ7XbnZbaLArbZE
7p6VM7boQbrfJ7IZ2afZEy2mGAERtaIMCf9XnvyQL7RR94Y2br7J/js7e8kLKH5uJxox605813I6
uHkZQDd9vcVNgbo7zy1cJyEmAivEqdY46eABFDTKx5LWu/szfZFwQ2G8IRbDzi/7o/Yv5Tc3fZRT
c1XLad5iHPiUnLjjqqAvBxXcHdm5pch69YYS2n9QrET65WyJ2AI22Y/xaA5Fm/BiqFsWW5h9v6sW
i6tAaXrEaGxIvgUm0/fgGg4MX8l3SyfeGCsI//+wfH2ijMMKpoLnkVEZ8UDqL/QzX810rx7tNwLx
G59oXe65gI2WKoSuBPBw2wvhrqp/NUkxiFbM+O8uylF59JiBSDYmUaBwpg2HkJ7LtLr9LVyNJ/xb
7/AMC6rCJqDxNvmxEjvLO5L53zWJBubFE4a4t7x59yc0DYdgxG/YPO0hVGVWgkYyDSsP8Ql7AcPR
0MdgWy5tjogbbe6H0vu1GkVQVhxdRp+lz+e1tw8/W1UtdJvay3bm8fOX2mWbEBVE12nk820+gpan
x9crDkCQJ7A/dgsHkG83XmcaQaLtCaVYTaTNgioOg97RewP7ZDwlB9yxcZFh0dHLymyTfa0O3U/K
eZTpHProdUOkhsva1t0KMyJMB22EiRXuMCNuSModSjeB28KI01RMfFwM6Is2aTSyWcMZxRUXMOWj
5idLlgU46d8LFWCLOR6JbG1or/aasjZMj7iuHNcy7lH49SxG9eleETqriXAcftVp8oA3+NJWxFeN
fHtQ9e25Ak3kX9Dnxq+hVA5xglUZKM3FIBxHsuP5FQbKE6AMi/BWmPMMuMII926zC+QIN3cr+RUR
HmbmyC2C0+z/Vt8IXB7WzWpyhUeZieh4xVIoUCqGgfTkWxHi3FCwPsZFyn1IEXsHUAYS/r3Tun1e
Cg+EsS1rUlu5pWQuResJdpTtN1SGryICHXtv7mitALZEAv6xPTOL2QL0hjUh92I30ZZohbr659U2
x7fBOQfetTwxatoOHK+OWe6Vyptrd1tIc4DeWeK5+cq5Gxn43Wtxe+XzlrOOGCmXroZXs+PQ6MCB
crE/syyhoXW7uyGVuIl3AMHapQmHSiFpNBvJDYkJj062WwP92SkfKbmDL8pQcoUCmX4f1oqhSUJW
YC/l/iU/KeyU1jn6gY9Wk/Zoi48QopUSlqcZv1u+FDm2e20DQKs2z3AWtMyWdMhu+3fPHsdM35yN
AufMEsCTDtbmbT28qdjOm2YwLSF9cRyRJCw8EnjbH1gwamtIl9inqHmepsqbRgXnk/yCdMwsnMng
hcbjNhOiTHjDX3Ych1TEIB259nwoglo6HrzVSYUdExWcT4PQ2r/6qtGWWISOvD3XLvnmkTvtnAeq
ZeNyaPCrRLZGWHekDbuJpRHuMjQGXjbCLOP/8ah4PsDVGL3yDwngSMQfFucE6chSIzoxjLBnAgWG
HfWi9tKm3N2xSrPxxAlpx4WOHDKulwE+EvCu+dcOfgBqv6dwrSZVX2OvYLw8CkTZ0Yk1i5pV5SXe
cwhCbQlgITeKrY8Rhb4Qivlz4/29zokxBhiU0ga05R36sL6q4rM4yY+tke/x5HcPX9EzaCzu3Ssx
44AwGfeWPT0dfq643zYvStfpNvDmkNOHbhtPlyOWvXR61jafIgyBSTqZejFxKaSaouYEXPTEZBw4
GFoPsUCI5k3MDizkjYgF4vCKs5egNtTXcS7/vspY+ksZipDjV9eqk4YG5U9fJ2bZV/8VPo0+vNDq
bttZMK6UaqNEMc+BUop9rmYCWOqeVLdX2a1bbX1VyzhdY3Ugy+bJOoQLIWuY/sSrGBtJ7pQ3DEBw
tMY6BmVF1YDdk00FOihuYcZYdKV6JwXQGuzqaWz04Kd4fQsoMMWOhCtfM0e3HNnuNE4NLJvCAI/n
j/JEj6RmaTom0N2pVHOh7o+605kaCt76wCKjTXTjEJ0cJd98tvayHceegQDeU5wewR25nwIWH4Mr
eBY2XLcAwx5xtEIdy4STPnrqBS7H4k5gKbV9GFCfHrQvEPgKnB3l1qO+bHlPQrLsA+1fF65t8bd1
RE6qSvR9ulNADmdiyNWeqMAILWmS8dbfKMJ8SbExIhG0Ha30c9xhC4jJrZodMS/lAJv6fyayGkhE
1zJEblCUDg9bRqdne0ktWv9HhB0wkntoyoMFIewLnpVqbqBA4qZOx/QRHnM1t9z8KzANFH4IfGA3
2C6qChEKUsXcoMikh3FDeLJfJnMJqdo11JB4GdQpNCfSASySfsqeC5sl5oobCNISvIO4p7Jx8u9X
i2ryMUZz1+9wpcXiLTd6f49fS1Ird2kSjIp4soxbQgynV+7+ayvUHPoDieDJOnTf5OTGKPd7ZUnp
Ixq/GaiLlnzCYYPAUN5znkYYrbSgRFWdu8qwVrRSz2ggUTL7PyulipabGQXrMhws8a5zQ17fM75Z
FKdH4sDpdMgr/HhLc5ooBrkXHepueoHKa0Cvjg3HRUfPZOVRk9yEtRIWYvYcWgVj7VygKsx1+Ueo
0VA4J6FsqFDuVyC/gp7tP9CwJlfZ/Bxk5a62QI8MKfvTFEw/nZp2kl+rw4bgXR9kVTDwAKO+wsu3
EE6UpsVLGnvYB6A3xRiiMFcjomRl6wvmA/23gmwG8URK8aiurF4gGunj4y5QcPBToeBqsVFFh9xo
V3t5pr2/Jv9xoeAMWYu7v6Qakmh9EhwldHFetztFMnrt8XmG1qSpQLHzcaFhJ3al0uLNEpiw9xwR
aMT9j/tYRSYo2eIXkw103Ljjd91S5lqBkSDY3kkPnAaiqPgDhsZVuk6KzDFkAj4B2v8yzTD5Sk1D
FuIEnuUkY82//sumsznA4mxjbzgj5EGzGrjEqK2/CUKBYIzrYlEVskyzb8o0hJNyM3cQg4dnm4Ef
7HBy0ZlmRSa/NPePysWUUM9nQhDCH7NZ4Jj3ox/5CQ8VdhpYq8ZWM9BDM/WfMAMkVWAqwV5dDZ0A
q8rao1yKN4DOJBHy+vO40Wi3coDSKQlsHihSlJqICMpby5adB+br7YmODILat7s+Oryujd2x2TWC
P2LAtDEzTfkliNgen3Nv3gx+CZBGIXh5yqa02NxeAr/6dA7ExHrq/7NUzkPt5Ka7UmW5QIVbuVzr
Ajdn8ph5QecAGf8bOD0J738EC4A6c83X+AH+2weAJ4TloZ60vFiwngzdCBXyRjuk42IDHhA0GeCX
8tWs8nTt63wy2776PHNW/YP5vidblk+X/RPE9LpwjaskPjN2CelnsQbm4hiYYhwZutjC0a4j3zgR
mjZGGQd20HORhMVSCR6kHjIZ+9hH1kTYCxyhcCnMOEEDVATxkm3806AHwbxpIEgfK5LXzmSdlBf2
YxKnUMNq/0cYtQuTG92g9Ok+3vyr+Pud20vRDUc6mRbp0bJcfTXtJLgfqJ5nvG2mjF3djISkeHv9
pzCr/Pon94Efu+hg0OwiSq8wV+3+F7CXp1t8EZNLfiI3WVHTqV7ikF4XU5sPSmjoOTHx/nuDXXH+
p106eyL6mfpa6YaNDZ5op6G+md+TysQMXVIDAf8nkT6CgYF11rjGrmMdifpob5fyHPx3+lt2R2sB
+yzCpJ0OvoSUylsFlv3eqclQY24eCuGENyeXXQ9OPnKfqT3KiPx+azhFhDwsrnOXGaKo8g6auZ2H
vd/a/JqOwSah2xv2A9pVRRT1YuOdFvf6CvQDU8FBcduSjutOiNzbzVBAwqYfTXZLg+CQCEzD+9U9
Q1d8LJ/RHZrNuMMERE9PuMBu4dV+HjwzcnlK9XwXKa1aK+zAipxiOjP/MKiJDqJAakB03OBu4C6g
zjodgoIjm4LFYQhIoBopZP4TQmFgNA1+Asrez9Bv+YLqrvyUs+HtabdTr7QszmQbLiTWut3GJQ54
Rk9o0N1Zsk46z6wE/AnTga4p7p9NDiR4aM08OxtixBHLT00hWxsvNOe7fBPI5DdCaZKcRnxqEVb3
mtvhRUZv6ZKGSSh1eP8DOgoc+1eOiwss4seSBAIW3ZuDIBUDCrYFA94qTp6Bj2j+zPyhk9D4O8qb
Sy6DM6hPXFQD5ZMOTuJNbdLAJNUa1tkj1zH1qtu64w7YjW6OcioO+tYUgHD90f9hXyEL98safixo
u4LTFSLz+WwF8DAmh7cCDdO8heBbfapjntnB6V6yswDhYmkyNdEVdlJkU0PldKXO378GUVXyhde8
6ST66bBUh8CGZWITnNMMzJf/xLYXfNHkF7qV80aH5TzbfG5ejIj058TdG+IZ4HVEOy+tei/TYfmg
WTDJNnaZr/ief+LbSvvRzjhMfXOger3eQBrvNrbm9SPJKSpvwFHiPoi1PDN+ekmIZ4mmHA+1FeYn
YxpISrQXcEwz8XC3iw1xYpcHJQOYAKLnBHk4z7PSO7CpJZYUF0Kxu8jJx0YABgwCzozFjJwJmn2h
MIvgMdDZTmCoNGmloaL0Xor02f4xcMjLkFi0C3dfIz5uFRU3nqmuVBgY54Jh4lQaX621Li0MZ4pd
c4AIFtE2vMS+MmPHmTvkjkpzP0t+EGwDivhuVuC/zd+YaZf+GaCDydMOzZipZAwTZRUklp3rvrVe
jSbmcr7PYPGeOuPcso84TpgY5uqLb9MhfXfmf8ujGVtD/FuUcs2+3KhepKgYyFnhukub0OPcuKpy
5K5CX+xsPyBDvwMUqAwnrzuS0MC0hrcYS0uiAHbMDKyEQeW6xEHGMEAF7MB+xzafXMqVNaVrmEmg
zHsze/FgYwaCMAk0f4i//p18OK/LqHiMtx91+mZ/09i4EXdEXV4g7z4tUSAS9hEChD1OnQKBg69f
DHz8cRsDO+SaDPsU+aCfQ6ptImvX56ewSomvJfOeGOpz/b6qeMKQb2p+gvjEZyJr28Mly9UUgcBE
DLMLjVuPHhnHmHj7AG5TBcPLHZ32XFKwOsbGYgGpOVRvSsQXBvEtShIS/zKkEWNwlWg7rrCXU8Fx
DBqpEAPWY4KsZAJJ/savIl9dBacrgtf9mIBRR7JzEbBvMWlhfzitHu+x2qfqJRJfEbSiAYbTx1yS
Ljm6Ro/GRsNBwdFN2+ScaSKUjAx4En1AyK+8EMy1gUMya59mUhyvVPrEnd7sDPqTzPpIb1X5Rxh0
VaQY0oU70oweEl++zhQ5eCOgV9LF5C70taXN7OpL07LulCg88LWCHGAXvmentb1qL1fAsBoGgCwD
jJ+VMo2/ht17OXecXP2Of7DXfWYQvA6IM79bLHJyZf1fUppMuHI/pi47HFaXX2fDna1Gyq+Rl68X
a/3gdAJMjTyF0gfjn2Vj/kcE55V/3soPW3hABeLV55JukdJYhc8AZgFYdTmCKbFGeYufsTEitp2P
gMv0Z+UxJzoNfev7qQiF00oekNer+mS+PJJBTteBd8iS1sjyLOhx582/D5tVeozm50aG+YvTOjdq
VZ7cLkabKQaNb0Zk55QkKkpFmbbY3pDjHyAsjzlrINvjAdjgzV0e0ppDQpMJZzyQB2XEM/Ixk9/A
OAATxFXoFzObng4H/7TNXjJqPH/f79zNwsnWOsuUHcGk4CUS3Z92uYDo57RCXUTXtSG27Qwzo1zV
F+cgIWhpFx6EEXRAjyDjefz6mQ96CSkGVqfv6D6M1ysq+BLzOFlwOJ1n3JIuTJUoG94MM8MRxUX4
j3+X0kLgg/jOdKQVjNWNx5hhoE8o4MoTP42o7ElbOEHUE+GfR9xt+n2Sjd0pf2Kk6Q4OTGKLP762
eVi6PI7t7pKwsZ25zOMjGUJyJa8Uha/A55NjB9JLiUkXLh7VJ9EDsCikJXjFtOaC+j1NqtAVK2NI
z0HbEZMV7Uj7XUHEhUOAzMLame6X/D/5NW9Yy/Fy9wPs1URloYEWnpqWqpSV4QCSEg03QkXZmPOk
3N5IDOMb+oK5fC8Se2KhrclHlgzUgO8ZxLdDb4H/xZQoFqp55tNei1Ky4PIS2m0JNLbEPbO2TNc2
Kb3jP0fhuIWqPevs0AT9BJYlUlsgxJB7u5XiE1WlOkHHCICbvracLL+L/K2iOj8kaHW2wnh0GdWS
aM8bg6E1FQOAZOPQp59a9gY3weidbOe3CBnfcEoPFlFulDtKipwB6t5SfJR4KLcozgUEuZcRyAHt
9SgJZcC12MUfBVX5CyOx87Fa7z7tALzr26kj0evJWP94kt/uxtl4VRAmN7E38Teu/OYHjuaId9My
9TH5sQkr1+WVK5n6huqo5Jq7fdpCBSPXHu1EnmP4bWHZpO2efh1yHmptDD529kesRYsndRIVb7Qq
q7DVE0ZvxTcMJ5UxD1QyLb4hC3KDQ8mvXcH+PQTFT6LkertKdGK4aaibv7nA0M5bUFwrhOKuri+x
yaSksq5mQEsPl3LNC26EURCZii3zh805brVWW8NvqLu34pRPGuNTZus3q/XzsMa1tCLy50TYrYAY
2gUPc/LHHmBb4GfVVAvaA/MHbzLIUKXtxle+WKVe+6hDU+oWbubvgiIHWy+tOo/ekq8yfFLxmznl
Yfj6ITCZ3EaRLq2yCTkYAIa9BickmLl4o3rNNjBBwlq+xrx7yz2n2ZkhB9VZSAD7FglSdATu2/1e
P6YHPAkV/Q3J4WaEtVf4tPnS96AVAncrtwTkbp+1/hlQkuU++5rxYRO3qGh22rJ5xAC0RCVju8tF
ILU3QLfSp10I4Ox0B1KGC66NHn27HyyuPIqrzzOW7epcN7jPHQid3NAEcQUEWQBhXNEdY9QUo0Qq
H2Ifp3VAPXj2lA7Zzc7ACr1iw1URA+bFSloJ+1CTsOEvGuEW7r1g5CtNCdEWXS21cn4eUmNH3IXe
fdjlPmQwb/NuSr+SNW6lOU+zulSDNW6n+S1uTpD/YHVSIiK/+10umnmComWWC24UyR4xU5RAUkbl
umNM8p3E9Ogo/W5RzA6pxQDnakakbx8HLlPFpv0PDBwyx/cN2FuVEAEvcyJo0nXomKvL6GUQcRuO
/AWyYr5dhrWVgAl0yhl4HsEnEISYm2TjTGkSxQXxuhKNvGifR9MYgcNrA3smzeH4VXWClgjEUapx
lrpx6Jn3Wn1vATo4hnMi6jiB60WMs05Xde6eA/9ZdHRwDxB9VnbKDjILHnUPlWRVr00Hs3j7m0t2
cp9udDU7rnfzPeFK4Ya6siFQt3dmyHIh3nRGzdiAR3HNWCLvMVaV+5MGb+YGAS4tBIUgMnf1sZNr
PIGboEp/dc67T9oeRcMYv1TFRyv+l3H8U65hhwVYhyKWUdjukcWhwgjvRw+iMHh2ofjcWcpxrptX
XqKdVHXirT4dDbM2pHZSw23I2h7JqY6bo9+hMSA7mB31U+9c0b0StQr5+CCSOfT+U1MkTPl/mLHx
2AaBkrhrYfR51k5OOLyH+OT7C7JezUhpmNcsnov4O4o1NdjrzMedPiay6E3/fH1dy9U9r+OWo7zd
YocwT12Ca6hcadHjgMw9JS6JeC1AJbPkoreMZnxKsN0kgGwL/iiaDBcc1ddQKYAae0MnxGsLmTKl
WpBFJP/E+Mg2bPNtcr6n/kyaPyo/DlapEAxOUh9md+iLrbKS1/tyYT1pxpXnIaTI6YiE8602tsUZ
LMpGOrfUVtjkNBR4/+2X5SIdnx/rGTmDH9K3kDGtZRtSshik9nYTUsaEvvMPUFh0WIYlf2jonCvw
T2aZ9zyIYXQPptHwhM9BREaTfvyYyzeDHwj2toh2i+i1saosrDW/2ZfujYhON55353ZRub6q7vi0
A70d0WSQnMyD+loAGub5Zq7k8E6q3dmrqbaAkZO3VWjQg3r06QRVGC1ntUKvdM1ZexwTTOhtsVAu
ZMXM73xaC8QBeNWAoF6IytFK4MkVPXb5PTlTSIqBMa/c+h4fBBCAVvBx2UUA0fk2mliGjQXw9Ig9
l6YEYq8urQCST0Kk2YtBgB+0y68thkhd9uoDpKMRX7JFVW4rqNqjC7XWVSPdEG3sASLjazqMMfkR
E4TsrCJMrXPd6CLrfPmHPiN8WdyLxj7f8Yx114ftxdx/Zk8QSDIYZZOcC/t12p8AmWa5E6X3zZeD
1K7pbYroH6Gr8r1/jkztCL4QV0ptWWr1BPSQiZlAN7VOvVEuaPB3GZ0YY1OXFv7ySOmdDfN7ZWiE
Op8HAyKugnSb/6awWKJhghvznerKr1PS1HmyeC42A405sh6CwGInR3ts/4fOwCdIpnRJroMmy/3y
xcr6aOoWVbhUEjDfyyoXeGnt0WAcEV7Um0O0AgwhFNEoU2STz2x+5yiv/dyFW2w6hcxiTvb8/qLR
LqB22ua6PC6hVH9M4qhN24Wipv1f5TOFVDK3dZ8mN4eJORkVxGGO2FMFfeBrWCHVIhnzwCePHLHH
zU6d2vgQajN1I102mX8PBRQ8U+nT0WCCjg51HxXm0jrNdqbpgAAD14GCo3OnLUhesaimXcpztlbP
bqayQHYXfmUJHSXkZsbpe4x3bm1w3aEY3ka7HaFvY5hSlmR6te3jKkSzh9UvdePM+YkgMk0chLCx
PBkZxd8uQsOpkkJLdVRx+krJJka2iStM1oVDLzknqbM3aoJG/mEArTqoIyHDexa+y9znE50IasUx
fJiN/kVWadQOlys3E+hs/ykEjiZPsZVf4UqJVqBqS3/DJuPTNazEyBdGy7NHpL1fvSF6LmZFKfa2
k1ojtgGwWHKuOK8wIoKlAsxmxpMWXoDMRfxzvYrBKWZeWqRc61b9+BwX2YARqyReU2tBdMBDhBfw
GZcsf++XKhJhY5mWFx0GjXtvNozzZaxoT0ngf//tV+wVCq0RE8ZmpMnXXcN4XkVYEHkNuuRTCeQp
eYW6k3SbBdBDOWI6Fra5qpfL31YgQu6LmRNSZp8Q10ozLJC/VfnLFewmdeCCyjeBZzC5beZHELVG
v3/ivF+w23TYAaONOP6XJOSdpEivf4Kbmc/fs7km+X5Dxqnt3ycEO+Cwt7LxIfP57JuvEd0M1Fxm
xFGbp9doEHdiJ1iVUY3Zy6iRGyOBhann8jBUuOoQTN/ZvsVbdxOmvfwcm5afHJ9GNWmtVjZ+qv2D
Syj6eD0PVQj1t8FW4EPzvqAJUEjEOdxyQNQY9qGG1zdlkJifWbJpiwJ7yfBXTqaazjxyfcxMnVkF
H0fog+cPnbEBTgt4seSn783qjjLIrkvNLYHDCiddamAzN5W+YcDrsASU2Wnr301irAwAsd5oNr7c
j9b9U95muzEEiC5s0IJ3d8zy5VMZpKueetr7Ws44+BO7kUqGBVA61FwbkEopQKG/7Rn1RzZOnEl6
LtzOAXFsdutnRRsaUG34g1Lli97Da6TT+cxG2e0qd1cb0aljm/oLM+xNAsPrGdI5qAFZKNE9hWpH
N4mAWrG7WDo/08oTrWmfLWD8jk4/IT3iuv33LnXvRBkDZKSRcT9aH9TuZrNlmppEOtCdL54/Pit5
oK35heyJAnCfM9DvlLVVYUzKXknNFK7kn1X1ZYFe4zpt4Oly+5GFWbMtGs/wXxOqDDM1J1N9siVA
ZJY2nmMpHCYepx+k+HfbiHH3hdz2LkefkHBgmk9QQVsm/LKFN3CdLtJ5zF+Ck/AxqN1gPRKMn5ob
tHXscY031Lqelc7keMA5+8j4HEbc3nJ1tpiicGZc++6arV1ZOUzyMbFkFE2H7Gw4SPsHGm7WAfn3
54qxaL4zR7dkyniq0rgp7FspXlPJ/AO5JupJ/43IEFcgktnHtCbMazYvxtLUyWpO4yEm+iY6XHvg
QyJXXAgh7+X1mwQXdS0ovSBuasaKQb8esY3XtlZKvB4tbaZEVpwG2WII+Rhb9tDTZy9rKGDL3tMz
16uFME32dPhvfdZGfq026G35pHYJrnIN9mFabaKvjtGHt7Cd1OjaSKUad2PxOowzR+YnUCDmiamz
pUseiMhfbr8bSlOSxdU2Vh36vDzuZbsDZ1PSFixIMOuuuPujj6MNnJlzxUeVzoYzk+1G0ts7FKyq
+I1g1yu1wZE6WLI0ms9mG41PM3XdXmy+pMf6TjlWZYs3phx2zHAQFpFfNdmaiBUduj02H5oB+sEf
XOjFGa++NXaWO9fM1cboJtQQ7VE0lqC6y08MliniA0uiaqytKOUP00afQv1AmgZxPPQl7KyqIt86
fN/J5AyKwAVDllVa0q2a9Pld+P+VeY5SHSNBGEg/LsEK/VumY1PdjGrtox1lW4DrJtmYL6MWXKdk
UDVhUQ1xms3upPv+/HxAY93IKPtlvUYOsRb9BcpRaF7h5oQ32R6MZ0cTO3LC4qlda8uq+uid6ykm
UMgqcwLz0KLb1O4QGzMwqru4B99ymIB6olq9sxdPB3NqvlotmSQoFWR8P6mconHP4g7ojulStNod
/1XMwVqmR8F6xjFfsIhhhyBx0TTcosL3P9lH0ApALRu1umN/N8HsKXKNKYTc84F6NJQwazHRo1T7
ydMyQW/8rDcIRTCAJaB7iOjg4/MUFjUSdVft3eX9P49fzmzYMCIrOqkhf531dej51wTU9x1adCjq
YObxwu4PnjZChL7RvK/AjspxPmw7dlD8Nf5qqMmpw9seDuJuI2LuxdnJLhML4eCFM7feUa1A6R7p
A/ue3A0Ythcw8WUAfCWPToaL9ZbibGJfIhGgs35GEopWrVtWqKC4lr70ri880FjmqrOgQNJGbdbT
8hVA/15/lvgmoTdipgIMMOAWZmjx4uFz10icmXlTOm/H73vkMyhtQGDTdQZUqvUGpC0nqCrr13mC
etQcr0HAa8PVQsiSaTvYxmtcoSIhSAw8aLCkjzxGtK5cK30Zs0KJ1zjFfR7tUxW89fx9a0lCzZ/7
ADA46scWqAcF/nDaG574Bfniczy5OjX45q5GPpxoFGS29E0bKZGJqSMR9pJ5YN1QAEeBQKJRUSp4
90ys6yWsHC/jGWMVpVsqptTphWLhXQYixS8AuR9AZEX2zrfnWRpKpDTQlpERpWzhKaZZqMw+aFbj
nc3i6I3ywNA/KPO7T7K4VfQ/6edq1O960shfNpMBC+cHv2sXd0G7ovqiFZpgzGjBV1yNsa//XmUf
Tu/Bd+3RRoUBjM+f+grCZP0K8PXiGao8crgbbysyP6oNGXqa2/7SrPIPo3acvopsy5KYkFK+OWYR
bxF9btZZuGKR7Tb1Z6nSXyiBF3ki9JXTyUSMhs3iTTULGhQPvZbgXBO/dmhloVfnqYGO7WYn2Nll
F5TGXHBlkrD+O9wvotWNmdMDt4eLddy9jNuFIWcs+qhNpDUDIAsSpHQ0cAXCJi9GMTYqyTZIsjz1
eJFZQ9TuLoIQTfeYCshEHD1V6hRqlvZ1lUcgciVQkNK1paoZuJuVzlOyxvtWEeF0gfL+lclQ3+Rt
LiPWUjj4Xe0z0OK29ImpzIbW1jpfiWYb5zyybBKjlYIo2EyJsDoC05+L11T02JJJB7qs1DnHWJNc
8uThKscUQ4XuNoUtQfhWGu8Wa5jRCaWtWM5vY8nBko+XI1aMTiloKlYEynydgLphB1+IOnMIbc1w
DMALnSBAFQ/UTjBW+0oh9h5TGxmCKzUTz99xybQA48KE0rAkELNwBO1WSN7IciZTWHOtljCO8yxN
m0VNlifO8a2oc0EJHgzsQxieumuwXOUTyeGx9XPESp8TE9yZIsWATFRoxe5HPCXCJbuoTf7+e924
Jy5h6EIQ4opACmkSu8HG8n7wrxky0lI81PoiTax1wNsx9eAPyxthO3u/2DQO6LmRhH5ceaTNX7fs
pbN1bOchIRaLlbPT6u8xffWLCdILkVAzyHhJo/smaC7aexdAoaYB5UWjHgxVcudCItEzWkYG1/Ms
pCBLSw6NQZDFAZzweZHm7ypuGN0bBgC8WYMNmcCnm044hYvZzPkBv7YhB9YKvrBZPxOKaU7g3HKi
PiqreAK1aVqoUv/PMpzUcHj7sMPnjtMEfV84FTRB2J6K48+091p4+EI9InVlY4ZAuegndRXEdNGr
mQ4WA9sIaYgjEBlW5rc9DkfqIVD8+cR1rrjzrRcoO79HmFG3S/mba+wCVb5NPDCvgI21seAde5d1
IJWunWiB/YNDseqGMDtJbg2YNSJTHtNTaqKYZgUlD748eDDHPjtA14JflQb8d/xvu3tuVTihOuNd
M8oWIX8o8OUxk7TJ+zoUjAGI7+yBRagCQgHa9MOMRMl2G1C/PXmID0a3rLHTtmx7DBngKek4uvdO
QpFM7DUB8nWbKe295mxlX/j+X02jKaIOZnSmlZBbHmhQadyQzZYhWOOTmHShHFq/O/xLDWtNsTKP
xudxLdMSQPIk27Tj/6zEwXLvc1peubmtgar+mw7C6ZHYPqwJ39Ft5g4esp8YqJRG0E56Wvn0RlI/
6x2Qd0psOt+ZHRmiAk5MlsnAV8pWiK824+kUeYA0WBbqbcOzRXhxLVC+PrB/dbZKc9uhmwisIGUY
lpvcTvNfl6s++mlZFDF40Tk9lTF5Rs7UpB5tncbvvrbPDkAf6css5kDYSdJimDwVBHUFjd83AlUS
HfLHnUjqhOQ3O9/zMQnPPGRZA9mg5rs5Wr9C3qugEnDLHYsNJU91ciw9EjFMy5EUy2QKfLBoqc/0
EmDFPoGh5JTstSQ9eRlEqCIWyfv1SnZhskJq/z/V6Rt3dpZoMxxX/Zcp1KJOPn0mRh0ZNtEWM14x
0lRwAyzVXKh6Fe2fW1ZoGIuY9wSjVw2CIJNH/d8h3AsboNLdSvRB8fiZQOYiROoeuIicvR1KkYA8
Zu+E+5wXHZdjza8mtM6mGFO8owBD3X07qXWD+QPs7CiSKaARnUz562zpI5bJ2rGliosBIFY9TiLz
e0iz3HnGQ0S5o4wTm32nATMomcKfYtlOOH9Azbl2EBtgbY36l0XbdRCamKPwgW3WurkYGNdNtLJt
z1nLPNoxTa1rM6Te5M52Frd9isnYZnwHOK0hCn7iGPWvdBxfhDBuYlBznjkTfbcB5pVT7N1erfRJ
x0wLo6ylk3FbvUTjuVTRd3Jvczq6M9x0gvsXcdvL568rnLvoCj6CS0jMpMHzea08DPnGoucjiOqg
T098Qy6pLKDN/fi7YFNmrE3+Ha6nyzcbDT/cBXm4YNHa9HYKD3lq7yZzt5Vzk76dyLS4RCDANbm9
NVJBQAwGf2cVsKPKqi4HUzxoYuAyK5+rW6B4tItHM7RRj097r3FR2fmi0KD3KgoL9VnXulWPCTYF
npWaXDD3GZehULFCFOQaDdG/4nEML7MbTGxM45yq0M1/j42TRcG0t/l9Fi/BG7uiWghuzb1+VTtq
fjHZ9t7niRSB8MnUbVOMLj/YtF3lrn6/jAYiMfac6ULwIfiArWFfu2huPOnfrR/kFv5SOsAazl+B
Fks3bkIDL4crLZ6SNX0D9mR6YWMDZgRPJtVy8sXKKR1UvnCoQKFjq4B7WHRqEsdDss/O5woiKDw5
LwKpy8FDfEDPIx9Syp0ZUfszvbMs39QpcrgJU29PmPQM2HYySmkwU/ZanG8vH2ZGWqCjCo1SCxIf
wrxpoLm1SyC9WKIbndmt9Gw63c51bE9md94UZ0OTVHAlvrnDvgfSA4JD0/DfC93MePTfyNhHMSFi
CulEzKh2Hb0npiPQOrCGH7dmCsduCK4CtgQxyQ5aDsKT68Rx4cIKTsXKnpUDWg7OpKH62XyUw4z2
UOK5RE5TIZ3JTMsujz2Guk/cFy3WlP6Xg65neXmu4M9rAmXk3/1Em2hq2NuRIQN66fTjOkX39NsM
hy6FSsrS0xwIy33JylaHsSI+wA/Wn6LaawPeYhOlBeBUlIbNxIm9EA53OjRRBqYNBpZdinxcOFe8
JhDAxQCP2VDuo2nCMzxg40Hpq9N3gevImJbtlA0/Kr3+Li3BYInY0tWccVVrBSATFnE6WHeUvJKO
l9zjl2eTnUzpwUqwHibJxbRYjOz3VMpgbgjyFbZ10xBh7bJ5L+tzwcCOm1WfpQM3v+GUo7rUJsY2
/siJQB4IfJ36jQSnAqKN9AvzA8L/3zn4Vvcs9ji2siVMAskWYhW62kK2+Il/0iWsdZsk8AnyzHV+
+QZX4Q2dxLe9lNef2KDicU0cMYGI9sajnAey4OIkpz6E1n5bynqy8WOVG5y4LzYF1KPO8jRoh2Nb
2yxD/YPLKwQ0ksHGS1eC1x68cotRzUB4YV8XpnOCccTLeOCsmkSiJPJx8yqj8fTvt7EiBcUmcCAU
rWbiResd7NfaLSaDNPT0jDUWcRIKqsBhtLFDoAoJrFLHpgVjdFub8Dp3FGm7xATyfcz54P+/5H8W
284p0lPwF8EKdKE0WxzRwWb8r2s1NPqNcjC5TfCUsDx0ieUhCmgLeXYgW9BXwmXBgzQF5w4b3tgJ
hkYfz5iO4ogTTSLy0snqUuyBcWItge8eTrLR+Nq5lDXBSLIjw1gGCR+OcQBNx03sbSJsdMnmA2+D
ws+QDINzq8J0G0vlMVLDtao/E6TIlLDqwCBNpCXa1BXRvHHuVo4IoGemXvXSjsbSSfkUV+zjzTmu
vQYzKx61lY2QqKyW29c5RS638HLD+MENo1idQf2iQJyCauvnwcVmQ99tljiC4ZgOTDibxdtdo8XC
+0BeUpNJjsW9ikn7iIuQ50OLzRy6U9pU0xtxDKN2vn5QmsXx25U+q5UO+nBMlE8YGSkKAukDkl18
7o+O7pQZw7ng0zUbaG8qJVdGfBKvUIcmg1OclfYnOAEiSCLJ2phnbRPfa95jmWaV7eFqFF9x4v9K
EoK7qGra2PqsZcqzUnFZ3iDETUubICMrc66S4S21HK7FMTFOHE1RvPl0Xz6nRCIA5Ly7fcsai+48
wHPF9yl7BTOXccWFh3objxHthPQYvEq07jt5Mg01jscp2GRxLp2IqGEwXp4uKyKwauGgMTXObiWS
T39q1CEysfb/YZbyFLw96vz85dlodl5e1gcR0/874qSgoVFjPUQcbkgzZ69KC038rM7/Lfbkt3u7
ksZinvZSB0fnAOcXrvpwleuEJiCuIAg4vg0LiRax37xqixebPl0WT1eyiH5B7O0WfP37IwCCgG8l
qP6urI2MwOuVwtMJ65SfYcA45H47BQOwTV3t9kQrxTjArt/LoJ33hkM0eXRZFsuPQg7ID0WbVlHC
joV75Aydr/2A090BcdeSqXtfVKDs9RpwRKV4lwkA8A34+eWH8EFu73zm0YGb6T7YwoOERmdCDFWT
cGSdS6hoX9vFHH9vkYK92fYmVmCMc7wq9egt726xPK4JelR5IsdbJD9i3JRHlNIfkJs9rmP9x/5M
4HU78XtFGQ/zByFSyJ+GHszW6aqyIzvQsXy5TxYvxm6EbTD8Pctzl5XdJdOdnaSP5V2yuXavhOhN
4GYM1pMXoX0YftXG8M6Y3j4axr7xO6tvdIbiqfaUA9XAjDamQRrII/ET6X3NOwMrge1sdPa7zQKF
ZzTy7NZn63s1Si+NWBvKM77w4cAH1PmFTbBwWV5joUf1Tx516x8gEaX5OguSw0rkTpB8gZz9BSu5
ylhrPyd9UneY37o5WfKPgHvJDdcPRt43JLL35pnKbfXIlYV3QKBGtTgtpUdpVVJsDyyGMGhdPt+I
sARogx++uqZ3F3XSV32G/1BPQ5pbdyezxBftxS63tLp18PprwEGDrOUoypHCBOURUIHBxXOYvCuF
gpDXWRK+/iO7pIB+Tlg+UDKlxYYry8RWw/NoAeH3KBgOBtZFhyFkbTCpune7rzc8gkSTCDWMr+Sl
s+swzwWSfmRRcJSswrLfvhBi8SAXoMEJFSW6tOLzf/VlmWP/8feHngua0fRZtq/n6b5eXohTwb6i
77jU9AyIyTG0+HAUU5ATduEXeEpu3bumhIw6WjOcXb65um1/xtsjStYi8rJyT4IPi/59I3LIsw/O
z4htV+desXrJu2JV8isKm+WhMC7LDgSWaAuIL/mkCEHmoVmxOdAKoFiJUdK8M1J6mZPhYUoK3z2Y
sXvNKGWzAFgqUA4mC8GNflhGVD4mlOX8pYAhtoQkLtPKG8E/vGLIZ+o7nZOKouJM9wQcNJ5qNNur
kzvBR8OmvYhD6bBRyjdue5iQLwS8JldpKLxVXLAferF4TA+WHMiog0BmdGml34N3tfbNZEEcdhFa
VfQ9GxQcgH0M5FoGc1rIgctC4+xhQX4XyWGPe9w4562TFLmalFmKRJXkzeQunGr5+oPu4z37T8lS
p4cPqJ3ZIyQt6UVqt85AeTgQSh7MKvzvv8X8dcRIFsHPKajSBfA1XuBK+CLT5RjIIatbQYKXqtVm
6o7aMVh2qk2dR/rlhx/qcRo1iuF9edSryUCbfOr4KSmyP7BP7wq0lA5gzkvjUdavqZPk8BC1XPxo
5jY/ya4dPdreUnzkvbj71CxJZvVl8GC2VkId82Mxqyn2id6qOMnl/2TaCzFlazfgLpsGTamTjWf4
X65zqFbs2P3eXqgW7UbBKNMPdMjfTrUfcz8lKETovcnqImehxbHRH4/mFoUvETHZfu8a4jEYCEQg
ZsV73om/h14I0nHs88yho4V1P9J8AzPIZ5w8JMRMhLnXaL5JjDtdg/WSbZ0FY0pv4eDFWoHr1Qdy
8aytQCED47lMBoxlqfsjse/YoULfvOMWrmSSdDkiIBrQLOvgt4xiJJU9yG/tp8xycwznWY3XKBOm
fB6kaQ9riA08j7afK/kTfgbUbYkSeK9dwNqPwysjNfgRcHCq965d2t4f8aD+DMgq7JWby2MUMu+B
wy6jNc+oPC1/1ZJFoaYI1CZDm3j2zxaWWm0lUGPBYl4uEu4YazoNDz2WyEoPgDc8vblQ6s/BFOr6
tLIZKIklYRF/bu11kfRPpM1ENezDF0SLCoW7IIiVFv75c5vEq8yg2u+tbekMgW7xL1OdP3iSOVTh
6E5dqlVtkFjFcWo6t4JOFxOqRFqqvAsL4PORT+iprLcuMDAlQe9YxMnx3iFrDqOs9/scqivuqCF/
L9SQmcDBlXhClQIlHtyAC3Rc3mzMUsFbCA2CAIEWAcBIsxezY4hqU7RvJiWNlfWCpjbOaytHtA1Z
cddvy7onlwN4/ejgk3xIgUvLYm/yEXDuql/m+XTsnhvQC7JEmm+Xqw58OJc5FJTi+gNUVoO6bIPb
FkTXQWZau2B4ORfiY6LcELCha0oCTCBClNwOCxHSCCn5E13FbxtHPYztRHiNASkHvLfCZA5QBPBx
/6OfSeEdcnXdOUWioD3DwdPKSh9G+ZV+6MULBGwWcMThm1LL94hR/uGyyWnCb1er9dIIIB21Tlio
tOZkuMwQWpN+iz065vONLlEylQF5K76G6HzsZWL9pXrsZfiT9drzKeCsQQ69ZwL8mT5Ii37JdVoX
LocFPE+QaMnFE2iO7/jSCRNfdrsBf2M8mnNFFEhuHw9myGWTJiUxisYhiyRgbJlorpXnt/mNrwZw
cDsFPrHYPaF0AtWVU/vpNqCamWMwm0NIMfxxw2pzBVxeypcnwGzzk+DN7DYlfNRYkETXWdKdeVxO
E2l/aoJucqpLMuIuX4uDkx2y0Z7sM+Z5PuIZZKD3t5Q8+I5y5TPM4ntu2YOL9VHtoXy6tskNbTrt
JB9wepyz4lEctJmKLbiH5X1o4V3gmTDiqG2XYSDUulvSfYbJ3Tm8or+RbOUDHsrFZW7Pan3e0wG8
vdV74uqiFMOk6K+7N0WFT5oP+ICRAnxPwmcmLH1U3o82I6Qlg5kD1dY3qPd/NZcTjTDUj84tAEfv
X60jTUiM5O9gA1Q2u2nvZt07lsNehh4JoW0+r5cXL68vWf5aJuHKfy+vzy+sRCGuJOcvnK0PwEj1
ihvMcFmwrUKkL8hdioTaLSUQoZSLAsSQVA5UStkDtXMRwl2uP8GOJs6CtthdHD1RMFAM2TnBbTOf
TWC3YzigRG4MBB+eiJq2e1ezxxnPEt2381KYzURnTgdFLeKfuvbc7MhPJSEyVbhEXQ+O1WZ06Wut
exj9uO3YUQEp/2MILLiNIFJC5qR7ij8frBVHf7ZhSWI5S+O4AeQT+ZPb3HVZ/pyIqtIpCdJRiEu4
GIS/UjxdC5h5LWSQ6eRvWjdWQkaZ8PH56gI0nVTFjwOtF6bu7u7qAWAD+08BT92GJjmOCpdV4d0I
Znxo9gvqTTVAChiSz8SOMdnFZ6y9TRYibnu/j370G0lnYBYmt30O79YVk+mU6wOv+B33CzK6f1EJ
ZTLjAdmmMwI2Av/4VtQRTqlLjWsNdw0ZuN67OBkolXZygMQ5zzwVlTMuthLO0hnMXJMzfXYOrEQl
UycEMWacuwlUn8sxfaPtR+3WrtB2mKJK+pimpArtceD4cCthtmu4ipGowb40odBBvo9nLlxN5tmB
E4AQV3+GBElEP6Mmmw8C92udlo3rHbr/Bb4axZq1luRPuaAPzmhbyrknB5ylNF2iCr/ShNI31tLf
peRyJfPcRFbqNA3IrZ7W2Iz4nsXs0tN/ZwTfRNPq8DbanwjO0EyxDxcUGf1aZO0SD5FWc6tgzmwj
5Q/GfNSLgFDXt0cHlag96DV+cezBSE0XlhAUokyF1bM2l0/3acX1tYp9nsofx483xxD4XeC3U+G5
NeotlidIyRVFvZ2GMtHiSlkVok85GHGC5uyYTTK740K+BCGAWd9/D09uZxZ5qZ91uI+huyveSyCu
WVyOS3wLhlPLZXdSffTplAqx8BC3qsqTJdCIk7Atw1Rblm8PviRZHs2GDS2LJIJzgWSSzzvBidY6
Wigc7xxxXhwV7p6nFHjySXMUjWhLdm9mn4AhQ+Ax71YH2lvHrNatjVkitaoWC3DkVJeblyjrIFrX
1Y3OiDEL8OJ3PBFdN+FdecJQ+KRjF10muX4mEqEmEwkTEHDhCn2KuXwdTdbHMEVOKsC1ojEhd/EF
7nmWHcjhTyQU4F8rFrI8jcUC0ewoC4IXTE4e8WfobymUW45TUw4vedrymS9SIrSZ+unRYHDWBqaF
0l3w8r2VzedYzQl+L5Vji1xr70eI1FfvvlE+gdBKEofsrHw7C+B59IZwbIvtN71+1KCzPK1KIYz3
LaelGpKhT+EDLKnBrANaTG9cxVPBtBIfo2TyOpnlXQxVG29YFoGMVHY6Oz1ERUKPHqnT1vYkgT33
QAwp4fv/tH2iwRAnlGFQXuYbkiwjIIQ7EAGIK9dF2mDqBkTXikZR+lRX722H00TDh6QtnwXg/+6M
y0RaJzJ1v44+a/tgSO4CaLsv7xdFRM2gDJRzD4M/tbtWixanKciH0CC/1od0Mfche5tT2bDOoZ9R
gopoht4Nn/kbvhbZZiDGkl+M4CjuqDXk52zbTBhSNdwaB+bFjmhccAlb1Of6i+BtgSz4pDc61Zv8
esulcyQkXS2XsU1Qk0yQFEunfFVsY5N3pSjlVc24HjbgGoLaLUj3NLYca6QuFQSVRloP1159ifpX
X/cEj7rRXWuTXIrjkQtXcz31KyjKW45gGpomwxNsoJbeNU/OVH+dABSyz3xBpCfcyhvzvG40Hsy6
xDmy5fsgDxnlZelLseL5fghkSKfY3Gceq/qvSdoEO/TWb6EHjCv+aplclWKGYMn6eiVRgqUvBk9B
obfYiaojY6t4F8JyRZwMQ6tqutRWNBnokaleKT7u0mUF+4X6Xt/wW+85PNX9IHPOgwgiYTsI5bt+
la/64Qi9ONRDcUPky4NmR7mArmGFygmUaY9H8Rz9bBnzHzR5Nu42naGLiMSoS7h9xwwl+mGDlbr+
bSJlZCVS1HA8o/yn0/UOLt5c8RUMaCghfnfwph8eyHJInlHx6lkJBO7fc4xnrNVUDBDYN6rH9u/Y
L43UH+IoNf11HUUSrjlRNy8PHynG6SHD00D722+vHtVOqAPbNhheT6AMuXMAo0kRFJis4Te0/6Ky
qsgUqSIUH4iIuqcjreuCweJlWR37evVOhXgA4zajiuz+lMkFAbUMGqLJU2bSX9XOl7JHvaZhcCQE
AcMSHDyw4p5GScPiUwrJoyF3nRm6IkxTOZJkEaB5FTsmx1dnm05xrTE0X/h+WHqus1flJFKA3RT0
OU8dp5fxvf3/hL/6YpjAuvgjyVHDKh7qtaBcB9H9DFT54HSSzMoRlaNIiqWAnByVIpINKABnWKom
RuN6sqq/rwmgTF2pREUotEcjJ3Y64CjdgAUOQb4ej4XpxRWW6rZIc38e303rzTQOnJLefhcfq/TA
csB8YJuZN39zJYkcHK3RIJLt+kfFF42f5mDBILXZrfN4hMYcKZRgSE2sClw3jD5PtruZWQMfLJpo
Y+mdTRjmsmFeG2FISkI0aEk4nZMoEK9MUvRRFIcEf5m+gKxzFnciaCB9jf8T02tQt0GAosUStbuS
46bhS+iHJC8mRDQLXlBPbpDfJ2r6+p4xApgZLvTuVVAFdtOC7WEXYrf7/G0r73PtqvobFY2ggiDh
2Yv0C0H+qvfYFozsSdfUYOxZN3375yCp6xeLEwdl2vylPuul+pe7a1Z4N0ULNYP+HafyZ8NI3aTA
dAu1gVy/yoU3+laYNjL15i1byo8MJAlRvS1blZYU2WWSwzQ9jxGrxNjOXhwTEl5bgHRBTCJo5ptW
iMzg+Yiim+5M+rZalVQHIp/8ZBu3mDIUQMsi8gZTe6sb6WtJHZyEf3JhW+jifee9O+XxCmI7ThJv
9XGAfWDA4tYeOTS5EWsIaU2d1srzHIr7jNfH7FnlGGE1WCST/tyk1EM+sLeDNZvgCasVgizvnzEd
pZYm034UrbZxIw/LUrD8BXbm3EK2HqLgQhkPyO2KWUKVCEABfffLlUb6GxVKE6ktnceQY/uSUale
/z6B9ZNSpY12pID+dDte6a74h8irYV7ZQHf2Q92UeHnbt+4QrApUoSEnsDnR3iSsZTHNDFgzf+M+
3ImjNoCpsRGuaHxPUZqhJeJdraZvoV+4qkmxCed4MhhH0h+mI+6FxjCqMVcOW8Ymm7C076USfcQz
T9/67baXuIhfqHrCbS/ojE12snEKl6bzhFIMzVU+Ah2A5K0t9UMw2s5T6EZttDCu9quHPeEZSspg
RhMrOUdwMpN1oSxbgOEAnrRGyWCeXiCdWkrjwwhCofHAUKLJRU8zi7CMAVcHbreNZYQW32G3K0gx
GfQFL4icRRjykiuOZYGeAD4KzaCN9HRI1LAdnauRvUBkzo53hGl2ydCUkFwPyqDrJZYSPvybf9xC
00m5GIaEbhNcNqumvIDq00TC86E0GF+Wj8Jj673I2MbiqqWA2JxO/LS09wYKxZHkWlUfyaG0vbTf
ObLGG5DzEYp85hS2Rt+fJo+26eFWWTPoc/rp16GudDfVB8K3ovpBgkoibCRDmThPrR/DpGd5TZfT
7QbRuZARCEPAnvqowrM1JFVM0bWq0VyOYbUjVuda6J2lQGIWdZV17fvJ4TG1xc1Pdaum2rL7JriZ
75Ym+fK/vB5tQOWVvbZGI+ofu9CtAMoEChQSW/lsO5U4mfdPZ/iMH5eQ5wgQ3N3FJYCbmCm5Ph65
OeL5v4rZtx0KSHr7Ye4AQaaejuAd7Hd/c1pYG/+j9+/2c4nOftL3BFgz9tUNFYtH5L/Wws3xIyej
1tqVuk4SMAWIw5WIKNs4CPcFNBu+vsrKzOtIO0bAtWlx7rlRmLh5j46hpnh5D+osPTwRbexC/naK
zDOUv8yhWn4h20nV24YPb2kZDmMeVrkt0I0ETn2qTzQcW4al+L+0/fqIgvOIL/GHXbCjEF0c9Ok5
kh8u73Psr8TRIq79bz+R6Y3tafxbFi4Do9vUug3nN9aGRzRx7bNVcVTPlR+HuqH6GM8qO4aE2rBv
EdlHb3H6zhbQWJkktkG4nhqq+oYGXd0ae1++EqL3v7Tn1f12Er8T3g4Yz2ZgnFh7mLUfCRza/g+2
MVrr6fDaYmWj855VAcmpEXurFPmryDbUzwIyd6c76/XZfPVzj4QT0J175gtPe/Evwi9lLNkTnGSU
UbLEWEmqG3lhqQ05SCQgArDEtSRXVMv0sa1QAHMsi7QjaqpiZZhAQePJ2xbilPVPeCee3yZTW5sb
xmx3G1J4vCR0Zy77EPG8d68cnlaU6l7/LIMRyYeUK+FeAF5UWfwhtT9LnVdCBmENgmWapoWUO5h6
vsqTkAbcCkXUAI9a8c7BVV+CwtP6Rva5R28wR8B6wf597NRKbVLRzEXgrAz6BSxwCbIzrPCI/Cit
C5zdmT3QdT5lklussjO9HetMFDeJ/foICyHE41vXEz8o4xiF2KnAPSzMpxn/3x+2apHkTPrIAdPw
/caV00fwLy7LHDF7rR3q+PGzHWBWbos/V+QOqaLsGLcJHAvQUmszVj09CU5X21/UVuxp29IEqhgB
jRtJ6l1vAp4wAoIIbK9wOH7TlJjbEjp98X+kqN7GmP2ylg9UU/hY9FTyi2OZgWCbyGtxaIbNYT2n
Vga7e67bsjtnRo2XzuhnO0ZdPVF34BtP7jAXI0uPeXumuXx7IebwxlUbkz4faju+rzbaqToaSxiT
vlYcnCSwpCUaB+vR+//cnSH5UBSpyymuDNWAfCCqcBwnw4v2Xhv0wt4COv+VoM8/AFE2mhQxk7pu
6wNBY6HdZ/gbPLVwJfpWuPuQ7sxTocWk6YReTUFj5hZbYN4ITZlliLE8A/zOtBRIb67ZcV4ivO+A
u4sa3ViQsTwOl9RMzFWPl665tL0QalVMGGBhoLqJ9K4L69fIvtHHogsRUEMQeRA+aDyBiAbmmiv5
LxFtGqnTODpEHSjzR31SLtIjYBVdfrLpAUdeZiYjugkJIK9YOBBxFeRAGx4sjIMihsRmaDD5fD9b
mrIH6O1MIf0TgntGyzfhklwL9gjUV8QBBxGo10Xtci4P3Y0MXzGvmXBrdYv+LYUfLGT79xOGrT2P
JD/NBuboq3XA0GjBUiVgMRBPt0SjsqsgCqpf1P851sOD9cK27tIbBtPOfFGsNwuXDIzYzmUvLj7e
HKW73tqE9L7J8vLiT1Zx1fl+ij4lOumUXr0kMVrzuJn2PbVs+4ly6hLu8L+2Oz+mHcIbAxZi60tA
lUUjqTDXDGJVOmtwBG3ZgvZ/nbLWW5zZyPBmAVsAyO8Ven0xpTK5rgrtWq/KNDNJb2pN5ztp5rZJ
FWGCLDCqFyHOGvAXZc/rk/3/7Uv2vZthXX1107tTW5TBToWpEInVAHbuGJKZH7YTbYlR03LrT1VC
iY/ybaNHPwlwkrFqjiqNhoO1wvMs93JZmX1B6oOj8laelwxEZ32V/cPEXXkNKev8SeOCTH36KIN5
1jp4xXtjt0Muyer+7OMnTteDzqRLh4Q2D0M++ZZkQsK2mNvx16d6BbwC8QNCwqyGoR2fWtn5RHSE
dS88WTznsPInpVLXhuSaGDZ0orzenFdluKS/rRxR3vV9IDgZ7q5NQmsBH50wFR84y4c6Wmso7Jb3
z8SRJ8fwLRkaGiuvgc+cNIRI1y803aYhukqUbUQcf4B5ep1d8SNvBjZvzW83/8anicINwzwktxHv
jrvwg1lsedQL4wuLcmAXtlNR8feJDO0uJBaxQo0ADnRmKWUqtY/UPSnCocJv5K9vBAJzmhthD9OJ
MuBB0JfPMaevyKv/+eidMzLHKsKoZaa6QM9jABtqAnjXeXVw9DYhS90UCPWGlLZI7pytHJoIbSpM
UktitGS2jjCImdGhncaQ32bTsM3pajDdHLwtO/F96veau3igpIDlOJyc4EFq2483vGpn99FMRUAB
hiB+J4EdJAqW281neuG5QHuUW33AeSwRCVYOD/oliCcLkpImeqDVN2DAnrtDF55vPo2tzEGZEdBL
mK1hWS3aUXAhZINmli2wFuTTLJuy3ahe/Krw0T4TiwQlNQ3tzC1XPelLkXjRdJNMVWK2xxvSdiSy
ZA0vYsKXXwafVPpYa9OH6tC4KbBRE/bg06d5cUTUQqiWkcN3f/8F/JwLzx7+j/IjhGT7OtahzEH6
rwX+vGvrdpttYQ3XRosReZ6AEa9aMQVBVfsHeOQ5hn9Cau8LmJBedWRhS5/QMOJjxjKU1x+jgpZU
6ZYhApcyPxxuK0LteNxDkFCGROC9jRtgmxdxVm5f6z4cBoQBGkSXlFK8Dq19155k3UNAx7KWLbUy
u0uuUzXCQr6UpN6IKAzt8q3tXbIhsnZ/Dw1PfMRcRARMQu0Ezdydt3h4QdHlZ3XHAppv06lcZEOl
tgmbWcktFubAuH/Y+JeIXtO7rkJDDIKiV/Z/bGZdbYqH8DA7/RzsdyBLk/sB1e+cjFMESUwex5R/
uBTdnkSscFsI1RUu3174+1T1luxEO7q6oTx6zzio45uznW1W1BA119PozxnY6la8okrWhr4hRJri
gk85e6iBBCsEc5UZ6n8MnBvu5zjMbRvLg60lh/S7InvkK0N8EgPTtNKbFTXe9C0Dyi1G+4QTobdN
NM4Is52o5veFMdLeQ1Jt1Yh8qxG8PpT/56x5gil8nCaZ5L0J+c3mP88/ARIod2FLfkyYfybCmxnS
BsRv0tMimATWU3AUByUJAo79wJQeJ/yFASAacfAW96MVSzczCBTHLQsVYLgv7sr1LjA2KLkmmuot
wSJfDIvalzV6CUrqsRLn+Gec8CjwgcQJLY0Cx1fRxSU7yqHQKltgzi8nsMEwQRSzmbEvbS84e1d6
xdxSmmesqNTlxomDvoB4Vi3IhLE5pJRdaj92pZdGY9sAt5gaxHKN7ZWUn5S/VMbDxuCd465AcrF8
2Ofcyq1Fs7/Xav4bMW6R6QdVn/2QQO/oNNTKz303N4fNwWIQFZJSSt1ByoW59OJlJ8VhPLbAy7fW
GlRbVl0NgPkkkB4ZKx+ZB5RIImSKzBEgXVRpesnSwneXKlsTyNHFoSc0bOFaRWRfoQYUurhA5LJA
vSmBISWrcCzoVzJoZ8jPgqYO4wRGNAikFmTkcRhSBhLBKlPa+ePV1kR+A7LnF86buXGJVcnDEStN
LOciK3zx/1lwM9gftpuRfJGiH7KzV199TtnFyM8kUHwX6HcFKHMM3467HIEtsp8bl7HGmbdDoJK8
C7I58PDUNO8FiGyovhbf4sDpKEci6/IxkQ3FASyI2TtvxWd8ypI4aWyP7YgJx2n52mD8ypzG5axh
5PTl4PBsls+ja2h0iKSq66A6tgyiR4kXf4omEHwzNVqtKg/aP4Smhiep+w9QnrTBhyeEIhVyvcmJ
PL97rrwFicXhVk2Bqe5oT8nw/0YBd3gpArsM9Uq0zK8Jks6Slm8HUOqMdsBhsD56i+2xn7hfGdXK
gfnB77fQCa8QtXrZHf9ieXpxATxKqAx3x4qM9fMfNHA4hVU8z80SU2Si4DkgAmXlwZDuY6RtN6rC
J1p+mBUJ8uzAC1mlKPLF7qM+2z/d2HzGylMqIsWTl381Ug118yhB4l77E5x+nz/E3idrOD6jwwuq
PzhiuxwCM/dgTxhQDPcXmDrKgSBPwP9ju6CjMNHVZu8DcQSxmTNjVLJkbFKbTVnwIuGcW+l85AxM
yS3Lqy5KKBjQ4JRzAhfOJccnOMdVLNCOC3lOq9ZVvYkY/cvOMf6CORPrruzrB/NWy5FfvDMAIsaj
Q2y8XlVi4qWCGjSV6y04z732+SYFiBD8t0K6N5gujPFDDjCDHJgch6DzNBPzd9XgBJKE7ze6gdfm
XaE/aExdsoU1+11pEvPk6yrsz6Q91cQO1ISb48gFoz9ltskoyxOim09sJ80Aun0p+tHBbW6FExYA
p5waVGLGcim0outRzDlJJNIwuyyMCBeLAtIXAF0VKFX+W1eIdmrrR7jgMfjjqMTs1ymqYe2lOHnk
NTzofV9L/WT6pU2zDgYL/BnlKBZtVrqxwg96apwb9nfGz4MNuTf/HvGh3ZDIZr7HxvIs06TEXXo3
LHCOgHsCB4G+1Uz4iX6CDSFi4hi6g+G8UyMeni+gUpwiW+gez8wBhkvccRDpLD/9JaNWR5X52uRr
w4DFu9VExnpNw1wRz+jB+mdYZMkdmVcv8rQFZJxzZ9qIUZBKd1MB0m+ZwJPTZYE7UaWQjZ814cuN
r+uJQh5ynQkJG/3sVGmVTjG7grkmfGS/wy/Xcqeh7gnx4nlgnvFlJKMZfwrxG0gwbQxHCD5kES/B
B1Q9Rz7jClgdJt5jfYG2iYzSFVvrBTBv2AAIv56MpsDIMNfufeskCCSooJdkrnIp0vON4FbfjZjL
MaiiymwWUFtVDnfVno2MKCEb5cGN/F0MHCfsEnD0DB+SFfVq4Na70QTuUFKJwYAE6D5CfWWfurqk
m1amgnnBUM3RBIAwnv6NnsjMmbWA37RcpLQPgj8Tji+Ykx2Kyjc9fyIPQcL1C3w0ylVXWD4X9Ux/
+k5Fqe+dCJrEJwE1ERWpw+MHoKrjl+ACH2Y23zJfixzp+1th1WlDHkI34AYcOiyz34UgeGpLRz6k
G+Dea4SgaosBLd78/LpAfnHR/If5LHHdRzxbzvM7PYojaqVwaWrF9MAKkSLP09I7Fm7AY354yLDp
NPfyFxdeeuymYKteRoJpiT1fSSqtknBJpgKxxm6tnjp940xqmZYFDZjdxPdpZfgE84sJRP2DQu/m
WJYeKwNp4JowUkhyP+FnLTFw7yZnjRKKUgxsw1Vje2esV7Udio730ou5ZtjsYOn270C+YE57FyKU
S+cmIvrk/RdXCINyX6PK9Ls802DxZgJdupIDtVTZBbkWYsfxK9sXEug2n0FaAhYugA4exqrVt897
L0nrnamAXWOTzAgQNFUPGDLahrOr4uW9P/l+dEW8gtTnjGu+sEsy4Zm7iIMklpWpNQ4fyB+HIwMq
SRvBCOAqApYkdvjG+egvajvS2GtfFZpHPSYJPWRjpXVm8nVw7jLtF8kWc8tst27dm4zty+PtMsMw
ViopoUIrus/VFtAPrATALTxlD72EDkx5F9F7PP3WA7bVaxkT9+NyuYpfACDelyXF9iLscNPgHuUC
1rpJ7eopHNUFXb2cL4QHiefavc3Vk5yshNcN8veIGxvm3hxneG55UA/VnQ6/kQVSjDatiXSipoN5
3eBCcyK4aW2GTQWzWjy3BjKmsKeIKN6zh6Z/oQohdZamD+2lrnp+NFPnrF58RZ82qlyMNgAM1jDp
YPt4HKcFO16yo51CpDl1gBLfHRWk3hi62kv5tUdzj8P7wCa+rxt7gV+IPICc69Yr9JsaZ84sIK3W
u71I0nEGIJms5P1v66zDvM8siGepF5ohKEEIWbfCPwDK2R8J2tQZx1ZFns7nboB7xqJrRc1hMSYV
Rm+6bo6CotuNBx46QpmI8cEGGd+t/pOCcTEzSeqD/z8Bq2dwfaPUG1HLphS/eZcO9SI7MVZw9UsI
dCm7Q0aF7qQBybbtnwvvTpse+Ur9WALzbV3KNMPz8JYl5jEu4TLNTWXTfcDZ0Fu3ioqRaD0wvhfv
5LRM2Fjc3dEr2cZC/inRw+SjXPYxKu/AeW+N8MxhefSN+y9Lf73Ffdeq3Ar1UvEyMh/cqib+qtHo
nmrju3kQldhOs+XV9TOlxf9qYKoPtC5TqTRZ3/FYcNAPt44vDFKrutJ2MTRZcV14WSh18hmHILH8
QsVQiWhl4ZrXPeI3g7sLULwMrJLZi6T4e/5Je850mFjCciVoNsJGuF6qaNy7REhQbYKWYsHYMx89
HoDaRZsjRB+9O/ny8vcaLHvpmk0zYA8j8znX1MFhRjlERox2lpK8+OWBlVVuJ2VLRBud0BHQuFrz
gBmDimSOjAMHaZLTgZo/nzGl5a93CdIk0yn9BNmWjtTjSDKXORXngVWu99xvMm9j/hzZD+poMSQ6
KDn+iYZpFQCYaTV1jMXSx0RpPhOpbJlvm0O5ABJLeYy+Jeo7c9VyEw0P54DizGTdy7DY3RPEc94R
DvNE/csyeb1uCEREYgVlosAkN9RzKnSTJK+kIuNZewXuZwVSYbbdC8aAVw4puU9fj8iS3i9nZDG5
60w5QSCFBsayfbwPrhdANw3LgnJVIgL9UmILrosggpkwiByuRwUJamYzaP+eAhPPT4mqMNgHvSnV
sS7F4v7LWGk/mWETj6jLgQRXxhY3KRF7aLxN1OlRYBE/HES4PV66jlSSERmgYe8Q/P25ObqdLS2d
zVGp5QFH4JytE1cE707VOxwo8cy+1rPtRteyeIsHlviSP3fRgCBOib+JugUqlnQrOt50cKFsdV/p
smcDOVjvOJQ78JvOKQwWdfB4JUtkoWAwPtaPSrQVRYdSe72HjfLXRNKmV3P4cbefenX6xNthyQlD
bvEsMLlgK8XBjzrBruopYjuc1pHzazNHEx7C5ZVKqeSjaEoXn4gHHP3feER9KZODl8htQC6AumI9
2Vt4+93ilF8AXnQ+sSEyuI+4SXiXqgDEJ4A34IQ6RRAALEJe1p5X1VBQo4pyLORiQr0+iWN6J56U
m3f7lgLnHw1yuFQX2xxblb12r7xolLCn/saXVDin2z41Tu3cigYOMnI8SmNWKCsEDkZ/t9jvwegO
ZxY/kNgMLfzBftjJd5BdVje9xjbzMJzvE8tg9WJkZVCCfKrH+SffWpUmaISaqQSMJ9wt6EeINMDd
KoEHFt8Qc0wTTlYNC5NsODRVL0WN/2veLuOryAaGCpy9Spd5N2zEb9FVo7GJgNlIexgaXLtYyJwZ
wA1k7RG+OpgqyqVkz3XsMGhlBYjJ2UZf3EF2lwOy8WPbY4kNXCLH3NBK+FZ1KM8UX7W8q+CwMWiB
lQhGDI3zn814ELWH+Qs04c56ERrf5mBHMl+KP5M5evjmiq90CQjcXFLjYbrG6xq/PVFBm82DcnMI
paVr3Iw65D5quoM5+5dOom9EoLCRhOvK+oh66RoZ9jPUE3ND2GYM9jcgZkkr7jkB/WnqH81B40yI
TVh6F+xLnXHT4bkQdSZaD2Cdt5s65zLnKOfkXQm2H+1uUThLCq1UC1qZ9k4tuQTMSuuONvBdB2UU
jrF8URkh7vmuwQmTkRWh6gjI8aF1i1N1kchcvnJS1upBlA5rlqwG0a9lPNOQfvJvFlY8EY2DybUq
dYqeMgHScnTXTmDREGZ86Xij9nX06hS7mZgAQng7s6zLOC/wEmX2TVeE6HQgqHC1bWTqBW5/iSTE
17yHMwTaIQ88ToHCRIO9IU7MtgXvQcTO43Ju6+ugaofTxnINi8Ny29+kjFpU/lt2jb7xG+RrKyDn
ZxtT2h0swoa4rwkqLPDjeGAsM8F/dzz1+uUU8BYF52i0QVafonsWVF1TKNPDFLkr2baLF+NLTMLP
X2l/NzpMCpsYTFD2QnxSShbGVu2XL7QKXOAjfx1vJ+A560qT+2h14xtAhcBH8gZREqcuZIDhDi12
GeIJrorEojUrfmcjS6SQAjJxUR/szJ9oj5bhR3wgDeRCp+Jml9dd9U2U3dNrCoqgwwDzu5igYo4R
27sSmEkMCymVh+LXJ+/mkhRhyCXh3aAYPjwDqxXOQpiLO03uzFcb8kf2C0E+Jvz5NagPlkoTaUCc
XWpE8Bk6thtLnhn5VrMDTEobrmMarRY85r0BxmEpcgX/gUljXQ3AOQH+isVoSwaaNb4cJDnrc12k
Gl/mgSOLHoUMq4cn+NBOjLE/ZBLias4M6ijNknW7yJ10utIvhcfspUzioXzI1Gx0FObEWM+1spCd
nF01zJgi5BeG6kYU8yKJDcyHJWB7xhSfqhawJnAFLbP1RWa5SxRIrGC22JSYdLk6NMyRTR3AesW1
CGjOAeoK4k+2/i/ftaYNoO4MB01UYGb9IuAw0yBKOGXr0+dKUWm/RZ5aTiAcLBKNJR9tH2TwWfrr
aEew+WsUje3KPRvUCYPD8j3hEWP9Uw1AZ86YtFQP4HoyKSoYja8DXKz6S7tyGZmZkSQLpF6ZuVjo
2vx3DTOMpnBuebMByV8/VNFSZP/IlSQqDwRqp/NZiztquiy6If8f7At7gdv44QmSgFqyWGrEi+8u
AX145vkk8QP6RQ9jmonIPm7noPk0LKd7djrulzoYUrMWLd9aUQgynZd1oWtuB1NDOKqUhTsA6C1u
pIcVOItzx0NNdlz6lFZOFXvm2DYeSBJG+2Rm019B0iQNWDJE291DxZDjOrwpwpKGYGZj+QAOi0H0
PCcuD0jWGFfMGH3CNj74+on0egxX59h+apTHmesv3385Z1T2mUIQrWbjQDiTDGun3DRNg6T/rvVP
xwDFrHlFd94wgoiZcufQEVlQvOTDi/euXwiST287WQTdiGwMTaPLPtfQkjYBxm239MP04bHf4TVx
Eg2/UboB8bidh+tposMotR1TTo7vINuqIr95nizEI9STpUIqeDp/jkmUCRwLci801JiCRM/yhr2G
zIlh5cl5S7atcysn21+WuAnZnkQ1MClXiTWiVDqApnNgJWv+Q24vENjK+rFLiA+qpqBuRxxLPcdJ
h7++ojuPuONIC/Qfpr2fUPqzd16xS5KYKK9Ui83pVjV+Wd5WrmGxkRgw+FndGLr6qc0Fl/iMCfmF
Kt2fb+K6o3ja7cjtM8+JCNXw4KsjmvrL/4fZOpIvPxa+ZxXvF4t0si4i/FsQWMDgepp3Xzz4A2P/
YgCt+6si37xcbZ2WN9hZo87pi1VTyi8SYUfdM/GnuDkAYifIah4GryXx3paeqXaixFv9HcJek8Xf
GA4VH1A0jEYdaGgjv2dhWeuehwQUouRJJ1Vlzov6rQQOlb5MR5CtO39tYFym+X7VZ0HadLrU//aS
nVzp5X5qazV/Bm4ZCWtJ3dFdMt6quDB3GOms3sqOI3q6kUrCpQ6xgd6ku02Wv1P/zhpEY9sdrqti
ZI7BfW689+xa8v02XMspp1OD5ZPTrB4cLphSwSXdiFBDKDNiimwtw39EmeHIdafE4kx23/ncSASk
Gf7VhBqykrWqxuELD6k5Py3UjB56LJ45eCKxcjXrnw63jww/Xx/mDt6VnM6pum1VTke/zwQo2FGx
OBqdAnskmPM1yGdBtY1OlJ/bdyCqHdOIwi2X2PkY1yVk6AlpYwQuWnqMOITzEr5OjVBS1oC8QNkx
dLAQb6BzSaZdUKZA/qiOoQM5KhHZ0fzb5AEmy40vYAuVVwzjLzjG/UVzMaQOTEpDfliSflmy9xTT
OWm/Sg1GBaBHwGKuxUs5n2TaQnW6PC5FLspr2IKGjScqJhxc9/1C4N7+Kwqt6n/gZ5dULGvjS/oo
2esTXnoaZCVfUN/WP122XX0W8864gkmTKYuKGkw2OSTM7+Colqk5xyAoIU/EYG/pbVG/o3JPVqa7
FiL/YLmXxgLJ99/klzdWhJ7SRaRldvYmI4YombLqapXBT0rw4ZfNSVVWfHQ0BF59/IFJvp2lhGfK
HVbBQPtSdx75S25qxYsjoE6WkSMewZcsnPu0B/e4XHkZPL+lgay2Fj0/IK8HZetsBVOg55gZb8sD
KlHofZ8/mamOx9MBhHT0EKSJcg7rRtaACtSigp99n3aJjgdTqPaeu50KivK37hGwLK4oPLeYeiSP
gWKePuS64esofT80ZU/xhc1iR1VeZeLQktqjL8kYjWQVXQV2h95IRMPRIcQ1ucStDo9mM4RSTjHZ
AhGWkE5e+9+0n6O1NjRj2ORWk9mdBzXLx/Gmn0x0aeXeqUfQDhKk8LMoM6vATUYlP4mT44QaFbri
e3ydf5lzzFVi2SurN/S6kuPXvsw0BvstgYLwjIcs/oHEGMDUH51Tbx4wDLgZm7Ew5Tg8jVhTCiIb
VYAfz9NFkfFJmflOkc6/mLUvCyEGlWGZtZqLtvmCRXRBA2GbIkw/WnhndCK4c45890b1rhFEBisw
q+N4hGEJH6h4J8mHLa4PC/Wv/ocuCiWbEOIEsRlojQj6nTxf+k1Rvd9QYMd3enmCNDdPUxDouwM0
OCACY+hYX9NQw2hvDOnsmMt0zIgBLqB2IkZqwzllFQ8Mi6zPE3+6jWWoVd0BENUJUKD0h1UHVnK9
U13ujrkyABM56GSY58GtDe+AkLVsIjLLrGuQ/hWqJfGJ596SrEDqKcmslhZeK4gDoZSUVZ6pS8Gl
2phvuHGaqSDHkHQcmdAwckMbSGQHMEM/fl1hxHjUGDqP5xPG24X8bit7aCD8p5DTlw4rJhARgjMl
iTvTxemmPx7eSHHxhlAt06rmKeg2JkfL+KptnhsCMcbtYDoWbiZ+nwGiaO4hlIF8ptJLeaZgQ3Wm
7Hx4t1CP+W0eEZImpz5Jl9OoGM4v8tz1wxLzv5e9J9wvvQ+mTYFQn19OlUXe9/909T5Nn2e66wuh
gaMMizBxFjmBaWFHZd8A2985ydqVq67ZFd+4JNoiJ7+hKjk4dkkTsEcVf6CCZBl97te/5cqvVJth
hz+72sood+Gkj5g2AMub13Jbg5FwoluJUbO7s1cvO3p/zXqYH8TNjOlN7Tza3WMnEjeTSAPhMPJn
RYVrjtXPd6yAfeF0ynw6TOmUFCp2P2h1Q7sblNGnWZeqaVWhKQCNcxdp3PPc40yAWFHBMjzhvEdN
9AmtnJXj895CF6KnP/kbwC7hmCNC3ZzmPPfWGqa7QBigPmYI6z4NfNI+7nk6Kmqyq0FJSid09rw0
lpBy+RhtSAROP41LtzfTUvS2573+aT8sZ5Oss5kNR4a5ocTOQ3MAFMxU/2qZFGxuLOYjQqfcEwUL
KdJQpqyqrNAMoqnx1K2OYpVxsfl6IIvzUdipWAhmb8bHV79urOrWAHPBiafN+VvbYibfKebi9Xsq
2n2KnpknTHQxAnwTuLcctbkXIpRpUgLJrDubRYO5dmTMB33F8lu5A0yoC5cPzZLR1M0JhUGBpmbd
HLpLgEVdkvyT24Gpsu4CDP6tzot0MFJyK8DVy32NIn7CdyHcAdz+ZBGu5voImug1TsJkCltf2nbh
YWwinsisS7cdf+kc97D/88n7YRgIEyH+olkzwroQ9nxPoifITu44r1pb4UL7AqnvbH731+AcCSVE
yoncA1UHxJ6t7AKeddJujjdZou+7MqTHshYnfKalWMsTGs7BoM/D3pl66kov/WHB1gE8T4RTl+/I
1YRNSo6+vo5PuC8V2HJglUZrtGxRSiei4csvONUb05n1yGmUDvsBJVUn5iYxZEpEknE6THRyw75D
bO+jtlIGzZ9o/c6DAmv9ohaYZvofw4b27sr69eV8RzB31htkNWuJk1O1K/cv580oubh7mrJTMMXz
/Bk/4iZe6I7II9qUN3ixGvmkpLFjdy1oVOgDPRom4JMdMkityaLFaeHirBGiJ9GjWDtWuMeG9ol3
3Ypxb4zP1PoRgflQ9rXnVf4d1+EKTzcnAf4uTGzBjYoF9uPEgoMKBP9ZMV+b9tnKfcXnDqjvbZHO
khxM2OcBB/lEJWBSMb/eJZOGi2EWp4nYWxr1bQ4QpWDH9V5HT0L2gZyheSWk8urBoCFNPdIylqHq
RJ86KN6LVNZ+kAylvDZ5DS1c4OOd4tcO3wH9PAZVxodHNPsQoAJgh0h9y5/6PPfSUrkKI5QFtecF
Sj01+VrEdQyJIYpdhHLYv46+4PFdayJdy49P1PrqD0yk+gKiztpJ6cI2WrD0FPLzGx1/RbcUHCsN
NoCuq1RiOZJwLaYY5mUp2UvmHoKHcEElJIBCkZLL7aWvdVCLmC0lOjTiwxzDFMrFTd/eJQ5aT+97
2Dx5HvIVwlxp2HUdigOG/U4nxxVdKtCW0oGkytdXpkseaqFCcF5qA93qYU8DK54q3IT4CeVQL8Qn
gQzNFpCmhHzRb4FywGqaL94uBFohP+KUSsmEQ/M1/hUaWXCeHiWgJeHkgwn11TB9uFbhLrqc3yXr
Z5ecdsnpoHfsmD8YABfLeuqLzasWNtVooZeJBN8k/Garl2WP/1KHxDktTdSrdSoZRCWxADohhyo7
kfJ2bxcrvVVbovIaCnF0SofjmjpEkftwFyC/6ZjlMs7WHjzu3NC5hCltihqaERnS2C5HICO7Tfmy
kZh/zDn1hoEh23UuxmjRcbCaba3+j4Ib5u0WVTIj9PSDCDdwN4tNd6t4JQTnLHdbJUsK0Uza+vQT
J2dZTn1wHNhEVhkl5Pbn8yJMg2R+rh0FoaPkXBd/k4Ds4sDV2a1eiuvDKlboRVyNpF/mNAcRYk8I
2QFrSGogNZJUTCZ/JwwWacEgHmxS3kD0DSlhPgrww9SQx8o9c9spsU3gTjY2nY1JfpPa2Fklo0uv
W/gNMqeNXhwhuwIS/nHcHAzhouPdIS2i+U6i1p0nZ+xIunbx7bfN5BH+mPV1zf7Zba5FL3OVg9Fs
5BhUZ9Vk1O46MJkuwSsRusao1Z6jPlyWX77wuQqCMgU0SttAG+C9fvx4U/zsBOvOgtq36z4QmWRO
o17d/m/zzoO4mgm042xXyQ1y1PLgr8gA42NE2P5MlybqhYBc8T3p7GsD4rB5kWyPr2FHMSZMuVkM
1yc9oRp/3Y21eA4mgRtLDlsCWKtPAcRVx6SENB3nCujKwKsRU8J/+jUMmJx2yPSOTnjTkbOyVEGW
twlZ1GSVIXBuRz3nnj8VswaeUTFs4ZDE1D9fOZLTMrzCTqvP4ztwuwAdJoOkktClX+I1I5WDsm4x
ECF/GLXXe+R0dyBqaAEwJdYhq49y9aHDQWqmUXPr/RaCfmFx8QsDGWkZ4lJZQpiJ97F+5S8XQ5r4
XhlUKUQtvSXpr1157BuKOHiYChk+2bJLjTCg1itZ2tP0zf+qlWY9i5NjZBzg1OpZ8Q2rPu2sPyyX
T57pP8MS4+8VKiwI4I1NJWV003LbGp/1CY0wjf7ToUa0s0f2Nv1LF6bvGatPPu9GQ/ZiNfUDgT+U
8qbkgOAEjAypR+RxE93i/IJfO2QOMR8k9s6D0T4EYaIE6bsPNq60GRZdOOlSmW/SSiqzB6CyajYl
QRM5/60H3de2rIjCjrCeNg7NSy4qZKAFpYixHvRFNKWR5R+SIrqctcIGLJZviEdHy7xfx5iFE3/t
VesS2IcloTD9vsSLdpH24CHM3mR3+rocltbFtYut7eBAUToSPKuqTJ9FhhTt0mm7ZY063JODmHdT
H0Hywajk6wz1K49+4Ve3+XEaDv0W6Aa0GQ4zZpJ7LVl74dJSEsEwYko6lVvB/hbEz1ru+hMf4gwd
JdVbVfe8kdi2PuR3idB5Eai5zkRht3eXzRR59906zaT2ztzATZMC8u3xqIv0TE5m5zevMk8o9ycw
CJIszCkiC2eu0cWr+EL8Cq3x39Lz2sxJQyf3wsk88X/3Jfa4RhvM4ypoJ56MHpUtrl3WxJJR+JdO
BFYAzYfjxpG/1xgTJog3sGtqYym1FyGlJr/4YVhYSHf1VAUqi0DnI1PdY4ANRo8uWp1nr897fwii
q9fwb15fXYEG5R14fDe7bgaUMYIw9Fklg+Ck4r3qaaCKY5Vd6pDNVajqwPj8UbIBoAfxN/RIQDSJ
SjF6GrNlFxv6YlXFVfS6ydyVxjorEpG0lrChq3vWy6sxK9xGxkdNzhmdZ4XNnk6K0r/V41V0Pgc3
8ZhmSvYmIQTKgHCYq+jBQ+rL0jYW4+nOmaNvHlfWBguz6mY7DvtPD4oyd6Z/eTRRORkX8FOCjZJ0
ZGEbMju2rk9PRcVnJiiE2pyRLV4yMTJWhE5GAjo12fTCJdaWREAeAJHchuqQXN6pmtvS0Pv2sfTx
sDu3/uiZyOuqoQljHv4MFWpz8RHCH/XDnjPkGXPesl8rtpjOkehixCyF9qBv8D7EWd1VuHCnaroL
0SXhtRiifPGjAXJ1WT+/c1xnOt4NmK8l1E9rKi6bCbFFxo6exPRAPlN+KNCcBT7kYZT8u87cPkdE
E15vEOATPFeMPOz4T11INNqgUns4O9WHWvIrNnUpC81NjLtUcaUwxVQcXSVkpUhUjWsUedXu8CpU
0Xnw5uqdAsO4KttjLL3UTsDiNVAZ2gHoFARUlpy7Gsqjaw8e/6kczgvC/oGogFlibl2d2EIMcxfG
nSkGfopzLd16+pAg7tK3XMjlT155t9ys2K9aDlMqXmKF2rKUo2IAbYdHIng+A1RA0/gAgUFarehq
AaJ36bx0C0231ZQb4jnRe6oft35Z9DqfoBDqeZ2DD0K5+3M4D9nn5v6GuVS1qAFuXKbBPFPitx23
DjOJlQgO6IXFcDMAzL6wPoKNVme0ob5wnf+118JFS0X9JT65ukLkWrgxTzQUzjFDdKndX7a+Opyt
Vk0eBxiTXSH+ok82n4rrgwmDQz1JPW2kqh7mXZlDG5TeKre9QIDr3a5gttC4ujf9MbZCx0VWeyeU
ED81joIkwuPhJQOY5qc3F6xDbiXSmeeS1QGJ+4+qA+nBf4Yh9gDV1h7UFQXt/nkAafUbe9FhRO7y
4WXU8ORvB8RJIm+RZNxDL6NgxsaK7t+rPEeNQAJrEHYkspYs4ZtclOLLj0fAABfpzgQYlGKSZGaD
jMIyvDWKqQ2Wpigm3BAIu7O+Fin4mV9Sra1J8o+zAkIXtgLCvw6nnQaCKXHG36M/vh6E+FOa/McN
8Z0DfMl7VRZUvA0/k6cCWV3/BTrsND9r4Yq6LZdDudDuHvDy/5T2ZpotZ0ppay4s9UqsyXPgUr3x
Cn2TFz3/SVraTcLcb+7RQDbN9ea2DVc9JlOxA+wuUAUIMSRU8siowvGwbI+7kUB2YV1TysyAqT0w
F3edanUy/XnjgXds7oQXHE7/yQ1bvrJEPungUmcQFYNF6tCbE64VNT+aZiX5+2ObRKtbhThZAgAP
A9GwN3J4yD5OjfY1GO38qUJP5M8Gq/cxw2DVqolvqn7tVkV2PFBZDlFw+0lHYDLsScmgNtqqFXU+
GD6Oo/VaOYpF294EzHC8Gb/AxNFnpu1NctlU+eNI77j6VIJIqHyx+tRd9nLqTon/WUHuAVUM/+1q
eF55Zq2hP0JZ39SOpjU9CkCC/Ky7xEGTyyXYce2hXHb6GY4FnVYckBD3O0wZrvQkZ45CGuCuYq/l
IR6vn51rS+Aq1yMTlh/2Dlm1XTf86DzAFttpWWd5om0NjV3U74goWelCJRuAUTxYWnAdnRxCWmEg
gLtoHGEaOC+Xy7ekPAcOkLFMe6HYdIK3LLkdytun0SaIHqhIV9It+wl0gqPN5cnB6cpElnD+thdY
kOyxLAt6dxk+fiqLBJbHHBs9I6nXVE4iuea6kMAtT1KGAibgdmsnSAo8chI8SdS7kURqJUW0/Fet
CiY4pIM/8lgmsM5caVifer6el+YMN+cEjKH00ZO+rMZXIMUHlJOrHuCo9mNPZYep337HJDak6083
fU8mtM0ZsPrlYsHD7+KYpBM9QKdDB4i0ACz5ds4vH7kh0N6tHXxOivXNPyhKQCw967KZxuUpG5uv
UvpiZaeGmWMgKOqdDbV/N0aIQc8uXzIg9cf1mU/2/KvB4wWGbrWbBvJ3JM7/Hy6tm0tQUekHuoq4
+fWBlODMNf3IlpuBFUVxbzM2b0wu2kwMBndyxKkp913XDL9agC7z2+IJXgjJLQHD2mlpeVQqvlgN
zVROmOgr2PcIvAGT6HyhBKmLSmsY7yLMJ0TLePy79uFOBjxIMS7Wgyn5pzloeX+AtfhwaxoVbWnj
kkmTM8UTbpcACP/bTeBqqlcfg4DyE/wX+3kdSDdG8+6CoWAf4pTrlKVkKe9WEnc8D/wRy0cvJ9TT
lxl253mbiTYCTlhkS9OrvLQkObRB5kUgOsRnJPmo1GT5djBqP6UTz78MKoe4aBM5zM+xaCbo9C3S
w7tzK2LrXLV27TNKp6K9uwmTgSBAmgQEfoLWnE+yciVXpQpLT3aLDKwfzCSBitQxQulFQ8UD6cpl
BgGCe2FY5Gm4w29GMo3hrrpI956+hNdcc2KTYtzGOO53kgPrWl1BHm1qbb73xqXeHs6MM6gOAzWO
xLjrryhuFA0P6PdNKTm2SG6Jq6TxqvrYZeX2WgHFZh9uG5ngWteUl0y9GCGZbJclQmpmFYcCtWOn
4SNBKSWIlii8opMmR5V945cYwjV3aAylBd9NPjIEk5qmoiqOQrNCCJvm3vE1q6xaSu4vGmQeiXFz
JZTNFE7gfJHoaVUFQ9Ps7Ssr3X1nku1kJv5xJ6R4xixXOIURaKbUjK800Z0+Vo72+Tl77lFmPDlh
HlFD/yaAskGeQKHwfNy2lGoj7rMuqUGfnJyp3id7lzD0j0Fslng/Klr8/hrnWTOeZgEBV7NxoFPF
QkHlKYlx1y6o9THbNhZ0ePEWUTAGtpc3FBjKLUvd4pfnA0F+aGssK8dfip1mcFELL6ZflAuePVTO
0pmsG0vIlVuQv/hww+kKzGvU4PVJNhSdPg6Df5Wj60mFSyg150z8iPAkBT8UFB0s4QMLqTOJX7sB
uFX5vXVdNq7sxdBeRFd2wcKFl4wRqURP8dTCL770mPgr8qHmE40FTnJMWWRjqu5UpladrqBT9wIl
6NFgT6C/DwybH0eKGAQxU3bB2hl7UKUtGb2dVF4kWK0GFoKNVsBeiTl10M6Mec0CSSK3BpB8t10v
YeMswVWwz1jVwYi1OSMK1iFC+Hwg4p7DVi7YC56NB8mz1CBZCYuOO5sWQF4EmB2wCgiNDsIsBb/j
G1jbWgPdPW8BJ1vms29V8grbyHLtP+CArywWJaPDsWOQ4TBm8Foc5ye7H7hT8vrjhgpkfNELlXd/
XtZGLkCNKZUx74AHkxqJPdLvQ1kF3agAnPP5894CoYlZ0t8j/nfrkPCtlVBUu1jahrtR1XZgh4xL
ziOeDepeToZX0Z3FtIN2eGmoChydocDLVauWZj2SjHStHg73v3Ap7Mebx/f4WpHudI9gTvrfiRxT
tZRDBnZIpsE81dedrxcCP9Yd+A51TRV1YF552QqWyuScBVuKKK2/xnKn8bpeHP7otQ/tBSC3ePC6
MWW8CLdftT3U1o/Pt93Hf9vVmbmzpTuvJU1eYOP7zhK2pdP9SkHwj5MuCYCt9/jOXpK5hILmNova
1BHYMCRIVBQXjErxkcEBu8+qAShddq08JOZtGdz/Vo3vhm6+nDsFrqXZnPTYvJyhHX3W/tcIhBEL
xnk1cbaHvQ33tx98LMi5WctAzryLshZK5C2wl36c88v8NCCSHE1nCZGlibQAD68Sgt7a+fGmE7+G
ZV+bCxH3TgIY/Qsi81up0zs6BEAouMR66yMID3sH7gs0pNF8p9rJqKTkufhs8cW98YVfxXnjD0jF
o6LaL7yUoni1G3is02dPOAmL8aTGjD3nkY2/3KvPA/+3tXV/VfNcBolPRBeUc26cduInnYT/nWQV
kfLj8UhreCVXwFGVM21nAf3s39JtoPSW06gouUY4UYjix37iq7glfPGRvGL1/A9PtrQUiu1/fzld
WPdHBxmD++jpjEH0/JL+2kkW8dWWUMxx9SRzAjOA9YnJupX4jAz7s2gXHh0eTl9C6lku2RtpSGl3
hG+II0xRt8pTK8VEg0KMjvY7wBlQhw2W537bld+X4W9RM57oJWFgBda8s42lfjV5B3ni0WKSPZfj
Cq2DszmMwckY9o58KJEL6zb6ei8sIrirf8LfX3rZrNB5ICoWT5XbZMeta63hp4Mv63J+eAtT2T8j
SG7eLaX8ObOpJYPIaz4h0SX4VZcFck9Xf1T1myKTcARrpbvpO56NfkAeWGzCS6BVcajNybQiTtrl
4rmwGag/MiXHb5VWJdtrNs94MmucGtO0bkV8aJoEIVozt8c6y1TetrWQcM/2M3NPGP8JBtNMINsQ
CJCWV3UDidLlrbA7/jfew2kJ2B83cuRqTPcepfAkD1H0RnDS5jFWO61ojE5iwfOo0blmvWSNm90G
+9vWwnV/j4vkigBwZesP6jcc7IYJprsOcrb9ZYsZ2f+QvKPfUbVHflryjinFJSjwTM3xp4rE+KmD
tBndsgc7u/va62RjlX87zZYI7prTb3ZgnxX+wVqHcr7GiPbwsvd2WVILJ0BbgpNJyPrLiTrKG4kp
mKoY06nyV6Hil7JA/m3mPB2h2ga0QKYFD/ZACTsjxuaSiuuEcNyyW9pgL7JjybKXq9nxpOF6UPT4
3oKlq/vMXvvUGvBNBhw/WLL9XXBBXrVkWuzUdmuokDGuo0pWanchCmSypGDeMQ6yfqP2yXadtgnN
s3qoCtD2V9Me+CwYBr3jHBSheQKRJjOsDFANm10cJ3+b3+tb4bXZ4/ancdDeRjco8S1vbAKmQUnw
qy0JbOJFc57aPFMGOt9CtnUXLZuOPmYyU5lv3tHfffYk2vdbCxGTFWVy+szmdtdUKOBXjK2XqDA7
6DQ1DsJ9tLouthYRgzgs8PRhopTqPjuhOJ/PJI4UfzFEfvPUTI97M7a78mUFqLYWmCjUF3DZlHr6
NWRKFJ3TEeHJPgfO/mg/x4xuHpx67eEhJNmJjvg+/pWJtMzU08/2ITfgbnyzG5hRZ25Uu4J1hzu5
3p2FmjL//IGUDYlV1sA4TOSn/YJIJauzH4mC2RTjd0f/l5wr4McOrK1vdSPpQKBvnTLTUtgiT6z7
nVmeWHmScH/u1Dlgv/JwpqyEVtTz/9ERo19UPUd8T/qX958LZnh/9CU4rb+EHHPVqU6gZ8HINkf6
itcyBorvSIldHHTl8+VFx9L5IfyV5ZIUBvbSDdUnF2MIPigimFs1Czk315e1bxXt3gcoaklaRLNT
AyKW5at7NzwlAAumyDKqKIWzt9gJ8m4/mvPwj9nCHJ1RXkFP5G9Iuy5ymYyK1bjtsQB7bwE9I0u4
msE+s2JevS0yNae8e2yT5bGtUSahjfGZalT/20XgWk89wwz/iTthqD8BBXVNJcIrOw0NIF32Rp4g
j/emnEFS0g+6X9paUSgLPB0JgofuMRPkiW5QoZgG8Z0Jg1fmL7K4RbOW+5pMfKoGblYapBdHxsOq
VLbeH2ANuJo0x66uLqQ+dNGvVRXyu4VDTfnqUv0wG2mYGEFfKJfqVihcxxHwJwLs6pPkZyY8/N9O
Js49lkQYnQhCG+Z4X4CXof4Whw+gcAMAWXQzPvznsUGvn7nkcJO37w9f3JS2I76qjX/MqTwNz8n7
BWomCEx1SraYo4a1MIf8wVnPEcNc2EHl+dEiyDK/i9IOdXQRbQvCXIJ7824O6smFJ9R7kvntxcB+
G5OCRkNzwS5y7KjzXU3PqT8KSwRfHW0L8V6xWX9BVjFpGxN94KxmB6xxYar/Wj9XbtaFzEYW6I1s
bAgO1vtbX9cswKkSA3azBDmZP38gvDZk4rMJOu2fGZ2rsNEx4f8JjtV30emtMDBFUsXyAHWWsdu2
gbxsSLKsBCk1jr7UgDTRXT4k1IwXVnktjuXpT1+Tg+r6+XPK7V4Oz55HcwpbEsV2v42Er8r772Mg
53jZrAz3KzQ7UYkI25UBYMWplnH1IR1jVRHOtuNPdrq6KbRhI6yTeyRtjqA5+IrEYYsDzUx1RvLl
sXYfe/O3KbxJunIwhZsUjBZdortwsYAJZ1zXySLShR6eIi4g1vNBOJ4g32H0kQ7Q92PHEdNeVIsT
Yc1ckA8deGB2rH65KcFssWQL7LKqYo3W3v/cJHG87RqI8tMm84zbExnaIACiDmlNNx1YB5wDb1dr
ISDSCic9Ml53vJ/nYQ+78jSBOjflinOwQNwoCs4vaPMvs0GnIfEQFoLliwpFSOW2QZFXJ1H+VaOq
ibBexNZ7nGsyWl9yrgFcWzznrJqvN3C5P373SFWn7tJu8nFG/Dl/gWcl9i6pJjESIkYhcU9pfwe+
pis4J5yhh7YnEfPww34wWcCwD8porXXUovTmON1BGs4o7rOnMHPFeiD00KSbRmFeP6QSL0Kj8Es2
R9ag4Jagc0Il7k6w19hox05GbgsBy2nMTtXL6PEuTyPBNjbL2SOXFHC/tHgB2rObQzafesu3XhG9
hFkGvUDuoL39Jzmiym1ytbBoKzapZa+XS9CyqV3v/FlKVxpSYgjqNXkhtpq38LVqmRTAExpc4/7T
QPgyAekyV5zvW1MNB0Uac+iuQyNKMSXtpWhr3/3YYrVGEJeOTJ/l/VPpBwbsTV6Ir6UkzCI0pIRB
EwIrr7aJWhO7Xo421koHqXH9SIhaSNLQh9DA36wUmYEgAq7fvATkWLo/T5cyCT8sw2wxv5n2/qsL
r50gs1ydvls2ThWoi+/mQ/X5Ent5DpVwct1HkK6sVbm9DeRcGaw8uew261TYudAk66mXFIcbs0wf
7NpZRfDx7eP3T10GvnaLS5Uq0pBXk+sqrTKBcKHyXI0fDM+7wfCsCziEGYyJN3GzHkaS9kSkQHM7
ohu85NIXy9NNq+hxvzoMXJronADM6tGKjr/D1VR5pe9hW3V7APaadfFS+97j5PpYJwrQSbVpvuWd
UUHgFBL6/Cf3oLXUZjU4UXI2VXfmLaJVUToDr82eW4Ab0DrswQehtthR4fjUbe5xOsp419hSXhPy
YrR7Tu7VBerqpKBUYJSzs9iG0V7y+z/Azcz79dP29u2kRPe8KA7tCYp688U+kjz/wXl6IhiNpU6h
G+hK7snb/F4TTrISE//lWwwYHPsuapamqgMpPs/1LUgMQMkugQjZgbPOV6tjjqg/ddKLDKS2OSb9
EQVR082zCZ+321ApNMw9dzTNBlxz8Q0WLU3Y/gZQBj9JMORkqpZEinBLyja3c97nDsg0D4AoncD2
An0qxgsjX0V+knHqJ/oOffPvx1EkfSF6hfri+F3FqCwjNiNGT7J52b/YvkHaNmJpiVh4dwqjdIbA
mgltwWwfalesBcJB/S2ioDFQbHpTs/D42AUVekEfcbaTlVr7+E4Xf8w9ZarIkAlISHJm8QtvbNH2
l+BIbHux4JSbzJFSUK0ang3oDVJoLDPpslDQya7+SKDuf04URIhsbCSYVDKo9mv4YJ882gLfoaGV
9iwefU10cm2Mt+gW2pE0BbG0/VXqfMMQs5K9j44tIiAMXEsx4CFAXcXmaBo1OAMi0rXRUPRMTPwI
tBp5rweYRcIt0MgfwvMjzX+ygA4ozSDR9N5XGvvv8zvQiDpX0nXghmPg5T603dlPxU/0uSsGRiUB
HRI2yizZSBGo6ksV3AGnBlRPqKyZgp8qBHRCCYwLJRIOlylrVZUkgz3vU9tNVRD/5hkhk7hwYuNb
Xwh8L4VCTuUA+U+keKgtEIclFfyHxpeCAsp4vbZTWK8UyKvAeMi0q3KzzPaEfPUZ6egxSiJmJpKl
3bIvSZ/xTxxH3TEk+ziDbpPR3ESXedWHfEFEElr+zm+s4MWBSVw3msN5Y9oNecfrD2HmGJU6xcvr
cG37KfoaLH1TloLpyCtI4EQ3a2jiNFh8eIQdtW+Scfi6wYwiOrMuALc7ckdhdNFfG8bz9AUI0Z6m
xvgut5A7Byro3A+DDVK1ZUOBGtkL5TcY/e4VvFTF36jObdbbE3ijCdQR5zkPJj6HpSXQzAz7FUjS
FnzS99BYd14dso+kN2xJ+n3lTG2q/VkexcledufAra+1FITQt/EF5T78hPkDecG03xqYrU1cAW3s
wZ9aWuRjWPhwdNp1/Al0NS+RfGoPo0neUYzAkAhoNQW0CVUC4DrIZJJZzlHK9BVvsRj8tRr59ty/
11i+gIvC4DxbxqMHmjLeKQUUmHLHReLgr1afQQsYROjPmjPdJb1hzzlHoPq6nUgFyMs9Fl/w/Qs5
y/rZ8/blx5WZezIy/96VIL0dTdjlilVnQCOvxVz0oWqYeVOdr5ijI8iDE1wF3XOjL8loqhT7u08x
cXn3E9L5+ps5U2nCDnbSidRgi4OICxxOuUT92vtfnlcFwCrkLrPOKtLsw0NHMP41NdI04oXkKlJz
FIDZAHW9pZNi9bKezehE6R//G0fn5mR+VbISk2/YxaNuVf16B7Jpp83RZEdLDSFt6AoNY3n7jwIo
wyGxTzCoDd3DOQoL34fdtV7sJ/IzErdl+hPLiexKJoCMv/N/axWGLmtOFBISiOotJ58kh0gLGdVn
5mJb8SrZlqYGIdUvSlJ3dSLsUadqPmLOJvfD1sWQ+NAKtJaZSH7/Pl8bK9/yCwsAXJpkT5SH8Oj9
aRwuH4+7f6KGuxFSbPx/zOeK2DzjoreD+HiJeRRMfL+CoU+oqLhO4RbDTRRd82KUNfiDLSS2t+k6
YhddDexcQvbPt2T2GTgK8V2bdzIH/WuGrxbnadpX0jLQdtDr4bhsnhCqTVOFqE79N5velySVYxNb
GnN6eg/u/S22c+INGEhoIRo5/nCAuEVK8jLQqwbdxK6EryTsjgt/FK09/3rcCj7BOh+2VPmoHlI7
b5gH2aUDI0HESs/HUgYBZFhSzFW+kmIjY9AanSliJOEAa04X+Ckyj3xodY1MD1ud+9CvLWfTLjQU
t39wuw/GLmvcX3D2KqJAVhydca7AiFjPq1frN5zw2QfcaJNR2lxNVIDWOQS03vh08L4iHwmOmKKA
TxaZV5ChfMYljtpCo7JsOk5RXzF8XIUC4RPIxXmM6WfUuWN8aI4TnqTQRlreESohGYCUaPqhEJ04
8Msaw6+DKC+ZyeiGGPcvevKtWx5yxR7OLOCAmAF9GeRasuErYDj4+5gzkkiqTUKyXi/r5R0u7zh2
I85GdXX6ksgI3sgEpxC1nR024rwLyZoPqXGH9Cm6tVQTWntCAkPHNJ6jjWLNn5OeE2TkfhiUzstE
RZb1XKyFW/8alkBsFQ3mHy8xH+4leUtbA3i3i67KQLchT3daTP3wp2fA0fnhUJbBcwd7cXWp6vkr
J6Ggs32wPLg6NGFGPxNZYl+Qv+z+u+8C4k+onBcCdkCNvdiVC5SBzv0Lnm7HwNSrlX7MCpkIXW6k
00CS+QjuXq9C1SP9+O383YJuYaaWAbGchWRu8OZcWbcvX1Dw7ZZlOKrCVir5LBa31dDIkpSStbD0
DI8xHjCEcYjfbvFNexIRXiTgwy4HzT5T0ZV+XAhZimi7U9UccQdTLLxfVOWjcB+S5eMJRxccqoyJ
HjbUkrDpdXrW+EMcve1t5i9f7ZNb/uc8o4A+ASz9Gn1WRQFfIzmJkBP4TNEpG3bYYG3FsL73bFaZ
rJGhQr6d5eGz8/VnOtDkY66Z7hKLfHil11w2eG16eAGk6XrZQzr/7y+92fNDcC4SEq579EiNFt0T
kxak95GXphevA3i57ngtGROc/lgmi4/J1UAb+A2Uwgek4wDZDRiHVh7kcZIANmfUygRa9ILtwD47
0XVYF00k8Rb6G6UJBAt96eH77vIm52+WUWLup3ER8Pvt6/ntTMvXd5qo62Oaxl86r4gWE3M/r8pr
VnMbSB41LHTYtYenJFD0/MTS9mTWulayI//uLLTZ3418Br0MNy1P1+lgLTE7PB/mULqZhcrn9xO+
Vc2IL0vczN5XinTN4w9tAWjCN1kQ9aiFM2mnPPgR0HrKfESSIDx/vKd2dr1hjaEnkC6Dm71iTIYY
BG9skX37UEnPvzU/xR3AS7hl7XOJHsXeZHVtleoNvFkPDEeTN+Q7LVH1RiPxHca4X2xIxIUSj2D7
NUKl0q4pzZer/eejEkoQQVNzEo6d8yICzPhhUKEse92du9ikXNwmm9fKuUN2EDKPfcij6VHWhyC6
EkwhPqr2CjdHot/HrnclhqHVfDzVdJjrOkzpaT4TZKZxx2PGe7i8EXlji6U4hD37PRAGMOM2kVSZ
pxpdyRH3Td9AQ9aB6cxsA7xUN5WaeycXqNTJj0ZbulkwiecsD2RzI6KD/OOzIPwxLWaQ3v0nTwLT
TmoHdBXhodSEKmNMsLJQ0yZTgAL0cy4Y+8ds0CvU+TU3Bz2fnn7d0FlL0gcJ6XhszHPtGRUD/+RY
P7pAyI0pab8qztWjen0PorwTw7dIpDt8KYEoww7XhqsB/v503i/ecSe/Cbm3rSVntqNI7CZxpDU4
Z60Lnta+3LkNGEThpDMn/mJQnRUmlRZOSxv/6csU0qFvTTbsEV+wSZSq9xyeCtE7584ANycVtyU9
RAPK2VAqiLtajISAt95if7KK79ZR4di2dSzADyh/CUPpZSJXpVSk5JRm6ml/Qcr7ogS13kLp/wnB
tu9RoPFg1zTm57ZHymGUm5+TQo6OC6UycQj7ziu7mrgo/5gM34V63ujlAxgX7Pj2OSSDRAtoyPX4
EtKoWlnQomAYz+aW785YUWdpAp9I1Uks4eijYRZO/V5N60EDqOp5LH8Lsc81zoIS1La+it99CKGN
0usPgYzcJEYYqYkR0WKifWOP/Ti63fCi7XLOthqQ7fvcSluN3b/sdDpzvBaomVhzFfE/N+/rFcP0
noBUujz5WJAOq8SmLhbJKC5WUlkrKN0wTvHgaQEsWez/p4kPua8GuDixRrRdzeUBVjI9t97ZdHis
mh4Ic7VySnWbgR3dE3VFWrYsDYDEs1N8LEd0eWPMCSu658+PgR7p2S1BReL8E5HtP8ayXh3bBGmv
2R2PLudDkiPuSQabaNzDVCOrqVy4DsKX9C9DH701SBpSUSvUM7ZN0yyV1i0w5MSNFaKW5jnjniDh
RlP3RwWmbCpBr4NBdaP0A/XNz15snjmUkVW/+hOfGSw8zhHImik9QwTrN3s8j8uQzrNBGjhnF7Mf
Ml9PksgTmxKx5KwcMEf9jqmv5f0Jr817dZu86+MoIjGELy8rzDEa0TmdDYLiLShvyUS92GFk2QJT
6Y/bjNd7oTLhVN/B26d8viTOPVrkPCpNL1q7BAZYfjv78mZp7ycqJfOlZgGEoTn8nH0Ys8EKs5yC
jWEiD0A9b4Vb3fgcPA6y5NN/wPoZzQgqxwFkuwwJIBrx2GOkc6Emu0tkWvrCiR8aigzxX+xToIx8
39E1R0cH1+gC+EiL25iRxE+3k3OqqahfWBft5BuGxfem/4Sd9rHf5cSBTDBDSM/RX+UeXnyTPnDd
RPQ21JNdr5FyqbU40ZjuWFNF8pWcFq9B4t3mZ3y9vm0qKyBf9mqgdKz0ggnmuKh/HqZOndyDH2qA
wE3mb64ZDH/zc+wJIrPRhIVd+iqnutV+Jz+iz0YXITHiM1tPVQbgjQ0ccL9+rc9I7dymsysFzAKQ
kc858up683bezJWApx/dV+wnVlGgwWOk2P/DHHtPjGx5edbsZVgGOiazXO/Ki42ArvGC05gI2f6U
YwBVDxbnfyppz8EDHahGWsl0aqdXqY+3PZMaGZHr8biRi5vGhXOMEQ+moyvRQB0oZ2wFi+mnbX6F
j29l6YlcMyzcKfqTK/prjteJRa3qryNKsxVgXdtoT68+hrp75cEkBZn/IwpaXLOZQZ8RD6wzxZNC
mV0zy9UmF/cJnTzig+jBLsd0C7YCWORIAdJqMlCWq5/XdqAcgVUdfX9IPnpwxhTYwYOTYR2Oduej
dykVYyhu/M/YxbSu/VqQMXrqqbKOtKfly2hPwvZkKm8cB1t1UryCpJRjdzexyMvuvCFTaxux/Q03
tyebvf+/UKfXMX/jO/YBZT/trRIkX71Iim4c6RM6nksCzqTLbCxAs+iViF1tJhyA6VywZj/81bvA
0jNsBPW9i6v8oBx5ZbD0vOdMoWu45Vl5jmbMw3F8Sj4LuOBWnlR8uX134PpKMOgWn11vVl0TCAtC
t+DyWhhgVBUpWfcP1YbNXqK7GkQyCRJtIU2mYCTv5RWAkAfbMkJY1DEeqZ7+/N7rAxknb/ScuRG1
xNhtgv+VzNLHqYOQNVA4/J+UHxD95fpmcvjsWxMv4r4EuPZ4+46prCv6MUiz2GbSYCM1l8KLQQlm
6tKzLoYHh6sG8u/arLC9vwSXSJrYrQlhcdn+KzchMsQMh5vIlyVQKHp7GuWhcjFRSXp0i46GPcG2
at0oFkWFnjqKSPon6rzIWbR3uEDEe/5zflaYhpL1akzFDsZN63OzBdN8wK0o12A2hQMbAsqFmU7x
NXOfXVOtrE/AwrdarFj/Ds+2+eeHFmHUrQyx45SS46sYqmdwTuJP7SmNCUFustZLHMbjSXNnRyiE
7mCV1eGjLfj8FPCg7r8/vsY++Y+fyQQtbPqd0rkE96n2zEixGp8gH7/lvlu6clQn7FPTm7jrB5wT
zov2lamCUPj0r6Wvjbchg5UGnlv8r46EdRgdNky8I8dTLBzCWxkZWq7XWpyZpBUyyG7OOj8pAJ74
Id5/ajfsdIULViz3zrs0f85Nqt6COAk1X+tPr8QkdFX8FND5U+OBgy6Y98U5pYJoAMIwx7DXu5TB
Vv3Q8T7gO1DGHjJJnaDa8w7DMm/MpJBFsRUxFX64otyopX2lL45u6phIo2aO25p6nYLWlVMvAqSW
l8suJMxcGd0Vnb5mfkMFNtCBfXNrg79UNgA9JA90k12BtVFI32NZCKWnUOqpnt+gjhWDuLKFBbMS
3o7pPaAJgNx+09PcrsIW3FI1eal7CS1miw/nv13mD9zC6tSzrD04rgHyWxxKOo3rF7C/1tGnoLNt
mIUz4FNV0T/kN85hClU8TwVKPzm8FpZDxc6TqRGiM5icjq+1akylCn6L66pHi4pxorRcOuUvgAEY
LmtI6JzkL8RY6GUQI5BD2IZuOqaXLr7WvlOVmywB9aojpRJYxkU1fzfhzElwG14GWKt39anbTBGG
PbAzy2sRUkf28WH7CUh1FyOpsyDbFSMJUYGVxYYdoiXrfdBsnAVLWh/VCYxX10jk+adSeVHEytOk
2c3aeeCkYE2mrmd9azBEA20uy2P+UYEGZfhD4G12tfmKypVjnUiP1fUOYTcAKrBT1ZfyAIu6Ju+r
ohkuqsp3wDNGbFkW/CR1CkY/etbVztEj32jP01lCjVuw5kQ/QCBAkIc3PegPl8NleQ9Qutr/Xi7P
tC97e8TOSWob3OzHBt4k4UaJrFRE1GY9xL0POFg5ragZUfLRQfNsiDKxmvS7BX2Lkiifup6rlO2w
RThF6u7DR/03ygY4K+nZstS3yA183sOXN/oW9/ghHSuUT7uhGdqdjLJndnX2TTsOzFRMv7BlaATN
7VQ0JHzV82W3em8ek6Dy0akV7r8BAaBOiRCq7vaaToFog2H+60DjlHX26rbG+5xWD/YFGMFXs5JT
/L9O+T2RMIFizG6F5Vt6McjE6tfs+gBYrRJe3iJcNZPnivf+iH9LeRwkcZni4BGY8dufHCeWcYx7
Huno95EvmDJT8sZbyVFMgQmZs81QZuU+1zqTa/h3Cgvf9x/iVK52gZ2mJL4XKBXyS4x4oGx1VWvb
YVmspmB+lV1RX4bNnLOpcHLjU0/Nj228IHInFV5m6tuIFpG42rPeBsf3I+Ct37jJ9jgxY7x2lMBJ
FYADN6DR+nxX7+s39E4PGNcAh5P2Qjz5eSpfnVtm6Ij6pL+3Y0JMAbd04/1yZVXuYVbozQK7eIn5
n228+XjnhaWgPYmr8vAJDlVFKAjtSWthZyxXYBFc3lpvKvKmNr6TeyISRK33iVs8TVnFN1NF/SSI
bIPjekIdqhQDDSecMpGMDNeXsSQ5rMGBvOxHBgmwbhi1vbRO3esoKAi9OFw3D5cCej24zKVg2YcL
4ptaM9r5pWiw0kpvJfZ52TiqMwEFKXy06QHn9q3BHcV8jAlHhRWMltGJQv/cUjHpMGUUz2PJy873
odTCBXL74SiV+sDAKWTCRokcYj46i5WNMPc1rGRLUFD+xWmm7vcqRwq1N+z8iZZ10Tq+cpK5jCOo
/5HLGnEkYoULMyMDQ0bSN9DEr1WaaVKsXWZSnKWM2Natk97i62NM/xvOYLUHzowfRt4g7v7CNsvZ
EYQCS+MH/rgnwwW9t2ZIXMpGICMGOv76dkUa425DgZpsm6jvx1XsEsqWwrQ0sAQW7FaN/MGSFvEB
uQntkNzqAC8KRnJ/DqUs6CiA8+44m9rb84hzenVxCnFPWHx8gUafXeM64X4ePt2ujMo/7uu1mdT4
D+VfOnlzXBl7VfRU0oOJ62eCJyyrAur0i0QyHup32bqwh1NRNtPL7sMqXqQNmg80vvcfdZ2CF4fY
zC7YWCeQYlpY7vKtSnmKoTAn1WSdQUs/tmPXN7CuTL+Vpl4eOZW9OKnyNr1475pr0p2OVa08hby4
+OAlc9g/VSYtWiAOiKSqqcgA0Og+1xOMdg4KZN0S6Fzjv4wRY+BpkYpVte0XR115yvckeZuSix/k
WNrNilIZG/JbbAvH45fJBsWv6srItFam+KVXKZPGdUQI8BomB8aIbV7cVU/XZYg2jWR5yXkD5BwP
XKZDJBMSa0lBpbs1zWCx1brySINdJcGTdIILOnr9bwrqzSPKNxk8YW83IIfpyIDvee23XhEGjUc2
XMvphNnzpk4+b8e/iRfpRraDiIEl4uHGWX1VAhxgcXilvq8fB63zq10m4W2zUa7/KsBMgB6f8I4N
niFbXUDYZzMPs2oKr3JDqT0bBDZN3IWHtbgKzamURDlNj++pHod80xe8QJ4h+s3Hs0NU0rdiYk0E
9bnkrCsHGVMTx7nj7huE+1etgnZWqJMfWi/IFZvdyLoYxfr0vyHvsbpXjbUOwfhJam/ib7qRQkpb
aF3XFNETJfkm9mVMeXtnc4ZPfkkjmIU1U1GIlAcpxlfh7t//C4dDkN/ZrYZIiff68AQ+wY26eSkF
1uQlRio9jtl9uezWRKOFyx3+Lp6wAHSV8wttpPdxrzkShhHv9Loyp7BCVgcXUMSlJsrYYFX5cVsX
Hk1k02HA54/Vau8tz/Dr8DM5mG3YEmoAQVEcZLjdBS1nleLQfjcFK+4zaq7KwkCAp6b6VPQc437t
9kjb6JFsgAYrYOTrlsrnoqvDQBCY3eyn37VbCKedmNxaBvwQQdpMLM6w7K0d6lOvB81Vf69iNIw2
mI72r79W9B3k9ETmaF/TspLvAuYw8RSYrkpzIXzFPjzC6fGSSL25GszxFMsmYjmqmeyXBAfV7zWd
sPrmcyWFe+Pyhut9PR9UOJJeb0nwHzpTZivKwWzd0CV7l6bwPhjjSgGUOkyspnlkWUWsDjZ/IIxq
7Wr7St+ZcytB6hhLyN/SyL+yjgQoIl/oUMguKeA5+AzUZfyPA8bvvGk6MKG48KMY6pF2BnxBWnaH
NT4t2fuCFjzDXUQ0V3pELeb5gcODdwdO3FCkazW7rRYLOu1Nzgc1g7uYlxLcI/R3WrltgVsp/UT4
ZZVeTQMphH6zABo21bhv1uIyLVqrQ+CQ7AxBBOtrg9lr20WbkpFDGp2u3JVKxWf14yrL2Zdsh2qZ
sy3uXzAUr4aaLvOLF32Z4kguegs96ZvNiZlC7V8l8Il4i0XLq2nBjnrGl1FhfquVayiagRr03u/Z
4ygf7TKlldABq7PuADfSfaBjhy0hiIzhvFSVMfFNlI93ZvQa12Y70pMeHWgvfbGBKKCxTQ5tt8j6
s/418BSeesxANWJqRlp+LfFKU6+xFzd/J7yNkoFVGuRPDLqVdHPrkEi4pocutZsTa09yEtutZPiq
R4uisBaLuuX3ZqVfDjZl2kgId5un0TtD4MllTXXzuuK1I/iP/hcVQchi1iKklORtgBrapduQz/7p
h0PQVlRATt3aRtFOG7vw/NXrRwLEYdsZXadIEWxNpTQbWFC0BTPdIqGEv2omJT0tKwfrdy0wP1Ol
e4zmuoo8siyy+aU1PLWt5F+j4rxuLuYHF+Fe8YMyrcX5uNrj/ussx5m7RYytlMWDPjNtiDEIBNLP
RIA/lSFWCPE1xXWq9PVJOTwMrqNVVYdcUObHnegzWGSuYEdBq/Hoiw9YXaB2apiZmvN0UXeCWbCr
NmDwzwpfofaeTP8M0HTYeKDYvmRwIJCnOi9Kb1w2Cyt/79G2kQ1jtz521TevAr41la2XkgCKTlYn
YHBssGEmN0AW1eEOu1qenOFg6XVy/0HcmgVPcLi5bUfs3gGnIC/pWokmgrHRKS4sSH9pMW5ReOCf
jfLFaQc38S+EwTVOtGHqJ+idp0moTtzK/nC8y95iwb2HaHVoGXWMX2/HaQIkEIGfzI1F/TObZnfY
oksf/sJcZMXeJxcUrPqFKpQu3wciK/6zfqas7vEUtR5pC0Fv03L4pTf6mEmjB5rGgbZUWW/mS/RV
N+lgXA3YG/4e/RVTLKf8mQtY+xb2U2P7QQM+6/rm7GFOOP56DVlvHNO/5kkoixOovATk59CBy1x0
sqQPfM0NLvuoY8ccUp6dgEgiB/Ioct+/cDeeTVqm0tJQAoutyUikLEY/Xdff/5DCBJlrP7m6r2jc
YEOMZiHnUIFIDWX04gOI0JVqiwZ0/0915rNpLPF9VHZK/YSdhxFkcfpqfBkXP5Ywjck79uZ8YbAM
Yz3NVQH3Pr05WpRHqsQcsvRmwCxll7C8h5pTKCRIqJyfg5NNBRE5Rr6uWn4cFYn204oREKNgYlR8
mng0kSsMoiAAA+ZvIhKsPoDi598bXBLxAg7F/YgnIBFZ1S3jo4A4vtBoOgni+vFR0SHFAC+RJTTe
ItYqS8LenxMIN8meaPal2rIdS0t7GSrgM3o8QQs9D1ZXhMFqVLyeHuzlfnjYbD8Ip06zkkSEnA+m
cuUyr2qmme+x/Yue57tewlQN5Pnyqm94aW462Vz2RaCGK2EsBmCpcHkFtBP8c1voZl42c/ODVFEF
2d2oVv9VL8B4+B2LCEdohwra6PW2KIrPyzso21OZrOKAqB69mw6KhuIn3KaiyEkJV7v81asn7L+8
8V2KhBNALO7KpuVREXS0uJymXt+o/0mzpirvLzRBjaj/uab8nBq1LQRmiymhwTjv/5t8xVN41aoz
XTEOouhvooqvnQCKc7q0XzsZ4imZMHFjuLlp2wx/Qu1Py/eRYjVvPrTZGI0TRxTOKdtk9cvj9qoH
AzoGayaxJjbnZMLyi1b+itL2qqTQAA1t4wkq+RvRJuoXGlzb2qJn0HhzIkT3kOKgpiajhOEQQFqQ
NhnQ7j5TrYXt0YbT6u9idjEyvADEO9Jy9rhWt81kN36wFcpc474Kci5vSju4ZqmnSmJhZ+WDXpTo
E58Ki/t2Yei2LbGiYUiYJo9UHro8ro1yf0ld4Moj8Rg0YxrUB6giYqLXePKMj9jXltI/Qi98sy9Z
EKjAt2j88N1GmKsGvrDdh9Uh/8D3NXWF2WwUXTXWbHsnEi49eE/p05T/BUA6oZBKW7k9PQ6g+UKI
C4rSRxpAhaW+8FRQob5VmMrgm9WpNPFp69fk4gHsxaVfC7/UtafzJqiytdDhAo/H0bdhOgtk6UF9
JN8cUenuH6KqA0ye1uOEXBFhkINsaMIuoMqTxZo2tYn5TAOaQYYf7OZxyDgwQv+Y6O1mtZ5NMtJE
FkAPeJLreOb0Sw/1/GBJOFGCxUlLz+XgRxPnSllIVgXWlxgCOp+KDexsrOSJi7TFlXvPmASz8WaE
3syM/+SxWn2dSwXvThsC9NM8VUp5R636eRPjDifqJY7UTERKTUUNPaRCHLfQ9DecR3IM9uxCSA2w
1TclObfC5jfei3oFDTdn425CDA10FA+fKC0rRrnBQsmKL/Z0Ov5kU5rRHRnW9/hHnJWkskdFryOx
voXUAW27zTmrkL4DEpYdul/UUQtVkNdy5uH6AjOZAVyHvMTlpKKLQrqAIcHPsMC3eywlGmRkVCyH
PbThjTZ1TnZa3SEg3//npZolR0O11oPtOharJnJbnZh645zzFzVxhhPIeLpwiqZAuxC0hfOwtF+K
s33PinX2i36I2UBeZip7ctwAzKl4kB3Qkcn7PeN5wXfzUoHzuN/t6w6K7HRIVwesfcNqQDYndq8U
ATVlw1JpmSXxScZnFLBFgiAhvGNylgnfTR3kwTTsXUEGeM1Kp0OljnNWNSaW9zKHrxWiPHDNBKh7
yl0MRhVrS/xBcNCYhwhNSCMgjKGpM+LGEcbAboqaUWzutHAokQdRU+gLRb7iRPUq6kPHhjwAf7AB
RLWYMilM4LWJEtgdgua80CjaxoXYprcPD1o/ItzaSMdhU/M6yPciQJfu5KDzWAkFIAq4ykBSaj11
2l+3lol3B20qI75ozrsmzir4XGV1swUaXbKXK+NzRRTI46964BwCoCy0c2KFGPp/b0MYtSKlFrvH
P8jkZrlWi5hxp2oGgprU6Q5HhMQm43CR7feadLxakp0tH0zFWaYME6qlpr51C0tbBTc1WHZNYfgs
B6Ut2RCpQww//rV1WC6kgxTaMvEYfJgi4oMCrMv2sPfKRrR9d1f4FnXHvqP0Yr6tVRAXFQCxX3lI
SsQ2fplejmFIIdZlhmV0x5ApqCx08QSMLT9iR8xMD31NUXveTEIvexoU9yQNHcMJravE43gkIJD5
AH9Ns/8wgx/i7yidwP4MzOG9X34Pu3CJ1NmkFldLM0UpmKT0OdIOhYG/1sGBHeHayZ7X4gv3Dbtg
lTlfroMnLgQ7190N4E7dczKXVv7+BDPA6V8KkVZkJLe9spr7J+ZDVsvMskfCEMjmxfuvI6SY0HZ/
SnVyFPLqDpK/6ws9gAftkrXepzIIlq6P0Obr+POo6sSt15nneUfhGz4v74rhNhbyoJATuDyDbpuo
VHQAHzezaYbkBAok74hLKX3eUrpTOhWLQX0sciuj1WWaano5QOFwon/14Yx78BlGJukIcAJWrtsw
1iAsv+ETokqdMvkOG4LAhstzi06h8G2komUzBEPF17UhXwXVqj0eNFl1e2lmz/Oak5g8qDHrdtiu
65i+VFhF+1t9slWk6uKSmBShwl11BviRtLdqC7T+KuFgM7BnJzSFE0UHHKLIxJ7vBlnRXLDFCyA5
fM7Rcmrqj9wxrDb7URDk1latXWIZfRc22TcuI6/ovAe9Dew1ESKf6YVusJmIK/JJik5NLiv719qv
4rexvaSr9Adn6mtH39tYHAJ2NnXxa41j5RrEAfw8Kbi6w36K0ULK59JDqRkm9tCBxvS2EepSyvF4
66AWabK64gE3PsRANF48iasuW38Uqbwgd+4iM9D7grEmhsW9loG6Atu+jYfMwBIHAwZ40nJGHd7S
N2jjKvr5h5sB8VZLVdi/9cIvl9Sn3iIX7YOQFGAyI7zfjIoG7drqfOKRqRAyJt3P7bncYgTKigVq
ZihDDgWcLP4pZEUZmzyVpCg6Ha/H4H4GSYS0OinrPWARd2ApeCcy0RRD7wnE6ER3HhEA0g1ifQGH
reQc7aDgEEyzjwGtQ3k6NJaobunofSxq9ocLtvlaBRy/uFTVZy7asQgvJbB94FHa6ye1tnBd+Acp
TjCncpSVf9x/lnHp+wAz4DOPTYhc55jmVEPXsM4jKy/0Po0efx0AyzyZGXnarE2Z+sWiBX6umsSy
f3S/xt17IfAUxAPRFBRTwY08AWXcd80Mqf3Rer7mW5QFtA/apzBeOgmM+i0L0tolv99truPrfJPY
7pKwTj2ZMsEcM+QTqHUHUbHAtOe6XIkNn2BDyL7+FbokcPHcXCdBqdVKa9pGL543176IeuSTgNtk
4oRXfYaRMygB/Rv7LZguhFTiTdiou97OgwkQTtPLlYxJhAzmP3QSXHtlSw3S8rXqTKhrmr6kgnMg
lXIKUBwINS9RP+ww0h15HWRJi6pf3kj3UdN6WIGKimYr8roeuZpEFCrBtFCjfkPLt7A7W7LaiW5p
VSy82vwZ41+pOsO5omOp0jBfvYl3E4v9Dcs0Iq9VHN6kxWc+248k8+CXT6pONNk9NztSxWDIFEXX
9EWeqZ+y7928QamG1SuI+Al/FmRoZtKoXoZoJK+PM8Dg0WP2hZIY650RyrTy6mn0SCTe12XGC8oC
zeIg+5kDA5pSN3fFNdQzws9j6+lksIxDtv+ILvUHiArj92a6DQBbGLHSwB8DUomGzbE8PypKtPuY
/bjdSUwt/nQQzP0d8LADc3DcbL2+yI7r+AnFLYlZ5u/0VoIILsDfbE8IFRP7IKkQhLAumw2AKvRR
/8wydzwOCZ8u6gjvA873/eIVhAdHKVOXwvnwn0LtLJMr/26r+etJXC13d7+c8e6I1X8S4fZgDI5D
wXN1sBw10SFghDI7GqVnbQ50gJAPXBOv2e6SMjhDPsz1Unc4qazQz6nXitfQy8ZmD0dFwRxAS/NG
iuQKH4vKcEcZ3pq3coU6wbij2Plkr1tVrO90o5GwNeDmdCOW8EUTizUBd2qc7BjoK1Wh7IrcVgWD
Nfs4RN/uahWaLB4h5bqsyOsz7g2XRPRH6ZI8aiJjH1Opskey7ZRfuMYbzF743JllCMpzt3BNHGmQ
cpMaT2Lm4f7bxN/8sP3QxjAB1noq7hHL4GED9ArLUkwdLlwymMCawJwopxqnkMPimQLz8nIfDLha
xWt0P2R3fxoZg+7IBEWJDU1n6ACjH4jz4XUN0zF/7OMzuqXFTGuUvkv8EdI8YrYuN874mpOcFWCS
3z6erxD09QBortJpw/+KwW/aA/W8g4e61dXQaS+WkdGwjW1X43fJSrdm6PUhTTJnNAipA43q70Gi
IabgzU1TG2L5UrlZukzFqG8KMYjgtQnFnmhNUjvhZSZHDWigyeUlMQfluphpt3UYFqLYMOjgL/CL
5uWoBBa6ehpKu9NkttZKTbLj6iCM4HIY9SrZ2ZriYW7EcjZGJZ57rkhR4ao0DKEoSbd7EiDttUkC
dN7+AjiQ11bJpHNQO8IaNkSmuFobt8nFs61ksTEmK8RaRrS5K3zjYCfnAjR1DbYtYOJ1UVbfockz
VpYwIBWw6CjsVEtqNVFA699JmbyXxjM8bJDB15AawstCZqzv/uhlFWgyvlQD8RUfQb+QYrOd9QW5
EttLRLym+zVJ7++Y2qOsMMaHQmHrqKE/FnLB+7FfQdY6SzJRSHE0wbGitAo2IRWstSXp79vXNCWX
NZJXQEq8UX+7SzGJSLqfvzl4uPo6XRDeTPeI+T9eJTovsJAKTW/KmKvoNfbm/NFdsngz/kkTMUac
gZyHlBZmKymj+4VenifEM/an25ljw+kulleCtBgEiYOprhvy0S5F3X6c5Oz3hNuyzi3YXCYAAVBY
RUTzljS9AFD6gf4NDyMFEJRobLngvHNrwE4tL4ncaHKsRLeeiL7uDsI8Fy/vUGK352vGfUp61ANH
Hy7V05mXrJELUZjVoO6OUJpi7tXNvfX3448Dy4o14JnhX1xshl21Kb8TkcWGtoiQ2+JRTCqMpMK/
/k/wJ4ABSnhed9pkAwLK4ZkHYDROlmZHFcDhVKL0Lzb4Z+J6omNziQTI2rBpntdEQvRSByIXHwZf
cfvUHhTaCCVB8EAQg2AwAK5Gu7hCyFmSPssIVOXQjEWa+z4SP4xKDLlD7JG6iF7k/jXGj6NXOt0+
If/riKyc8CY0lbG0QQm/fDK4t15y6d1iM0q/Tc06Z9KWp8pWpKYuNAPuACfdb4/cYxZN1gOpabkZ
U0rebMttZEnmvPCkEdVyOf54Hi6glFaiTl0QkpdYnCh76hit9W0fXFeTx3OX+oGiNjRNj8C1fkMJ
fkNZUtXAL5/EnGGibLtRKkhL26dx36Po2MsAWWEHDVVALZq6ouIVD3EDGq1rM7xNA1OQLzOSNoOl
f0IYxA8fiwIwXMEde7OJMYwo54SGkctnt5aYsVtDZn9wfmSv9JpI3BO9Wq40lbGzMHbf15r5JFi8
uy62AGbs6GLK4ZJXOmbbLKBrXsgWG8+Rw5RTp0gMUx2qWIGJnIGBakFTXqpNMxfuXAe8yU1oyrxC
XB/YrDbnkZ0QW5/FlmeV7G2NgMaTAEWyxmy+PFif7agOgtt4JsYnLkfsqC5t5s1cVtna3Dp6bD0A
hpaTaIIC4EEzT8rMsRT8LtX28v8eyE8t7Rwl2w3mnJ8xhzecyIwpaJkY91PB7Evqfnpz8qhGCGxK
m6kaZ5v6fr+XEkvNeHgeNkYZQNIxWv12pnHX2qMwRH0GW7ceKNf/jFzZQ/C8DudNqpq3aIp7kpZE
TUGt7KrNSh7F+i0x2dpVnWurSDx5Wd/PDYZz/GtjRbTDIc48NfXm6Mg4eH6UB0PmbwbeH+sICT/C
g6ovjxSlT3XXfzkLXSMWlenxDFUMa4eim04UDt/ccRUJAO0AmOTTiYF/wuATFRupdS/hcs7RUsFE
YH5sIeEC/gYYhbXfFVCOQN9t+5rWaBYIaxRUO1GF79TCfbey8CDeze3Q3sApLFvqB152zBxCdr6h
6uRXhGEbBl3I7NiVg5XlfUhIdZvkK+yle5ckozyNnm0pHIXdhIcFC3wWCWc5KkeMJUqQmHAA3XeX
kGbD3WznCGCMF0siyPo/LJ+fJrfl+0LZej7kmGgsAzcxwFzrO3WdAGNbh+6hQX6i9c19pvSh4DEh
dY8As04c04VG8VCnPiKB8iQRmDDQwvo6FAgtgMhFZ92SR7NWRnSlheo7OQ8vZm84DSeWtryXO3W+
eH9SUPY+4+asOdUkAIhHj0A6zyWCZ8lEVBuhHHjlZ++JzQYI270DwQSkmgWfAyZxjO5fkfniCy0H
3P5K8L3gOmf/B8rSVebf4splszkwLakkE4u+HhJCVi6r0s6YssqJmMzkmAPzv0LQyAI5es9kftgz
D/SxpUjObGvI8dYk3hrkoAcFCnI/0TYz+C9NBD//DFi4lqu7HPaRk5tqaFHCvOeY8K4lzL4l1+wH
Ryiyl93v4fcMFzgewq284ad8G8bebpaU9rqIRIpgernyz4VsQap7DBrsUgj2tf5WvPFUhFHr7gUt
scIVL9SjBrfA5LBbaDVAnwy6G/rz05s74BukcS2HakYhIF5/3aIQj32+1Ig4Y3Zl5bfB6+wrDq/9
5wsh7Kp1j5wQqc+me3asE5VWTrQoemHHX8vTDqzYM7icz8hS4MnLRuvtsp0X4yewY2uJ6S/KHAJI
aCKG71rIWkrMHnEopVFPTbA8dKYRTOYSoUtcJXTi7cqxEawlpAenyh2bZVbZPXtLHscqTXnmGzR7
Lf0Odpl7YRopCmk9rOF65o9oJ3aWduj55RAiVFylSb2aL3k6+HoPaovBiBYt/GxVBDn6ZW9fs/gw
itg5G2XkYQ0+HNsI25751KxXfeZ6QTPCvlCBwOQ4DGhEmwt6s31RmVGbzrJneDQfH6x8kg0Z/qtX
oLIMIT8FegyESKjta+uTmOfC3j+MiK6RyilMxDk+Id8G1iw1ZdO0FP6SdordHILeh2j85pvnbp9K
dLxOv2NKh4vWUosqeBq2GD0ACTF9jd7MUa1ZPzrwf24eBHTp8yn9kW2+P3IQtX+IKbG9ElM8oHsJ
UKp4wt0kqRCT6Ag/g4r7qfHsepeEMa/EoLJuCgPhQOzRHJYgPD1kFZrbz5e2RxGuFTkj4SW59RF1
cCYpIfJ9liwrBZhfcQFtB8cAe/9mJQhZOo9dfWmQ8Q+DbWAj740DRTo5pxa5ZSRrgotJt/b69A1p
H2R89jxpMEv0pKpHcXnitP5ZjGUpW5eQC/IrVZZgOnYncGI+QPezP32n1Yy3TipKFkql8xMBRns0
ksqa05khrhXbiWHGYPus+V3mx6smqk065ttdCjvNjcFcPCn3nfCM0HEVzGG8oXk4NdAXYr2FtyjN
X3w1+fx05u+sDySc2neCiVDm3KKqHcIvYuE7ccCNDhjbRCs6sSIb4oi0ImrpVgkOElfY1zUmBUDd
J9Qgaf7ZsGPGhZbXBX9OG01bTzS/lwESBWXyvbvtuiqsIipEAbaXKTjyrCNCF6M8x7Zj2GFO2g65
j6bB13Dv2Q3c/i3yc9XvDmdRZAJzEC3Z58kazVER20Vl8zIGajwnhvKBGhrls+4eLB8JWcjcyPoJ
EBYiAlsr0nB06xMCNHekiT09ug2U+YsxkMVzcv9S9YVfnd6jEX/KoYoVAsk8UNOZYbUBiwtfryR0
YDLK7bMwz154CJL7ylG9VZGlHmo40t2idtRcMCZpkdWUb4K0wnLmG2pHiUdxM7Ms+mbaDdY4Delg
SP8pcRAA8nCSDqGe/SbqD2YzudTtK3b5jFDD5+UBAKwwuL27rjOmvF8vu86j+uA2h3V/xq/zusjm
ThR5XgQ2flMe7Rzi5kAWItQXe+mi51hESr/Q3xbgNbYcBt5A5sV2IklwC3h/37VBIAkXHl1dBWHM
Kw4yqOm/jVP3bNdJYkb86/GQy37Yq41fDh8fiPmnYrZz7Y5suN6MYllqlXkVh+1Fxjc11n8NvErh
LWbd1g+Xnh0aTsSHHw1FdDHbELufTLoNCMenmOHi+P1xxo67eQ5fKU8iy7HK9NOB8tD0ch/VXOg+
H1Jl62rHfxHUnWQpOoRBt8mPoJw+1LQHaVfxrelUWsog1CvBtU/cD/DH1tTxacomEq8oB12dawn0
DdOPmZX3IFyIv/VQ9cFzNOInx2ntJ4wPj3PmQleMxJKfwFua91VzTVVJGCXcPk7edXwZNTRltnrq
ctsHOwKG/6AMSq1vbaZsZBDjcDxwdA7Fny+EwyfvJhGaJKuYtepcrEaPv18ecUrzcQVxwsTwahRF
1Xer6RTYQF1+XMmuLUt9uQrz2MdIn0EMGOKUczP0JiGN5JHgEo5UO8aACXe4LoVVNekOJ8lNsbc3
qORwUXcjry/8uwfDjRqlVjvNxffo+FsJZ1Qh14vFE0YlIGMIFuemvB5YY4n+6ySEN76JP3CER2Ip
jmAsNiP0LdSkcvcrkfBy2MC8tqP/DsHl7L+6f4dOH29pNQsysB5GDJhoiLV3KPFx9vVwwW9JSJbw
XgGy03rCtqi3eLDPdX3zChYt74jNPucuj0JQPiwdgbnco2juvF+4yCp/XO3j2WuEmxH8KIKhTkIi
vPxYftIDjEHu00y5yu5lVADZX+ghmi+0IFu6ruiM0fFpEo8lrl/Xlyz7CYSlUoimVGS7EKuTLJve
Bs+GoG6h+Bfq9C15pmRJmzw9lFpFXb2pchgW60X19+vJSdX60+yvDA+5y6gKQQP5IIirJYlzJvZd
+z1dXsNFkM7RKloqJHO9Ud8xT+uUCSgO8by7lGC7BhNXJN4k6OWkvjpoqinC7BA6zZWapjA4XCl4
BF14700eS4rqto1O6Y/AZAFcVsqC6+VV2a338xroNYxhFecaSEYnhtE3GaK+Ue5Jue8cetso8KHS
mBVRdxkHAGniWJpraWIyZHH9gUdAoJgH2jNza7OjPqiAZ8McMb7/iZOnPEPF8C1w9goqqGNb4sAw
LNN+54/fRYWOZPqA/BH2YK0oaSNOW/V5hHxrcHoC433E48ToTrPHWKT0uAZdQqCZLG9sU9AAHslp
SBLUuUAEuL9+LmPAL6ResEskxhfMTycipopglJNSEagaJbkJQKj/tqW4sXKhHXwX5FxGf/ONXvBe
yD67YU1Y+XckL0Imij2Ar6lSQhPxfMxmpmohoe89ukLH/4gyWe/m4bicjkYdpZAsTx2Bj8nIwVTt
4jgkRHfi8w18h0GRqaImxNtX/ujRE48JrVmnyUCu8R/WcYKLbxsKmXWgGnjKIL59rBiNw1Z70QgP
5gswVWHU5KCGj8xctdtp+oSo0M1GENtX9Yf7y3ni1hmE3sAGS2pVJhXDR0gwB/oFUUsc8hNgOI6i
pfjU+EvaVdQwP4j8jpjneFIHSI/rXGG0vusJ8VqkS0rfntMugY2q02nN5jmGClhP8HSQ55FziXpV
eTn5qPX5uKhUiwb8Z+QeIxFdX0BOVNQEFJqVsF3Z9ZwS+ClXm03vniAzeHoR26PCfhS+yGPIvzC2
8rzo7edQyEDPN1cGnobTr8EvSGD+n5wHa6K7k73V+YM2XFIw5bLaDCSFxBSX/rH/yZB+IdrHINU/
dgenYrW5LK8Qsu1bc0xZXXzkRCEJ1USn8t38jNue33ekXUr79hxQtpDVJvzYt3g516EcEOD+Hpju
Q9WfJek3/4oP8lTPHD5GyyNRgpygkyJ3C+twANsdt5MnAmGsqZGEWL4VRbyFVpQyR2LtPgAGO+GB
GlyJyXLxRDwwKhpafzXkB2J26YeN5t1LNRCxiXUVnePk0WyxglADuZzZfZIZTWuEBF9YaxLX7Yas
+pxRm1s64+BGPdVwbmqSGelOBnKY6zXbtGTvFAKSUHKjJ+LYDyplL9HXAM6Ex++NeoSnolhcSw72
5ML7ArJAumkHWG4iL0COSOHJOcLlrIhwZ5xrr9N47VchcNq9vwMYKcBVLfpX4OkUT5yF97smsBno
fi0R7cM/kT4iz8B+5nt509ASE0RHupIBE/4FFcjDlK4WejRhzbbvfQ845gVEgL3ZZfCloJrc5lOd
n1EHe3JibXbe2+e5OeQ/oyvZ9CRx/+Lw31usc4wUpZp1Esz1erW9Zr2MJl6LepTLzuns7ff9VbEb
uReT8t3z0sWrtE2Y28XmIRbCOdySGFeJ0roGsRro6UNwKK7vZH4qa/4ZBmsDnxRVSjHZulEnKHj6
VEH/UUSkig9dpmV8boU80Iima9ncustYHA+cwHfNH5Nolo86+ijYOS5f1bCOfrxqwAXVf0AaUCPO
Ku4nUWl82j5H+OlnOGAsdtFw2bywvNJxFNUD6MNN741tsTJ6UZ9FkwJw8WNuowdDxvS+X6Vsw8/W
cfoWOOg+8VHWj2wqDoDOqjXTkZZ0K+sYBq09IyiP32bsbrTUCq5Te9aZ4i7PDoICfFS1zUunN+n6
aPvwwxPpBH6U9QO5HNgs/0A4h6rXFrsuHZAI6UqrGVNPLdr9BPFDeM4HD848wAwlNjcg2lw2RC5X
GrL4ELMlVjydM4SwqGsAo6zrR3Zf1ECtf8AYix+1XK00g9zpQrjZmu10MHqbkk1Qhoutz6Zvl2RX
7IiDDZI1rJgpvxld8T+q9qGVsAjGTTCj+a29jcxWSCzpAh1rqIhECXe9VLgMqpJ/kpsPwfC7aM44
g8MgmrGRkjHB34FD3kMDR53XWH1wLmvpJdFEEIQOtasCGn1eNy7/LnY4HOevAMCnFVQQFQHG6Ems
fIF9JXW+sDd1R09YbVEl3RHFy1euc6t6GfCP5TvvK7F7Xt1fb9vUa+qBMZH1gcBB0GB9cA9CVK5s
kjVxbIAzZpWnoT0JsXVEbibLIGfL2v29rq8JFleMyszIE81YBWmrENhYRwHXga4b22vRLdWv/hfX
6hgBUwerlAcHYM/oa8iZc6XU2wTJy4q1qnEdvOksQubUgW9dEsna29LTjaJjMnk/KwqOAgo1VGoJ
Ar6MODGLGExKaJaVKXr/fhF8q9NteWOjRjvex6niPiVzxxm/o9r4jzNo6IsQ4UbxHEfVldA0kp7A
R9Mpt+Y14p6YcsZ6SIbJU+zZ/iymapoAh7Z1UYGOHZ1rhvbl3gL1UCO3JbdhLhCgHZ6+XH3Pp7sG
/XpjMF6mjwm/y9jo7p9fNYy40WvCrHAyvAjAjeE9aadSk+WaxFR1bWUJkKNKGqKTWlu7oaCB0bfL
XiaNC+UV3ZjpP8HqVdl/Gox2d7Ctqdqso8rIsO88tK/r5B0EOMiErzhnQQGpnH5718D+iFtqjQUq
rB1L6U4wSLfImZqjwRO5aAVrQBLvwKE3H71/qAKeXw2NfL+qOMoctUYBlLUYEMmGZk4RRPIOXIaw
7WkJSJqJwHarVsOSebVXKoIVYO7iHZKrm8NcdiQxC8iOYD2IaZVMOyRWBVWmdWnf8pemYG93V1UH
Kki6IVr7g9UQcug4vIDZFEDDblYxANS9AnniBROoXvZVGd2SW6erjcjVr0Ci11T4QxVmtOd0jihV
uPRRIKAqYsD74UT8Nq8Dcsz5n/h4HIBBeVR/4+oxgIrtChC3iVsiuPqZ5W28foi6TNoNqaYJAVzZ
uAmn4zRuJhzVLco4EMUGHJ5arprqMJw63MSubDvbaeAyuOOrxIJxJxXlkucDvy2ia5r7wwG9X2QV
Vj1aYr3wrJJua01PxFfytWs7HpnMGtT3rAW4UaVpOGKiBYxVpH45tO/dGvQxF4UDzGAFp1boS/+5
/3ZLN4UBgSGYC35/9DmQ9fLcrS4OfDMMUr7YuKfSlDn4nFxczRkeNEBpphUX9z4UWFFCW9WcUPyO
42eOAqNoV5oJsVjV0EvcGoZ86URRw64HP9vuUIYsY7FGskyl+YhjFJI/WgNNd+uv5XyCuuHHikwI
WBt1MGNiQRgajtdZJ37/Z6lMJ9FY8CVqkdkkDY854HyO86IR5mW1E5F+Di80dD2PYx87gNRmzEwb
X47PwYm6uI9kf+Q+afnj38KDWZJ+WV88SD2T7KjgYuDIZPmtoAcK1KGX14f4dBOhP1LXuOeXQjbf
8mbXxp4e5EG6tvML/8ilMez4WGe7DQJYpRZtEvBluJGxvpMMm5YtTG1NC6Ks8fB6y9G3AnaxR5YG
AJOT7b2P00q9pPgnx/oiDn+HhcvW/qwisbHxBT0VHzgads76oaaXw8Lfh+quBLp5woXrZnLvH3rR
MtTW+R83CYA7TUT79lByzYEgxgjy65McSguawrH5mw923wpUdFs0EwRWg68IB/20p1LmhbAYJDWu
uquoymgqSOogEmYaj76zZY7/df1WjVXHTFkd7AYBbfKlCcy2InzpQeWgVvRFCf0WKqv55RdaEOtl
mZnEoiaYJ3w5UNMJFGogTt0VUuYW/mi8lL1Y4HYA3yuM+3dRSh90+pXtKp21I+J8qSqM71YxT1Lt
VYg0NAW/Gp5mSw1WFa36Qc1zYBZ7kxUarmF+HohLrYrwAWt2R9h8IfIOn4Nxg2Ha3oOIFPrSn0F/
t/JKahtDBhmvoj0GTDFjNn0RJiqcbZCWEeilS9ZMjKvqZKTzBuXCc17Vqtyb37XvA/nIa7GCRThb
vIAcQYKkYvFVfmmfaeCcUsUOwRFPAEI3aRdhAWKK26eVUepkDJ1sqHLWhJz7oLapXyEZEQ4CEPbF
U54A9dTkBDbOW9rTCs5uktlrxaQCFzIFjzHiaSucwkgIsrqtHJ26FuKfk7U84YbHWXCM81AVmyQj
KSFurlVlOdX0UbrJNN6JRXifeZDjP12noBraEYxys7Oem0t8BU715CkwaWnVXV3CvtoFH/Ztpks+
09R9bV2jQwPxyjpLMhdiUCAcb+CM25SedhZzzg/LcMle1JX7XrmKMl1HnkMx7xuamJdpAXW2hCtZ
oInGaJunb9lU1+kmWzQAFbdr8TLJkooI9WDqjTYI+11woh3+DtSlQtxc3m8XjKk8SdlsanMOtSMa
KFZ74FyBCq1DVM59p25jFLitsJUNEKe1Dx20zHbQNGfmzS7yjKS70/Zu4/Of2/JJGRsQrn1C3zvW
a/osMkrbrzcxNNRRlWXfOyJLg8eG/Vws5/1nMva7MZ3CFlQKwgTiIfXRLRp800KGFM5cjdtydC+d
+S6hvOKkRMctOJazQGE+EJRfValHvDzniQiRzUH1RzlN+ybKqwLFY3Zfcy3GBEBVPJdS0e5gM4UV
TJsmYpt+qoufMX+mqp3QhH0+ktMxFhrx4JbdR2gY8k4kvzLGL34xcO/Oy6g0hB3KgHrDpy61+eFj
VW6iD+lWqf5Yi9pkC5ezIhsGuERyVIgeFFU85vtaToixXxaVLBdlwGcuekKpVbImL4M7JREE8LyJ
0K9Ysr7pIH6gyo5NZre6+wZfAivuhQ3YWv0iwtPQVpDIvL1KyMV3as92dUtFoVjnjxnDSI42EmAM
JijYx6fCE9rZkifBp2TWAeFs4XzAuJ1D0k14wsKNV6HDKdvlJogOA90YA9XdMa56/uRe+K7DJMTc
HFweu2NQyAredGlUGE7FiSL3QY9RhaNsZOjnUVDfZgyplcy4XATLcWuQ7PnaozWiBMY5n3yI+GF0
76lTgpGom5H+ouPDPvutUGlsUuGFkl+o5+Uk2n1R8+P4guWzXVsxk80AK8YPwLhR5j4JzI5sed69
kUZXIJhrwfDaJ2V/4L7HP5N+ysQ3J7L5onIpHvFBvAwjK3U5shUZhCdS5IB59MgwrKcyxmaptU3S
PjtFelaOPaP7Ze96rjsTMZ4Mh+v1trdy4g1c4ItuUMW2Kap34LLC2G7V9EPjN/WilqYFrRxS13Fz
1Jy0YLS/iRDQUwuQGrY65YE72Kw3C3WAsnYgy19wHVrfhUfLiWxbz/cqNwnt7E1SZ5wEomVTGt4L
EfMAufRCB4RYsSHQFP/ShGf2/yrxgX1onpGQmbbiyMsJ524tN2vtEEge6J9AbdqhG26C4SprXklA
4rx8ct+8e8UfQSwrBa8UxiQbCWsUL5dxLu2TMmzJyb0FODP8IR3x/I939bDxjW7wvDolEnvdvttF
pglvuNB4Y8ECkHJGvx9ca+V7IepSDxleWjFBVMjPMi7lDMKwNJHPCyaphZtVNKVtPf2Hwz/zjrsL
ViWluhR3BXWlI0c4zqHvuvd9Xoa6LxddMhXEzUkdvApRfKsPWpVFahwFEHsqGRcQbeENewKHcUe3
OUyF6NTXWgj2lnwcI/H93F9pUJl/NzQMNVdpYwso/9tue+01bYpLvcIZIvkfq51xCOMnhREt96fJ
QfG/Xa8DDUzLouWlSPsXiv3iCCS0IlNFKGEKSS++TTVSAop3/KizK8OtXTOGaXLZJ9b8gifWMxjl
X1igcMmufm3E7KM6ZgXD7lteMZWxMGyFKZJIN8adCt8W+gupUBP5QywQhmYOSd6nzJmjMXG2l8qc
+j5DlsSJnZPYA2aAC0XNQ9+LsYkknj2RHPRwY4hRzYZirLSg2SFd6qHqlw8VIrN/C7yQyBW/wfe0
A1V6km1V2Gfou9JnrZAzmUqUA2QsJtjOjGBpdXe0pGAN7ZkxXxWSDVEsY+ZR3ggtBFuQI4pzc/h9
HrjcSYTdK4/0f2ecS9dO3GHzx9kAnEtRlnJpXf3rMiCGEFZdeR1AwM2QdfFL3r0p+d7G2T0K5WGF
fNRbU1/gLXxLw6qk+uuOfIlvV7gKXUTh3y1JmGYqwEI9QR+0fv7//453GNUgm5RitVlSRdccyz3V
Tz4iHhmk7vv2lJjojvUgIAtMHzEVJgYECksXzuw6PrDQuGvzdMKOTHMjM/ivgN3CpzFtzlBHRuNM
lHgdPXatiAv9FKNuIp1LAkE+Pjg1EZOtiBpt6pBNImdjzy7eVnOq22yBgtBXfPqWP3WMoRzcX9/2
q7/YQ0NBBbpqRGcJA0RLMGCKbRR/hdQcEfK9ccppoxq5y+m7wtHjb04KfgLH4My1RpUSqA9sDn7x
who8UxmsaGqE6cIjEplNG43xbhcCFochXjNhY6HZbtyLSFRc3cVb0ooJKDjiM42p0WB9aulzt6ZC
xreq8Cvs0OvCUZHND6X+Zxykx66pHRVpQ8GEO5fHwFX6Js8JWTKAfBYBe2KPCOY4JZ9whZM11Wxd
IUhD7O4cJjKmj6njdHbEOmBV/smjptjz5mfkLO1RXF3vnbn/SRRZiS5ulaHRfC1U2iQJsCVqYV6r
eJMxo+RHKVOitOu5oJFaHheuTlYlQR+fNcIsMvNMN/P3MqlYiEVXKgzykLutUE0QOxu/onfQmufk
7n5rQ5V5rFxFHuY6YYpqlbuNrjtS6sv85QB5c2KU4C9StKhrwcyDNro79UH5stnv7ws3xmwB+mmI
au7MQkr0c3/3ZI/4+zu7PG6Bp5f+PgRh/e8+ZAKL26gzdGlS2IejyCECAmkAcV0lFYV3/mU48dCy
BW3zgVTl17ppMAdfI5lnS/oTimUQqguEiVHCLuunPIUcSpucHMymd1ls8jbB7TJyyqndqjRoi/7f
TL9Yj+vrfCXJkvbkBzPKEKx0mHwLZr7TLXQFnPxXpTYpL5MmbMZ1sV4sU4c1Iif18UWri03qW3an
Ndj6EcOXllKVT6n6GSlE/tjqRG38SvSzWigYBSL232WyT8Z9bhTFUJWiZVS2qQ1yuLHrU2+a4McU
semWpxQw2r0gkYyjcMjH/YDvFXa4aOksbBjo2PEzBCt1G/wldrWfFLMuMR0ZSPCQqlwOhgbje70s
daiqExAJ28noHMqZnToezQ1Hm/zW1Pmq8peWgYNrY9P0H0ptmCcA0whAFtwKAIcZeM1hKo0EdeL8
1fgXWfxGbmIUvrv/0kxh9eoKdw3kq2/wuEvfiuXhG7hVygqpzNPyEi7zq07eAWYaqVfdZHVMgBiH
T7cvjI7FHpW3TBEWOiM9k3zwwq0BIeO//NaLcIU674jyHnenH47yY98koQSj2VALophdY2BKViFl
S7NQF7cEUR5Zkc6DBu7SNY5+ueqHlCmMcf/9oOc8SMWVqkz8lN35gTIM08/do10dh9gou+5vb1WF
siiFiW5zd8meMnrpVwalG6dEnU5t3fiTi9D99cYVPwIIbm5QbzUtvmj2Ytpk7fgrf26BMW4lDquv
gzl07guCHGuleRzj4IyTZJP1Nbjv0dVyvXGfaCdVXQynqKziWIOj8Qg9YUapBY/7cRXpgemJr0Vl
fWSruaj9Y9blBISBV/0BzYSosbowE354+LJJb3X6rwEGPBR91maxg473GMG6maV4GX/JaKbxycDO
GdgHLVCuyrM0t0UHEn03sDGp9iM+Mx/81MPzI/044taAe7swXKidQrjUt5WeHCvfySOjio2UcgSS
OvVpEM2af5AT1xJg4FaTPFbpKU+Viiq9kj/B7hbmqpDCHG9b9abLVjPCKoIj56S4dWGOoUZ9xwxw
CmWGLeyje8qcvp/jcmnS1yZrV8vVTz+5G7LGYq/OijPDzMNbi31ir7+8QU856PQALmome2Ewfa1m
h9n7XhDhb+vF62pT0dtXrb78IlaIPyZEQ8Msks4k4UiTT29h/ez35+E0c6JLPJrPEXsSFQHAT7zq
NFUXA3MYtYqhjl1kgYShIOgGMGurzbYGEaH9NopsSwVgJB7cUyPjKG9msw0RiuK9ZcbIwZd5O8aF
acmNOyCECTjk0uFQruqyQUGW3bFO8aVOcv4qKIFXXjQxd2ion4em0PXYcd/OfsvCsvjfj24O6GIu
NOKjdTm2N3m3fT3Voa7BkrxnyzjVj98wUFIvZ+pIFuWyu8tTfBvHZoEpZ3jk0Et0xJnO0v3yDzTb
CeNv1z6N2gMa6+Yo2kZ8zKZwXZ2wgDl/L50B3YCd/6L0d0WtOC16DIbfDHVIiZZt5xwbuaK/Sa6I
kPhHSpP9J9uRwnLGTXL7zdtzgqHCiwkEQVHhCO7l7vWneLzLWo0lgD0GGzoV2ZXOI3Z9HOIUIcK5
IUXm8kb22bSe/ZZY4x0osxtj8ITSFFCvs46JAgMcDApilQcwlRqRB9yrSei0NntDD16h5d+tIosu
NqLUj26mq5EmZof3Ymjgg7fdkygNswQ3KRvZ53QmNo9UwqscQ9g8BDKdH5+AlBsKHpUu5gSCd0kO
25Urjpmk8suzmp0CAJavonq3/76Baf9vIL1+siRGDXylRopypR6Ne1hQ/Ecc5fcYeVimDaRqJ6wD
eCeoTl64c/8ynqHrSK50N/2N5LW58Kel9zrJW6rB/+a3WB24SvZ/+pJc5WlEk1CLPg7JldWccggE
d7VTt+qDuEa3CeDyviJjLMiefHAHibZWbitKCYxewoS4+4YET0jjny5/JzyxCJ5rhZuKg6Fcj3Bd
W4sNIGKzzd8RRsds/HFfwvrs9JAGMm9Dm396jDxRUZ8aV6vZQ7I+VgnXT98NhnNWQ5vAEQdX6Rgs
jNJtmqVbZUsau9aP0RDvIg88M0DOSF6vcyvDlu4B4ZLSwW0u4roolz4K2Fop+ZIuinCi3rFKov0j
QjVOYSf3NFYnrmpbS1XhqzWMDTqOWNVIJ68ChdVC4P+3GeXw5wBGNo+6eSq9gyQgrj0a1tZ1OdZi
9wWG1Ao9oUrnCOqw6Sght+bkn9w6+wytck19NbtWJCzxgOQi7KxIVczXdzGA7UbLTeS7PHGJ9FAz
w9vS356L4/qP1iWcRYJ9Oya0gFpxe0l+hNVadmh2MrTCJdD/Rhs067c7wdiGq6Ly9IUeCy/rONEV
kCO1wXgzM3wmFoPNNfHJiSC1U4uqVtLHv4oJrtkcXX/oEWyKklUWc6Xtvkj+d6xiIDoaGIoIH1Rt
eX+jNDsxcTbWRCh73PkHPpObcDPZPjOnCTPFBnv1TjwjDmhCq9vyAO5m8KqoNDXW8rATdOQiKhia
pJWkaSUCyHVhhGW9Oy8R0m8wwaIeT3I54mPnxKrVAe1mmTdcg/3x6yTSxiFrmIzLKIdN5uOPPQ1B
CIRqkuWG0cG6DZstK6/HyM8rSEQWUsh5OM/GCYM0ebmSyAzonrakCGlR1bkFaOG6ozsO9oVFusqH
qdstdAMkBsRq1eRXWhpQNjZjHTCREX+kPeDg8GQd4ZEkRcLnxUQEH2MCZ10Ox+AbCMDrDbakZ5g4
/uw44x/HPxIPOp5geu2LePtCz60gQ4yX7bBwBgXo7OlVI/El3CXVkHc02EOFf/KIVRt+o/gFSwBe
EvGbkGpzwnDNQ86+OmUoUzwk+Y47tfqGn//D4y3cqcrIfjtVycC4JxjkkFgzEercUbAUu2H5aCo3
bkstRo2c52nNXtJRFpPRMgRfZJWRLMIKZi9R58j0vwv6HQPwq6xHd5nf5o6Xb5Cmh9GJgVt6N4ry
pWTEm6wDfZmDBYrwYOVEFXyysGeEPousTWkzHoqzhXjZ3PQAWhkbyHn5g2kfRXTXwy2gS6N+4YA7
rGJgt/Aa3OudXwCgb4NeUyM6hBv5Mkqly21tn2dv1WJ4Kb6sJ5FkapbDC9M1X8WzZcFZf9cQHfD/
RTHGScBoTeCuCbnVoh9p5axwhqpMyZdAUwo0ZMl2Z6K48xJEfptQtRNl+rAFaIZHtKOFABA2gtuR
g18a1c+aRYVNwovqq0VatwvAEzsEiVIrdaDL0IUZQFBDBTr/UGMvP3nGdVQSxp1wXfHCerR9KwWK
m4psxfnzrcdDQBUxcn6ir9PbORgHApGHYC6hzWwADVs4+uyhpn8/FP8HeXhZ4k1bFEDOELeXmp2m
5VYYFAQHqLrG7nzFi5mks9mjks2O2AjD1f3gGEK6kSw+1aNDWkgg7fbyahpHSlwzMfdM34Aot4I3
+zM24MLZSFqL4f8YNHAo0Pk7C6e6Q4gm+TIKouPgnFWftr1lDG9yST5f/Hdj5gtq1IXiJS2sryUF
LKJGGtUl/mZgRo+/2DZs3392eonrEVR12r+zYGrL7ajRNEOsl4maW8GczgL8Qzk2eILaLlkrMN3p
DUK6rQ2XH7rvEDjy8X7/U0OfGQKi/1ZMMrkrnd95iG0mKdZSnXdCpSXqESibA2cO2AjSxaWK+4XJ
yas4ciWU/DmzTD+sOsVlJgqOP0Iu1/IiNecreTrEX3n1+8W3zN5wEZm/0/lWirVdLnrnR1Y5TU33
0wfZzNSAnwS9ARXolZVWjADuyp3YewTuDp2QRLdSwcGwMa5in/wvRddpckdRf+GgW4lzxQou6fT+
3uDBudecjfsXrJhUX51DLQQglC3vAGkmqb1T3LG8x8a0bpzsVOdkd3ytvCN2jb+5j4xVOCrtg9JS
Bt1lhZm8xmKXk6e3mjSp+lCwQ6XAzA88naPvsp5rN2Q+m5J4zMzLU1dWTLeVAYrmSCLlsz9o1Sv2
SvHOL/2EVB0+5yasn7buL+fCLkbgisg7d6Fu6kF4mQM0HXWHqsldwcZB2oeonOk08Y5cfET1pSgh
itUa/2LmPU3smzh+aXxYziqwnDhBDMzSEK2UynKKqx6uC7HHdHOSeBvYSDiVc9dR9p7iTdxeNbdF
mxGaSU2dtoy3kH7gK9/U/VvD/LevXxAx0MhDOx5ALBo86ZdCn+yVtHIiSSaj/oLEUXptF4xiCI9k
Di7xsr6rC3GELdnNirDHwX0ONIkR7F0u1FMr0fg2YLnML74D5KN1ZtkNy4quO/sJqqjSwoLwy3WR
uwlWJ5WkWCJTm8WnMAHJIgav8k9N59zKI9ANHjKeHQhS90iAdbGydpAaUzfvlPekgTz8dD7fJLSH
4LOydHAuDb+yJX68OYMtPBhmXlV5MVcbvYF8cHYK96vm+9UBpT/3lANKiAUYTqZjlYHPfQNTVBKV
13q0LyV6+2c3ITn55DZSxWAPAVvAqujm76yJxT4hqZwz/2+wNnM9XLkn2NC9A6xvjiTlSKcSEMeD
wung3XIC3FwNU6aC015WnSCS+wpX7xMD7Wz1PFfyC2S3cRcQ871b/bu7wTDZmtXTcShfpaYdIm/N
eOoByW2MuM3/xxJ7OxkwOrGVn1/3sW/t1GD7jm7dxrbcmeb/BXqPV50eW1gDff5oBBRfVv6lzBGE
nUBuHFNokIL7gdVu0Cvb+bdKbw1Zu62exnUGpmWQRd9HzNNHN9d6/bJ1GR7K29aOp9Xsm1U4WMwa
5JzT2qgghXpszVXDfmjyvvPLCszgWYozu/LsoFPzvTVZpTISgfhaFvaKDCYNV21AfRP3x/PGaodg
JWCk6C+VbfokS/rAtysxD6b8Stzre6eeRulvJNaLhcs7V51XMkluLWQ6wINNvc0ebVzDIaP9teND
hm14CEsDhkSEVDOqFRXcfVDL4y83PCeKYMAaWnyWdlJaDAbJl7X10tPi45kOQrgp56ZpcTUq+lfO
k8Dsh/mfvRO9lE5Ij1w9Umbx6MZwfvvS9HjQoo7IrhZnMzPnzauMhucFspDYDpUem/Vy5V22aEM0
4RD75Fo500Ia26HDR4zZj8r16/CzPuSniRYoj89wd2YF38gYEDieLWtg3s6Pf4fj9I0FM0ZzPXGU
jGeTRsvSqyEmIBb2g+syq75zmal9oZcj6sNOJzzb1l+P6cfZBpimAfIWgXHgJI5aa1YIJjGnw19H
hvEeAnuGdjyFDhHaUafVsrlp97l5jP9S5B0LDZbRe5YqoAQrdKhnCXCIlpNp1jw/hM256Bc7Wjwo
EEaiUUF39ZTomtWwbORFNIW64NYLFFmLi9B1hN0sCcoeWZaYMzdm6lsu45d/3WTRPEatei4D50hT
AYh94Pxb0tgW9qWhTsU4xMuTgvfw0Cjqpf/ZVhBdxaJBT7DJ+BfaSvr15ZvPchQWiqe9dqnzYjwQ
lYP4m94L4yOqDutfmEWeXFZXVeoKYz2fBwI0I74a3K75kFDrwPGqt3f/tbTzEAWZM1zb8wiEM3us
gH9DE1r4eNMvuewfHhVlk2EdcjR19UUYGv6lRq+UeICAnXwYeO0DlcBPG0YCjYJgymKoiO7EARF5
iXFpqIg1UOghzsMN3NZqSGtDifMKHLCUPoY4eAWjmXSx/mm4MDPiQU4H3yBqv2UVOE7EnEZenkaw
i+kU3RUSRuJKvnyMWMlozrnKLCZ7fKr3f+Q8p8EUPxhdZabn8xsU8c4efcd5Ux4CDBHCXbBETPtL
QwEyn7YXSGez1j45N4pRpeT5Cux/pRckZxJrWy4fN+xaLAzBm0x4TFnJ8ltgWYEwPlPWidrGecz2
XEUJJ+Pqnsu+coCbS3ZPqbvjwhgqDXlji5bzlWzYTU5qee+A5jb0sjd2A3q8/IOvBK0SA19Gocxe
x3AS72qrTjbsMuSi7gctG4TRaNKzA/KDOCt9XnK72DwtwwEv4Rq3uIxjFtStBZwGVNMEAlwDysc/
OM7QtrtbrleONNDh5OlQWsErpR0FmA/mM1mq8d7HcOE/TsYI4GuZdYEl/tAAeX7lRqaIMjaAI2rN
jiTye2XACiVfVj+XD88q2x+Tj8ZYdSg2LWZdBjox57GZQq+ZkOL40aX6pbxpG9EUVvTt3CTYgP1u
0cBfh4qjjilnh4GbBSnuTeN/FpRoUp0jBFiJf1MIhWVtowUHw6yZk33CEIqIwZPQK68GvDmLQ4fK
56vP/O+aIDMQvgRxJKdfSv9qxb2ysN+6yx/UUQN+kNSqmTpyCezrOQtsweFnslBLJXQYDOJ6OsdO
vtGHtHs2eDjTbyoNlSrkv0xi5t7N+VYntr7AywMz3Bvl6p83lKXKo4ILe3OAEL0nPAek6aHb96aA
v1xpRYYh+6xOQMs88BwUPtKc0J3XLpEQ7uVjMIVQEg86L7RaPRGNx86HvWP3zCvveil5XwbTkmuE
aAHONgEkdp0FU9O4t2SsWbdar9ZXSSzjuUobTPk2yOVL1XoAt0ARuT3STe0HTrJQmHCB/K9JG34B
c6FmP1IQBlJXzShWJCZCqsLfQGG9yfVpduTZg20gf5xH4ukubcG56gpKHLvJhP5Iu9ngpiCzLSx+
Y5V25NKqdvFmyxw2MeD0ubvoAEIbziad4CV2nXRYRO4S93p5qPRtVUc3prg/1rqU57kqBT+02z48
+FB5aUfsFmpGwgdYw0ASDG5vd1u5cqBjJDf4PbDYQf6nkDT31EIrphbTnfMet3SB4I1b24AjxV1J
SaV0WkiEGtddh/vGrgzlrGB53bsLI9YNdcK8n6sIuB6WxtjuIhQCSpQkl/CkrGznkJTOXln2pxIO
bKErSn3eEE/ty+IFIiMLdDXhYhN06uDzah535pbNyGQdSMqoI8Mg2pg23OYByyf2v7i6FGxfsHEL
B8yAX/u26pxyv2T3IEAqgDgAhyEtf/TX5mqL/tC+XlfyL6V+bWtNMd1y9xd7JVOQIjw8gvVRrncz
Sx9sqG/5geMnkUv6LA5MeFkgMZrb7jAnvoJE6dyCjWtqZBRcUNRUrsQKlFuIHpNXDMT/YGIOKSsm
wWCeLzddNTGFb/ImOQ25jF8uJwHHjh0el4DImlv00ko1lu8utPmfsDdkt656RoehBOPnIH3AU0wI
aHYjacMBNA+fVbXAXE6KnbREuBxqVpy4MIBA8/yfumjjaPKWknrhLE0QuoVh9QjOTfZQYTghrnUK
th6TGJroMSfxbpLjYn35Iz9vgLzR/Eg3ELXBC4cBWSQTrXUL3GpVZmmiQPQbrtxN2cmY7f6N4/2o
cIZ5tB44R+8bjDMaXARwq/gnTfgchGEjD3tSQtYU+qV6BxzkihvfcE7Qc6E3mSt2L38xUyQv7ZwH
Q3O9kxn3/5va/YKJul9DalxmjJ5sxJRsBKVrT2esIYAL0HT8r/juTdn//5F6T4fM41UnbeJZWfyd
AHHm+tQpWRFvMyanurFAMVwbXrzxhihRjD8J6MzkpOF6vZDoYaRU1oiEz6xeG9B9ODFYeIvyCh3d
tXKcJIIOS+drm8nEKY8GwGmhFelJRGi/0nimJm0Z9TYq0EhlD/5otNWCYj1/rG3JxSCwenojR4eE
lneibum3j+mv7Evd6HePl9a/YRBSCifqTUq7npxeL5Juziss0NT8XQPOQtZupLUj3YS/4U5sRTqe
IDbyr8lkTmbLxKxBVVIe+G96GJivYv/YELy5/chgDEvhWvwui1dRAK0CiSbHZXjbwn8ffr/g/YN6
Sb0za7ozT04mf0rs+tmyxMG3DNGskwCjdnbHZYVAxrg8B1a4Elp+zOng30DtTZ91V7SyEdu1EAK1
wLrgIFv5QsA0HQEtXaGGAK7Of5jgWMo3CynXWj0zNbq3DhJJj83gCLtFk/QOYM4MRzmtV9wENlkk
lUglVJKKoykUt/On89qgLPMLhQw6Baam6Dja48nyjkoCbpHl1yFynMLOaW3kAXJLUsq4bzP9qaCO
akyjIprlSlqGXvnzD3Br/SiJgnXfLXqhCUKRAKlSjw9OqjGuF3R1Ohv6FnpJ543x77DsLRkBMSRC
1guGG8tTk6tyF7SJ+7hWfI3iWdTydcTqhB9ajVWF9T1ebnd8wdMW7N+ES8+bvQ5SyspODXCmPbVU
1SHk+uU/JR0JktDtZcx2GRYoPKDcgcu/ECaQdr7VetVQwXOI+BAchcPPy7INzOG9DQ8ZFxI+tuDc
Bdp4img+iWOmKaw4WI5xgm/AGsRBnEsbrnZ/+ar+G8vJQzRZ4BIEsL/Py1mGxU+gtHsNYF+2LZ8i
u5B/QdwtNUCUA83tMEF6sWAs1fQlqmmUaQN4XqFBmo3mP7oqx9aeIBlCSn4Oit3gqTurBaPlkNk2
gQpxQzmv8ugW5FLKJ9JH/5EjX9rTWOVbYwmian/rzSOeY05nSjBosHubVxc0Z2J9Soghe2XEkqws
hbp8SCRyOa+AQ5NkcW+X8MJsy6cT0GTo3zYYFI7G2/AxomyaPBmhtOKKwUX5VO48nEJPDBbQ2duS
yDLSkPomzV4HsKbwGmBnTzmYsY4l8kAXsWkUipmdcij1JQKSESiDjYTaWQHZFCnqerrl8z4Q052n
rwh+nc8melTyf7lFIGXy9LpZuFFuHF103NF1kJpDWk0AaTdueHTMhf/5ODtlXR8U32M8aIPUyO8W
fNcRmWbZjVksYA+4VZWV1kxMzrEyd+DHR0b/jq3GugJzkayieGRK41Qw+sN9FSTshsx8ltK+wqlr
e6HgRCzE+0bjxohgKMeHUd0TStBBdlD7SdL4fjPMEKRxiEevZyJ2a+t+UpD3i8kLlRuDS86biuUK
lVFrwQMdBDhkYChYwpK99Ar7Xih/iJXKbwsJnK5/X1OE+Gu+ISxo5it9FZEZwR6nVg83ZiytDJBM
zGjsCA6POI+zAFRnKMf7NsQyP0T/G1Yfj830Iginl9cFOr//HR/3D7rMtCJTX6UqZSSeuZtNT1Xz
AsZkor+Fbz2o7YP/CkoM3nS8hrEEKqb8xMCApGFPZ8DivtyDnb6KKQUMDfpaUmJhdt+zoT3a4Qf+
jjebBGELzU/krb7IP2mD+WARfbnLhly+3mVVn5oMIt4lIc/mtJR6SfyQBpCDnnw6H+mww3lxWEJJ
L0PMgK9L91MRTn5UBX2ONYp6e57/O6sdJHfDj5pQ0JnyDbPh3cORGdi2rDx7quk/JwEyAa6IBH56
ORmDIEsW868sJJrtJ0G75C/4Gv/MtcyoqbbYpCTpeyDHmmoZnDVNR0hppoXcuD5YbjDvb3CEh5xx
yDLw7q19gTgOKRIKRR+Ex+trNF0WS4+0HsfiTMNj8xVEC4P0KB65COPDw2U5yXSotqNgC6u2stdb
P5akVa9/qp0S3z2qJoZ/mLLlpLVTDd7gJ+0Vv8BaLjzY4aEP628sd3yplMgjxIlBa+wkgGaOUJRT
B/k9xi/1RsP8IEg11B5VT9LzSYx2OntTWJg2uCy4uBrwcWngm5sXOfQBgcHOiCNV1r28U+wGVMZ4
tLlyM/QiU6JHZLFZJr1pxuHy7GHWJ8H7lQ0Vm5TQ7ESYQ2Mu5g+jaHdTsALEaeVFPn3nPrSalRGT
GTf0ZC1wOg6p4yblwHX71tbnvDKo8Jng29/Y2J5v5I9/U+wMD+um0EXZSSTnJ5VcYUR9a7+/2SfZ
4/BW7Cby21A9rTnniip0dbNCrA6n387MRh0y8GaHqBWdDoKMzgr9DMxfA1AA4KB+ioCjWkEiQFeP
D8k5a3BLTngsw6cpw5THOvSW9HOnaRldA57axN0aALUrAraM8VrunTnZTAuiXfjwTSDbETZEVU7G
5XmabMVAv1xHIKFK7JonKPIkwpL3BnCzLsGyVsK7wHthcHJbJZHiiE85FIEYbb5NnVaSfG9yQnsd
U2I/aeeGwHg17JZo8wDQO8lZatylVpti19xUe6shnstQFHbkrsbdEx3sgDLQqRsGBHCAvkQwE+FQ
QzRWjtvPTKo0hpjp60+cfyjSGckMw4FAxusOrSAeBGXK35KWgrehTTbjEocdcJtyHG57kxYU/+eS
YABnJYulmd5mIbCl1ubPuj/hNPYcPP5aGdsgQVxgM72e911NoJbYLjVXp5S45LmlcAPSwidJpvFz
SDjsq2DwoniwFhphFVRKhS+mxhaun5+U6VtAiMrAzOn4rSkOdYxF9pqpKHAoFsakj5HsspKWRCGZ
DnTJkb0sYIkVJBGnNRfp9B8yjXNJkWWUGr01GWIPOocd0dT6zfgSnTV6F96QN/1qFYeuqAnNWEmV
91isGPfJCLtZo+PVAFXrleL5cjS3Kbe7XLF4dvHylep4z/U8ATpRNhsBbFDEPDo0euhX9LkWYRHJ
CztJe7+xCRDNRs6WTb/89vwRWGzYRDE6y+v5C0/2exiDig1HqtAMeoChbXAZlkrv6Xt85Vz/ayKR
3tuqY5gsfdGlPzNqx3gywY48bGvoXLR0k2FBuUr+s0Z91kfZVVP9WSdm0E9LAMEGwqBrc5pk8buf
Wc6VXxXq2tOXM79aFhzburZh+D1t4+PqRfERXyFIXMeACPIMkzkG1ApCLv5zmbi7Eq0zuxVNPKJc
nnj9WWdBmbVSCOXlkiLFUL4edU35xF+IWyElezugZ/I6LWQDAdjxMkL3SiYPSPDDhdrqwLAHBs+X
0rRpow2EDMbfKeTv8yGGbYYwsnYWcna++0kCIdrmK9RXhSK7eo4PG93sSdwNxTVWEK7uufj2PZUn
vdK4JfM1mCX8FX/qt9OSeCu2LXVxLu8wP2IWqfCKplllrlone5Q/5Zk4TID21Wu7u/QelYpcIxZh
9WzGTsEfKC0CjRPDECzXiPZlRjLdCKKjuwTMDFaKhfEQo+Gx+QrJR9UZBOfIrbviFerBhFMVjvPk
XVlydmh/0wyewxcDZ+J87VOAaF2W2N8zk8cmruKEjUD5NTsoL9AetzzKPSNUv2p79KEW132fWU40
5Xjgo3Wx4JxCVOesS8WTAFTD0xmIqPQLSCwn5wOnZc11apzUODlv1arxRVniyfFrJXxIczOdikTh
S/XBuSeLWWeuKWn5nR3VaBa/oYFareEomA7YlMEGwb1wGtqsXraTL7iCZkFAn/Fbba4wBAz8febs
J5W369rfPTTIEf8EuUY40KrkYp+L3qrp0vPvCnuMRswUQj4GhRGIvSPq77LqlqQLUK8vrNelNmbS
VjrsIU7hTRbr2hjg3qe9aefWK+UDaNhqP8OkNaVtyvTYy6noZy9+xpmKyOOqBWgJzefOyr/twc9p
RZXH4o8VqoKW/QzZElnQaprpHtU8xo4U3319uh12PUwIBus/RSTytM/nL0+SOM7qdhCQdS04rvL5
BPGgAZg+ORQk5JBvMvLAb2+7RrHZLZ5zfalJYDngq8ovZfJ6JYzd7Q9tAbQQwNv5ZyKyHuYHLhe0
KgGshuUx6r6y0HcoQo0XlHrUilOcgEc0rxFSAwwfn8e03EkD4N7oPgBBCj14b3toKmi/IguyhhjL
2B9IKi6VHFgwOYBzkjTNPrm0s+Sd/GsR9e1MvsQRPaejKKMLQDNID0ia26rD3oKz6X/EG7i+b4ED
4V3B36SXfgxEp6j3Pu7Dhw+8AVldaPuFYluaCCjFAlH+UyJt6pgE0bqYH7u8z1nHKV7D8QzyDxXL
GlOnggrzBb7E+/DkE4KEVddCsh3c3Uq7yZLN/Oh896M+F9aNK3x0ULRf3HwmNnQVgvuZEs+dKJbO
2v1xnX4yXmzH1qALGEKufW/S20BUMmfhTcaB/nd7NpVAMxqUtW/I963AMP/15vnpnciwQYun8Hx7
DegJeOdoqT4JzV8oU2QNbo+GktyobQca49BmSyhQT88N59Q37oida3gZzwo9TDqyMYfWDHqe8brN
ypnkh+xNyjbHYIYZ3A0ZMGQ2to0J7HKR47bRVTHMMlqe1LcEo6Vzi9LqcanNRXBCTAxWmPv6XuKc
2W4DVs02zX4ZaFgPV/PkwhDnjuRmO7rq741tqwmjL9HAII9P76RvWWFCRFIJ2S5w5AcLUfAkMUjD
dheC7dIU9+oN0wvis1Ij4Th2qzYwNUJ5fEiefxjMrSs6/YvoD5Oyvy4HTt22zCI8DOTJwFWfiTlb
NlKVj76+ukI9WKl8r7ruyt4T7YdZ+fBVYb+jkDpk1C1bYcLagImk78McCGzhOHW36hkbWK/A8vfX
MjeucgZ4Umn1CQ7o/XmsTMS8mlsscVdDTLJselYu2PR78cBYAWPFPfpwFztE0sU4SLjQSkKtTWE0
AHHzt5wvj+1eRDsoC5JiD2a3sfYcYYXtXYe5aTDqSXsu+ZfmcvRie98tMZRnP1rn1wVCNTRnmlOR
YrvYUIH8WgjT2e81J6itTASdPWCF7rjLE53xYVokj1rk79wtPfLcT3qeANkhlwlJ08AfEp0A1DVa
qoFltQ2JMz1Vkjl3adKnZJZpKQED0l4JI7X+qFTmvpZHxRPwMk6FwLNBxBZTxcjqxatA/uLZ6hCp
r7W2NdFVKKVbqZVyF2ha3ZV8HPaSJKdgm19UP4asL0FuUnQ1jovim8LOd+X+vfPztbRDLUhVEf6h
JTX07tVPLAv637DGOhM41pYBxOjpY7lbxKbV0QjE0jzHiESB9XniFJTwUyFdKYQKE5lbvXOZfQ8V
D0unWLn7MlDLWrRJZO2bwYIU26zIvXV1rQnoY1QwnNSqCqYKQAQaK/SqffE3Pt5IvVMbQWakhggF
s8RaeSMUB4kuK5La0BQ9VcSF085Lhxq9LJFNnki7rnhmyt3/np6rIF7TbXu0to1IxTAiHQj4iDF/
yfFYELqJjKlJLthpj3xxkc0zOMX8TwyqK+lrksEv2q9ckawyQIzi/V1M+DZYBUI1yk7jR9UCKPKK
ysd35BiHxwEFqsapf3UX6S9ADl/BlHdN2/Za0KbIGeFO1TuSmgM5fbJX5RyPSuu13RGqulDMOvFl
kCneGz8mO/1wMV5inbiIxHMjnDa/Kbct8XloSpnzcCd/DOxv+W/Tm/9srls7wmwKzb1209bTSFRC
D5gCcw2cS/ElFUI83mQ3CFKoY88en/niDDOT2i20CBwKnf9Hun4XriRAVDERgCJNaixP4FD4Sbdk
aDo+JkAMfautwyCAONU4pKCG0IKzMQf3FXbJWq9NlJXnW9iO6+/QhtFwqCNXX18R2Lz1mMhbfSGi
govguJWpGWrZx8pUkGZjpZfUmuIGFTU1o6pcBK+RmSy7BBUZXFEPUvlwFBhc35iWGQwoI1JYdXQX
pyLw7MMYrGue8Gzb26mC/Em3OwSYMMYUL7Nbia/9aFEWBL0zKSwQwTA/yCmni4u0ANZRVI/voHuO
qRdXmDKJ0st2XYpQteveFH+ddA3oEeSciDghEmqCUXeTlruU7jIa8ntKy28VcgCBMHqiNC2L3d9b
pthNcn65EZ8nWHQAJaPKNpbv7xzpPD3scXGJjCyNtrn7BN3Y719IlR7MIMAu7G0lJj7b8+ktpANr
CqKPWR8hmmTE2qVwWPh2v3IsPEulAOYLf2Fi4oCuRTz1LgoPbTZX5pIiSvKZhocaPhKrLyMaTxmY
GQhStkjJVkbmVBX1HMW+tLK9bXCkQD+et4sv7gUxlZL7x8z/us6hnY0u1tWtOkkR7yHnZpGb8A0y
Z3KtETO5Rb3wSKdShIxv40JnaxokSvjhNcdBW++ztYI4WBTB/RNTR2Fews6prJqCFng+HRUmdFPI
A+UcyBZYElT+bv6yQ2FCJl8Ue1W7LmFt0smTUfsHDKevqJUqpD1P2zdyCj58gHb++s0zT4aNRZup
lj88eloUCloGXZ/3QtWBKFE23/tzJi+SFgbbuUUPIPaD/UfIqtONrIUxnJKj9tPKgAVTzi5Tz4z5
7uMKDGCtlFedeeC+omF5z+xy05GNsIagjzSzrYIaiyTuOyby/nSyMNmKP4fA0BJqoZeSTaLwkHOS
FG+e3bC/0Swx5kWnXbHTSNhoCOjx2j30QA1Xp+nokn6SD9ICs3evq/Jdm5LfgJuQwsbZ2/LohBdm
H3xhS9FPNfFxkzONBf4ghx0t50fVHdqpu/+b/pUjIaOMfoOBTZ02Ie03JQ2b9/OqkgOJd/CrMEgy
zCVdXtKdGlwZQECYLm+xgINWqHROCf/oZwtYTtNU1+FSZmLKpN3FvFb5x1fnSPlPfhR3qLCTE8WP
G2eXVBNZBCzITLxuQzWM3ZKmc4q6YJriwjmu/bWX0+6rZiQxwuOJZr06I9j8GbDGgQRQSrjkkyVA
uAdKe3YbVHCSbgRBUZgjZRCF8ZSNpZ9Duy1abjdLqbRibInokAb43l1Iqx3r96VkJDwwWDfpkwU4
so36RJ1EBJl+WZqc6425vkeMS2AA1AnXfcq3Z/QmKfjCurZwDrjdZI7I/K1Gb4xpqEWcEnj2stWR
9bb4+XWKiwKK4hn+lY0uX1zZkIg087mWtkCTG2wDX6IZmOvvbhR/lcPzKwDXvgfRrUxe1jdnMAjh
UJT/jgJDwH9xWm+g/s8r960h2i/c0sXK45y7IFBu8uEa7tMUDvNYoUMq0ipHr0+OrO2Y6mjFGdW+
SRPOWKGHTi/NWSyLOaEQMwvfrsR/Jc8TkrAm787ePvLpI54QLkBamkmE/kF7O9yjY7XHTCRjItSg
PrfFbCesUQiayTD01/VNsFaOOkJh7UZzu5jTo1H62Ig7xMBidNKP6bHVNTcVEkGRls4aBWJ++WOZ
FNou5qlT/2b+jtmkDJNhINkyLvILIEZak3mJ1zgggm7G/rcqsREyrOWWcJ+4efY3+j4zcTODnzeB
Ksi1gLM+R8LwFV/8FzxECnCkT6j2p7qmRLv4b675uGftudWP2y8k9PHZyaySyyIbq+s2GfsGCzzX
qFc22RBLeCxWFvlT1Yn8xRv8Xh24/YsI5JvSWoCce8i12ixmkfMleY+mwedbS3+sFNEGlc9OiFDP
iCJAZ7dSOljmroz+AmICsK2Q4NQyFw+hrEou+Ir8G0n9hidgxySZoYjqOHxJoFbZUGiJz81ErUeO
an8XY6D5Mtjs79RAivNolCXpmYHWsBuHaM5YHF9wQnmuTD0nrQhskYYOq+FNE9J1+tvTxnjKEVC6
HaEQrWdwaC6/KV6E3M1O6Uqj140JdAagvDoILYJ29lADLhRL2L9N1XosDezisjFX2IQfN1GCwiGE
NeKTIhXhO9KSFrr9M0EFUmG3n7WkkI5NoopojvZlUJeOfcHzRqDH5PfgoqXYdqa4PloaRarE10Qq
1nZqq/GifOLLcX/WXlv5/awyD5t5v2h/KuR2zbG4jkefag+LK1T6XXhePDFv9uYqFvYJhBxMmQwp
uevokk+M2QDGz0gE5o90hQL1Tj4bPmeoHtC/NfJuWITguiA4DcFtnnSBcZSk5EGMc/Ca8WweQwxt
9872u8NoUUMJQcDaVdIqSeOcrZHcnG6+k/03WggMxE9kuNOKRiywdM30arQvczm3wO3yQ2McgC7u
KQQIBWd36gBvZILqEcp7NE0IDJrOJ2/ErcqgUX+Mq29rgkuVFQMIY+O/imbyvFUU7OuTW9nFCCra
8k5zUBFaKZju/xCtJQY/BrFz2T6he3V+Y5BdrDvKditsjAQYk5C4UBVZe9iW4mn7S9B88x7sUmyz
5yrTM3JrqikqoLOCQm05+LqEpZ9Qq8qYxJ7TG9u/FtvwLK5Aqx60cW7MUzg0kyIj5cqLuz3OSvvf
9NLsvlfhqaUyurAxrMApjo3WXRBmaHWCzKPzztQ/zj78GsAsgF3ftv6rJsYqA2sdgKAEEQNH6olX
b37XFqy30TiJ6OxlRs8x41XL+yn0XeJ8kaZ0XlbDmhbhUKpQU+fxJHs58h9v+G1AaKEsViijWWtS
TrmG0LE/22zjzmoDTjvuLH8CdDCTxnfu6Vjqo9J1/aukVkDzZ74YJzDMC8jk9oVumaq1LGVy2xwK
1yk8mW3H9S1L66PGfyF/4WFQnGoP1LG6qV9TRaFNorPfXXfs230SMFhgrASVraM7prh+e7EIMlKz
/YUUqKp5g+XmcuAOXgPOTjLS9FxyWnSk0mcqQfPHsNTDx3r+J5dQDU5vmeJp6f8aWAbI9Wdy0Hal
fJnsWLqOzSQIXrKQ5o4HjesyOhN+5nKAflGthwEL4dpPJty7V5cWAO8klJcK/+2hXBV/HiK+mGvD
srbibRLSePdVsbxQPCl+0tjJllN3SUTrEIG5AFixiDWmxHE61oOMmb80OcRIQNAjcLarHkD+jcBX
qm3g7h2y33cASkCMGQMbHCwFGjhCrrKx0R8Ws2DRoWQWZxONvREohZKf09Y97Rip9oWbK7o2I80Y
3F5GxrPE0ALyjPWYP/D/IVktTk2ZmeWjHkymDdg2I5gH4LBjstSq1jcBh4FKflPZlv8YSblZbeet
DBDjetqg2Dtn/Ga7v/v4eiTdBD1mrNULiL17qRX7nH5OsmQ2zTXgPkXN6Kp14rdEYi4PZn1gnsS6
LPoXBHuQcm5ooCOm4VL1bYkxwtC9SyXgkywyPyuXvkbPa/hVxNKPNDP7f/aX9ccSZ9gdoRX7VyY3
EzC2XZ37xstlBNhTod9ia3349t44Hp0pNFaPq+o6lziB9v9ruGsLYEc0msUWPhMa0YU06DomQu8k
FBjNQBMD66/9zhoeDhh4lRlqfU3vVTytLJ+2weNXbOtIcm/v/0D0XyUFJnnTSV5+63Ki47pSHuH2
m85BAECHJZxPa4Dn0687LJHzdQ7O2zjiaHFmUj8pga1fEg7ghsR+oxrHDPeMFRWom6rs7ZBafGOQ
BF/GU4Xuc04IYOTrlTPbK75AtdFDwz9BUP6bsdgCy5EkkfAX1iVLSVQiUJi5r03ANAZt5OEK6VRU
2FXMPmGaU73KzB2a4bseCzG0DvTl1DkXMSM+sTEql78TO+Bz7e9L5NXsbxr5MfuO0R+cCiahzzJP
7twynpR8pmVN5Vq5UK0j5/wF/tiZ3gpHVSU+TbhVMuv7pP1xHrOnZiw02nZnc2U5Bj261XzuBfDW
FYO8rktoC1U8MCjMAzbfZBOFAAQHpCEibOfcKrXxXTw9VK44Jz8ZNlBKMki7DyQzJMSjzHDMI20x
nCpqzldW1Dk4W6DZOKlanwBCW4Luxdn1SmeSLBS+dHZzuGy5hoO4gRCQV855SzzsbuEiLXE5Uwd0
+pl2o9ISBQiahibhCb0h9TJQ3ZoqLCsnnNYnNWWaKIsk2PTqEMjmzys6+8cdmJJueAE14emBzzOW
W9w6vrF8UrpBjXhtOVK1GkRJujmMcmh9WQhd4igRWg6Rqg7s5sNROPvuFGtjFcuCyU+BInsQIKji
2M+xYC7Z3VK0ifPdQiNrbQba2w8NGKb+TrOVpt6Y7h+vxs5c22s/w7cPNu89ZkwAq9k7WamFJmVZ
ce/Ay3L/TXkWJ9myO50FsNGoDf26a8I5uyDrRdWCQ4o22Qy+qenAkwJGy/53DW9oI4FZCUuOk5kx
ZeADTpRG66LY0RuozBf27ypET+nmgYl05V8/YWAbTfyMOuVraCYjoysLSBOmBmt7hmybB+oxsSSi
Jy1scyJsYIn3BMAGiHN5XRj6ZtHFGlucNLHbNirPT4llWbDz0ypf73pFI80YfrKYOAP0SbmMC1zi
7akTxC6YpCywVE9mTiZCefUBNRXo3z1jYhiQqPNSjBLlG+Et19ExePgil+1NC2HroQ0Zw/3xHuLq
vdjrcrJ57Ya6JKfckpu76m9pCnHcg6xu5SzeM6u3OGpFI30hmf3t6UX57EttiakBxYjmohxvIQpM
3t8caGLZtLFSVolJ57gtqUbrjTleeqmCx1KM2nYlBbQxmYLZga1T+um7/ZdzNy1dTzpXeq4pBeLe
Osdbwp3+VCiWxnb2wZyLUh9rvXh6x6n3BJ/WVFYkGK7fIx7DpwL+7zH49Cg/HAGPNESDE1DSO+us
ljEbKDlwWXmykCjMf/aJzOBYTiFEkFbrBFfx4OsQFPeQwRufj+WW+jhRAtAbJRziLMU6jQdoc2JV
m+qkecewqgikISudADF1Xp+C4yG4Wh3QTkSUksYv+8WLzdygPv8gUwf12OMg5DXYnT9wCaCNqMgf
9fRWVFiF7f1FHCsP3h64lsQAvt9gf78BnPXwfZQKnkgKs7ij0OX33AAGGOykY0K2l26lQ8hta+H+
96RHFLCsoyt4PbMeZ5YbxEC3cdodHyMJGVZ7lbq/CaasHOP7npSwU38hNpr5NWqjwsPoIdKRnTfk
gvz8R8NvjbMKwt0KiXnUrNes1stuU37Xxk7XlTuL7OzzfnA8VqeRwdCggSXK4IabLKhM+JlFkrYg
jnudO4O28ccOhtQmO0+IH8Q9/2zkLTEfFahrd/cGIs9Lw8U5/Id/gdnQ7XIjw6PwvqwCqNUYhcF1
9lnc0aNKsrIwuhGiITB6yJrgro38+2QM/6BwyFrSuA0y7xJ4c2WjQ6c/4bWQblfkBEvRnki9ZDSI
kheFi69k/KtknAD4orcx5Nsg+kjeQRsE2hqfVxclSabAdz0Golah0hE3Im3L5pWjYX4IYXOeIe4a
9fYXAbBqgDnyKzM5mv6xZeU0bb1y5olQng/QmkOpK5dCVSCCtcTjo5+qY4FcHAIye15mqARpolY2
vOpTF3riS/001EFQwLcRFK8ODrUtKY1NAQ1Nabr1fMkvj3m4dbw5kLKjJrxsFV7EEBq92M+6WGXj
8PZD+cIqqiHmXn79mhnxoz0fv9bbvimTCjuYUtyPeBiVmjDSz23pfvUgHp1C9s5JdQ1BI2MLsokW
eDti1zEtBsydsKnoGOYG8J056DxsGOhXkdIEBF13uC6NjywZWOdfByVcIRqUCbxrQ2lEZI2dMYHg
2WYckfxvtrOyoRs2IbaBRo7xMdG4o1iuwqTAL8imbfFvKBYu+QXCvdXJDQgrssiTxCxpFYabnOU4
DDdrQYg8Uy+dnpcBa4YBV0qsHJqNnQac757+LxRg4PFk95YIMXKfBzULy7kW1x489t8NyazhFwBL
0h5Cg89zcKExePb3zR6coc8y6OoQXYHDDOrD9L++c3gUea/EcmRYD3UuVVuODTBLcCvzl1f9yc5t
xDay2i3z3vaBUlV7QYjgazwiQYLrwbLVzSifhfnyN+e1lRSMxnZRuXYeFVQfNcHSpMyTqceESeCc
LW3zilFFE0ra/uaQ+yJ42dLS5c3lF+gK7VRFyTg1VV+btF1+A0hH88pnUIBio9onUU4pDqXVR59a
88rez+HuEPs7eF/U4RrQ9r1Fz76yH8p84/MXn24aq0FqyQjhYDYFSNoME6i4ggWtfjZw+4xtPWT7
wNgvRM0WLL1t/J1u5vnxRLkUP23PpaZ36rq3U1gMugDvmrUMs2u+z1pALxm3jeR4ZfouCoR2A/dl
QoLJUC6l5RN83BfW4iO2y9KFW8GgNrb6bhEVaCJtNXCU2HHYAqFEAnFg2ZvKCniGCN0P2BCCxZFx
gpwS2xawePLG6QbKJAtc//YBzRB2sOlt47O3S3RBNOT8PZkHkjJ/yP7E2uPCwqxtT+0rDz/wKFY2
+C3b+6tteWW33mOmPpC6x59wIb4pSOI9+9xiwuWcrz/5nE2RldSoIckZ8Vm8BfhHQcK6KziLWwQ2
8kqUw2ykAgGjeqm9vwtXlbHfB/VdLfbdpR1CEPNPG5HeLHQiwyOwx8aS4+/d3ZTSglrPr9YkaNy0
ByMP3OpR81Ahidnu5xBqg7WndRSxSsKzCjZxI8aRFlx1rjUnuJ/yzSiTzUinkDESr4lew+LMZcUT
dC6Ny0Rb7RtqdTF9RGjsLjyoxWCslPOcT2oxe001+rhOTE8vL8I8chvQvIXJ3plzPKIA3O//bmvd
Tjq8J5gVC03H6xA1aWqGcWOkg3W33nEIz4bBebTF10uFA0J7D2LF8bYkFChWQHb87GXBBxKOlcDR
w88vHJAeY1L9M1Vv058ebCpSdjgIsPbDCMPgZELxGXJUSmHePH4xt5DkYFCC+wvP+V/XMctVMvZ0
jSF1Zz+IFuQvAH4feTKoELWYYMwCGtG5/DWNdjPpB9XklPpqr9W04dDOWz00FBjW8pdKQyo0U35R
7JgMrfS7azqjTXD4pIokcKUe1zvf0OME/ZKWH09G0uBFvuwpWSKzIdwRJthEhqXiEoPNr5W34KpN
H32NJYeYIMQNs4DVkWndQ0kIj51kTUsSrN98uRh68SmulWc3bx7sraBOpHOJ0cyANDvyblPjleB3
9f6rnIwDKe4aZnX9a72MNTOzoZPxuZy+mvarpEWxvOl3FR1xjmKXRUO11MYdQCYdyAwgl7psVTdl
zveYLZg/EnmcjshUJ+DmGrj7OxDo3Mxj/ckUWqQbnbAL8nql8qhinTO6lWOcjrcHe0EEhYne0Qog
4INK8evLDRJd3n4lqmInftcun6dhoiN8tOWc1eKYroLC/FAE+2k1I8j0myEOw++3TtRANHd0bp8P
axTYTbxoR3729MoqATSyrSSuqvUTLjUvNzisppawPoOKySTSfcfGTd+rMAc4tjRG3IQVOsBuaDIq
cqw0xC8elePkFPv/pBBdqwR0kotTDeT3TJY0I/5t5kiRHK+UEFNJuC6F+QJr+5+Ngj/xyCk2d7BW
sh00SeNJezx4WWPIT5I3xJH6sWnQJQoNAnrCaqG9IXpdplhZ4A3iDjJ7am9X8NwU1Kj5x/AgaW9c
4M38ejnSFXI/RtnNU9Gwwsrce4LwoGvs05yxgO8R7AWTzURwwFueHIhB5t31juM7oO8GX9rqQIus
s9N4/s72e0aX048T6Cv1dtXZRzV8K5tf2mSVNn54WE7z2r7IvBlEx9cNBnc3fOZgm0l+s21/UIor
RPe8u7xwEXxHgm3KLIaoiqZMjns3QEMrmNCVs40sOkRu1vCG+JAEcvb9QPG6jOqW6oiz1l1Psug8
hl3JfP+OVYH7/8kIPPNuFkdppEAattyVEWk+dycSEZIyOlL4tuT1h8vOSyzamUbWkfKj42gdH1Ax
Wu2Q1Plg2UG9a0muItyXhr1OJWM04Z21SOhVFSHJKNNB5TLlpdQxanYgalvwDo+V4rXevpWqcUw9
wl3xlq8Pf1+V24tHM3BOq0CpRTplBbLZxsXeDdxn1mvCp/DHP+ZIX78+Gx/ABLe/2hDPlyxTY+LC
FmSvmP5jxaBrZVYNBZuvXpVr5OwIzBITt6Rq+PMO5f6vGHVBzr8t60jYSW/ZorOHFbWHpV5u5g/M
vspBPqp0VBP+4eYsi2+/Ftc8ZtxxQxtLcYqj3JK9B8vpNCZ0KGwiXsQsy5I5XMTFQmveWGgtk1H3
B/hKd7YR173jw7mjICe6P9f1BDhP/gmp8kh90QhvIFC2AVnlsajtFjjohUbpK0pkC/lX3g+0Gmk0
4qwytFbYIAvbrZgRZwX5PX1rAcQ96+fGe71QyS+dMmOoIWLLN25l+59Yjui4XAjTwwWn2+PoUk4k
XbdaIoNIkDaDc3kfswweglpf9wJtFS/4G8n79Mx5ozU6UM6MeEQfeuP03hw0seFZ74viBLto9xBN
YfXBEgdjUtNHV84smgqtkgc2L35g8wLfUo102Qpiu6zgYgDcb15YvjqE2liBZhi3EXydt68p9EAy
sG4EceaoaQH2MbibuaoISrY217vKNZY53ryxyU37E+dO3sopUgOS45d9QAjbi7iz/kagLOUjOIJu
iOwXe+ALVIk8f8mXApMalJI2akoK0wHS5sru2nsuWh1Ss/mbfgK2RUmZYe/wJEbHrWjRDr5ehf6S
bxpwfWZVIc/PAyDiAq9tawFEUpNaCXfdOvEZJzwszZHYcW1ToOZxPQyhXMYtd2b1J1vt4qZNdxP8
GS1I3Vi1nHVrFQQrBYxhVPTUL7uYrQGXPVgzdRgY/nvcRVD2NhvPicnJogn4hFlnh85Wzilli8b1
8bXTlni9qvJoXubfXSw10A3mGxtYE4TsXrRXJvpqtNZr7mPtZd+mKoECdKCcIFaQEWKq+57zqD3c
F9rWwfIpLkmqch3twfGHvdUUMOGSW/6NwSEsgp2a+eLG7jDaY7FEClMOpv7cESIi4MaQylFD8VFG
q/iy1wqugi8uv7mpnYon+ofYjyr+AN06M1xyXKaDzekQXNBM1aBLt8jh/z6JFAjAySHyiO3kHRyu
0fkxh1+3UHZDtFXpC6AXNvcko6TlT1X+3dlVtA8yV+qJkApH/8GMGZUII6bWKZE31VT8ly+oik/G
MisRKeNdkp8eMXKGWmp41xp7n4oJpmXZv6/h52L2He+59VIt/8rAblZuVWUSidQ6eN7hJZWWtRYn
9cFq0A3k3bCn9LIP/LWtCBCtDrHdr0Wb8xeMhdZL8Sv06DJqSqTpT7l1WGsQzv0hmXvYu4noa9TS
D4PYbFkf8rh0Qv+nbTeu6o2TERkf7rUOcyy48uQryRTpwadzpaE3mzaO6PRb2BjBTZIhRedexFxW
XIq4EU9vWYvGBBP00nfr8ZfwqaxpZCtvTLJFCzcmaPEO6UJseuSSCRHXifHu3nufCeOcmcpxL8Yi
bFqr+sTChIm7v8rV/LLEE8C8ni8aIEBmmgBJXGp5nzk4kuvCpLux5ojhNEgnFxkPPGCBFIXV7bAf
pua93eE8Bgz5sJK54TZG0CVmsHjpkiXAzEduC2d06NskGBWhxFIMyE7sEGlQvsFGMRXVtnhapRDg
KkpDNCaQpVdrVVac4XXw+BqwbrYY+1jNroBQ9UbM+o75w+cDCXF7Xh0bkUJFS6dVCb1mEHVEDSEY
6JwUOXIcZzVq6dU3c5byJLaC638HOLCUpGPKfizRTReJiGCHBgoUBZ3p4qIke8T3VDSa5UdsgWSL
9CaEjAusaC2HKEV4bbTDRoUpSXziWySP/Xc6yYpxZjB37vEkFLPK3jJ7TJiio86PfsM9x6lNP+cF
cNCH9/AMwiHt41dWMhNdGBDPn0aOEVyzv2oIQjsXta908NLhjHZ4uAM4cutFZsM9HK5ijHlpmM0m
u9amgWDvTqEPA8SCurEFDrrZN3xE5oGcGzg5o+wTdDLSqZs+D1sOotRdcVvO7BN6TL8RlkfY/IdF
dnDqzOlUG3nXJMm1kFJDbF8BF9QEpZqVT8YyBCplxBMWnJOSnhd2I5N7UN5mcNkivxTvt/KnOgyG
UtvAEdJ5w1C/CCxyvwghor3ibAX22MjfSnw47i405RvFDRfh/eikr057cxvnEyIn3OJe3we34ZJw
B34iDzVaoLLZa7BcQyvl5+Ch70+8RKB8qx/cXTn24Y6U33qmPign0afZVgSOtcDhn0Cz1cZuiF2z
Agbal6NtxEGTBMVl1twhUcBSosgA4UujVZxIwg5h1+3Yo532mtq4f5si6jEqvEEdGfHQO3yu5GyR
fZjTCAWdFPCU3m2J/BWOh/RUtLsQr+7uzmq3v9vK8s72WnHl8rQ/tQweNHcqHZh0gUx88V9JIfZ8
b7qG0nWOoSUa1pJJTZBSmcL93nV6V/VOvBVF3H2zyW2exJhV0dLcC5P3ueh3siJrKfw+WSvDwG0n
w46+jKM0vwOAt8wAbk9sWYn1/ZzwAc36G6/KoomEV5a8pe6J2dpDxeI3SY8VQ61aRR7GIyVAbdwq
KmYm3xgnLDHtnH4Uzn01nFzBy9oNuAGLOnWszZ3hvOmIS1hDR21YSDTdryRUe9giibS2ebdpNRVh
WQsu+4iUTmfSZR5G6+5ppaZ3F2JL1OAwER/WW1mzmFj1nXCy1eUtJs+DNP95UcAc+QOxSKnoUTXk
VX6brGDYSxgS4SBpP7tA8wuz2F4/n5Qj0Z6UBKD4fpNvtzqDrH5LCtA6VD5hlAlVp4jerw4UZzAL
9UJ4tKRt3vpWvD5P97FhT8f9ctPt6gCMg5nUd5YbUrxx5dS1QB6jaldt7q3qqL01xNBdwwkwQnoA
BxUmR/LHOZflTuZ7Dxz6nZ9KPP+Fib00G4pxUzx4kBFrZjS/5pgCJfa4vuhYUn1X/NQuFYI8oNWC
6b8RoMf1zTrrpurmVFNEeBBsDrgYkix1eYKCPBnGEoyRz1/wlolP7uvqkGtHayO+TUzqu6yt0fNi
5vPt0DvSqQ9Y7uKtYhwg83p1Qcxmm1xQHW9YsQLRcizQOFNHp+rsbBj+G6Xd40q8KH8KLHYJ8lxN
nL0/E3ebVSmwXHjlflwAsrXdgwKYoCTt6ct5iLl2sumGz5dpkNIVXxwZmYfWhvUKU58fGdqzk4bZ
UMCGvQHoEnX49BU95q+GLLC7pRMJfZ5HZI5f5M2y/yHh1Ep8ia4pVcwxe47jJcqkP3fJ7+SMjuzu
ZcHKin6TX8dQU6XYFxciz/gVHqQgXomkzhFBt+7VDb4dbAAlhqdhdSUs8syRVT8E8I8Tv+QmQC7c
3Pb1YeruwUma7cCEsaE59VMSJBBKNZB/j52K6y8i1bhPcLLJTGbjxcYTF0FPHnAmk9Vk/Jp29gJD
mJF1lB77zALmORbjDbWPTRgvkWFXfPRZY86Kq4zete7o8VEf/88qkwAaIQ3FL7/avGpNzyI9r4o6
rsXI+ljl9//jjk788xPnw4tv+EuJE/22xcDhQJpuuJJyVitoITgJb9SPzKHk5/PVN2Gw4ImngAMs
mNKR2pNDqMatXKTGZi+8F90Ik00jGUUwEpB7uaqhtqjkHjLeVwCg2ynGKousGZ5eiPu+0e8JoWQY
NiJKsNsDy9gmsO8D8znfUh/qD2+apJK6w+Gd9Y79yjXrB7fCS8mnLL7tZyfnCto7smZSF3nmWxEH
KlHP1DortT5flttb4+2Fo1ztKNTAKG8gYW4z5S3WXi9Me8ETw5zRjgFR19SLisxAdn3S44BMYCwv
l37iTDiLhxfM+ZAfJTMny/nZvZ3vukWlYTxwMckh1fTFgK5wp19tvRWstboFDHPrfBcNYh1Xj7jq
QqFRGbHvwnbLZHXMWZu7weHrfT0jyM/aAOJ8s1Kum0Lcox4gdaKa/ZBz/CBayU6Nu84PX7OxTOXR
XwzkX8IYuV9+p0MKDk+t6Vpa88XN+HdKiwDZMZTpBcKopTrbGatBbqxGoZRVy8E8nuWB9bBpwKpR
MHJ20ASVPOOR8lj9gC2Uvc/Ez0Ky4VyD1cOa1yZ7c9BclSe/Bu9MGLC/RTqxEHIIDoBF23WgCgK+
PHj0Av8AdMbMQ3eM2Wcca3TOlnyhh7kw25LMhu4AmPtjB/oBPY2qFF12FZNKPBOUeqzA72psZWmT
qymMXBaNqgBw/nVpcKYMDYsS43AQ24XYxvILBGIB9G9vNAFbUxugjccrw8XdJhIbNGgh+Ra4LtoJ
NGEn4sysmEZd+5UjFgeokyC9MRvGWHiEIb9xrx+N0+moXSBVoTxs8fJftROq/QqNBKROlzPx62yH
h82PISq3SydOElBgUuSetLUYz7gRLIAG/H1QBIHbLgqAFW+mqwsf8Nrj2/SHSn4SHMTiyDfUwvDR
DTp7Go8nSylpunf41g+AqyJa3LAP/C9aTaPa5OpTPITZTka3Uizp6OIuElWspCF0fbtuAP/wOF5B
SyyFdpZYLONSt1uy1pm3cV3AFW1TbfpHdENSpBplSA6ltruN8hHwDN+XHnTc3mtaHQtmAqyfA3wi
L4kP5SFlP/Kz0MHSdHeUvkkjGaWl6FcPqKJ1q+exH6T2aSh9JiB2GpiTdbZZhhRmvOccbMmEPkq6
P/001l6X8xEM+u0xugBM0RCYZ8vxoffDYBQRdFW2akbnpUmCYxZZ3Wzi+2TPojbQS+si1u2s3qfX
dnC7GugKM3ZvZ3MxgVQwNR9oNGSDUxbKpx4jA9y06WI8HwMqCjuUOUpz3F+ZpTVgTxnTyPUK0FD8
7Jr2NVkpCleTuKYkRajdAjhJtU8n/QYDOTWlLEClG6byB3Vg25oMBXLV/I+omckDguryUKKNhONO
j8aNYjojLwUTVhJ2hARP4UlVwP8qV8UbKAJ7E/9zMKb6VHZgo8vMU8FNyi5ceZQZ9hi9zHb8MrhI
KH2H+dfPEdUOC27Lkt9kYRzsP29qGEiufbTZwGZDExRJGORhNNPk6rMZ1/dqGtcoYkzVJaNzg3f4
ELdPEX/mHJCkhySuCaOoRyjR623cOnaCZt3l7rnClNOBbwpqhgBPtyjCAfdh3Uan9mHVTZnz/8sB
A/Hk5Iw+18MpnLakPmi065Qa4HvMw9E3pcUYyIsS3nhabjU1YUmHsZ6rVQD9UHKa21+B7YEl48tX
3SmDmZbCtnrLKnwRCGNfLRaLzXfIt1WE95flaehZHlla2RG1dM3SadssTVF/eySU6eRBw3xxwXmk
Px9gfHCo3w7m64Lkya3ha4NITrDMMUja57Fm3NhjEXTfUqOIEIOA8LHtm8sz4GOnJvtb1Fy8Wu0l
7EhUK5F1GfTkglf/6867/4vjAZE7WO86fmZ81e8NonzPn2DQTfjOvPz+XM0GeWdD6BnwGBTKiq+w
eJ87JZtgiA8KqYrUY9lhe1XwT1DK0TC/Gsd3Uc0cdt+jnKLWkmZqouXNyCurCN5/lrNfg72Bknk0
hwR4YR4C77BVpNlcCP1g8h581o82yi/RH0Q31Y2DHIOZTgtQB72YhuWENUbrJvgjjm+cpKT0b/Wn
D9zqmVWDe4ZjAINtSAYjEpAsxm8yMg1kPEu7aH+F1T8FlqMdqfJ1hUEEGR/Wu4I8yEaSgAT246sI
00Co+rMhpavfYM9lyiVyKsiQyHTpXcaUJhIzCIYo4Il40MFNCXngsdu0Z+RzQ4yEVefU6aohb51c
nxJBq+NyIX24jkDC1XLYLov9kLINlsdQ+duO/WBHImuPieGznig31ZZmfdfcrl8HIwcVafUi+4lb
Y7XRDVjM2gxVlnraW4ocGsC9+xYjmWCc46885qsNucRC0m/RKIuzWKOofaAmJtbx4GXoeqPvzaV6
xwusmxQV9Ww9m2NO4JvR0fyIwlRVMpotjmGlJHJRlQJJGq4KUP+ISSSrZVOTkViFS4qf93cpZu1F
Ykb+Ol+rtm/6WS+UqXUKzrBv4jkBFNUIm7og5n0e3wGWn0zzGniG8S/LmzV26yWdMWANip5spYkM
NU6ZAjK3NGCWwDdSAop1lYX0e57MenqLBQaydP07PIqRh7Tc29BZiWa6OwG27FUFd016KUcnRkOh
5GW3esOx3cSzSC0jLtPnV9cWAlinIBai+c5k50cXkwMK6ETPGjj3vMN2i99j9ZX60im7xYLTzGTe
R9Dp6keMRuRpU8Yr9utftOtM+lQZIgwUsg/h6tL86Qu97TMV6C20TR7ucjCbmmTG/L0cXvxESA+2
nhGdikQMKIeFt5KPb+TzDJqbXFOaD/ScKIlzRKBawskQAydeYxEoKjeMvxOugMTGKgxQFU/HTTJT
fxEXvBcCiuRQyUJ/Zrx+ssXidGgCUvXW1fGIMxTCgjJb5p7aLUoX0LCHQ/M3Te1IPIJWgx8JdI0f
vkbbS+AnwV8YkIBrWf2lqXAImmqVNL/GKW8GaE214218Yr0zmQ9IThQPbAnoyP8slQcHFDVWd+fz
piWUV/XbyJe08hdnhyu7D6wym4BCakNfdmrxNXCgK3RopAc4fMxcax3DfjmSwwj6m4dhTqj68Qw5
Hfcs3eoni3A0FtLGupbcQCQyCdP/TwgQCHSTLAMUeKl5ftI3MY4S3VQHrJwMt6N4MC3vqstvf0Lz
wmnHfZtAOFBRA0iQvJeQ7Gw6ISDFoY6Wt/fs68bWEHlm0r10WI87t1wXpJF2fXDSSzDpqKeX3NTE
aS/pAQlkM/hboiM8pWCQEaJF7D0KlnQzVMkR5Hlm5o2DB73Tr9Zd/q56cbAyvkUwf7rebR8Z3u3O
megxxyu+vHXKYsWGoMbgYxIw94q3WRUvZdPvL8Ujpsrh4qu/SqeqfNTxBd9IbqwosfdUTXk92+nU
5CfoCAyXuLFK0IvufE2ynlLI9dFaVj4tjZbH7WgMY31Hho1pXbZqd9kBs5QH1T+899cCVMDqkMEB
QAEW6FGR/VY+wQedUV0zNIWDmdXPhk//J7JjtutCYoWQmdtDelSMQOI/nkT8LH+s6VvnRn/pAxps
50n4WktSZ3gYc1FGKGgOu+q8+wYr5IApGUY6Txy45dbrCPvAVGy6pZwcKNaqCah8Y8F1I9ZKqvrM
5WEFoOVURTIiYYo9HjYjeDzsmHbYVNhhDdoxoAb5HOxAl1C6UXVZUiIa6v/eEeEXmwbUqZQGgDoy
fbR1DGixktcRxXrbLwkXzRA86VY+5WuktbZynE9b0u4ER6H/S2r3MfOUrNbJUJw5N8IxBdVCV3hd
PE4ccCaojhnvRfebtf+v2HGdnDS+uWHMsdqFgy2FgNcf+nbSslhck8nTkdBgAM8OcdJWt/N5s4m4
+f1RPy49u9+2YPK0X27yeBQXvbhYfAvrnSU1cZHuwcT1TnWkboIKe+5f35eoWghYRBrwfk9ExueJ
iSxtChB1Q0DjurqsutHaLQ1PUa5vfifdfT9b8c1yGpaGZRJsD/X7u7xGxIX650hkng8JmZqEjSqn
WUxfqyQ3pS378Dkd2Qlv7QzIqoAIlTLnTpvqmR0dVj2887P4d60+eQQHLPT6ck63xsxCWOisRfRz
a7xunUiXVVXrxnWAJsL0fQa9fI9jItePM7XpB39aOCf+Xy9OGc7lVeEoITSv69gMSLxovL3vY/ru
Vdq4sdWXX/Q85xlDqTnkpTKa4WCzcU6fRYawdI5XuMBu69O5L+49qYhwINTbeJgtF9HpJ0CcbIEZ
qtfd6u7pxAnCY5pE8pjGyOHHX2j0k1sTrFr1HD97MXn9LV+3bBthniE/mILvSiOE9XLQoRLmEyBD
sYpLJzpjKjZtWVCIQ5CDwBksvlZW7z42z+PCm5kpruUN2cQ+LHkWnHp37xl72IL+NwmrmXjMSJz1
8JClFFOgOQ/4ADPN5UcspErlxjboBnWgPOj5Y9eaZhzcRP+bHquMbNfxbLjM74kBbNiHHDncJODm
bqrY9iHg8FCMXtaCIxv21QAM0KOeRVznFnAYGBB3UgTY2YNaEpN5Sn8Xt2ciM6f/sLbevFwxWzGe
zrQJ27tAXYjylpixVnM2/UeMyFUUpefYk7qXfxoeynXx/G6oJ1iH6VxUa5jOwesb2s3+R8VUAT14
qVwco84OWS+joZUiK5dDF7b2MWAcNU7a18RNTGLyFk47V9kcwDhH66CkHIlyIJqb3JCRJpECGSSN
hjvp+5GiWeueZDqhn8TuYSO+Hm/C4Bw95rXuFUGebNxXxJRTUO0tPRm1JePaG3VtHU1HqGkFDovz
guwmpc2JI/dKFalUsM9uv0UpJ5Zz5Gp9Fpj2FaeBBBa52VOJV4W7sibGKBsFgGShoSEEywN9uML7
cIvMcHUhdtSjOfdNR37Sny4JEJaiNL18Kp7FFDobEfyPVpkqoqHslPmnGia+4rYoG6u0PzRSSrK4
ONEorKVINYsRxo+yO/fkT3s6ivEYm9wOkecB3C4GJJyKlrhSMGVeA4L35ChqI0twwTVopgwQGihn
+EQcKsH9q81NXrVrnFmPpeIm6MyXDuVng1IkC5oJmWotNEGG5wuIhtHf7QchSGc/JBNS1xXi94OV
A81PmMApoKHn7ZscP00jtjwPQkPEdzAc1Tubms79TGjnibiB7NqFhjjUFqiXDO0vmqyzoD55MVPn
N2cbbhfMORYJlxXkaUmM+IPZCIIWMxCXOP6/qhVGlKGDDXUiJkemmrtGp5HIvjCBWHWPfzAF8rKu
e0gGONpsBcbcpMvjuasJ6CKCqzh3ZVVIiJURcFZ4Ds4RvxmW2lWbyPEA6sSs5VzQwlB7WejBPzjl
22abyakLuwLjMG9CkV5C05VRtQ0cyvz+nF/mPUSrufPSWCw3/n7/u/wDM2jYTjrj6gCs4j0R4cfL
5sh4M8xJphg4ibQKKNk+3Ww5oE0QIYgqzPfOH8xCjacCkeSOORnxroCbuJrUkH67K29n4kOaLy2I
flPLi/5oS1iNLOlOWOe7v6ssDvZ8HpdGL/PQ2+FKuUWe3zi9k4SUi5q84eEW+enqK+hQtwTPynNs
4df0HKuwL9WmTr7/xcXrQm5E3Y8SXtvv1toQfR9ViDMhAgdXLLMijAUCoGP2X2iaV0d21kkLEft4
arBuO5qeh6ooENg/CwBYVhHlQ9loOQN3bzSAqPGY2862igxmeqcHijc+rmNSiC70d+4zSbpTD/fM
mxrxA8ptiQ2Bb3HwTc8xcaEQ7eacRThtBrC+sfO1nqEZQRg+aIgZAVMjiGNAlHXNqPp1n/zIJeP4
Znso2QtGuMpVSf+Y6ZIHT2Rj2Qaqhkf1ulwNrCZ3k8WNZGdfH3WP1yZ8HAqPHL/LVDYH68leJdVd
souG5CEvoFpr9tpB5Uae6tBqYKhP6X1oqO3TFwAPC2rPINyuMaaWHzopOjICWfh4oYJn6m45gKHP
E89RBeAvPtkX8lASKIWPsmJKcbDhWuHS4gMSEUnNYPeuTpAYeMjGLeXs+9E/ssA3fm7VrN1U4N33
1GF4yYw69VY9HqhQv9zSKGehipPt3fceg1pPQksQ1+2LFsqw5SqsfQw1c3CQ2k2GEmYKK5n/m52T
CRjurKKTan7wy2pNnoweIQ0gtj6MZ+SMM5KOfINA+ULk4oGjriHMp29F9TYnfkxB5bEi4UgcLVPc
rHrvJVPw4dskTsA105TEZKRxbteD6prWScSooNah3AQbIohWcEmhUJbodAAmJIJNTsoBNUPALTFa
pG45l8qzgjEKdYXzeuG1O58Onnjt3cMY8xxSVnEhGcRrb4ePTQpy0U+X03A6awk9OevY0vQjv084
08FrZK4zyb6wqYDxMOz1P6M1TmEHsoVXQsbNWlS0UHuvKGKFTcp26ohuaK3KrAI4JmI6QNW5VulR
bGtd6NA5ZFk1ka6QosvxHkS7fRQHA1HCOF26bUzdkUCS+1qocDsjVMQU9mmdYkGVdyF1CgGXiv1C
0JZFI06xSVbfyRhOuPxeZv/anx9RiEveoI5jlS6LDv864+Yzvdto5cfvfJEyMzWnmEwPLqw+8hOn
83uag7EYHmA9JNuKbXNY1ek1mBVzg5x4x0eO1wWKUgsoozGrkK+pMY6H8XSGl0pTgyLPqKMPGNWt
DYVCcmrWwGphRkocOJ/4gOUU9kXalAzi9BSGFzfAYttJ83wDWVLKq6i9mGMNJDysVRw7Xh+GFHg6
YryQKnZrepzZINwWqOvn6BgDuBfd8xX4xdu/XptVT5avz6nM88zKAXnZJQTz0Jr9fMUxcEiglpSE
tzP5x74E/UDuMB29e/4u1aG0PHgu56NZin1QacxU+sEuFg6OiclGnCWNMYDT8JfXi2dshqzubb1r
NeHROridzCTLg5wXB19CbWLnqf3IfTmQuhktaxk30BELqqM54T8Suxqi4rFs6luYRGOFzq2XIvrw
2U8feRm9dRRjKPQ0oa6Dyh/UC1QT9HnNrMqH272wwJz4G5xkrPJlh5nU1deiXQMUGzlpewZf0O9x
Ai7USnfmjA9LUKRqQuw8RlE+LH5KvxAL3mS3w1/qprK8sdw3AYuRQAEZeUdSKH7oYp6OUdcAdc9O
t4X9Aa088bBWicjBSKj+9W2vi6xkG2R/rq/iU133EtGH+bIGwFs+O+DG8S3p8FPeF4HnrVhLBEN4
fMfw9NAQjZ1pC/IhUPGsV+lfTTRrQtRNv9ltTdXMC8SWdLZuExW3fHYVctidDHrUHtcRnqUgLqt0
UYk0X56rRgL/gk7x7NepFc4Yzbwk/dcM8o8R/ClYzTe7qi15B/jSFWMJ5Ris3+0i1+99BYwkjUsH
gx2bKR/4EHIybGpENxc/gd2rQ6RHM8Kj+2kqMH9tXakcIXhc67HaJ6mYNtPh8+wLpL9lQOj5kSF3
beLK9+ha7cfe8+FwHaVsZz/K4abjBX8eFzAWsQZRHsPwoVMD6tRjaLNcgarUHch6/EO3k7x11/Qv
QVgbBB6bZlZXrtIv8TZ63D0tq2qhX0DB0bI0mPDnFAU4nWEQNEKoEk3Q3FU3dgrmNqv7RYhDhaIx
myXwzIpIK342vtdc6cVio2GUXAamCgBQq8ZjuliwGhXUJArtctro2NCtbXQnev/bdei51mjTsScm
UeWhq3pF/IFUe5HmyWlO/h2J1YKsDgTlSsD9EBQKbEQ4ShDZ0OJniESG8mcdLdV2cYVlpPHXqbpp
Kl/qrlr37kIPdP2BuMFzEyg0zae8zDvhqkyUvzblBTBGX1YycvdSawve59CyRcqGZa4JpJkt67hM
e28nYJyI5aHK7yErqtKEGo+Hj+x/Axd5fFCqD8Z5GUh1MH5fTHEizbb0BV7XlKlOIURN7d2XJEmR
4IURWXnP8gUijIvR80r7eL1K9a5B1O0KenpDUXwAKrpdA4nAg9cWnnRLG1a6h5gW4G4+DeARxeJu
reJyatK2XukOaLzZcCTEFfUabK8R4p/DDX0fVm8a6rqc/mIdSdhUAyrK4FtmbwTKb9v1NusYpUZ9
cAH7rDusW9Y5WSSR8G5EvU4yuBkRRnaNQAJyzJxlqZZOf5X+D1RQvl++LvxDGJRlAmcT+h4SLTrS
HybcBQjorZttxBOoNADwETUe5cNrWvT4wd/5fXWyRkopw6vwKZLVMIYTpRggUfK00PzRbyrQhOKg
1PKmyAcqSv8wq95Bn4sj8NAVPx4AxzCdtu7Lu96Xpi0mbmbkw/1OWSB5RuikB9fVS+f772dYA91y
9nVmjj9a2HFLrr4hnNAyN7/sDw46e8wGubBWn8zfSJAc6w4jIpOX1ruAUG/pJeC+UHQ/UMrDawpm
1lnaeX0Iv3+JeAKS7w66lwWI59qFhkj2IiuXw82LI+UL0fADz7tWzolSv5nLG6WycKCvLmD++P0+
+v1z4qsoBGHCPI29iDDLo75t5HMgtv5jnCjwvBooSaIOWFfMsIK+yyu7rkbX3Q9+aGs58c26dpIW
ewjJOanAUlY+u4AllikeFg/M8cLAMFGjwuuUPyX36Qv2UWG6LI3fESDzmF+wYbLjGZ9EI9KH+efm
D7hFk/QR868GIZsUtBsLNKNAjfekoRg/UWyDP2HHabridST8ObZ/SUcCkL0AQu7+iz60Jv+A4TqY
mMI2oP15xLNXyAUBVS95tk0a16YN4SeTxbE5F4GrPQFz7r8YeuZe+RgsS8lOB/UX8rgh/ZPUPCFe
l08i2WssgZ9QWIJSIoPQuxJZpZ+I8m+a4c2OEzt/Y6doeVHSdHaR99sF0RJEfnlO9n+mc4VA78Zb
xd40Ay8MlQOgPSNFjeM9Nd8H/J3yKgi+P21wX5qiuKnZhSpJ02TwRpnNRS3sJMlGuQli+qTLYly8
WUuWlhWG9TK/o//Z7hJXGy5qndFWI5m63bI15LeV/OlkUULD+VxlXD9Mb71qqjskm6bVEaGueWwl
fp1rmHeyRxxh6x/Ld5mFLzlr1ZmX8JDgBDXqo6XC0NgID0Hkgpsls1v/viPLzLthaQwcuLO/P1vw
I1U6sJE5YUHcVElLY+PXfCUdJuHN0K/Mj4Ibok9Bs+rxROLrUV+ZGyF9N6bd+Muj8fUaHwvT8lZS
va4sOunl4Gn1fQsPIHpVhVloz3wmGPFjtZjFwvw=
`protect end_protected
