-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XrZKu3tnpDCnYk3YDE55jNSGjJGCxqufinh2lZTbk+OHegfvvBLP66YsTayA5SuQ4HOZHWOOQFLu
qY9rT26xt5D1SWLfwcfVCWqQqLnRdlttyPh7+1yRSfWmC61YTlrGOzw1WsV/aeb0t0ji9NmaVkCV
6nK8OFzPXSUR5BuxnXzMM6v2puqFjYZR0NulVRuKj49ciCJbfIlRuJIMNZI+EqjolyOBVPgP0kOn
B09kbEbUXaj6BN3JSHJYqin7JPEfXayyvdJ8MudTXXA2O19kEGkgCSAmKWKSgBtH/YNqqYmnGynW
2UyAYZAEoM4jomYNoWqQvuSlJn5h+umZg56t1g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
SPl/qLHeAvoqH7TWuMSSJbZVDyNAp3oMXkDvCyTt0GnlAgWwECyb81cZ8Gk/xj59T300zp8NvaPl
el1g1o56e2/rCZa6JmYYgAu2gm88ka6Kym+mk2ORttCqOhRUHaEx0MwzCa7/ImWVrhw0i+L/fgKK
/qzm9aLOboBoVWqLKBhCZrblyNmlPvwbPAAAAaCb53QjZiLC7JmxWsv5IOWNT94WycwgAsFe0Q/u
yCuu2WefRGqAoSjp0nP3RE3UMq271ezzK+LbdxuQ9Uyt+059BGWszjXORqNYyToV1dLjb9CGSiVM
+E9Lf/sI/qo0GDPCieDDcz+Vkj/KHrWQja0r69i81IVVTp0wiJwzFISUgKmKVcA7tzhlrkZXRoQ5
+RbnlDmOsWT37uH4UZOvGBeT9fAGc56LU9DBeNhLb9GQ2H7+Xa1gkizbQRlnAAtmLA7t9ZkMQazQ
Ly+fFw/+IlHjclG7qZisI2Kbkl8/NH8pKj8x1LyOplm40Y6+bKwiNmOW5f6w4ZMWOl1wiISotxLQ
vz2fip1RqpAM5+PdAiDsEppyeeUIGtMeTJkmmnXdc/MUSrI5RFm8fCw9pnX1laSzkvA5XJSpHd1w
RG4AGrT5uTRKuCFHMVcY8dn3VMQWuQHu4yHY8HMeLWD5LWQNSA+lV9SwcTX6qmpK1g4X/6p6hruT
lAoDJtf4znQC5T3ibwDwX68iX9fdhqD3aLblbctoQ4STjQaJJQLJuryPQs/WvQAhEBjMVy+f2uMG
c9z6urzwyCy5p4dZ4g9R2lcQogktZZdkAHgz435Nb24E8bNDOUikIjrG5ThocSIKp3G4HsCRl/Hh
gLk6DQTvN06CuOzAZtuU+UiHVYQjE+o7XS17IxbaP7CR7FvHmWkZ31bmlfk4YWtvwyROsJ6mNga/
zgBd5A0l7WOu86IU9BhuEoQzMMjcEe8f0l0Qgcmu5BPF03nYgIYN7+iG4M+aFT5kjYajI3oTS6Lf
0UCIqYQbdnfZubnC/55Y04Q/3KOmnK03uKnLXhRydBGhxHZ4vuV80scrWtju6SztI8Dfq4JmU6GS
IzagMKVjkRKs0Fjpfe28nWb1Tt6N5qvqiuJJ2O5OcwfvxLe5bS6wgG6zISAyJl3fy3qZaao24puo
yabTtPyTxpydeWmeYjGpUyI48qt6PFk8zI+/oi+RXKTaIAgU1gMlohw78KAgthlkAFTQwF0T4H0G
rJRRK6CTMI+XBzHKzhdShFoZolB7rAGEVaK8FDrZDslssRKOI02v6EK9yiI1FPKlEyTdk1oKRFd9
x4kFTVG41E2W1x/Q7A2NHSU7W1eb96bMhpyOnQDfk4zcIB+TIwvp/1/egiyymcPXmd2CBAv7muvM
5JDfq1mBtg0iSa4RTmYIVWjkR+qd6gTECOjpXBl+yEqW3o1LTsO2DQ3B64hCg9eaqz6YpivJ6bci
kJZfiVUpnLeG0lyoyUJ1tWnHADbZl0jcpWAqDnr+ATv6VtzLuRAHljdEG2WoxftPkLORnpqkTx35
mhN+cO/45kkfIplyDcWwHO/R2Xk5B8MuR7LAuNCmjTqkgA4NZM/HoJ89AbwGxoMAFbvmxQTycqRX
6AV4bk5NRpRDVGXMB5vcLVUYbStOkYWiz30AXo72Yebwv1RWYVoLDR2jVJy1nIbggVQZ+QF812wY
EslWVpKAh3au4U57rC5RcfoA6FK4sp7k+nxCE9JSBa4qoXSqm/XhqiTkccUp2r/jsioDiUAUWxV9
eE5rCaaMNxbTpjLF2UVJEE1DTfQYvDodp6yDcwcxWlVq3yI04olWy4JnA9S7/ySJH6w5VbIozMLp
rFYSLXFXSEPsXkX7elVCkxeCcL+I6r2ypoMCluMyPefJ3wEj9/D+ZbtswmoWS9Snu59HmU1/2aEn
RLFg5xZHp7omjaqpW4FqIw4OYOogU1FRwlEdhWCBQYMIMJZcfS2O0xxIBnJCqAKZ25xi9LLMFqJp
5ldeNesHJNjLWR/LS+t7c5v0ZxLB1Hrt8iltZqhsb7R6c99iwF1VG+fHkoN2eUW0RxWsyJRbaHY4
1KaVSF7HrDQy6iTKr7HV652fvYWTb1ox1Vgi+XA0SMSaFZYnXb/CKC8iNaG2ElDHpC2GXxsO0Fz8
3vpSXTNiEd5B/T7IuFqwWEie1AaxttPYvID2GcnCDiX6vpbh2rhtrjjKQbk03Tv6XQRwwlOPrrhw
JAg7YDJ5GCqfwwDlVsicH+IKgFPW6t6BRX1MgeFws4V8RyzcY93ty4/9xSUwKRAZgAhn2YlxJbF+
KIw25djv9wBIxGb/23EeOTkmfQLlYZBss9smNV/lVUnmiUGgEAfC8B7fGTsAOPM6p7J7aRxFQiFK
bqbgMTWRsxljMv22UwpHQ9ihnD43VuJFdpF9FE4a+vZoWRttinm0rlZMArcBCrvJVdL2+PI42ocb
aeGHg6sNXlutd2qg/8cq8o9dMfYYXsgy+U/KFdjXrU4ILsxVGnKeFeNZM1i+XlhmQ7W7pxhjyEKD
On8jDCZJo2RzzUs2XcSPLYNOk7H91GsfBT0m4sPvQ+b3qayyyOoUzpYMuaanUJPPeOx6j2+uzuBO
xwk2xIK1qlIwGRL1APVt2jIHKPFgPXhdhc9sXwnkmuJpGaP6JnP4cPuU3GH8RgTgNwwTupm10VgX
DJylJgvkEoXhiDsdlwqa9zH061C0TEwonYa1Bw8x9Z2kvYtorGBZqK/cofx3EpM9sVTxDTEnu9bb
8KAxrTfqY6Fn9fNa9TcgVPp19/f5h5yHP/68stcBuMR79jJEEmPx1upgCkQ4sf3gTq6O9LtpUL69
VkLKEkymXtMqHL2cRI/xAUOyAMDFqpaap/ltvHCu+rxaWvv6VWavbuF3qLZHiUPsvM68ZQ9jci8M
YoteNsLwxWD8clKvCB0vunxCRAJhAaRU+Qz/FQFt5iX8Gsy/JytatQuf9/9Jp7L8qcT72k75Aohk
N+MM9nisvrMAw9lSm9/gnlS7iPp5cguKcNH9MgbeaCyyMpfZyexMZqM12n1O/kIdvYQ/eu2aReHD
jMwKgmjZpJCUo5R522xpaCyq9GuePERhH76mtIf3IaNdPlbaVvlVCpALblXQWYg7Tpa6cTl6EvJR
ui5Me3vcedFz+vAJu8x48vaJqxazRevtLnBbE5Op1XruqLuBIFCPpYzcsy8kHAzKQyaOHMRhrIpM
6nOwGbizx9ai33HW8B6VcWxt05EbPMW9+8V0/Kc2Gcv2IPBO2rOpkodvjrL3TQ3fNWeeIc85CVSk
PsJwbvCJKNK1RPB5A9FrkfzX+VcVkFQ+Fr6AXuDLyDEypge8NE7zwGPUv0b9qL0ZjKQbRM4eSafS
iiqaihuBmVkP6u4eCvvtG3vxij56EvuzWyWsmIIcI4ZWBmuXj6/M/GDUR03k0cCU9rHV+7kKj9cx
Hb9kexkQyH0V43YIRjFfssilu8OQnBCUy9rlSgUnc2q41A7/MCYsq+11uBkenQHXEfecOLtb9/p7
GAlFo05bAe8TeW4oXvjoS2TwbXXfQ+ZYBccXvFKB/fzYScquP4zdqRF+XvRo5jBgM2DExk2DYdUG
7nmKz6YwjzTfqPx6WafsMLsoCCDeY1UsARccmrzALcOt0eUb3iGrfejO23cV0VVb3HJlpOn6nGUJ
pvFfRbW7ukMrK8loYaC+8TR8Ft746b1cymhfGsr1bQ1/SNlo1KFEujcmo8EcNjkqh9EKei0W1zRO
/nqpKzL4SFC2ygJiquPX2wpVZ7Gm3gxC0twE5Rzpq7KD6erer1xXXo/AaOLfoxge2MlJepiycMy8
cB7+D/L/1+V8O16sJhot2sW67Vt7uh6L/W9G9DwNUh85+5VIltzQwcozTvPrlFDX6iS8jyouNxeZ
0XsaOb1rLz62LXLtjc+gJ0AxZrLN3YnaJxcDZ65+UVUY21BeMNIUsswdsaBiO3v0r1PwOAFNw8zj
w7ixBD2aeqQJQJOdgtJNTyNuSrW/MDrFV9m7Rh2TowA+DvjaxCQPmAJUMtaloG+6LQAxqgm9RSfE
PM+RbACG4WLyzEob6F0S3k5bhmhIXT9WxcV8y9OUslx6uLDw2tfQB4PL16thMh88YxEzyNAJPcK4
VpUjOXX1qcXaNFKShdUFYOAAbmmmI8dC3GVWsT315WvJd5ToDDRFV1BWhlf4ZqgbJ57EIpM7qXI7
At2k+bOiDfdrD0s0+D9HZTejQ6O1v/B1ggP2JiWBBL8OkNEwx2zkr1sWwjMTqtA1xxKg+0sjfe/M
ugO9WmUfEFj3etMTPu+YNN1mnO6Ey04cIhF0ssmoCTKSjl8ahLd7SCguGBV9MBehKc2FP6CDXbvJ
AApf0VxBf53Hzsn5vmZb/ITyGEG7O0xEtc93YfV3nlu/WyniVhPnOxyZjNPZGYTZLjL0n+P7VoI8
GkLqERWKlzp+7veHy3q+BrSRjicss+teXN8GESXl6Oq9C997TAcp8IXqqi1s/O6zWykedIm2mkPc
fpQfCJ+GBeWDT/TPpqv46vviWDYEoPueU0N8jpemESCivbWsCkoa0NXIYHeZdV6m8JDCIc5wusxd
QdCtPg1dVkxytox8pFK13mhudYhM5G7ywcDf4nv2tLGOwJTI3dYvZbdZI9if8wH0lZcPNwW6vS9a
L9KQ3MDM3wO/zj9M6ePEkuiHsly7AlM164BrZhdj5ru+Tul3Md2yWQ+UoV0c7MM7txsjwHvcpkYg
bwo4WZ+ytUVFG3IWWVzsdRC68yjx2Nkh+GLYEPmV+scGrbow6yEVKz9HvNlVZUL4WJjLML3EZQqo
CtK6Y3DycbqfITwtpH/ll1bBD8pPjgYqDKAfqa/FPWfkDiggui6b3SxO4dB9lhmmE5ZW6LVW3g6r
q9AE1i6PNO8eRhwq7MSuJw44nafR7C7aAcp/Yf5IQZL3Q79IubISVpSPgy97uOdEaqm6ceQ1loIS
sT0BkLNCoE1xEKj9Qnw+TH4OmhDVwBn2pXlaDULKhZtN+NyJVp5IAyD7G7X31wrXchWwTlMU7bnm
2viBgxZZQrmsCmHn7DkoVTq8T/zVVZdsPV8mNdnN8y7Cu9RqiKXpvPQjFeE6JgHXGfeRya9A/Erj
IdBog91tpclJqgbxdQMkpUa9deV14iX+fbw/tMBDHWB+6zu7J1U9tG5AQ05CPbyZaa1nqDpsiCFI
hfUziuCbLkStH9YjJuzpEWdGkCuky0yFJv5jyt82RgzyIo/BFJruz/M+dzzBNDCGBOjsdYK/PIRO
TvXdF1BAajCR8KlryaoiqT5SBJpOiuPpFpXxXfwgyUyK0koukxctoMzw/2DXJDcQKunA4ruji915
Nkt17WR1ShhXn8/I9PClSVZ/jLvW/WecDbJ4RNgE3jsxRO+lj/VET1rEFEbbXoblebVUw0xlf7Ke
x30Ye1geOQVS2OIjOlR8SWRl9IqV/sEAshjvRnchLk3TCzOm2nR66UVJDBfPNlgYdz7QIBRVKOTg
cSvbHyoMZL9XGVJ81W6R3G+W0Eddnakxmwp+wz/oSURYnURzez8Pq/iZjxExA60agZ8TUw1IolC+
LDdyJ3IceEVSs3ah9mmJkyrPYawulyPcAmXpphoB3epkxZcTePlm9dKVAIEuZ9uZZ2DiYStRkViV
+F7j84WcWnJx9fllFBlffi/oBimvn17lr2V4vuA3qQo7KSZ50KdyvlxbGrJygChUMPHnwLSAutrS
lKepXIkz893++lxGQOWYYL1y/DzCyicD+O0nz6gP7luCb6JuFzR9xuykF7Db/p1+cjHrT/plwWkr
Hjwz2DAieJ8cl/PlBe5y3SFxMcJN5+E3VTEIjB/KNSHGNlmUge/c8wd2dBkaRJjcafYoBuZS3uvM
eYn2MIRAzwNZMRzQhesYKuJFg2SOrFHewMerwcv/VVLQmBTAoXvLLZc6P30MYyvB6MQ/8n+y/T1H
E477zSW89l7ZAW6osTWS96Gx4XN14NsQET/j3CzUA+EeNxPgpO/OBcpJSd2BmGqtWAaA1fU6ACZS
c9iGpz0izyMpz6etjt0xWeERLqAkV9muxNL61WyCFXLgmsav/3hvFcJmFDx70u9qiwpx+i//j7og
2VbwAKQEk9VyPQTgSee91JmzIw8RrjsurOklR2/uNAmw/YCZhBeTcwDXWarHLUSYSSD0mhYu+TkS
q4bcOWbtNShHeN6OjwY1i+fotVSDArb2cKWSwbmIBcScjLTos5HRNE1W5wN3ZyAkeVflKWdlsY50
7+dEw+GY/sDBGCb65WzN0cHwSvr51j/ycqUuO2NnnPTQzEHfKkJiwgLb5JqDLJZRCS084OZeaqq5
SAhtO8Zz20deh95wM/+O7wuU6COtarAZ0+fl8Gk7JLXntK2ZXppWHEgsuLOYKN9kFYzsF88MARyn
6CAN1ExacReFGnXIOZ0xd7pYQv4ZXASWh2+u46XG4Zfp56zrqe3RCabul6AbuEeu6s/QmBer+BPR
7TsBGC0m+yi17GsNIGVu1ftFXuvLfe0wUmysGy24thTqv7s/XoHqzI7NqP4ISgBf6zEv0yBlRgW/
+QpBVdfuCthqhgecopCL7NaBNH4iYoj0WBs36BsI/VZsKcPbyLLhiLnEYS+MaG3NWRe8lqt4KM8I
n7As0ju3Fxgm97OFdpDQORyFeiR4XBnS6RJkD//MRpK/DW8/Z8oiwVTa7i7QFPGyvOrVfOncMj4X
v+IVT0XhG6VDS9gjY3zm8dKgkX90/7s4ioILDjiYxeIRoG1RwKvyHByWfA/4Sxo2YwQQ1grSI+mm
mNtIhp+Teo6dK7SCHVf97eWDOMM+vZ1l210sPAL8uej3JSy38dF6OByMnqlw2I1KT53r2brDH9SS
/+MFQ1xg9sNsH4kBKt8oaIBzb5X/RD5/3ef0updwbjqxC5fxM7KcZVqUIKj54eX93JCPx2J2p8H2
az4a9YxdLR5T+apJtsgIxqfovorq4MMBRfUJlU5ZCVVUFRlBmruXABeN0d4lrx8xtSPSa3MdRWu2
iqi9Us0MkxXK3oPuAUIwMTOCE2fhFbcezy9KBkaPBdoKBGdDtPA8ORPztfUvTVWNAb1fAno4NQAC
JT+82wPyM2X9CXlbyZ5hQ9jiKUr8w+m81OMZJ4ogEOI1kwTCrxfdMA+cMS4adr3QiRp9eb4Gl/dI
ypbk/VW+QW3alk8GbX32dJBg1GW6judXguD1bergtl9v5wrDgBlUXtFSdWsZppaPnieqLyqIlGav
rg+lVsSf2LYdYpRoO7TGHaqb4XTzKQ7RdPyamL8SZHVBItCpgsCWxD6akZ2nkkqTWfbKFEG+S/Uk
ceiD9siAq/BfZQ+kI/xpCkNV/5xpcpVMSbK9WnRdVjFQjdi2YRUN3hYe0ISDaMfs4cI5mKRW0kIj
50D3IBMqpRW1YjHl2KHGtAhPK6+YUZU10bSqjggmd2NmSpXUPf6BoZOctOeXfUK+9O9cOmI3Ij2Z
vzJLrgJz+w7gKyhsDCAnn9gd00yP9bkqnocze9jToBoIEqeCG5odd1BQS3U7RZLFr1+Gc017ab0I
oGu6spt1923IroB1sY1Tu/nRmPM+BEkPqivb4BwlL0phJvrV+U2z2ZLidSzRU3RPOTNMwspwQHQe
kWorAWWGixqVgOZDA81IsNlfRQeYwAC+91BSclHWOXcxd8/oAF+ngzm+jVKxEicjhzOEwghYmZod
TwE8CQMMA8jNqfCjObEiAaYFRf0phIPf/eifgqwM5FqfaDdNqGfoQowj+4S7ZNFCuiljibBQaBCb
Vncyx7L9kmmkGhwgYAwn/aY90DzRTgUTHyFvB0cwrVryXNpD8hbj8H5Jf1/FZDm+lPj3FJ5MT9F2
j/qoFHEeriSlmvYe93FGaTGkirBoDJVYkwDcHPInkMyiCH6gQZVjb9YR6VDEiDmRprg+wpsPHIGF
eOlxRiznMELF1mYLVFO9Yyyc0hWcfwCGxzHHZ/kzCQYLStF+zg70Tj987XTdycrjL5PmmZoFZbsU
NH6ATb32tAP9b2pONzTNZHmeb6dR5dDaKl1AmsRnyY/0vFapb6mXyuhzsfHOSa7hOdrs/f373SQW
qhqEZKUxHBVA4Z3zCdj2COLDRY/Q97TLO9LrtKfVS36vA+J/wDaXGazsp4Vg3R9RNLae9z+mL34w
07R4jzaXNQN3GdBJ0lPx1zhxqzMVUc/x0N30V2aMJb7vfTsZ3MMj97QFDe5tpxElcVp6TDg4Kxa8
69YxfYEpQqYp8HzHCLwlQwbXunqv93ctJ3WPJch/wmYMPFEYilI9PZ9LGC8nG7Ivrg4Nw+GNEamy
o0VneUtsHmBkOnC/vB4pzGZ4yPuv44Q+z5ORAPD+//h53SWMb08+a6wyFcqKpJh1OHGCYD8WNKZw
kdOdCvVm2ngy2HspwVxHAKKH2VH8xe7ibXVXiMMm1JSVuzN6kbEgAAW/lFkvY4e8jl24/ZOPtdHM
prJ78lBlF+jaJLEH8tViOHdEOXlgIYIQR2GNnCBEePjKcOghepSQ9tj4Bz5lbJSxNxzesrgP/e1T
JxdcpuHdlCEwgaDbO/T2I9EBevG/MV6o/+NWbVyS53AC+GgHFuUuuNXygSt7KLe/kAHoEaS1MB1K
Wkflwk8TE6cTXE7hZ6bWui0aZ1IGpdU7qVRoamxDcc0iNLTNm4srhqTAFlSFRguueZuhbnhIJJPI
FP0OjQZER76CTc14TmjUrcNbzCJFDtGjfaKV2xP372htEgfA/ni5yHlX5XR3mrc1mloWOtYjrsF3
8BkW5xJaF+iuqX5YBCYY1RyuQNUtceekh7F0Ee3gqM/+FrYXP7x9HiPoRtN9jQE9P38wrzbOdyZr
Gbmh3qDDi5LdIwAUXhuuSvCPUxU7Hpu0ZxiEw/M6N9mCxfo0E75X+H0LhLIcGb84UAyp/ZhN2zhi
Fl22zqywxoy/ZViXccAJd2VvEoYrvYl7cq+x0bCPSKEcK9UBhjka+A9XJQOfT4SbwBe112zEV/He
jBMBUjfhnh0AXl9jJl79DC1A4ldKUjb7cHKM9S8zJONsQ5xMlzaQtF+ABIRZBO6yl5BBrj03a5Jv
Huq/Xsooj/leAln4OxQ+dv8kAfJOVjK4d+srhrWaKmN+a9TJNhK01r2++PHIoYpYwvH3d2LVpuF1
hcmqOVgbXM5ovdevbbUt42e3h/UmQUg9IIema53ihJsoy4rSLypOfOPNeT2M89AUhbnTSwEEXidq
K8KSZiWGXF3o5L67VFX4yEou07OIVklep9VuCg9qBGeMQGas11R+2GjV1ql4czYnfP2M6YUZkj2j
dslsqhIOYoC+hJBuw2B/cDwtmbnN1dvPewncNxIFJkxT4ZO1+yjLqilx15loLv8zUqCDicBNba1X
Weqg8ljNQjxmvVSgy2AsEF7bw8BMxBaGsKcXrBp4fk8rFr13+Z4VKKS3jUaXHdW1CYgjraGHNeuQ
ApPl4i4u2umV/dB2xgvizAxh5ch+qdB0f248X+NSejZQfVyxT+Z7ER0uLdWUjbD5Wtf7ujjhnmJx
/yRla4C8d/GYOhHAHAiiSHr9XMuRXcyfQ6A2oOLSceZKTtJg3GCg02KzJxzxT2JlA5pB9wQ/IuuE
FT3R6riEMP7DQHdk3EZEZMsGPdL6fH8mxejs+srwsqc9r2dWFNK3IVmsil6hFjlbyGyYtvveEXbC
yGa8+3HfdD3KtRypqkSTkv/BIHZUf05lvIvOiGbqmiGKEwW1pD+sG/c4DFFS/+MXZFaqvoapOWRu
9ho0bSU09cEC1fAU9hjaTm70/UjLy06jCrJgozgYJX8gHwBZHkpeeWv2Zyz6uRHFZ4UOtNUmoHFU
P08bSIEQA453Iq/oHrOG73WTT9s/4JROIbmwK0lhloYJAVrJs2zqmhGbTHUHGCcA17UnnEIf62B3
3wXAJqCllf8ifnirmOv7nyHzWvBJsnAIqNP0jIyk12dVpCeV3kB3YFJOphczLPRU7iq6vJuRSe9R
PsXknFGIIisY0UHeOgVaOj9HlRMm+u93juiBtIDjhIPCja8Ot+wsWkWrzzB5P5KRoboQhqNgtjju
+NTdZee4Hsq5bR49eEibnPjhwzgkIveyYnK/q44ayujZqwjTNxhFr/iqHmit8uqB+kxdSud0fI7W
XQXLId077jzK0B7mbnVwiyX5MZNqtbqNB3tlM1b7SpssF+IwnBdCtP3uorkgNz87WF0Lyp7fjpb4
xaoWsCl1rPYQeK/f8q1Omuo2Wl8Ef2bh4LKLU4PJodH+rv9pWcEYPFkVfaNu6KhcHLkn+gWAAKM2
lOp3M3MmoG5MpzxwEKYJoyrFX3aU8vswbJkvUBaQOAZMyB5Zxc2t/Tu68huoXAZS4YbKDD3Udcov
jrQYBn4OH99hdDZpBDHw4URg1qPA8c2hf9Kwx/vCs27NGSNE/lbfcKB99HsljbKDc83NuDBzYxyT
/aT21z6Lw0Ob59Pkh3BYqdzjZq1KMSrCtYaffa7UFMp8PPKYCnKGPQhNVUoo3NgFsgqhoip6Y7uB
Phi058XGsrNgV5kT9N8PreKhWGExhHzWu8e2uZxfh/n/fsu6eldbdp+6KjFBrcUPpbB7Q6qANuY+
cpTMnLBxMdaDCaooikXfVEa62vG84O89LIXpNyAcbwSQ3smXAYOHlZXlAFE891jb+bgrA+Ia+Sdv
pClJGud1BUe14ZGAT+efjKiTCBVN/cIKuRmErF258bhEwG/7s63jfN8VzizJb7g9PUqp81P95U8O
R2ufSbCYeKQdvpoHOuyIuBr4C+0FJDEhVOs8Xdu+tqpMqu0pa5iI/vInMR9Q4m2njxb2Q3tKoz9x
OwVUSTOVs4U1jEdAYTvDS9mBLcHAuajAa8XKdVmgRc92v/VnTCH7SWtjn6HrQrAl+aqNe4TqmYcy
hpJMNluHasUT3niXkGCkP/QqxGqR2vj5cLr8p9PRxmdV3hKZfdsEMGVKF/u/yiUd+YpaND6f27QD
YnaQgIywP4vICCt/1AImkZAp7IwELd3hvzUY7VjTr0eMOzZrAouTIPTNJjBHURxpjM+yjRtDC4X9
4Yei3GQiYcB2XTxAEQZuFjwKDsjW4paz5Mb3Rejy/S9aWF4+nwrU1AxRY3tmAMfxkBqPbN9UbsQO
V5vX0tfiyz2aAQxXhk7sM6Rco4QGx/dfVvWSHLKIZwHr544zd+JpKVTLaHoyEzGPvdNpgWMS+Yhi
4UiRveMner7aom9+N/oDKUkcqcOFuUdam4GYQRZ5Mq0laZ8Fcd1pFGFcIOVQ50Bwy5PSxEF9q3/V
TnsPd8NwTqilMOn/QezyqvOQLby8q4WpNaZVQXTNir0F7eSlOzwXK22jSWLKg6ESOFqltwxtHNW5
EPN4NKo9Z3wayERkX4obl3tfrWvGbRJ+KlG5YQ0/d8ph7pSdpKS9RzsIcYI7LKpZ9f3/n2rGH9u8
eJNUFOo5U4Vsp1F6lnmyXyfOvmJ/GdoyvHAQbnuBYLt2NPX3rAg3LOd5Q8L3sqX2g3d1up0C5eHs
RMclaCkaWOepBY7Hxg+FPYcoruyWSgoNrMbKEXAX+gBnBHUnDQbHXm1mzomtHXmj7W65Vgn8/NXR
0/Tw+E+i+a5epG0CU55aVLyIOh7p/aBTx9TI9wEzCcJf36QzUzWgSkvr4Jvd7Krg32fKkkToxYxg
hqDF9ySQqZuU5BMMYbtWUPgiPdXhvFwPexQtP9LZtsxbynwUH6TYm8V8MqcfIKz7ItE8v/N4YM34
fGawqDyfMt3vhnCEZu443+U7cRyTlPobYB6rPzY0FSwegoZbvbeN3aR8nN5d0ANLwQt1tR/103kn
qHbsuZSqfQodYrHzxThsJHxtvgOqjkz++Ff6AeYa0NW8pzx7Y5ga3yRuhKT0bIi75o8+Ruyd7c+2
vdrLDp/ID8mYhkrjh+LWWjbrlsTq9JJFcbfR98JH146Kb+dluP2JP0/DIvQEGAbO28/d/ifjaZDZ
0jftotDch43E49u1bSI5aT/NMfcjO0MKjaD2EYqbU38yUOELUIHoRsv7kep9SFYraRe8wjWaYHBt
VnGcv5EXECHTZ2OVjZLAxCI3+hBzb9t+AMbEOumNQGcL9d4/eIlLV92BQEtqc6b2cHnx57ubwzZP
bkPhsogA41tGr8roPtsp1hJAJXcL/eWMIiVUqq7CY4Bfi3DRrPBK6wsn/J03FNgbhr+5eKEIavUT
tVG9z/ZUTTKSEqemhM+0FArgG89zbn0ZjCpDOdbLIWSDOxkz3qtnneiVbtavMmLI8ck703wGsaM9
EyGj6CFdw6rtHIGm5c0lmuFPZZIq/9j4s4obDG1Qun06hJczoEmrSxttWqRDN0FvKwoSawRDHJRh
Acw7QC8Ul1UIePp3t3g5r2eYeiQLcuUs33Gg20nm5EqOZKtRFOdSYmKQNLhGBiMUky5uk+AsMrGD
HCWxHNB8HRjCa5BLte3LsKOhDamRDu12whk931sSHlkm5XzX9vxfI3csLJOuJgjtjrtIF2UfLl5V
KNY+XcJ+BcvXPQPZnFUn6xa5fuZM4Ig/tfzxHt9vmwdvmb5zvswtkbs8RBuIV2DhU4KyMrf1VS92
h2XsidbW6+fkQOKUE1Q5NouiwLaMhK9quactmdC4VwJl+z4opXYok8Br59XiwRuG/4KXhi0ZfnCp
7rWI1sv3ign+oaokkEeSQdQYTKVvmsDcRsIQhDwFQmo8hwZqE/z8CCizuTdiK62W+Kp2gilZlZKl
0NxuMGoeqXO0U3fWzsgxSXvYP/zNY4aO9jCx4ch4qUzsYCRTyFHh5KTvybi9WRfHxNsfaZOxaPqM
FS8lJE92Fo4/h0HufI78DrXjnq82GyUQMOc957nCvLjDAVmLKHm1zKIobXrduouqgcHSol40W5FJ
dZxEPC3uJwoaSC53wxqRva4LQX+Qy8Yg337ImIZ4GfhkR1GZuT7jCEEWFZJbuNhQFOAIxEMdL9+e
kDC1bhSMxjkEfcGuNdwIlTSJABLJkbMGi1gsKoOgTM3eCO/3ug0=
`protect end_protected
