��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	;�׋��oV�cŕ��w(;PFt/����NZ@N��H�����x .?(�D֮�8�y#l(;|� I��&�8 �� ��?4�}�n�u��D7���z�dּuCe��+��{�vRէ�;j���Bcl�Ʋ�U]oM#w����9.@��/�N�!�^�DI��T1���İ��+�c9����.mhu��R�C�s����cGF�Y*�ʇ;�0YLx~��b�J!��&�J�{#l_$��`�;�m圬�Jw'j����H���s)!�~K=���褣�`!�ds��)dk�U(�<��xO���>��Wu��\o~z�
��_�5�b;J�ـ��R0:'�ɾj�[�oČsk
32m��l�A3nz��l��Yt�֙շ����"E�!�r��CZ1,���G�}$urun��@D��-�X��e�2��%�j�Q�C	���&�j�Y��Y9�p��bY������*�c�� �k["� ���bI�{ʚ�k�7����Ӗ�l\iI�!�2 ��t��9�+�a[o�����5~̈$�`т�!;� ~�*`A@�� ���d��w����+��X���x��F����*~4�NO�b���������pD�'��9gݩ�c%��6&�E���-i§��W��ݼ��s�sZ���aJ�"1�Nj����A
�1 �d�����t���!��46�7�%J�"S0��d�Ir8�M�!#<?u$j�@q��&�����$�v	t���1��PSْ�A�Ga�Z�	H|�h��"��2��O4N��!��%�NV�i�c+w�����0|���\���F�"������x�qܷw����뫥��ŌxL}�J�1���HzD$������<���/߱\?FA��t+h�ė�GG®�maHqW�]�qÌ��a<�����[�k�����$�6���߇zᆦ��y6����Nܓ^��	�	.׀U�T�3�^Lc��<'��#�)6��J��޿��<��^�Շ���q��d�?_�&����CgIѧe ��6߷�'�ѣr�d�h�.���^(i�L��Ic\�2��
[}�&��}���	�*x�YCc�"�Io�Oè�-{�e�`:E%Mq���Xi�Vų2��̅��,#.�Ϻl[��d��vzW�0dxj�sx�H5���k��M<��-�A��E�����R�kǨ���n/�S.��bm���4ʁC�"p����=� ��A����' �J6�]Q}��������	7 ��@h�؆��mv��ڀ$LcM>�F�ٓ�7$c�����Ao�@�1wr��bV�VgU���C��ܳy�w�� D��O���$˺s�H�y�q�Y�n�K&/��@�L��T⣚L;*[���1`�F����f��nU��DW��+���mh�M�������f�~�^�\���NE[�Fio�O���`d�N���:gce�9������a�%��C�oH�Zs�"JG��&#o��A��M�4�����@�6�����������<�(���p]=Y�2(J߸���Ct��5��;d�F��d�C~��G�i�Bt����_a$?.{��Zl��ɇװ)�|�z�Nb��>��@p��t���]��*��[Ӕ�M�����G5U;��g��%�{7�s�L����9嗩�"����ҍ�j�����*o�����g�]�B�By>�)��[H�=&�^Dr�g�N2K�.vB���,��Is]b��u3k���$���-�̚�Hݜ�uf��0��"4-N�uK/o���Z�<�
��B���7�U�B��:N��y�gRE^�s�xZq�>?T,F'�mqx�v6I�f4�v��@�.��YW����cC	fn���ql��s��rפN���s�<�d�<)aPR�k����� �u�>�hA��c�UO5�/W��T����w椑j}B2���(�W*�^9{�t�2
�]pq�gi��+�{����.���7v��$Ni7�qY{e�N{+a*�R,�^�'���{�Hn����=t!��\�:EOd�g�ba7�C�h��Pӓ�C���E���L%����ko����k��h�|���-�A0�7]g�Z��==eh��dM@v�}8'hG�"P�K�����*��Oz���{12�̍����:(�L\�x����@���-) ���r�]���������`�G6Z�����g�&�笈K]��%�%ѱ��DVK�6��K!�,��,�ی
���ﴴ�n
 �xyꋔf>�9���n�ꜱ[L�J�ֶ8^����Ӕ/����e��	}�1Ȉ��7��.Fg�J�>X�]�������8$�U��&����+��;�x�>Qx������
���@%�������d5=0��A���|rm��qG����i=�g@�,�u^���&�<��Pi�ڒ\j�7���������EH|�����~5pq|O�.��_�SV�ޝL�Z��������6=���`�..)l���^����G��Kn�V�{�_�T�{��a����=#O��;C�cL'���VOƸ�9�j��D}p�C�=�Z6��Mi..�(a�'���e,P��@��3 �/�2_/y���ײ�l<:��֧�]\�,���ƪ��?�F�_��w�$ԥ���흳�5�ڮ'	F�(p
#�d �mF�;��h���5'"΁�����
J�{���M�)�b� he ^�vݚ}�ұl��dl����/#�N	�ɡ+[MN�&N����r^걁��\n��t�NE�=s����+�Y��XYN�ܫ���`Ķ���u\��������N��r�k"?S��X/�+�����<: @�*X;�s�3b�KP��X��������<&7?����"9��+mOPM�J�oЙ˪�m{���Y4��,�=P���F�� $Z1�)=Ѓ]�� M��W�":��8��yߠ�U��W��Z�v���q�Z�g���*��=I4��I�A��;�B�|0�9���2���ݜ�F,
~�tf8\_C��A�~h�x�<��~ gay�h�;��+�&*�F���)w������i��.,vE�	( /���J[�WiP�z�K厽8�(�.!O�U\���{�j����ӿ���g�i�0��T�ͅ>��V��&�U���"#�أ2j�a���'z�2���=-�z_�Җd�]}K�w��(���7�<OEC�r��5�Fv� �h�PM�/��	H��`�z��a���#�/X"��'e"#1$ AS×���P����F��-�Kjf���Қ܇��Kͅ�4���	Z���g��xXQ�r�}%6;��'�F���D��Q�}ܾ�������қ9��C qs����ɺ���5]C��+�ɑ)����9@�~'x^l��iw4�gI& ��
_����,�)ћ��~�f��L��H��VW��4��p� G�痠�H�N��tt�ox"���K�B�?����]�D��fJ�@���Ny�e�/]���b����
��v9��7^�K�[ч�R�L��X(�YJ�sl�Mq��=MU6�GV}P����f��Ŷ^閁��D�gݤm	ma�XQ�vyrʜ�[��&v$VvC����F���u�������zux�&���7��tS�Y���8jTu�����o$,�p��������.�1Z � ̆��N�}87�0<��	�7�����X�����L��%�����xa!2 W&���0C�@&D�Y����b�@@��oC��FhZ~-��A��ױ?_�֭�U�sCl_�w�4ry�ϖ&�(nhן� I�a��=��D��a� ��\��*��:��(#1�����&1�vG(��$�&�̙��ib����6ݡ��2�1�D;�)�`�� � 𔰏�?{��TF���j'l@3�;�"�ҧ1
�~Jy��
;$\�=��yH:���u9w�����	�_�
��$����&��~����r"<eκ��ްfm4p��x���9,����8��𠻓�q[Q�!J�0[��gR�Q���:���/�kKÉ�Z���5�<��_]u��t}�^�;�;�N�]Q���0���v�Y��S��xb	)��Ie�<�FQV�[D�KtQ�!��EDPX�/.�Ӯ,8b�V��o4��WPk��~�����!~��g	S�r���?�O
���YƱa�=O�FĲu�ckV֚����w��)�} 7�y����/�N����y�_^i�1fM�<fNG88�h_wZ��f[A��DK0�o�9sV�x��!�r6�U�[ئ��z
�N�/j�n�a�7'��
����қc�츍��%b��:�������)[{Md�4�Ox��3R�mJ��6B�<q�o�_���Ij�nF�op|���/�Ջ���/u��5�ٺ�wl���w!9_�c�D����}����wi��1o�A�.!Κt.�b E���_�����e�y���T��3�S����B���r�T~���{i���"�_��#M.�ȭ����fΦ��
>�<�p�Af%i�c`�h�"�s4'����f����M��vQ~�f6�;� �vُr���o�nT]3Z�X�[n��}B(?f[��:��E��sL��M�pPzk�B^��c�-��[~����ň
r4�Zf(jǿ`�*��,�����8���мK�~�YH�?��]2�t�l"sl2�x��`���O~J<��"b�:`��|PIנ�Mb��;���0'��B������<+��׀z��Iw�ߵ��Jب��Q����E!�{#B����w:J2UQ,i��5{��*����#!��׼K�]#��Ku�����nD�"��D�Ebㅾna|I;<��3b�x7�i_�a���I�"?rO�ic����]7�L�e�c���I�Q�Ot 4�lD�.�yn���u5�З�����˱���&�6�-������
PYJ1jq�u��մ�Tz/\�3�P��7[H��oY�}$'��֧vFy�s��
d<Ӝ�>)�����7Ia��Y�V%��@B��[���^���V`u-ĭϒ���?����`2ɦG�?Xuӈ]��/ؔ
Q�p�
9��a��|O��U���_<�Ѥ$�k��6Ʀ��������Q =`D��wĎݼ�[lYq5���G���W~��?�F�l��Cd�о�.�$��*�i
�r.��/��f�
#�S[:6�>DNܨg-�3���s�R9̓l_$����ܛ*���\�[f�vݴ���Q�H�^�?�Oa�"�KTS�xp%
���u��;�vp�^���B��k�`Z	�_E��b���Zgʛ]&%DIH�{1Hǉ݉�LlJo���$Q�����V���1���G��V���7�)���/��h(�@?�ѝuʐZ��n!�s�_�7h�����i�B�I���P��v�Ά9^��H�b�t[�}��#s�FUU�׺�0[r	�ZLn���� ~1��0������W�g��;��x�M��h�9�,��5��V.�3�o��H��I^�S 7� K	w5����x]�q��;��V76Rn�� n����pc~5�JQ׺y�2xV�����C�3}�1�|
8��vx��K���9l�X�/'�V�78Ji�n[
0��/�����u��V�T˖�b�|5��0�!�/�'��w�x�+D�%�+�7��!�`j$�%���2ǻ�I�z���)gC��N�(@�&d#�F2�\�������}d�pm)YO�Хy��fjp��q�J��v��n��U�J� g20R9��d3G���$�="�:^9�ӡ�{�Pr�e(M5|��ܑފbn�o���&^�D޴�/����"�(݊u��M��O[����L�B��}Ȃ�*@�r���I�2屑*�Ч�?(',����s����0��Uۓ��{��#&�q\��oʂi>��.1�
���"�Y\Ό�,��63>���uցq��[6��`WaZrә(�D�q�#O0����q���s�ޜ^�T(|����_�3m0XM�,T�/�ߛ
>^K����A�1�Vq�`P�y����ym��6;����s�g��!]+���8�*�1�JS�w�_R���N�����d�'`��l���»0:*��B�����<���F�ޑQ�)�oF���_�#�h8o˥�R�rY�=�U��
��[ uq�AU��ֽ�:�覃�z���J��J&���O����a���К�?����0��|.po[������^{��z��g�>����R��"E���2�9�6���KAI|u4��N@�S~B� %n*_%gM�P�lDюnH55�$|�*9a��#�{���|�MЋ���~7q�S�E��*��A�d�1|$�#1f6�)i�Xe�U�&�h�GG��4�B���ܚ�>��!�,�e�N��X���=���1��\%yY_.�rJ=�,��Rl[�4��+ohp���*�=r`������*`qڕ��'4R�=���D2(	y��=��60>�	m� A���#!�OA�np7�d����f��$�O*��mE����9^���b`�� A��(��di�)���)0����G⹥��\�������n�ɮm(iM,ԀV�H�kJwY܉o\U��,$�ވ?h�ɻU��A^���9�Ml�fc������&�^�,�
�?�MAK}A����7��3���K�;��ߥ�c%#)� ��b��RR�����K��r���O�_W����#�Y�W�6L�V,2��h�����~Z���!�ZRF<��D1��Q�ٽ�"�~�E�zp��������TZ�(�g�2.�s��+��r�'��E't��[֊������>V4��h:�h��E�-e��d�@2�]���Z�" I;�FL]�B���l�q\���x����+�S�����ҏZ��DC(��x���aPf�/�P���z�-�ni
K�(�r���ԓdc�L_�b�Ω ���8��K�)+Wd�7�86�Ţ���N]���$$L��7�#%I<���[8�{%�U��Ы�+�m�p���/�a|���R��3������ ]�+��wr]�+t�{h쟀�F��ڻ�Vݺ�Cٌ+�N������y���htZ~��tU��;�"J�*3s-~R���L���WeJ����M�cθ";�Rtw[?���>v�S�z�������Qm��j{#�������)a~8�� &�b�� �9�J�@��j�14[�o: �[�����>�sg릺aA��.��hn�[1Q=\��X���D�$���P�k-�s�H�h���#� mI�ɿ;��|�e9�������q\�qXtU�.�l�-DG Ȝ�Þ{�?��6M���\�DM�f�ܤw��R����P�����$�%AVP{���6���5W�=���j�2�z��s�:)f�i<��c�p-�g���%��߳@��Bz��ǶHV�gΞUr�v@.�>�9��7���,�2%F���e>���i{��؛8J�1b��n

�� w�|v�^'����G`ڽ+�Q.K:;%��7�H񸬬f�9�#	�ioGh�}q��J��L|ۭ�c�g%>��!���"	3�,���N4���-��_�~���P���﷕���1��|�����E}����Ԛ�>����D�G�AZ�!I�ŕm�1ˀႫWu�.
�����i��7z���G%8���/�˻�O�h���?����5҆Oi�&a�A�mOz� �6Їʱ��6�d�c�L_p�#p�\�~rGR�G�����=��Co�㱛M��:���qA
��j���w�_�(RQRp���de/]O�����Q���7L�>*=?����b�	���_�
1s.�G�O��#5��'�P���9���Q�z���l��9�r@tt8h�fݬ�y��19����'J]���3�;|]��[��"���jO� ܏�ӷ����b�Mnz�m��v�����(V`Ԏ�6^j%Mq���"��J�;�tC��8���1�"�����Z����Wa�	a%���RH;���͒n���䴽�9#�����EB��
�3+U�LW��l[yZr�^P��K���&/��u� �v	/.�����#Um"X�ʡ� "���bS�n~��"�� ��L��b��J�W%� ��#WxV(.0~�q�Z��O栱?� V�h�EU�t��+��!Y�ǫ�j T]�4@��jJ]Y<1�_�'�sћ�R:�/D�J���Z�&sY���`�����8�YCms���ыZ���Tӿ0E��|�)?�Mב����b��0���U�bD����Y3�P���τ��匌e��M�sJj�ݏw�"��X���������	�f!���I�j���b����2+����"��������<�8qb$4j�<�QB@T۸R��������'�`��8yl�vc�y��&x��%��W�@N������f�(<�\gP6�����UP��v�IΦAKx�%^�{x5�+��2T㋥	L|���E�>�}��aՈٞ�'�?�=,_C���6������"�"�35=6VN`���l|.��X�w������	�K��a�Ի��	j�#m5.�N�'�>��W�.�P�b�^!��'b����210w5��4�J,MJFdt�Fr�E�D��� �z��\�qQ�
��0Ϗ@��\��V����ZFǺ;���`�l�^�)�����`%�<��e�)99�H�+��B��i�Ø������6�w���xZ�E�����o���	H���m4��y�p�=>�UΘ/�)v�oS�����9"�8#�A���u2�����iY?2�����ܘܕ<5�|OQ
�$txI_��K����nDO�F���<��Ԁ�?�v�yC��{$���}�Ѳ�� [' ��X�'�H|�P���j���!K�Έ�h���y�)���u��Я N<e^�Hk{e8pe�(�2�d�3;R|Yc�_z��@
�$�C#�}��4#�x7����YE��>
��Ʃso�(�ʚ}JW�����2r�rn!�����k��dY&�:3|i�^��:��V����R,)��lr�A�M�a*�����{`2B�S�/H�˸�Y�}��:®�Ë}x)i�=6�@���;H�O�3?���}�ekt#}u�������Ѥ0t6�?��Xe�n@���� s�sG��;�3s��Hҵ:�������	#�V�5�+��X��T�E`�-԰���g���bx�o��|�D:�^�!ŷp��Ur!Q(
)�F6z�-1����i��.�Y��Q���1ߖ�y�١��l'��|�]ʑaU�)Śi�9�=��i���N7{x\�BJ��y�Wg��eqFb"u���H�~���x�{������;S�f��y�KrO�gS���6@VȘUbT,�C������B㩧z�K�+S!�8,��ճ������~(ɼ-�����)��K�ʦOsYb�G�@���]�Tda[%r����/Î���_[�R:��6^�N��k�}�C��t����щJ�B��X1ъ���Fr.��(���8��&��l��'�N���m��iN`���)�4ۜ���c�^8.:u��`(�I*����)Ɔ:+T�e@�7o�:����b�zSN?!����)c�C#���bM���3<1o�7TL���E+��,Q���P�\I^SRW��x�hIW�]�"ɑ� ݸc�m �Pks�^�Դ=��D���E�P����t�<�?�m!��F�?�szA��� �@F�as�T
O�[&�������t�*k������N���^7��j�ϝC]��c�rq�+�� VX����\���k��� K3* Vce㎢�_��a}�L(.k�"/����:��̸=5Ð��}L������Γ:4{'�K�	�fǰ�u������]��>�K��)=�΍d���R6 B/C���Sͪz�U<V���)�5��aw;$�C6BT��������G PD�z� Gt#�$�ơ����e���PF���<}���L �+��4�� U\�P���J��j���p��m\8ͭ�������8r��H^����(D���Ԁ�{���wkRڌ�ψ�#�T���S�Z����1V��Φv��K
q\aN�vEd��CVZ.Q�<�âxi&�m������|`�}d� �ńd �=ns05�8�qTT�j�XO܀˖W��|<�֊���#�H�Qi%��6�}쬝b��KM`.�^$=p�<�_��#�nC�.n�7�����X�z2�Z��<�>��r+��-;H��C0�a��l�,*\��>�9�1�$jr�@�6���熊���X�;q�B���9�w�q8�\����|�$�nn��KzI6@U����SI����iʩ���B��G��*Z8����Y��U�>��G&��a�}�-���%�ף�%۶��[�k�Vkʃ���n�������Π��B��ȧV*u%��%~o�i�Q���uQ��+�}皋�i����[)e3�.��=A����B��1מb�3o����_v4�n�&:�G؁K��� ��i3}�P���=C`2��f�Eh��qz=��f$�FkG��i�C��P�Uw�rϑ��Jf�5�R�{�m���5� �L_G/�G�$����d�=�8*-�/�b�KM3����bgk�K�@[�讜��n�(�8�6|8(�%*Nt�h��J`w�8*��~m?>K�a��:	���5���K�mć���Y�qj�s�WM(oq�A֤�����S�3>��x�~����:�tL�h���K�1v�v��Y�`��}�x^X'��~xN����>vC�(tPY|&����"Jk���� ro�4��J=L����Nu�l�%R��E9�%��*���`4rP�n���a�w[@��o��W?�u�7W���Ŭ�-&�5�������5�
8n\��w�����7Vy~�����\�g�+�ɗ�Il��љH�HR�tu�b_��69{���{֩�ZԮ�Xdh������mY���M���%�%d����T0V�!j��b����(Ϊ~K|l�A��A(�:6WpC�����7ǃ�(��_������vC�`r�'#^E���W'�$�s(a��K ���U\~hm��r��U�g�c��\I�]`y^�cx��)���y��, �fp��=[�}�����~�g�þ����%�U�h7�v
��*�~�'EUv\e�A\W��?n�M-dY��=��@�o�\:�D_8��!\�I�JTfLg4 �������mȳ�����E������v	p�u-}�h��V�4U�S5�1������;��"b��o)q�%�%|%�'&�����d�=G���k�����5(���̓��L݊�%s� �Hx�+Ѡȓ �7x<H�Xqj�H݇/^�>�`sJ���p=�L�J�#P���,�'���&FS�c�	w��̣���#7��ec���dWR�.���(($�9�Q.)8x+/�p5$齒���(I�A ��Nm�i�M���y�O]��9����-�yv�F�|���ċ�������ɑ�R;l'�A�¤s�`�P�����'su^��X|�(ϔ1C,����"P;juA�4{
�,ᆷ���U@Ğr�9`%��syDi���<]�JR}V��m鼴��&��/sQwd�ـ�J������G�UE�Y����h�L����7��'k:ϕ
���E������[�fq��0F�"�x�^����r�[�7��\�M�4�o�����kᥭ�\U���73���(��(!���OL���Ί�J��4_�PHG����i�`uI�G?��v�c��A�
�F�G���>�̹���V��U�|���@TT��hR�a!p6�`ވ���"T�D�1͸TFks}/�@�zeFH=:_UT�[CvU��|>pH����=��Xn&�5E�:���j��2�uP
��ܙ���|����ǂK����ߚ���lE����W�(Z��3�b�Ex�i �A�b0'�~;!n}���˟�Zփo��׭�(�!�W�M�Xc���\^��
���[m�wdǷY|�/��)_` �$n�j��ɵ�D����*�_��v��eW��XФ��WC�����<
��i�,#]m
F�_�L�2eF�2w!���%�� ��a@��m��y�:.%]ݥ�Ş�?ޱ�H;�S�k��Լ�>XYsb�T隚f�Ց���*�2��'=������s�/����&ʖ�pK��c��H����BJ��r��O�ƸM?F�<���4'�����r[�-KL���`��e��m ?�T8>B�A#�g4�9���*e����	Z����<����5����2�MJ�q�Ȅ@�T(�
�_?j��ɸ��Q$\�3�yp��/@J�R��TgOG���J�P�ė��V���7������
����=��|�lK����!uD
� JW���Тe5�'��"�q)�#!�+�F�
W�pͦ>�E�Xޙ��T�1}P�WJ��ؚ��t�������5J�d�j	�&0L�/7����|^3�D�_�'��R-��oC��:󊗊��&�s�bq>���, �_��CR���|��"����^/�K�����%vi!�/��e=t� ��
��_6D�ZK�w�jo���sz�?��ˆ
bU�`���zJ{�WEI�N�YW)w}yv��`������ւ�O�G@9����5�8���4�����@�÷\7�@Wï):��IO��6]��	+ ���U���9<��G��_�:m֨I*�����V�bq7t9Z��fnܸ���Pg�x�4`S\�: ��4�r0r��q��h��Q��{��m�	h�b��� �� ���St�YA���hd����zС{��ne#�ɺ���"+�F]9mis������HL�.��@዆5� g+�nͮNҖ\͕�)�n=c*��L\ )����]�]�{3�&΢�q������4D���N��nj��a��N�$,Y1�9�̧�tj��{��o��6�Ȉ��V���})��I�5ǙI�Wp�X�~ZA���5�Dm�ś�avy�JQ���"7�H�p�dE�p��oD�h��و̺E�B=QiF��ŭ�b٪����,�;c�=9D51����W�P�ŝ)�V:G�Q��L�/S��Nuށ��F��%�e�jx��h�"t���Rs/�����T��J��24	Y�;�hU��.7p��/'$7)�pJw�)r%�����5�c�4�f���m�0��H��Ã�UL1��.�g���i�,W�5�F����������mc�����9�-"��'ͨ�2mύ�x}�� �6��(w�;�[0O��%2��0 ���t؝�<���&��F�.	s�k�Dݿ��ε9�dc\D��*N�u;��/�A���7G��t���1�y�ּ)����G�܃��ٓ�;n�d+���Ft�g�B��eޭZn���qI�L21m|�	E�L(�n̛,)�c;��rx2`���4@��Z��Z�����c�	��#P}w��Yzu��7=�8�rYm���k�@6RC:g|d}37��e��e��C�h2��H6����R��a��"�!��	ʠ��w�E$)E<��-�Q�˫��MA�������J����bb��vDJ Amu-��D!懶eFN�h��{��T{�*Ղ']����Iӽ���T�l�!�����.D��pr��Mz��*=�B���3�p?旰�uy�h}� R���
���[w��9d��#S������}>��3iQ*t���.~ݵ�B
�,V���.���������DuS�'�붯e& �h{c,��,��y:CF��ep��ˉ-���o\��r����*
C�aĪ��
��3h?{ �Ua�7΄;p"Tr$��p����B�JY�>��r�����y�j@�1ccS�i��J0o���0��&���֥��:�U����n�sPm�v��QC<�=���^LP0�5x fF��D�9(�S�u5��K@OK���Ʒ}�)�P�D)�!�3#�ì\�s�E��C���[�4���e ��p;D��->@�	w�<�?�b�������գ��h_:���M6zO��Є�%	{"��%�j��D
�ae��ќ�&���&��/�\S�@Ab?/ARs͋��Z�(��l�"��ʚ�Ź݆!uWRz���g��g}���뵕WG��iN%��̂I�`��%q�k�q�$.��hď����]� �-�~�*!��VLI{�F�G(w���KLT@����R��|d1J����N���]>/�4�k�p}6�A1��r��=�s����	 V(qDw��5C��L����v��*dk6,1�zQwZkb�8�Z�ڣ;��2�W4��w�PT?�T{	��,����e9/�@T���B-�c�`�,��a�?�	m%��_�C�]�/).)m�JurOs�t�,��y��4W����\#G���� ܧt�^�Hs߬P4B�"U�*Pb����\�A�/a	 ����,YT���5�� *4�z�W��\�PJ�$?�?3k��_�ܚ�F8\{#��(=����O�a��jo�����,�>�'��(�����G��ӌ4���z�}�lע�0����C���(*����+��Ըv�
�� ��d$�
�K]�B6K�)��l%��������g�#�Y�S%��|���2��.P��d�Ҥ�Cm<�����
q�LϴG�`�Q{�����D]b�pK#N����r얶�Z�1���o�kZY��9��o�}&�S�&�+�y�M���cZ���BƐ�ĽP C��~'��I�S��lX��҃�����qi���gO���$��`m�!;y����oc@}ꗕ �f�_T���|��ئ���A���=�+����؞�l�A�vIdy�ot\池�2B/�%t�6�w��	{=���O8|����{��E|��kiX���hO����7�:"���0ğdJq�U\�5��l�)\�x�)�0��n��W����g��3쨵�6����>=&�4�j�=й�n�G.o�&'}3���h��'/m�?��{��%���Vv^��gG�M�o�Ҽ� �	"L���]TQ��)�D����=\�(��fܖ{I3�M�]�8��W�C�f(����G�d%9�N>IȖqsX9�/]Y�7�śiY���J����A�������%������e���r�R"M�i
cB�R�5�Q��`4���|���ڌ��m����iA�m��G4(.u�<.'=���\ �Tu�LN��Xg�m�D`,w���N���vA��Z�t6�@B�:�(]o�"�9Fϐ����$�L'�.L޹$J��<$ɇ�Q[W/��t�m#�-h���hzt?��wx���e�}��U28�=ǌ,#M�I�xRLh�5^�p�����΂��  ��w�S*�!�HSdј$�d=#G�D����2�<��>7�Rr\��O��b�L��  ��y,��l��}*�SZ,vc%��~�j~`��4�d!0�K�B�E�+eIr�B��90�C��Z�� �,�n)����G�	tp�*Iұ�ѧ+5Z��*Ե;~�BKF���t.�\�#1�lI�R*�ކH7Q�mSI��NF����'�t�Q��l���E�cz���V��b�j΂n�븡<����1X/l�u��^ِU�Aq��B��+d�ͧ�7+6It�������3������e���JR/4em;�)F~SJcMZ����]:�@����*?XhɜLҽ��}-�dj����Tf���8��rW]gM;b�n	G�@�Go[jqh����.�t���c|G�"�FeN�j�ū�q!�_7Gy�b�T
��,�����a�/����7�G�6f[ܴ�	�/�3{�!�k?�d[�3���2-_-��Í����yU�!m�#���S>�L��9�V�,�O?z�p!f�8������hb���<#E�݇�O	<�5j12�K��_:��=P�'��"�M�G���r��mM�
�ݥ+u9�ߖ3}����l�@P?y/��G�c�vi�m_p�����g�M��M���������m�[��˞G�-�ԁ��B�0��r�%�[R�I~6���QE�.Ku*�g��Y����"z5m�B�
7e�q�� ā��g���	L�EmMl�0���|�`�aE�V���es�)�y١�Q�ָ�lX 9u��`p�DNR�Y:������ɗ�,WmcGT�zێ{�������-u�C��c]��4�s(��P��kDϽ�NMIza�B�Omu�/+��~>_�h��a��d<2_��s�3&��溷y��=��3���er�H�t��푚��kx�u.1�O5��!�{�l]y��@h�p��-�lB3@j��v4��4��<%���y�JX��V�VuW�Dk�Fc��&��$Z��d�TkE�pa:��H�:a�iO�d� �9,�ԓ�\m�@�X���p�g�!(E��%���ta���~�=nDX�����p6*����i��2��0��ݏ9��>��@+\�ӯӔ��R����Wk�n��c3q�od�ȵc`�_� 銋}e�Ԅ"�ėsn�����ģ���=������ᾐ@�k5`�����Ӝ���.��D�f�)Ց��Q��EKԶ{K��q�h�:��`������'�����f�m}��PU'��gUv͢;�U����>����}t����C%PL�#ʪ7�D�Q+��X~S�[��̇�S��t��{�+�_+O)O#���새x�`Y1�9���v�>DY���9����{��p���ɗ*S�G��<f�����4몜ͮ�M�}��
���BǍ7%���Z�T�2Ѕ�E�,����B=e�Ʉ>��,>S7��b��6tg�P��	��T���|��6�h��V g^R|��xǵRzf^��=jr�h\�_ޞ������=U���bAiL�6� 黻PI���O���;s������-��aT"�p������\`���F�oyA2��Z��&|}���!>�>���$����������%����nPVu_t�O{���6��I׹����Ok-拤�┇�Uۇj�n�֛Y����v����"f�\3�X;�B���L�-�2&�X�ޡO�Bet7X��u�"m2;���UX�k��RϬ.��#Ja��)*kE���O�2ڶ&s�m���
5����lA ����K90�Vq��k}�wq���Y�Ho'�Z���j�YӨ���3)����J����d�
��$�X�
�7�Հ���Eѕ
d���h�V��Rt8�ࢬC����r�$�QoX�i2!���E���ϩ�#�vW��Jw�1�c����'��Bh����x:o6��u)�t˷v�1L�-ol|�`H=|V}��&�4���S�"�?e:b�N*b�E�[yѦ��pp��O�N�*JS&��\�3�4��̞��s�Z���Z��!v��0}yL�P\1B���H����y1��Pu�;��C�r�<��?9l���O���Yu5=M�^å�a�W�����'����}E�2���L%~����6�����n{�Č�'�cG�f'u��O��i�u�Ȭ�I�H���R@B]a+�Ə��L�:}���կ��#�Hx�<�F�T��0�l˞�h���[f���7���,,����|h¤�� �E0��=l�Q<�k�ZDʨ�YƆ��
��=G'��.6ȝ�'�jjhk�;��:�ck>*��x˻]����x�c�Õ����<q�a*���u�l��9繌!]����!'V�N�`��w��r��� ��83��_�%�݋�L2gv��T�8~r">���3���. f��Y��F�@h��tg?�.Jg�'�oX�&��ɛ��K��Joc���l�Ê���b�#c��:G8	�����m��7k�o�Tw�[�Y�)M�õu:kq� ��[�I0�3�Mq�Ÿ]D��\���b��i��y�^5��� �O|C�%�����;Ge��cC�:��(�D����p��W�廑�߷�;����`�R#��Js>N�h����I����3x*$�c���pt�~�^ �Dq�	Z�5�E~��熠2�5J=\XQS�$��[0�CT