-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S62qGjn5MHK638EK/RBQPDJVFqN+pVpT0XsbHHUuuF6N0nv2/Ph/BX36TfRHL+oY0iVK7nq+3v/1
nDhGL1/WQStvSrX/JW+921XgFnpix/ecEn6mKHpOylvbdUt58Q2EA/RKp/YRv5wzQ8JJpAQIn5h6
yvBQ6iyRYCRRCQ/R6HEMLoRXEaW4zJ4Liv05aRAKJIbWtrJXFeP/JMdGq3xqeFp5cPOlpisJdQ7T
RTmhf/7Dj4sa80vCjwhIbizK8QEVmt1MyG1eot7ktMcze/NSwTsRMpSZdpPmAgQjb9ahI4YylZco
P3TFJfe0jn28EYUljsxNVP6J0jLk73CeaolJiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
8Vt7AXXO9aLJmNg6TfYApH0/WnGUT8SlX5gDQ4wxPpjUZu0I1Hl+h4101C6oD0NFNM2x6Vm1xj7P
QRbdP2K0MB1jjWPOFn0i/IzZSso+fx0KltT9+Vfia+q9a8l7CzbpyrdMW3Pllqjk8LUIaH7X3PUa
WTe/7bYPB9qht85LnL+LBhAy0wBnYI95e0VjVYBYrLxJMh1Pf9lyVL3jhTGY0VNnQXVdGvLIiNDY
flJH/h9U9/6Veb03j1P59cUmf+a6CmzcmXSLueuZi24Q+ayzsuLi07dc2gOrrntzJP53b0kMhVJH
JZ3M8D367EA01YllaNi3529o/+kEBKbdEVT9C7hb/9lAPyxCIeaAwl/xti2l/y88Iu1T9o/TGQA9
J85BM80QLUdORlWNckqNmOJhERg17bqpfhruFTNfgrfUWYaBWT8g2/dbOrQUk6bvZTlRQWRiitrg
XojzJuRK4sYPe7JhHmT3JENeyc3hD9q+dgppJ6pbuNV5iIbof0MxUcVzAR9AC5Usk98NRaMEMlgQ
r3X0E9Kdl7OX5tzwGd4nghNqxzInUQ66aTLKwAVyFwDYgSRUbyQb2o7A9qNVbFYcQ8srL+eiqE7t
gAdZ9AJV+tbevGUxQi8OtLaz0pzLWB9KL6XkXDu9A4qVgVtA7lmOslknykKi5yANAT8QAO2bMZ6a
Z7jdCU3Ke2UqRY5iy76BnptRyrvxAoUQ+6LiPvBcm0gElZhuNz1gAFm95TJ9mO3iu+sVo3DHjl5N
zQxFo0UFgqbvnLVNOC2GReVXEuuKsH+D1m3PlOE0KWO/VOLBKBH4fP8XyZ1O10AuLiebKWoRwRy2
PWzrmdaQw866nQWf2Fn3StEXP21oMvh5PgNh/L4yAA3yS663ug9/OJYNoOaUh4HvZDvbDFLhHnKA
mg1S6lBwQTPx7ktqdaTlxV6eN6+jVdjtQgOk+DcUh/OTc4/zF5kRA2nS1jSzhyq7uvHHbauSxrnn
US/uHqdmVuUuULmpfHbHJVqNKNoi68lgbWPksKEEuLKkZ8d6sJ4vO0mfnCYi4tePJbkqD5b1BalG
SSlwoIHTg18MHSW9Nh/vrlCfx6pAKKVLPHjpttjJMzTydOXtdjMXmKnJX/MOprMnjd8+fb9KqKW1
V+kkKScZLp5+OSSdxXuKaI2t0h0k8hJou1SYPD4MpAX4+0GzXReY0Af5h2fVbZCFhFXHYyhoaznx
fTqaJO+3Ea5fhUZkV1h0D29IqhoJ6BgBra34MgQz7ZQSkclB9/2j+iFGBm94dgoZQKpZ1ypRml1V
56It53nQNDld/N6ozEZrLaK+qVgk0KlKYFFL/UmLg2/7ail2nwMEzx8zbz468iS6VmI1CxsfHedW
D5r2Zj3vqGRtc29dm0bHWBY/FFs7bR1TQGfm367w1v3xieI7dp9ukacQVaQktKPmGfQnal+24V+v
drfVBemTsqrEt1iR9Z3bCWObYc3YaTHsnlz/ghAaB3I+9hBF+v9VfBRnCO0r/Xdhm3jhMRm91kZG
8KFFkrv6vvENOyLrAC0JWICJuRf/qVY9Jj7Ty4SHaaniGbnE6HAqpf9IG2sZURdyS3hfkbqex8tk
68KAA10vvOdTv98O28QxMU6xxxoDQW9Wop3AToy0PQPJBEG2u9p+3Co7ggKCnFeSvrodEURkyXq2
N3P3c1QN2SvibpKqQNaiTEqhs9KXq0evWaejdPysnxhDHbU5GP8bAB7Ozl1oRi1qXHED3ABpYLXe
bTqSN+3F7EOJlIP9rN9XpS3l+gVU4GWREDRAXgHfH2yMjqrctG74AF9CeU91URWJEJL8lMPEXZLW
vnjXoqxlYNwYToxBdQuNJYBf/BCO9/5ILgVoGuPDpVi4XlCf9Dr5oR0VGw0kEb6Z8nageMAvf63m
U5Ybdh/jy4zY4vIwxE0TxLnAJ/BlvhoCGu1qf98vwJHuc96K3bFZhr7dT8Bdkgo7kYH3AaJxhd95
8lunR7KYfQCuPff/IeExVgqonFR5gJdaJXX6IqdMWrhECr/IqPfu0S6CrFUkluGs8nztHJdGblUZ
yDxzi5qpRywSnKawyjmol7R/W0CwH2TFQXi6KNbFVLNeaiezSXeEovd/r1gz841ZfTnxRwpjVJGe
C/PqNIm9ecJ6U5zdNMvfSLjJkflgqyt8/MGsI2H+2LGeFIgyAbNUFn8nZ4ymiyikm9KR+WJrr83D
U39mYLeYseP5/GBPl7S5P5MfWflfEHyLw73o88ihkCGyg2B9MPnP6kufxDTIwKLG4q0Ik1lOhpUE
jNtYPEzhnHeN68UBltRYhyS2Rcons/tOMbVbHRO8L72Eb/GA0dsHHv10IwjG0mIX/qOPK4OYsWVO
3l7a4CY1OIJkP38BgCfL3c7FRJqenyaUdaQd8nMUiZCt4Iq13zq+cYjUV59n4zdJVkBNcgD4gb7y
zRzzBj+VAejFKHiv+YbAozAyefxyUm0ZBvpKXnrHVq5qA3vbIDD71tteJyg7SUeiMKfQUq9bf7ZP
SoE8ji8XZPMXmkzXjoli+XAapeJPH95kf7WzBiFo46pSp25WCcBWaGL586x0ew3AiKgdqsBGKoV0
cyQ0lgkkr7+FdP5D0P7IvS7MLaOzFD4KklAlpEWOysL8Y3J29CEllGiVVPzScd/HiHXWb90twMZC
XiCmt4kzmVz7+cbDDLpLcHAeCzaGSWgL8rb8oEDCdm/0LlpkrlJ83tiUa3xrc6t4EFyGz6qfGqDD
8OdgmpovB6/AICvtv8CtzpoOzBK/rAtU842paBVQIhJS8ehgSXVFeTY9No0TlcAyame1mKGqCIvx
7ZX42TQZTO3iWnP8nZjlk9Qs4DPQWMSCpaghunQJ3zWPqr9wK6xu0uZsIZQpvLMF0AVmnt0LFqbJ
dOJyLziGfmPYdNp4JiR+eVx0MePSMsp0wBuBEEh/PfJfbssUA3pytpUveXjLyeEiefxQDSX6Yz/1
FrPVXFmquWrb1YqDhyKD7cRuIUOIL9aU863r5v2z6QfU8r0D0hrni+EEx2gC+/AmXb3CLblid80i
MPEyxn/W+4icJW0sKQHr7E1cBq6nAGsDWpzLslMQwwQWhuULjZakVwy3SXp0j/XDfoZKaFuZLiWX
GHWpr+wPp44vtfop4xYl/38CSQGKtIVhsUcFGXXtINt2Jv+mKUz4zRnVoo7TwY5rV8+8561EROFR
H1108fGapum10wp2L8CfwKWUXCBdLD2rSzvUwcbsrpEg+xVUin+JbSPoxQajbV8TlytWAIok0A91
bGXJ+YLGzFwb4kJSlfHpzUwWRZKHy4Vq8By3YJQQYFZs/0lt+TqNCabfS1JnBGxbFxKDvfbrtl5e
+VC6YtS/SVHTsLH/8X9dXiHjJSrvVTHy7PrWC50nzw5JaBqL9mTIbimt6ASEL7r6SENfGN5Ga6kY
j0ZhLTTSLQRcZXkrn5H31hPGyrXdEHfP5GVI02d5tctchBx1CPyRTNvYPYoXtTr0rhaCngWnvuGj
0d32dc2x6v/E8op5UmFL9dIpG4FQMqqqNVjL898X4z9gkYIxAiD9AoY2B0Q6BEbhg1XCzIvxzcyu
m98j2lIUee6guZLjK+vsgn65MTCUdWdSNnVxSWC/Gwr+yAcC+XCqlq7MyCKWUuu4d33RFS3h31PS
Uf/Hks9+iaQkkUmCpBym3CS6ojLA9BNzv2k9ibcewLbY9IeaCDpVbmGYk53d12N9Qvo+kG8SbcQ+
yvln6jHExmr3eyfNg9ZkAYq8ELuD4+SNhyxZ6D357G2gIGNwPjCDFTpkhGIii/dAAWw8+w0hL04r
OdA0T4Lo6At8RyoiteWk7yDP+orj5kOXzMpTGFFygPcKvriIeiEKILjyzkFZRxTuPrCB9aMZaaLH
hYKcHNg27tW+6ByQ7eFJpaC1fhiebPt9O6d1XtANF8HQMuA4xOIGq7Os1mu3TrynBhGsggHJlZ4Y
lUiYgpOjBYpRt4dou3vJghme8dK8anWnx56kfaip12/3+Z58kdfSjMz4Cm9Pww16AFvJy5EVA9VV
ERYJGm5Te1VbfS89Yy6V0kiD17tJ3BgMdiY/rD1mxLP69ITqTu0eiDI3NdfX7Nxb/QZDOcMHrELL
pLJUts3OavuMgU03srqqGjmDIL9VB9MjP8+jXxRIdkHMLcoXW2ym0HgWQu0JOjm8xSakzUzW3gpB
Mi4h/oK+oCqhA2qnLyo6m0+AYsnH8TlQEN0TiLL9mB5ZiTh5rvBSakEji3z8Jxe5Ms2xsdXanmw6
X04qLRjyNYaG2Yi8H8Kuasxjn0rrl91AoertokxNo3FbdmEAbBZzLzBMe6V07TntvMHMHc6VuQ6x
OFX+o+9BPPqdjlh+r5dbOwpu73IeUFrTGpYRCFXrdUr+7FqS3OF6c3a9hkjXxdW5+ZFD6KPa+LSq
6klEAg3P3i6Ukhef4fTalwvgyV4c+BA8VPz7J6zb+Ltunu85evnx7Mh/ed6hpBhfsu7EAqUoAPmO
/5anvreqLrdFZIMgji/F57ygzrh9EQnnljXXJZ2DtHKV6ZRk9MB76Iho+c2MIoBvH6s/zJFV24Oo
Vy1EDTGMlacHfDo+dXEZtlnnT5PaoktzKyM2zEehF3NTWZjM14GTbriVNavuqiux5l9Q5GXEZuHU
Zve6nv0s8P2L9nzdWoST3jiYtyGni/wnrDrTJdw9sFDOnNFEqzL62QbY9m4mlCd9WCj4IH39+WWh
3MbWeqwo7puhR9gUL9Y51Rjury8vrkcD7qYNhJJu8ullsPUrflojtdhQhb2q4+7oOS5qYH4bjFcM
VliuwOWkwl4ETftg/uUGU04T8uHA0XNnUY8DnIGUJmVFLlLemHxNsdY0eAqDJez99gVqhadffG3C
ALd+MZBxX3bMSRnhcZeugYhtmqXJIhZnnaRYo2JJE8iaNOiM4HWJTLli+LOFtkLfpqLPWZpUooUH
d47YOsb5VpmY4Mig0odIRiIM5hjgA04+x8Q/BTDY42GMSPfPW/PEvGD3F5s1j7lFddq3mSPhNtUS
rjpfjIukXq0YCBgaxPad2EvflBCe/+sMtTQHfQRM7nz0KjhiMSCgPBcdxEgWSZ3IIYsof5Bpiiho
bkfnnf65WzRZ03lm08or842wiASSK25Z55Wx3ThcJkvV61mBnBKWfjJSoxn+L+oahi6tdGhKOZzK
QGT6yxb5XNOerAG3xwsywgfAkj16O26oiatgbeEofkLBoJifTgDt66w8/yyAZ+FbY9UjQM+Kby8U
71VtfddWfByZPlaGT7XPFv2JsyenNGmfdvS3J34p4Hd3qTNNY9MGOYGr81IDT6eEhWPm76nxr4Kn
R4rhNNUFLZh+Hn6COUykN76N9mdKCx1xlp1d6UwKEwzYDac2yiffVw5rwzygF8NkWId5nRvr7z6J
pkWnZWWtNoAVmEgc5AyNxMJvb0TMPfZGISu+Z6soBR17xnYKlb4oRrtDIdzUD5XC+uff7Rfwffsx
wHwirlZP2dffY0BBJfhRUr6zTfbzJk9PnsAzQHDnDg+MYQPGLXOc0MtMZ7c2VsAxq6+dkFUs2NX7
hgh/jOr1wCOe6n0nE9ctVI6NNDvKyJQePSbK6Tg2dskCsNalJ9w7rsPH2hlCAPv9390L12UJQmkW
t/Pr+3k9C3XgvUWRssDiLEozbId8/PreHopYmEcqwJpleOWEnuWSntFQ5F1Dn5oPsC5AGV8ATFPF
ZzKh8yFiLKGCuoDVliz+QD2aD3ezcse5E450X8l8zGnCI35rcBS8BUx5k0PC8ZNOolZpoALydfxs
UL96tMznnC/1wNkK3PgC+JVTdOXrS3BsLTt4tcs4TP70RzFBz3CLsAYrVSEX+PuYWrTCdrlVzPiq
YlLj5NHHEfm9Q6Y52qEec5a5k3csihfrgkU07VAwNqBZe0cZxOKNhssciTohgu7epORyfF69PmFq
1l5oeIu4lZE6rotYyJu3tFANzwlCwS3a0QgguA8KiLT32/HgrMD84PLJeaYKW583y/rrjXrnL3M+
/ha4Gcb8PowLX206uCQkNm/zTTnoh5MdrkNrtH5UsNHZjS+Z8Whs4ieeZ+EIk2hj4rmNIRvHgHNR
tfG3Q5lITWVY7aTdTr/JUxJ0gXWwUj73D5LZKx9ye0NlaZH4X4hbMMXvNSWyTjL5B1T22GT5cJ/+
sW8s32NvXaX5g3pQZgqPCJ5+BdH6c0KmCulZC5lKcIFQ+aoe5mV04KdGE6xxLBHYrJX5Lu7KPhBC
FvdUQbfcDCVBw2togsjz0DYLoKD5x7nXgz++K4cs1bBWGtkcd76ORv46bE111s52O7KrBHbcmLsI
3jfIQAiy5tAFqneAoR1itYmKA6/5Fj9bvHBmJCMxd4mQ10Nb4E24fplX0qfyHp0SfJp9IQOE7urQ
B7b61dL60uSFtyuvOH9Q1IHwRUff+koR3Eildr9wqt+HPKL+/UY2mgc6O4ous2S3S3po2ikF9vIs
whyWbbTVfHQeEB28uOpDR1SAFZhZCkigIA/hlOM3HhbQAWnKj7vSyseSvIJM8tWnPwoUs4IvYjSN
YEOHTTMieqv5wLkxIQ9e2esCMrX/iFwxwJjIwnhGES7F+vIBpisJMvglscGU4L08zW5dK/F8fFBR
njvRNpghL7/60V1t0CNlZvdNJ94UyVy1cl1kDgTCPkMpwoAHjn2Fdi7hlTmg9HiJPEdN75c4TIQf
algHkaMvxozIuf/pAJR+jSxpobai9UPwZOnN43CZV4flF8u12dAPGxo11KYNvovuGdDbFopsWYER
oJqEHBmnstfpuOFN/KjTtmd0+LjY9W5JaFlkVXmL+bMK8lopugS4ILunZN32W9PUVASKmvuf0agZ
XwayS2trcRvpx43wgLJXiI7WE+QKmqhzs6UkueFyAac1cClo3MN2nmhmah+fHb64dyWyyJ+LhHgd
ADGMKeX1GC180MqYYd74wf3/lhKfD1A8fxV+KeAlZqBwLdwxKIN93c9JvFy4wB3q7xf9FlkDi0pX
4mdmcJhT05POuTzpweKMX0tu9vIcpZLALnK5WtRISWDEp2hnF1AITYVQ7fgVawK7rd2Bdi9GdDOL
quzPsM57IDf7+aBUHeEzXLpYewKQDM4UuokaSd3RfGtW3/YN0sZnlXlJutkrgkE3+HPU377oDb5W
mttiGAZKnSBjI/zEPxtjSCgQGc800GjXzyNzvGLPuqyC6Nfl9siLeGA48FbDBxZ8AEQNfgAIxCaD
TwAOo7WWom1lZd2iGrAXtTRAcdP+gFIGlMPCHs6TvYiOpKWtbq6SIa7h4pcbLMv4nvNfWx6zYBeP
PKdXVUIl2I/NS9RlBRlgh0U8Y1y79FNK38NLBFX5VHF1l6keMkc9uJkDaUTsBzcETRDG4nzed1q9
JdL32JFh+6tF82nUEW9nxApWZK4IEHSWTOBrrPDE20MmFF7qm496bxniWAxUCMtDt2WYk+y2W6gd
YvPzpf2PcirNn4qwPZRtZ0+BG6I6Mptr2rKWyyUUzRJXAX/e2n36YZ6zPZqnv9xot+Ch/dD4opEy
y09EbWr2nWZppj/3o5qZ9O/1ZpnhTrmQmbFB/3VdTc3QkaOYAnVJH4wMUFNfPdcqYdmAZB/UkzTG
ZO6MuPzvucvcOXQu+Inr78CFeo4nNtIJsXMei0OfpiLwc0GYeTiLmbLSCF/2v5cbvGLAJIoSygxB
HzBiXLkY1TRZniA8QQhkjAJqRioC7oY0uMnbQEn7B/BUJkWNLXK1bJqMRtRzUjDC1By/k6iIQWk4
4qbtREB9FwAL3XpgZIuSH1LFASdj67VMD8wliW5Pyh7/ME+BGok9EZi8LvDMv8pX494tGLLJyDb5
YEMal0/z+ODRZKVeEtoQ3XaEzAYq7PwvsBJGQxEv6yqeOJ+NiQOHxoCRrVsMeIn6pMSPFHqgSBWh
/GoxpKgkncAgemSunRVZZivTO16Uecx1jZ1H59b0m+zI5m7PIUAa0DzZWQ3UTpNksjgdQlqb28Vj
5sDkt5EaMAxUH+HViGD7G4rg0IlQBoqJSpTt6EY4C5Zv7X6QHx4OELyrw6e9eFDmyhNczRSbKaeB
PanlZ9mZNKECAy0iXjVJuRHzqqeEH1zI4QrwnUPfV4Wt2nuoDJP87Sk8lT25vgzQqXX0GWL2kIsE
ptYI/iLc3wqRcgH5jukG+Itg8LxcpfhyI0qhRdvRIjFPrL+g4341g4qmKayy5EKTHaftPCR9c0UG
VboeMGaZiFfslIWs8oN6yXic/oRBpZBxuVx/FeCj62D/FMErQFrB9MuGcoGQ4lNNXcYbqYy7E2/v
tldEIzgShkB/RCIPku6wg6O+m9Y90xXCGdHIlmbW07WXWUFNXlVu8omae303FEV4YihvCjVgBq+k
yWekwX060BuEiVE8C4GaKUCDtMhOcQx48WWIu5BcEgh0Lumq7/wwQXvBPDtqOP1N98K6vrOVMjr9
S+oeQEPo2mgXrz3aQQkIz5FYPvOg2r5sNk6ZJbT7hP03sGEw915R5FL/5EOzN0S5zP5e5F0wUWNG
bCiSqro4RSFNoMxJcsvYZjeij0VJAETQ6IQ+9gUXWaS0gwLB9XQMJ2bNhbOTLioJi2wMrj0BYIC1
ZddsvhnH+QsQV0oHvxsuKyJn/EDE5dnvOrnQN1b0rVxzIJ5C3cL1mSpoIn+1/6jrPKj7VI38LK0q
b3YR2y+WqUyP7RX18n/ogjtWrzw4vocfiiSbwgqcxLwT8HgVQ/O6LOkS0AXtgcYin9ownmLb0uXA
vODEUfQgmFQ8ZuX4cxKNH9z3MBd8JaqAKGMd94rijpkz56/J9B6qW1+tPeOhpm7dYM4/vpyZn4f+
Q3wpJErFPFRVc9A1plGKxufWihd/wdLx3tA/lBsJ64DPGXnEC69ZAgBrR5NRxaA9x++PuGSZt47a
IbWUon7t3NPQDloG18wcH6jnwiX0g/+c05IxC6XjNOkFdRKktzmmQY6kAA4y7qx1cKZBvepQDEo/
DA+4QUJ5xbaBImyi7Xj5tQl5WAPMMqQf/ha6D8TU/W1s5DV/FKxtu6zqA0AjCMmukm9TLbRHiepF
BFP2SuRaGCTOmoWXQX6IEmKQYLlq5nrPp6cigV8KQWNSvhAZT4vx1bkQf75XmvsX3H3Ix+zYgqW6
UjGkQQiozO0w0p7bDc/TslPLzYhKz9Ll1Xm81NMnFWg9L/DfB90Xyo144qmueTVvvfE8rXXkygKv
CtPvVY+/ycvGfgkzuoz14SYmTq0/cmkmHXldv7LZfmbs2fyBptisEQ14AhELMhaKoVug1vbzWngd
0ec93dlaUINEg+pAGp+9bR6DRChKc5DNMhjOqa8nmlFDb/CQVrwdn5Sv4jHgbvKsb2aD+7BGfU9H
bfV6vDKVThI10Kvb+IUVM2cGinCw69acQX+WU/CmgzWg4yVi+vDGVz3JWGe2ZOApCgo3iJZBRPvv
968HwQFxEzOhTPFBZYK2fxpt5oyD+u9UNN5fU1llrbqlZIx6YJ5H7k89INGoyvDTIBjYA2O5gC3f
o6142RsjVott+rJwOaSlBVF51Y7EnrNaGuUFzwMXOlkLXzXDTyhWjW4jgXgysYpunnaM1Mg4vcs6
uNZel/bUdH1WfvfJH5B+CcGWP6D5E3bckXBUqHa5R+EP5JcDVVMP0gtQApkVhgyd+uaSGSUW+m/5
0ST5BTTEPfuTBGlInsSvL5z2pdOv9tseQ6tW9SdnJF5NJgl/hMxyK9KMVmaXcNVOEN/beiVT86Nb
xVnj53FkPG27COak3mD4LuTnrYBc1Z7D8abwRiwFP7VZpTX80ezV9JpofvYTByR3dZVIOi7FPdks
RmeCqouahVwGLcPJekn10C8JjeJv3i9mzbAuazQ/mP4HAPmYL2noAxVCIUo/uldw7s/s4uwM4BX/
Z/5FqHYzx20aOiOKtSnGUK90rRbYUAf7O7R9H1LqQqw22MkdfAxqaSNccxVZGsSLoAiOFncMWNBA
nssZ0OXDyTzBXJ4YV89fddqa2vicVQxG+NGx5cFlKE5bvOjyBSJTLJvMFDEj6OuYAJTlmpqHXLGF
WesF0uVwwY+KbDT5u8sbgjk/FP/0OYJtRRHyvnhkFBWPJeZmMxqO6SnaE07XG4g2UqjZQ8e6TuiK
s2SmgE04RKWfWakhGtL3VMX3Jg33S0M69+DIvb0xvmBwsMPs3nGSfZMoFlcYqvcoDcOfH0mY94f7
wbcpPplLy1tu3+ykheXeM+sum6DcJC/Eniy1sr4LtiUBOChOBI9McCzkdyECTBEBgkt68TPCWpHF
/xN7JalUPoLfmRFz2Rt0OT7fCJpHou5/262dNshf8k3pAZYHxWclzuiuyeWdRKSCJ3+DRHCTpFEu
JLyztA1CmlT7vqnWq19BUrxNaW2a9ObM6tvpOuM0OCa7b1u7aurKZz9FgXpV1OK8IyqPoJLSCN1U
lSAWpSjAwteDCFxxWi+vhwX/dOP+ulQSjoiIUhpH6a+POMHpHA0pzUF298LlpJsOKOt06z5KkOIP
CNYF/tO2yT4CshsRDwaMakEjQDi5joEimrynar55M2ebTlyBMJS6zBrxHJ0eRM1VBY5pn4Hua7RK
7NvBnRzk8CBrOMrvt2NoaGvu1cxPPskuWyS0/qBpnDskrU5dmhw4MmzWboehnLYO+fmieDMJ+CPe
MEh5BfH/SAn07/cqfh929IGZgVQevlUOsBiq9zAxOtvcia7izA9hNkxU+QtWJMB3D/InEu+CsW3s
WpgKp61qgbMty5m5//9jjJo91bwKoZ0U+hJdwRXaSsIoTnVDuGnmusCejwCXtun2wzn8r/xvZA2E
MlXaEGcMo9WPs3dMLBAOseNpQ0e+jgQ2iXqPMQs37hwxeT1vxwJuuTfFfGUKSddJALS4pFUsI/z7
ZqDxIg8K3PiBW4q02lzv7Xf25q6oeUNNoEs/2H7QqVk1upKud39eYJ0HGsD29dH5MCXRaDrxe6Lv
HeEGqYOKHN5agBwtMo1ORHNWC189eyuUCarWNs2Kc54FHnal21wDSJJeQ4d/XCvoptPpDmZhUXhw
lFnJyP5E46ZlJ0PcJvf14C9DnNrivHasacImg/yN7Bj8IlSOVJxiaOo0vFvUH1sD9oqG97bf4u5f
Q0UR+ptloQlXHp/0wXLTs/5kqLFO2jTcoMiUx3agmBrmbtBFmtgmw6VQ45GgyAxVtAgVib/29B7e
gatNVF4kaEHnr93VekZjZko00gjbUBgZXQ/yhtDpwZl6UY54rKOuAJzuusPrMvkSjccPlQDn9Lvi
SAjj4Q55dfPOu6qONMpvAGy4lT09rpR2Txi3ZTwb2WlVPwWADEJv759GMnqqa2XCTVEwUQo7eguS
EKm3MpA7LyrniqgBScGV8Mx8QpwwREyoAEP58tDD5aQydkcIrnGN08dS0P8U0QSEST5yoQtJbC0O
iv/cR0O/fOwbCs/evEqHFZ2fe8eJkxuR8XlEfAXfgaBi/1eURFnF86fmcfvk8A40/Ya7uN6EJ5HK
z66DsqsqhERgQUjMrJGw/941K7sELBrnjTx5yYY+z8yAVKXnp/uJP+ytWxYkvaznY+AFI7QcszUP
zkoeTYKiig/AOKUhZkzRGXDxspPuFjazU2t+WJiNWpDWC+KrG2vReDlLb1keGRmCP+al3WU8hFFP
96EyrXOmVB74k26iDmY1zY34dRMhLIJz4QbbIdvNZ3qBoIOyaLiX2JPT9st0BO72oM+e7w7V/sp1
1ttremX2jLivvxDaNftHQfAKpaBtFd/9JJBFLwiwpUV2mjON/h2sRt5wOXueYyuGi9rAmCEVejnz
14J/s/WXKfaN27GVBVQLZopzd4ahcx0FgA1uTrryfVi7ax9mtqGjTp8vouN7wLswvu9nzF9HacBf
FEpFA5PNGRmpWaqX68kBZL5F9Q2kF28Fszm/nuJIMZGtoPQhm4tyooC/Uqh8KAzqNsHPAFj3y3eK
G61NE7fsomSIeqFqt+WVDPgNtEE76Q/vlfK84U0A6e3byIxvkaivKc927FhYZoHphfdERaUPV4U/
c87I1JufGUxBAkfbFO8dfXIAtF4tVfQpZM7txxxqfx40sMNOYW0DIQavMNIQuiT68DptKPxQ1P0A
cuvYI+Of9gdgw+XU7gTMRcrcRWtLtQ8lrWr2cg74QpHGpZ8nlsJOyVgACafFVdD3Ot12PLTzKs1Q
Q+hl6Uta7A0ifLXFRjMLKDQLbODAY886DJNKxOcbJZ9LpRVvp8BQrtFOJhZCTKlzHZjVKUydKWsR
ecpmXzzSG9u1dXJjOdzMNsUkLZVNXsmQkN+nznmtjR86GVhgq37uGiNC1bhjisF34yzNrIkExGhI
99p4CWlPFt7ohe9nXWvazmLMyhjry9kcRQr1woeXKBGqoth9orRPi0hg5oZ3tsgqzYrTAhKBMj+X
d2of3BTqRx9HmH/F4cgT/7Sz6woWLWY1XN8ROTnOrLzwkAwcQwJMHDETBCALNp3dT4gVXEos6j17
rKYYD6XPAkX0V1B4+0gnfM7IiwOZhdmZiZ7l53vUdlVSJa6RHZcf9iI3kTWOrMs+yoW52sG5/JSY
+QzTnbdsA6Y2La625vHQerxXezDYNauSVajhdwhFuTXCeEzRQkF6BRmb5VDDGzKYve44MA6qwYvj
iDJVdlRy+U/l5tbpMC8yqptQVMMRmzP0X9KkuDIB33OMdQw8ZuRXF9NagTOIxOCuHAThK/33QptA
y5Ii5BA6C+io3tjQiyIEPmi9BrEfTvrcgda5tLcLGWQHHGtmFc+KB5E8BAUEcvdH61ujlPefysX9
tswvSSt2UzkDJuXlK8C03ZOhsDL5oA2HoYlEZ7H7a0qXXq+9s7insaY4RuGdpViQEj5gucQcaDO5
rOPdpBYflXa+IsjKHWfsu4+YPaUQIbBTcC+xL4f+FaDtHC5KUBqTgXnZ1xzqLy4tzreK59Sevltr
IXrJpdsOY1ng8ANUU/DKzl94mNkfSOtPJFXt0VCAYroE3HCkiOxZ+p+ZRhPp3TnAHBgGfTqmTGlP
PHUq/H6MgQrjugVfV0/zNozaImx4vut4UQHPIW63O8patgrWw3qEi/OOjFMzEGuz3r0hV1t5Z+pd
ILW4zLBaRxJ07++k69BfHZJpEI1J8vh9wHTz0NWDGEO6i+C02dJTxi+/pQjQfMeh1vQtSac2UlgP
ma8IpJoni0VOP6jB9YLytKvkILsJOlHXf/iBtm0wFGvMvPw5ci5tST8xyLF1VrENJa1v68YtIQgA
saJl6O3X3V7IHM6NjBdW0yonQs0O5S21ryo+dyQlu8wzPgmWSyu/FWFqPWeZ4dWj/Lt9bnQCokW3
Fk2Uz1E8q/GftYxkCBIh471iM5dTIjtDbGCHKon4Un34JDDockjnC6Ph5IOXeAWTyV6yLOMWfoAg
eJmITmgHr+ZOBQvAr/zGQbbCQTEfP8uoVsYrxMrW+45gFcjozJooMdvhIT+ThvqsjFuvgRCxDqCi
o57BuCdgdYS8lOz5E4vJ8hvlGhbyhO5Zw/paVAI2m8b1xW5wlkdDgcQ6v8bkh2Lx4qGvPkC+7esT
uihy9jAznnCD7qP/iboAhQg3Ym8dIrKeqyH9+ShYTYX0m89z1NcMzlFMGvXYuc/07z9v4XZiHTGZ
FBQPMW9LGr6Pm/5JNmUO8w4LEs3pFVnxwrJQXev/BJTYrMMBASyaxnkxjhEWEEt88UO8t1EjFwku
wKSGgEgk0zudiiHnGYN/lcZ8HVNH1WFLXXEhzEnr7RrnLnsXot98onRCZPO51J/5ygJB+/pZwGnT
fJ4uvfpeqUzv5mzpFHSwBCo4F72kY6lAOjfuh02a90P1LmTyyDZTi9kPCPqznpkEQIK9i1cPi3iP
YMM7z77IBllD/tw0qG9A6nJkjJRycGlcPW2QQsFavi6pZTBBwAvHYbrNaovpmljTi6fW+thZ2j9z
TcxGf/2/onycJwVGykFrTtD+PRV/u1rmZzThdMN7jNV2KZpgE9e/1ENBd7x750Is9GcTLEfDs4GO
+LG/Sf6QKv9qeDDBlie2dNB32OBu4O70K8DEzqk9sPpTY+RIWOEQZr+u2HYzdssmqO09hOlH0nz8
JoogouP/wTZOi2AIsYXWfk38GeC/MF5GZd/MzDtlTvO0sQdA2iMDVAg8A/Qbn1K5vK/UXzw7ZVUF
1aPUiHPfNi3T3UGPL7Rruz/fa/dA/9QKKAG+ot/iQc1QDlXtgZWohyXRxLcf7RiBdBcPrgZ36IVh
WLomgNzEfUeZsYak7AzANNVE35xABcDmzaJ2DMiMskKenNzb+6sMNFTgrLEBSg4tntPo0xJ3y9nv
LkpKfwi9n15Us89Po9ZqNTXd8Je4yFenveZoIsc6haIQgfuzJJxLSSvVgtf2TXLKbFo2+ZUTRKm0
i+zjvG1aDcAqHJMM9l8icHNXU6whfFwEkBfnFUpGZraEolo5xVJQYHayFybpkyOzMiwGt6yqqWAh
uQGMo2rhaVzbIe10sZuMum6wA+ATDHPYyOGUMi/kB7SeklKP2kEMqpvUrNLtdsRYpANeCtHj2DgA
mq7Kg/pDzsaijLvGOYwhXdrdBhadoiZeq94HQATgqTaxiUKO/NdTi+zJnBZBpTT3OvN8n0SeG538
5k9Is8JOnSe71asNtmd99CPyQoMstXgCzOnho9L7EkwfgntGzALNdztD56Hf4ujTT16hyL+5AGHh
soPw4sJJ2urywyeFagR4S3nNXHINPUcLcal9gnzpDr2L0D7iMFJZxCx71pDBu8498syDs5c5bEXI
CfdqHnpcYu5UvmpyQfvytYx5RhnEU+VCFRSryGPbyEv6Rk7sLqGTzJv4+cbvCq11pOUuwocfGNUj
ehNxAyGUWcsg7unRxxrvEMeEPRgmjOv/6mafi6RLHIymNyl7H/8iTdIov69maJ4PCNyv/wAaCMI4
zm/KdHZNMc2Ss58BSvuWFJkuB+fmwHtgbujpHsL0Qd7Liwbjll79gnRLl3Rd1hEhGmRzGSADObdP
wiO8K9LSt7bYvQBsOsUg5pdnmWibCxy+eXty/7Pl7XEpuTblkh84Yl1VgdHz7X5TVWEehoc7+9yr
PxLmgowHh1BB019QXFqEJs8Av7PC1fygvjezsTIYZ/6YdzPWQL2FgZJxF1GT85b4eSzJTpzGFM/r
GSANCgLVIJ71INWicWahjLOtG4LVJUZbyrHdnAY94DMTDkpKCUonJNHfxfX0NOmA6ofTuRYkWc0x
FxszdLZTeM+5weJvRuBlEPeUuUaYTfa9Sj80MdKXo9wUh3YXQ2Raq2CwsWRh5+0n+IHLhkFkVFiL
wjgMGK3aOD/GQBxc9pdIuAxtLDqH0pUmFapSHk4Zt+Bph75OsE4y013llmDHcLr2exr/GbdDASf5
LapaMYtQT9CxvmN1Dxjz6RJYci2RWM15/CJN4kTWmlFVZG58kBbIMmtYykfK43NMQIUsyDFE8D19
NvIyAjjkkCGTXi34QvRU/9b6/rgE4Ewiu6xBiYaZm4YZyao4Gbq81D9DNEkYLk/lDCXmBkapBrJl
a9I/wjihCFR11SBF5bgzgNKQriGc9q9fw72h1AswDLqgmX51NQOA3M+KkYjM+L49lkW1l14Q6jFk
yMcXo/pabVng+QT2qowffWo/QQ1XQVoAhXib4BgeQXmfjSUp68pTvkOgXSUrDoayD+a6yq4H0p5r
TtP2FZN+L64+G8AlAC2PxYpc0DuUB5dLOHrOAEPA0qJHi93ZpjzOfVa2bPPSdb5lWd6PORRhmppE
cwSxzcHn7uHxUjXjmXfkSgnVXtXliYbqrhVdgjY97BLtKmN8Qa63c+Zt/icfwRiWLr8x6tpas1Rj
En0GC6kvLicM6SgDrYnv/1hwKkYroWKLG+unH07DjawEaalMswNSF5ix18pfqKO3Dhls0eLSwhrJ
G9mPE3IxqrMu/N3LdmSS8uoEZvHD0KYDY3k3XFAkupUh+emrA1iNHCA5p3va4O7JFOboVNhrCvsV
EZeTAAsoLXTo6bO8xrl1e+ERQwXvJKDj0qSSd6RW0EF7/CkdnduL8XqIhyFhVb6um9mkWkXr2e7Z
Ccn9qRN3hGuvQNnQ5k6QTL3rDc8jEnRdS6etHO4cAdHvt9fOIfip/ZXGXaoCnDljt2LQJUE413Ul
/tHBb9D0Q/a6b7MFRoUKA/7LzbWCXugrZGInLSdZLulSu5E75drbzeahR7ZYYA3sEjr+rgQKo+Z9
YjRqCAho90LBuecP75hbmjALYTxxH5Ad8iSTqkred6xw/prviPdFblpUIMJo+ZVio6SOAjMlWtoS
X6L2VtQR0zAXZmxY7RfIPMd5fb7xTxz1EkGHCou11vjbn8umjxCWmp99QvEfZmmAOIuAHW7E89eM
cV5umbnZkEJKAEqm5yTqLOkmVkSyOX5dpmMy4YYsYOQsa7jNEKfBckvaYIiBZS8gXofDWc7BgfuT
kkDBoryI7+K7grTPZpnVN7Ddv/TT4FF2EIVFxyTHeVZ5acSh5LBnhlp+UrZYMlD/bcYhjXy/TcIw
hCLkeaBH7HyKXs2LeNGO/Y+/Z32x8hl+URvMZWeB2ZZsSiQI55t08cxEvg8yr8SOT3ZZTr43UnaX
6Ebk5AcRUQ/ywfqg0Xz2bq3zFe8GklOutoTdiSPDsLiRAvW2eMeSWtJnAOJ48yMMsi3TCuKV02yF
EeehpaXfHBurxVa2Ky4FFcC+uV48oNE1uzTgMbeqNZ7u5UVYFsAT3GHsW5zdyC8m2OdHr/ACzUKg
LGS1QGkYdEJ2hJjZ8u437wOi+5we4p/Dvi29j3GM5SZehbFRDUUIWZ03wDPojhPKUzHiXw5QmTZC
02hSQxXJe214CsP/gJ52Gt/vZaPkj83avLQuxdviiy6Rsax+9WoIu/k+RMP16tJhl2bnVOfoECvm
uA3nEcj2K0P7XXg0pkvUVUZ/viz6VLSUEfXXgyJUm9TYVSIJRUwuJjEF4Q0ys5WafwCcWl/cg18m
HwMaoRmYi2pXCGAc+gRR9MykSWsSb6T9U14Pq431dR7LJURZ9cd2OAXzMCgIS9/FaD08Yy25hwke
r3WO2RuyP2J8t+PN5ppmh7R5MQSAz2I7D/zn5oOaTlk1p72hl/tP2pkeavzspSU9QG3e9CUhPFD0
6CICKNYoeD1MTBw+1cd5nSQXmJnmXNgdXB7rHvvzCUQEkULWJCF4uALbVIiIRfZzmDo2w2QTo4N+
1FAiDBqP0uJE/E6QfXQvKcOEkpS0GWDXMOAOP4hv8TfS5omYCr8YP3Z/E+p3x+JJI/HjSqt2+tn2
YSmvYGt4oDLIfKdwzSbURGmtnCQlOmvqWMQ/raIzSjusBYOYOtsnYTBYz1WdyQD0Zt/epie3y6t9
5nNYdSKLgsfreVbXPmbARvf99N3nVtiXpL8Q5JZPHPEgIVv7nHmntleFmX5l75uOlXQNIx8+0jtD
TSYBeFWbjT11VbsfT/Oa5Tqeq8BH/fDHeybFr86OZC2SeGGxzmht013oAWONgsXZ9sx0beO+ucvi
gYL2ZTVVqrPN8HNHmC6w+8THKTpzpd469k0zXNS0yFAQDmD4wTy/6Mja4x9+WCXeQtXH2buV+X3S
ecUTqjfdro0Wax9mZWuGWzzwy3O8RsuxhiX3zM9uBAOQ9JT7XZM2BqxGgWl0fde96fI74wdMDjPi
TnXe6mK7xPsr3LkE8kuFg08GoK3zXriDsXiY+2GbgnbBf8ZX+S0GgGsiDX5Qy7xQdiVD8Hcgs+jv
f0ykPatNazahbIivjUma
`protect end_protected
