��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	B�1Ƥ�.��ʱT;�HM���������B)E�3\a;t+�lr�uY�H�J�,<laL2/���_أ�t�%���d��bݓ�Z\i[�<{�eҔ4u�m�̮�Nj�Ü�4����4�&}��BXk��_q�QL$m}&�S�s��1MX�eGr4�1�{Ꮙ38�/Dl��Sr�����7��k�[�"�;;NX�:��gL:�p��E�>���� �P��iT��`�{=��/�ۇ�t��w�?�N�.�/i���E�7�Y���b�&֤T|w �0�B��6F�?�L�V��W��x�@���"�vT�P�*�1���I�SVung��2<TS*A��
�m�I��j]�R<	�N�Xk��L��	3����f�>.��ZĨ՜����~7R��;@�"`�l��}�Ҧm-ޙ��d����n�Y����F����?6nhԞ��;�m�Z�]B��z>N����5���Q��� ��2A[8��4�J�����H�C��E�-��7	��1�rqcI9�����2�CDs��s��*��d
�m�E�yw��]x�{[�HGB�A̍qy���kf�<ȟ�wh��̻y�HԾ��s/��O,�_}Mv�8,ӱ-�SZH��lU7N9����x�� ���,�8����i�0������fF��T���NZ;��V婘�pa��h�5��
��t푅=��B�2�l����ݛ�����ND�v8�bѺ/�*x�ʡA����i!O��v�X�7�����:òr�GQ 5���\�7�q�]x�����4���o�h�
�I����g��K=I����ܫ{�#Mo荡*3����#��r[�=��5�3!��i�j�&(	y�V��`m���Iʅ��A�#����`��v9A���W%�]�ځGhI��<<��şf((	�#n����7lT]h�/�Б_k�Մaq,?�|���j�TE�4l����E�:��5�j��Û!Y�p���Y��8P���֐';R���0� }=���"y���� 8���� ��f�q^sIA°vA���c��T {+u���{����(�{���Q���
�p�ǝÈ�n~��L#�֥	rKV��\se��be���3tl�V25@�_�붵[��LM6� ��=�J��OY�,�;�ה*���icHI��Ar�E�i���FO4��ᅑ˜Y������i����A� V��"{�r�.hL����I��_S`���IB?�|F��~r��c��Ǜ��~��G������D�{7~�-"���"�|�([]��,1���z�:���Pd�p2��wI���|�с~</�o^�bI#�{�a���]� Hh��@��������s�E���X#j�=�iυy��V
��rv�Ur( ǈK-a���sk������}�V�]��i��uo_R8F��LŌ���WF�,�h0�sH�����������؄�m���������X�y��O%��9PV2lV]ΟK�JCi�zf��]G<L�I�Js��ы{� ?�J����^9<}x����u����
��ʩ�`���P��p��A�����#��[SB�>�0z$i�X؍^,�����S�fp;�d�+�T��z\.硓I'�|6�����DJ� �O��#C�'�Q�k�� F��6�=������N�	T�ѷ��� �����&�bi�iIY�=B�2��l���M���Y� ^+w#B�lU�䦖����{ p:]�9��n�s^\H5�	������"���EJ�~�K��Dw�p\��v�q�:���~'�x���p���>�Bts<�*eO����O0Hx�Ξ\�'�a� ��TIq�|#k�-�U�c�7I�����z�e�r������TwX���_�YP��Ս� G@n᝞�tw�oZC)vCL_��Qx�WU��`��e��{^�����Ť��J�L�dkS�~ӝ� v��8��:>ҷ���lP,��``~��fQdy��uM<�W�>��!�~�ʋ$�W��%XgS hRC\�r�	JM#RD4��J�x���m�5���%o��������$��\Aǧ�}�!�;�������rj�=rӒ~�B ��]?����n��}�z�E�l��͞T�H�;8��nfE�3��W�n%��w�/P5���G>6Y�p�<Q��&��%+(�)��p�#j��]9���#5�C,b��8��dc�B�>��|bt81���}�gIl.�W�4�w Hɀ��Q)��Zf،�Dr�H�?KQѶ7L�{��\�`������v�J�[���}�pGx��a��*���CQVxO!ض����M��;7�]53�K�_h˺���g���o�[�� ,���Vn�ʁbвѳ�T��P�I��j#tj�����̂7���i��~��l��
�C�a�����p"��暐(6��ۍE����z�d�W���A���K����.˗�oZ�B��Ŏ��Ǯ�i��&��2nK�O�7^�'n�ob��gs�$�,_������Z.�"��f.f\~��Z�C�p,a�N�H��f���4lNnv(�a�����>}k�V:�#*Þc#�o��[��w�`���߫�Y�KTM� ��?d]Ҍ�(3|+����
���K�[���3�i�ﱙ��E7�_�E�~rpQF�������O_
����ӍC���z�Ri��]��R�}ջ_![��杴�$��J���A�9���x�d&r�8�e��nx�c6S�(�� -���LO�V�M��m�x�?�z�z��ɰOj��0Ϋ�_�	v���.�,�-�͈^��i�� �Dݯ�q�fc$���(V�i����[5�����z^�fO����1���,h�Z�CM�����L���>k��jE5�(ƒ�uo�1�*�6��X����ܿa�gjTF�wN���i�~'U�^�O���*�x'�[E�=R�/
�x��Pf�S�[�+{�k�29��	��!�#�����o `1
I��J�DZ��|~����:r���Y��/p�l����t�n�Np�-⦳M`�@YRf�����y�������QG�JR���di �?s������R�0�^�Ok�-&��:��_�*���e��7Ү�+׏J����J������XZ	?}iO1mɢxT0���{�v,6VB�g�j!��7B����N����� JD�f��$؀F2ܢ��<���AWѷM$�!�Dp	����%�0KV���ZÌ�Neb��5��@���-��irQ*�@�x�/�X�R�vz'�yY$l*�e����֎٣C���6�DA�.�X\Ҩ����,�׈���7�Ů0��&�[Y;ڤ�	�
'���VB��<�C�6r�{5c�}eZ�$)�Y@��n����qe�����&%l�A) ��X9h�]���H�6^L�Ǧc�t�V�TL۴In�}�A�D4�J`|;�`��k�X��O5��X#�������φ}>%�-�M�R�4����T4
�H�"�PI�UE2�{<����K�x�W:�������sU\���<���]f*�j�'��ׯ��֯K����@�F��e�c�-r�]:C��ђw�ҁ	mxzp��iF�5]+��,g�]�d�S�q��i�%�b��������`�I�#�9����2��8�t��}�o\C6hL� ==h|����;���U���G�[ܽ���#����c�i����=�[B<�4#;��2i�ф%О�l|���)�H�Z�2��g���RZf�N���Y�M��//�I{�����uѾW�׺��ʆ5�9���U𴎃�#k�y��t�$�Jd�Z��ѹ�̥KQm�u�ĉ�׹/*Q�t\_	i��+E��*�τ��e�4h�^�鋵���7��W���6�.��ŭ�1~ctW��2稍���9��d5s���F�q!݆�����?��]��%��ܭ�H�R�L�9:�3Q�D����A�Մ ���U�~�brdR#��i�l"�U"<q �`��KZ$]oӏ������{���%�!�S��cH9�>3%��j���J)��^"ހs/�����`��=l�-�<U$���oT�Œ Z�>E��h��Yu�|gO ��E$#����_D�?�~����
ϧ�Qztl��3�e�C�@���!��^� e��qF��5F6*,���\�5AU<>�i�m��vH� suU^�a�J�x��1��K{}��(�֍�޲J|@�� �4z���b�qF?e��"��!�*�0_�/�n�Έ{�a8��6�Ό�s�0s3��׀b��.�g�%Yg]�'���-YHo�4��YL�ve����r9�hm�EChh���c 9��ˑ�Jo����M���oMJ�T^�u��h�% �����T�	e#�i���{�w�4�r��9����X+����PA�<mQ]}byH�$>��;~�XoV���Ѱ��~	�Ȝ�w��M�V*��)����ۤ��m��6@���� J�N�!�I޻`���l6*���^K%Yo�)n�V"(t+'ً٫�`�
.�}�@���4���B{r�H��s�moث�D����!�.�Ȥ����e���S��Ӛ;�xTn/����'��׋<��g]"ʢ���A��[-�jP�줗��9k�u5��0��t����	L�@D�	_u���а8��Q�47s�7��7��{b�S![�^��(�E.b� $C��:���h��hk���R7t7ކ���yr��9 <L}zI�A� ��N�#\�]��'�k�ex�%0���j�^�z����0�/�z4k��ѪUа�==��m9:�_��ګ��ω�1���Q�W
�������kVu8"����Z폟g�H��,���2�0���:b��oؒ�tx�V�E/1���/��1��R��o�<��q�	^HG";qW��d�,W�<��׮����?�Q����.������c�g��r��z�ҍ�^���	��T��*�"�U�o�Cl����ʗ�-<�i=�������'��s������:]�Y�n7�|����*�9���5MUhP?t��y!`n}���ij�/�A�"�?v�F�?�j�!������f��S�_��ˉ��c���$c̈�a��ݢ�^Q�~P�F9�zB7ߜ�O�9a^��7���ey�
��_ �5y[ၧ���sq8��Yg
��w����)E�uv�2c��d����h6E��#�1/�m7��_Ee�d~L��=��~g {������*�PI	aP_��.��=Sy��ȩ$�	!Y?�8�����G���v��D::X��J�j:���n��k��tQ�����~I���n�����Qg��*���@wZz?�/ћ��rP���U�s����)܀�e��q��f��n�O��lq-�+(�	;�T<�I%ڀ8� �2�ú�t�L�R�7tfMX����\�	0^Aך+��B��Än1�Ct�ؒw<�>#E���8�D��̖�3�9���E8ۤ��V����d͂b[��m�S	��yX��̤���Kd�ΰyFY%X�/l���*z˿m0� �������o9�597���ih*���d�Bc]@�MIz���o=W�^
�ע�g�'E�?��`$UGC��k����o�h/(��z֦+�2�V>����a-m��?�����ڇa�P�*�	s)V���L�$���ܷ�^��jzh���dw*+�&�Vz>�H)vJ>:����H�gh��?���]u�4{�I��`�z#����A gp�JOf9�uD�zw<�MP��M~�"]��r�6Ey���>1��M���$?_�F SI�h�y��/�f}�֧�7FW���3���g=ڏ_P����	TS8��$.�^~��F���I��<�4Z���/;u�f��O�T�tK_�L�l|ʩ��B?�l���6����S2�e0����F�b�l�[Ȩљ��Q|_�2b�;��s��l�C�a�cZ#/FJ��!K;='��)�.�����K'L�e�xL$sí�'w����
�#��%1�	:a  ��1����T��5F�/g$|��{.������G�.>?�?o�j~�XN�17�]�d�쑅�|> E��̸�MF1W[ǻ�%�cr�qB���VE�� �tj�W�~���%���w��`�5l}(��#�sE_b�kЗp�	]�r��Ms�6��#\�2��4H��'�$�|8�X/�)d�l\�v�27}`R����k5I#�),�o;3�!T)կӁO/�}IHD�˨b���&�)������Y�!k��D�L�q���1{9�l�*�ӖZ~>#bHE�_;� >,^4��M�ψ� ��b� Q��u���n�qSg㇍��p�6�@��>L���XP����?-���I"��F�����>�/,
����>���i� ��9��˷�K)��,��_|�#�[�(�OAtY캺ab��E�T��3`8��O-�-\��ջg��vϕQ����s�7�$����6�ی{C���4����k�^]�bz��Զ3Oy�g���i���;/.���8
͹gM���]T�訰�o�Js4��=��,�-������@�[�=G�}TG�j�PH�3�|{�d�k�B����W��ir.<O�zy_[�X������rk֖Ԭ-E5��'���&��{���ݚ�[%C��+<a�����ތA�pr0WB�ٰ�T��*N�}C+2��C��J ���*��W�%N��l�/ e�Э�=�Sط�ܤ�#�K�?��E�Iv���?���m�9R^��#�?�k���<���Z/t�FƠ�xǴ^��$	��Gn���"Kc���(�cܲ')W.�@�F7�����F>	]\~�yA�/D7f�hy܈�.$����
�{;G�`�z�E�B_F\�G�F{ǖ�Sw�$�W��ޓ:�#;훕�,Y�:��n�
2��7��7?YPcC qOtj�X��"�r$�Es{�H�������s�4��_#���km��F��.7@A"������:�|����;��� ��ϔkw��Xw!c��[FT����O��Q�o����E�e��]������L0Csp�-v8r�s��h>u5y�'�#��f�@|�j�%B�UdQ%�Z��eT�z+�4�
x�.k��.e޺B5�Z� �\m�:�uF-?Ұ�z�~���U ��eE=wF����/t?>Ð�[.���d�߶�� �45��8�ߚ������eʗ��u���k:A�d%vB��dO�^�����v[y+Q q��ݭ���*����қ�WS�.F�)��;�a��Y!;:sim��x�y=��i,3w+��l�_��	,��<���,2M���Ea�0S���"=:k1�8'78�)(-���fݪn%'����rI7K �}z6�d{��'�����(�D�2z+4Gef��<� ��w6eI��n�N� đl��-� �z�d�A�`�H�$&�O��Z�:X��Q���=
8��Z��a�������I7�=�BFp3>3$;�������!7'2��g��F�p8���4� �ӓ�k���Ռ@�D��
b$)�P{ܦ��� �A2�Q�#���č톾���o��THu�جk�`��=jVY�+v�˺���CN������2�-��3��*�XK�;��fu6���2tC�)����qT����%s�׭���!f	�dۄ�y������Z;~�?�U��ϖ��9����B9���63>H�Y ��w�]Z����k�fy����P\����Y�)}@9��>C��S�cP]r&	�{(��'�zԆL/Z�64��=%ip��s�h����B����7���$ǉ!�g2xӘ�n��⃬6�f�P0doj2xC�!��	|إ�@>3���U��[�j��t��f�9jGq_��r�f,œ��5F�p��������_IN��R�E��J��.w�)�����#��7��#��Y-i0c��� ĄhB�v4w��m��#暺6(/L>�!�TG.�-Lz��*g�{��^�LV`�`�T��h�Z�uK��d����@S�8'�$<�KG���vѼh�2
rr�͏MZi���a��8��������ˌY,��ȑ�����5�KJ@���D��ʬ��С�����hT�֗��!�l�'����q��c�Gv�w@sڭכ�Ma/���G��G��.r!ݓ����A��7��2KƇ�)�^�n?)Ƞ�&u�?�N���=ς��pnي0�>9-���:��]f26Kqu����>�5#���#A�(��m	�C���ލ�Y�[H2�T��]�d�բ�f�Th�X?z-)]6ۉ��蠸���f%V9?«TYoȂp�A�2����cB��MDj�hA^��M,�Mh&]�ɳ0/��R��<�F�y���z���l9����p\��5~���ts���!��k��k�D�|6�˱�Z�_m�u�>�a)�=�c�� ѳr��
���/b���w ��n-}B'k��r�2_��ޮ9��/W߈�X�I�w��c;��*�-]\��a���H�@�� �ab[��	U{� �a���QҢ97	��ރ1�R7��p��5 ��	����tc��_��B�"hä�w�����	c�R�\�'����lW���k�DPy<�,='o%���?y���4�A��Nv��ga��K�%���1�A[d�����F

�4+��^�\�$ l7�q��䳬���K�I� 0'|�"���0��f��ď�>(�`n�qG���JE�/i�B4�7E>_1���5G#j�*�MDq��)�혝�` i�o�����BU�o�U�)�:�D��S䕹wTx!������II����7Z�����