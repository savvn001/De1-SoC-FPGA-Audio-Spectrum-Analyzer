��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	K���r��"0	�@��-2�|#+"��V<5�gs�Z���	~�+5rp�Ur�͘�����_
FÝ��PZs�\?�qU���q�>x&D��c�M�	]��X5"yd��Qӌ،��R��|ʔ�ڻ�LQ
��v�;V�q鈳JO�*W��?���s�1|9GMȦ���|7ϰs�(����7G�׃l�GF��*��7u��"Bur֓�sշ�.�����	�:}�K.��vz����H�Q����@���P9g �d��z���Y��<��)=���{X��x�~q��Ⱦ�*h���n�Ҽ+�r]?�sNv�b�1�
��˂x����N��oap�Woj�N~�`�_�������?u ��� �[6�*Z7�9a@���xy���� 4�o�f��_D�Xu	NGhj�F:%���!���Q���P��������Q$��i�G��m d��S���@?"���ȲV��zA�*�U2�,]� �(�,��͎��r������6dY-M�3<�������FJ�U��g�!�|Kp�Ҧ��l���A+`�p��T�^85�/����q�5�%CE�Z֞g�\�O_AJp�*�J�^k����0dȦYbtZ!򪀖�䉴Y"����S���f��l-����X�!v��y^��b�@F�dD
��ӿ��p��w\~�� i�/�"�o\��~e�I݆jYnK~�
\��|i��-�L��9zJ�L�d>���Ո�j��c�����zj�Χk�	�QB ���F��
��uړ������ia;T���P��A$C�r�ʅ豧���2x�\W�;����,˸d��jq�x-D��H0�N*��'u14��;��B��qoя��,����"��wm.��H��ߴr*�H� �r�+ ��7���A+i�����.)n�Ң"D������ϒ��f<��r�I�|j�X^�g���3耻�5%i�,����f�k6�3z4�ׯX{�9���� �C�~R�e����!�V��>c�&�j�eN�
,�鹞H��;N�pw�:��9�x�&�T*q�by�3;����ńe�>�oC�.XJ7Q�0s�na�LEv��Ƿ��؍de��v����C��0x��S�{%����E�sa�/C�/�m�1!~����P�(���ì���1#Y��z�d��`��̀vP�4���AVx;ǿ�N�rs�ţ�O��x���,�F*��Σ)!0�k3�:�z��E]���ʖߢ�J/�ře�hX��ծmҍ��)���6���~�x3^�)��}ѕq7旆a�d-�#�v#EK�nU���vG�Ը��k�C.�Bi��@\Z�)]��I{�ѫJ0&o�̥���o�T�qj�f8n�F��huͣ"R`4�Nb]��kG���/w������cѴ� &�D�~3��Q�5�O�Y���Zd��m�F��kdx���ENX��.٤�"�����=zUF�?�!�[im����(�[�(����8Q1v���s��an�9�d�',v� 2iP��Z�vC�x�D���e�۠Q��M�*,����g<�aK�O�<=�7�O��U4��fb��.�-b`�.�I#��;�HV��͇#�g�!�J�:��&sdч5�%Tu�*o��a���pT52�� z���CSq�8	���s�*o�]Kl��ZsL�X�����O=7w{6�*ħ�`�^��&�|�*�в�S�o�Tk��o��̚��*D�4Ky=2�b�qY��e[c��g��Z�d�� �b�r��(#���������G�[o�o8uv�,�Z� �[�LȜ'Yx�؇��ap�{�m݋d_�7j�iלo3�