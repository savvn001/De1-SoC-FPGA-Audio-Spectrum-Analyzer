��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D�8��t�]�&{����F��V{��8��0�b��P���o���,�<<�tͱ���:�4�Wqśv� (;G�����Kvn楯<^��1�	ҡ�8?���'o�|�pl��s-)��朏�j����-9�����<�y�e:n����
�LM��\�Z�T�'��1á�b�on�I.-���# �K�T��G	>\���[�:N5���&i�_HQ�^���Ux����q�������)�j��Q0�"w�����Y�����.�^u-߽N�#&^�Ԋ����Q�t����U����,�s���W	A .4�k�)*]&q3r��(T�ӎ�_�c��)6�8��p����,���[C˛�-��3&H�Li����ꏬ4՗�����:��m���]P�Q�tq΂�����N,9�=g���R'�(;����w�G�y`�3���㵹L��H�Ey�\�c�'��S��8��IM$L�kK�=�I���n��4�{��?��λ9��'��t�1�_]�M�+͑"
�N����<����׽	���k��tn�����GN�8��]�F�@���%N��U�x,8�5[�r��3�%O�����^�����3�J��L��h؝S�����LN�����
8w�6�VK�훮x������5A�Ec ����w�lIR	L��������Q_��<������7,���|��;V6����DK�1��O�k�~���j.��Lk����LՏ]�_��{@�6��4�3lŷ\ ���mT�5D�E:9�� =��׮�r?�� �����#�������G֣{��=�#�����5i?���Wj��9UI�,�~J���l��x��r7�Tscl��R�oN��j�&����C3[w�(�W����*���gm�vE��d���5�r�T�0^�s�1��`bh���aK/���yW��ۼ�[��8��kǼ�CyP.��$SHwnO��p%k��];iZ;�4I���95����P����n�}�^�ً��"��*/��He=�h����d���D�����GYW�c� &	dx)�&F��i��8��4����^hA�{�@6o�s��^A�L���=U��>�"5i3�Q���!pFy\#D�o p0iQ�#lmiZO�}'��ǃ�	mk��R5�؝X!��>���W@w�Jp�t���;F�l�&�qQ���s��ۀ���#�E֊�;"�A��%Ƿ�6
��U�B=�$�s�f�c�W��Z.�hz��z�" 4]�/�����j�r� ��C�n5^��h�B(�p����zYv,�@֖��c���eEv!a�嬠�k7�%-����Og4�)���\0�}wF}�G���&֎.eE�8!�a��5MK������
c��Y�8M>�>DI��36�0�Z��1tq�C^�U(Lw�7�V�+��)9+��������C@�}�OWF�G���Ӏj�S�-���ۣ������[ڙi�����;j0I�s/k�7m����5- �z�
S��8X�1����2�z��n��[Ōs?�4^?a�<�}IWZ<{�>�uSw}XmYΡ��n`-_r6
]���x���\m���@�b�Q����Z����ͯ����$���!$��C-�M7���Jk�*B�r�cʡf���}��@i�q����Ȋ�\d������ޠ�;�`vU<C���Ic�-�B��c�(�r+�1M�0�0+����}�������'H�E۬r����,N�����i'�*)�W8�{+�a�j7��jk,Ea�o�\NS}��������y���G�%�?�<<*GP����-V[�{���,����ݶ|/zxѯ��Ƃ�������Y��T�U���,-U�T� S<y7ᣂ�n5�J%����ʒ�/��6<7���7�c��;�N3�<K��>c�=I�~X�Gߎ;�Q�%A���* ��O�����}B�e�vV��b���ؽ���i�/?�$�LjҸ���u/�����]�&dT&2��x]s5Ώ�Յ�*.~ګ���-l	HF��l��d�T�����$�>HQ� 2�&�&ӹX{[u�!{�GA?y�~�x/H�Ng�0s�w�<ǽ[ d)į*f"i@)ђm��9����b�rpa��� �r�{�RVփ8Ϊ#Y��j|ṣ�g��W^'���"�)d��a�!uN/&�n�z*1}a��l�V׋�^0Y"�.��";�%}7Fs�\�[D�r-b�i��G�Aq�dD�Ӳy�!{��촡��f5S�H$w+jG\�*u�,���������/@�&���)*�����;�ITh��aL@���x�K��t{�0k��F�Z��j����J�E�"�l��6��㎩��<ze��}�ǈ/���>FQ+����e/�f˺�����z���.ƞ-��e�� #��K�q��1�iI���H�~�;�g��I�Ɇk��b�}I�x�#��%^��K���:��[����o�q��:��/bЕ��:ޑ�8Ⴘ��˥�h���:˙�ח;� ��7������}��B%���]����W��Fl�X	�s��<�z�]��u�1X���n$�*ؗH����|����Q��ctu��KƕS����l���9��
��E��1�i�t��у�(C�k��Ĉ��M��7�D4.�H	�e� ����g���tM��.��'d�*������F�վ���\X�wO����1���Em�s���{U���(��^0���Ҡ���6��2+3��f�� ��.M���#PR���NF���D2�W�*1Ϧ
�8� -`fn��۶�^߱��������٧�Ԝ��KM���_ΡtY�-[�s�C�HU�W~6Nb	@~���ܗ5@$H���2���B��{qcY�Jԥ���irw �Y�cL��
�z5,L6��>�!��3걪����7�V� �G3�FB�\<��O�;MkJ 3�-b�hۨ�6t��L�(�f��0W�Jo]��!�B9��9�N�����!Y_��ni�pc��i="����1B���K��1��Q7��Ƃ��M!XB�L�>m�:��$u��¦���,������{�&�4z�K`T�r����1�`;�e���A��?�y&�WE⊶�|�ad�H�T~��;<���A�qUD��ш�1�r��hDY�5]CN��4�bS1j��4�J]o�.z� �d٤�a�6�b�[R�M�;!������@o��t
�źS�+����E��zȜ���IBA�ٛ{!��7���k�{���:��A6X�� ����g�`��i�(��� u:�X�$w��w}�|W<���o�^�q%}�eӓ$�h�����=���r#t��G��ums�>v��|���:�P��~�'"nd�`W��J�c��&��}�ҡ0.�B�ͮJ/&����n�=]�5ά`e�m��ܦ���%~���=q���d668lL�<9Z
7݂��7~�����x��#ԝ�3���`o��\̋�mQ�?"�,x�������dv��9>��d���� $N������V��c{��S����3�k"%S㑤:��t
4⟍T��s�Y1�V��u��f����~���+���r�}#��j�\z��d&Wt2�.��'�r�-s2�Q���Y�{�ė�7	��l�e�=���lޜ�!��t�%��d�v{R���+2�&<�/�\����bi���	�7L-@�ī:�R�${�B�W��Z����Տ;8�t�f��C���|�?�Ej�쁈�.9�i�]���}�s�c�Z��s3'9�k�VQ����q��л�Q0��}���}����%D:��4��>�����ۉj�����b`�S*l�'6&*@A[X���r�b�b���퇯U�6�P���TNV6�i��S�mܴx�tV������O�o��D_7�4L(��S 5�����ٙ*J��h������Bo�uQ\ ��X_c�I�"נ��R�SX�T6{�+�a-J�����'%�,6-*9�q�<��F����O�J��:N��_��4���z� ��y����ԥa�×L�}����Ǵ~g�>���RA�st��4����0ny`XeF�\]Sj��	�Xh֩%�Ov��|(���3R]���G�����=i�!Gx���@��yEWKV�,��K�a-�W��KV��������0~�Q}pK��q�tO����N��iÏᅤ��O�Om�xX��N� �]�����@\�aX`N-��ʜ�4"R��M��v�!�"���4:Gz��g��=�[oFyy��tG��R[}Z�1\8F5F1�8����K���f<���>��~����,I�YI�/t�?0T��X�f��6�,��zQ����k�ۏ��R����PM��h�jp3�>�Og�xw7(�^v�\�]�8Y�M�r���=��:�yd��x(��Q��z���@��*��=�~{JM���PMȟ�*H��\f%�츇�ws����C@s�ґ��#JH��6��ѸŰ��j�{&���r��~J.ܑ���ki�Hp
���ڞЖ�w�rv�6!#d�j+��pf��FjU���k��n���[�0��8 ��(�;��Aqw��s�y������� ���ٓ��B��<����kZ���ֽ*/���r<�d���gk��7��~�bWW��%q%�c�7��j���)� �ҏ+@��0	�d.I6���[�H��2�4���v���^�������ݛ=�����}:��O�EJ^�y,��-<�THj�R�&�.2>�%{3u�ƫ �x�Ͼwr���������`�h.���N��٨}�DKw����kyʋc��� �t#
%\c�Q��:fE��@�uG����V�*�Exɋ߃�6ċ؇]�Kh�C@���R��2�a͊R�Х�G���f��4��B�j��zU�����7BzFĈ����J����ܒ��
��|]D��wW��j:[)FD�4@�C��*�mFrE��Gq�>���g����[EA��j]u�O�A�ۿ:��Ug7�M����ӓܗ@8Yq}��M���*~ox_�����598��6?��g�8])S���d/�B���b5{�.�IL�ԃ肸�T- ��a��jM����|�l���p
$m Ԍ(t��ģ��%��k�2q1d�(��b�k�ux%6��DC���w�u�)VLꝒ�k�4x��Z�~k�v��"���ӥ�«E�5X�����>�k(F�,+�f�U�O�
Y��/fE:���g6��5%�Bo8��M6�̣ˀ= �2Ah�"��*�B��C��75�Η?�d�T���ʄv5�hL&k�:�#]�d�FX���H�C���/���E_8
��;�8�J*�Ω���6S)Ä�ɯ����\�27	����-n�N�ZЖ���z�oN�AR[�͚����G���ě�I�r��i�@S=���|'÷��}N�vj/��wU��m�I�+�(4]�P�y�ti0�+���
y������06�2Rz6�M�d����)� ��늁n>���{x�/,��Sk{O�QjCAHwi���*�_�ՏZtvc��~�+e�%�3uHsB>�.�p����&���T��R{=1{&�L΅�ƭ�Ѱ��m��ַOQ��эVg�VT6�k��$Gpy��s/L1^����d3uF�j����*?ȣ��#�UQh�ڍ��}	4�%�׿�SK����	�}�}���Jf�"�$�
�ަ�c	+6|'�����O��i�X@��:LU�Mq�팚�}�|��c?��9駱���q����",]�����h6����%E������D�Z�7�(֔ ����u��]��Ro(]�y�&���50!҉e�cd=� Ï�s�q�ԃ�,/3�)�Z���/¤�"��\	�`:x��4�O��P�g�r�A\�H�n��#t>�{�^N�=]�ʗ�udI%.��=�R���Y���� 7nn��.���?��V�}����[�l�"����<����Мz/1��t����*����lp �y��h)EM�\�Ȧ��O�*�Ĝ�]��K".9Z�P��v*df�i�'���P�n1�@�S��[��j޵�YՏ~+r��,e�Ўb�˯ae��u!��x�K����Lu̡/n�{�6Iy�C��+ٜOk��ѝ��,Q���e���*��N6_�����fwU��� �%�\�{��r��,�4HL��
�`ʀ�ϗIx�B�Uxd�|���ݡ's��;u������j1�J:�)_M�?�dj��*�����[m<ږ0�͵����WO;2��c��W��U���X�"h�]�N�U��P8�g��Stq�S/��]��ϣ����=u�������r!�P���
��6,���ű3�쿠K��z�Q�J-�>7�֪p��|�k�^����s��E�N��¶�J�~��$<����v��\��'��4Lh\Rk��AQ^�	3���ۻ���*h���e�-���$m��PU�,�
���û�M�烜��SCB9<���ZlV�kέ�vF�(�+��`	ٕ�]."��/��1� n���_���<o&$i�\_LA-5�AhF*A�&V�lGGH��2����l��ԧ�I�b�Ue�
�j�S�^��T��U�k���@S{��O(h�����	}3��Z,0ǋc�q���B���ٶ��$øs3�U?F��q�`���(�U���ΏQ�9t�2ц�z8���*BW+`{=M1����Bt��������I�O°�����G񀹒g�����40��G�OTo`��qT�6��p[�;�&	q[*�,�Q�N�|32~�ڐ2)����� ���]�K@u��q��}�/���P4�`���do�|/
�%_����=���{8��kiI���9�sYi�c��䱟o,�p��s�Q}�C�.S@;c/fK��`�����	���r^�[zҾ`�Q+ШJ�N��#����U0�Q&���jq�4�'�wW���M|htP����ƌ�^Q,�I��
����&ՠj�̪��ǖ�g�Fj��
%W���Nz	(��2([,�&���=�o��8����\FS�/s;����/�>Ud��:����T�i�8Fxw+.���Y�P,S���|����!k���|���<����ٍn���A�ک�Z7�h1V��w�7�&�C��\�3�@2�C�l�4r����#�q��>�.G_�g�s:q7Z��W�I�;x80��)MP�X#�O
�_����Cp�)g�����2�E��H�� ��Z4���!��'�k� ��ظ��rW�d?����(E�*"��k*NE�qu��{�AfIK����v��ǬU�Jq�U�'�/���O��0����0]�2К�9l�8-��u�*JΘ@8Ĳ�HѼJ������4���:��c�e=��B���[����F��ƫT�B�o�D��x��;���A�ۤ%���\"_�&�Ȇf՝�����`��^�)��x�U�b�v�y��k��5����qQ	St����nE�QVt�L]	6|s��ܻ��@ib���J�a���
���'�\��`H v��ѣ&eN�F�b�>:�JAq�cE���l5-����;��-�����n��F�yu����}f��Ɛ8�
����
�L�QT6���C�}N�:|SW�m�����
�CDa��X?�2b��wW|��^�9���J��m`D�-�cF~T��84�v���	���ũ��y���K�V�J�C5�-gܠ�ŝ_��|lp��S}�cyv{_�J� w;�R�?YC�8s��ԣp��Y���;�T�o
��z�J2U��
��E��nߥvV�Аg�u�tb�.�&��0E?�?�\'��+#��>��3G����u��/\B��d{�q�@���
UW�����x�a[�P&�N���e���l҅�C�^�(Lh=��
V��˙���w*j�-�&@	�\�4���zC�����1r6����B�����#bwZ,�KQ��>.�v�o��c@2|YҐx |N�a��#Ā���S���}�q���D��5���� ���4a^X9R�;Ы������H+�X�-^��|}�͜5=���T�[x�xok3Li:����,�{�&U�����'q���՚���2Z�5ܛf �Io�ѽ���ɩ}=ﵪ>�/V���|\e8spz]����޼���,�^�7��t@+�5r`����=�L�d����a6��W�3���ò�	7d�[�L��I�-�U��`MI�%i_п$�/Gt|S��L����� �x�
N�D6�4D��W���,QWu�����`���Ew,�9-�����
�E�d���.e���_�k��|�Ҋ��^��aC���=_o��pܬ�c��=��ЭZ[l��a��E��e.GM�Xn�6an�Q~U��q�[6�����ĩ���@G���0�%�$��z��Z;ߕ!�V���:��U���R�­��P�J*=�)��@>
���a��7���,���%��\��}jg���X!yk$Wa���Y���.	�Y�N�����}V���dW�^ă�C<�f��u�M(&T�IK�B����]ݑ�����88�Jn>�����J�o˾Y�V�b�Tq���!ĩʎͤ�ث$W���SKI��Wg������^��h�n��b�G���k��?�1��ZM�ne�&�yI�?'� ]fI{&��!�'k�5D_�'��y�e�+�b�S��U�Q{�'���!wӟ8͊�T�I�^_�!|\'E�u;��Wg]p�� ��]ud�x`"5C�9��7��8Y��"��N���������X+�%@�p���W"L�"bZ���;�l�t��B@��G�t��<����P��G8;6�>;�yTH������F"��S���iQG��e���W�	���U�j�م���*���,kRd�y�?��c[�1�G:1u��FK���B�]�N�,[�e�,���pxp�x��9o�/�	��I��Kn?��6�jOv����X���WZk�����,� �T:7R2��t��e�Ӧ�?i;����]���A�j�"S��i�f��W3��k2���kbA�|�x�~ݝ��W(|��J�m� U�<f�(@֎Ģ?�D�1�c�Htw�ˏo顝�����:���[��(b+c T���
*o_E�b�s��9K�Y�����@P)75�=�T��*iI��_��o[~�Q�iMm��tG 	�N��1Ni.5`a�TI>3�	+�3;A@ND;�,@���)@���eF0�8Ƥ9e6 
mi�g�7���?n5W-��K6X�D�"��x�J,m�v"�m�C������(Z'&K���ݫ�:�ys�[�f%�YcOz魡���ލ۔O�� s��חV�S�9mn���e!o�?�W��W�w%�|K��8\j`L���g�t��j�Ϩ͢1�� a�{�Èh�y쨕�Zk�mg���y���3#�H�*�6��%����d�n~:����2/�x�s��]3L@�?O<J8�/�	���M�� �X�!�D���-�,���� �\�v���Oѭ�"���m� k�h~^et��[/��bZE�lʌ<�k_��׉�����>�~A������tt8�g�������������%��W��D�����j	��c]V�]g�"����}�������w�&k��+�����y�)����h����.���L��˚H��B�I�;�,>��|���9��O���N^���(@��RC�|�oa�f�`����u����V�O�� �MX=���S�.5���u�<�>Z�-Ŏ?�����y(l_����5Na�&9�v���ո�0�s�b�/jk⇁�,���T�W�Dt�z:D��GW�96/W�$�NΗ�l��4<=j�P�������CO(�ۣ�t_`ed� "�˹Zw��3�� ��}Wwy�PU�\r� iaN�ak7�́�qGnP���[�6��#��A�ê:c�v�&��I�]]�������G �+�Q|�#�*�C�i�n���%�5����Fa��ڢ;Oż��oXm�1�p���!Es�@�Q��#�؁��������/^��Ѳ�Z"�:����� ��˞-|[�'�ܻx��SM�	����8��(�D����M���Я�::_�*ʗ�DJ��;bq=H�cZ��K�����e�/Թ�Z��jx���({���~�XRb}T&�#O��*P�x ���a��7�o�ͬ�]I���3�ah�G��qn�A�+!�s��Þ�����%��՝#��E��H��d��ntmp��&,sح��(6�m�>�&����/2�Bl���l����V_���h%m��Pd���\vvk�E᭤� � aq�k�;��D���)�ɧ������g&������`�����w(#�wP��.����;AQ��,ݵ�$i��"�����3L^��I�Wae"�Č�_f�N�F"� �l���%�y1�	��u����}˴����!ȭru˴���k!SC����f�j�4�^ׯ���$��j�9�����������%ܾ/GD�y'=�l*��:�
V)zk����+z$�c.�S�Y
�sB�2<q588��~��_!�5]� &�32��EH��2��$N����pn0Rj߽��{ �'�O��Fe�}`�����Q�8�:V��Îi,�W�(~ZE���3a7��*U+�����v(bA�(�27����6Gh-���o++Tpn���]�^ϭ��RZ�RD�=�)���k��q��۝ϧ8��h��`��gꟌ�*2y!>ݥ�b�x`�@��_$1���8{������g�&��_���}X��^ﲃі8�=�pQQ�aaMe��*GZ��*��$��Rn�q܉T*�?7����� P�j���<�+���ċ�A��@�����CI��BfEfz�m��lʍO3A,W+�Vn]r|�.�,�R��$�VBʈ��
?�r�8O��1��{u2�U����ne�%�f����*����Z�l�h"j�3�h�1ȸ�b����%���qiRϲH�s��]O�@����:�3�� ρ7�Cl��MGT<AP��U��|v��i����P��d��v�5�bp:��;-@�WkztZ[�Fy�K���3":M����]�xy�5��Y��/[��b%���?�?��(�a9z@[��βo?ϰ<h�\�'��զ��5�ަ��_�$m�!ɨ��6�5��A�����p�a���'�X�����;]�Z���2�Z^eԮ�ʚ�ayP�O��e�^�Qn���-�Q'�1�zO�7�"c��B����ğ-d*�4�B�>���y�OEwz�ó@��+��� ��fk�l�0�֊Yʆ�;~B��o�ҩY�=7�n/T��M�7���4Jq�dO����.��D�Qr"8��о������$-��{X��c=�&d)j������d>ϳ��[���3�Y���y��t���v�\Lō2��RI;�{�v�-����Z���6+_��6�E�j���ᶰ�qvI0�=A-+4�"{@oGl��������&N�xr��T|h5r/�W�{M��.���Ju��ǉ�B� ���¼8>��M������6/w�CH�/s	`1�ދ�݌2@`?���jK�_����XA��XI���J�S����X��Ę��v�K^��E�U�)��v�'na�<�k �A�^{��g�:r����g�W�aD�Avn���>��}���4}�s{r�N�4�Sa�t$a���f�.x��sm?���m�I�b�����Z�&x��#��h�I2��Kb��yV,Xs�C�R/|�0)!4m����̆�{����R���g�K*|$����1�C��7� g� 1��x���_���c����{#ƨ�`^N�i���$����~�3J�2ƂI�76��j�E����O����uF�ޤ�o�q��ې��*�w#�s���e�H�U��6طT[�:C����fp��Rs3����E,-ID4\���Q�/�� 0���}F�q��|�e1NÊw����p�SzDn��٘��ь�~ϪY��"�b��JO����lnr�6�a���҄��͐��d����ZW8a�$��l���%��Z�*�1	td�XHΠ�a4&X(�OG��rU�u�L�]��i}�^a�'^ƺ|~�;G�ďzi�Ml����n�} �ಣE3�i����]?�B�&��	��᭓/v����]l��)&__�߁h��籜�o��g4*��LM[���s�^��֢T�4�|���Cľ3c�0�!ܼ��o��[�^���f��I���P���Bd�U��T˹�����U	�*���`;PM�3��R�p�2K���s��8@0���Ŕ��#�9[�ط�A�	�mXuތ)1O'�	c�g��hV}�\����a�S���V}|�(�i�̱���G�q�h6���j,�Z����@�@K���Q��vJ���[HXaz�ʟ%�bWc0��J�����d<�.�z�	S0�:}��v��9��h����҂�0�����|w�����H	�1:j&�2&��bh�B��٥x�4+D4�U� �]�y*�Cs	��w����b<����i�R�}�ƳamN�[µ����-� �����&u��|Ƿ�W,�Ȉ�*�E�)MF�hv"ġ�Tk��*?��dW�Y�p���|Q����>��3궕o�s�b��Y� ������PlOV×(k\+9�k�6���v8�P�A���
��6R�~�y<�Zv�8 v�o��4��!$Ґ��JU�=�p󉨷Ps&0-^�r�}g�7����QF�w�)6#/f����c�g�-7���S��L	{Y����0鰻A���i-wmsL��B1@{/���.����v�lx�d-��;�&����*d8��>g�I�'�]m����Y�@��*��bA���m����\��Ċt�@�h+"��JI����K�A��n����r��>:&�  �;�`�'��|����6��p~���N�f) ����ǒ��9�d!ƈ����'x����cX���p/��������e��z�>��
?��)��x��{�ڬ��j8,-��m\�0!Ԝ�mVCX�w�k�Dz"���B�]�)�e$��}�x�^�f��Or7���8�g�a�E�-��?���u)X}=�Y��������F��U&��,�� ڲ�|����/�v$=�	v�HuB��#���'��Ū%��Ptl>��^Zl)|��ڝ�����;W��@s"�(�TX_Y�AR�01���܇��)a���NiN��G����.�K-�� A'�m��&���y����{xC9܋�Y�U}2�w���d�E�]����hG-��:�p5�4L�Z�1
�ыfW݈
�KwU��+���O�8��[��qͧ_f�x�n�:�br�w�|�|:�1At��L�/�tO{U��ZЃ��B �m�,��k��?�\�eWn{M��#?�P�,�t-�����5�����0X�WL��7�Ȕ��H�-���o	���#��I̷]E�G�;7�*d����3�ݯ܆��-"j�a��r�k�g?B)�	������7���!��:�Q\��6�I60���[[Kg�<x!I�m�e�K�(�Y�-C��o�z �&3n?�l��>�^>AƇ.�V�6�+���A��௅!	l��*F*���Q���ó���$I�/`.�Vf=V�5R��A蠀`��U��k��=V�:i�e�:X���9�"����aS1v�(�o?߻O9!���b]�b	��\��BC�},��8��{����9�+U`��ߨ_�2zƳ�V�F~ �^�_���eOO!��[�������)�̚9G��X�Cp��eb��s��01��/!Xΐ�:�|�Ҩ�<��ؠ�CA^�F�	LLA鐙tq#�J	���\ׯ�I䲝�)Z7���0���A��U	�����7j91}!�Lp�:�=��vЈ8��]+S2���L�9-jDʧ���U�*��Nk{������43�w�Β��Jh�Y86z���_r��# �'�A��U� ��!I���
��V�C���y$����8�[=)�?���}һ����O6���Bζ��47BFw�S��7�L�fӻ�y���r�mD�Z�~��C���l��`vSqՊњw�m����6̏�GmyBprς���ֳE�B��v��u�p�XHt�+Y?�+��Tu���SU\#�]i���w,�Ӟ�sAR��<HYƆ�q���i�8�]6����G騢��x�+b?9T<��!V�1��Y-,�d=7$"^:3{���sP���89�$F�"����Q��|��a�����|r�ߍ�[��l2�	q�祲DI��&��e�fV��G�iv�����Ty��r���1�?��deD8Wg�'�7K Υ��;��.��]2E���sґ L�����8U;�YoC-�PRpY�o��Շ��x��/q��f.)��@ð�vr߯����I���!mz�&��C���*ޤ��O��@~�bt�.f!�'0�b��MGF�x��w8<�vd� 6T/��PY��\����{Af���Z�S�7-�����)����C�ޠ]c� �'�q;
��^!錭�~L�iA���k��T�Hp�(-=ۂ7������q�7*t��8�eWan%���+M^0��u�\_�+,�=�ht���&2�.�qM�L~�JC�H��N�F�^	r���1�\��g�w��
�ĳd�� �{Bv�{�V2G_�Q�~BaϐЊ�<������A<Z�7{�S��.��Q��U��F�"Ua��޳E �|�B�͜�"+�R*���Z��R%�B^��C���4�fp&���_q�.WLx�}�}�m�K���z0mE�n��������_
K�G2>��j雦^1+,�~L���`a)x���d�����wB2JNX��&G���]���6�<1Ȩ�Q���LŪ%���]�ÎS�.&�ֶ�g��;�^��*I��P��\� 	���j�޽���
֒H������V��#w���������c|-��1�)`��xp~*f�xM��|ű9ɾ[�Az��b/��c/Vn}����V�/FḞ���Al%@m��t�E���}�#EM���el�9?���Ӊ)Pj�?�=�Z�U �ǹw@n�ܭ���d�L>>�`����_U�~;���~�ՄJd�3�	k0)�6-YȈ�UPS[�2�/C�7�ݺb�N������@9.����=<�+J�����Tu����^�g�D������C,��9��\�k�����Ѐ��ٝ�ew>a�⟳��s���SŤ���ڙ2��i��� x�����b��i�|�i�Q�����	Z�`�Z��x©�51=����u�JX(����A˅�������M���D���?A(s`�j���K�g�Mj��8���k������M��\��봇��!�G��)щf7��k����^����6���U�9��NC�L�o�W[�Q��+��N�(i>�U���@�!��ך��g��
�cc�nX�:	_&����Qٍ>hj���E�to�� ᔎkv��Ws�6��X� I�7.�p��M�Q�tho|��_C+6	t*��ʒ�Z)�*�I�!���r�b������<t����j�C�]~Ɓ⃗���W�W�m��f+�~걂 /��c|[d���\qU���K���sR���7�j�4R��'���<z���ggD�^��sF����o��HBs�^L���{Q�9��2 �<$��7�Q3�9dm8*|���Ƭ�ťf�]�r�M�r���������׈�c�g�9�mg�m����}G�Hk��3��Q�V�r�[�K����#s>�m�h
D���!|����lLN��� F���f��9=�y�R�v����~�]���6͕J-�c{֖�Y���g8���Չ��G�X���G:U%�{l~f2�q�ea2��NҾK,���N/δ��|ဌ�d;��fd(��d�����jU!�
+Ov��U3[3�C���@ں���W��\�APj���}�Q�E��Uܲiۄ_���L;��J
U��(��t&@������O�T���7���<m�1���>+���&P�P�OjB��TY�De�R�2	�׵t�&F
���[ę��Y�b����<t�M���M�*�	�_�J,���c�Q}�K%�=�sXT�Eqx�闖�#�Y�{�*Ί��*ס<�2OߋBuE$���> ?Fg	�%�l��.���۲O��S!���.��E��j���������������g�w��XM=��+�E� ���c22����0z�M�?1i���)A�����x夰o�(��3��N]0���6�-m�$B$���IA�¦,6.ADI /���
D׶�Br]�e�����0�=boX��D�ށ9����u���|�;y�Ň+S�i�Ȓ���|}�<sϸ���=���8�������m���<ĮS�D)�j)W�}C"�pΟ`9�f��\ʓ�@�-X�5���� ���! t�
��%�ձ֖��(3����G=D�#�&'��<U=0��]$�:{���Li���"O�B��F�X>�3�x���*��< 8���l���>h�ҏ!�iH�����]ށ���O]%�G7��ΐ9���X|_wgSWa�?�h6�~�?�k�EW�?��ՁݞJy�%���:�u�Q^�/g��0�\)��w��M�����>i\�M��BǨ$�CXw�H�mݞS d-A9R���S.�`�U�d�m�6�E�aG�G-Vɑw��6pL֡�z�\?�؇~1Eޞ5��<duv֘��$⒁W�Kq=x�����T^!%P��5�2���]�'�Jfm�-G�=5Q�2�ʱ��Y�nR�o��_��Z%�\K�)x3�^��ǀQQ�AC������cx�(��Z �a�v[���ءp�:�de,�eFxA��"��O�����h�ޯª���({'�\i��,x�0�[�Ye~�=�(ȧw(> !K���m�o���f�PR�qx���[⣺4� Dn�t�ɀ���HB.%+ΈOȲOJ7�7���s2��)��q�� !��l*i��+/9�cDMvX���k~>�8I?��ϑ{�E>��a��TSO��H���?S�qR� �p��Y6i�}��@D+b�%��@/z0�(��#Il�Z�%D�����onQq>V������c��>4O>R7YH�e���8��>�6` ��V�Fѫ���!^6�Oi@Œ���G���_X˩/���]��"8�K�1h���2����ИaS����: �j��2�iQ��穤��f�ö�|���;5�ϲ�7��Ӓ��d�B�<��y��Kz�T"��\���.��80��a��\��
����n�7��&��m�U�3Y;��cd;����
y�9����^ֶ0�1z\4Eاp��c��������؍���k��? �y\����/9<���\��VaL��'�|c��<9r ���ݞ|��������Q$��Ǯ�1V�ld.{D�&r���H/ 4�
�ֻB���Z�@���N^�o�;�V�E���Iiz���/�E�<�L�ׂ�J�C�.\��}�I]dH�St��L/���8[+n�T��K�DN9 �u<�Cӏ�>﨓�Cg�Y��<}�V��y���tG���hQI�����-ꭜ�E�0�����Y~�0�rjb`�g�#R�Q���h�^!�;�9���	�^��S7�K,��t�T����Z��(zx$��<�,�lr�&����ǯ2x���6F i���7��$�E����n�=4mHU@k}%���.�������,u�])� x�r^8r�>����زd-��+{Þ�% ˭��˛@��~�3,ݢ���R���M��3p������9� 4����~VS�٪�6�*�q��R�Ao��ɣ� "v�F��Zg��F��N;"7����8Qil�~p�$"�GM�rL�)*����R�ڧY�.@ҊaN�W2)���a�����ͫT|fhd��3"�ފ��:��Z58)�A[9)�����s���G�En��3��2(�	YڿO*�B�E�yu�#�d����2�i����Z6�M'��@%�%�?�%��������Y�ٗ8.VJ(�Ӣ��<�F�
�;�eP<����1���-<�������K�oމ��^�v+Ɛ�y����>և��W{JX�e��������<>AJ�"B����ls�+Я���]���<]4�l�3|�I�A�ᇅS�c��`Z��?���0�<�c5�	*��W��[Hr���f]4�^��!e�?�Gmݤw�;Q&�7���}]G�e�'K</�L�#��ƘG��������j�/vG�͝��z��"^ڕ�7�C���(�ʢefr��z�(���?KI)(I�����}5�ۄz���F�S�xl�$_`����+瞒�jA�*�?�jAm4�)�cT�N�[K*��JU�c 5Ŕ
̭����?�;���j��V�ה���ui�Ʊ�]���VI�q~�	�tm�����G�Hi�i�m���	DQzc�k���S_R��/Q3Oh.1n&���vq>����������:��#p�2V��n�����h�L��n~M�LZ���Ӆ��Ġ���q�e\�{� f����؅���V���ۭ�+������=�B�T��~�Y��h=_Q�$��m:>d�;&�Բ��Iԗ��f�>�W�������o�c���*y�Ȱ��|g�Ƶ@ƈ��;\���L�(����,=�C0�1�����p1ڒ�B��h.Q��Kd�7f�М[�=ʪ�l���j��p����ر	pa�|�K���V��N%kӪ74��9�x �{���6Ɓ�z<������ܺ;xs>Ѱ��^$t��~|H�Nt�~W��5)�&si������# �x6�vv�����o���u���v�gk�';�(b�-bj]����������#�XoK���� �+����='d�3��Ff4�|�r�ml�cB����vj�6Ű-��T�6�<5��6:59��ߏJ�W��e}��)>c?x��6$� �� D�7,S�j|�� ��Z����JS���}��kϴ�^��P�1�rl`�?В?S�.
-�(L�%���Y#
[��k�����O���G6jx�S�en���kk����Tt���G�ǧx�1��%(�M5]�Al�<�p�iP\ d�����E�ñ�T#y�H���L6g� �w9��a�2 DEa>t���Ѩ;��{$�n�'N/�F��B��a�#7G���X�)6�fZe;��V"��[;˓��>Mo�9N�,_���:����j-'={DzsQ������2��z�g���-]B��%q%A�~r��Q%�����ζ�"	#8�ҍ�R%୽0(��%����h�]�v�͆����b�μ~ρ@E��\��;���R��%��󫋂tS�}�u�O�\ԙUU�ʩ̮0��Ȗ��Cg����X(]�R��,k5�eC���R��ڂf�h!&�m��dN��g0L�H�&#-e�DF�gؾ�'34��^k�I&B O���CjQ|l7�z&�ㄸԚ�S��
Ρ��,�}I�vR������>1\���E��T�ƥ4���VJ�/�'����yW؆Ų��)�%lߐ����m�c��t�Z
2'W{l���`?���]G[c�Eb�犍R�a��ǉ���w��[�bq�`Ў���ߓqY����h��h~D�j��:�=\Q�������-�&�wH�.1���Y�ʦ�#�SXuP��ύ{,Q�T� ��2�H<�\Îq8p9(��v�G��x��W�Dh �����T�r2Z�jn�@M��q���R]k�]ޗxݝ�&כ$�J}'W(�E�%����1 �	[�X�/M��X�=~qϕ�������	��JĴ�n�@�h�l^�&Yd^S�7�Uw׬�������e4�~3꼈b4���с��E�4�ܿ]L�̡f|�N-#�ܝ�M�<��|X�Ko�z�͞A1��=�=��S�U(~Z��W�Rƪ��1�5���;#q�q]��`�Q����3�>�.��bPW�x��Չ�ZU�-��e�W�z��U�G�A���H��a!�}�@Y+]�8���Z�N����R�!�Yy�1����J,atDU���@��#�����?�����H(}�}� 1sb<׆��ԙ�Q�͝*�wC{��MS|�3ߦ dN&��u����f�Pf|�\ߔ5ڈ�;yGD��8��.��+ِ��:)���SL�ED�� ��^�0��2�;*�����3M 4B����ޓJF��5�Y}�|iY��<�x�T5����⣷'��*�1���p������l	�S�y��5���A�L,���a���.	t��^�H����_��U�b�ߣ�z�'�AY�j�z�PS5��M���aAeɽ�@@�xq{л�C~�C�
6w�A�!v�dp =�j���}�W�u`q�#zxQ�hhT���Fd���oV���=����,�#�����ߘ����9b��!%[���v���@��4^%;�.��y��e�n�̤ab9����g��8�f�z(i'Z�C�Di�yA٪�0}:B؄��*��)<�6k��D�5�+
t��Q�v�9ۍx_>y�
�x��h�\%�6�߀E��'�	Ŀ�n^����`3��;qfW���zWwt��f3\�z�-8�,}��sߺ>w����]ԢK�J>���X_�G�$ �S��c_���+Yd�U�Gq/x��j&#&tZ�n��p�� ��%�=ߓN��l)KP��1ħ(�|7fg	f2xWE��u�XR(Q��w��6��%�����^h	U	)	f�:ǋ��X���ޯ��9���^�F��c�jD��q~�RL���(���n ӌ�tI#�5VM�B�/X?W�*�ڨ}X���/���9͠k���C��T&~B1m��8 4�t��)"�gg����ҏ� ��&�by���lN�K��~�!��@x�TM�D��i{ǀ��6ɮ%�1�X��^�1#�T%{�M�:Ȯ�a��j��UX�	)�T8$4u9Os�S��dI��J�"����k������9��9��rHX�u�����9˰�/��4m*,�o��Ji�����|��4:��d����-��U*#M�b�&O����x�����Eu9���_m����=�7	�"����>iN�:�U	�*�g�& 0)�G�"Q�f�O:S���8��	7̺/��"'0����A_Cc`C~�D8���,jA�B6bE�]��n|�����(S�$�(fSg�(���-�1����`.�"��L��\sbw��^��0���eha�R?h�H왏�8dk�n�����$ƫ���y�j�Q��V\cC�M�Ї�M��J9Ws-�ȴ�t�Q�;�#?]x����{�<:�I��8�|�~yI�8[1����47�@�l�~Ԝ�;�V��"����XTLG�n������?j��QJ"Z
�0p�z�m�#�)���qO�~
E�
ݪ��ؼ�8α1�/|#Z_��_֮N����^Oa��n����T�h���S�Z8Tz��� �Q{'�&)��&�^x����E�z�?w%��-$���?��i��c�dqG�G�����n]R��i�J�O˼i-�T���_��J	�c�NN>�Ρ����VOʆ�[� x�jD��.Cd��î���ܮ�\)Z ��z��M	��,{�������{<H҄�+`Pc�+i�(�F�0D�����{=�?vA���BZr��V]Y5�;H%��s�[*��bQP������æa�_+�W�(V���X����Q~��&�d
�W����\�z�2";I�XX_�@�0��zHkV�-�*흥���Y���9�G_Bĵ��A��7����΃��tn͋��]&�,��l���A4����9-#�_<��;�l�����ȉ�'E|�>$�	��t��W�~�U���GX��Svuf�}���N|��u��s"�=�m�o�L��m�ʑ�ܹD���AWX,_��Ĵ�o}D�|U����+|l��e�̘5I�ɮ�o=+���q�q�Tb-P�`�.�Eq��1��Wgp��e���aX�AhE0p�F����D��!e^�	��*�#،�����{d--NJ����>��f _�l3Lȯ���6X  ���~e� �@J����0���[�W��F�Y\-�}��8��)���/�k����oE;�%⨃�xɔS������k���-Z��ZIW��G`���B���{�e��S.M>ޠ^/�=-3ǒ �M A]a\}��C�<B�e0�|�o�V&gv%U�4bc�S&�!�>��(|H�L�فԹ;V�\>��?���+*�2����EaB����%͝�S��z�d&��W��(�#l ���?�\h*�]�u��,��_"��|�=i�z�{�4=Q��p�J�2goT�{�Ǹ@<����P%l]i��'������*�F�0&�P�M��=�R[h�����2F�>����T@�If5�ܙ�і�B��CoT� b;�v��S`�}]��;�M.mH?_��,|����#�����K���H('���VJ��/��G����l�U<;K��H}�B��ze��%Tn1��$���� �)z���bJ��F:V9�<��>=a;�/�y�]֔ӭ���?��ߒ�?6�)�߆��l���S�,d������0*�!�T3��I�P�k��?��~��UP1�N���\|�f�v�N>\ߦJ�e��4���hh�������,*�v!�z���б?H*�UÓM�;1����'��#�N����"���-�d��)�<~�t��������pW�������sM��Z��mm�0�G[�o� զ�9F�	&�W!�#�u����*��$w�Ȣ�z6_���"�,���-���-5F��T,���J�eJTX"�$[bOyȬO�gh{��"%����)�ћ�D�k��PC�J���M	.�|����}c��~��\���u�<<PK���'�.kon�YNx�E�MOF3�����@�yVM�N�W.#+4���*a��6���i��K�1��<ޒ�Zs��'��"w�
V3a^��HI[Μ&C[����T3;�)VX�H&�R�POr�Z��$T&����cɞG:�+R0tĬ����� #5�3���#��3{�̸��>W�A,Ƶ�2Q�q2w3єk���&���7���=��/���M���B̨r,��7���g�LNȆ�#S��GR��g:2a��nrPYS�*6�_m�9$U!��� 8�w����6�A�w��n'}��>7��m�o0��p�U�G���]�k<B��8�w�~SO��)�aϑ�1�&uL`TM!c�Sh��kN��3���^�ie|��	���E%�c=Jr ����[�H�|l�(���L�0m�S<ci�Tp�،n�5�D �f�Bn��#��Ӡx�}�Wjd`F��rwQ�Q
Ψ���&N����tJ����y�����c�/N�ӑz�����R���0V�����oI�e�ʹ�7;����8��G�/=�A����������L�Ͳ3.�Y$�B��h�������i��4��4T�vh���g1�>�q8?��`�&��9��Vg�!��?����zPB=IJm3�d��DҜ�U0]Mg�M�e��x��vL���21S% ��VX��t;�����r�����v��k��C�Bx/���',������u����� ҝ�0���CK����W�e��x�&���s��*��#r/�6�Z]0��:���*����#|��kף�A�h�Q���JB\|ԯDގ5N�p�v�p�|�ĭrd�D �i�%D*��f9��'Ų�c��d10~7�(5���=Oۢ�A�����ȅ�%��~�����i5Lڿ�z��}��A3�'�~�7�p��`C������Sa�gIzb�δ�.�՝�E����b�%���O�<|�q]?O���k�g�������2~7Dt�qe!���t�L ���A'���y�(`��"��Dg�;Q��~�i�y
����}�J\�NGv�4�hsC�o�5[ÁY��<b�Y�hp�����^�qa�`����ʹ�U���8�(W��M�/咷?2�~d���JRWZx~�c���w��;�|�HG�p�FEY�'�H���ԩ��G����`C���4�v�gI<h�GF�夔?�y�>�a�`�M�^5����l�KVL��o]�V� �_&��w�,D9 �-�H�n�J�9] (�����Kh���T�U��A�C��H������W����U����<z�?yb�'
rZE�Ź�^����fi��f��YH�0��Ҝ�q";rf����]y��If[�]A���Cx�R5F�*��M[�����z����t�Vi"�4Qd!�H]�_��"�����JO���0R�-ľ@����5MI��m�>���e���b���d��ud+~��.]e� N9B��Ww,�f��7:��pr(�=�հU�YU�Q�ھ������ܩ� 3��#����kלC�.n,û߬��_N���Gv����c Z��Խ���wA""�d�����(��v�; =�9S�E��S~���sa����P-�OQ]^t�.2���q���- w�ٓ�H��J�BU��W��+G�ލ F�&4�2�xd�(�۬�l���?Zǡ�'�s7��]���ׅ\�O�\F��)%���������H�V�q��B�8#KUl5��VnYh����p���l�ꖤ�����z��3����W��Y߽n�~׷7���LD&����;рXL5M�����A�v�Ϥ���̡.o���l�e>D����C\�Ÿ�t�`Ɛ������	i�a[��A?���҅����sѾZ{��?�_�X��2i�����]n�������Ǿ��p��x���������և�Hq��%�1��w�
�K��x�2oTR�G�`I^U�=b�7d����|�N��9� �j�A�s��Iߴ}�'�(�����)@f��W �$��f|�S�,��>b�ZZ���=s8;���ꑂ���(�Sӳ�k��h�5#�e�9�A�޶��8犧�����	�.�a��Bh�i{9���K�xG�M�/�������¨%��6 z8�|t�P�[�"5k��q�+��G��p{�"n��0�<�:�G-}6�������g�gFNWV�����} �b�Bf%ړ8�����J4�y���_ܳ�	ݙ��S��!�:�����\\e�4d�5�7ho��۞ �ynu99ţ p���ӢO-���hu��t��@O������LxZ����WF[8�ʫ����J�qz���+	��s��[U)�E��E���k:F�!���:�ag |M'h� �W�K=�ʙ�K�g�u���K�$��7�j���p����D�~� �����H5�l����и� �̟t�2@��1� ���eg�j�n��&�@��4Vl���U�����?~5�9����I"�o��������@���w���)oE����W�D�a#pr�����p�'�9vt�у�Ѝ"����8�*3� iz��R\�;8���c�i��ζ���c�M��Q}�mjڴđ�qD�:�Qqm�?Ӫ�����(�j+T,r|F� �G����p��{�ٽpI�����O��-�ӟ�\0iO�$5���d�`'+��VLLL������`�s���U!�j���-A>�Rf֭��܊��L�R��3:L~����ꁋ�����Z兇m��ʍ�?*�!���͟UZr,z ��ģ��Eqڙq����3�t�� �f!X���C>h&��o�/�I�>i*+��l�K��lm7S�6�E3Z���ڗ��N�z#��A��߿���9�yf��*�>����BÝ	�VF��h#�I��D��q������b�'-4��,�yU��;�E̋q�X銱VZ��\{��̷Q��E�i���p�?��Na��Z#>�i��{�@�B��w'�v�1��׺�f���Fm���Ҡ�Q�)UJ}���mv�<6�tsQ��s�Γ(�9V���eZL�!R�.o�k
!.T��S��wf^�f�
�Z[_�BEU�|ʞ~:3�n��g2]�$�9}�l2q��ʲ�Sإ��6C�{��?�l�I������&qx��?�I�Us�Vt�(�|���O������x���rԻM+QԤ�q���_Ź�_I�S6~�G}�;��,iz86g��h�
���;w�PA��Zt�tJ6��c���#�_�#C��HpnʼMP�U̽ߖw֦BS��Þ����MD���t�wz�2t����QZ�u
�;�X3*pL��[O����v���M6(TS�#KV&@N; ��E��Zw�1aT���왏������;P8r(T�F}�3��,�u�7�J-��tlr�!����4ƽ��)��8���k�?1�]O��k�)�8P ��Wx�f`	v((46H���Ǩ~�0�:�'���M���S6B�����ނ�u�\��_�_��8�����y��I�q���I"���o)��[#�\>6���ËhLh��d�[_O��2���H> ����o�9�rZz��q��E;������}����g��O9�a���	������j�Q9�x����\��0g�`��D���|��d�E|�>H^ɛ�:%��މ�o��G숍:(�ڇr"@/�2�/C��gxxB�-��C|��8&`�d����Y����_��t�@.s�}5bbŊ0`*huq�CW8{���_�R_ULO �I��?e5��Sp?�0��|?,����)��Z�L�/����a	T���}�%%Zj�� ��������=�����y'J�H|W�cP��ڀE�E��6WczS�� �
�q��խ�%3�?c��N��c��Ěo����P����6�+�͘�9�|�S�~H�cG[8�5�eUX������?1��7ii��gt�>��,l����&m�@�g�s��N���a^�p���g����.m�J_=���zҌGi幈����ln0uڳ�7�J�#p7�#�$?����'�qX-c�N�� �L�U~]���r3
וk�R�`� f���F4�~�xm��7�=Q��Jr.�Ja #���L���M���~��@�Ұz�o1��7�v ��8��5[�vex1�gk���q�mP�tJ�Z��v%��h<|#�[w`�p�`����q\#������!c�*������İ>�#~������e�aAl���x^�0��˂^�$j�]/�ѳ��Vg
��C�A��xT��J�w������ߑ�Z<j���l��d�O�b�I�s��)f89���k��"Lz�Y؉݊d�-	���3����N[Q�\�$k�6�e��~��i�tN��O��_v��A@C��<�c��weɑ���Y�2�>sF3ݢ]����t��Ȟ��V�ԝ�9����?Їm�%��Vw�ǻ�Dν�*~�b��*�c,7Pd��>hj3�����Wg��_�Z��n�iӮ^G�h�54C�/+IB_eC�h+�^D%(��>�n�6!n7�<>7ɡ��9c�B�lQi��Xy��h�q[��E���;^\(	iC勔��DY�x���;��3Aj<P
�|���B��� �8U�A��5ܣ�?kC��e,jd�����p���"�^p4i�R����f;&��3c���v�Q�	A�0�����?�-�?)ˣzPG�q��1|�v������o���y>��.���L}���\U��E�Z���jӪϫ�n3 X�.�A����qg�fm�o7��:qQ���^�2md�=�/�>� ^���nac�l�_�a\M�$��~�����.	ٲG�]��[r�#�b�����17�c�1�x��Waۨ+g�EY�x뼃�W�%g*����B��-|�b����9׎�����g�U0�2��(���=��v�+B�HԬrbs�o��~���?
A�I��U��.�g\���������E�/��愼�0��"����pǶ��(����-�FIQ5�M��M`mJ��t�!���4H��V�JCY�ne���־��z~�E5�[?�渏@/5~�S8I� #�9����z@�^�C��U�0v�k3)�E�LK1�G=�3��H�i|J6����^�Dj�9 ��s�G�B��3i�p��1��OWDH�5m����4�Yj�>b�$NC�}�;C~��j�9���\�����~i,һ�����s.�ڨ鍂��g(��\��AR,;Lqr�B}>S���F�Jʺt�r��-L�(m3���N�J��x��B�]��MES�9PhZ�u(���pY5��;�U�����C=�
Ÿ0]9��S7\�J#�ٛ���a�Xkx��}��>�y�q��@�n@��ʕĴ&��+@1T�+�p�{�&Dj5�I��C;'�{$�:Q����F$3�ȟ�x�c��륃�W�m�c�lL+�;±����`ǣ1ea�L��W��n��L�Fm����;�*�a"�V���y	]	
_^ �
�
~k'J\ Ln�d8��9�S )ُq3����ri�@��I�
�VB��u˗��d��2�`��Wf'zwJ��<��~w�(�/$F���܎���U)���]Zy����G�T�:��<��:b�M�Y
R+�+rQ��I	<���b�4u�'��<�vH؛��ABO��L�+�@�Yp����k|��0�9�A�3M��� �v�xδK̆(���a�oא�����k�}fr{~�G�
�ڸ��l ��e.�K���9�}Β�� ������x�I����"�Գ�+%?���dmg.��"��7׫�đE=�\�{ �A]�z�!��7 ���ਖ਼ (�:θk#�U\ӓ/oe5ێ�E�-�R꧎`�0{��9@�ox�{#U?���g�B<ٻLd r�W��r��Dc���=�0|��"E�q�,$���zc��-:�/�X��k��M��s��Ȣ�JI~h`"���E�����������N��e�1v]�u1��"38��FSv {-��1B�W7��lE��6@Hw��U	���\.Z���c?T���1�!}Hw�>h���!Ѕ��2��C9�iZA`A9[Z뙢���3f�4J��LKv���Ujd@k46��7��x�A��t�Z]!.u^�j�I�B�z��_4�M�k��o�C� |'����*ُI��6��-�?ܬԈc�Se���c���5�C��<a
�>�Z�r4'����zAE�o���q!Ed��2��륣��O����2�_�<�T�j�'DA��_�|@��fW�"��"T:^����Eg�N��q����oj�����:x�k��������P�f+���pQ�}����4��r=��ț�E(��Z����B�����~�|�����2Ӻ�eP;��GYBF��w�<��d�H�$
��h;p���n;�>I��ёs�r�7/a`�i�R�+� _:�;s;�)Ӌ������ r�\�F���:w�.~���g�s��ik�ؗ*����I�N\�V���/��}��=X �c�p����ܦ�j�d}1=����K���ҳ�4v�q7h�(�g�FX]5q>CKC�����Z�CT�r���?�Olnj�n�_.Iy�襫 %U���ʫ����m��~1e?{ �w*�����77�����[�`cN�S4�L�MΪB����c�������*d�(_���1z�o|�[^�3~�a!�j�څ��J��kǳv�pNvkHG�S���,�y���}4��8�눞�W���X���t$���y3�h�K|7�͟o �?qS;e�u�0�>{2g|X�G)'���W� B�8XuWD�k"E]�)���rr��>q#�-��enC��@�k҅����p�w�CW�𛇾ѱ�EÍW(��]�!�F+)���B�auP�^����O�ӒzH�13�Q�����V�y���M<iy@��z��]�e𑦃��-p�4I���>�����-k�RA*���Ƣ[ù�m�uA����_u���r�*�tgs��EQZ��\m��� φf�(����z'6�E�`O꣭-?[�6aK��`�9�6%<�ΠJ����^ n�و_ʣ~l1�:Sp�*SKK� R%P�V�ҊQ�����[�Tp{�N��V�K$��d�.n��_�����ϪZ\��ѥ���edr���E��߱�Aرq�LMN'�8:�x%�j��i[����uyþb/e��!Q*0kIo��{���GOC{�l��ߴ���lj��!Z��3�K ��e:<�ߞ2�_R�������8:����s�V�,�ERw������ ���i2)�!�ܾ׬�/Sl��)f����4�s(��(;����<��y�wj9�� �6u��9EB� �sJ���C���O�/dIA�D� q���v��2'9
_�ꊗ[vd��j͡�Ȱb�]�_�U�!��*-{)����k��(UBjDs��"�#��r�؃O�N�Ļ��Y���`�O���M��2�A��YtY9>sJ@X�{�㗒�x���~�OT��;>^£0�h��QW��0�o�`��}��{�D��t/�|�8� l�T�N���"�L�Mf�58�Ŵ�k�M�T0vhuz�Ʀ�ە"�>����=Ь�|a
 �*�Q�T��lS��@B�N��;�'3G'��1���N
	%�����g�܏Z[���[��7�Χ��#��b����(�h�S��-�D/�5�X� ��DS�<�_�G�e�/�	�:K��++=�Ԁ���8�Ҹ%���e���|�۷[�]���-�1g���
wNV��X�^I���~��G\5�A���_��y� "=�+�6l�b[ >U�7F�����ߑ��H�$[[4�����N�� ��X݌��py��	.�߻�r-�l2�d�ғ��i`1v�\?�`��d#Jt�����%�oǜ9�%�cމ-s�<���h�2Ry����b;����6�V����.6��E)�X�璷Lm������`E��,�+��Y��S�
%���[HF�ē��-V�����x���8�Ts����5��o0�n�0$��4ӻ�3B��Q]�H�Fx]��!>v�F�j��Z��hzD�d���3����v�;쀞r�8�,��/�_�&Z����1� A3��xc��㠝����T4��K6�A{����@�d�o�~|��?�I���Ʃ�+���8K�S�܂��r�pK�g�ו%8�IZ2���q<�1�S^�� ����$����\X.ロG.��kaHfE��-��&��YFiz��;��)�Hd\�V�C<��p��bK
q���beD�<U���NNkX�6�3\�~4�$8�L���c۔+��gO�;5��KO+��0G(���!�Gp�� Zc)2�d���d(��3�j1����iT8��k�3��i�\�qc����Yԇ�n��W�+����?J�� �{��m��YĻ����[C��Y�Ỷ�~y����ڨi���R��U�.��,|ҙī�/�~�1�O
QH˟�%{�m��e��u�N	�Î:���TT��Ճ�a{�}8�*�v{w�E� ��]�[�C�_s�,ʉh��I\��ð<�_awT&��������F�Ӊ�*\��L@�l�{��^4�q�Z=eo�o��?	\w��>ϗN�`G�L̍�"eB�����"�M	>h��~^]��PI�J�%�n���3��e�넦We ~¿���aPi<�7�\3��w9`K�۳嚰���s�q]��#�/;�N�'�!+~�u��T�������:�Vl�F�o+��x�����o��f��;Y��f*��Zڊ��9��r�>��m��Ga՘@U��8��"���BR����'jKJ�ɯ'8|�5����y|���*U/\�q3?�kRbK0����
*N�P�	�B�X"JL�����Β��/�DF!�"��gyAn�@	�����nfn���n�_���Vo����d�U�����E���^;��R�x� FkYq`KWw��*A�
�9�E�x}�m�!�Ex�GZ����͆���0���`�t��S:���߁swN+.�<Ҫ"�>���|���q\�g�M:�i
���<5EڙR�]PL� ����ʊ��`pT�\F���yz�?���^��>��<Ǝ+qY4���V�p��*�QG>�YX�K|��W����m�ɺ��"P���uf����=k)�]oB�D����j�+a���w��-�b$�J��������H�YN�!ڎ>X9F�0¥�)��C�ֱ%� Pq�/֖3��+�G�.�~z�����������p�Kt�~�߈���S��ۇ��VP�C�((\��o��|��׈?w*u��ߴ>h_�
�=���
c�X��rt���kVB��rE����C�q�|7�������?1x)a�+O�8O�����fe����O;&�~Aq^�U�����E�Ň�6B�H�D��c���c�2�d[�僽��kD��~��d�G{�^4��=�B^Gi�C�E��?/!b��)���/
���!ۜ&�<��pe��[YWyB�o�c��mnQ�oHG�Zm�/:�� �$�Ţ��I¿SHW��	��Uqn�.���ʂK��ec��S����Ȅ�zuI�QDG������QX�g�|�Y�j��}�zI5qd1�@c��{ry��b����mR-{�B���aa5���Xl�z��P�|z�wO�>
����;J��ƕ�@�H��(/�=Yv��p�-c�h>.�!�����Sm�\��2�Q'_��@٨H��T���N8ˢ~�V�?�-[6x��&���/� �0SLTL�Ҳ����L���ϥ�{f��c�|c�ߵ�^I?���u������ԇ{[L���5?7
�U��]�
��U����v��\M�D,��~�Pw���{Ƈ���Ǵ]��U��˖qQh'��ǩ��e={��,���u�:�f�h�;}y̎�}z�~��;��v)9Q''{��ˀ"�9/,����N��ĕ^2X�֫��1��b��פ_��%t�#����]����$@tA�]�pC\>�([���	�l�&mpfX�~�H�g�&��!�NU����eƢ����֜2Ky$�x,~�BW���}cwbfb�7�#8M�*=1cLrh�COѤ�X��·Ot���\A�2N����´�����L�Hb�* u�>��X�$�m�wc*���O�}@�����m@!�����~)�_�鉖���KL#����_����(�Ȳ�i������b�T^���/D�7Y?�6���r�o��>�g�}�>�B���ڡls0��g/��t�D#Xi�כ�_��`�LlitB��!a��_Ǡ
i�<��
��9���d3u����K��o��!�)y�I���	�hrF �H����j���J�\�m��i�E�z�ױ��ӈ����R�����l�����LS�8��uP8:Q�ϰ�M�H>�	1(���\�j@���f��36#�/��D&g����8?�{���:-���݋�7�~�j�/?DC���;�ً3a�wA4a�ի���v<^����l�EjGV,{h�D�|We��>�����k��՜��_�_M�9��O�xC���2?�ōFmd�kw��=�q6���.��V�=���U�5S���4Vo%`�q�Y��
l��P7oS y�͒�����oFc����B�J.���&�5��N�J�O�3hP���Oh9���k>_�Q�`�>A�f��Znm�����}`K#l�]zq�E�|���5\M�1�½�Y3�=��l��kE#��9��̡Q���`�+ܬ��	Ί��������Y����>f���Lg�.Y �i��_���d�sb�� '"���y����(�����56��ay��S���=���hMk~���rԶ���g��$�?�v��,�U�ܠ��Π�"�t�wsb�:Y]Ly�i13<�Cx646D�[��P�:f��r�F�:a���6�h�9�����7�=x�X����>?v6f2�+��Q���t���U�^�50�"�5�A�V��0<]��i��\v�`�5��U���8�M?�F0ǀTj�Ŋ#v�۸E�����%�_��_L��A�p^z�-��T�A+�w�:@�M�'wo���F�c�BM��ht�05`�[ �������J:�A�O�$����\r�7�:����Eŵ�� n�D��Ph��+6	[����Gբ�r�iڗj ��mx?���� U������.����5�<�11694v�$ ,
����W�NǞҖ.(�E�&�D/������T�:�kC�^��5m��E�9�5�xˍ/v	����!L{�Gd׍�yڛ�z����]C���^S��&�Y�� q�\~����0��p�\1�Q�Q�l�8��U��.lRyJ`��H��s�1ȸ��-pԡ�a��<�@}�W5セM�Rkv�%�����?��^���Da@}2�4��xR��Ͷ3�	j��[  ��D�x�
��IY��
�	V��~�(���������Nb�{(���[�Y�ZO �Iz���cT9
ؕ�����m�ֈ�����$eq��A�
�z��]H?����&�����)������ �cN��"��� V�)7˹M7�@��ԜqT"�;�T��v/�n��LC��r$��	5�v�7�Tr�2�`OL�ڟbHQ�(�WR�P��
��f�cѰ���$i�7ǝ��	�@�Urו����jA��Ψ¡���+4�����.�%j�ߛ0�]���^���c�LB��b3�p}�"�`�t�)�hf�/�� �c�P��XP8 ���x�Q�,�!s����))PWyM���;o���>R/���ւr���}C��IS}��]
�4q�ۖvc�}�μe=�`u6��{ �{z�В�Y��UqC��DǑ����Fa��Mk1_͆l�����b#��o�Qؕ��q�t��.C0 ��Ɖkɾ�<�
mY�
o���V�F��\�VY�L^@t��l����N��*����J����/c��#�O�,��� ��7��Xv�k�*��ݰ�h�nf�F~#J>Ŭo&���P2B�)C	���D8f�DȈ�!��nΛY�_�|���v^B�K�oFq���u7��Pf�YD����&�I=��e>�xiM�^���2 ��^��hO]�3���?��e��-�+��m�����6O3�e�)��s����h�;��no�/��K11�
Lǋ��W����T�����.��hU�E��Ul	��PC�D�g����8�i�
,Ƿ!i��\!1�;���]r^λۢs	�hB"������P���L��R�U"��Bt\�����@�T~�������8u�w�,M�3���a��6(��1����k�.��Ңe�,�����+�|��:9���-¤����GWaɡP�x�3�^�%Ȏ�_[�kvk�٭g�LE0Q�H��;�y���C��-x���;�iֽ��A4���s����Э��E-����ᮙG���s^��Z�'�:E4��#��mJ�BO�́�5mhOU
��orۍ.�U{��s���k�=�{�}��Sr�J���m2���u}Ƣ=/��)d�KA�]tIBN��in����}w�k���zJ�%�D"C�����.�W-�_0j	uـ�m;���}�q7c��	\ %����/��Ȼ�;ƘL�O)�2m;��y�T�⷇�j�u�X��Ѥ�~��$ʃ��u^������ ;lc۶A��(��]�+%��U���F�̘�ŁS;ځH�ι'�/b⥬D·�>l�v�|ꘜ�PUbV�>	B#	՞&f��.��>~*bLZ��L�c�`}LV��>s��B.�h@�9R`�g��>��=�F�:m��H5e���BV�d��A?Y5 ��X��fܘ^��	����)����޵��|�j�]��-�������,Z�|K!��s��!�=xS�D �A��a�=�j���+��G6/�3�,ě��^�9.6��M�YVhgbzȀ8	����,1�i�^nʲ��r��$ܻnt�.�k�aL�o�U���ؑg�~�vtI�	�G,?w;��7_����� W�:��n-�鶜k>!�2�m�����mTvR�?�D)27u�|�J�m!0�:�c=�]�ȹS4��.��%�/�b�I��f�P8j(3Yo$��8����L�����s��}JJ���
��%��Zq����(�s�x�ta0�,����A]7oH�������kݴ�b�뚐�f�xƅ�7b_`	��,�I���	o�1#գ;�ƪ!ҫT�H����Ɋ�&�脻B�L%�/
^�P������lNRP�%�l��`&����-�p��`��ma鐋\d��b]��J���P���H�W[���rM؆���n��͠=[I��6����wx�Ag�J���4p�>CD^7H#�+������Z����+؀��a�q��<I�o b�nę1n7!!��٨�Э%��3YS�R���q�	<	��i��Ԡ4��>v噧)P�����=6�u0RG����{��y�P`�'Ywx*�#�mw�X-����D�h���O���
U���Qs�i =�s��O�#�l:��`e��ğ����S
�z CO��_K?փf�k����O�5-]&��9� (�u��՘ö��2J�;�Q;�/0KQ�%$MI��K�����
��q?Ff���9U�/����O$ 3"���>��NqF��2�ixl�
41����[�j-	�
�ꆅ�����^0~U+���a{@�.~���^���b&3��hxY��-�$5�������+�u�i~��T���?e�il�MR����gO��p�@��!l��*��̸ᶩ�LD��@�I	�f%�dx���SG(�s���b��1*�����'���"���e�娵�����,���$m�c��T�n�|t��d��?��ū�w�ѻnXHc�x��li%��጑뽉-���0��3�!�:"`T ��n�7� ���-��M�˼������N��I�@�I�5���I;�[�vVs)�CG���{$gǰ|=��Ԭ�v��z}TW��e���͢�?�f���C�JY�n�NE
e�N�[��UJ��*z����X�o���?�V�]km]��~sT�,�B��P71h�A!)�<�����tbV�F������wF�._;�I'5��y]�>�$I�#��o&G
�c�f/s܅��t�CN�d�V#�������yO��/2����c�o��(�:8ʡ֫4�[�T�-̋�ǝ�v���Au_ ����^R=����puE����O\{���-"m�x�.^U��16��@�+��
}�V�T:��
x�5е��eo���K�Ť��Mc��n<���J
��G
�m"��>��B&6a�����4%�aX{�p#P��Ԭ~i�=�\�t��
Fo{��ג�ɘ��i�b�Nر��<�I���4!��w���5��9���S;����cbb�A�P`g.C�n��� �b�=��t�� ���-�Hc�R-�z�:�g?坳���q���E��T��DM�nL$������
`�3 I��''O�@ �3m���	*������=�U�T���+$$��ॽ�]��
�=��:Y���Iu�P��6Ge�&&n�vj�}��5�84D���T�p*V�2���I������r��k~W6�����￟��D:�r�3q	�s{�N�2U	��#��������"i�7>m~I4Z����n�'^��9�,�D����
@�Z���bD�"A����mWj9�i�~�I6��7ƿ�;����퉮�� X�:ئ�A߱���UEJ�x�di�P�������O;�Vx��z�o�C��n�T|P��ӿz#�Ryp���P/P��\kk{dcJ�B�L~��nR��S0���8��0s4\֜������"��JL6'�u�.�3t9�;06��yL��le���*��~x���D:�_����9.��.`��\���a�.7 ���Fx��lTA<fɓV.������ߔ�5K��.Yo-7�d8m�#�`�l����d��͝�'�M>:���dڐ|h&����7[�w�L�OE@C�d��_��'��
>U����~n��<l:͇�K�ɳ-Y`jq.�I�z>��]g�`_�a������)�L�׵łmF1󘚊��i8�!B2Z��B�a��"��y����SrA�J��29z�~��I3�|�PA� ��=<�����>_�~޸�m��W�s8��0�<�J
]�3�@:�^�%s]���0���$ � ^�W�HoS�)RF�l�UC`���U+��XCA�?E~�"科��m0��X�qu��f�7W�T���U�����my�}��!��Ѿ�|L0 �c�Wz�JM�9�V�%H	S����D;Au�ck-�_���9��@��Q��K	l���K�|g�[ιwx�"�"]�l9s��e�B����
i_cvg����V�m#�Yś͂������Ҝ�d �t��{g�ɤ�P�a��a���������_�F Z����BC��~c=Ǵ��C�/+)?�g+cS�X��tPI�||{�y��-"R&���Ֆ�:�lH��@��!�><�9@�5�0�d�Tډ��Dg?�^X�<���������B���b�5��ɊF��G$<S_m�4g�(������WC�Aή9����^"��')��I�w)_u�����w���~�3+�ִLY��(�"���������eG��9����L��t�E2x�3�ɐ��uT=�_"�\���i�o�����u�({LOQ�8��	�u�(��~����
ƫ�ݙ@,�??h�Dhcɑ2�c�y�.i��M�{+��/�eE�bZޅ�Q���_���m}�u�L�AǕ���q��p���~����;_:ꍼ*�����z�i�����V���4Rz��袏���,�<��O�OE�̩�ֺ~��E�c��M��"�ĕS�r ��=�W(�H(�C��N�.7�%���o1��vu�(8䲳A���X 6C7ʛf�xX���Y��:�r.z���~�5�v�(c5Ϊ#?�Oe��8T��~��ɵ+�fQ�vѹ�C�9�P��7���	���E�����|�:Q�E�P�}0(�@����|�a�Y>���Ur<�P;Kb���wÍ��l�y�[4��k脪Gs*P�9,$�b�r��܎6w{�if���`̻)*�к�d�B���(��HN��:"h���B�O��� �79[~�}����p@��� f���wZ!�1Tc���ם���|�U���F\7�qr�������@&������Տݥ�'-&�om���9�s�D��%H���{P?�P��oܛ�+�>�E.,�őc�w�jOV���9T4&VK��rw�o�,���T��o8���J���MN̍�P�e�	���P���������g��R���ƥw���"�[iu\�L��*�hY�xy�s����G����?���D�G�:��?�����{��=4�n���������Æ�����dL]����;��Eڗf�1<1�$���C��ǘ���tWB�PZ��������R�ε�Xt{����G|S}���=�����P��V�]�6��	ř��y�e�s�#��
a�yh�� �|~�[%x�Ul�9�%f�K�j"��aUe�ְ��k&��,j���n��e��0ǁR&��h�3Z�e�iy�zxt�v���-�!�.?H��U�����uۀ���3t��Ơ�+�iO��}~3]���Q/��a�մ�y&�`_�O�Ն �%��T�&�JK��O���.�����l�0��*-s��R(J�߈a��0�TZ;h� �|��%D��!�9g��Yh���YT{���b�y�ԏ�׮�s5�?*�4 i.+�7���~����d���x��G)/T����oI�a��8�ͽ�ug����S� �BIbϘG�sd���'�ܼ�VE�����B�7�\'�E��m�i1 ���u�&L�#���kϟ!�pżL��{[4}s����}[}��b�͉4��b�!���Ĺ�� '�������D�XZ��爖L\l�'=�mn �=P<�Z�-�YJŐ	w�K�5?���)��>��tD	�,<p����4m�y�c�ӧh��4>A��ٛ7��^�O��c���h�hVPPeX��HX�BQ�L�m�N�|auf����VS?�)�G|E3������n�u C,!��5��	�x�j
�X�b��!�q܇���16������*��b�4|m��ITA���6�H˾�
�� =�[%����8�J��X(���'%�V,���iE֎�
�4�极���M��Ec��ǃ��0E��ҩ�H�pD�\����f(�����	{1u��_j���	{f>�{��b���o������t�v�@�V�(\��Ң6m�BhK����[��'R��z�)��f��;y^ ��3��gw�����l�.d{MhX��_�����_�4)_7C���+�XH|'�6;N͞����c^q��
L��Y����*����Y!)3��� �a�
�śܓ���f7��_?��ؿ������V��&����h_6`�fn�P�T�rjhV0K�FP��(�y��8H��;�_��� ϣϨ�gN�X���؞sv5����_U�h�HM��ٷu���D����ZJA
�>I�iy��ҙ���^�$k�;���M�d�k�ż���ny,"���d�����bWu"O"�D:;�F7ӫ\|؋L�!ɔZ�*CdE���n�j��4�w{��p�,���ex8���61���y��&¸�8�~��0��7�!�I+���n-c)Z֊�~
ՈJ[�df�Im�2C껟T(��_í��=��'TX! �[~�_v}	�ܷ�Sh����솦JXE0:j��3�d7�m��U�Y���_���ZI �B��G�\W��Bn�NO&�r�����G�q��5����P�Ƅ��i^�^�A�`+ŞҶI�m2.�s�U�k �(��ٵ���7� éꑜn����a�M�۟���ws�H�[�V>KvU�m�6����P&�I�VI�L=�w6=5��9��!N3D����	�~o��/U�w�Q�A���f_)�ycA���'_ۼ�Ƣ�ץ��������S�O�]i�@���������C���e�bs��L��J�A��>7��햹��t*������A��vU�����="���)�gp�Jj���:�H���C��+[i =�Ji�Spʝ�%����+AeMr�T �Gb�zN2(�y�����\��ʊӴU�VX�q]ڂQ������a��WBt�Fy��Nh|>��c���878��Bz��؆�F2�{=|��?ɭ��p�K`�曺�LL��^u�̔����s�q�~@�������\�dġ%I��`I"y�x��yG\X��c%����y$b\�bbn1*�=9Ѽ��@1qhi�P�޳q���odT�ޤY�Ժ�ӡ���m���//Y�k�����F�k-��=6]|f+���L��/�଩c���nū�>	�%�i3�.�=H���ٜװ�p�@.ڍѮ����t��>�iP$&ܾأ����֧��~��|ϺƋE%K�Ĉ�=�7u?��q��n
�
'�aо�T��0w�=M7�8���u'ڳ�џ����/�V���o2��+>�#|�<�{1�͹�fi~f�Č�rA�Ȩ�؊1l����8[����)+�@���\�n�\=����?`(�&X�h?�\� nd>����Kt�������P����l����;K�:��K{���.�4�N�5��"N )��jm&r�4�㸳�#,�� �YoK:غ9ư�	�	aٰx��kUC���v��߂w\�!�����K�n]P�e�/I�~=�׷�׉_�%cf�֌\!%׸��ʑ���C&��џ�Z�fS"�%Y3�_�b�1b4�����\t��Myv��h��a3�w�zЫ�,Zo�ﾀ4�����ǋ�}�%짴���L�%#���A:O��˔~��%D���U�K(I��H�Q�4�F��z-���",�A�Sm�����G���w��a�~���q;F �8�o.#u-�KPO��1T�f�mI]b,C(�6�@���_��j!�ГeXe�-��
����\VE2�T�'�m����� o�s�M�G�1��<nZ�X��Ĭ�,F4Y�:Q[_*q{{*�K%;���:�m0�!�� �=�OE�9��ښ��Q��UfpȚN;�����Z ����+$S�d|ã�i�O��%��?Ӫ�K��¶��o*tV����bu��U�ּ(�3�ރCϋ�������_g8�O�~�}��{�B.��O!���W�o�>͈1lB�^�qEl�����.Կ1�m�|�Xƨ=��4]�U�/��7�#�{��2��tJ���h���p��!�)uKi�lng�����`5Qu��C�eZ����wn���K�A	5	s�CKqv孺�1�^��kZ2�:�Gt+�)��u����&�
H�8~)�߻X�=���V�I gE��}ʂs��O6�u�J�LՇ�����s���$�9S�7�n5���b�7�;K� �-T�%"�X�*��i�'ءP��e.���;A!�ۇ��E��U�zC��hU]����f�G.���&��Ȑ��"5�H��� �ď�F�_�����V�޿h�a'ZC��I�fO�HZ�"\m^��^�Զ��*�T�'4D�p,^��# }ET,l]�MU��=����M�G:bcBJm���'mx�K&��q��uu�Y���k�vL}� #&r�4$R�Xp�4߱k	>>��P̀�WN���ؐ;20����íj�z`�DؙA-i$�@�O��\bdf���/�p��S��T���k϶.����|Fma!�6�飚�h���lh��\9�v���T<�D��)������r�7o�bz]��� �.�qZH�+�ܵ������1F�>#�?�G�x�@�PK�\adP#$��oY}e�ȋa�	�qk3�<�A��Y�x��G�Ǻ�Y�`f�Wܥ*�(YT	!I��Cow�o@Z�0��{�n`�kC��k��L�uv��������Շg��_>�@/w��l%��2�G�O�M4���@��(������z&�F���֪h+E|v�ь��C������?�pTo�&u�v ��I�P�p�#����L,��1_�99���j�w��B�a߯��N�7S�������`R5߭�g-b�aJ�ߺ������K�t���Y�p�-��m瞃�j�Gwx���/���RʎK������A��C���N@u����f�f���L��lDh��%4�]����:��+�g���b�e��.	���/� &Hc��7��~.��ե-[`�T�ݍi�uh�t�-ZLen���8qQ��~r�W)�qML���򏚘y����3c~aigY�o4X��f���+�Ll�����"�!Qd��8�ړ��2��7��7���]�׵�(�K}Q5�4JTޡ��w�����s�=��H;�D��J*l0��M� �C�ӽ��Ul;�n���al��)�������Qа���2��̋���H�� �������{��s�?lcS�1��Xx�����)�|	�s$�D�ծY�0#�Ax��ޕ$���ώ�f�}>�}����U���7�>lm�� S�2:O�nC��Dp����0)d*ϙ�hC�N!6�P9�%�{&�m��Z��ؔp�����>a?Ŷ�C||21CQn02��aOxA(���0<?)h�GJ��N_�ܾ}�'��ө�$ߑ�T��P��O��8n���Mq"&��r��M܃d�oI�"n�`x٬�FFa���e������07�\ �%Re����]�`N��q���4{J��;�i�LY����,=����%n�P�ir�� ��3���r�9X�?�����^ �褏��i�+�Xd�-Q��4�˦(8�}t�-�}��)�mY�j����mevׁ(�%~�o��S/��񼅡ي�o�1���L�p�e����� с�E��{�>����U)k'v'lT	b�e��� 4�l��e�{z�!~��%h���`��D��y�fv�,�� �#f�^T��""y�N+����F��r@�UcQ,�Jun�f�]d�X�����Cy��+��\�3�]� �zx�j��-�t��HZ��q�!+c0=�E� �\��	���VҀ}K�c	�o�O���qk�i�_F�4mn�Ì^�$U[z:�:@Rz/I�󕞔�i�}e��l(��Q������ۨ	|X�dP(_�+�N�As��Y3��Yy ���P��_tb<�A3B����u*���Z���1m�?2)1㢀��O������"�RG�[��R=����u-�I��i,}I��5��j>`��戚��r|��X�M�s�s���z�����u�p�]aNE�T�3UuR�[���_�Pwh?����mz�8
���e����E���%i[9G'Hu��'���,��X���7
�N`��ˁ�(p����M��xFԨ�"�.8@�ڌ��y�c+���T;˲��I
�^$Gj�D��ޛ����F��s���_��D�K
�L�cf*O�ҸKq�I��t�H�t^�QoQ�K��+��)��_�bȫ���8���I����[����� V�������ŧ�D����F2�@�?���A�/�����u�F��D(��UQU�hC:u}`����<�/��6��V���`eÝ�.�ͱB�$�jXO�	�F�xeX`'����3D֚N�ܯ<i��2��t�L���H[n)���2Y��E�Ĭ�Jo<�^H��Cjtv&WP�S/�L�㗱31Y/��������r�v��y�'��m�{�n���!D8W�O��	�*(�$�8�}I?`x+
�+�{�6�Ja��vf��QR�I��bextdz�[W�;G�ƙ�3Wn�,���y������x+�1�ޛ�2R��T�G�2Y�N��}dk���������.���>q3)�:E�@���f���J&�`!ʠ������:�1<�t�z%�l�v-�O+�.x�m#���l��Ի�(� ^�s��Q@@��'���Ag䤜KM�C��	8��pA���}��TS����s��'��>���Ac��V�f��(g�����Ś��Ɨ!��9�ꝷ.��NI�/���lB!��pg�{��R�z0�����h��)ܭ��O[�놜%��Z�?�#X��$6�S6�<|��M�۴��v�3��k�K�<r�IL�.�qU�������n��[��2���MR�/T��6�˸o;���B�i�Z���E+o��1�,x�f��@��+�2Z�)pU�<��e�I�ď)�9�v�E͖�C�'�*4�K$��A�O$E�ta !I�Sf���K�5�9��z��B���)���%�Gtߤ%�wT�$�)w����9|+�x�ο� �#	i��:Z��ߖ���*?������ڹ��M��w��m��K�f-۬j����8*-�rj��On��T �������5�����6�L��|�)�#���Z�����T��x�^��3�<YEu���8�n��B<���4$=S*���7��v�|!�1���g����T˥�rF�Ҫu�V�|��t��do<z.ԇ��b}��(��*�|j�yv��E)�&�-�K�T��=�+�j�8|���Fv�W@ߠ-oz.��Z��OճK�ƶ�����4��⟋%���nА9V)�z-9?@�2UA�Sy��j�n2��&�L@��U�7֏��|9���p�����'�ZL���ӪyGM�d�|x�~O����6��K���(�S��k�Х�~"�����p��z�A�Y.�x�v!fM^g����yG���s�]��|}b+(�y ��d��kBpHD9t�*}�7��(F��Hƒ��G���g�±�����e`��JE�6�ܒn�
~�s�r�]�@a�I�����6�����E���t�7��I�[�pﳶ�a�A|�m�3� Pǡ}�� ���j0�Z��+�R�u��4�̏|��n:����'��Q������K���c�L��+4��jo�`��K��c,���:��C�F��}ڶE^T��n��/}S��-x}k��:�K�Y�
F�� �b�Ӗ�:s�[6k�W��i�1M|��/��d<{NJ�ӴV?�QL,m/�Ԣ�	�Nv��� E�*f<��3S\.�<�m������d��p��r��xr��I/�+����9�����Up����/4�����O* �o��6K�2�!oḲ̌DE:}��%���>"�mΝ�"�Hi�ؿP}˟�s<�auW9PZ�&%9�jUx+��X��v@M���m��3Е<	0wK41T����	�#�3��#�[	�
H;lN��E\��em��{�]��J[<����@Ƌ��G�ݙ���00�uy(4�,^B���T*֧� ��	�u_�����ګ�,�T�!�e��c�-P����,V^�`R:Ɇ%�%۾R��w�TƄ�?�"&�Ӂ�(s�0��D�(�'�|-i3Ũ��/I�E����~�𥃰�S�����\,1���������� �M����FqOqQ�^ɟy	��4�1i�w�j����@���{2��R�&e���^�!n%RD͘�ם��f�F@�1 ��W&�=I��F�<0o �qNVw����z$�1s�	�S���Z��S��?$�^���fM-�8o���ܚ���)�d�8Z\��;<܎���os�u:�j�PR�Cz����Ϻ.�8�4�)���ĺ:��/s} -v'Ykᩜ�Ò��#V]�=��T?�����j���:54���D �٭c��Bš�O�|t���l���_��^X.@�3W�O�����2)���K-W�^�/���[�o���DgS�K �4 m�����œ�uFG���(}Y\g_֬H�ĨQn2�P��Ny��=�A����\��űo��mH�|s-I��X�
�>�wG�$�s_��֏�*��hF�Cfp/Qͅə@�l�ǟ l����d#Ed	��&�t�=�����\
^(�cDk{	c���M_��u�9�`GN���L/:`���<�����	m�1���qea��j���^����T�� _8���5=��a���U��[֐)���5�&ij�`�[EP��~(��!�.o�ja0�����f�|�~��f�չ�*)�ə�i/R���I��:�6k/��w�_]����!�O��V�:Ȉ�6qѿ���`=;�\�|��2S��n�ti�PΪ�.��o$b��kcV�� �d��Vu�+�}����H�>MF|�-O��!�]� �/���������"	ljX�#Sl&��*t�����JR.����E���J�JO}�h�k�f�;��6^���m�@{����Yo�'�+�
����-��	�`~����G~�b���k4�9w��a���9CP����Y�Oq�Kj���s�Ĳ��ߥ�"l�� ��R�������C�H�8O�_87���,���b���ŽK;q`c�]T ���}�MX��;��fw� ���ۢ����Wa���j;U��@��+�	n�ip�'��<�AT������9��-)�KS��d���n����m�t]���x\�;��'(C�����{�x�O^P � �j  0W�t0c�c��BP/����8��D�����|V��ֆ��eݶ��d� �9"�A�T1�h=[�h*Aa�4��S\6�Q �㦥�:������;Tq�Cı�{��!O��,/�,���m�N��ҧ�Z}��:���
.�A�d��Q ���P���H�HtLvþ ���7a�Z�ғ�D����U�5� �F���C����Y�]�TkŻq��ߏʅ�����tސT&-�H����PNp�;� �T��y�����VM�Mo��&�`�9�r��u*��9/8-�4+�ڎ%����=����1��{"M/���1u}�V4��D�/8	�q�Y*.� �\�/$�>�����Z
YQ�%�8f7��'d���B���r<m�ך��ؤq��������ݟq�O4�WI���@� {�hAW�rj���z�$�>�u��+������xD����"@d���=��j��U�`G�	�̴63T��h��F����L�P����e�+?GZ�A	�5J�*�v<�"���B�}�%ӳv4'V�Dk�N(\&����ŝ�-N��v� ��dle�o��w�PQ.hh�aTA�TIo5�.f�a����j�=��LXe�oz:Lt�Tb��}�zU�ԗ����f�{��ٖ�(s��(�k%�3��X���������N2��'��2<|A���+ף��T���r !��a��b �Q�0�.����]aGFE��j}�?��i��'mB��4�Mj���������^L������(��㐊�D��Cв��FQhlm"��3��m�ݺ�@� ��v�nգ�
cJ}�)sfa�:g��6A_��0��f�D:V��"*�����%���`���u�$�.f9�V~i�>l2���9�Ⴣq�����$/9gw�$� !�D�����K�����	��^�Hի�:5�
��E��ч_q�c���wpS������^ە��hMƀ\�
7��
o��KV��FC�T�=���I+kXԐ���$��<Z�zkbQԔp�O�)�7km}'���f�'qѨi'�Y��e���z�ͨ�q���0�CC̺�J�C�;�0�&%�������rQ�L6�H?�R�	{�Ցٙ�j���7�yO�y��9'$ңȝ����ۇ����;��Q��vsf�I�x'��s���˶�p�H��*e�@u�M@�n=����䪫�B)�f2�i(�N���~(�T���z��#3iǭ�۷��}
�sЙx���=���w�"P(_y`�8v�f)f-�pJ=PS`	��&}?|ڞϙS<�\�v�ｔl(ZZ��	M��"A%��L�|��࠾?
K��U��Nyt�Y�O�>��X�_�y��'��(�812�7���I����$�q���K%>�8�Q�
V��������0�2C)ɓq�Qa���#�2�6�*l�I.�4�[�_{�N2������L8{�t�Ц݅�ba�^	�s��KU��n�'��#SI_r�(]l��H%���J{�1�d	�s��nlB,����� 3�DASk�����@�kN�s�sv�,�>�]�n�/4J���ް$(2)��gv�r7��}b�Oߣ?>�]%wib��3��ǵbM�%���0�^@9՚��3?\Ɗ�s,�b���9k�p���.����N�`��G�ŗ�L<���aꑊ"�N[���<}���k먼��Am���;19ww�c󢠕�
�Fэ�5I��,�p�]�L�7g�VQ��[{��V:���v
��S��#��z���?t*(��.����
d�#���XeP��1 ��1G�����\���Zc�T=�,��'R+��	�ⵡǳt��'�(�˖�2��"ߩƠ$Q�H��qaRx2T7��C�,�M�:*�+"ڋw��W1�+VJB�o�5V��l��y����/Kn�[�꿤��b"��G��_g5TľF�a�تO�hՓ���B��!W`�pܧ<C0S��ȹ�hW�<3W� l7�� ����mI��,���0@�Gs��
I�?�}�@��͛�I���]~�l@���p،O�s��f��w�"u�(�e����^Vz��|�5|���ݞ��BD�y�$�ђ �ڏ�j�s��3,-N5��YX��z�bh�xGGj���	A�X/*�m6�u���m�Ӗ�=S׷Mw{�k������#(���o67q�h{�~��*�i�	�����6e���s+~wŹ��Wjm�`���A���E$LU�2����:�����S��?����BU!�8,��RQ�<,z`<��f��ZJ�'C_Vy����psڲ�P�e����SP��J2�����Q6��R�Ixk�	���T�į��$�b`a��Գ�v���uf1�	ߞ�D��OK�3G*�J�)�V���+�jӅ�w]L�!�v��H�<B��:�> i�$�͟ͬ�87\GFJ�eE�1���[�!�<�l�^�B�4�[��v�:�0:�w�夫=��}E�Z%/S_Í�9O�k�a��耡�����ce�O��=�0�c|���}\�u6q�r7'+,Q9����F��@7x�^?���r�b�k4w^�M�k3�ގ}���Ïx��n��}AуktDo ������ �����,:��j��郞/+m!�sMDyb/z�Cg���H�\��#>�X;�P9�1^����t�B�";z�����	� ������D���z�0&o,:3�&�[��sh��@�r=D��JU?$��V3��	[_fmC�����S�DL�8~�Y���\�[-&��y��( 2��m{�U3r���Gb��� Z���P5�6�N3:2�͠u0gu�n�io�{@OgU�a�K��:Cl���#�-����X��أ��v�J��p�o9l�&���t�Ϳ����X�r��W�e�be
�1n���S�+||�ě:�݅/!�#)Șۅٰw(Y�V��h� n��s�`^_�/ۋ�F�
ހ��Tõ�W���<�b��\��	��=¼)��$u̍a�ѧ����ϝzi�L�У/��R����(�<R�w9����2nvH���Ａy@f�^�HW:G��p��{Ɣ��аah}S�LK�QX-���Zf��j�p�PІ�X����Qp��u�{���Y�?�9'�m6�|����t��Q�8�4������S9,����]�P/D���r�B��\�<�v��zڙ��g�PGpA!�O7ɹa�wΰ �E���R��|���D6�l楏�t�fr�"CS�$�[<��A��s��z�O�Lj�v%e��/��'4Y`��F,���~6c֤�[�Ĺ��V��	�W�˔�k����ۜ`4����n[�4cf�����Ճ��.;�(�U=�6i˵�Z8�n�sZ�M�@�~F�ܖ��ˌd�I�=�͖+WQd!٩B�d-f�;}*�)�aߺ�����ū�nF{ϗ�.!YT�q�vT]��ʉ���lQo��7��`f�0S��M�+9���m�h�&�xp�������8�r�&#���F馒?w/�7���V����|q� �yrOU�������SZ%�ͷ*�j��jt��X4�u���-{b	�7xj�zN�f�� f��d�Ќ�F�z��U��Ȥ�V�#K,����ۀ��ˀ�����m�MDÀ𪿆���,ܚ�)�j�T��G�& ��(����WSby�����gҖ�y�v/�@�x�E��Q~[�tj$�D�.���V-=
}}Ϋ����~�������5��`L��a�ly��H��y2É��$Ia�S�|��t����o_��c+�yR���^V������T�S��e�f��� I�� ���tT����f���{�o��T�L�-`.��=�7h�x�g��h��+���X���N����
���"e����Z�a�G�:(�vs�����N6ɦO��]�<\��Rs�m�V):^�fCA��XR�3*(�ۉ'Զ�r�{���1 ��{��!i2Ue��R����62��(�~b���6'
�w�M���������j��:E����y�[�p�E-_؏��cϐv�}ēh0��MY7u~Ȗ��Q��
�,8*A2ȏ�R�
G����W��ib8s��T�;�H�CU�~?a�Rj�z'��$�B����:m*s�|��������%F�!EaT���]��9�;�����>��:��4��hX��;�Ԉ:-�(�$4+�IԔm�2�(g���d#�;�pA��,�G��(o�:�,![�_�֡>�@~�p�4h��Q�%�c���{�m'�����h�x�Q�mԖ�h9�SIk�R�?��ة.�_ue�e+߹�o��y����Gz|�:Y�3,�F�6)hIZ%F�?���a�:)cʧ����h��H���9ݷ���.Y@���ĺ�O��Ƌ�m��*�}ܽ$��x��rÆU\m���	M�'K"�x� #Y�E�~�D(T�Y�vc�9�=P��|���a�א"�Z5U��kR,�C2UWk���D��wm��PT�&��K ZVqKP��*�䌎s��7=����K���;qV���w�BH������m�|�+UosW�>\l����x�1�:���F�F/�ÿ]S:�����i�G[~ȗ}�����Xf��kM�66
;�Zw7d����4���Hy����+c��X,�3�M����R�E��Ή�*���0��y�Dywp�i�g�|g�BH��/_�<ۅ�P��N��\������j��E֧�qH�Fkۖ��
�(T)PJ��+�GE/�Ű7$���h�g~y�9��_/S",MC�[ַ���Z�U qH�WΏŋp=�hU	��fI*�;`���f�\�q�i�Zэ��4�P�8�j�rV�a��8Y�YZU��Y!tr	=�)���_��H!R������-.���\�!Ma�%�ٞ>����-�V^*֌쮚�G�����Ǜ�Ou迼}
�����k�d�	;��(  
!�tf榖��kDrN2����#�L�-bi�%3k�燛�1s!��G�p�«5�����s�������{ ���C��pW�h�u��J�_&?��r�2��.�E�#N�{��N�
Ù�,�˧�Z-&��k?s�&��iQ�X%��
�=E#]������S7:�8"z����g��4S��]A�Oc��ҜIܦ�3�$��m�Vl�rd͇1�����I�j��@�(�w�ĩ�E~������V�L�(�gtJ�};�j3�T)�M���4*]ez��^����Wȥ2�l��F:+�1�/&G��h�Լ���T�<���:��K��<4��O���Ѯ�N�@�������kb�Jǌ7�����JNo{)]�c@d�4���rƢ�y*y��-����;�|��%���d(�\Q|��Y$jM9�p��|:��ӄI�m���V�h۳3ҫ�R-�׀N��,շ׮Z��v��(��d�y�<����1����ܢӣm�s����w�OC_��$��֤H�o������I*ZyQ	5ծ��9���Fۻ�46ZP2��~��_�0I�/���N0\=j�6S6�؜ڇ��a/�!��Е;��%�4]Ֆ->�������q�*��1-O:?�OY�9�n}��-w,��~�i�/���3��`��/O6���x�{;�Pp:��y�0S���W�*�Y��q��oX�B'u�9���~�����q\N��Yqd��m֞�d�4{1����f���Iٻ����˩����◍�i�B#yi�7��U㙾s���V��ά A���!xL�'�ނ����ET�}���&�9tq,0:j�A���I�p�C��Ԝ�y	�(F���	�u��Y�=�@S�t�|��N�|ω^պ���U��S�<X����"2���R����2���k3����B�.�@������
��v5ں�c
�%p��Mt�k���5
��6���f��f|�ԇ���.j%N)�r�i���si��wK�k�����/$\��I�	��.��U86kbˑ�QՏ�	d��7�|WRw=4���KH��,��P���#��$�y/�<X�X�#����I��+@����t��<,F���N��^����ǫbKP����J�)��C$iE#�y�(��@�ߏ7Q߈��!��N��l��d����3��TwA<��T��E+MK�q2���#R�'v��`�+6v��8{z��T'�����1��mD�$	A̅�`��+�ʀ��ȑ���B�n�d���^\�6������h��C����|"_9��'��~60�:�� �߭��z
�pht�1����Q��4��gCG�%2"-3��E��·���=�
�'?�$�d��`q)�&]V ��Qk̎M�c�Hܔ�D�����S���0F�K^��2��Tx�g]��ꦱ^wz8��=e*��3�8i
��}C�Ɋ=�G��aKϲ��!4�v�yo�LK����@�dJ��L:dΰ�Ժy��?>�������@"gU�3�jَ�j�"�5)��`� ��l�����������YᒛE�Y�4q�!��ӌ���M�	$��hS�{�q��e��)[��M�4V���£iI�S@��u��bN	�r]���a���O��r���
�[��Z0hYT?[�i��#���� ړ�tCBn��QQ:9F.ӡ� +y�}g%�Fr���bHCXM�%A(>�j�i`5S遃��}�+V��!!���R��׹ �� ��B��o��}�X�a�O��>ߌ�M4<�|�:�&�+k~: Bov�4^�>D��)�Vb�*n�;gZ�X+�����[b�
U����+�u.�/�'�8���nu7�Z��)v�C;0��ph5bx����y͐C���.���/�����kb������E�a�R���Nr�ۯ���*��'��b����l ��-YP�ߤ��ۣp}%l*�r�e��a��W?b�7)o����D�� (Lǣ�,w��vc�o�esFd��D�zD�G�o!�� Z`V,j�n|L�;�b��K2��2���x��1p�r��Ɗ�?��*�����Uk��`��q2��D����B�G�<u�~�m�Ǝ('Nb��;F��.�q����� �4j�LYZ�j��H��HB�7��.~R�iD�N=s_*n���M�������Ҭ�ڠ`�<�nn��9	���ڙbf��h������ a!;Q�X;��Q�m����5��7�t��#,-�#��V�]�O@��=����@p%1<o?Gͨ�Ê)�92�H}��󪈿���C��?vd���P9�_�g�}���tɅ��a��lJ���O;g!�����%�Oe���%ĈŅ�����)~Fn�_�d�IN]����	�E�^��X;蔱��=�Tof`��4�XsAj��
�f�o�^�}����-%8���k	��V����vc�:`�k2\�Ý�7�	Yw�T�uxk�%��{�<,z�s��������:!�o��QQW�h�F�%g�PB�hv�~1�Gk�ŷ&t��O�8>m���SQ��'��A�p�7P��?�'f�qZn"X��Ez����P�b�4�E�ڴ+Ü:�>��s�`.���6^���튣�u���b����PrE���;�>rC������	o?�m�":�������w�=Za�>�3a�GXSNƑ����
�g:Y* n��ZX!�<��
vs�ĻiftVOl�/)�(�uZ���;� � ���Ba:z%�򰦞ŽԺ^{ �Jn��(�tH��~F�I�>�����! ��u��G��K��O��
Qw+�e��������m�ހ�#43���A��H�NJJ�W������AC�NƠb��b�e����΄>�[�̀�6��ZV|?�l�:&���y�Ex�<O�?U�E� D�Z���s?X0�	�$�H-���c���Tx�
�X���Lo#�+c*�\z��㗏��~��������`]M�uܥ��bq���)���A�z���hC�Ԓ�-j`�윆�~��Q3H;���L��yKa�0�w�`�����Eag��B2�!������H��sD��{��Ne��W<�D�ҡ��̜����Z��/h�(U��s��8������UH%����g2.Q@T��;F�{�r��ye�"��K�L�Sc�~5;�6�7k��c���ş%x��g���.�+:��xJCg4�G*zԡ�o�� ս�*�8�^��B�dS��ߩ0נr���tT�xf�1Z�q�;������Ȼx��E7P��{�q����t'"�$W�:7��#�0~��v1�J����Z=B�~b�2M�&����%o�)���
Ҍ��1�R�X�Hd��6�[2-�J��]B%��WA�[����p�B��n���ie��z����TB�	:	��O0�s�� ��&g/���;R|d/�n`�'��9�0�Δb�&���-�=�M(�U���������S�u���Z��)�2��p��@n4@L��!]�Tc�i�xI����7�{�Q���<N���m%�8��Fp���X'<��*��М��`�~��dP������x-����6����k�C�����q�O9�ߍ�~S�ѣ�J6�rc�ԇF�2����ϭ����J{�>wii�^XB��cn�.+�eOي���E��ڄ��T�=�V	C ���4ą��vم�ӯ98��RT�J� o�Ba%~����Bl� eS�ʩ1"9�N�����X~lݱ�B&+yc�ؿK��'DQ�>�L�&Ț��v&�~L&��xM�O���c5��]f-�7�z�yi4��!��Z��ɛТ˭w?,�L��Ϸ�[A�� �ߟ����"4�!0�!���'�e$Q�.�P�E�.�(�}�U�"r�M��.�U6�2m�<no3�s��k<���1$�:�J,�<Sd䰋�2�-����N��2��w��)��]c4��O�$����}�%�<�^W.+�|�*}��	��82a�+����&�g�>���)w�_�'�D�tˤ���z^�݉=��rTP�XxnGS�Ȕ���x?�W{KTN�wF?e�1��ٱ��U�'���A�k��!>��[�I��S§�a��*c����$���>շ��]Wk�ʣe�F`��izlDU�i�����փ�TX��iUbTW��#�ľrxϱy�%��[-s�މ��ErҶ �M�xf�O&��D�P7'�H�
����^����F�u��y{�e�3�A������­3ȝ�<c��u˂`�v� �ՂH�H��Lq�f���������:�)��I�̊��]�i^���RO	'p� �(8iJ�9ka�'m�3���T��W&S��.�Ny��#��2��L���������
^KC�p���_iV�v(	GP=�0�}Ŕ;0���[���{rj!Pb�*X��~:c��h�g�s<:�QK�yCB�N���OIѥ��wPh`�T���"���M�朼^b;ANU�q���c�C�#��"�� ������C����(Dh�~�S� �O�RDd�S�o�JA|RV�h����t�H�ˊl ��4�ɳ/#�C�������T��/<�"�Q�C��O�)�EOh�U_��� �f+gGg���a=�v\��`u$�I��y[8�D� ����^�I��EZƽ��{
C�6�l.�W�-V�h�w���+7V��"�vߓ��(]82���)s 2X��,9qP��ր�}�1�Wf6��3sK��4JJ�2�VQdXΩ�scq��!�~F%�l�=��:U��kC
:�y�[�G��뮵�����nr��L���G��hh�/��h�q��A�l%��}N�(if5U�77�Y|� �	T�Zf,��ᡂ��g`�LN%Etm�;Du���H)C�n��-�02�FeTR��nz}�#䶧�jВ��Ӄ�\h.�'n���L,�C����}��&��vA{�k�b�~�2�1���t�j�EF���MK�%���#.�D��ۀq��q}Fa�͆@鐹�f .5�}�8�����u�l�w����:q=�6  s�`=@t�{i]�W~�6�G~M�B�f�0ۨ:�pz,�����\ǥ��������&b=��Y�����LDÄ�����Ѯκi*Zԭ�`��s$�x��m%���K[	+wMո�� �Q���{�8�J���b�( ��M��n�O��˨Q�_h4}��yA;k����j�x��e��fwj������S�4�����м��=�J�LŶ>��?�:1�Q�(�Of�ћ��l'\|�ZE�?J�� C��{�����|�ޖ�G屵��HI
�o<�v��<�2V]�I���y?�sUMl�4a��v�.���U�#���%؋����r�/�7��ydh�k�����=Ock�u'S*����=��Ck�lD�yZO|�:~����,��q.����'���WM0�T��m)x���d�w	�p8�f�~f�YЗ��G�ŧ�����Ò꠸me~M�f�й��t�z.�3���_G�Y�>Ϋ�N1��x�kZ�����_�D�����<׸׈;&��-����<[�p���%���hS!z$����gc_��B!A�;?E��!����D6Mm�l�{�+D�C�u(h�jW�0��䁣s,�;eG.V���H�$g����t��f��o_$�֢t�)<{��u^�]���ZQx��sfi�B|PDlCD��bDSH����%�O�xG�?�j���ĊH6���4�(�^6W��3Oo�����\^{���0���-��,����0����DB�t�G{����丢/�"�y���:�Me�.��.
�A(�!CnL��
���S����z���|@��YW�����h��X\�2�/,�ZꗿD��r<c��c�Qס�0σ�V�M���lvl���N1�����]�Ʀ�bC-��7��K.1Xs�!��Id?�>$ظ��g[m��Y��P��U�ϝ/Q�|D�_e�/D�_D���nv����W-�$��$���|�RS��z�|��`ѯ�b�;U�J'��_v��{�[�Z��l/��砨��;A�\t�Va����}±
y��?G3\�4�_DX���=�U��ʛ5O}�bQ�>�?%�s��Q�����R�h�������3�d�ʼBN=Om���!�>�c?���Q֠�S������(*��6��D+ܒD�K7)����k���q��a���{���l豞?�)Z����Sw�ފ�'�Y���aԙC�XW6u#���)�1�j��.R-�����>!m���f7��3��@N�e�8��r���'�#����P$u��CN�L�m��;;��b�7�*�������c2,���X����G?��H��7Q��g�]i��*�C��( ���/��S�wA��j��b�1"
�S-��h\E�n]l���#Te�����k���������䤯9Jf�>�1$�4��-g�ؠ�o���Q_k����+@r�i�E}��ak���6�w��n��&u�U�0�WsA�ɗos 4�8q��b�	��mf�qSgZ�y
�cR�k���݄8���޸h@��oa�����]5����Z6�H�4��(c��gţ�CQG�Ļ��J0M��yd��m�������Z�EIû��I16{Y���Uޑ1���>ߙ�N���}�Ɓ�Ԛ��t�1B��q�H��X�ĻC�T��
��Qm�jSM�A���YSӃ����j|&�A�Yv�-�	+=cŞV������9nd�4���A���E�zKv���l���+'��L�䤬N���Sò�<-�[^z����4��w��
⽜����6O�G��/���k�������ԺF2�hS~+��)��'�BX��p�Qߧ�:2��OXC�a��8h��##����K	���j�K����s�u�"N�7)�X:r��HἾ��3P���,1]}�����/lE��/aP����[��5�*�>!W
�S���-�cY�A�?t˨��[R��솮] ��x�}�k|��sM�jHL�j�T8��텝�i��KH�N;���y�m	\�svH��rnd�b�ơ"Vb�X6��c)ƴ��#�b8C�����E�ɪ{���{��}�,�)M�^T&E���傴�KL٩� �]4^�����Q݀��ă�ؒ��ΑG) l԰i����W�
�j�/��[_@�o�,}��؞iߡtisK����aUŌ��
��npB,$����q�k���u;��?{��8�5���% e�?e�HGU�:y���\����!Lt?�X���'�!�bm���I�~�\��y�U���.��WU��[vo�a����D��yv�*2�xd�.�����w�]��S?�k��UIM0���焑���>��<��ipp8��ϟ�}�'�8h#ύ��5���Y�Ԋ���)��F���Νv�	?�I5AZ�m�ؘ߆bÂN�Z�BHF��*���מf$��ʏ�\B�7!SRl�i���̮;~/��R^�	f� �\Go��
�y�&��J	ء<����!���{x��l�(�������_͞ح[���(S�ח�B�m�����`��"$R��� �v�O�j1�&����:��j���N�[�6=����fI�H5F���]%i,Ǜ��I�O���"�$��n����Z�!����L��1��x�g�8�HI��o,n�N��],Xe6����YK,W�gaBd&��s��&�e�E��򻉕�Y����/����`���P��9K��9�&]y�����&o"w56�l.2j���O����AUࡷ%�<��9�i�E�T��6Njɘ��+���b�o��H�ꥊ@�M��k�L��o�<�5.>�5�n�����)U%njl�ʚ �+�z���м�p��.�����C��:�X\~�o_��gs����5��77�-Y��RQ��7n1>�`�pڏ�ؖ��x(���AAc+.��5�������ԭF���<O9�����ƺ�� ~,����~bD�D�ƒD/W��K�0p�M�����Й�I���;�Q���c!#3���V�@�E'���dg�K(��c��i��|�Z��0NoezP�=���>�M`'|�h�H���n��PJ���9f%I��;�{Ć�VC�r���<�?h�N��F!�P?x���3Ζ�7B^�Ieg���
�*O/�[��ɮM��a���m�d؏C����M�� ��\��9��� B��n~ WѨ9�A;:f%KK/!�J8��Ld�y	(���[L<�SX�HB�| E���J���Ӓ@Z9a��c{W�Q�i�z��Ϡ�,��}͕��m[..�9��[��.�V���sÕl�K��'.�����K��y^[�۸����
\O�*���Ԫk��8��or�[L>�'ȻΘ����}�
z8E�0~B�Z��}�y�*z��㻪9�#c�,a�i��φ��s����֞&5j�s�~Co����rھ�Y8�3J|쳜��*�����>P ܝ���k<�*�_F|�#tSĮ��~G��Q���j��7KB�v�k�t�D��CL����J)�1ا�
�E@S�-�c�P8Ǣֱ2�v��Q5tOaF~���K���h�g`��宁A�Kn9�Aڠ�>ε�cbi�* s2��	I04E��Ʈǅ�����Ue��P\T^�-V��vb��C���:���)�ԦH]�gF�T�A�ygu�{�k��R\���!�j@��I�y��3����_ש%��=4�M�g��~��aY`"�Ra�-詴�	��
|�� dl������H�'�P�ٰҴ�q���@Y�r�vV�{�]P�D��99x�_�0�LQ�S�j��hӧ��F�������w@d��q���
 ���E0�F�V�o��%�q	��|S�N���}��8F�v0����{=J��+{B�Ԩ�7��]�q�蝲�*����.��[�6�&�)O/*��?B��t��d:�xW=�!����"�YFК����Q�[��4a�#��5��n&�����+�i'52���V�\����O�%�/����+����j��I�	�+F���[7d��^�N�+8`�����[��	�	����._��F;����%��%�2���f��_1[2�ggZh�$�	,�ڎ|P�6jU�V�7h�8G��� �>��[����|8�U��ejĚ�o���mpnߨ�z幾g^*aK� Z��\��.�����"!��<�I���k%��˽v0]/��eٻ�n~�N�����������I�*o#.m7U+�5�8����b6@�s���ï��c�HQ�����U�w��9������= ���Ef�@E�f5���f�qO���x�ʰ����bA����	�sf��^|�=�b&��`~ǲ������;�Z$�.�qj���:���.?�B���h� ��~��PI�F������߯(�����t�n�9�,��[�{�
�uLk�Ibi �P��:[OB\z���ӤUG�`���2m�}�4�n��{d!���aR� �z��7si��-�9�~�) 1��c}|�ݱ�%��SB�����v�F�ˁ��*��8���k�O��!�C�ZV`���!�ښ}�L[/ʿ��ڐm�Y�ю�D �,V�ݖO��S�-8���黬������Q���{�eG1�G��sn,2ܬ�+��z����_[��m�%�ܑ��}��KM)(�b�5�q�+���)1k�ۓ��խ��nM��tN#��ޜ�%n�̘\�<�e]��6����T�oR�JJ�ᰞ�B<l��`�9a}Dd��7�~
��8H�y��m�7Tϓ��Q�x=���H�(�mL��a��cq�֞���d1B�N_,�+7Fe��b�^�Q�&;��Q*�0��08�w�sw0��Z6m!��'��U)����]H��TX�\Q�AVB[���w��u�7�Q'�U�%>��?�G�A�S�]F�7N_��*�.��s����&��ֈ8��2��[����Nc&g�Yxl9�JE3�4���%_�7��h�b�����&Tj�5
/�4�Pa�RI�,j����`�ꄶh��ٍ�K�]��}[���:R���2�2�2й��۬.�@�cs~�Sz��<~�c>�$��k8���낭�W~I�˲N��S�(4��΋�<��n0��;�����.�lފ�9�wr#c�d�)9�{ْX~��`|��O���nZ�eP�L�|���>t^�:EX�S����D�Ό����nqҧ
�)��ٹ)eL�T�B�T �"�2��5u|b�J����;G�fg#8Q�h����D�| �VҰ���RA��0}K��ol�ACIW�o��z�x�=�e�	Aݭ2�^�ӷ-��bɓy��9��{{���Ε����+�����s���T�:��?�D�z�E���YG���?�ѳ�=�����'S�H��(����M�o8S�q kC�� 	$�ҰB��sR�%�t��䲤��?b�[ȯqJ�0J�	����琧e}R��:
�DX�ksU�ܙ��zE�옾.,�p�9i������pD�I=�5�=0�Uծ�������p�1�DL��Ȉ�laD	w-	��GS�9��"��4bER�
I�5��)�I�ܞ��@7b�	���Hw�=P-�@	��p��uU��!�Za�ۀ��u���CH�ȖEG;�?�� ,\���=zTg+E�����+.-�T����.�1�R�SU!����M�Cʖ�|��u��S�2(ߑ�뷂1����S����g�+�)�	Mf�u����qR,A��L��
������`A˹�l.}��j�z����ec����`�������)�F-�'���C��x�s�56W����ڷ���B�2�h�����]�Hx������ :]�}�I�WlsYN
�\�-�Ϻfle'�6]����m�Hb�J����`�En� n�ŷ͎��Yzf����q�q���8L +7����;].�س��c� b�j��u��ħ�]j��t�.�X�������:f��t��(��. |�&6W"]!���0t��Ċ�A[w�̜��by�&��L�s���LkF�@��GָI0�7��� �l��vn�d*y\\]���eM6+��:����;nR
���L�c#��i�^� ��u�t��*4@V��h=p���?W��+eH���#���r9�y ��ݷ��Kڹ���f�
�K��������8�b�QDAE��Y<�D�䰲�NB�Xb�';�N����x����J*�S��������9*V��clbq.�n a3�]o>	�=�%/2�4ڞڈ�g���e�
釾��"|=��ZC�
Xʧ&ͥT�{r��_�_d_�<Z�C�F H`$��S����s�t����sm0B�|;��e
��5#�mxKp�����H�|��b[>1;�Jd��2XjY�9�d�=ë�檶۬0�ƶ8rƄqMf�ęX�쁸��*1h�0�8A��c$V<*$Uy�J�q�n�9	���{� ��8B;��%��gj@�[Q��3�ZI$��bef���ZR]�����M��{�-c!n*��C����(��!�o
4�J��8��: X�2��]���J("�+����t�,IOc}Yxĥ�l����&_�xF��"��w��_�3Bn�:k�>*=
���mA�w�N�Ea�Y.�΁��G�	��+�0�w\�`���"]�mZo�2�)�,����$㰸Mz���A�����VDX�j]��ek3k�d�T�/VT;]=9(M���R�����]pn�����y�����r2�;�'��8k��_�Q��o�?$0�ח��d]�X1Xq� ������X�]�H��K����ö����0<*��t�u-}�,���!�\��x>�7s�b
K�8y��?�A�_w6v_*�L�q�~:���%��]T���h,�ݻa�X��ֱ@3o�*1\	[�(�Z6IQY��k�]b���w���<)�a��Ns�$�	����p)Ł'bd�2mR�T���H����3��\�׃So�`6^eu��Bڈ�>� �uaHx���s7)ڒ�Y8�-�+g����YU��>U�Λ�q���:-���R��R[`S?�?]=7��_dZRwHˉͫHR���)��^T�Wj#��H����Y:	��xp��ܸ��=l�t�J���}�r: +�I�Ү�>��jU[�9�筀���3�UJ�f�Tmb���0�j���VSQ���Ω���10���#nl���V ���e��Ԭ·���~6I?-�h�0kp�$�r�u��3-��7~��H�N��8����կR�#�>0aY����I��l�7���wCKyq��a%�v��1K\(�	���<tA�6��M#���K�=��A�"g��z�_�[�"9*&�Z�B�?�7��'�
�v�Q��Ʈ���J��)BQ�8�-�bl^&��Vc^�I���#� ���tț���Cx�k (?]��b��	qG�N�v�*������&V6�S�D��k �x��v�d�K-����*����m�an��� /�+B�C�·ruѾ�R��E�4�1�f�a��P��h1��-{b����X:�}<�m�LT��qp';�4�q������#��T�"�2�W�> �팸w,��$:��#�FȈA��/�_}.D�/t4t�Ǭ��Τ^(N�g�dV�����v�����	�Lk�����	^7�)�_��i?���{}�8���� 6-���K�{C��w¦���ӧ�2��"Gһ��+�4�I?O?�nޟ�w����~:�V�����|A*d��:�]lvr>� �,N��-)�l}]Q8���s|�������>���$u�����_�UC���F�&!Iq��*%��Fމ$d��d�&���_O����[o���a)ZØ=�zQj�ljy6�x���=�49↘�J�w�S����Wy���a1?���l_p��^�������ۙH̞�j�!�a����J���u�+���5�j��~��E�7H�';����% �M�� O'�h��bu~��4tbj"L����!Z����u��Z�J>�KsaliB�A|��-9� �b,U�����wD�3�< �`vt� ������֚��j���@٫!�]@��I�E7�s�ʿ�&���U�����)ߤu��ੁ2.�:u���2�sl��j�"%���=�^*s��cс�TX����$��e9E��?E�`�9e��o���� U�R?��v+ ��>GT�1��RX6p���j.Qo�j}�D9Ȳx˓ދn7z�2���%!U���(�v��щ�����[�)�rh�YR��3;;���`P��*�*J�}��\�x�3��v�J�%*q�-I���)����m�߷�@��~��@vL��JY ��������Eæ���������i�0Y��0h]���Mv�g��ܻFm���ӏ�hz��y��7t�_�*���;�Ü�>��&���'o�lE��m�� �Z�z�~�k�[d�g#�i�YP��nҐ����-�����_���-��S��Vw,� *kW�'@.+��΋��P�3~S�j t�s�H�!��@���#��b3����^�s�'hѺ�Ϣ-v������b�3�x����,ʷ@Ť��-�)
Ţ�p,1�E�m�"g��Tyf��~�DWΟlB,B��R^�rY�BO�0w�%��E��cn�ü�'����H�υΝ�[-*�iɹQ������v�s;?|�%P��T:�'��SE�_�0t�ɀIzpG�2fxq��[�A�ú��0���Dܡ�wc����"Bi��Xa#ōd���d� h��(P��qd�eL"]SY�� �I���d����B]���$~v4KƩ�
"��zن\ch�b�8Ȟ� T�eC}��kS�k�)E���G�@	 u<Z�e��Sd�3A���,�A��_zԤ�~��S/9v��=��f1����fê��7��	䐨:m�Dh`?�pK�/5+#����-��b� �1���GP�^ku*�.*�(�K.�c�:$#{>aC؅���}���T4{�\��q�][e���MJH�d��`,t��>f ��1%��A��4��eW�A�\��~�R�������k�	C��;tD�;0@L���N�Ė{�n�����%8��I"&;.c�¡�U�`aΣ��.�S6��f�@Z�����ܗ�)="g�Z�Hz���v<֠�yy͐��b�²F�#�� �S5�B�Ҙ�9���+�h�T�q��@L�����i���9D s@D ?W���B+m9���|�����N~�k�G����g�R�RX�S�D'�F��뺢ȟ5�AJ�Ob��|�8N��/By���`���G���93�Ƿ��H�,�9d �u{`�)�ـlه��))D�Y����Z�3��	���Ͽb�w����q�́))��D���2�{�� ߤˈ�^�)�4�4��m���������}�F/��N \�F�x�A�S�D��dZ81�m�z��Г&m���'���B}	�ʡ3�5X>Řb+��zO�gR���V&���7i�N��|1��3�H34��3;������?�V&_�T��f���5��:ۛ�t���o�d��B�͠]�8��!�2e!�G�2�X*(�Ix�P��C
�aU����8���Kl�J �ݟP���t�f�rל��q/�h��2��y�����)n���S��K�T�i=C��w%�2���M!�'�T`�X�E�Lr�ߥҋ��yd鄵 CN)�U�H��js��U�, f�R��LC����	f	�5X��s��-�dl�y��**C�c�3B`s��ҽ�Š�6�~i2��JN�<[�3���{̻s��h~��ի�Y�U^�D�q]]E�M��� [mE�%�1��0w��*|��ksm��Ch�L��vo�%"8�����k �-�D$} �
��,�)���z��#� L"$�y�	�^���9S�~��N���Z�t0���+��8�=2S+���淌]C�X�b-KT�:�:�^��r�����L�&�Q>� ���n銎1��e6_��傉��!+�Oh��ԍ׸c/c7h�R����#���M��"�O�/7��=8�Q���3w�G]�R;��ٙ<O��\'������$?{m4�j�?:�vTRW[gv�bC� ��8$���N\?��[(�����tdM��7�bʒ�MT�%��.ա<u4�X�t����C����Ҏ�n.���d�}#e��~*�u�Q��8d�C�e�
�"mߊ`�Ԑ�:�i<\#�\�����H��>�������<�Z��>5&+�|�k����E)o�h2�Z^j"��pr�*+����`��G�FO"�b~�a1/�K��nȥԍM���*�J�!u�dt��	2������;��	�5��84b�H��'���xߨk�Xx�1+��Q.�ò�ք�=Vav��f/�����O��방�g���(���}��A(�E!E܈���K�v��YT-;��]8ϼ?\���}�޿t�s,�J�r�+�P�ƣ��.E�L�����N��g۞b��>Tҡ��d�?n���+5¨,�����I�7o�=���|�+]���a?�PA�!��hR�(+RF�IL�PD��{l�}o�)�~�к���n���-���UCS�Y24�߷�<���TM�����4������+D����/!�,z~�WO�R_1�Y�\Ǜ!���D�a��5�F��3|8?`hO�qM��+Jl߼�Zl�G�[Esi�r�A��v��r���-;LO�08��&{%Dt���C��}8|�!nz������N朧wf6Ȓ^� ��������:�H_@y�SrH�����GL1k��x�6,�����@z���ʻ��C�����-8(s��K�!ƭQA�+.(���q���7a���4k�LGs��"���I�Ƭ�ғ�W�q[1,ə�DN� 0�0�A�O��?[�=mx��i����vl9cn��� ����*�yte�b���D��z���a�IلgX��<��t��U�3�Y�9) �o:�:���K�%
92E_�h��l�ԕ�6ѼΔ?kT�2	4Pg�j�J�g2̦�G�g5o��ĽqT�N���dm�	|n}�W��y+m����W@���41��i��!f�M�)1^��zQ�|-�O@
'mB=0Rq�`�xt�E{r;c�nV�������c�ɘ	�xP�S�4~���˺�rT+�N
?PI'����w�����Զ��I\$L���1]xz�r�_���ƬS]�g㓜/v�j!�W���;�ykH�����݆Q�Հ6)6h�W��.T���Z�&�?�z����Lxl,3L�x�$?^<�2������M���4�i��$�p������MM�0Ω�!A>9
=�tV8߆��"��li���Q�;/���6�b
�gpS26D%m&�l�Zܭ'wW�Z�Y��3�uj�O�q:�pjQZs������ͷ�Q����٨�1�ȏV�{��6��A6[���O׆dc�]3'��?��%@ǰxH��r!U}\����P�@G��(ڜ@��u5$Q��?�������r�n�����O%
W��0Z���/g-����O�<�e�1�-�g��\��m.��7}%7�}�{���|{jC��W!���Ȩ�� x��O3��3,{�kM-h�%;��ŋ~[���pe0���Z��h���S�8��L
�"��(�[xڹ\tyd����HQ�c��h�wvK�����4��b��o����)��Ó�,Po�����ӄyY۲��3�.I?����4u�I�U�VG��"�ɩ} �x�	��~0��S�PTӗ'O0�����zQ���V?>ϙ�»2Ca�@����3v�����-�8���v5t�os����+<n2����6;
�$:�K�yp���4."W�@�<�E ;������OkF�G�Wh���d\M����B��A*z(��4)Jc>g6�3<�#CU|��b90z�%�s�a�x���HA�O��9�WV�������I�e{���L�d N�!41����3E�SR${�`�/(��� �*)������fl�V@���qeh:a� π�P|�oM`6.7�������^�Xc��!��j;�Zvm�!H��9����>��Z8����RXf �խ{v�t����0�z��q#�iԊ�h���Z��?�^[��$�6����ND��wY�����?�q�С��,�AP�z�����p�N���@^B���9�?b/>���w�v����&^r?j���Aæb]�r�J�0�X}�S�*k�f�ι�z�Y�,���q���
�!�Bw
�ڕ⸭�Y	!�ۦ�g�P;~�!�	��i�p�ݶA��h#� n2��D}q"]nq����q��I�hi��׀�)jI�<q�ϴ1�C;�-(J�T���V�<.�@��� SHL�
��3�V�V��en��4Pl .�a���OZ�$���U�RmY�Ywr��*Զ�ubl)`��j7�v�|'��>����	З7@��|���<+_�Y.y����/H�!Y�z6�j�c��(t���B��v�	�d�A�|�$���s�$1�7/�O;3�'�T�?j5�(5*���ӷ*���j,ݢiB�Z�������j��?�ΖDi�y�8T+!�O��9ǖ!.�R��^��~oU��q��W4^���R�̡$W+0G���2f�QT��Z�:��s�|��kV�dY�T_Ɲ7��x<^Dy��g���'�A>$#�\5���]b��5ʮ�@3{�v5�-������F- ���G�M��W�]��״<�O������P��֐7�e�Z�F=�?xz���suD��w�B#MҺ�+ٮ��TB�2��ŧ��ڝh�&9a1��[Mt<�Bǚ��'��� �(~�-ޗy��zLr]�g	>�-b��C�z�$�_|?�H�Q��������bC
n�X�����t��]{=s���C�C�ª��MV�2�w��8�z�$��9��{���=�]��׺%}�����$�+�W���#��NMǩ��w��݁P�Κ�<,*xp�@D7���w�"�Ͷa�դ���C���w�/2������=������Tbz�F}T$��]en�R��˼"GEh P����v'3�0;2=�ߨ�<���m�u���ڟ@��mr�v1�j�ݶ h�/��=����'��
b����^�M��U�mHU�dJ*~��#&�0%�Ӏyr�y�z�M�5��6ƈ��o="'���9��-w�>�ձ���WKK��5�&�⥒��QM�l��۸O254zw��-G0��ħ,��U�M����o�_n��á�R�ME� ��-F����R��֞7'&Gr��pe%���#h��?���7\Z�j�H�� u���%%�3Hn�)ĪD3a����Ś��Y�b�݁Q�¹�K�=�A�=�v�<���W�k�c�]B�V-����D5�N����[,���I�h:Yc1�]L���&4�5.��"-o�G˩���!č�K�F�zɮ���nDs\�8Y���.[V��1S�ru����du����*>�rŗ��ox�/��X��~�0|��hI��������ԝ�ߣ��!ܹ,a���81К�G����1e�K��Z
�D�i{yB�f@h�i�@���%Xt����<��WM����x�P=��e��~��KS����K�]P�4��Pl�m���� Q����	��9.��dzވ��L."<��#���ҙ3���N�:�u�Ʃ���Y	?g���j9$h��L9�7��uћ�-���3+ȒQ)���:N����,�@�&�I ��w�3��t��i0/�z�\⤺
��V�.��	r���7�K���[��ܱ"iF���q�:�D�)w�����d|�٣*ijb�f�aҍʏ�<jM|R]U��1�pU��n����f8�6�Q��E@��s:+�Ϥ/+��\K�[!�����#�и��̇`�(�[<�_k74.1	�]~��nY ��ۂ�a��s��ޒ���'Vu�O���j�s�1�������w�=f�G�6k���Ǳks2�O���宭���Ѐ�H4h����ε����\4���V0���nQ!5��������um����Xo��:�J����B\��]�=��RDȡf<,	Xێr˜��y�)S��d��z����Z�b8��kt�X�����5E�&��葚$���|�Z ��mK��WK��#��Oe�v���}�Ks�[W1�-/� �R#������>ӳ�b����P��G����
�z���B� ����
 �Y��[~�����-�늽9f�۸�]B<�Ȍ-���BE^hg5����u��)Jg��q��`�<EOGyO^���}�N3�S)���(�s��e��"4�<p0���6�H]��Z�_��8~��6��:L�_�?�y�(Eݮ'W�ہJ!�E�h��t���9��7�SG$�}�VH�@	��"�����x�6	�%����*|�d8u�+I����D�����o��j���p�ϵ`o*!*[��"�-Q��a1bj�*F�܉K��0fD��CT�Cc�mqO ���&�=�eDtG�$��D m,Qz��Lr�>H�!OEg���F3��舋Q�+)>�!�<�r��Z�a��`�$�?6Z���L�����v��a��[�F��|�;�g�`!���?��� A�9|l��PA��,FO�O3��fs�q ���
��=\�=��2 ��s�4�MȈ}.�*A۶�y��������;���"��I�{�TaluXP6W�W¬N���6Y�
؝��!Iq�n�ΣI��M �g��C�C�� CC��2�#�{�+3�UҮ��s����䪾)*�	�ʱ�>i�l-�wn�_���ն�~��4q(�^A{��p�RQz%�C�ъ��2��{$��>��m�g߃)�o��r-��ԇKd:M�
��!��kB����"���Էu�����66�7-a�p��$�%=�����"�*�9 ��<�a��-�`zD.%���DL�IY)U�C���K(M���cL�7���~Tc$x���h�ܒ��-��	Y�����8Q�<{��R����soG��ܝ�Ӯ��-�Cnx�T�d_�æ�>_����;�!�pӼO�!<�	߅�5�_�JW��C:��ٮ����b��F��Ouq�2�n�MϘ5:v�i�o�V��Vt��v�,��Q\�W����^%_�T;a��,�u���s��R�zJ2��3s�V/#�NY��������8h��*zV���Йz+��VH}�9a~|A��b]��~E��iÕd]�\����BDI� `�9w��d�er����I�$�#����er^)��Q�^C���gݍq��@����������W����_\�<h3j��V���y�hw��UF-���zɼDɄ�[sI���QF�(�uV�1ϕ����xr?p�t<Y�U�\��ga���_^::Հ^�4_�bӘz��!�"��H�j�z�����/�y�S'��$f��u~���f����F��!���E%�3O���ŕ�N���^*֋�PY:P7/R�D�LD�J�cŨ���Lsk_s_�5� t��@����>V��1�H�T���H�x �ӟ������C6h`���
!<6ƃ?E��d��ȏ�"��n�úr�/���08�p�'��K �4�!�c�6�6�z�չ����Q-^�%~�
S��+�t���������N�A�e:Z�c���X0�C{�����@�������M�#M�(m�?�
�H׉�6lq����D˺����E_�d�|n�n5�0�Lu _(�G"�B�p�g�� �q��q�K��`�^���]�B���8���Am������X��s� ��dpL�^PV��o�)��9�"d<^�����9�k(A�B��+{��+��߇�R��Ȍ7��4S]2�]�*ɔ�ŷ-�ޞ�˷��&��q؟B��O�B�q����y� U��ޣwT��#�:V�����E&�q�/�/)��+���<��^��By�d2
Ӫ�tjr���*�S��FY�	��~�=����P0,_��n��fH�����Jd[1�7��O����n�V,���"*��Q���M ����%7�x�!F�𷧐�ոSz��(0Hl�ˉ�
F�#����P��E'���0�54k��f���L�>,D�a��3����&�;�H��֐�H��^�x������'���" t�%q\�A��������j542d��:6�K|*DȪ>T��V���P0�<_��.�2����:���y��}�����YN��$�X�L���M�Z�fş���L��Ҿ�ǒd9�nE{-^}kiTo��]�Af�#Og�3%�l�uf�Yq�ۧ�8Ä���$���2��L�1c�OPj�;[�Y���J�@��Ɠ�����~�>72��X�9�L�� ���^D��ƉFݟ��[Ԏ�"���ue)j[�Z �Y��@�y��K��q��*c���������&�6����/�ҩT^�n4!Ce=�d�����+���������e\4����ft.��*&���
q�ۨ;����Q�+"�#ms �Xy�0w�w�����w	����m�@gMNj�<�`#�LyD�������ŊG�Cj�����jѳ-�E9�����q�i,�$��~η����p��PZ?���.`����Gc�N.W�j��Zׇq+�2G�v���R�K�q�5U�Cޞ�����cD1�S�p�8�9���寡ȃu�7�	4��6|$����~~�ʴ�7A�N�ay�	���m�}��I,�lA�#z'��;}hxEt5���Nd�F�d{���r'L��%���r��w�2�1�43�0�_}���X�/��ѷ���Ps�-�z������R��i&���Э�2�*�/c[��??�y9P*�'��p�K`�H��HE(���Q��z��h.zi�	��oq���|ϔ���y楰�y���S��/Tn"�"��I����!(�r�V�g{#�#(3e�8F��e w㨬v1�:�{�cV�%��/R�.�a�`�<μ�|����Rin݌t�r�x���Q�����zLk�ؔ�˨,U�C��;�,�:7�rz��hB�Q��A83��JubK+�QP�
��4he��UU*IT��M*_,�����j98�b��z��]�WγI�b��'���2ڔ��>:��8,���0�cE�LE=W�JS*��LVx��Mv��p�x@���r,$�{���Kw:!�4��Gɯ�nwR?���?
��n�r���å�ݔ!bg���������glk�z��_�ik���\�e
9[�ۍR�����1��q b���W~[+���/U��T�LIw���^��	\n-󬍢�}I��)<�_;'��f�iC2�[>�S�� s�T�	/��wOs��ӛ}�6��A�{�$�:A�ҹt���LfA
0Ջ���A��t��8�iղ��e���1��'9�Wea�����d�ُ���0�4s>��]��i�������YJR��D~x��Yt`��D �6f�a/חjh�%h*����7;��Kx2es�̺r�Ҥ0RJ�,�����(�H���a���sϭ�,''n��g��*%������g��Ʊ�U�5Y.P�~�[;j-��;zR����-9Ku����Tk���d\R>֡���ӳ�ݾ��!I	��^�B1��� 0����x�\�m�^�4��K�C�{
�XD|^�����(3� I�o�����6n��=:���m���ܯ��qƚ�p.pfPL��!c��	+�Z���Y����z�*+eg��(�q��[�F:C�)5:�,��}Ք��و4'�r�1��p%��F�o̸��WM�U!Ġ���b���1��S�����G�+i��&B n��S���N�$�1���9����r��$_��<Yi�G^PYW��l �<	|F�Yf�;�?���W�q}��])������h�-78�&�x;d�E&�v����<,u�je�_�[Zft4�pY1���̹�MD	�~8=Q��!��+�f�����B�Y �r�^n�c.�gu�U����Uܚ`qb�sVkv��q�p:�^YC�;���u7�ݐ~�x�ՂOզ9�7�J���7ڸE��M�e��[x��S�a��k���W줃y�Z��B�'i ��<4xxi�ͦ.szdl�ʦ���!k?����ZQ-V�iG����a���5���>�"Y��r��I��槫�'fV%R/�Z@İ�3$֣_�.��P����t�֨��E�Y��Ey^�֕�i��AթWZ/i
�#�M�Kԕ�l*BF=����Gx�~\9`�6��)=����	�Y&��1C��0� �P�� B�W�!ܽ6AN1��N�X�vHx0)�&��(Rk�ƣ�O���#�ي)&#x��"��i����|u�%CVs�m�e�����
��h�YVj����2�U2)U���E���&N�C����`��E`O.F���(��1��DⵁO���2ZP�;�t�����F:#��^���V�	�D��n%ȖF���!ݴ���H��W�א�%iu�U�{�b�����~[�{�f�+�����6{��ߐ�ZX�?�K $��+t#�&ev��K�S��j�Y)���§��?���1ڰujC���t�>k�� 2�Z"Nv��=��<0��?�����DhC~���Sb�8D�lJ�ʈdBQ�"W�4y�$��}����΄�-�V<Lb~d�to����^^q���3\K
ȷ� P�"�h`2�[�ǫ��8�/b�X��eD ��W��uȇ>��X�a��.a�R_�6��3ޓ��wW�� Z8�ߛ�bz����
Ӂ��HB�;l�YkR���:����9�CV�N~GU�$�<j�uۉde4�{�2{vlÿK�,Tm��@�����+��m��"�I3l�����/d����y%�?~:
�ǫb��~�1-���Z>���Ĕ<�ύ.���j뙝Z�y�/�|��֖�������wg���s�x4��L����	��|�5ƍ�ק�)�k<�CPcJ\J~�d�Mo����h^�T�����L_������h�FO����W���i�����2�]�3pѐO�A>\����!�w�'�EƜ���A=�1��_l��%B|\|J�:��;�L�ƈ��0��gY1\�׾)���]����~��*�b\��s~`3h�`�-�����f�p��d���	�AM�� ��c��
�y�<��[/W�{�f�6ys�`�$�-�'2�N�����o�QNP�v�- �v���9��<BWH	�4�1�P��׾IQ�(��C�?7�$z�v�esu˖�����)9uI��0[mND0�PO�F��ܠ�7T�`��n#����R50B4#��G�(�׼j�z�ș�����!�,3$�B�!����'O
�B�Y0��}�6��Vm�_d�/�&�3ap�C�i���[�D�؞ؗ�x�{3�$�N*�N�Ko������Z��R�FG�5�⺢�1�A�9�I���O7�n 81��I���w7x��- [�1ܤ�ei�J���	%-�-Y�iGp�x�)����m�W@�z�9���M��n�s;R�öF*[����T�`������/�(.u��F����*����JN?���B��ϱ�.F��O��ݸ���y�n��Mm)I�8<� z3D8@���0Z������0 16�me%=ʆjF){�?W=�Z Y��鿹�I����}L)�G���T�lW^���o7jw�c���� &��]�\eH_���W�]����1V�3��̈�YG�;������֑��W>W�pa��`�҂.˸����^m幀��`|W�8�B�oo��u7hU���B�\�2'�a�:x(����fT�<2w4Gî��s>j7��5�I��5���ȼ��_h�Z�r_ˉL_<��\�~�6����h>���i2����{��k���%#X��D�e�W˼s}�k{WC�P��
��;��d��.R'(M�Cr���*�A��-�O��B�ǐ��)��d���:7���62���l��y� �SeZ�c�=O4D(�H�!t��%�/���E ��7��{�v��$����zd�}�W�ĆQ%�zKb�����ܷ8N�]cx]�?� �Q@t��&��t��Q���Z��Ph@�`�54F=��H�L�r�K�ՙ�LYU��*53��g,�tf��n�i�<�>�5%�,^�(Oi	p�K%,�&ۜ�1��`ᣃqF��'���WB��W�ӣz��&j���\��)�C�+3��#pA`�ٷ�ӣ��	��Օ�NN!��4b}+�k�i�{�����X���6��W�`o��H[MZ�$��{2�����O�^��16�R��<��M#q���kyz���C���l�zY�i:\����C<�}g�°�(���|�k��5��b�ah_���1���4��)����&�a�a�*����`�0�@�4	Er�`'�Qv�18��qwWC��33U�h�aG��Z�;G��tf���$@��9r��eţ��(���F�Po���9�Q{|��A؀��'r�E�����<ǎ6K�*�������L��Y�t��� 0��� �+E�2�.��=왦�ӭ�s����ht�׋�����*���Q+�1x�:��i��ye�?s|̼��_Q:dz�R(T��g����4*l�1]V�*���(�4��E���0C����ނ��J����z#D����3��IufV"�^�!��G;a��ť���n�0��[�-��tL���},��)iʛ3�|Q�	��!e�n ���6���-�&�j�yG6��q��i�(�����-AH�J>[�Ef˙��A��DYח� ܿ`�?C���� a�Wpt�%bl҉���B���3{�XhX H
.._��Wv�m5��bT���[>�$�@DF$�l|~iDi��;!��w4�aq�&+��KQ�N������gtu|��fj��xg:���N�$;�tA�&��6���*D�G�������+��5?�����82�d��W�N����Vqz��`� V�̭ ��G��E��m��X$����I� 3k�nc�KLa�0�Ƨ�v�"��!HRmO˴��cWDQ��o�\�2�_��H	�ך\����:4�ìNKD�6�Y3�<�����&�ܝ>t����l�5ԑ(p���Ӡ^�������[8�(��ۥpP���()y���}2i����qİRԅg��ֆ���v��C�z.���,{�}�xy�C�N��j����-��Vt7Ļ0ӥ"6 ڷ{�5F
�;.�8u���;f���;is&}��G!̵R��CA{��֏�Au��.�0��PP��g 㥐28�9�c�Y��{�o�ӈ��T���%�/y>�yL�YY~�4C}�EYbϠ���9v�_�p�����ɹ7o���aɼ����C���2޵+9��X~������cm~��e�C���t����F��٢���^b�|��&��~��'�~���#A�������`���n.�n��|��et�ksS�I�<�/jϫ���-v�KW����
���K��/�h�~7��}8�nǷ����Ы���2L�4����XK�>EH^����([�g������R��D85�q�p�~dS�V��
�1����X�o,ä�o�Y�s�F�.�hm�ߝWC���qFm�y���g�|D��q�!s��3�1����3��'hLEE�Z��t!.�������cC��N����nǂ6��*�c\�gZ\���I�s��V~K�Ҝ-���q�#��J��J7�:�z�'3�4W��XP*����C|5��>Խb��]k#�,]��J�� �k��{�'b�z�o�'�n��^��{4����q1V=�v�w=2#!{B=3�B���G��
C�'[y� ����7߈�3�.#��܄l�j��H�������c�_�T��D�ʄ[s���LX��Xa�����r>4��H�hgC�04=F�h+Z#_^��@�����q��&O�!}o�!�+b	v]���#��4�XJ��g�2�()����~sѴ.S��&�X��X�M�=8��C8�eYo{����rJ��f�>�QѬ� �j��>��u��03e�����#��G�Ѷ�x�Yak�u:�����l�Xt�������!U����B.̸+�(����oyf-�����ج��Io��W9�G��po 3N6'����C�G5�a�~�԰c����y��-�9o�][��K�Z2
8���|�]d�=�����r�M����XKx'�r�k
��op2�?�~�Na��+|�>0�|v+J˴(u�M�~.�bDc�"'����w�>�C8��F�����l�U��8��|�c�<��4���}Q���[�fd����m���[a��Phm�z{�t�Zm��(�sd`����i��j���6���6�6�n1e#Z?�����6�Z�E1�0į����f:�BΫ+=?��o�p�M�n`���ķ�auR�͸M����YѦ�QVI3 n.Uo�W��m���	0���M]������yM@t7��O��13��.�w��\�^B	~4�8��bѼ� ��R��LB湰��������n*�it3�sN~>��v�fPi�`|M���HJ:���$2��Y�񒶆b���Щ������Lp&�.��]"%<��;�͇2��t�.eM�-f�ξޗ�up��LD��#�Rt&�(�����f[�M�`;�{R�
o#�[/t��j���5ƿa5]!��\�͏��D��AQ�)����,���+o��s���E�rH�9�y���"ZlR�ˈ�^I�3��%\k�
X�ʂ���~��&�ԕ�hU̐�j�#���Z�n'c��DO��ǎ��>�?�B�ʫF��h�,�l�O�=8\�����og6L:[����=B*4�u��e"���������ψ1/v5�N�?�-)3���:0�r��"Å�׬C������4�%A'��v�P��Q;��Ǜ�C�p��C�,.�xF��O:�t�J�ΟU����/Ѡ���85Ʀ� U����e&1f�Jɘ�!�y�j�N��S��ajv�f�~���Q�����b��5�\�����܀|FE8���N�j�ɉ��/o�C�����+�4Z+'�d�U�d�hХ��|����5n��WG�I��5�yT����T�uwTkMy^µ��Ϲ���-76KJ��*Y��a����j�}��&�m	��lJlk��a�y�/�A$��?�޾��KU���3	�6�fޞ�k�Fԭµ�ұ���2.}W�s��z\bzX�,KL'UH�?^ɠ�u�AK 1d+�s�e��pw�Q,5�Y�FR2$� �5��Zy|%��QS����\P�9�8%�_.q}�+�t0l��蚋\E�<rO��ak+�[�p�$;E�@����ƀE�6bQ �Ⱥ�Y!7q~i4CCTfy��#��h0m��p�;"Ҧ�K�,�zi��'�/���,�x��e�Q�_81�, ��s�����\F�,B)�Lؒ�,��rwÅZ]�62ל� 	���C#elru�HEw�p�D�d�l��K��5"�$'�ߤ`����Y�cyi��\d}��ف!�-��Uo̴ߜh�T��A|:��b���|I۟dtF�e�	�H��DKߞ��N1x^�W���	��bi�[p��b&�� c�G���oq�Fƥ��}������X��Im6�|�;:WX�4{<�����ԍ���S'-wW�7��S����i[�aH�H�e�0�>Z	����D̩��ܘ�b?<ȗ��	���W��nI��	�Z��+m/kZ���f�ftD���Is�ď�J�e��P ����&����MLY�x �uЭIҚN�q�`�i=TI^�%���)��?/�e2 D�l��V--]�����8�.�?����o���M�l7H�= ��n7��zX��^v5� z���M
Yt ���h����ԧ�~�Ѓ|+���ňs�I�WYmo_\]J�������+а��I�$1:]�V��z���օ�� W�I�Wvieؼ�|�����z�0��s����nv{�/0]c��]��}3�j�
m� ������#���P<�ڽl�� 0�1$4�2�YOp�m�?���f�Yrn�@:v��Q���e��ݨ�����=�S(��x$}'<]�F
aRzX2��74Ss���ejyS,��T��&gn�7%X���:C�{�*�[L
���UR��|��Vd:�g��u�ʸ��2U�yC�����_�i��ߐ(��+wC���傂��[�a�+'����Wr��"Gs����p��,z���j�ws�������|�����H+�bw��+BU��-�ޕС��k|��z��O�5O-L�����~vf�ZM��WF�H�X��(�<8��3��GSߥ!�C<tZF�Z˞�&�a��^q$���%����dP�J��j�UzP����cE����y!Z��>�!�.+������ґ��N;�-�Rf�\iք��=X|��.��]5�
�M)��(��6T]B�Ж4�S�HEz�Zc�]�\��E$c�Y/�~CJ~��+��,S�O��'��7u�S�q��1����g�q�A�}���m��8� Ƕ1��S�	�x��M]itkXv`v>�S|�`��9xS�L��J��`����q.D�eT* �C���PB��h�1�����j���Ps�����OĚ�W��P�0 �a�D�s�aw�V��[.�@���G|8� ��?�d����>4�FZ�W-.����q:Z��bk���ܤ��;����/kB[�m�'��X�j1���b�����nɥ��+ɂ����3MSQ��e7�֙������0��թ���zԮ�3o*��.�u���]/0�Ϊm(T��<8������.���z~�������1�����^;<�?�E�L�g�CU$ˏ ������h��5^�=�������aS�O�h���Kt�6��08��n}r�g���1^yr�\m2/�O���'teN�9�~��r��g�u����%��<VJ��`l�{��D(_%E�G]0c��B��c���a1
�Έ@"�`�N�T�:�h��r6=�Q��,��J��kd"��\�/�^R�2
���뾰m@���h �'W�I/%݌M:����@%BN�X�M����X�k���w1�t�Lӑ�1L�	}��$n�/��f��s,�����:_�X�.1�**���̩H��o����_R�h���4g��Y�3�ws7�Zb_$aV����ux2����Q�C�LϦ��8�CB��]���N�ҁ�z�h�T��C�Y\�������r\��ƈ_�Wܮb�v5�}�>�+�xr�	����d��Z�(���a���3@�#C�ӯ�bc���
e����!!�w�M1��*�O�-$��/u�6<���Z�ϫnwʚ���cj�Ĳ�d�2�"26EA�}�N��P����:{���a��L����U�{��-��4��O�TW���[p�_��8']�\���DR����-���>����2��s�^Y'��V^4�%���5�}�ydt6Yr��:$�~ݟ���ђjuu���%�ݔ a�$,/Ѹ�o�	�L���s��r٫,���	�E3�B):���v�N�+_"��Q\�>/�}�����Hfh�#���3�@M�͍w����Bt���[��aLi�S\Ҫ��]�憽����~��!I���Y�bN�*����OK_�Ѵ'��~L�zVf/�V�J�gX36ǾT��b���U��I�V�Gl=��t�@t���ҟ(�esN�>�l�4.C�Ě7x|CH�7/Uo�5��z,F���ࣾ��X�ve�~ض�.�|�K�Iiܱð�5}�ŇK[IhXI��L���w�0a�� U0uf�ͱx$u7�C�"�yN��؞LRS���(�tW�cŸ��[jj�}�!��#�E�ϰl_:z��f S�G�6/n2PY+AVr��`�NUz_y�;GRD-�IVQ|#\;�]��l��R��[qcO���6G���i#1C<�Q�i��Nߓ��})XJg�CtEm���D��!�p��!���_@�P-�D\C������6�P�8���J��nMѧ��kq픟s��~Dp:	��)^�,2t
1�w	�Bf]�;���F�qM��>>=�ժX��1@u�zz%�OӹХԞ7mW. �?Ӣ���Y]=�:W˅ ���µX�ڈC�x��*wĠh��g;��}	hC�}�	�0��k���y�*�$C܏��_�ypQ��Q�͸nB���Հ
c	��W�hS�_�3��bL����+��ǯ���O�M�\1el��k�ޗ��9�;h�Q��A��!q���[e_La:�q�� 9;��� U0���l�Пiu,��,-!�J�9�d	z���q���;��{�)<D���}�����hw�-��~�۶���a�k!5�b����)�"B�uee����t��9x��B��؇	�L��j���J� �V XG,Ɏ;�r�!>�n�������&�{Ɔ��R/<DO��p�L�����w��YX��#�S�x��b6��cGmЪ�f[0���e�a�(15ø/
(̤��Ǘ�Ȳ��)/.�ԅ��4lwn���%����Neу��:EZ��8���!s�AR�%�/��/�cdϜJ���  8:?�W�&�c-��*Ĝ0rZ[;�X͉ ��`߰s�!�b�xȼ�W�	nwE��|g���˽���Mm�����,}oف����G)�%B�׿��Ҋ���\������u6Z�ɠ���Q�"�ZY��"4����>��{Yhu�� ƀYq8��8�e;�b��?Տ�D�0(2-�W�2���Ŏ�Ѧ��lns����z0n�_"�����c>�L���1�c@I�3xQ9Pu'� ��x|e���+X�[�&������X�g�>���iy�)��2�w�z���?���Z��K�ؖ��&l�wBd�L,E�oz>�u���	-��Ʉ�+�9��H�ڦ�42��<kD��j���_y�S"��ȋx�fQ�
�i�	�
z�
�J�Of�ZƉ�,@@+����2�6�����R?=Lw�|�����o��#T:+�-��<���w��AR��99��Oj~�	X�H�A:x��]$=��"jX�qk�]����+FS~RM�5���hDv��`0[5�����Ы��h}-�������,H������P�5R�l���� ��4�&�k����P�W�^����~�{��b��=Jg.f���x�.�i�k`��Q�I��`�Wj850�G����di�8�,Fy'Z��WbM]��' ��C��G��0�l-$��6�
K��H�	�k���`�X%�
�Mc���ܜ~֧72˴�"���������SA~I�F؍���Lo�ڍ�|zŀ�=CU���N���]Ppĸ�9���f��=z����\�2O���t�g8@��Лe��Y��Z�]WEoR�A��A����<fA��,�Ȅ��0���J ��:q�a�;n������b,� B_�{b�Z�b�q�ŦcH�'�����Z�A1m�0�{H���K�q�{�C����3�*�Ja�_�����w����[�2�ߦ�u"�,��D��C�������%�gS�����'���#<����<����_j�.2E�J߀G�g��Ny�}}?;.&����X�n��
���+�g1n�9b#��=�p���U�'�
W���ƃ�6A��^�:��U��5��y�&4S������Տ7�6s�9F���6�K�	/�y�PW�,�
�{�9�N��-��X�@0*il%�$��x�>cU���1�)hv(��M�^v�v��V���"l:���>IMhʾ�M8�' ��	����Z8�:(ouL��^1&�����)�g^�c�e�Ŀ@��<����i�6���&�7��
$lE�,i4A�V'򏠳��QgY�E*�h�����̪בԝF��3�,U�0%�ͦ�h��$W���ġ3������9�H�)L�^J=.=o�����XyQ��!����E��8=%Zp������rC�����ڸ S1�z*�c��B`�2�3�m{��L4��3p֗ys.Ž�Jՙ�,�܅�L��gVI(M���d�Ȥ�>�Ffȟ����)\{� K7I�r	+�|^�/=