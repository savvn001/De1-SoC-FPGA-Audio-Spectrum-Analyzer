-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FHMxNUZyk5tUaqeJS4pObnBGmvfIPnWR5hzxijJosR3a1P6JXj4kOZwMAB5BI0Bnl1drbAdUk4gd
zDJQaPi/F3Be+0BaRqF6dW8cHzqRjTkw8KArS+ksFdCQ3bYQUyKFIUb8nPO8+SExlPciSIhSEwqT
CpO+2otWc4FktYj2UajZPi+nvt+O5qLWAYMp7wMnsvUYQ+yDRbw1QBNrxEtwUkzDOGihZqrj0I3l
9Gq1CX6Z3FPoeHEAmbjW1t8rGm8itFOo4fhqzTwOQY30IJPYYwOnHNj+YIg0Qirw6SF+3UqsFSyD
Cz4eC2eW7zovImjhZBgMbNRxr/GKYnuHc4NRYg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
Jo2gRQvYWDJsBR481Hu+O8h6Rtv0GWykHOvmQK18N9esGd28WDwtnnHWr6ux7P+KpNSAe+IQCxUt
c1KXA1xjGZum4gzR6NueerirAM0cRlgQWP8fb4Zjk1QeqXQvyK12wYwydE2SgtwwK6RGRzFNEjuo
QbSREtNG7Aapb1mkhk95IDX6KNFBEWHR1KMEnwcLqM6ZekXHQMw8caPj1Dik5CHRly373KgQi/Fn
+uWEzU7tN7ibJFSX2W1ez4mZAaHZlnjq/Bmm7xC4rUiOICx6TUXYnE1IIqKq7j9OoFu0GO9NCVlU
aeLIAjh5wHFhOYG3sRhdQTIlRLQuer5H0IV2tlz4eVK4rE1UTGci0+q+Qyd7jTRMtGnSHqTdrukx
H1KmoOaiCoQ4/487pbEwrJKseEJsbj37o5fXvv023TKltA46OfLaPBtBsnNQdwZlzGpUpJF7/BDY
cLeeXCeJAfwLtMc1UxBU8C0NY9JGSVyXZmy81+7DdsMXcC2/Mu+skrBvTCV/wpk1f0gEOuzI+73a
F9J7qrqcpGf+GagG14auJrUREf7N8tHdsu4EwY8PYrF9/qdxAIJ5Os9nRX0M9s/6jz+afeAzRTlv
InNbs1d/xRB7fTbEAvBWZAq5EKVzmGRd36PKCFrrNtJURNHS8sXU6qnPgOKO8E3FgoPFZWvsfLUs
8Q55vHgE1Dft9wNGdcCRpQGimXcnARQ7aY+v9PGyVHzT+c4PwVqALpoHopA9h7EaJsR6y8M4Q+j3
PegxwuQR+MrFtDtIoOb8px1tElwka9o8zy+r+on45pXWIG7LJ/ylyIF7YCf3hRXBJfXgiLBBHPdU
uLaP652aYm3i4ZFoVmAn09fA1ikAmOOa22VYKERYTGvUaqvC31QcKVTizdqd4j6fT7MURUBFD8S5
c9wMC8KhrYbyDHpXdN9QCuLBO1ZcKX6XPB7Cl5/edGbCd8G5duyphche4/yReQknayKMrm4vt15e
YDleBTr4415+CXB2LPpPS7VvjVc8PMYGCZHBI1tyo4UR15x0WBYVOVB94p2ifM2sVQtgIkkhc8Wp
zGOiGHdxxUt818XFEIUsck7090A9KF7HXT1sZZKcFvx/9GDAlT4f7l9jMslZTQ5Rl9uZmYJHU2Cm
cccp2nVf57we1l/Kb84GbWwZNCslTE0cgyQ2bi9T1z1OnkMk+RBPNZM36p/BKezXDLGgKACrE1O0
WDhkFEAK6w+tbAD5vFIGZC3i9w7xZ9SLsrSQgLD8G9bDGg9kuKSWggQK6/brDHTv5nU+Jmyfb+Xw
xdOG3uS2IxFRoU9dsLgy1pJL1s0Ec3CJPOCa0Cak7pf5/eD3F69iWXTzsxombaEeFndV4Ve1MSCa
jAi+mrVkt+fZBW4kgI+C6b7xSI9ypRrtUKfEx3WeR7IVoeDCrpLpwlvp5Cgo85XMHciLLBtH8qS4
2d+t+51J1YHlF7HKdxltVfQJlcKY6uHRof94mJs5mjK0Y73uAuUtJFfONWTADJQf9zPdSSMEBEPD
xwafsFpfNqS0N3TO3jq7VRwuHmszStfXzAAV80YO6A2KmQ+Ui2u7vuTIbsNUwnnVODgra2dEknSM
Ef2ePXmmizr45chMdWDJqFLnd1JoRy5UD0UjhR1B1eMHYznCPlaahJHXDiykM1tMjHA4vTGVSxsb
a6mfpaIdiGHIh3mU/lt+jx3qEFEp3tOGPJ5ZFtilP3o+84Wv2zpbP6qjYk9Llyogk3tygl61xMfH
L+GFp9poqU2+lG13olxUmEK143ltEHvdnhF7zsWqvMIkuH4b4YV6XoZYbhpDak08qOKDAVs46Vg8
BHlee+1T48ubQUeNvkk3VJ/7pKihAMZDw3v6KEYu2jNMnhd5/VfhqaExW3h34L/PVLZjaIoj7BvO
YKsayW2+f/r+1S/h/fMapmOL/Dordu69SVrEqyCBsW2olQ1ZB+QwqC1Sr5W6nQ3PaGZOt0x7x859
gLQFZA1dSXDLMkEbQWyA2xgTVEnY1Bv3Y+P8HaymoTxWrkJWMAaWmOP2DemWYnIeFieLUCWBBPqE
s+s9ZrHuMoxhGcE7T8eEIyplQxeBQIWKvehU3J2xKRw8+3eVTpE+ZQVc2UprWlJpdubuMzOniRW3
jR3j+1JrkV3ZSW/pnDv1E84+iIZeZLhkmuL50/Jv2sHjgp508CIJvhGX/ejqcGoUHAZLwjO2NXyw
HOsxgonpcmqdE+FAP9WQyGhXW8C+HQhdeGwQMzXT6gUJstVZjI81waLCQulhljcMnMRUjRWGi4WK
REJkvftcRBkiet/7HnBkueo/IFcRxc8Oxcw3RY4eMlEg7jSxiiu+BKqBI5b+PZU+YxZa3+ZmfjuP
JhPhh2KeotT1brDhua/ifNWvTyIjxjFSnbufAH/E6QgnIrePWhauKwPhAEZ5Ul0jOlioJT8fOQi9
jwrO0q06mbKdO8CXjkXbsS4L0X3Tr6QG0MupuW5b0u8ILkzEnJbOksBQXuB4GN6/XLmaM+8xAPdQ
55iVo2j/mNLw8FOcczVeBGxDc0b/3VOebgda922S01Ess/9u5EfcH6dgvgp06k22ZN5XUHkIgOUH
XwqASXmyGfBej5oKIuy0hel7swIqe85MBYiMnBYamHqylYEzWrDj1wY0S3NJjjT2vCRw+YEQLWyS
DqPL9JlUkUeEOpJRVh+Z6JfFHanHaxh2VMxna5rAAkBpSqVGb9pSPHCaBy92BwXwezltzje06m7T
HN2vbJg8PimalOUiFkDa9aHCMRQEnMFg7fZ9gQU0hWe+TRf95+iyPsU1CVKeA7y9DWMzaApg40RY
7shu9koIJa6EJDLUmYhkG8D5FwvkiShhn682WJlAU6YFavMaB+GH8OXkTU2pDtJOWEGz6nqPcO+T
ZUkzffcl8QM+UTCdtQBKnyMOs3CaUsHSVJHoPBtNKLT1VSIgBdyY+LAAt9tbr6mSOUOe7/JWgxsR
E+TUhX8+e5GZjFfelRw473keOb7ZOQl/aRQq2oRDoIwsvJg+Lc6ahwsfflXIuFU6dFzHJWxTeSW6
GG/kDhWvGvW0g53Hl6n3JvIRiW1NsBPMxhtcYZm322jhVOLgFtMLyGnbz76gg1QxcqGRVWUXF8DB
Yt0zatLu9OzKNVkVT47j0EFRNTAkGBph/Oq0L8FO4FbslF30prYB1vhJGJuBzZUwikCf9EZ5Bx/T
ECtvv8QW3d0cyQ8S9oqWPI2ojFY+qJZkx6EqP8GCqCeooDBxa+bkJR6Io9OCt600g2dmBXg9d9Ca
ucx+IoYi4y68J8/nO8JSYQrmgTmIok3MTfxdAZPQouae+3+chfN6DS8GBUJk+iFw9vQABt7e3f6D
yyrtsYTA5mytTVmV9+swe5wA1yWeKvODYbs3K1MP10vsyn+LtoaWGWa3tJjZ5hAmFYz8cZXM3QmF
ttee+S3/N+//ARmqePLlzzFcTELx9ctZuRGjU6sg7Dwu7Fsq1V8a7iQBSYZco+3YgdDxJAPxPttH
oF9GfceIO4YreI86uv5MtSrL+9kKsfLDJrPeOH/kZZZbJ8gaWKo0gryE6FqDzMFQEvGQMZCXssnj
g/n3a55ljCaDnAo0y+Dda56lp6JutFnZeF97Z32nEkY/Hecg+tvpPSUlyJlu09fMNO8czZgT5cLl
uWGa4d2BWd94jPiDWZLR5AGddPYFtLeCZxD6D4PhZwNq2md1ardFjHIeIfITVfEVfQ5SF7wo4jLd
n0aa/SZKoghK+huZ9OAoJrM0jVUV8uZKfRvHoA/0dAzk1BOj7NmOyH6m/OYplDTFb9vwBvYvmubr
FZqzVyDhQ1bMCwGtudsls1BEV7ZOZ27aAXanj3NzlCReT7dItcAlXYFtydPHSLBDtMFXm807ydW/
eEL8zk2YyuLLRv85bl9Db/TfKlRIURsANfCPsz8YGRlyMdDsADb4IUVRwYq/ZtKhaTLbLVtya25v
cHv1WLoKSAFQbx+6au+edVuarYqIBFrwaZxe7hmDkSxVepMkw7SUEtjVQ3y3EkWmeHaV4syF2w8Z
J8NfvQ7tVu6NF/bD0tuRYI9R0TiJ08M2vk/M13RmfR+5aYx3/ptadfhMEbZHMpprg6g4wSw38KRB
AE2kwAspGjX53uybFVl2Xy/eY1wzoTyNR5LvZdv7DiLlNv9QdQ1lmYn/Vtkb4yBkIc6xHq7pz2XU
7G11n9OpMWGP6QtG2ZIN4TF+AxTzrbmFW9qHCY1FRK+45rbb7tI5qVH4E17z4ZhUCXHWZpt38XRD
Wbp7wjhhQhLjm+zJbx6nfHNFr0q8j0J081c86bK/2ay30IwAlBFC3NrRr7XswNYhdQKqjlkjAmqT
OWMirv1Bmayct/SoT7K2+4Ep9zpSxctIdpRpfomUUUk34ZVWEDnaB2+ihvPnTfFI9D8sjhgPoH6Q
R399KDHMBkEqUN1zohCaQCS9U5PRxNtk2exHWAAQXsChL+zRnwzXCy7mUepImTY15feKUPfCZOZe
jxro9TiqMtkXPvuyQ8TzMSSIU1BI1LjQBb0pjJNINfV6aGZ9SK1S9PIuVQwq5G+hS6yK638LT0XB
KqY9O7NEfOScxbBqZzuLDRfQGqDk0kJfAYdSylFxcI3k5bOlsUPxg/z4TUWv+poguThP9oGBzSxa
jKf5dlQGaOxhO90j/HwPCcvS8GmKmFPVSJVEe+Fq8O/4ncU57GTDkUfsC0vej2bNWDj+JPPFljp3
sl1G5/vz3DFXmmI5kYB0G+5Xy5L0Nm01nsAs3tZbBUz6hJ109FzrtqqnJNpBGrV1+6haOKz60w9F
IYVZ71lYvX+i7SpoWpdz8Ux+yHWb1eHAGD4OTKavqmuzW+WKIoFQC+qWpyZ5dNaIarTAYcf7J6xX
9rTesYSIbieTHVmBe3HSGA+9ni7XvowOmgSeEMlYMZVMA5D0x0rsYN+4e8WpLRQ1S+CZRC5NVIKk
dITw9wHFGTPuEd7PXjIF6Xvr6AG66WiA4HjXd/2KH5tU4syL+jqvA99GA0Ej0IiTSSnh6mcMIw0C
DACWPgebn+2ZBAnyV+xz5FDmQTs36tNamj7UPzccFJIgJWpxdscb0H6ZdVYlEkol+Z7rIQpGmsmn
cfE7PTChq640Lem+F5xltkUIx1EamB8HGVzFNFhx7nt4yz5ZU7RePDv8hOt0f/1JJc1ucRlGEFa5
Tig4GQ5vkE13KZBwe19mw8lgnZmr0yQAf2PwyjDnA058/SgReEOxI6cMpK2EyUsGmcKMrExMwYow
Q8P3kbEC+0PjxR2xp9LC1GFVrCtb6Xs1oLjlOCi2PtZ0gBdvdsIHVbNpb8nODvCOmF2WI5IQyFEs
oS0qH2de160OfgmMr8yiUi1gOLAUXt+fhOOTrgZ1O3yuVZM8jYqlynazfVr9rD/HuWlo8XOK/u3S
u3W9+g84KDjaSUk45t7m9Ygdoo1dn6egQwb/UR4Z7qe/q0HM24SHX68Pn4xKFsRRpvFt/rxidx28
KOYskdcbNxtBImKZhVivhmSdMN9FiiZmT7WIZgK0Rgyc2YlR48kYbdmMrMeORnajj26BMxDxvHCB
Nqm8pdO3q2ZxJwzakm+gk2g/y4Lmul9XeHMPEshosC3DavWXDJT7zHdX9eKZW4zv1b6wu0xeL7ng
w0IdF0jrMtM/WF2hCn3qAvhcX8oUHc/cxlDelPC77eO9Krat08SSmAIzQVEn4in/pjn36UT28blD
BVksafOe3GV8gcDrXk0wVYFdaMLSqXNNN0rDhXzukXZxGbfWQBNk2jhA/GXD3v1unFMC6JHGWEbO
FiAQaNZWPo3u185I2iFtkgF9kBUcTrPnlYaJEWbceY4DpEtgevyX4T4LKUtLeX/ilWbG1L90mog3
Hs5CvJATj9DigrLQXCiXkmwJ7IfKZRuUy4pUIBMxYJxCqbLmpqCIa+6PzIEGILDxdtiOL16NsNU3
ltvWt5c2pznxwo2ThFcLz6HTAYOq2ZJXMJBdGjY7imvE2aemcKuDk3NYyZmtycVSNg2CJ94GfbdN
+R9yk5sN7iUTFxceZbM4Nkj6gmv6ISuQQ7CSX0IMIRqKkOk0JbGT7xBPBhhyNbE3WU4wQpEtnmU4
ozLpZVqD4nxoVdAmL4sUY/eGtxu7lky9dfvbWWIRpxpYX+36fsm4W09qX0hU+V0eDj6bnbNXXr9q
VRrZemy3uF/c8fab8Qvs8iDqZ79BeLYfF+d14pMu3LF5XC0Sqwm5x1S4Bg7bqUtLCMq+6EDv54KQ
CFWc5FOOLDuBRM/ibx4i0FkiRN1dnKOKdqvOEt0JdMg9woHQ4cBCazZmwz/IfsLYuQllh8bd1PUr
E2nDY1hZCLeGgGg3gTE85ZSmzfahsMAng2/6SN90AzJ9XCmsHm+shqpL4GxhklBukVhIfqgoZaDO
ASO0ObvYpfKLREtMCod4Gl/qMIfMnLKQfaQqbo5Yat8myRRiKaylSBDn7KkjD6UXS1vfbtz5Tcgf
h4X/dQ2XJzjCHgiyLxfgPIuSk+UjETMOx5uJAJ/p/Hq1SwWPEt3SNebcZX1JQJkx3OiGp4QUDZwO
Wbv7nQrQlwklrbPnXFU9JieiM6AEBIr3vGuLr/iaUZSx3ryvocaIDSITeO6/1/Zp0B7w5jEtWUdw
v6c2h3oVDAUBwAlPsg7YzgiBwsa9Xg9zuwXZ9XTiL4cZNFkEmPoi5ZOmoPs5Avr8tQaZm1bCYng6
aF8JL1rGaf45Kj0b84Tvq5UpKEWPOyz/MMK2JKm7zHdai/wBPlmDsdC5oFNlSK6MuoBNmod5Nvft
bZkmNbOaYzWvzmF076b+fNE9LgvZzRraWxGAo41GzKT+C4oPURHsaOtGMGJanZoBr2iENiKvupm7
ykgz2qMxFpZdE+i9h6aJ4QaxdfzAqE4PSyj+sfsypswNrpLuG9aLBH57K4yf7hYhXyyfUKpTwXOI
kmYa36B6Ea16VCa9+pJsM4MPRhmRe/KTtGOChil0Shf49OJZygGCjMrKpagY2CqD5pvhkhvgVrfh
58lpKV3RUkmnRpchF1DbQ8GP1VixqP9ZhOJe+1C10UG0Bd9aG3bLmUgxKVeEGw1KWB3nJm70uggy
ArUzW2AVUpmUvMGHfYb65KFBwHekqB5G3gFG6r+z8X/6gJ//HU4nF/eQzChty23tJqsIKU41ygWE
3xwOXxUC6OvIuF++XXJvVxS6o67tbA07hwkHS51wSD8z62MxMy5lcJUBOssmtWHfGiV90d7dZxJl
MSh9L+q1IAHtbkjeypPcJyAE75ZxCp3TzhvKYp8ss0M2DHP57f4nAz58MAJTn/d8CDG7eZzY79a4
nyClwJpQVjm187jCiu8uuKBT9RFZCN4QKfdUj2smk0IzwPds4taVViHDUwk7YlfBBSOzUspNF7JH
yq3PhfpgAMKDXylm93c4JlQDV2n+5R+bMIGumiHC2MgWwzhsVvxpb35gaW8NhgCi7qE0ALCKLQDk
9DPQs66RmrcIRSr4qZFtVBqhaAGgNNMyiwH7FplY8TiqpGUz8l1YWkWhvFnvnHrOQ16Zq2x5VK+P
rnqZwEAOk3SiSNuHxTca28DVK5WbnBO8d+DUO+MMIuhOMWDiiBQmrrTxELPfprxeZly9Ua8xAYGY
TdqSaEgnByZ2N1uWCFQcQnS6Sm/LZp34W7S8dt+TBoAQhxKs7xgDt4euU9UoEj9dDj+EiC3KQBBh
FKtXLjDldJuCKgrxx9ndHMCJ6a05ABMQbkvT7BAVv6R51qvFeSk9R3CbyySitR3vY9OPgNUNKi01
h5dgBFA8dxvSJYeu6lfADN+NHdI3YoYNQCi7wRUO+sExQkO4Kr1g0BUJZTUIbmT0JtIL0sgEIkCV
eWhPOMI+e6p2ssYToVsWRu4hwT8aJ1IJbN6kYvcWdcdT0qrcyepsbrvevZKH4aCLXd/GaT9SnYcf
tKBt2Vs0KhMA8ZtHHtYDmGUlfVJSfj5Qek/r2myRXEFB94nXDObaQHt01GMRcFyr7aL8JmT0/ybn
UlNFVFlHxeOA2izbGIWlu4GodZyfAtJqrEG9hxu8bnd1FuhDMQnW6C50AB1iIk9Sa6ThiqT7KMiW
iDoQ+1sEQUz1m3Tlww70ohR1XprT51OvFm9NhdmMnknYxNW32n3wqpI0dUw4cMzjKWh1uV0aEsVO
tLgIYExRjUs1qCmS69DFV931oY8nALnLyJqcvI+hkcL+qmApZenaf6ZEexFlB0hMaDkVybPTc6lu
64fuHksb6ohJXd1SpOM6YXBXr2yHWvdrfSDpZhZTmhaewcguO1HteiV9QQjdkx5RSol5CIDUL72q
/UtBfixXyQTxtrD2xrhCYsZUmfRAsTSuDj++QUCu/mEyuKr325ZlExitpq+yp64x31ef1PQ30lzx
ptkduW8gZmovWsuR0aZQEDw8Ptl9D3VnF5G/vq6R2s32d0CTo65NlOXLUxCG8H5w/iwR6tzylBLZ
KQYGCpfO4lW8iIgazKON5Fi1HIzp+RBJIeg1uSOAfXenhdeREBhGirCHHvW8N1swLlMsui68AwQz
H+SrNpIX7imN63e9be4vqowtI96cbM644Kcn52m1S6EqMxMHwf5ux5gJSFbn/eKyvpb06Re7Ktuo
TgT8YpHfBn45tX9AFdur1ykz5d8LB6CwmdVuBCg7FQhAqPTYp3OhCoZ8bxYag7ysFeN2NAMWXxOc
YH9YS9QYNKoNTBEzqYI4KNtzSONk9JptMV9njT/sNnvD6qA4WujIuzX2YwXT8PPgGRXSk7T0DZ7+
U7iHl5csl4cahmva/UL5b1f7U/a2iJ+/vcFTLOSvoQrOhEcUdf1MjFWG69gXfh837rffqSw8qrgk
oe6PB+VI8FukDJsizSTAC+whbVRoDvHBgpwvU9Yg8DQZH0QcUU8szO32bW/4V4aOPLdUptvrKjA+
G4/IZ528q+o247Lg+zCiJAxRiEM17UMkVrmOng4qOTnRb9c82EfcvB6seC1MP7k2u8x6VPaDEihJ
03VqSZXdYxXkSDyUlVzFpmWGO1s5rIkce2m53L3MqU32RgLJQHtxZCXF4esR0u9bzo4cMstDWB53
1hfVIipPWGKc8BbeXd6LdDmQU28sgn6vT2D8zTwdbpIorOvJFpn50aralCIOj0SiUQlEWI9aARhQ
SJP7i7jlNJr7Rq7irCm/NKWzo5TuiWB2FgW4lxvCQzEXRA4RJeqQAXPf2uuXRZlF2Ec/f9CBg/++
5gTxdtRzQRUbZsfvbLWtMVyEyTfyicH1ekugg+4Pwmk8K+MOSdS/Qgpxlh3y/Uygmq5hsHOfocvt
xoeNOD4Y5kj+fVyPWzgMONEAt0k0rSHmY7vEDq2LLWAmvWLwegq3fK3eTExOE5nFHMCbqBt+jvDX
gCQCvS/LMBZ4VLmHcxC2PvP3DLgNxvyivBz696vpj+Jdi5D9Ai3iVTIHhErQNUWhKDMkIPPcb078
hRCe96g1RZd2k6x4NTXv3jCZxWxq0aq/5HoFKQXFXwRqnPfTdCru0++nd9yiq0IL9c+ZYEj1G5EN
PclXmvGDPr4Z5YdHI54ldmob+JqKYMcTCMJlwwAdhJ0/mOkDh27CnkpbCvfJRKCp3E6CSl/K44Nq
hJw2+9GexFnvvSLYKqyJqD1IOJS7GWUXQ71ZnrJ4RPD+GMEqs3ZAKNp0kn221DH5HxdWqqJZ2G//
qgdqscUIFWPpjHFOUxsTcWGcoS+2UJ5qzA54cc9dmwF3anOLkUoM1A2hcXFzyLHYwX501DsMJgsu
QE1j0amJVB2834Js1tRcXU2bCutL7ejlU5wgup0Age3MTkm1jn/VL2wd1dTnG8xMiQFn8R6B4wah
M3W8p8VlNlGbDju7gSIvy8P6D0DKIpctm+M5JWwd7rwY4cw68Ua+ZmqAi5s3jfdA5BxW0flyev6q
+LkYZJMgaOQyjq0Ruh2dSf3kB4y5+i/9XhnI4WdrkuN+cyZOtlF1XFYZAVQG2ibscA6BSQ9GseUi
KZkvq0FnRodYhKtO7uNg0n2sZzy0Hg+PYmVj5aWE7CGvAGKbCwDyNjlmDWh6MyoRcyDICVomrPD2
gJeJMsafbkqVWnnfd+dphIP8heSZg6SlHxF/P7nMIGxxeyytRhTVB92nFGQVOGHMOL8cmO9kDc/Y
oeecL5i2j3ro19eVnwkdpe/3ruUxGq/2X8qA616py47Q0IyP508hvr/0Ad5tbA5GYbEFJUbYTz+D
THLNtI3eboP0yx58jkE1g6FYVICTz/XKCqaW8KBqP4ZKV5x9ARWZf3OqY+7fEO/nIa8EqgBx2tGI
jvOXCxPnellrfdpGvkSoHAxDLzFp14k3nVXSwtYqYHT0Vtk7VtjHCqbefW+VgUnUolBUkulRMWLA
N5z+s5vvLxk7uYpo5tBTs9zkSAHoBuXyTOBojH1MfSktihb5uLabxe6wpvhVacKI5rhiYgVqRw42
F/qYg45eVEJNORVkkXYxzq4HRAVGNRmvehTbpwwAEgLkQKcQM7e0+T1y/lCa5dC7vZvXzL3+NKt4
pNPg1KgHl1jRfO140Au6XS72g0FCgV2eIQ/GN71wHd44yD3ntzCpC9P9Pd0xkRcA4phMnA5xgkhn
bSKFackDQGEczw3NmvQOwNq53B/HfguvYydIw7F01Fd56EF/6fJ6yTYli32mbiax7zSs+DqIy2at
P6n8aCuKf25rGHpfPni1qS0fV4GkQgXsRDIceEgScN/yLF2+i77Jdh2UMoy9sokyUfyvyNtMfQMy
kctN0IyGFed4ue5zKOt57J8L2EEwnr/1KIeqi48AFBkREXdtt+2Xywxn/g5cY2Sfpbv5rXvMUeKK
AD73xjXtBXKlgH5kp1fMjfPZXaa4c1lZ2gBg+9g3fodDRiRbwq9yJVYUkpogOBMfo7UY/qg9xKKr
Zo11p9XRQoKUNYPRgD3tAFp5QdDcMw2GFPT0MMYI6khgx2quTvf9NgIqP6jz7Zxpm1Q43c3uHIl5
ePrFedZvFg0oYG1UCy0Px26D/MwjE5UoRxfktKnnuqX3DNOHP5QgVFB2lOsUDX2meDU3cMqY2uU3
KA+VelESI13oSvbegBawzn5zPXtEWNji+FlpXhcJ+edcm5whVMFgCEzs3s3oGDR8l3QYlPvfVsMS
r0YGwGubOqsZtzTPkIkyPDot0YC/pzxI8vNMoMMzeSPj90CF3rBd5j3L3Aq8VFuHZOY5hUkxG9zf
aRAz3k4dUfTYOpOA8+5tvQamjVdsdIlUjbXcY5XfI4z2A7coDcN/vWZGNxnOFkUqw3zKKBX4rTQs
TGYVX9PTa1NY7Qv+4XfNwp0CF5L7ID5K5l4+zCFRFycFbb76BD9qcV/bZ1GrK8emROc43SD2ALcl
2yitpsxdveBLZHzKSKoXh7s4OrDLrlI+Jc8CUjyBfUJGlREFJUrLKFAP+oDRs0nUQLiPCHmmZKdT
Fh2AifnVNLwRV/kI7OslBhh8XNaV8pht+qu+pQYFw5zahuU4ZlAQrpzOYaAYMX8QNZatab0KhXz9
5DwrL+/A7fMkxYH7J+Zm0KqNodn1mNHj/sTKQwJSmmii4N4Xk8QYRMe14gxYUEodt5qBkqICiJsd
7qPr2zkqKRklxQzOTTArQqVF22oeLLMYe6A2wiIa69R1EPuUrBw5bZeK01uTMeoSlesLKSWGQuFU
LSQCIah7Q+Bw46ohkwcv7kAGy2WLJEIq1lHDLUtiy4lmelzIMXHRjcoKsXYgF+rG22H0cVP60KXT
QIFY/YHlUURl5dhBSok7qRS1jaNRHo9E7PMsU2z4tYxTMpmPGhtNrNmOZLBs0H1kNzlEDv8yzKpj
CL0LfVY2bPqoThH9ell+dl+rnhwTgIGxOlub9KeobWdAdtIUjjWnAnmYEg0Ch26Uh/8N9pZUPzct
Gre5drRjAHNuHDuRNIlcccHtQPFn5pFJDJ1pJUPOdq+ZCATX3EI6T+5QBbz9WB5sjR78tsaGryYF
i1tQTriL9ROaEFo0VtIb4zOfyZfma2mJrsVACdUiH9TN5FoDjSCe0Dwh/t1oboCJSDUE23ZWF7zo
06nPLECUFyBrpSTz0MuZdugkaBKWYH4QeyXi66G16xTkbY8bX4ql/jjkm68CfBYskJ8/msDeZ7Ps
KUAUqsiv/6f+rquOwz2iPevppdez2Jp5Ji0znBkbwTaA82aQhsxh7G429ljTUs1LLVblDVzWezlN
a3g55I36Pw3aY1bv0bw1ZUDHrbvNvzyPwL1/5hy0k2a4dFQqNB74q/y9kiSf96B4jo+GgIojJjo2
TXGO03dTxivktELRlCS1iBhxZdBCi+oa37ANiovmhFVbW36qm131tXvJlkxumursHeP80Ce3LMMa
GI4Cuds1LcxdYl/hBnWmST36UPwfOfxwO4MrKBVEFYuewKnf9TdWO5TTWrUUYWmDKZyhRiMdKNv2
GRqEczzSwDBsaIUoqxxjSB1PRYjN22b5IAIVSxn3ExnI9+EgAORMfsKmOMU8ajSAh08A3Kbtr7br
km1/r3m8Z3+IvNKqf5bPJoCRM5jbfA6wesLdn8e5OdZxRu0qrQHGvA/ObGpRx1cXfurS0nqvcnpa
bJr+ojWwq+ly0mp/ECNmoAIEwg9xVX0BT0R494RDOZyJX3+U3Uj+f5XvBdA5DjImkVbj1ZG2vzhc
K3l5OTExsEDb3BY6rVQnkSOlVytNnTux/daGJ/vu20wuf95+TH5/UnYpNnBrKyLDM5PnP84a75+Y
HLs5wlNM7Ev1W+ZOyhdfQJnCU3D6bJEg2KCxP7nmeyUrZTKyjyr7y8fH1VhLVG+7OwJPoLcOIIuV
PsCbWcg6o68m9w0GihIkinETG97O1yFuTbA3jouJEcrSb/ml0bqu8tVx7kiEkpvM3H4lFiZrWHUG
9GmqUJ6TmU6jmuZZWkr0dFpasOxVXxbZsbpurUiLH7xLHrsjvxNXWZ5qwqJKPeID7YHnD33w2qNn
aW1Xq3z69dk5M4NSsIsOq7jWZ/BItHsNfV+trzgu/LI4JqWTCgLOTPK0vgP1xsMhRAAym/xYwZer
BdGFzQ8p9/2zuN9eqEsDsNJUsoXdCZCePV+sECxapOAVqTufzuehliXPuWRYq7SszH9MRpl2nibA
OfiLc78lVuFLVR9RdcOn+nXNk5RGa5zWy5FggDpJg5WceXHbjKWsYelLwTGWpRXFVKIpKZSsWZxU
qjnxn1F1d6lULUruHZTFRJF+jRysD1ZS3B+cWE8DvtHfKaM3miEXpztxgiHhrbwt0Rv6HcjkmIxS
UmgNo74Nh5JvHnHyMFVnPhEs8v2DLp2Pt9rYiS391Ka3t0qdJOh2gN1th6eXEtFCVbT2CydxAGnB
/1UpE6UiMoj6TcX4P6t6FH80IFhxMVY2EeWS3mNMomGm7WCyzwxAoZZW5FKmYzGJmSk7W2iOlxni
5u8iGEOPA2RJRM3EzknAqcAWJ4oWkLtKZPEikt2h729UjYkEMRE4huRvtnmPlVvaAO4Q/JbgGoEY
K6dgscjQMpYh59mV4q/q1FDEwQ6QUqWthIHl7OTbwPxwmaQIC4AIyJTU35TKu/l2+Ul7Mpc6cc4p
Y1zl/xZJmK778168aLpYBs4I1ydNsy0GI4G1WP8zme91PONYe2b6J03gCByxorPTlAYvWJtJMisu
blMsgNCXmIY6zncPldZtbByk1/RwxBfhgwVtqzi4cZPGpUtPuNQcov45ZXbIqSUkujm/YcwLb+Wd
K+vfxbRBthzrwSCK4MtabzvFdO12lFe9r0jheHM2RSTvOaS9jGuHescVUh21GTldJ5nWdbNqj7us
0YwEhZp/QQPNyvLXt5kS3DzPj/EahsNerPvDW0e4cbyj2vLCyNGsyMLkwaW6NsuTwq34mGBOX2GX
aFVGicgi1H03gujbJs8mVb1EM6CrodicN5U/SLIcuii3izvB5duU43NzEDbMbJMu2eMwi37mmYLW
EetVFGjLl9ZJTjDh6FaDCuc7zqltovf9a8zBaEOAiAJH/ZheEwNTzGkizMI1wUy2vGuC7nkpqCfF
AiXzJTkoB+nNDYbEJxc+nTGCKw7ikbhpnV1q/jcy5/6Vbats0Tm3W8qL4qNY12AL7NEqTp06f0AJ
S37Ga/+BsqbZJHncs0vBMVk6BUZmOKAFa5OucKQeV/gLrz1LXXYDNathKQCtrJlaI1dPgLBw633a
ySSXJSCapwYTQ0B1YnR7HZlE0F9kgLZr0/kXGvbloJ64vhkdJdL90a75rT2OLn5913FLSouLChXa
XPWoUt6y9R9GeE2SawrN7pJQL0w3t6yJzqJOlupq44+e2fX9UPlziJ5xeQLwyAMyLbNexEIQnuX+
l7Wv5tz8QRQdGCFU5m2eJotJVS/MqUjoY6TrUu8c4JtEZ75sojQCF8mivNLCY3JGQ/lyo+Mhc7sw
sSbk+BHQzxhmOPAKIIh8GOiTd0qRo9Mr2oAJUORO/qVVYwVQDSjh9WBtYNYd+KawMVA6iXHT3Pge
EqcWdk55BcDxkneqgj7T2SX0mzSN37PCVJtXP8JpujejZVzWqUWbxYP/mQyaZYg3g3TGEysXWg7c
cOnJsE1SET1eZgM2aDt3os+jJv82alG7AyHdF9X4lUmDe2GF2mFWW7ZG1L/hmZ7ksCjrmgrjRvwY
Zc9lpky+BnCoA2Hll9mzdUY3E0Qmq0eIdVNSkHKJUkm+1P2HI9A/2sAXDn2vCMudZeTtivQ51v2g
8tReL7b1geeGcqCwlO6n8HX/MqiDrBY3EjvQ1Kz96f81KtWfQi1xNGwbWo3Nhp4whvYAPp06ujVO
psGnYxagXndaKTZ8xYkVJ9R2iWGHBT6YgXMqrOcR0PSltPY7aSC8o6gpE5tvcha7lzDEXPadBBl3
hWXcvSdqiKOcOdKFpcyn+hWLFWc0InZthUPP3RngE8IpnZj/fJFHhJ3nfZrQhtpn0vImDcGJIrjM
ezEErwfD9yGOtNmQdZxxMlKaFrKRk7bAi2ORtiReXmFUFmgoDr79sMuQ9IpX0oVOWXwyo4/AJAo/
0BiXMK7miGS5fIV1gd/MGlbDFr6x/Fz9Ozbxge+YkF5de8Dfh+5WVziO3h8/6m0KLk5a0l0RYf/E
iTdep0PGgcB98XAMv0cpnrBAeUfSqZdz4tPadRjg0wURPgGKBP/UKp2MdVgIwQVwmDq1JTmHlyq1
00iEol6hWhkjfSxXPI6g//2s+AXSb+XQ7lbD7SnVnHleZktAjoTuHWGQipaLv3U4qroCKjzVROcV
w47BOG6k19HlXzoJbNK9JvbkwTI9PiFyd92I0OOWq8I/CJCm4RTm3ro0v3kCWUPcn2FUfK63oa0s
yigIYbov/ENqWp5+QioYBKPecfHVSBhhhvsTeUR2pOpL27Z0V+d0a9H4DQy46y1xkzWG59bNgrLo
wTgmHcOCfY0wknVyWstIN5sTQvQhFhY3IbAuLwAnW7HiWpFE4lx0aUrqndMowk7LIdX7++yMLRrw
0jWToL0+mRqVAXFYqUWCBNik0fhbhUJOgbtHoymBoSIrK3052cxk/vns0082oInI1EMSp1PZZXte
Q5fkBzo1HfmgJQn11VWYcM1s64LwRExr/Mg5E3ikBmkPNyDqswupDypij0pVITRKgYlaMWaRF8wf
v3sZEsVCng/1ZEX50BmnxPgfBI0ZR73kR/nSha0A/JdXhGbZF576bXG83NOpZ6foffl3awAfyOkq
+pDZOchpE6m5d9FjUd05b93kehxtXtglkFlE4pmw7G88krDh+Ioc2a2VT4qDa8H8eK5tkdRH4rdj
HK7qYCPBhEfKiB3aI/wYfI+wkL7xeVXXBfM+A9aMeOEj7cKAyFUhMA0uu+C3lD4Xd53FTMpdFro2
/vV5GiWw0M6vXIpCP2AHBtIrqHmVYEzxFHPLf9i78rjbQ1shHcvw7zT755AfyouFrPWapsFMMn2l
BNzHHifXI8v7iG0LtHTLAlp+HlGNcryrqDWgWJeKTyb/lDaHqSnRUKW5Zq1kpx5Gm0Lh3N9oMgzO
KAYVQUB0eNpHCd7J9i2rKa1YGUseNjKvICJ4Mr+8s5P4VItCs7fCq14awserB/OIbknREY4lE7wQ
dtUwcCM1AYsjL+D/kN2SWtCGvpeIsY4XjBltlx6VF4MmAgYsGXS8uSvQBqd6zFQ1bcRFDaDCzh1V
pCZOsA/+yotcdRPW3aczhGmjE8Q8QzEd3AAC+6/x1AtTo+GDEb6gKYIgrWcNBOS+szj1U5Dmm0ls
LlErQpStCL6bdUpGl4G/jCBLKB1ebnpTvnCoi7saVTSnKnbhPFUR6d2xa276SmBitcLKPLL33mIT
koEBHGieEN+X1GbflZ+w0/9yBuKSJfdPQToKQvfIkQF5lBJsmmjb2ziRSgPlMhFYDMfRz68a4wja
se7pmMSL/FeoBMuJ04JzaNPHpPBQHfGCG0zldK87WgXBv7OtSR0fKTdpXto20p3psI7KeNcLcK2U
Ik5t8boEaHLzTp3dhbe/93PAHPdWdjInmR/oXTHiCAhmp1F1gJ4Yf1CedT+/LtunHVI9iRbhRlkE
wtgUyaG55SSREg8THuloh3nrJHgyT+mk4Siib4u/lbESgfjzyuK5WzxjbQijwL33BMhktylMQX+H
hdTdaqS/rsXE+9hoK5wiKfRzGaJqMHypE2roaMMIhKiftrhPXdUT75vnsNAiPc8SL6DXgUIH8mhP
wObjlXYcEINT0nC2Uic0DUvz8i63b0k1tWLcj4aSgWMWsRUh+DVVhbjiO6gVqWeBf43w48SmsZ1p
RnP6IZbMRDKQzMpWFBnNcbDlZI/8mDShkAyOXoYxRBDsgixSi+08ScihHk0F+Xn+gTj6WN6fyCGo
GLUwb4OqsP8Gyv5fALiT2dRzUTmAI5J5Lu/0h58e9JxA6yyGqYJ9Ln6edFq6gaYiDM29DwBuV7Z7
gANbexW0ERF2FhbqX6rALP15zxLm30VHp3lKdimFyskgYwmORZ/CECysj1RdVxQCwcV/qV2R7tj4
46CxYYx8OvvGFdw9Yp9rjR775QTvaX0uUzzDf9DqzLp5Az4VF9tpzB4dHuaqgjbkljxCrDgxbnWS
4d7l7XpCMaxMxzUU/MyYUF1w3YAumfC1N+jbvZXeMvxfPXQ3DJQNVdxBsxuzKqQeXBTOs3bqAQzc
C+ehuT4eoOgYIK3ZznwZNWyIZ12LIXipJC6i1+B9iEjTIQpiSex0C3N7YO+zc6d7v36WBykz4roR
9esX8jXazrj6mVCuQYVio2PaEfSYE5RX0i0/8AWvEoVjP0VNstsWvpY+WtpTd/FvrLrgsLUbabGX
jMuUffSnz5so3CD+4NVgSpK87GluybDAS+wULK3UQcpl/zfjkjgk/yL7gSz2vZQ/HtYUdmPKWpa7
Xb174w4KOgtb+T2PG3x2qbC/i2CRaVueuT1bLyzXUTvavjH44WINn9GW3qREQ47OZh8e7mQRhQyR
9bvSJiOTKjbNQZ6LtW/Z8dn4Mh1t6tcDblu7PcX/oD4W9Af6wC5JEqKBwLQ5bUWm05OWs6Bwe+Le
FfzIvk53qUJpm5CjkpoG9i9Xx4/0pD1tPDRS3dCdSfVm9o1BdTl8eyNq+LuItOvmBGXMEjuadP90
K9cY8HF25M8iGaCRSc38w9ZjqRpV0qESiM7cWHYCjlaKMd0kC9dci2x/naNwxhOe/duIlDOZ/PPz
qXeCyIGCfqKWVKRKRdpGR9ywx7adza5Pqk7stcpLoEgt2Xw64+xD6gVuwzVft1wC4EpukJ/R7bXr
z/RzIXnkOJ2d3JncrL0vFWK7XqS1C4Vf/LYvZr74VN/me+YBsn0OMexJdCMVKXeJYJWRlzT1JhDy
FNGjptnvVBO3GOqS3HZZX02RuWlA9ksvZ+3+djgTK+jtVvtZkhj1t4QO8Mar6CBUAc/gSDZjk5K+
w8SDXbbNZy51l1whYXVorrakP11EdIvV9UdJNyHIx6aJFq5fwOvJ1vSz+m33sFmFSifFNY/5O9Dy
DIzU9AVz3w+rwKhGAVFPLlSImx33CdR3wqKt1NPgxrdZ1c6/+LkSdQe01VI83XZJgaWMj7/xvb6B
ibzvSTwYcvIYsQ3xoqHf8MvfY1JDnDv6+mndk1zElNDC+1OEP2jt7l1lJYK9HqUE4fz0Hf9c+rRc
TUSOjKcExKu7XvNwDpA7dN2dXqjfG0wHMzdh0FBA/GPMEWE0MibxzMuPVVjIclvNfC+YW3mUJQ1X
oSDNIKj3rbLhWYxJlfBtZMsaj51WYw/lI0eF11GTw21xOlE+BWDjrN9fcC5Yc8qc5eUEMbYOrDmS
sEAy5c90HY2gbfpakSxyCjApeCVDFTGVDNB8MxWgrFGdo8EtS41SxTqSSHNt7vN9azWierSulFgv
29tganINQe+mqJP7DQLDhFrF81hu4N9vZ1aS607VLXpkWASONbMsQhYGz0oFAtJ0iSDPm6VuIUj3
gAbLUHUSSb/ABqC9bLa1CIeKMCo/Me6YxK8PHmGisL9hFUOlTaYOKkLLe33bNVT+/5yWtDrAIrWW
xAryBQh1RtRmByd+/8TJLWbAeJ0BpvWH3YDNC+fdbNc6Hx8FP2fqWi2UZyavc54tmqe071c+UMx3
JcJeLohTnnq34b6JOvCsPzyAQ/Quj72uPX9AG0hbrHzTzlKmdrEdJON0O+1cGV52Dm+l9N03eeoD
6yOIqme1TYkRsAnRg1t5T0Jop6wnpIZi077hLuM1lSAABCouRNlPmEv6vXSzwZxPThKY4d4qZt96
WZHJwD9NppoGeViebS5usm8Q13ZAjri5mUQjQkLEIdFn5J9s1CCc85ZM7um/xEMI9ZfJjUQJLl1G
oRw/yox3rNWuLNQ/QT0Cqh2G9EPx3FUe4sgPXJlEr7JJk2kPiNcv6aIwM6zObKfzgTXkhNVaibyK
2pBpZQLbY0XYI6D8XIZJWxzjGD8JkqJHARPIBeFbaq3Xo6FSCm3cTVtFinsGtai05g5+OMKa9Nau
SMLgGjbLMPeqqfyOQIYP9NUNfjKYi7NQOACPyoOdsDbdPeWoBLA+oDl815Oq5MKY5rIywlmqbovW
821oOD0gwGKvqC0fq1p3JwQrZBcdcFY1HWbgdE7tayq/M5GPeE9U4pOKe7GOaZnS69y6JnaEreMz
3g4I5U8SRVcr9Nv9z5qubcil8l48qzMvBm3b83FMSCskilk8dvut93+rzPeq/CksbsuhAHFyXu9k
xG46yE94sJDkvNMCZ8Ob//gCkFwvGQ/xDVy4WYmcbRKa1pMeKx8zo1/p39JP2m0ir3saP+kqqkyx
eEisRj8sesCkuWaHns1p4NkaX8CPNNwCRbr9rX5UP9WZkv13Ha3wsJqm6lgWLC+EkZpCBAi5JpzD
PO96JUbbuYbhDwx5px0gVd1QMpJBV+fSdIHqpNlzMe1cpsP7kzUdpGdwWaS5DvvPPZSxH2ldMfJd
ozt5ajcO5ccy79xZSMQ7GtGssPoPY801PxGXGHFgdtiXFwT/XNsuibzVZUHcujNLdCiN3Oeob+dd
oSCJDKdIFKhFRvsf8GchR8xianMzIYKujTFvWlN3+D+Rgj24GTtoBzFwO9CgSzcxDM4jJ5/wouc1
fuFY9hcDpYFlk5pD+Ds6XGT+u8LYqjCucjPCNZDazIWcSs9+7O03oEWZxWveWRBPJkyp0E6lNNmE
nJZLf5DXb0K8BNzkdof+C2evDNy9j+WcFKvbmBtJnZ65rIfGhGncV5pMgt+agXEl7JDI8WuDX4aP
AVNfb0iCNFOu9QtgXf2YeBH8Imztqms16AbvLHSJn6MF6ulqOyGsG0P3+b3IwfsiUkS7YmuKw7GL
mG0z6aAGxSflMRhpRZeXek9svgXn7MZ3LsmMmh+Feu/XTmF7svwymlQ62rK1qj+i4ByLcx7KC0OA
fG2YmgXpLHTsTC6IkS/n7MrLRaTN4By97eIit80O5BKkce7EGuMQyQ5Xj93wu9Q2z0chSCXHa2dy
fqWJXnvNln5PXbZyvPXE4eqn27/YoovdX8CifIjkBCVIepEaJwVlEMNl2qfa+GxCs6Nt6GDpl7n7
uD3Uy2Qyac27NrS1hUlGGMJ4UPoGLg7uyZqd6yunyVFlk6SIVHOGwDPW+vEfgf5DhEJ0KQwhBOHw
GdUvz2e4OQSfj87iGJE+SMvP6haLre/WrkKz8RMh/bjWvR34ZcguMGqh3L63upuOCmEr7DNNiYVn
L2ia5R6genNTJ9dI/UqJGKn/SlaTve1MDUavhoUSOXqYfhwLcEv63szCqkG4Fx6bkJq13yZyZdPh
Wty628q4uB/810wpBS4TtOtLHYdILhdzp3fgp3WSTJG0m8t2Gt0J+RaUf2JSgl819zShZ2MXHaBb
Wo297Q+TDvm5kkw9CwTmRTH9ODRhRygGaz5sIv95ZAcLnSeo4ADZZhcHazss5YvVgc0Wf8LthGI1
AcsZFiekblGCdmQ8QS/HR86VHfHAm2QzbivCuZfaWEw8UPIACZsZtDTbq+UohzOfHJlo0MqtEB8w
2S+l4DDK/KYSQmyt1skXXhUZ5WPgnO6dkzuzhSxamAWWbniiazm99rud7h8+Ee16ESHEdOg6cJVa
Fd76CnsuMWHzL1/+0dARMMixkKz5Hzh02VEyFbyJq99a4jZJZXTbvifiAvhZU9Lnt43dJrGGNhMB
/5jC/Tq78Q8NI2CJ7VO+nQihQJ9o2Howysqj56NwVHo2lus2rA8Zv+VWhjpAZ/yHK8KHOOHcsFQS
TRlIWI59aRKXrirU37bMZBXyKfPYQ4XaL/PDz98HsD3CS8+zvj51E8J9EV1XsWxsFNhbUwO8owxC
1M0+CbwdLxCZjUJeYmSWPZxys7k//dc37myY4Uycep7v2Lnm1n7KKiciVTnzj802SEnUzCRcZorW
qHn/CXEPB96mBpWxoizUIOOkYUCz0cj9u6qYGMclGAkNsJzBAuQrN4Hkh37kGOYfFgpLAtdZYC8N
PIzoS6NyxG+sU3PQCE8QBFGnOFU67w+V0QLHdnOtG7lMo3SPkKyg7dQBhLyMIoDXSD6EV1vMCpFF
dC1QysTA+eQ9ugjt5XX7yynnbUMt4W5Hm3PqaI/PUIsDEqkPv8gZU3led2LEAKaP4KUZBNXf2YoK
3F8p1ITtHR9nPb37U/adB5UMh+7En9qynKLcFgkQCGEd3kT9+gUd/nOQdmsJbBwvryh8rE1dATng
IU6O3Sf3d4qDASlIcyTYJ9XJ0lEq5vezjbSI3fh0G8FdELBcepyYawaKpBiOF9mkYVQuSbGMVsBO
MRFY8UE+hR5BpWMvnPXMONAv0SB5noGdAKv4zBy5Z41QjSfnWf5lB8Jk8TfaP2cfALC9exvBV3Af
3V5rEif7+DWBTv69+8vw9IoZkxXb0MXvN5HIdppENf1YHTZ3FjJ0lnP0LUrKd154cXjSlt7Q597a
4d/dzzizFNq41U/0Qu+UaELHTuq9sSpZEo2HT06Jr6edEzv4o/xAyJEYFsxtjTu5cQvKSL3rRmXm
uuzt5gwzm6aww9UFLwV3shnFOjUyrkORALywkve4uXF+YBa+tx6JXERCJMBJx3QEFPL0NFwDH03D
s6D3dnYpv26Z46cjQ7I/1qVLWAzW7y3fpFuajuV2U1PEX4ZmehF6YTKxlVt9WKB8XyfdHdphTQkj
O1qBiWxkQpnnVIISqm5Zu7NaBqeTYE8kaMWBjlda424Q7O5tE0w6sxFaQsmudX5a3ES2p0jSXls5
IGPcCNa8IQCneI+gcUl5ENmmaKSGRPpGLoaKafC8szZTX1t+yRF+R3HnEip32T9DRIwBMxkS+8iW
AnrllD4ZJJ12BGmEM7vB0oI70O4543rB1zffyDl7QmvmHSr2EQssfYZxuXo1OpdXCUr37Z0C/p98
oT1S3OvfyQdKOztK8oYadFu5hYiQv62luKFgf+rUztAbTOecX4oLX7r9iHkxFI5MhJJxbPOM/a5W
bcujtV+aGHADw7zpV1GNI8gpPDfQQPrLP0GR5s3DyhbkXwxcmQzcnqPcfqoCHUj6h9NhJ8fcyYk4
2tk/y46Vk0/rLQyBcjykZZk7cnwlH75bYNLMJZlb4vIe73wNISPWtNM6Suv1j9SOVJ1/mKMqrrm8
tqlJe98XMnTnIx4Y2uBLiZ0vOTzRq3efYNZnQSDklCkyPeQ6F/96cYya4Or481qbTFuSFACI5k7y
1e8TtMTVjbvpI64bQ0mjZtNRR5UCvXSyG04fBm9Mf1ZyV1h5BGFiJ+uDFhhToUKvUdOklkbqP5Ju
9EZXKShrrUNymNy8pS7yuHtjac+CYMvKAOlo6nZw+xpamxgulk3TLRHeO9r9VFlNmpSlaP5b7bal
L8ilV6oQgkuQNaEqkhuA9CXn0wqpkdvVi40Uwj6XgFkvE3TPN/jwaFb1CT+iVXrK5iyri7DExtf5
b2a/4fqJRaqsROXZPNzo295Jepg4qvQEVj9sTTYkUWy+M4MGCXlLxcFVeNvocmikT6xzUPfn8+ws
8BqNJSOdHUjpuK8d496eOXuW10p31wt9xWMTTIxD4A4EeShZVmmyNFU0Z70EoultwnxFYrVmrGfx
eR5Ln4G9184kLLEdF9jKrSXmYM59r8amAxQIH0PivuzdeMyHQOwyfHUoGsjfkbac1TOoBXHUr1hA
Xuay5+3wctUlqjE/G+Vqw4iWdzmOcxSwtkDEh4yrGaC8VmIPHeUSK8+BTl0bOiPTnen3kIRQRlN+
RnxupQiUPy5f0EVsYGZqphD87h+3uCnTrqETSCtDHOquEHGwEDeKOMAA+WL7p5Rd0+2g3/1cQd0l
JjrX7kp2IByRNpC9KPRcBGqT3uvVbXp61aqe8awYZf+JDAa8Yg7PKaDONa5dur3J7okEOmTa7AQq
O1pz5gVIlrqCTuHeEQlFk10PUuTlbqg7QcciPlkgOuQq63LojZI24pi/cwCHjrvkdes1HPO8i2et
NP6r2oDCsCbgnO1mrcmo6SqrnxR8v+gK8vfqQvm/gZs4Ixd4kN8ywwORXzj/tU8xm5HG+PmoAYqR
T05ex390er9FVxXYY4SbIVR47AjSa+wUtSXJs/e4JfDiudShKoInO2KZ5SEWAW2iorNLS6aYdhTC
ZXscAQnEUHb0VOnk3n8llSKG0XD4qEgJ46AbJkyuj+3cyuH6vUL1phyJnqYttOcgpVrEhxOwR3h+
C16H9as+J9R/SQqPOrEX5auelQw5FfgGb/oPUqWvYMaDE0ZfCihCDiueDtGkNjX3hMabcwruowMq
zwBZjS/4bo7uACjfyfxK+RzUMFuLKEyfFLfsyGtdbRXLGG/nelYR009M1I0s/8x/ATV0e6FkG0TG
MbBZXrRTWKv4Et+fKQgYHrc/1grQDeJXNFoZRvmDXOhPgPea1iupdCnzAvtd2Nm2M+CWwBZYwsMr
1rZ2PebDISbFXoPTjz4eICYOetHzwTIhWue9WArUz7ASF6YUMUgzyh6TbeC+YpTKoqeV6ZmzAoMA
M/b0EUnGB5YZiPgfkOhVRBwhtnlASDsOMhhvfNA6mN+DfuQU6f1CrO0Chz7jlFnu3WSfvnm+6feT
LJSiTQdh9AB9qCBCgIKU4wgoae3uJ14ccB9YieIKPKVeAVRi65y4pI1ED9mmYTnaHdsquDfcNUC3
zKyUqZyFEKOPewz1dZAgEWXg311A/nTQw/OewJ9jhB1Pqi9tEAMPavA8XW+0jRGs6Fmhz4u+72N5
9hjyskinU3Y5T0cTkTFjsutuy3ZlFerPe4SaIUy0XJPIHoouZqFwco2cXsbyr8rLK11FNiFAdA4+
MH7T06iiw862r+3lbg02vCoE4u5k1E/nvot5xe9hex4Y8VJHOg193zGsvSU81tlYFrLIOgyN68SC
QWzChk04B4RQqcMDbFGFCOMitIXSMahJBdVn4g0JE6u0Ht9A/D9dLydhGvsy2tNbwIAkhNW5YdOl
8ghwrmAFhQZq7jaPVfsdahAkWP5IKRIHZmjH6y4t57/s0Y6fKpsAXqyotWzTWK3bXze5UHU3oAo7
g1l/mwJhgmjhekTuS7wIdgL2JaiUTnf2F/PP9CEmebpSh1vJB88wFL/iWAgnAs4v0f4VKaWSdS1b
x9JEkD5/3hFOkncJP420gq2EMTsCG5Y+4XH0Apmqc0dy3hUll2Ws/F/IOtDUbq7b/IE+tkwrfe1w
2ycq0zdtwkDBiL8sbpUFtAqmZ/AX84x04Xav1MmyOaoVZtT2T0FDY0iOU3xKpSFxHKEVvXMc4p5k
W2VgLk/Jqz8gBEKwxa4kMmf6v9MEop1BX9JQgHnubdvUxDFTUBp54GBerDqE+JeLL39BEI+yKNsL
PyEG44XWcyBtxVwyVo4OIR3B3OQQy2bpyumyv7hEWI2yR0bd58/6k+Geqw1RZuqjgHvla0Re8IhH
B1XAuS26ctfR5ve/Ux1AsnHZocvo1HvHA8pdX9/ZFlJEQGaXdURimNudqkJeF3Efh29irMrobbr2
X38f8R1yO9QQlkGO+TnXbD9DoagjcfZSJ18O5gSsPV7Y04yYx+OInz9JkJN5djizL0yap+Q+4QK7
8CIvj2uEkb/Gp8UIesx7Bb/6haH8vT4QpfKhUyes+foNgz3xZE5sG4BiFcAWUl5XXYySCvGJHKfk
bSmdIV24vuvPeaKHv5kdOJ1QWboo0yvvDGi62BtPg4Hm8D62uZXsCPLRThkgklVYorQZID3NsBSg
AWsGtqWlvQ+fOoyNChCRX86X9pClH7zqZQ3wtzfT/Y/YH1zugHWy1jeYEjT3vDwIiNYUNlnEcXpd
VIG0Qaqg+u/3ogHd+3uxffTrOsSW2ADxsjr8WOibhY133CNMOgd9tez4+E+530xjthL9MOUePRSx
XCzTh1TP0yLf+psVB/mCiNAe2Wf+SeI4kw4mDxplDwrc4F7+sgwiE9ZpeQSXODTk8ImjDO6JARvL
s63DlLtEVT6Uu7ab2Mhy4ETyjf+O+7ym/9HOKOJvE1RlCHCDdaf+tcBd31mASv5U+vTDWE+aaR7U
JCUuo5lMtIVRkTYuhFGr1dTlcQpkr2IpFG5V2DK/6XL4Si+UjodgMd5FWRGDiHutb30lXtT4z7BP
8s4kQS1vq+8D6xoSx3pNRZa+zg2DJXDS2KC2mhNixfG0hFYFyx1Khprn4K60gQsWcrTyV4NJYXWs
VNURHDzW1ivxbj2zGIVJ0bMByE2pfUSB+Ra5bH3FBlKmoRnRzvzekVzgOFNHk74u/SJHaAr9dihk
c4g3M09zTDjDZDvI98Fp3Zk6yoc2Ev4JXtguH3g/CO4oXnR8VxEq31rBkh2zg7w40+FGGj3OpeLQ
iiCsUoiYet9470O6cIhGRuemYsNqstEob+IYL0i8HfxFkg3ZXM8YeIuEuCkM+bWSaekTlLHCloN0
iBrUCk1/YoIjQw67rYkzQXP2bX2Ys+c9/9rax/OgQuYH9k/n+BeSTQbE1JM6S2xa7povD0h8ycI3
WwsnBAxqjcPMCcSVojqRJ2Nws+XPQ7bdYCsflXzpeH25A9TV7l6c/RnvL1VcME/YWruE54bQu6Th
WHQB/Yj5xoTTnszIvaMtu4hnpNTfVtlADjbCusf4jkXH9TJ3PnkibOJmCMBwo2MSN5hyDMlRzVrV
5gDKrn2AwssRICWrmtW+b/OOdSSRhj3mmCj/NyTNePW5bkxTzvALXu6p0TQWChyT0fPLMAqh0IX+
gPEk8n5hY3rR32QNBJXnzKGoMFmfDigBRBDsMsm80Kj4Xn4qdaNaIW5SGRPcOwU3FrY2IEdfwQUV
lsCStvedlQKL/pWRf65UNCcxXqW26IoIefM8RVKRoHitL5B22fwVHERWupdpvu4JzEPvCaggbIyY
ngDmvJolnySsqQT+96JOZ06kOTFG684r15+MNhSq4udrTCmoOu50PcJ4/I527oPXE/yaAiAhDLTu
gL3E0GJDYOo08mRj4wNY6V/Vh50zxL9+bdQlVU2j4NymF6dFfdJQDG+c2F8IWEZ/kWkhYLM0QH3j
Xr2/4L3npizrpzTxQ/cSEh3PyUbWyNgwguRJlzDewucXSiCNIybFtz6WaqrDQ8cJykDcgUgmYPnI
BPbLSYscn4edNukZ5cqQdRsIoieZpj8kEUVSc9m8OYuXwEhxY+szxsue4FdfGkBRJU0C9imbrJJP
2+eT6wJOCrNGFC8lTOHgGvfAJ1dpA+qhqCOM+uxJ077P5Gr0Pv68Sau07wCEfDzGw+pwjYzvmJrM
PU/fJrshrcGnkueLyDhojbXutRg29kd0yqGWbrdLPlVhiara2SiKSOkNLQf+oZYykNBjTpukFvni
Ni6Sr36cTjCo34aSxk2KvoivZwQAUFTpxFJLHuWEnfJMs8C7hdhR9RZdXvtQ8zcmHForNpOj2JLa
NF4VSiqvq3QiZiStIqoNHCwsD6c+Zbp/YnQNsG4kEDVT74CQZQ7NxpT6DQamQuS0vcVydq9JUT9G
tzbyBVg7VjlolSVr5aYgR/olYgRz71UCEI29xyGR91fW+4OCwOugQbPFeNXw/U5feSb4+EbuYS5f
g03Mljv+51zp6k9xIAFaImmyY1CwX8Z1Evf421efOPPMMR4SN4m42XYHTUJH/6taOYGUVTlLJOMr
zhEx+/vWzzYWc8vWS++er+7/Am7ZcWzSxgS6awQQeZMDmwibFCYsM030hmJIwaJbXnxPU0AmgmFl
lcr9QqTOsz73qf4dEQMsY1SQtnoZp36qyKZ+FqeJ+UquTl9+OlAyA5CEf8KsAYTFBS4DgT8tWuoj
dwI/rjIKSjdh7eAin30svBpXgrSH4bHAdUaApMGB0AptqgzE5LHaCFNqJ/1LfIr9wK9/hczCBJIX
F3dTATw7IUV26L4opxDueXIPD+gkeSvY0L7n3DRw63Xq5DHzdXenlS2mLY9R+2aJhHQgNtDWH42z
WoXXea6stSAMU9SenF1ZjwhTkbZwhvFDcARjUBiNtw+o2GbKKYqHJBAj7g2yN90d5Wrt/c6Oc3FU
7fiLraazg7ZpIWn/to7f7z6XBX6bQyo4lRcuEDb9cU9xAdETtPlpRcTZX5Wwpb8KvGMuTpLvHFFh
h9qVVXlPT+LZD5ADpVnXPsO1F6/7ytMZ2gfqbV0V72WxcmR4wF7tpkaim9ozVW73uIzGEwDz/at5
X+RSGG0JGQ+ao47SPIfF49ydA8ARwcfitRKKn5y0KrckO7fC2B8xl/jNojHL1kLRHI8o1VgFnt3Q
+TBpf9+oumR7v/UUshJlfXyNw/JKvZfrwrqLiF5EenbxOIUaEB3WI5Bdjvq4O5rK+VXVKSSkd4fg
Mt/HKdi8HGeL1ELgMbiufSgkTjR/onJ+rJIDB7QHajlbmPskLnlueP4Ra3OXohGFW8l28ZMDWl7R
QHgvTTt47TUZNVP4BmoGbVnM43gIlt9AGUcZcvqY5lrADxmDrhivBkxoE63zy89VGhJ91tvLocy1
WQgcH6vHXHFlT9WoE8Qu9KxDQq/fkAg2f0HJyMtXWYTtzoHJqb0a2TyI1/MJnHjSgxUCFFsQCJjR
c4swI2XO6k+oRNPr9Y7Y0Diq12XjhyQjk24cPRr9G41gplAKhiqshTiEITHSqlkRm9IV8oG3mLRm
y6zT1E4eyQiR0zqPYUsVfFYf4wYw9S8Jw1bfMHtZ8tI4a5wi059TqSwpr3ye7HsK5sNK2q9YnQuD
KJS5An65XoadVt5mmt0x6aLc3jsRiAtfpTAzwVejVTqvw5rlzc8q+2Q6IqNA7JnX2FPInxH6bjM/
4e6HlD/WBsNaj1SIhSf5Ggk2U4hT+pLNXiPuZuC3TQcYi/fIk1xjUkrsCy6Kojc7GIiPYDbA69K7
rNXbiZjdVs8eq7MSG5NjBlfEIuqJNClzS4IPJG/U1h7bB2nSLuKY6bjsjX4mtbxiIr26yMDyFgxU
Qsz3MhrAASHRFGh0uyJU89ZN1WOxt+rriMiRSNBT+E8po54b3UWxVfVJG/GlE+KH/mGq2irUyrby
94DeM/eb4fpzDVES7bXK1yUOwaLeiYzfyBeDXOy0z6IIwLewdwL/4+1g/ff/a8XKKyWoVUjQdo+O
ahaU/puoIWLcA4mNRQpJAWhUrpSb1RdQvbclwjjYnkWB2uA3ttHDBmMNqP5i1fPojjG158w1UUV4
R0pdYsHZHMvpLRRbTic4jebAM47TDYNiv3UyS6QMCR6xKjAk86iEQoybU3cEM37ZmQ6LqJL08+Jc
oL4+g32L00QI11SB9BTVLrIy4p4oGt12k4L3RSQTxtIE6igxgbscEcyoOCH7gmNtdQfk3Va/zhXY
7U1uvi6Ua/fVRbHRoLqE3rOwhBcqWnMRPYTaNDBmsJjNjvZwlY/t6wCuTejM3CW0ElhM0346WTtI
n7xsq3xbkXvVCM+KAE4HZeuLSg1ZqCTPjuYJKsz9GYrjdbuThzWl7/JpWQmUHrclmz42enjW701B
K8Fc0qWt9MkIEAVOebR6QTAW7HLl8VlFfjOWhPmVZM1NbUKvvkKgytnM194ogbXmEs/nd8rY7GiQ
zlpJEcA1Jd2GhmQuJ4QP/Tjz+cW252dFdU06kDPsiYHDbfBPKnn360ShQVKcwJghBqR29DHq4z1g
wDjeqxd7XFkBOQSc3IRDyyjiuQncNcJ6nx6nvyYuVlPREAyFNZSeN/muBm4fg+0Uqq0+KWRoVdzB
CwrwM8vYrm13YDoEWpNN80xtQjxlQ/yrqN9eVZvo18Z4M9KOtCGR0jBr8EPWeouhi47QX9gtqeOV
mf1HFxACPh9fbRc9RDsf9wR2u9CZlmcPIjfU214TDodsAvP6smyeGJVuTMZHXwoDxz61xFaIHAvH
DvkoTcSpeicz6d6PYSr7uBBqnUWq2VEOYRFT7Xj3uzeZE9GEXUFk46YQo7+QK9gSJ0x4E1YvuQgX
Sp7Ujy/6ByHbRCBG/FlBsRgxXDFjEIjW4D1MOi/9GrAvTDp8pnEnf+07sayg+SO5KrB0px22XvMD
vbRDb1fbMUi41Zm0Y0CXrDeGQswtLk+S+wurpNd91CE+GH5zi9K+QSfm/gP0E+EaPHkLNnpR9WOS
q/YzrZKcyCD7G5iGTCnFfHN4zdrlqEEj1/JCgRG4Ifpu1r1ZeyZf9Jz1b+BdPjnb0P4katph7+2G
+jE8JDZtbcVgqG+VG4HihlrvUBlOyzsOKUzAFotcd97Dzc46dPurKyBx4cTIkMR1gto8mdVjCyl2
h4XN7mYdj564dx6UApPRBexvnP5iwgF2m/CoeBLNHgvVicAcjyZUBdJJ7sFtNtQ0IHOM0CfAhdF9
C6z0rvx1JPC7UrOaU8Q4fn6l2oaGk0Y6M7nxguSJx31bX88s/s2UnT/T6jXy+TpNdkg5rZWEhtRf
q1S1WrmB+3eCQGy+jHypdGojNbvWMyjcXHPcp1K0AjvmbE+KIKKTIRubCBDe28vIdjDuuWZ0uFYg
U6gwZ5p3JnVfejlqI2nC81yt2xM4EqVFmRmemWkViB7MhQLGTTXl5+gBL3aEes9i6NXrhtpkI7XF
qabinbYsgSQktzTW1jcnIfjN9kA3suOw3dXryZHckC5r+uov6Yi8F99BnD1U0DtGPKfjXtrYKKFi
ve0iJtVRlptIGJQeGo/BFMr4ce/o5PKlwROA/eXiQDQaW1eSlMlz/wCz1meG6ZXVONWO9c3akmM9
AdGXpv8305GtXnxNppMJP/c5lxknt+UlZmkoJvLdgpoI9RS0/X4F7yv5j6DX0feoZcPfTItXLojJ
D/MPo/Yr36+R2+2JJjtZdd091deg9PQDtM0LZ9PCgcxbHZOBVnCsyCZMV+sGG52ixqcs09h6rap4
Njiei1agVxauf0AQ1iIJT4EELV4VXKt+TxZimDW0XgVuFhDrbOEU2uEU//ddUg+O6aR6VB+e0914
U0LiH/d2jxOTSwhRQOxMHnNzYd+HxSzUeJSnVJe0psBkZIhvkM2toZZh1qpjyCmHFAqhbdVqk+SZ
VQPOJM80AWiMvAE9uIlHyOTAY7GxuxFl8H6GJ7zBPqjOQ6cz0wOK4e2ODfedLZuSvrCmt90vV5cc
QAVDSZG28ae/Vcemh/u3X1gWALfK///s2/99Ps673aHF7IXqgYqCQ+anknVrxvCUb9ulnVSk6NRr
9HEkDJKyMRSSW5vxdz9PbL7K0i2dIOAIMvfd4PIkb/tLp5v0NlboHwEzFGsshxOJY7AMCaapePBo
yVaYX8DVTL/929DBDJFpb/5qDZoRZWzMgA24XPRvWW5EzPBA3jyQN2hlkQWOLTaIn8uyTIXO9UkA
brktxOTqv/QEbYXGuJtX56Kt/UxHBBu4z/JQt2DUhaaf5knuL1UlrkP6tv8DBdP59O7H+NDPmgvG
HGW+sMdqel0Od5yX3k+e6uwto6XDvYS83RLG7sk1RwLSsB7rDGv/yqhVO2JTjCsegJRXPdsfZd/S
R9fzerCUVzEkl20AelmPOAPqFoLLCyQbEiUlq6lQnymvR+lMgA0ObMNIfIqZzm0YpGP8+jRO6Uo3
zUvz2ZgAv++9jdHPyHGzeN/QGvi3pJaAl0Z+vwoPr8wneWz4acSoleqkO3zP4vNz2RLxf9AVVd/p
izER+oHcFW90UelsUsV3XPTFDAbhAf9WkNA4YJcoR9qIQJ9HuiOYgG013EciSQu4YwW1C+4PhSbc
5rxG5/65Wm5fBFAgYqNsmNX8hPhb1Z26rb5NbFETMgq5kEYQJ4qsTLdDAIHgoMvtPnxzA+IWtf9D
PDHj9rjelRu0fytr9Rby9u41Iq8FQGBOyJq+5npaAW0zk6V1hNXabYPS9VLWWWvsS0v7PpNnR4qI
ax7ZniccmGeaGqlF1F50kYCn+rVLuSKsmuorqhg8uzxzKsnLj2NcKsxH2MH2VLVX8t/ElaGGoAny
WhUhkD77RFcNL1x6v56aGH09AfDHs5p94MOY5gjoHVh9k5+U08r6hPEyzmyvtjfCwKrIBQwfePNE
IHq6h5A+BUoZiTvzqSSUQwekEI4DprZvwiC5z0N3YVdjcSyXRXQ+JJqJsqRZdKVBC4coZkg899tI
5pvZv+IZxtoj2KcSopUCnMAOehMYNnGflRas04JQX1nxdFDmZCwQhA2Ea36wJfeXV0Yo/Y0nrjQO
DXGArmOJHXpv0IMgQ0gXV2KHZIUtDOxHCC6GtdvUXTTejd/v5PenuQTIK80iJKIUiA/6fBlciYkh
iNoz4/ZboFPyCA2hZjm+r5BLEv5UwKJs1jDNPnzBZP/Af0UfjBN8JHCm6rRe+vr2PiRlpnBkg2ZT
XcDrPD2WJXeNfXFxXf8IdKX/3xT12+dMy3EYah5NUmUHxPtQANGBToHgXKGMoq+7iDWTFLxwOwD9
AP+/zKeE4jd4UM8JPcfKn13gPU+Lt8N+SNtoVq+YUKWY/IYTi/7p+mE0mmExxYGZjPjByiEWMiAe
GFWVzuUAqVRuoam4Sz46IKe3I1ygW8eDKVhlvsXoCOhvOJBJ8V28AqB2xkPdkllk5wr8dTtxnaaW
kb5kJE7jBDYlcr5/Jys3j0ysj6DP83WsirMtenj1DUqb8W9pJAQX8KxU8I6uc4n/rGef+qGLl0Ry
h+hqyP5sQKyvM1hMIrxlJGX5RbPnlahE6nSs82E/RSgueVdUICl9uOMAwGBC1a2vwRtRbU1Kx2dq
x5NeZDnSMxMVKbohpnN4F4uz28eyHYuWRuZE/f77kaNhUSJtkNzdrWk7jcettAXMlBwYxOJQCmqS
QMTokPtdFa1opWlc/sxLkTd/uePDgIEALcG586PaDFv6FzSkrL4L0R7H9HkXm0wSXINUS8OVqvCs
cbsuGgJwhtnJquPRiZ6Bk9j/TSc2yccUvFxS4icWon0A+6N92oY+JkJSUJBqCKJWLf45CeJRh9/I
jWQSxMxKI3EeXaAp7HtxpictwbvmZ4Haee1c1eFOTbgogE3vs7650ly5B7eLekKcp3TiDm+Nc4HV
tCY72WRVGA/qdAiOLjVJul6/TWwIpTqszKOm5Z4HRaL+Jx5Jks7oW+6PiYfLL+Mpn2H6+EfYJfRZ
BxgO5pFQasRJIhWzrjgC37W1WQE/IlW099gsGyMbtqb7F0SnqbjGxKLzuK2ua8zm/hCWamxh1fdL
okwqugERFPXDCtJcGNqZDzoRxpIwomtdpomT8GSoK25EmZip8ruU9IQ2L24SZeV6CnEid10qdlOs
MsoNUhFqUr+6LebXoNcsC4slX4klUU73u/GwCKjXQv872elJsueTCHhpMM3xTHmkUx56VCc7r5Av
ZSMMCrfEIg4PA8lre8wT626S2ILJ6nZ4j4IV9tcH0SDbn9LcfZy7EOdSN9FX7P8rNpO/HNsZNKY9
DRaSn5kHImU3AsaadsxGvcfU/vwYJ0+UIi3wdumgBYZfAE/7XdRxumg/VFuNwF8N7Mh3j8usWG+8
F7DJENshX8+asQjbVeVyjP7IvAPushkGzkBvoM7iks88hJon55bhQopaHudsTm0P55+tInz8bViN
xTBcF6AnjrC5q4Y13AxiozfCX6LcYRcwJE9EPxPrpQ2T2Jri2MCoLA+KVL/MO6nJRiapiZd/bSqq
XoALYqpxm8W7L60X9fp+f+mO/C17bcLvTd4fN1DeFXnNgQDzllgP2QdIGxlKxE7x5GlL8bgIHNC3
lLqMpxn4lW9OFQtP+OFbBsZGK0zjPfBQO28tQmi6RBsqT8n823sHoIyaBIMcIOX1T30/yd+4/n6Y
assZr0/yAh+NkVjGoS6ZGPkrTg34Lbn0zZ9IE+uoyWhsmnvsLv/n2aUT8nNXLwUEMBBhJSadeKzV
UqsDEdGDVA+5M626wBjFp5cBAzCPZWQgAoDGtpJAWXDpAnDi2AJmn7ExEtLK7/0+OU6dUGgWwWlR
TkxQ9jXPS2D3uTE5g0Ex/2AlHtKnLYyCoSxud5d7OK1p7Z6ydnmDW1Wp0Yd8P3OUjSod+0JfdCzj
MYipFEjR9s7+ryKyffvhPtDEAdDIxBcy+AQ7mrL5o90k0xXIqwd5rCng7m4bj2oyna3jbdrAYwsq
H6EUus5zjoxC3k/v+5WW1AqwDqmQpoQgvjkRxFP0nli7QEtKpi7VwnIDsG4McyLyRYUfRHkEM8Ju
MmFvCgabmEmuRtiK7FTKO9WwT1236PqzZabzshHSfw9roExc9R5/SaVpX0dOXB9hGdirddON782/
G6CLFkItIvENV0C25khEwpr4/F1D+9xULX06dzfjUrvbdkXSpzVFkkwZiykxz10gk5cFN3TZ8NYv
Axk1Ycs/57YI07fK096T6qNjYjy3V+HbqNih8rQx2rlzY7OsY6uIjTxQeXXB/UzVDh9UTGeQfVeE
2x17W9J6hHjKOLuJmGaNuDg8HR4vzt8VuQH/etoybgM/+F0XEPBzDWfSzZCzZxATWo03mjBN3f8Y
ANSC7MprNlhTWKVkWLe3bDJirdWirdKdBLsNkp2a8TYpA+bBbU+Y/OcSPBhkIiOmJ8y3Q0QnoYQv
dVsiQRK4JM2LN0hxlTOUfdxIXds9z5yRtVpxxAZr6DkxDzVmw+Ol9yKe3x2BTGV43qV+gpUgMqcs
LcFN2iQNiT5csvgApQq9WTHx1bNE+cnQNXT6PxucFKTT4C+kDyjDQlofdfWZG2uaIixPZgzW5rN3
liq+nC9QgVIL/AdVYCSfAhv/2pEtLOCYq6hHZGxZTleG1OK7um3+LQwyhG82Z69e/tZAUiL75fih
jIvKl5cA74hPvZnX3SBCJUIFaPXObsjE+XexCWmTk7DGvQP08qoy9/rV8H+Fvdrsj/4EX02noqsd
k/wcGJ5m3A5Kal/w/AzdRIG3g0dfh5EtTr8ku0qd1tmVG90ztpughfbwyiadIxra4G1dDiUp42RQ
MFixjjypIJJBYbkYwQbhCKgqFJeHwo5xEZ76tdCaaM2+qWJ8jK4FBzka46lf+u71nMHEpfmdr10f
iRH806ebAKoKRgPkhTtivrbkL0AArUoK6frvUe4tQMLwLL3QTlB2tbkvX/rIHKLwjCuZOkoMdPtT
Px5N8vCBxj2rWoWfLIwAwlRP3v9u+HU92z6RlFne6om2K+oSWHqx4wmqsInMb/RjmIw6Idop3Yas
AM6MeVw6nBopYEZVBuVknCaHfeFloetJYAwcGsU7rpc/JqLPcRQhaHX+YQd1KcMpDLZLybFBdVRM
1bQWa+ESKvYYCy1rwFaX0eFWwKUeL/c79r1nrMdswHAbEVmB4zXVS4HJO4GamuORgW2F4rfmSiiA
12WBTQWLNkYrWD6GLF+U94dXwkgT3rJflkLBaKPGLbfC2xyLv/swsJ8ehvOEWArfUPXmdNMj4y03
uY+Ds/GpGCg6Db0JZhWIKz+lQ8YxtU/wIr8NPymNe8IDLwqx7YgzpuMISRz4+ImsW8Nyj4398dXV
mIR+SxmJ7RjcCLf8rCIiRBUeTngpcw7T+GKv4Pf399WSoGs54dhgvzEaydCNxYjPdqoPKs7O5anq
8eC3qqWKevZrF7a0upkjPv1Vr4ANPvlQgNP0kAo0QwfLeN/OmyHFpJzVmrLYC9nB+VomlGiHmQF/
352Z+rQxDgZkRdWEOE68bUmTGdScNPmxcJXTpqPTXUMcSM3c/b7Qj8n48w4Y/baWoD/hzFdlOoh3
jkH0SvDh9VabHNS3c3UbUZCU8U9foLlM8GUr8SLo02sRmCA08JmYkd8yhB6qKH/uWvzXttftURaY
Tiedwp2JCSDtRnfRfjfQs7ejpmjBZfBw1hcbSN/ciphqFkjUFOy3drdkpMuk1XcqDrhA8ym4u+bo
OLQQ+8jNndVU3/ZhbMwTRZmJ6Oxxa2IHA0zTKO2r8caYrDOi304wGlrK7iCloCyRn7bmPdaA9Puz
wvTJNajjeSzacnsuChpHDLi6iBXGiNEvpJcVwgdPI9e5yFxuAyPgOHg7VKy2popegqGcgYIPfqpX
lsilUouK0mmNlyu67Axy0TctxtcbpobCMFU5sZLPAqudrAGxBr5NqjDWexjcG7KjBouC9VtBBTmx
WkGDTPbaKTUn5hfVigscBsHeJqkfgShtr6QQB1nQUcPdbndg1LneXvg1q1KomWmTMBkmBHzelG8/
Cumm77rRu6zcAfWXwiKu7PwIf0nR/pRQRT97e4O1fg49TMF4Ip/0sL54UG+MPGyH9kY9Lz8gmqfZ
XrZwRvnWxlQ4op7zQPjDpZe5fTccVMqI2zHFhJJxTwVBy55T4PGlbsw/NKA/UfO8dUb2Fjj+lVyT
ds5c0BZnXgF5sSTF0CtsCZXNYHT8F1CdYPH2+JRsGAlYgsusOos++xr35Ig6ixUHi34g/NbQnqLT
0O1nJDK3giz/zavV55qRKC8MsCoBr+hdvPfwgXFQUKlq2k6gIn5LQQBhL6yk3CKznGeF+om1Ustc
tLyyXs0jBKEuiHuF9Yjo+n/zTLW9DuIic2IO5Rj0w7mBjFteDtPiVT3kNnBLssgWkzbKKsqfkHeB
3TfKTPlrU2l0yX4U8CmMMW1mWnF+XF2BsRfJ2sIPSgEhq8AvWth7yLAuvaP2I5Bdu8aHMvWzPO+Z
h5WrMwV1eiuoq5gsvsGAIORVya3T6qneL1kwovFgl2iahhL7NoK8sMOP65Zah0jflIKpcqz9VucZ
S24jxsysvXckcWogZ8g1tmWQjCym+2KDegUa06ERQJV+QsGpFHOjA4+taMkfi4POHn8+82J7rr7L
FxVD9I2I6mju5Yxr9NZWY9O1hfOB8oPkCZjHr7AOmL+a3I06meC5pyrmS6iv5jbfyAIvLvdU9Voo
QzH+1pJSeSAvFxpjOuxqUuQbUzt3MgyJyTiTi++4iSHgPRYsNaJKZO9YmA8VmLd0n8pDzt2MZFv6
ed7NxQA3EF8mFbKrauv2OD/Wh64nr0fypd7a3HjTW40fdZWQiDSq3EhoxnDkUoZE3tKcJZA9mQ6T
AbIDVXXd69pyMQI9O1gWrGbUY8kD4MhwsdQEVg8Ge9xt8NqvlfAkoHlSSOlIsU0fDTaDeChZTfaw
v8eKT4Y78pKqSEEKg4M68nMOC4NT4ogC20GPryLeCfmj2fGtZff48lBdnLHjfQj1LhQMfCl8qk0s
03205Pk2jCnvc7UueWb/DnVWp/aAkgk26Ywi7itNfNuzuepVox0kbPvlDGrrbXpjZnPRVnTZpGGy
W9actC3IZibJoax+X5I4A51nvuW+NOlM+xBWt8pHNr5+hWIB0KdhnNnayxrukezkZju4RaJQQTAp
qFuccdJHp+fK3MlVB2Bbb9lrrDqNjNwiA2Ywonk83PMD1nIQcdgzLwVvLzuv3H6rJtvYPng8bKsi
ADbWiOFEx1L39HYWY8VkKBZib51DcSumX/KYi6rlkw2o9hAEpyZqqpGy+vONAVDklrcjDjfdLOUX
ebAjzNrVLA2h0oH0v3SvvMnwmHg4VQIHdsyRuCeNJZvWX0QwB+3xjYsWFQsANzFLkp+ww7t10TTE
UTvRE+nDLrZaJjHtj23Q0HKtnn4egIPp4GzaDA0LfsSKSjA+D5KJeOlMmblRf6SAIhNUjWzggmHs
hpqOcgT60LpZUfd2BoZDvKSBxQg9Lor7ffzMHTcAq0K85Dq6ysBDOibujGeRpmAvWECvZmdfFbIW
TqSb7x7l30Sd7ZaYV2a6HT826fagIpQwYLwdJcIIVX/GBI+vUZUle54wAgzMP6YeIKTTLo7xuq6E
yKrto51raR81xAtVKtGZ9iXhx/n8QrJJg0hWNBi8/SPE8SsJFfVrnLv5azPiZPubSwk73E8AFn7w
UH+W5J8ryvtAMfwmGp8Ydmg3yn7jbtW5eyXUS7y9IS/ORnxNzIWphy7FicROiJylw7iEpP6inHuj
RksJqasg5PUQ58C0OFNFWfG6UBoVIEPXjxjrKWe/KwzgQUDe50sb9++QxMN8yl7ByvwGwn7Zqfw4
4QX5GbAieUXD9zrRZNBTRQLHv/uYcfPZNOmzNNIJSerwKH9aRVTbGnhvKWHzQO0CwavpS2rAIr7g
XwlRAhNaNdzj/U2LU7S7d0L5BBb50tLFIs0a/d5W3IcWdVagWeFxTaSY7QTpKV/NMAH+vGt5kSaT
un43q/Tyq/JDRZwaHYBxxyqegMhMnMNwUrIu0zNlDOFnnnwbpxTohFAsg+6AzGALZXDVEufDVSvc
wi/xjKnfMcsWOd4Ehtt9dtbxIwMsULLav9fsibzalaVopoFNdP8ddjJR6LkPtbYBZk02qbHjUhiq
vXdj0DCPoT2DtPazGsaIkltEh3qLZDHbiGSHugrX9pxFrkEAHJ8FiyZx3VdXJv528Fo3Z2HxLEMS
ou5MU6OmwmDLlvckp0z8v2fVyOItB/suful6adeeObKTV6CxvKEOxfobd3VUANGf1MD/iPdDHCeP
epRLP26aaZSSkO3Zg9IOAAfARIwI532SFkcZDfqhV0+jaUId8pKEtWTql8LJWuxLC3BDA6XlZTNp
ndHUJvmmj3ZaVdkZlq/PeBVM+Dpa1+sVzOyqf+oFZLi62aA5culMPkHQuxW9PCH6a9GnAR1X9j/I
BpsnRUQGBsdqi63ZquEJwjnzSincrjEk1ikxv/PjE7OG1447u3sMDlsA1VsvlQP+ffmzqpgqwfYX
aLx/PKLnwdpwQYRyhDfBb5eZ6fpKxLSWlVZ6QdofPDTWGWLiWv1vn+Z/JPG8oKr13dhQoMuFMtAt
bczOT9YUIVcahD8M9NBsqqDTe5ChpzPglppP5DS8X9g/s0+FWSJO7j2f/Fn1PcCd05V9g241brii
OSkzlv1nKqtfwxUMnAeSPb0i4MSXB4AD4mxrthUo4NXUb9CiZdAQLD6V/zS8c5Pvj5W1pJ51rz+e
K6yoEforS35+XollBEK3S7AY3HccbBmy3bGJ4U4cVN+l35ip5Ctq5dmLaLKFUPxCRgBLWLZGCJ4M
hF+IKO6RO6rgNZkt/m26Gci7jXrLLaK4w4rkMxLNQWs0y9vhAMWDckFraB+3b8nvGX4H8jDQFWt+
tufaHKv22n8aV82W+W0+k1MvsOaBI+8dsOfMDaG/qMBKCyXa4w4B6cyBv8YZRU0u/BEqpQCGCYTu
XvLHykYoAuLv8m0ponlPimSU7ESyCY3Ykpmy6UUQgaFR+2RsK3KR2/WtbTbB3B9vyAfxSdxxMH+u
9+1IXpw5ClcGHVc/Uf3rFqRzfuXdkS6EokL/HwKKTbf+R2QJg6suzMck3C2pUnYU4bKnNECtllsh
xvy9mkP83y7RO0TNtdc5pZ0sbsuiX7w87zQ80e383lVcbqBhtXpcTBlfKXZjvXnX50So+WmJQW1P
9T2lItuTr1jjAByi605mcZgmx8LshOOhAP0pv3zx+bjaWRd4uKaKfzLfaGNhg+mu97Ap4Keoyy5x
HU9wqSwRPAVE06kKpSU/s74KgxpwZdTS4JpHUXtlKwY9r3IQwvu91/L1llAM9DDEf7epjLM80sRO
cq+vVrC8c5LYc0TBbRzqmWS51fJZ6LobNlu9cN7XqL41gm/ThLtOfHwftlaU2UJifpr8XlVUXCZ7
x9odhjzmch6mzMe/u/rYTLDdUNvgEPdQumBdfXr8RrySbf1tcBjxcqCnojdcNE+vuRi+DqekeEDB
vvCZQpcTrd8Xi4zjOc0eH6iuVfg63GPOOn93EviYjRAPGyxV7cXeuHjwunaJig8x4kF9lXP56cwo
OJW9fstVSPAm7MwVQSfdVKLK8qICcR7NH9B9wVl1B6U4IH1hPJZo1Q+i4/YgZ5n71zMTmOZCZIMd
YjIW80vR9x1pS5p2IAIik8trPSux4wRnCxDcOFS60Xc3rdkBJVojNPhqqCFhY2mHUrAKk81O69pt
qSMoQhxEmU59J+5mdxyj1L3bABnhNUplMP4GKZ6oAFLB5Y0U9IU0dV73VDeHi6gEmXDfPU8BLyPG
+NyBMeCA+H1FwBlPyiT5dDMHFqJV0oizTxdXUUa7l/DBQgeLmA2NdAvCRC0WUTl0JC4ynxTdSqiW
ewayB2llnU4L1+JSAF/gTb6eYf7uzbQzu/OgjAfTsefU+rf4HRP0bdBczWmDIMxjRw9Zne94GxDo
yfcnL6ycwFf5s+lZOc315oOjcW42F5K52j5/7ALohqZAOMjRjT+/h+8Gz56LnBcahezRmwUsat3j
tw2g3E7w3dS7ObUjPdKJE5FZAy/sYcvsLu1X42YFh8A0IOKegUBTabAINEm9qGWsnZ9aoi+RWFu0
h1upLmNcck72gnsrJq/Ve4+M7WUujzRLdZKjwUxJS8jXo9dh2MsRdji4Q2wAA7R35xl3Poc3PeuQ
jOVgL0aTzjAyEkGdFHdr+3OaIH+rXhzNAfl7Sof4aRoKIKd/m7T3e4koR9McOisMLV14Fvmehyve
U48QNL5obtSfLbneCS2v0CINIH4nE85bUT/2QkV5Ea5gn25srQd14Pl9CpAO2uYdCoWWgEm0APtM
/d4R2jJAmSE3ZrEIZKDY1ep4uq2+0GzOJbX1uaXUT3tdrhWT//521kQOkDszr6jo27feOqwogMXm
lx17EDNFT2E1stuxWdOjder+xrr56e5GU07h1DJ1PWKIB+90V2MsqWcVN6UJ/4ii6G4BrHnilQtw
lkj46paBG8KyEiOnp8SGl6IcORUN78AA1brWL1CT3mBkAWTiFYTvt3I/EO1ddX4u8BMlNAD+Tn5u
X0HG+3AUszaOGsW12vTk2giyYQrDEiWYd9cJEscq2qGMQTf8xtA6MBd/th4XUoTgKxnoYR7WS+Wi
XY3MTMaiURCQCRmDUiQK2wvoPVxcNW+qn/gtb/sAEx25jKQ5OP4rkUHa18oTJyUDHmEKiih4jE06
bQPDaeWTPI9u7D4IHvkAFmLC/NNEtmIr5dCy2mYxn0DrtncvL/1+VZBsWzRaGE7HE6Ga0c8uXGmP
C2fWbViclS8hFqvKR55ThCReko0rL68slMFKP7XdWw/yLXH8SdhvmKmZgV6aRyxmFEUpd8+L2I8o
E5Fk7HgMHU/Mi+u0ivGSOXM04u31J9F1eRY8k8oEwYklsacpjr3QmbRMWvLWcR7Rvrcj5T5W17MZ
vL3W5cTCyl0+rW1LjRPH2dkcWH7bKg+sfHaQ7ZVoViKZ5ncogyzbwLeT3Ei4tg6/cJRMA2+cWLUa
XFpaja9EgKTX39qEOiy/8oSdVpNmu6pgFR0JL9RqYOlsh3htMVvq6wxccMzrn+tPpAWlULRBZpir
rxwXbEEsfT1mhh17bAuucFGk7awtoKRlP/2I2xi3+sg4Be70qXAmdXJO0pGL3qW4hVSIPRQb++y5
CD2rCIh9QxM6za10QG4WIgnmTLMC9fJBDCTvIXCAGAFRT/+v46iXjcx7nODQidvrXvmPWHLpmGOi
670WWm45y1we4jSDUjdJVau59iHhExVkAGOVlbVRqSWLj7+WFlZHZ9Zr/IeKmgum18zOYs8bF1JZ
Xpyi8OFg8KGFNpin8gaq1sewF29cQRB4vhHS+DJjFJE5FU0JVXyZSGVgcmAYLUuNDyhhGgN55vXL
Ew92hABPxNViPhK0bqKv683F9gHdKkqT5SS6XT6gkvm7j6thVA4Dvle2NXgbW/bKy72kLfcRsZo3
IXwD4IQkzLic289gQ9z11A2HxEuNkZnFuz4Csz+oIY4AucK+g0olKDO5aFHIDNe+/boulIfxVTZK
RHfkpStaA/UtZkHw2WcJH1tOIyuaBSEZcsAYQ4gavyFnOLss/jCWmPfsgbYdVJueEhU39j5SEWCq
941tWx1+vusttbhlDkO92R8R5QvoVmsDIcTkwDKkSMBOq2M1OPz8edJW98/gFA6D/Anw2nMScwma
j0HfbRQD3IJkF3EG/b7LHLyqbwKfjDSUpfVfXTUnHOjrboA0Kl6DIj7SFRIJhgO1+rLGBvchPj0x
0f/02NQHM5125/Lv8bzM3opzKvpP06/M1qOmr2lXXNGV7TGJGJtSkkSIgBNHguEJi+R5xEIEdTPA
9zG6rn/HElYVWldfiCIKhizdk6H6nvwilTNvMZh3Y/lBE4ZUZUZL75rvS9JZWkfJFZePlo4JBXe+
12FJyO1CJ13/+nslLTRK8Bg0I9DcTq2I7cxCLqgpE+N4XpJ9ZIlK/Zewhy37txW6RrnWisgt7Qq1
turgAAq56ABowR26J3TfWby1LjaAxFEM+yaf3ByFpoHFcSWtZEss+1pFS3WMPS+BiNSvFWD+v9xw
TdKvix7fAH1kPMydCafp6EYCZulvzri4tvejyCiKmVUlv53nKd6QLgLCH/U5JniOQa5FGzlVsv6t
iUSfNG7mBMODRE4lRhulCUopjK+jihEMPaa58Ag9MWbMP3rp7qc1cAILf0ujHDHhzaYUn90bGeCE
+2NkR5ST/9H0PRM/2B/Jlu9UY24ZWQELXs3w7IQj5sLv1u6t14hq6uCKtjAfWC9rfw6Xf2CeCbyK
MjabOUtOwZCWju4dsvDZDF3waGQUL6xSLIJ8ofhiILleJ5f1Bdk5R/+hJQHu0SlGzuKv8KCj7dNZ
EIdP6foXTH7fYLfna5fRSYBQoCvYFSAJflBXZkTJk3LAj3NKDPRSmlZV/3U1R8eq3l5jGToenD/Y
1VbMSASKYO6pE7SxU4FGpl0OQj2Y5tLrRzEamxHDMNil6ul+T6ogpi1gGmcjiG/5mEgsAZnDVC/D
2goDGO9lTffCUlP2fCQaSXmZ0GdJNIiI4fAmxL9YXaLu298vOPuxW7GgzdvfliUWfe+OnsZzToxC
sCe5qDsH/V8kms58G5QOm0vH9Kdszb8v38vLwcsP4Yt7VNI1/qzTVR0PRTxnwhPR75kk2ec6SvWm
9GPgQ2Hyr22LVxjj5nukUAoxCFhEI0uyDUnwNrCl4Rpw6sD99PWV095MIpQ+LSC7uoV14m7dtveA
CBKI6uT54V3Ofc/4oPF6keYe4hUMIg37scODCFOTYIX6kuvfvWsNuH783NLyBeA0EP9bmA8Agx9b
PLQZRvtxjz4z+4KANRD+2bwSEwhGaAsD/h6AmL75HMNgSVYr4dbWjcOzG+ZyFkkbEle/yrqB+/bI
7zPGE5YxQtdkqFHDURTDnvXV/sOGXmVujAdNhvinMEyoMIYcNdt4Hg8j7JC/ys7K8mqPZcQi2VyE
Sl/aKnP0fq+x1g0eETKgQfFlEyi4kJ7j21p3Jhc9IHPSERFPJ4ehWkKyuJHCK5pVR7j0PT3trdsd
jsE5G75hJPAN/c5zARvwlyegwiHSBU2kM4xJe0TrAn53z+RMjVNv8tJQ8e6fAWgzw/oK4J9VqSQ1
GPkDKzU8aEY6/Bd6sD2WuN4W8ofWrHV0UFwl2ZBnDtUFLLmO/HypFqfsKlI1rPYJKknamhBKkUA4
QHx79cFEhhzUc5lbRUJHTDjUtcIGzPerknBePrVBWONY8AuCi1ioNhm37Lvp1BMzgxbQm1OZIttv
xNdXbZ29+g/vJ18P0FiXpK/Gt7PhX63hbAwbvJ7GVT9v4pyVSWs/w8QaTN1Hb7ihPe6lielhU2jw
gs9zPMPKL10OCAyFhLOflrIIQFL7VJqyy+6Fr3sd42I5zioGiiBiWCB2zE4y2sWGynUJt9MnYUC5
TSblWqGjHyF4XXbdAAdzIivF4q8l6mDxNWKW5Mn4Sq2DyecNCK/O6DBOSKykLmQ0E9Oh4QzMj2G7
vfcbAoTuHTlhrLei+ShF+4vBaDigBgSpp79J4hPksEpfALeQmK2dlu/LBTi/FctEavk5gKmiNHgx
0x5klZCA17WrbIaCOha3waTztUKPwYZQdU8wulrUzLLpnv9gq9wWyWufLCG7fE6dIBgwbP7x/P++
aQMEqDtOfP9BhwLKAu2wBnH8iejcm2VTQzLSQKt+2jjzu5nP0O2Y9r3pDQ0iGx6zNe9BWinpudhB
woiunLgVoLY5r5feV1zITObw4Llf42ocMbHtiKLkdYNCqpwxXjlFa0Ise6xThYdp8zgFKeaCfNTK
fu9gsPvMXqASRBeJY0OuDp53mxK6Fmy3kKcgpJBgVivdfbq+Oi0ew3oPNshyZKFBgbq3uBqbzQE6
Q5DaLH5wDgiThpe2KEEqBVWP61Wwih1dV+0HiKF/6afa1wYz8Ua5XDL5UAyDKj63Duzv1S6c68k1
bFt19PzzxzcNj8LteVD0zweZ2vSJIgnFBrQZrk8o5CcjAttwnlwpoTwBkHyaJXBp7tX8aD4fvPXI
vQsnCEte42kSNf8vwe2mwmqLoGv2nH+d8pSil1WpbO0NJNo6eFbmMW/tIz31SiigLADlCROfiqbB
s/NZtNY5JY1oOrPggSO0Ag+T6OYXrKKhHjNfrHfLeRBMW3Yht0rGiGDSfRbEMxEvljdzbPwyI1ST
u3w4xMoIR2TMllrXAg1ZoV5C3cGiNsB041p4abRpvz+0/CrGiVY0iUlrYTErFndeFwS9RsNFQkeY
6gelzp+m19yh/8S5wP4rKGS46Zbu1WVuPeOsxREcLBlIutnrFUyQhU7QJOXH1CJRxppLLAOz2ZRB
w+S3NPwdGx+rN8lt1mBHOEAPx7wYt6VjprkqcXvwjiwiJq9BokQG6sA2uVLjXt0WO+KIEsj8/JoY
ng5dshvmyZNfce7YHwIn9T8O155r8PsnpHFh+J9Ps8B1sRwdV1SvULel6LWdyQivSEkI+XY2zLuh
s3PUlyxRFL4tn6AP8NslPUM8iTZfEwDkXlxkOpVYV7FlSolmQbp7emCg+rn7Bo1y72LoVmd9WPlT
vBX/44jKeuWcGTC46sIGvtOtM2N7G3tI8LJJv1ifFgqd75/4sZRJ4NcaZrX4DD1hjUU7PK8/rugY
HFYVAuV5Wa9oS73vHd+l9HEfPgv9+A9F8eAXTrymi4pEEZLh7wkTWH7ruqEu0pdxcqA7GKlUf3sI
ncslFPAzYrSApzBW55YQt8uzHspEcPyJ1wKld50VAjc9xco6Wc7TNKmdn3JMPRxjbCjnvroRpJuY
vhTw2Nr1JVFO4zY9ylIu3BegAADsHj2U25yhy1KGfW3a0M33+xxb4RcTgGEJTpIl0P/g5Lacs+qb
QftwqiniIXHSu+/avYdjanm84pf9/Oyky/dCTr9WpJrpTom83vpca2mIav3EXhS/9wKj3HFJWmEx
WIrVktyXAuRGlU156wEdILmvh2BMFQDlCZWyBmyiTdZbCSbExCm1kQHnHw6Ko8813HHJy4CEIydg
VfHhCwzx2B79mewTSpHzEamLqVp2TzB6D3NBsGChFTkmWWEKpAyvL0UXERcRQIQHkga26J0pPZfM
WlWQApddD/18sKuRZF5EOY7dqBMTBEkKadOY29hDdjZbvkxY86HCzFwRdLF7TSN+zSgt7x7OCJUl
h1ZHFmQBmrj2WSunLmIRj7ZlqoyM+eLbR4htBpvncCuq0zH1f4Vd4WQq1X4/DFZ3OHbaWXX51tLF
pzPUmuUyoq5eGNmXve3xgbcI+vZccK6xnTXlHQT8qCAxWfig6nKElJCmLkiqXrpKIOHprpF9iSrU
hdVz7qNnLaJRllBH5LOyfBWTVRyVUwJUR4X2BfCy5m/9xZY9rXFQr5YSFgX5eVfdNQKchlfZyYOU
CNzydVVWCZbmUbMnI6TVEyOoIqHDiOn+8DHQuWbR+Qz7t3FpujZqxu71IQYsUO2dFcfeIj8xX9UN
vY3dTRscVaNbJABrcqPOWqGLfz0zxf9JPrE421zsTeENEXhQWfyJ0KvC4iYH1C52Uk4/N8UTzlxt
tEj/JhH4xvYe+lCpMiaJD3c+59sqic07w7j5EtwqujaMz4vWR8qc42DEkOS0pFwLqjDVSLHzTOPy
pWzWbA3FYtWuC00hCx3GUBH90qFD3i4BqnbjsD4hybJZhtFEkcTohrmnpR+pxboJoe/Xn/yneqXF
CImK3XOM3wmdYFU+zZ68t7qJsQtZGb3ZPXlaxjNG2bBNdp2uwh7AJw9fK5cYAtJPIZgrgCPgkAHB
78lguOknCRqaIzJkInSEL01Bb3RqeisjrVJZN49m4uY65JLQBORnA9jWhpbTjoiiPCDTwq/xfVfw
GTr86MyurSRq2CVshsUlhTHFO4zmK5nzCbFDp2Fk0Lo2iuODVG0Hru5E9X633GxRgogjUIDJjnGJ
GwH9ktLxBLDFhyAjFMGzs75vb177kZb1zfi8z8QUe3q06uQ05/Xsrz+pi6UO7bBOHyH03QN8M8M6
kHCJjiV18Dt0EyMtG/NYpKSyGSkkVy1wgL5WMrnw5tvcfrXkVY5h0cvcxOcLt4/2cSr8SrOuKCyt
eGBJc43+S+vXMCOW/Gjibk4E5k2ZGwB35VzapeJOmlzBUnnGKFHvQ3K4wiVie51SvLqEx4zAYnbS
WOXPfEoNi15xlwV223twnNleXDkdZ8IaOy+gr00S8HZYEweGy9toFApoo/++yxWRgrFBzvOOsyjD
orRHlPry/lyzZWJ2C4gQF5ToSO65zCPctm+9ORn7iBBEaevQZIgiczAKgs6br1P6++NiKyErpx0g
6zTHfoK6u5sApp+aIvMqAet7oeBX9GMdXnChx3lg8jLZkI0HAOLflgqWmhPlVfA+AYAtLQKoPg0s
LR0ZPd8EiIOd2fNvGCks/qHqnwFJVLPoVln8WK7I9XEnjrVf1F5PBUtCzlUVJo8HSo6TcBT6auyD
ySABbrimluKTu4Wts6Ei2gtTBLqpw9+NRG9h50lIbAL5O9zIA9r1N/PTy8iM9zpLA5JQlbhfRtcP
nu5aauO9KHMJLlLS2ZpPAJVE3Z8ky0KSPvlEnaLXBmZtNkD10hz5Gr722YtJNsb/5xHFDRzsDDYi
U0xRBIWs7P05zYg1kYU4rTKCmNorKtdLC9p86USpu35Y+iiPor7ij1Ff6Mk/OiNFrk2wIVLk/e5n
T/9PxdkVj6Qjd3W8sa7qq9FMcTRVDn32hy3wHEtX1FIMwSxXhqFV38Yq0bZzURHAydiLn11HjGwL
cbqVTEYeljiDQ5Vzyte58FK286ohPNs0V3L1+X+In7PI0foXr2xjNzbyO/8Wa6xvl4a/XHXTr6wz
jo5OZ2pHX4t+PFFUoArp3kpR37KAKTXBVNRd7z4thdy+J7YVr8UbHy9Fk/HBKJJZ05ct8D844A2F
A/ytp/+U2/dmMuSly9Odeg/Xy8rE1gLqKB7mDjhmSXonhXE8SXFVTlAexrmUIda0J7TJ50nyj2le
89jZNfGEwfP4x5GJpRcbMGBDHnprZ+8b5Epw9+On17UZsRZy+qxu4/qxbDDRKqu87KApQ2jLfZ/n
6H9adQJHgWNbjQudX8izUbJVmKdlkvgRhP5rqPmB4MAb0+zapcXvllSqV1ix7oIXdMoklvsYWnej
pR/JK0ce7C4FBoqGnrCVLaEKimRudWM7DTEOit66dpTf/SfpIXg3jI0KDhxlrCM0WQwpZzNs/YCT
o85AOFQK1/3x7mrVmONAxyvlYYr87KTg4ygsXtifQzPm9Z0uz5vrU0FOh9UfWwJe/omYiFjJ47+4
w4NlL+1S0bwDYLU/id4Mrx6rnmiounx+JBdwR4Y3yAeAJN8yo5BdZ8RDE4s54tM3wxObiZNWdL4y
LPW1ZAJDLcpul9pj66c425vrI2MbYQtU+XOXfNmW7TstNjDME87F8q1OwF+X3pJuS4qDlaJnPdmy
16Hflyr2DSzvwF/v2rfomHFRfr1W6VNoENTzw89QDJRwgJeYKG5YRdfUNvOEZZP5GWfWDg9ZGYXT
worcopY2MsKtrbN9wk7Xs9LUhkS6OdVMXELcnmYi5d5XfAkf4SAzP1IgwPBQ6XO+uIsp9YRUtKw5
uA4/e98kRNr0pf5Ud0zjzeAKuA6Jm38ivoViWl8prxL/Z4drl7Rh92QU7SXChbtsuKHLgAW8dBB6
HlBt2WX5YDMf4a5sud8xEfigoY7peT88Y5SfIjccYX3SDn24p/tHmv6e0wf3gjjHQw3Drf6LgwMw
ttKTbI+uxwNwMFplu0zKHus7gN1e5hqahjhEJ2qj1239bLWNL2znA2UE1aipkP4Mr27rRnrbL9rV
zgIye85HFQmIlCCwA+vpi+WcLd0gY4/oKGAn2ICDkya8Jp70LpC/UpbSQOdWstKfaBJlBQkQLMmm
X5xl5PGgwLW7VMstutq+TTgeFcxc3BWlhzgC/t5U5eEgCE8GNtgitwy/QNNGnS9x5nQbUvuN6emI
cp3XVj8mgWwYbY+dd6melvvC1fNQXCK7VuPW2pKff/RlhXfek8z5NGrYdb22ozcwp1lnvpaCbHLq
+3eMN5jcQBo6Mt0bTogyz62PMBo0eJaw/QQoSBBmUDPWjSgTGuLu2TQrPTIXlWwMiwsJ5MBlRLfJ
4AAZvhfBICc4JYRCP36eqZ7xY/oQ+T9q2VVmvrtFq7M1s4cfUjvOuNye+7GZkP19iTQA5f0M9Zon
sDWEs0i8KvjK24tAx51tA35tCSncjvRWdhGM6DgMJ0zsg5NxZ6X0Sak9wa3GLanpAqLHrxDGazAi
L/ZJr5NDebqYgfzGWPAcreuhVE8vUAQ6iOZh7z4DEZ+je0l1rm0sq2Ri688Ez6XtqUpOvlHN9jne
gw2n2Bu+R4Bg1zeh/vbEYvypAR4zhdeYRZ3jxuTi05UBvjdyO9G61rAXMpBxGLQEWWojBP59+QxP
PwDXi/Mbac9oRA143iIPdHTyADbQfAWnehrA9TAmmS66b++dBe7EpEq40l+YeRZxAjKWBnnFVC4A
37RKZ7T630uA3t/ABEXyY3Kk2DcQDMfJxAvfxPmxU6/gDKfMlRefaPAMOH9ClJZUblsI55hdZYPm
Xic7YOPWRkVMBgCk64PD18xXUvr3M256NgVelpIXyt5BnanaJkh+JsN4GVkMbPSA1G7uRojtNr4a
Rypi6W817mD1yACmzGTq+wseHJVGcKuuMjo6gBwew9WTrJtwXCGA7rbG3IQ6mEiS1Xq5YvEU1BPP
JHuaO60CsexGfJhaVMBeOYGQySqH/zzobCCX0NrD0gX85OhXa4B/oLldbtyjMWzQXW7x4KDS6i6V
D+Hypu/uskP5H4IpgMaslij5ynHNG4UeVrjjTTMrm+HOQOpfRuXly2wDydBrfTG2XQT/Yu/Gbw5q
/8kV7dWTK1pZR7fcIa1xNiOepyyemz7/J5lI1u1aInkWfW0wtSwLCPFrg5UMd/6nNnRaUVxiT98v
b3ugg7fmIgyb+b/lHztMHDoM368R5DPtsOu87W0olTyAegA+Tq5VBgf7/+JN0tiD34BQZ3VqYg2P
ylsFXFQnoqncYkiY8wydMBsNmQ2mIO0I0kUoVLw7n6nUIU3OLDIcEQfneiC9iALa3xMixMyg81Qw
TxJW+pAyuem0dGEW9eWHaTIu2m2bZItxjgH0UzdeICmRIzsjfDZ3U2I/Dow/mjMNe38cWevwXH9W
EFwPBdg3CTuA8Tt6aB13mbKVUglskpmyFY0P/yLeXOUxmXmKKwru3sa9bJHr3mJ9qES0tIQV3Oey
x4hGS1+wGGCxkKyLb2xR+aQDWJcKgeoC+DUygNrl2fCwuci+Ezer7we3DOVSpyBnz/0Lc0G9OpmL
OUi78xI3ALBwg5EO+KAfXiHyIi60cUUj6HQ97zCPL6t9D8DgLfdMRRmw7dgiy7UKH7sqUvKH3pIm
WqCHrUWKWtDC04V1Ji2ZnB2moBw/WGHy4Papo+9XtDpb42ah2CK3CD4tY866OKkRai9jCvcC3eui
DV2caHK24SPV0FxLHq/blF13uV9AfxGefn+GLv5ZkYj8BL5xUGCGe05QzTcgHhS6FCT7Ae5aM7P6
k0CcCbGQztbTj8bdkYwKestkYvyldNPo3e94w2is+j35rzImwwvdkZLGR/SVGoV+cUevh8ODRP27
zf4kzcKqbI2+Xln2dgBiC6V/+AOkAILLl3Gvy6Pbh9MCbrCghBujTQzr0ucXPSxdxN7YIvuuUNIf
NcnvJVw1E4jjIRxqTUVIYpj8uvdOoMtYR7IylyjUX3x1x9q+Y7xxlv4iriaIBlEeitC34QZbyYuE
iUSprNe/GHFIdE9vOHniDxudVqtYC18GEFpa+VLYu5aNKFDweyQMCEXMZE55F9uw8F4ugbBUzS/A
jNVl18kt/wewncGEEtaK3Sor1uCm/VuYaxYdhsZ7PONkn4muvO+n6JoCnYkWDsO62yznzivE7jC+
g6APbbMklcFOAVy/j6cgeHqNKqwuhnemubFDk0fkSEqHPqfT8z5C5U+aHT8UWfNQn/BkCH+tHuhm
NvMxJb7exeqCCtPrLQZZ74R9/j4SjrLqeufcH2ovNKpA71TEQ7sCDVR3LmIFUxA0fA2BGsMsTBin
sQP5e4uQ1H0EMF2EiyvoM8/hDPn9vtcJoqDBGv5F7u4034JCJt3ibrb+xu6Y3IzCV1SrCBvT3V1d
8PIQb2TOxUR2V0f1yq7MuxTVj224X3Ayokqmr1I66oqpKgT+waqHBktAoMvDyo4fIk1mrfKrtnYO
1aTWOlLmjViKtgPeh85MGW+qaq7W1jFqkPQt7AVgKPsvJFO8k+VZwJQAthAe9SVBjsFVRK88QuJz
FZygmTn9COjrHVVaFtVASHu/FcG9QOvIVYkDdVbqzq/feLNSiMFzZibVZIOQ9aViE6jfAgPKyEMP
UlPHpl1myBmyNjAROsaw5BMu9csx+ZytSor1X5SVLJ/R6kXPUwHgogpJB51AUMHIHArnrxpJRPmc
MGaNV272q+8DzzUHorVjZp2dQTI4xT/FXSvsDSqT9YEiuF1AMWdfl60BD8o9DoKuFCwrIo1UT9eO
+dNHWJjQgba4odEuFMRAv7uiPdilDaLwy9YHGdj9+nZDKYi3RhTpeZtOoHoVDssCwXUJfOAyttiV
9RWAiEeJWzOEhkroDs0CvZ4s8bVWS01WHT86igL6Dk8Uq/MsGpBfhCnUMGvGkK63/gb5UXx7NI1/
0Xp6uJC8lb+xREwvvi347zaE9jZ0E6/ZX4F85iJ/7M2yVOf2ejjBsXFsz5pDdt6yXxm789vWo8rW
YV8heCkGBar7uMKTaCdbIULA6qnc/Ie5rheTiVGX9VOqfaDFDzbNXF/2xFD4XjWdN5yIlvHetnm6
vtUS8+CRYwcXH5yrBBxsaN2iNLF2EUen8+9USCFlaB6XlbhdWJIq0CYmwEoWcUF5YzULCsyYLEf/
0m4f6Smajx6YJC49L+UOKKdL2xPK21fU3+oB1hP+Kz5+fD4RND0dsgy8Wvedhx8OSv8gfzX0TkNH
aSDUoawlohdvhgDYXPEof0XgH/YP0cTj6U1JTwtX87zmfMdvMssBhwmcSck7q54j24S9ClzaHOam
qxjAnu053Iv7wPZ4oH8A2F9JdoMKBrE3rbtD8Q2uXeQfcqKk1JuDGjG1T9RbJaOmWlrkbcGFaP7J
HlOofaFm5oeTiL9TWFh7YiP3SNCIdU0uPK/ccnEzUPdqeisSWkgfnb8B7njihUXaqdM2ZSJzFR4M
XCv8uKg9Y0NjteuPGMEnbEaCtprTy4+cvZxl1BYSIsaTNJc/wtokUcbG4gs3uYRa2OACt8XZzZ2S
NvEVr4P0gckJ21peONputWqnerwK8XV3Lx5Wu20oCcaqwG8kUASLW6F8yA9GnmAesaFYwpMEcH33
8gVTQA6LZyF6dOoik1JHphMMhVBxISyu0x7p+5ePNx66vQiI881pqlOrmhABUeqSUl35AHa/sJD1
rJHU38LP03XU/ky8udjR7bQYc8Dqgi8pwVTdpoXce0+pg+DF9rSAS0LGEEFWYcNS2iAISIL4w6rM
JBarPWVCHILCqYeGF+XFM/db8jWa7IKGvWWh6ldsCWEOg2wRQvpFtcLurBpLZ/sQXZssk+R9pnKy
Qs/kIHa3CFGr9gWue0LCloW96W73ISyan+PVtbxlW669I6d18GS4OXqQu2o44w/zZay20pQ7pmCk
nF1WCYMB416k8MV8hea9joEhST/G43Lluggh3Ghe9GZRD2Bsk1dH8glO9XqmQBu4GbpFbWjNSFKz
rF8jjlVWHRjNb7lyZO0vPYf42Fr9QU4qSrJKe2bBIBFoc6798pK+07D8XxzGx95buIb78X7N31mk
rvMr81qDj6GT9nV0UdSVBcyqP3m88VVw08IfX0/1REKOlHtgijU+DmgzVVbl2EvA4V5vq3NR+q6C
PceF5Ybva4JaVjpqB+fHy+zAiHhWIHuY+VBRTDxPdpHmmPn3HPUoHGRmIdRDrqomsALGhUihntN9
8jU+cyJghsxnhKRXsrl5qgSF29pRvcuxO3eC+pG8yGqxTLiSdSNTrriDIpdOhIGOkMRttK6BeC9B
IKZ85PHapYz6MJcLdgu3SCtzAvevu72WfMRkYw1YxqHuDkwro16Vxg5SUaoJfvXNI6eZcT1t+OKD
jCHkJjOdzyaf/Rd9zp7WawEO9N1C6y4NzBH+rXqaq6mVWNQJvRr9FStvfbZ8VHt75QCQb0lhg+BX
c0Q6BYtKAowyiwmCN0kjGP5N2jmuybWptgM/Ot2tglZ5l96/dlS3oxG8G+abKrlfPjHEmi7XrAal
YSm4stZnNFtiebqZCaWj44Zn9U0N13jl1dRWo5RK5BNJjRmKnN1DsqhF7ePZ60qyxv0ZWUmAFjo4
c2EdnzuBLhFowGcYXEoI4nHe8xm0ByZsV0w6kDKOiv+4gKdzLHTQJryFhae6RDt5MrH474OTqAEs
Dk3wuJZRr/qYATlxyYA9hnpmoRxetYtfJ8wgf0tRlAbpjFHJn5luR21NAP/IPIyRc2k24D2PJJ3K
SbkVguaaF9ntbCAozE4O3upuz1lm6JsUjYTd0kAw5oX4zR4kYkKHpt1QC8gABGpmQMmyJ6w4UBHk
Q0ItqbrIa1xZHHW+fdHe7mTErNUCAz2LU8YNHa9JgsDuRUjGI/iIbTFJtMNuFNvGTei27YT+3NXd
KRb8dYOTdUQuLr9snuRWHzMtwrqH/S54YZ55+ASBmYWWEEYYySRA/voE/sNk8mTh2WvCcIG9FwA3
43QYVn8z7oJmkBqMGm+lm3PYOfKJdF82FLl4SCLOxjcapKlrRdhih3OzUVURHlp+y/zXR/LGesUB
VtUgG+pVBPrRBRzhklX7dTFUHsCFUM2H/kprgmpPMF3LeFqy3MHbEtPUb5g3wboF/Ch/tfr06HEE
Z87TtURuwljDSwxX8GoWuxnFJaz6R/TptqkfjadCNwBliI0+MkTj6EwB/Q6vgOOleYXBh5dGnVcn
jiuUEMQHII6CJsDnNrA/p+Wr3F8RvrzfbSAK6yt1QA+YHg0iShY9WFNL2bIAYv2tPFjXdBrLydWj
uomxE2URUGvFEUACSJcnbLuiPU48qd/j2LsuuGrdepM842X8vg9oeegjoduZsL2Sszd/trk8dCP5
dUzgvnm2sdgrTiqjJ24W/bhcGeR/EffYRIJyfVQkiJ8FNai6Wi6cu2WCIe3OfWM2m0O+uDmTwaEM
ZUDGjNIWUsUJSvip9dRL9MMoIdeSmqTEl/vfcyZbGwhZYa58Bqce0lLkmG8RUy0rxi6ua+hpt2+s
DBFh9WSNOWzOUwHG1lmcNshYdQyxLo3P4yG1SccTy9Y180XEPrf/vsgmbgQrYFU/EeiF0JyeB832
3fMRSTZ3hCideMo+yIVjnh8Guv4aYziQne0mUsXXXGXGdIcTLcCcdcxY05W5bY1AIZTKFDjnIMge
B8aSg6oYoQHAnH9mO18Ngx+KcN+AedIt18ydE1Rq1IK0ovrMw2OSYHKriKWQCuPcIjL3iBY1RScX
7KSW0KzuM5Ea334YOhBnf8X4MPO97fQIslW+8TigCIqlhR22c5BL5Fp/AmIOxFLXIaFJyY1M8bhM
bVOWPYSwUOjEu2zfwy7UUqEY1l/G0RnDIebnZdgZvO82XYsa0/DWnf+S2J5JfCpWZzGTCe7Tq4EC
buboXctq/GXvPPz2TGhgTbaBWcOBdyVIfK3x8//A+/ZFQL+MDRm70RFlT5HGAFOerqzqL1r8V09J
+pIuS9FvWINYWhtWPtEdcOsoWv/myCQJk/mHcGqT4DDdNYkv2Gh5Ti66rI+vLKLLE7em1JX3R82R
6A3Geg7ZxAAcOYmlDPuC/L9NS9ZhRIeo0pGOzUp0VsNoB/xwKWzk3r6f8qyaxABd7N37cl3ZYvU1
xlvvfK9p+IN9aDii4Cv7xySKzevgwzTm3ELyIj+fl0pgCGX7zuGiLHkhRQpBZfJb9ou350XvVvnc
L/MN5ccYePJJKepas/ncxHgiKQxNxNgcFSPaEV7ojojOxCns8oaUDH4g911UOicPvtZaCdLQKanE
kYaEva+1Iywc6lpgGbQvf4Pe3vknTbtGXKH1E008FMhkTcX3+/2LsGNmSTu+aGt/9kaEyWYqFips
Ipj4+EUglHFMB3rFUdHLByuAhBx6Y7NDPqnoOklJEZ4Lk2SJdspNgRwspHcpe5GobpcBwYi77SBZ
dWtw2fcTwonmxPzjeKLNtc/ck0p5+YpwX8MfWLqrXtD6CQs/6smEulCpz7eOfwzUVVliv1VvkXD4
bFuXn4dgi8TGTMtTgRGjJqxlsphb/X5yZXA4UddKbKXRX6A9xnQHEzn/n6Ub2hT3CR4Op7l+z2er
W2IC8APwr5IqJL2uJMoz2IhaPN6yDkmINSvgLW/xnpn9sUqaLPYKDWRhK+cFnb4xN9qfeF0bop5q
4HPp32n/sB7I8TUyCJzEra/9XykcqOopfz9L2sGRVMJpZqDZHqI5lmUFri3GkbN2RkFU0d7pgPws
oXmeiJHEH1sSpfhtf2j2yTpBX6sfAg93opAwbO6wJd3a4dfOqwxp/RVpoWD0wsD4g9MFcjsxyOyH
CIrsxvkHBL+UA4qF4ZbjJcPLhnVY7IVrokZ2+dY5U3dcryA3ZO6K9XJrVzRhSTd/o6ma1UUhgedI
1Vikhif5FbSuUnczsdnyEVO2U9AOhlE0it0Z5ZoZxditeD56whDddij4nxBnvU3LTgdFOGGQ5Xdl
xF0G7OK6fvfkaGVP/xVsk+uFDLjL0NMYbQrAU/QB++b/uNp/5iqH5ouk5I0IDTHciqZJlDr+kh9w
cigbxfDvxOb5mq0XP4C6t5r9NP8uWzeN2SNyJ0ruNqJo/BbJG5tWco0BUVIs7nbxj9Ii/Sj6mib4
ApQ9QfdtDUSZ5ukg4DkVYkG5a7Wu4zIK7llb04zKoE2gkQ+ZSkJJI4zLX6lxVrk9ko1m6eyVJ75e
RBM3iYzt2Mk2X+kw4Al7iHDlfd4xQZj9Lx1H0N0hINZ+d5PShZ2xlpnCGINCwZVusRaZpGORV2yl
cS1nMTcsh8rucw1OT+JwVoUPhKy9MKXMHNK4AhbBGPqjS4pQkuAEcYzNwj/gfpj5s1MNY/zPYWwg
JaVCGC5yO+khrMCSGUuxzU4s7cUnEwUufMfrK7mKR2goORY+fGZu4qJO1I6sAaPqAIIvsv4QKA9j
YT73QdmH+lKwFndZX8FsG0N+WBH7w8BSch8CvGS+p5AYKw9Z0Coy5eS1NM0pKpGxXFCBPFdxD7Z/
lVYfN0/2mQ5i5qFZtz4NJ2tHTDpQdrYDuHiu9Eyo3KsnAEMWuKLQDLTb09/7yFJ1AS9JPiQXT0fg
OdUw1qoGKzd8ZzX9+emaniRgciBRTE1mxRgc7WyY6b2E+GBAf8V55FS3hgsodhjWd96V5CFMX59+
6yn4b+nM4mT7N9vdvfkbfj00dMb/rUk32pIHyMwnDfTAFKwCo+xUdj+dKHKvcZITRanVHXF+0n6T
JoOnIepb+vEFG8HMrPhMR+BJ/5QqY/12KCdr8T69TtPu7UjVR+LQFh5Xljs5oBfBeYQLe7UtCwPa
xD+0DS6SkX19+pYDi7mpF8fmOzPrRtlVRpW8dtPkoEFx7Ufm26U3sOBe03vkCxRCGNXoyo8gkRnM
HUVSdu1nCJwWr4vMP5chAsQ/llYV3+NtZmwqv5m8ygw+uxEjGg9/D+RpkVW9CsYJBWIm2eWSZbS5
LWFqn70dBRJy3jbpmYcgL6skkY4FIcdm851SLyLChXyXWRW+Dx2nhrexYxxGjtVluq2n8v6Rvils
cC6Ma9uaEf9ml3cmyz00qFu5hPBLfFMH+gA9DhrF0otrvetOjY6niTxTvLl59190H3IQuAd4joQW
tw5l5E/FYc3JU9L1+WovkPPL6hpfhoYrt4WDbG592tGXocpmOGf5CxO5tqF/MShx8FRP1EFQ/NcU
r42Is3Jgu5USUsJYT7LaAzo4sf0pXIktN8/d9pW7Rds94HC98DEMGNUrb4NeGXe7Vypsllq2y0GD
zYLYTnZuIGwlxX9figvy8hdPbnr+oITtNN5Z0qpiGd57qf6CIBbIZNoCwCCr9onVvnOwR5eBpbYB
UtN9+JmMrvAcIMuEtz2277sp+XD15BnDTHKhAa8XKjPZIRXgBsGN1RSklqabwihSYrcCXFA5zljp
FubMdTU+dyerxhZFaZnk4Frb6tqWupRkGfuwSZW7W4k8TuNdyaHtEFuSMd1/DliaPa/HcQcJnbIs
hh2eG0khfrJG4BwFvbcYIPeg1Z11r4SYYYqQ75lhDk/fJWyFOtaJJc/Y8abYvvbux4Gh8FVLltKS
nFDSMXlLFOkQqG0CRDi9euH1lwBhAuJVDnquKz5JYulIXWw2bSzCBKc2SziFK8tdgY3jxVJnJOJn
UFj1taoyX2hZjG3v0pNAC+r6K53+cGixkHSnQuwxLSWO0pBDXIGHlx88zENBIkLJEhJMjDRg/+/G
D8f3pmGbZ5ME9k16pKLwa6H8lPRutS1/DUIK9+JmaomuC84cpE1iFQsfzum3PEw1Bs7z+paaF6vk
fCwy6ZfygVbQkCYcRW9zXWPeN3/P8vtUI7bYHR2yzByDg/8ARqllJ+JkzDyhhcAZ+4xg+REr3hnx
Fpd1NDsV6awprOVaA9R0xPM1M56HrBpQvJ5KundPERpEsPIF0dId4yvPLZQXxGjTaFuHDKniM/X7
G9BoRoLUpysXUreoVb6CkJrT8MJ5nXAY/MLnUjmNzB9cKbkvJTyRShlOtxEKt5jqNjSiZKzJmf7k
Sf8FoYUk04OeaQJt0HPaFs/o06pX64hgAeBZIArOYpcB2XmYwZ6sSaf0cYnh9dQgiwPbu36mObR9
z5h3+adKdvDrMQJjXdOGdikRa4/x1NF4hQTU1lum/ka/LfodtmU8T2082CvHIiGqNtd2uqGFtwXS
ezfIn6FBqhqG0P9nmT6hO68uYpXoY2ZIBG8qzasAZSu59yWjQgvxyTD4XyclFZrdVk5XetAA+GnS
NZE744yl6nm08t3J0iY14+RHUPZNtZsIo0dOnv67wa0PqhRZj9BStfxLI1lqWF6Xjso4dVEG0GII
ZOyO5EgTHKfHxvqJ0XJsQWiwsSmBzQtCaw+ZhL7YVoxOssYKpHRl/IK5vrdM8Cd90M00Xrd7tFbL
gCyW2y88E6iwq8CD/tH2/1HSP1rjq3cyy4TPH0ifUdetSDWT9KvLJtHq0s7T2JCOnXdGu3+2cVQR
gqxV1ZX5Evlir7QQ4WC3WLnPlQmvITsR1mEQYX9ctxFJ2FIHJDY4PTHk1XFHoMTjidQZ1M/xxcyT
6pKKxEr0RKE7HQx/KaHaMfsRYft0AahHWVx+qUDVy5soOOcYVeWjkGiXVs/ZiBjAeZvRseuc3j5t
pWSvdtaEtDQAlPZpaf1+do9CL9sGcGxAbPg0J1J0rYVctln1+fVZf9DHPmv+hnzUot//7rmlq2a5
Tnv4KE0CP8R7lD9llRamkafYiCB918IyWWIY+qa/1+1A1rvUpGomrPQqvYX7QSAdmGzx4hxrJQWU
/jFsIy4I7Mz2twjaWHNKfjMGUENEB2QrvaMQGWBezbbHNabn3hjuEVI0enWsbLKq13ESrGJaZsnY
5RBmELVG6ZFAWwtSDa6Yr7IcNGFMhY+sfUO+TEikvoU6JNx3gttbEli7jHOG05y040L16lFcF9K1
Fnz2rAxZdwMwiFdEpnVLFehv9kiDcoOMjsbuPVcDdc9qGfXWp/j+5C4ZSR/qf3DEIMcRjMhQUNd7
LZ/HIJqrViYqmB3fZQ6X74VNBjQs9hfxRAlJRgz6hh3ivSadid4tkz8lP6Wum5Xwerl7ac6CeJWH
zZdbwhPmhkH9ugoJ1KLnvnYhwNSZQGsUEfYjiW1TfA9rfH0F07rJJSIVPn4OwsbPJzlbmXtOVASM
dTyUBOG9Y+dmsZQeJYhKlP1NOEZkCEhVRdwB8dROGWF++JmWuUaTGNuJl2slqgILGNX5bknB3ojQ
tYxoSay+tft3UiGT9nei0nsX9vvmgL0CQmn8Bs8LR75k0ZFvowa7tiOeE59Ka0d9X5hFtaVRRs3+
M5tjy6QpPr8hQ0h6rABHZkHdd5/JLFgxld82TyQC7vF13GU3zCYXYcXH4Msixh4cduKB5bAEWjw7
W0ew8umJOED7fHxI76FkFLKAoGaRQp7UGm2kAAQBxtT+XBN35Vb7hjpIdsRvfipCTdIDd1I0V80x
odn8QtrxR+L2k6pHRSrEpWUvri6oRBVETrMx2OLztmNbTy2qMSCz3tEQqCfzx0TLtcKp70EMmxWm
HpCa7Kyx3NahgGZGdbb0FMqG0ZxixNoYKAyaxDytkciNFISFyyUpO2Dfic4xnmibe2+e+T3yn2YP
FQyqnDnvfl1T+3Wl3/mXEavwaCiNSpcGGU3lgG5NMBVMuiNPiYjBHkkGBhCpm4p7tYM9ynbv5YC2
YYB/lxzwQrcVmV/lEDyWgllJFtCd4CLr8at1xi98fVJP5E6KO6wXVbvI/S8V/vhzhIf5rbfe5sCc
jvFlQhcV7fx1xusvPEaGxleQx0fJm2jcYXmbUDJEpcpPLPrwynkOErX6ogcL0SNW0t5VOxR+ZGuU
/YebCMkv1crdCLdzMbTm3LE2+5peqGf/nAIzgTcuN1/miFN+NYbwH/W3mXRoRXRdBMC0oFnjYGd7
n8m68q5Ss6FNtvixNa4bvFB74ENwNzPj2/pvlZH8pn/eUUjuNL+OykoSEn+XD37zckpvBxQ5Y4sw
jU2AV4qohGHrIakKWTa8nEUtic7eyurUy/ACbWgj/4qEEKZQEy05nLHZ+dKH1LjupW7D0CB7ceS3
Knc1F2hvGYpaRxR3oZ+KkJhLXNmE2uZUY9HwQL7ucqWZaQY759TI7KbKjk08I2alRv7+bPytOUWD
GRygevtnxzQfbptrvgIGoNwdXVPxybSg17B+5GCvtFGw7Ufcev481ayJEovfzHL7LvH+49yHffyw
zYvQ2O4YMelOwPuc1Ov+1l95XrWI/ma/s/9q0Gou7N6hxs+1SlqtsBt6klwbvZFBJiceXXa+hVCJ
+sEBgqconNMUsFVYCbZbtiqEECeJjdeoSL5ZW7yZJAR4kg9yNSDubrD/Pum0pjgYX3Sbm1hbsAUx
fOrA8KHC9JqQXS4yyMa7Oio7xT3gjmsYnyYxv/PDlSAXLJQBk+Xeco4ZmQY0wfWCQQTKlb3pBROM
oJBRo2pr3dVhS0yncMb/SwKfMNSsUq6cwBRB2g3N1/eAC84EgEB4E5zmnNXIkY7cf2rcRxgGebMY
nbiKncuqQmpwL+/4qUMkUe+Cwp1XDEsISiN7SHtRmEYaL88UtUmm5a1Tia4MiOIMS0R+fQt06dcZ
kZHwgwZp4ACqJw9SwHiFI3shPOplsf6WlGzQ3iSLVg6mFWCmkYSn0aPrnBgSgXOp9IB3zaXCDNd7
QcI/mJ21BzsY0mu2NMPV5tjP04WL+Kz994YUgXwpaUCN1+fg58J1+bij6jByvaBif99vGcw22k0D
r9YRxBk4Fa/yuF2/Utl6x3fol9yGHNq0E41tpgqAauxV0nvf/zqTbsIuoaJPVMZjgQojDR56HxSZ
sY6vkhjBclqT6lAitf8jkdzoeyENOR9myTmEiwqdNSn+FNNP9ijFRa+xjSzO4itRRi9Gz3rsoYwV
fnQjpixkvCldHLP3iW9XOI/d4FC0n/a7TF8Y72atctZoR8seEwTrpSUlDiIgrtf2mw0EVkRaGxqd
mkL0+bhOBlk+NxtI97SPx3ACsJE4fRGBiMoF9DNXaCzQdNCh8kgbCV72xYMz2rA/cv955fiutw+r
E2uh04D6Yicz2O3Q+HRSbb7iVzTWLDrJ4gSmkuAJF2En2iA/jQMVv+I1sn//Vk90qLYGUipIpSyu
f7WxjELqqCPGJCaJ4HRCWXkJGzF10uNmkiXIaAV2g3pEYjNAwUUABhR8acjnMWH8FDewb7MZ6/BD
Y9UFRkJDVuO2t60Q4iGIwD/qd8I6DlF1b7+FBwWtiVTnEER1tF3aS/hu59/pS/hN0rvj0v8MhpAJ
w/BlHsRhf3yukIrwO0nUfJXlO3zVnUHWHv+kasRW0T0A6oxGJutt9vghq0KxP4avnrjm55N3S8Fm
Wc+we+2fpYx+N0JyxrtDlm3mtEgFcXA4KNy/apJ3a/+agOAWMOb4lz3KkVVoCtPEdKSZ5Fg0eqwY
x16kwKJhh6WSErAGxzwXU1npeqYAHjs4PAOTc2oyF9dPIbyvwQWx1mKC3mbPzmhTol5kdDoC/lav
H4B8NIlJZfWeDySjquyx+90aNwh8oOI6Wie5SCWOocFsVLB9z3yGA5qJXD9GdrXBjse5e69UxLxI
g8hiXUWvMf566cRnLMdX4Tn5Ft4xfbrqE6CeiioLWYqZ87moA+nwOc7qZYvBsciRbyNumWgFL1Zm
bkQyEnseiRb+rqOBOHs2BANgCWUHWT4wZSnCDQhKfSBL97sRPZ83r5MxLt4PL3n0e6L8j3Rb51J3
fh3odC7dund5j1iMwW/+wv/+U14lF7X/hZ63fdsg/3A6GRyRkJxl+dPe7V1onqnIVfSnLg6W8JMd
+nWA0sfITrYN92wN8u8LWixsBt2XFVFEGd8nBDhULGAwr9IcD28xCntTJ+ZEH86gQqEN4LL27z2R
+junuoJ1gUDL2dNBzldswdsflldI4oSingKJF0VxU13ju9akUtKwBa5u2xWgnoMVK05Z6kNykEV8
rCm/xho1h1WQmXwAuTpcNncyg/+VALfB8gnf1fPSsxy8g6OdEUls7TW0hCVecbrPq0GXlPbIoIis
9iTt9LeDgqCiR5/3+H+MrTPpxXSGPP7V6giqyoY1u3pCxlo4wKVAG1ZNfIAd0HPLvqq7kAi4ksoE
k1MSp7XDd53hFHKAEGz5VQ2gbXb31i3rjIJGh+fZA8TEPar83MBAukDltlhx/TtSsO6h+9xSe4Za
Z2k0xk0g/0IFvSjHzNkJQV62Pyq0E9hpaiH3vIxqVcpndKUe5Z+kse5xFHPNH92iuNv0bhfqNX3x
7IfGWmpVOWkePbOKIgd5d1rEBaq2do6jewIpszx29zauXBmKagpLlqwIKVhFagFHmc54tUGDHlio
vHtclRcY8lf9hw8yJsXea+yO2b2aZ47g0KbXvAAUiRWwpLhm3/OIJ3pQuNDsRIKyZm9q7aIeiXzM
1nTj6zIlIwIwBZaQ2E8d7hy87O/4U8aCk4KGlm0q0uSkwfPVxHqKXMfw4Ctjg85Mjb5GfvDs55Bz
MB6q09GkvcLxaDcuLmUI4Lwx0fQk0hVwbcskYBZPADYdVv6X5BinaLXA4uJRsNfi9Kzy7r6IIybj
C8LrOBsb2HVx8KLyxPnxTH2Jpm/8m+DBc7/q2ji3w3/JxKE4NehngL9SCoRM4gs8zh6iD5n7fcUH
beAxb/Z5SFdxwFLsiNVO8Fo4iIXCIY0bosIp6sUGcNJZuauR8Bo/PYLKR6zgbIQ0ibIf/Srul4XD
IeAqJbwmBcOCgaSilhxcgYKsUZZZiYoNnL6S/xvDHMJyBoLuCRmYZuNFLq1mZEWGK9tRC6xc+9Sm
bciPruPNJdu6AsyWNF4PZfzREEO0T4GuaBc4pQwcJ7tk6P/0qdNF63XeY2SJN9fAT+J5YY2kALXA
3QGb3eUz5x9c2ma6iruxYwgsnCfkSFFkQORvbXGLGZdYE0EVcOeq9cBwErEw+f7gSvzn8xXuOgq4
EfjyLwngDMeRtHtgWzp0IM8Kxak9LIDE0JUgrMen9FigMrRDJgi8G6aqEt5be6jCjhHb5w6sLZcB
IyMOKvYCqMuMnhbXYjU3OPW2deaDk5OUp8D9eJ3XM8s57WihcemgNX/5Jnehm48igN55kIrWK1J2
LjCLV/kOPbqowt95yB01+22ce2nXfWLGkW3WDraH9+XDtwH/4yGDUav+vfGaqjgpW23bk60JvSYY
p7yOp5M3SrljYy5gHTedqnYqE1g7qx+tYhzlljGO0yUCjSjyTSkIIKG24BAAuLmXk5M/61r6IJkU
9s7Jdx+ImidNIm1Jj9DRu2xRXiJWbgiZN2e1TMLpIL0cgzKyTbWuZAZp0SPfA0xjupNs7rLCz1QJ
8hm7EOkmD4JfeD22TTpJ5tNqqrutJoegB5N8jTv2cEgvu2MYeAaJJMImeuTTq8F92frtQk7fAwYj
Ojn9K5xH14yPuxbmO3b9C6W5EuAKkjNhZGt49xfUtI2nl8fyPC2MLGKRTYJd5fSGltsO6iFsXjy4
RlD2WVEhplCSbBHygbC3cBw36ci0PDnG/5uJk/JbnPiGHjNt6qzCo/Gr688GShskxcXSZ+8hBbOb
S6R7RkgE2IMWSwKpTbNZoTIiddx2qBP/ostzJgt3B22fn/SU+z5tRVrRRED7LSLVoYJpQ+2hQ17W
UFTiNuHeMHzOhZrlWB7qBjUPyORU5BbfnGrfqu1vYr/6AvFzIN8TJkY+Z3BN0Ezb1RXYkvZ01cIi
wd3qnAOx1FF3nDvhTb7BYXWfLCDqieMQTtMQWip6cF8uUKLg9Sbs42dTKZn23468UHCLA4wre4+u
QJAAQQYnsX41idj/q1iu7nVIHOnX/EZZFkUGM/87MS/IXsKdAeHX+J5Ci+X5GRrsX+RF2sLyIVXQ
tNoKCb0GEvt+7TJGv0MVobY+yF5wq9JA/ZBhSGBru3FO7bF1whyhXh+4xt/2OXfvsJQtZ/A8nBdE
q6Kn319GUUu4uvStdmw4P2RfLKJ7dmBbe8ITHBdHNIcYeXnAeKale649o1cdudTDmngZqKM1xhNK
lF4lqh6VduJkAH8Jh27mASOSJtcouShY6c5vZ8dufL+2aiqoP5SGdsfdBgQTu0k5fyvxnldtoROU
h6/Eo9koI9UFV0TGJVfMyqOYF+qyEpZF79IUCgah/gdRLuJMABSxVoKSTiWdr9++6MAREcwqdQGn
U0X1XTlF4vgO6DnAHIUSC28OdU0TwwQbc2/qSY5YC/sqUIy2ceZcCWq3dLYbLbSkGWmlt0t8XZng
ztA0WU2fVkbWsXsHk0I/f09qvtLthYoVHfzxIvNfA/VPHKSkmVIKIHMhvD2QPkd38W1Pv4zvHStl
LMblufInOzEzQWR2Pn4BwDFkJvZc47s4U+Fcc+ImyQaumDhkxtP8HFf2UdpMHXF2jZfrsotKtpXn
+w0zsIaCW1hYB2AdXh16SOgbMRXhOjljiQpArL5uq4UjdKuGvCXiz6wzS+yXhsPWzoeC0T9DqYfa
t7+KDC0EHbVYPIBt6C5hRq0IfIK94IsHHOBFJG1UNJyiPhuyqBGn1pjRA/3VE35WKRDe/EULgVq1
7xEmPcUdd/sT6vdK2iNEplLoJ/zDlExaEzLJP9t3MWVQ59rGncpIMuJjUpWDVnc9VedcheisER3A
hirCXsyu3ANq+j5NX/8akAzTlHAfMDKkXTaWg7fJP3pkrvsI6QHwZNgQ749RgjPjhE8NwO+ZguSp
ouyKlhbvWF+bk0AK+Or6aODc4ZsjQh39tipk98PJwTfl22D72UPKq5oDmemR3jSqxF7ScyVcwmOp
/lvdFti8Z7HTKXfn9LNzPEtOWzYo0RjhdEDLEaza9Knna98kIlydqQt+gJ77eloA0UeWWavkvDJB
H41jP8JTBXVoaZyiSWlaSpp7Y8PmtmB0fAbk1fwYU/oUIfItjInXthfIZlLbp0wmef/flMT1wFGd
Osf4UE1tFlbisxxaIWbeWSylnEnQZv+nau58rYH4WRLb2LF4ZL0aRV005kam4HLpXLw6//M0RkCg
RlmB1Ja/B/SuqCDHhvaXlIdk62sxr97qAUAr80bc+yJ8YVWl4FdoYN4me3gEI7oSCEHkpkDFfejd
o5kL6pyFALUvVEwS4zzteKlDqHfSxpEjaxxPn8QOeA7UI6bASpqDlv/Ci+jkImoMKwm0SDE5KpgQ
6Ee5ltnSuUydRPW2OMi49kmNTQQU9kbxkH0fUH+iblmXvp067eHDs0sw9+F6+ByJFqwIAIIdoU/M
FZex5CbN7wHDfwqO4jtnkv/Ila6BoWKK2jeG94t1TgFf9svUieRKZBsIk9tWvcGlrjDtV7i+cek+
tJ6PlzJTV27s3DXcyFZJHgMtI6zcsGb4QxtzZeghrg9whsnXkjXZIuzsSjUjO+/M4RstvuR2q4hk
qhhmLLLGL0wqMEdk04+uUe5dcKrgixkTroVJMHhddYb0E3MLCHOEPpUhuH8FGbOKfcseuW5r7qLH
CqqiYxmRgkdzklkqEm8M0SGhteNN/rTOWw/+RttSf0Wmk82nXMbOc9ybr+oGQL4gx6BdPkDonBq0
KeK6jrFBir+wehDgrUUCKEJnhC7csWpJ5yEkzCIN1cBAGssPsPPfvvXxHsJzAaOQfzPoyWB41AOM
71FC8s/by63fkCnnqZmPkWTyeGOajh9qwVxFvwDEhsD1gKx03SrtjkBDHqYyVHJ5s+OBacAWKByc
WtnrQdK5gDeDy4Q66+i7jAwClSNAK4TO0T6yeCerR3X9e+5m7l+FLEjJ8t9Gq/7WT8e99stpyuqZ
a/Q4yzlfP/BhvtIFSo5ug0eS5dUQOZrU/xEIv+EdMX9zZ/P4aaUqSxt9G2al/R7crnV2v1mrzbYj
w1N4msCMLxL8ySFq05MlYU+DzQL9vdBToY9FP3IE79ZLB9RkwAnFIpRUvm0wiv7wZ/2DBzvmKNq2
O5i+51ujoykAAJ7ZR9hdVgYAS+wgrWFwk6GlhYI/t1o4D4eWPSGw68tNhYh6Z6mRiuUyNT90DOAf
CNozVBSOjJJ5hKMt2eZVo+J+FCa49q2+reQqWhl/Z+xxh1mtE0tQFdOIaeO3XdUccuDeiiWpuFfH
vsSkbecL2xq4zvKe4eonZShrF28FlgOVGeqzGpqJo3xrUnD/o13YSbOb2U5piOAXpyb+j0BacxCV
QV0TiKt48hkDYGwfzZOQ2uArOoePeY8IRkiW9mFI4rWKRynrX3DfEhZ/aDeF9yp0BlNk25HXsW+/
WkL3XLAHTnyn4g8NlBItEhc55usHL/Zcquy4Pn8FEx+Wzr9RJk9Wa5ovsYL5HLnFk/VVbCTftZYb
WvW8p8Wgo9vscX+9nMM7ugczP5C92O0SNqa27jCu2Ojww4U1KHz2HgcK8p1eiLQOeOsq1S68O7tK
BNeQQYxjlRjlhhSoMKo03bSyF+z4pVl4SEqpRo85C2L1bW9Yh0+N7R8UMsWBR5nIfskeTtTWao/v
coLS8PeIQw3f0AdqjF3YJPeEa1NPHRflC1VN5FmJknQaB14ucS1jXiFqLuVj7Rp7C6iCtkeYfk49
SakivlQvNmBIR9hWpdfvVWMQNCtdOS/18Y8RcwMG2pFD68S0XTsg/bJZ88kBf4QOhWd/MmQp+D2n
HgYQbMU4h7s7OuG7BY9mVQIddds8T+CSet/r2F5zRfFirUVRBzCApXzmAS6avxiv2FZjcfD0Oioc
BEN5M/VLH0xb6xuBODl2wQU+moBjw6oObF3EvqXpxwnyKPmHyRVPSznag13JMZ8LpxOrMj5SDgI2
M/PBHy05M77Sb9fOfprP0OjWvSaPwFsu2i9HKP3480hV3JtV0WKNUPZXlE4AsE3BXLADb1eeBEGj
nRujT5hNqdaBI+1kGo7q0Mz7SEtIMloMAlxsmH5R5XFJQOjwJKLeuB3uBWjYXX7563OSuHjQS1LP
m8N6uRx8libWRI/ReRdDgj4rMIWuczuk7y2ESgIkzHrw6UptgdWaldkMljDJBiuY44LiVfC4k9vY
DFl3AAc4MIz5tyvdmKXvqAWG3YhFgvlfe8Wfll7PIkvpTS19Mh590nEH0qqNyFX9m9PgAB0pt2q/
TVjie8Q7UayCHhd2QPqnMSaZtNqlz2HRTHpzB/6sA3geAj9wOeER3GMgAsenO1HaohBiENrVwBhJ
4qF7DL701sfN8dbJ+j7/8amJW6uP5qTrBoKy9vqatLZbAMRumjHNpzb2vlJOKEm/EExAdEpCt9ZS
DWeSlUra6ipTPKIP8CVkoInGdeJZoxgvmievvQYiCJJ34+IxL1b8hPQikabBv1bYdYwJZDKslAKr
B7uWmLzqlmWPot+RK1azTuPP2QJI3OFFur1b09/wkrQMtboe3nyubkxfYqi+jsQ1ZdNZObqCzzwC
0PkJ2PrXnSTMXAF3aef0Bh9dzajrheeMjgrM6yVgKTAiIfvfnxB56nNo7+BdKJsIJ0d/Hs2CHUsJ
OVZP6e8KyVlFkA6NmBwJrg1H3d4oXwXQ2WKyqgCYTXQMcFC7+D5ZYVm+jxuXzT8DW2xgfLV5UuyU
kxS1L/eb5tBy9XT7kRKgFOH0kQY+/v77F2ay8P1rKQHGAz5b9AfJSeQK4SSf6REkNPeXBNUe1y92
TnPXgQs6L5t1D6rFHDwtEQcYVPtU5LkliyD3hvuA2JSskOBIcUw+d0CWaRdG24C56DrVkY1pvMAK
AbQpZKW7BQCe2QuUH8amTVKuUyiDFJ+jH0DQ296vMOpuzacZQO8ImlkpSZI4O+aTzObNu5k9vhbv
0zzecy+4AEZXAapSRSFDc+dbWLCIol3/cNdNU4xCjr6688EFjkQS79MWRxXmMw0ViYs0MTFeFnWF
1BS1aA2Zp8pKuOmqHpvccDzAhYOJY0iJGjAIkC0e3YBlHISXDaiIy1OZReQ+1TAimlF1GqzyLQyf
5x2ZjJNBMvPAybAgd+MSUvbxxSVDagQoGEHksKo63lsNNdTpHB18WrHviOl75k5VdcB8EQw7uIbg
ecuG6tl9C+M/1uqKMGFcpF6SxYGjTdHE/6OrQTk8RKMiUFkevr0oNQiaxA+fCdScTdwT1fKQz+gH
EBxx24wbr406Ygl00gR2s889Mjft40uMOPDikMBoAvQLiQ3qf0TsaoKMLMPVRaJqxKZS/f4PasHw
8GYVLds2HIt5yQBGKWjK9Cr0iki/aGWqwyxWR1HgV5ZQkrFYXUYSc9bjTQCTdeDMHigvazKVyDMg
WGSefQBykri1YZGu7HhDr4f30JkuhS23K46w9m50kXsB6/6Lml+Cydjemjfi9fZECNU5amduofE5
MMHTeuewaCdZelH7rONdatrUYZwdca/n3dB2WuhInlfZxBYUYPBmRKXW1JWg9C6ltfkGxcp8wtFr
BUmIEM29S0peIJCnlpsAcM7zQH8ueas5nyFDlTDcrZQ1VVggWPmBYEY8mvd3dkm5Ez1NCQAvvi+m
dmn3hTiJj/RfFvAm3Ty5L1smwjd3B6dqK9VEA9v2IfqYuSQnd3jFQeTH3vMiShZsvZGxbYeYfa2f
xj6yjUjF0U+FACgz32SxwKW+R2gixM0d+K6/gzckRGK/6vegCwgAwncWb5UXWUGkz9+iPzlZJ9za
elVm3wlNmVLGh4VdziPGfdYKZqiBTPGkdVupuIVZEZMOYiDFhb2R8Bd5wWEvC950hZrVAk12xH6Z
9NLo75jVUte86ZhyXo8yEu+VTW+EMbn//mvv4U9eedOc88PCqgKhkGZh30sNxqwOaadMcjLBUDEz
IslTyAmwcnBTDmzFXbCf/n9hC6CUuqhNxNApNrApcrgiYNv1jAr0Vu4v9T243HS1lfFXH1CQXLsn
7eDsmIrbQi/uqUicuUdKoHhHuZ5STkldbnigKg7JPu0CjorREDxwXfu48ZkXERVqZ1g2MEFwbhPz
64omZKrhN4dtpfJKmCuWYpC5+T9Hgo8c3iPrsvHpwHcUxTCluiQAozB8ZB6MwULpCMGv2Rh2LSJW
j6X4EPTFOPndM6lRC2O2/oT+IEt0fXGncZWd+uQiht6dimuMVFc1qrHpMKx7/wSuUIsyqUOBAYmI
lxFQROECpBfJVxtA3azxnK5IHdZ4xYbNPRB+zAEiaWJ79Nx7Ko75AegEOqqOJ811LrKsCzXFJZWb
NUVCh6qhhocNCLfVSnRuoWLPRWhcQkIqK6eNosqfvG0rCPmCDnahhJWxHT541vRGYnWdrqAYB7nV
qANnu9GPDZN5aHsRljv1+De2QcI5HEwIWXCM8c/vJ/8Y+TfQI/4deZgk15R0jpnbwkeW3FQfKQ9Y
HI5z+PYRB+BjrCxx/fZBNh1QQrfqSOmryJm3oYphSWasuGSS9OQDJcQPwJzbahTtOXdgRP8UdOnP
xCjC1dD3oX6wqYcL6wL5e6ze0Uqvqc+MLRD7rTCLNr5i8iyXN4Fl0+J5Ij8E8jR8MuMpbFK9vIF2
1rkb2N+rRiJSEk2DqTPKiBqP1ZU8kGyvsT243AV9qi0mlLa0hHY7LH+6pZEXDUko67IORv8+B1bx
687RH63f3Kz56rVQJNwG2owuwhspprZm7PifoHrW6HZp6NemNLOthQZeWRG6EvGHRFjqh9dNh1HE
7i6htYUD34O5tWAaiawKEKF1kP0srW2eUWhlGc8GyYF9IGLHnTf/WmKMXaVW3NPS4/ojQgErCXI1
BglaNzymoWMlVjhN6bh8pjUN5o6hIIQyjnl/fkGzy6rtckeOtTot5L9jrWufcNLZFbGDdCHlxWbk
a5txWvm3tuu3AEBhsbQWlGhhbheBS71BhKHUNcznQQzR8+zLxrMkx00vRXOHji5smXtXj3DXeBaQ
stm+l7I0dSM3hikQAAweYkvDVvSZQSil0Uju27v/VhKu1uxskNjy+Jcom2dGfnbNS+XKRzEJyejb
cVqO7FxM3sxgCyNSz1++/8JnIDj6Y29+rCS/8A/H6fyBjk7esggU+e6rnEF9YXJkbU4Fwitw0TVR
a55Nmb5pYRHfcVeQDIlBdjSKFUrvzwkIC72Y0XY8y8yOhDkdnBurF2Tt8OP/xpfwvplDoaYe0STt
85WDdGDnrcuf65cA9JiC4LNBC8HqKctk8/lQs3nUkKyQvuy0ysVJbfrbfDkicJvKe5mEUet9WSDi
x0qKoCGbnZzmHKBc1GtOzna1LjsKthaMksgAFvoNIlcScDcPI5/ae2gdq1cAD1LCS/ptZkJOoZSX
yLi3CQFQJoWOJLYrO0279oLM807rRNwtHjdnBOnr7C0GjtrG92HoZ+NaKSiNb/pMzjPrD3bN+23V
/r3BQPzAZ4w4Opjw+LGYROQw2JOJZM649ul0SRv2vfQXd7F+a/LahE9bgpZJEXFK9WswQmXBs4Ge
tTFbTBIuByXoY3tTsxIhKJC+Y1Jpo8HgrLCsr+b9AJpver157+LXq9ofmC2eH3NpXjVzit7nqu40
SdLbQNy8NK4xX1w6VGeWbtcDz17kZn8VhZvPm9CEZ9dtL/u07UVm8IKdeNM0GwYeevHvUliQyvQj
s5O0OFaOSC5clddm4j/tUh4OpagaDQ1cdQSIZBTPPti112cgiwAQowTVicdLwwMCZHbMK/0StdGB
IHSam87j1yj+rJfvbKGKgKDyN093dc3RbTwYMHfali8zCGvzmC9MDmxTkyJcKs5elH/yHowatMu0
BWSncMr/iNiYGCaAV6ECYWn6nOSLAsrededG1+eXsMoRl+NHxD10YwfqRaKEP5z78Mfoy1EJtcBZ
Wdvoa7bKcePg2s3cDRkEo4VGN458nOttVlhWc4N+NMZ76Z8olzKVSzlctUyTFwVeOVDIxP2j+kay
S5dLi/r2ZoJklQCbcM4Hnj1j2ep6UZkRWg91nzPOYMOaPIYcubZ/6HSNF5qDqhWws+W1zRGGAnNt
49ShpsPYtNkMTaGVnmP8M8NSmj46MFcVQoLLVRappR+ffiHkS2eLfP7VWUBKBXAjKEHrMKJuIJ8F
unzm7UQvvGIWv6hiHuWS5BLAhxrZ4VyXtuOmbr+ApRMqrkzLszk+wSjDJYvQjsti9GuUbUsGNUTP
P81m1iOhaSFoErvDXwc3za3fT71tpI71Hcj148AJW3jhipB5cKOTtqX7ZBs6aReZAp6MOSMs2THp
QAprcfZx4XRMCORk2wMxgfLAaJuzVAn9JMd3CHLJwM/pNxe4sdgbPQugtlexsnxfiKDv2dxISKVu
7WlrZADhNP/VqEfE1D53Kjula8i2FShpu3bJ1XwFaIBmdffVSJvxtiXmCl8DZtaEHRXwkx5ZFX5y
jmhTP1jPHql7MInru7FgdXk+3dyOohrB9xxzxeUhfh/qCDT0w5rfZRcgPQYXKs7/SreD5R0Q2pZk
K0fXenLKoh1UfXJVQ1SBZVDZK6U5qeFm/plOoU+2S2AkSu0L0uR1mPntEgAmjxPzFHS8uS+Xm7yw
BIZ3D3cvpF4vWXtGPh3E+dEVsjlJx9tdApKGeBRDKh0Bvuc9clO8X67JwrmGhPn7HszTb4wAj2QX
1X47yJ2X4XayerQBVhmjygtddtfb/sfTlBv8YJBtzhxF5EhEpnuD2k7uf1OK2WAl2+F15sDWDeug
8WaSkjOxHwaiLSOSYUyZbLHN6caIQHmF71XxDfcTC6U2Px6kXxJhT0LzZ1uwkwuHquApJLhnxWQW
wllfnsNjl8O2k+YcsMo1dXNc+8OxfDcj8unEFExU5++7g0ESLxLstxzEwA27OhnwuSWrWPLDQQEB
WCnTLssCCTD3x/O7fPS+uSlimNKTHD7gEBDo6pjvv1CxDD7JTGgOufTzTEahLZi8mlmuee+Z7Jin
Fb3xeVlOXQg0vmZpl5KYjHNMj16zzqfl//1DK636aSW6H/CDoCcvyl8EmyDoXDcziawbd9vaIQtW
dvXR0yxTtMOHGwkcaq4rl0mq7O3SSAR+eDI0yd0dxU/EwCmTY0ymcFftEzIoMNqTDCc7c78LveS/
8c+BgYLq+0esits9uzN3Q1rHLMfLwu9czA57SMj195XGiIveGyr/yxqtsaxB8H8p1JKfMnzmUPZC
GLiQsmOeRvoynQwO2wQf3UDOfj5GRJ7t8/O4cHvVqU8Cau8W49vPrZvm8pjiOjYfYEA1+KrritXY
bc0O4n92ZeN/qG/nAH10MndnHeNHsDp5bjfLLELZRIK5gdtED/NvS/OUsuoY848sq3no50ZG+ZbZ
CsCFp1TSrehW6qPcI6A7mh7URs89AmV0yWi8xViMBii3kyGZwCTue7fVw4JD8EvxDvNexLl4iXbz
1QeI8O3qkLNmRjb2K9ndO+ZUXmSGtq9ZMrWA6/l5+cjoG3/LgYgnf8K1it/IHfeMXCvGpOLWajzs
e5U2YuJrsXMZxSSodZRHxLg6zvxAV9BLCnm4GvG9FHPvE7EcjJ4Yt8xKOnFPiLBMD5Em+K4GixDB
2qOytWJDIthFarDPThhOnDYzNwyor85STwipvx2mitDKW0il1os8SigEgo9lyc2X3dvdo76WhTjT
PYjKOsLV7g+Oyy+MV1x3DQd0kg2e668xzpxwMR6Ms46qTlXEyhALOOnCHY+z95v/BllBcloC8k/H
Coqm+A1wn2k6CdJEjpcB9FnW5weZjjllxSBkR21knUbBEgpfeD7lcksvHLymWTUZ/XvBWJu0LURI
h4LTc6GYrqUTJ5dgIvryL+O0FK4tP84oCBdtnKeS7Y8guo6HV29T3WZdwTjHs6ZXEhX35BM2xMJV
YvmvbzmECJi/Z3ViF0lxQFs++D4q3sMB41lkY0/xyb2Nmpbz6X/7vvduAhAcwTdFi3aWYONgp2Gc
sH3MUMYEdSkN26L63tHFD20v2IH0K26ybfxizDO97aCfg6+5G+SiokWvQCXuCRSj2iJh4vc39QMb
kLR/3Yi5ZUle+72fMElcTWQ3tRynLA+5CdEJHe3J5PEQ5dwF5/02JvD8PA57401YiyS1fN8JEocZ
npXuOSdwzlqxeZiuo+in8j1KDEGIfL0VMdF97TOEbaSPoCYBK9kkPEzMBFRwsCwYFvyvZAAc1BGo
mne5MdTSCR5H8Osm4++kqGJUmY8nwPd6VuoLVmQ8qlfyV1pkUAcSLgOvwN6VW7at0b4MAFMFy0q3
dLfaT3qNVPbIoAx/0xvv6mBE/kRZY0tleujcTy0UJQHRoo3ifHMqfWnqIP0pQ8FyAH5yUgA+YrIc
xocqFW8swzv4R0TdUdK3C73CLmHtLy+ZRmDCjPBMmSvmyhAh8RdsyfM6ndwlZrQy8GC9izcXjLJP
jCSA7R80CKlM2rnKeYcVf04I7iHswXj+V5VfWD9E28JXcPW4VUC2K0p3kjmKVC0Cf9Khxc+xPC0m
SyZzwSExMlocQNnD+eSxKWxeu3pCVJAm/cJsaBfgScY7sgS32mPINoN9PSiaixRtCUu2AYb7NWD3
8aa7VHr1GN9HloZBLzqFE5acNWsxoh/IGqSGYLjkQU5s8e7Wca1IeCkJ5GBiuhrXxIOiHQDj8oed
IVeLFONzAkA6WbmQ8h7TiJzpruX7Ts2di/grQMscfWRXFmf0a7cUT16faz3xEAi4K8obaWuXjTd5
M3okrj/38by/0KUv8/JFH88AlR0KWJFyaOj9qBv7npnHfkYNBewcXlkohykRZk/jU3jOfjDzwQ5B
gqvGetxTb1V8pzew5qT7vKgqLY9kDX9AW8yaaU7jwj8b8yPvrSTML6s250dsbbM0KeLYeN7c/kil
HsLS6P8h3kx7aKn7D+2eqMTQa1O4HZClCUhC4FLBvMRDjSyLMuqmOBxCW2vBChsGdpgnVC2mJOf2
i1WZ1JN6vXPVy2C8P9vPmlAV8TwYxIPwc6UYncApx7P66usnNaxQG/+9orl0qHEMTbUrMWMveMPX
al0fOI2gyw29aHbFLVLibxd1IRBWrMmRCQfCNx9Ic8Y3G6j79ukGeVBXrO8E1LH+yoJ2EabFbFB7
PkybZBhqUeXpx6CfL158jZ6uwBI3cOkP+33cPwBL8ie4GtJkvezz63aB/hcYvc41WowW7c7q+Yt7
AsmQqMJgx7PNwDVxo4Iah+90TTeB20h07uSwz8QEdMtfCX3ZX7J0lGAIS9mmBnz6oHvXRTqpnyt3
bJYlAwuorjuqH6tL2TiZjiGOI24cn4PUhJEDKuLTarUTpIYvdNWfy1GlMblKD5KUmcVfImyAXkSQ
DHyR1ezmHGmVAJr9WAzny1LBdXNHh1aNQ9BQzp8IcVZQR7QcCTcHUvd7z2WldB6EPgmW+B+wIDF5
SpdaG/UHppltT0Tq9FjDuUmjC94Th2dbm+ntKiZVeOvsNWo+tGYvQZJY4PNaX6vsWA0mQvj7crAN
LTzNB5rhoT6hQqy9tYDXe4Q4a5rRKkJWXhMmduiqUniC723u7GPnthSio1ur3GbZrk12FTsTpIgE
UsDz4Ht2DiGIK2OYsy5GtWMJ7RHQBXAvsaRlDcBi2b4/jPl6PNBQIyTvpKdcbkurVYkgnQlqfEMZ
TAQU9fohhPZZ5MAMznUN3rPHO67C4QC9+8pfYo9e0ERSDXGH5S3HAienRhZMK/QrgCM2RppzHuv2
xihaLiizkXimakd+BGcEpPxP/QPT2VZZDaZtYMqtuEI5n0wAtbf3HoxgvJwgF2FoWZwgqmjLsjMh
48TcBJFYKsnM/6TDdS1Xfrnq00DS2e/d1JS2bzvFI42PdGwhOgUXyKF7h1ZQ3hATfVBAhZJCSApx
aY5ECEVZU4N1IXQhLzji6B+/MRAYlLQt3vgjpaKNeW6fwsKBOWWUQerzpviyzmDXTx3r9b+ss8Eu
fu1cc9Wce/gbSN5XdvyJqS9gQeHXtjCFQAOxpTWyxUGet/nGl3I5Lk1Cyhnmgv1nbwvLfgf0pBND
C6S8mFivqDO7CHbxiBWWS9R3mz194N4FGfcST+K3buL15MNfbAGa4UPI7TNKgCKF1E2fsG8pPUIs
ylD7kRwhpaFPaBhPbYXrjV6TYEziGKi/WKiqU2skli+pnPPaxlrCagRovYvOjkHNsy63HWtPKEXl
IS6LcDYTFqOzZMNTda+YQ7jTk2IlcfGWt5Em2rNtprBMF2+8PrFGN7OfHzDfa+6kT3pY7Qaq/Anv
B0YVag6ZPLoFrQUpzS9CCnkvYZuXMFL/p4gwfhFrNn4Z6q75PRTlpoNt5q+bq5McArnBPdwKcbMB
DYX7/zYsw1nnBI1yT2bOX1NADrAE0FPd0BaNSGQBzXRwHXExSvEgs5sNJzXPPA+c5hbVIEGsdCaz
arxuZ9wMYKBcMewgLTPTyRFiTJnG62HdTJF8Uv0WGZfGTOa9oEfMZfE5Di70fR+WTQsPGsf5ZSTC
IHX6yMIYHM174GFGV384ixa9KoYtqS407DEg/IwYI5zXQT9T9zrmJ6eieRITB3nyUEAELsD6pMqK
3muREEa3pl1Q+DxsJE/0A1qkXUXisS+dOewQZkHmDopy+3kYplzNlfLhR9B2PJyvT/jvjpNo84qb
ZCc0DQKViq1M+7S4RE5WoCUJsStySVeVVZxwoJp49OKvHvVqkCnBg99F/nfy9J7Uu3JEnNZ/lgCP
TwvpbePJSMB1a5b1Vc4O2DBudrxfsONGqWycPKMZTyqfttV3bdf8+OZaIeRgs6qy4T0gU2YLCdC9
9yr9fgLEc+vRLbNi8t9Qf/D4FpVGRRTrJ697oxF5zTycNf8Pxz6iZZpbA1Ao1Q5LGLLvRRtSQ9/b
ZMH/YsZf9nCNwnjXBtpnvy4zJuAMaz9u60B9MNWRxDsrzVbMeewLWfR0xoOVDFjU8UlyGj7CXaq4
6v6UClujOSNSJ3J8o3CRHwwmoeWg/Fh9jlYn2K+M5KhDtvWa58mkhEr22oV8lGZVurMvx7m4pPi2
UFABivicTvoBuw9raXXxSSJ77rbdX8nO5Zx25MsDQEeQN1QdrnL2+ATh81oxfDCSMUqkLzaihbhP
6eZV6pbGqPT+cJ7zmrm4HMcu4MhVNcaNJBZKqYWMgkQVI/fP+qGBMfTzop1r2E+onfRFPodWysP9
Pa2tTKOx43eFfLptLy7dk/conevZNFEmUGh9UM68h8OflY1aj6VOPkqDtf5NhpV4YGVY8CqBsuFm
MOMyRmmALuKCYJfhHLLAO5XY4IBaKI+UySGO3cDxN8h1CLrtJfcqr+STFTgM9RNCqdaf9DAeCnSV
eGWl5gLZxWRkFNiEwyWtCyfUpWtt42eYjqewRSMg87d+I31lzTYussGyFppdN6jUn4CFm6Wiu4Zz
B9vbPUsj+BSBsij42dRMqngc5vQh14zscv+zRg77HCv2/rGI5FNHRztF8M61DiXq0QyfUy3N7cyV
DuNiKz1xfbLHUp2cAmo0Mcbu8KADLD5Dmhsz0lyUqgtVTxWCMe2iWKQeatf68tPFSShCYwYKij9f
iAHImqBaXLfk2P/M4nSF4Ef+f6dJ4XW0yD/x/qSMAU1ILYGZbQYjphWmDJzQA/o/int1LX72Yq7f
mG4eBRtaHQADeElIJaTUKIwTArN8e5TsWjXBubJhNgV2nSh+ZxljIFACT1dKq7WxDWrS4BWWMQgz
4ACI3I6RAGz04i0f2N1VkJPy+qfITv/BBSa3XQ5v/MRnefjIr+VvVwfW6xwdxtl6U6yXXIXdpGsZ
YkVAPZZbBN4h+dZRnOAI+b66e3eAkL1Q/ZWTSbDrta6RGaVX/6O8ZT7CB+XEhxYe7jikchPR4tL6
kBsNstw+dM8lLXv2+XSoHjDp2Ozl+Alz1qYnA2jfAkbAq5stB0acLPMxQF60f0b6Jb2DFivwVZjZ
92TCqOXIdAPrVR7kGoD7KFZzQfn0L1uZ7H9bXgY2VuGVrOks/VKsz4iahfikVbuomyivCw2qfvBP
lETqucDEkrzDmAItB9VnvDbpABj9AbUZtQpoV/nvPXZVwcbql5VBdbnUJwSKVbIu2bN1960Tv488
LkjMLvmynDk9Dyum/5HQg+C/S20ny+uEm4RuVVhin18pByAU8o7r5h6cbTG89588/edpdjoEIOfp
iFMwR42w3AqSyzFZooTUXw/J5Rnq+YSfiHH3JXfqqnX7LzhVwDHgs/TgHXKGGYFKO4emUulT5wai
UhDEKdbRxwycbMxxCycz8iRZ8MDR3hqn96OFEFW+gl8k6IGr35VLHtCtTUKDoiHyWL8ihAqe044C
Er6v2HLYH6mf3tcWCi8E3aaJzcCuCmRLnud0xTUE1+inOU6z4UeJj5ChOuApGCod27cW52y6Louc
Rs38B0kKOUy7X00arUYlDahxo74fBJxuNSZ8EQxRDzF2zReYHiPTD6L1HkKVswaNwT3TLSnSwcfZ
zOILTiYyqXVFbMHyPWJzkZdwE9wdvhC0SDL/Yy+NzXWNOqToeAGEkLDUxP1vzLxqw3Ugb9Loh+Zo
gTNOJVCuUERThh+anZBmRCrrTUplAREa6DcrD9qIQ5WSnxqu+RVjJZ9j0WaTmLVnEBXuSFi4sQVU
6DEfROcf86yQh4p8OW/cBxEv6e9+AVlVktqHRoylWd3LKSo/PAlQsfVU7Yl7qtDVl2DQ4bpZ9IAL
R1Gv/Fdpi9GDjoGdMuhRpdpdVsYUFZ9bkInQD9EE1NWF4wXrO+GkFfnQOIpVTuS/TUT7anwxYNla
7uRcIp4xKNZLTZlOhM8uQFxtfHcgW8a7FLTbjU+9cuxGbkHpZKiSlZhbp5B4md4h+QsVyoTHPkNT
Rv66I5v7ZXotz9nTrvRcjPT5Zz7lKOkRcmZyovJ8Efyas2ONpZsOZ9/0AHSwdzv+gtUF9X90cIIb
rnOHzQx5j7l5XfTHqKiPjaiUXWMJvSvYLEkInyHc8qm1B5O79mvhVU6Iq6pvgC3ng+KjCLE2rciE
6+PjJkvkFYaAnCJZ/500SDT3t3ZHTGnGGMq2CO2bHXJ6Eq8KKYnoUnvKtZbpE5423pLkqvD0nrK/
mPFhF+1xr4hv6MWcslthLadpY0CwgkFsSOX8rmJKSvpGMPSCKVIDhW0BoAiG/Klil3P8aG3wIOH6
l1/MqOwexBVpHpaTSXEzoI4eVIkFHprRM+1P3G06jDnabgtRWOjdxKoWyDFPt3544PuwX8p2Z9SN
z+6wA6eULNyIswNtw6aKCnMfVn+Q1y0g9/GKHUyIlS0+sIGI7Mg/9oafuQcpeeRgaDHwc+j2PAT/
gxG+bT03Hkge+2j96U8JGcgdWuRjl4JO6G3Wkxs8PZkQ84oEV9+jOMl8TZpuRjgHcedrNnmsqBRm
2DI7c6rIj2S0D7uAW47KwXq3VNcwhZEGsZuFNNU/D5IwOCWLLaQaIcNZQ/InIdGFgTCTu0o1RWE9
CVaAn69t5AXSyHwd56p9ZwuKGYXCGxy3XlwddZFbH53dv854LDXYoP/WI/BxVnXiomXEU3FDVcat
Cj36ZJJVWW33nepoaryIY93FFouCd4+T3mJJhRcHcXQ8AtAMMPaZQsalqXf1WHBaI4MS0XaFHU+d
aa3zk/taSjOO0cQy0X7o1DOx+wZSNZKt1mFtc0RvD9pjg4ckuuZOGYhHU1uf26Y4aF+16HwCV70m
TtKKuhxyDO7mKIFd8VXy7xsADaWn60JZOmrswF9AprMqSrHT5SURzQi8ER1nTMVTjTTFUXzlGLhh
s4v0IoYDJA40TH2nkO7dFhFh4O64t4hNwfktnjZ/etrg9embPrCTbcHpEoShlb/OLbalCY0YU86q
Dt2V9RrSdMpi7LiUCTjA4r6mUXtEpvFu5UYcSIOdrNTuX2YQFuLhpZQYMoeWFmQOMX89u4ekHo1U
kfVJUojY2F+E8OGHTUBU4E2edPDTw2z55uOBfPPpw+yvjBXMKAJcJI+3PLMPEBwDem/veJom3lSH
pjc9EEqTAvd8r+mcAeZzIOLbwoa9/u7MrYyJkOz+3gitd1wMl6WhJ3gQBhGYYshhPYKTL5EhLSPU
Y38GxlvZ733j81FvfJEjkzGFSOiUqDAjOIZCY5oHJS6I/qnDABnDvhYTX7KVM6AU0GpcUFSX4sGM
V4nwaYpFOSvYIpmhtfTA71Unc7qnJphpoOq4elFTPnCgqYGcC1XsmTzbm4PXqooRBskXQnduFr+D
CzFXpGgQi07uY5EBl86wpLBX6EpsP7GDk+te56Mj9qb/5CanCX85AnTOxcRwRWv+t++ZYFku1Pw5
X/A149FK2H/8RApg8HQ1tufOHRBFLE4/hRSkuK7KF+eoCk5+FBqnA64MV2J1iVhmKiHYLDIEkX8X
U6N0yb3oJbMW1yZZZzqdO/THMjGpLJnu3kYgD/kIyHE3wcHtDKU8XnCc+pzLSdohV4e4bxKjFYX0
NGgamCmJ+LVIbMCq2iFsL7Ai8ZB+Uh94kgtVBgtlcuTkEfzV7/d2hV7E9yAZeFEkHEgwGyaYblFj
BGzNJLTYPdIXni7EHbaONkmg2LRRzktsaoLl3HgISeQV5JEvdKjhzdoKnbs1KfyI4w0YZNTdxCP7
gg3nlfPaUWc2wc/6lT5Z4RuVtgGyJU8OtzGXoWgnfaRvRZJk2mciT7SBmuf5iUrsq1NHBXePvwUH
rfAw6wPQ86L1P6T/y3ndVXfIRrDEwnf08GJG02B1Eoi8SEii2Tb4lMiHT8PLGQkHDSFSubpFUctc
1P5Hs2bnfcYZJuLURQmU1Efxi7HDhf5L+M5cWMZ94YqevHrEnowMrNYobElljWTOMy9RCk0/kAFu
PnQlAjj7aNyYPuUW42AyUBy8x0wLXaoGGHH9WthA/o5tcjruujCWn2ksykeID3v8bcvBCTKFtvzM
o6NzjhX37X5RSqsDeEWSzoB+dJUYWxYhInmZ4hDxPqal+n23MRWjHyweYAY+7jvn26vkF/0wqjdN
JRhRrqtsyH1QRyRg3zQ0JW3MmwGJeZvCmp10Bi30MWhQXapZDRlKS2+lkk1O1AsetqsDcUjWJ817
YrlzNewHpGSeqrdPXjIlunF47a+JcqW8TYqpTBNpQ/O7LuPr+LDKOpJLC/p1LaaYsoYTnJi+HQQz
1orC8Y0VsD+Ziygp4S1Fj9SIhm04sCjEzKOT+0lma45Nm9IUiLa5/9YpCRaVO1oNwsCX58VOxe+X
iokINa1VdJbInqhA87WtB9cbZl0BnfWsNSrKqimj5KviLCUTipS3ERl2iDdhA3PhJ0wrjvUA1fER
JgNJPUGyGPJkmYKwULCvTCjvIL1ZGmBYxJQBK9pWkv57W0qDLx2NUv2MyBkIwQzj8UxbLVRm4PM6
zHOL53W8TXU0sdd6fGvFgWdpAHTCXrovrl2WMIEAEVF/IUijUVzw/wjjOOSeTlaeDsch+jrdch5l
cYT3ml18G6sRVy4AYx0+a0p0UDg+aJ3ugrYNE5GfpJ7wB/3zXxh8jTkavjwYNp+uaRR9heL9ShX/
kG37GLWbxt3mRqWNtHKocxv5lRf6jAviFnmcvTlCgNfVnRb7tOy9japRifB1ezb8H9ltdlUqNTBC
JBIW3kis02wp/9xzJbPwan3jbP0iZQ4D8HdKDaZ32sY/Yq1VxM4DVmoynfFxTgTjo6zxj7GGOT3Y
LUj9TNk4j9kVR46ysdEd+RbR18J5whT94wxHfI8EoNdnSQkwehrjM1DrfGk5ha5Gk2Dr73Ay01l/
SBCD/U7ID8ifGJ8ZIdj+3+nG2wL+dSRI/Mgy0g43EAQsuZupNqQ93LwguYvvRBNgMMs0tRR9n5dp
OkH8ZFDHxW7t8rolMmBCMD9if9vtcKsc90PRd4sZ1BOkDzNIO2wfNj5aE/ehuGzwq5p47LAw9lrf
zqx1ZlFFnIbaTFSJJiprNV7g6RskFwYOjykfPjjUSGe11Ic3Zx1P5N6Awrs1VEsWlVf2qLY/+Uh/
xQVFPSGsbsv0K8pksCXZYi0zHteIayi3VIzXITLH7VQpzppztGd3ppleRM+D/9ppKrbCN/t+37Bu
Anv6ZJsmMR5/PUcg3soqauFuv1R3TNM1znW84e/9EsiSRAOQ7ARv1+Z89vy7hWaIBC7co1BvORSX
Fs+n+a/kv+ojZ1WbIWljJ0cypVGDSbZduZv/HjW98JaMh5zr/GqvolagLQtzIVw3LSWOHKawhIDg
30iYR8JNH7PDs8Jae5YSzxAzzhbBxEz2oN0qRd6NQyx6BIv3DIu1H0p8zIEvJZBZNol3F3u8jgHa
+Jp09lxPTBt3kGwPJ5x+B3EMFs8P3GVLG/a3EhCe5dUdinCmxv+vBn3HAf4376kTVWO7NzY/TbHw
5p4mNFY4Jv8bWNQynzp2pzugffJbbVg6vGzZcLzZTQc0jf5KYNYD0qnBgMsJCBM9alHk1sCWYjjB
Cu0coxKhMB4e5fSXoZ/xJeJbs+L6qqXGxxYlkBeFsn0b1SR1t4EWkg0T/DIDnIrKa5TJCxL5PNts
tbYZ7kPaq7rOfJsCdLYw5E0np7ZBzZkL8Ci0w+zkh7VHmYEgNPVz1l7tx/+oKcPPA1ZoKf+kWMuq
RNlhqI5gUSjbaVkjbRIb3RI2mdsrMOTuEO2G80N+rMyJtqunrsPiYzqdmHQsbE/tV5AjZBEJseNl
RDrs5TsFlLzTnb0AU5vqcZyh53uhabmaF7HVQY9ey8DBZtV+s6+MUFOwVfWT3DqO94zdRJBlZ0ja
7JBTwwRK+cG+7GYMgVHe9rpxIqQZY2b0hJBLVVmhW9PDWiPj4zmmLR8evkY3/d3Xl0wkl9HdKZQu
I8bOM5zuhXQHPyBqkjZJ8HjGJR55LegSbphS6pR/aSmm3IB/nUf+IQW0cxAlWeOtrCsvwgNUsTgr
EngeVgjVVcMIr7CqQhFFGYFEimwkDLH+dsxAwQgpy3WsAFLVHis4VDiDt2xoGAR31TaIZ8ORP7aH
/blxnggp2uqFHI1Jb2QWSs1v0AzQ35wptXqvjC5CuDJB9qfd9hPUY55ESF4ogwFgZj2RzlH6zswe
R1kOrnDnxSMfjXWtezAB57gfCVbttnPlH4LTE8N8zkgNlpQ2ShQHvaPYyrDNmjF+zkuAqAPTEWPg
D7SeNiJX4p+NqmEnK8QE0DyxNJtWNSoN3rwoefh2YX12R5Mpj9ZjrFJaCx2cTPW1ER6LqQ+fwSXk
TQmyL7xGtDD+LrJSEooKvh4A8wPJHQMrKNTq7lSGEefU6rfr1DbuUZzCgW7rY/tqyfEALu3hPMkz
T9y3pGS3a8KhHNyCdepMZ0s8O9oIKHapiGMyLPz8hbZZPY2HtrUl2dfZV9TUYNJ+nhlhfFs3yQsI
fjidJYAUl5YpqlLDdcjWyQO/4li75Tz9eIOyN00BsbABR2KPnpAS8UQEP1FSea+mVONQbM7s1EgY
vzMc46i58AQVRDKOPf93+OuNa7V5U8l+LqbDm6nuCmNH6YkBWIeo3ilCIFc7sOmdlYCS/PjAA2V0
d+1A3NTw3vARTsDvfpH8IrImquWGmi6NN0ooYqEPRXQod6GCwJ2S4LAZ8ZsZDQU19kNa4M7U/hXo
ophS3ldj9AdXk7DdVcJ805nal+cc2gDFczM2667kanN9fHp2x7Ka0HgHDaf75DhgwDYobQ1f+2FK
PoZxYhfEHYwo+66yaYAJkUTikkh644hHT/jBTox2qxG0cg9KeRC2LQe2BZ12WlNaNncMkS/7InrT
5NgRzqbUnYMzh/oQHD/otEHFQ1OTFGvjWYUWryWYYca2ScRYt+yQ/llLUR65q6y6Eq28gJeSBYM0
1+0Fp24e1c0iJph1IJ2dSsIVgxpz1jy5L/dPwYPr3kjZsMRLGfrfEpD/aNdghYNB8z6slv+ZAxB8
0U6DhVJwYw4u2VTxYp/uqebQRuaRgT8u6h6S6PpJl0r1OD8TNSlp9YM8g+siIp/JC7X9gONP461q
VHu73DOe4tqzLn0dkg5AogYWXjGYJsurTof3KApsmtgFUtf6/fjaEXqJcMY/3OooJbuaAv4jhuft
p7tF/kkUXe+jKFciGN7OmJFFldavmPBONLNM6v/7qwF/0s8j7Fx/2W3uTA4T+ZsxW4odZ56WdDvr
rBSY/FL4Dt/ar+/olP+KdGDwd3GoxP+o5e3BMNsOFLXBjmZIMmtqn7RPO/Gz6OvK3kFgZpdz6ek+
eZNVBnnRCmldpweYR2oM2HeKCfU9U/SaAROxyzLbcO0tkb/HLRdwyphG86Nvx8pHbhOlue3oD3rw
uOZ+nfcOlYwary/PiXze+pI4MJKTSk6nkv2Qcm73ypDUTsO8VjVDsSFFBw4bMZGeEMHynuTWOcmL
i5dOF4VmXwFFZ8r+lfKRujtIiYxmpxAJuV63Y8ykIvRMP9nCMGXYzt1rKno1qEBng2lZGJQpIHxF
5vab/SgJ3V7PP60RsOwruAiGAEgSuD0M8EKtcgddzbtQDvQs80+eZrftAYTeiKEDISSye7lug/53
AAy5nN+0zJW9/bk+bJ0T45bzIUJoZmVYgElV7uVzoA7+PulrQ6iSEf2SlIIyxLj0faQfWEEUOpDd
4eaFGccj74y+07kH4/iUntTG7sJAll9hoz/K/hcctjSGAXG9V/XMZrV2XRAWXraBDfte9ikYj+lx
9wTzh02zwc28I2YgZBJa55Z/0xrbOVi6v8HY/O3ZkCNJCMoFuk6TIJ7J4ALqO8YuPNpYWGOrGVIc
72nvE4XYZs9XStKTUheB04ZzbB6mamq/rXcAHoeTaKwd+/Ys75GKffxYb0BUeRJ2X9+bR0VlgE1C
Micv/FY46v5fgTYuHeSuzG0jiN+/bWwtT90r/K3s1b/8biQy+PJdTeMmm13lxPq5UBL4OlrYW4uw
rt14s3FhaV9gpYY0E+UFnnG5RSZ+CAWnlGD3ryW4C4JX8pXmKQBMVSPIDzUXmHImX09aPlJj4vbO
DIG7dzg2/2zK64FkKMvz8zlY0/nBXEswQTY6r6zClAwJw/3272mYDrPKVmi91uCSLfJz612zoTgV
9j8qsRRmwtwg1WS20stWHzSoH/dhpd85NkbvzePNSegPwQePsboK8oBFjsZm+4KPXqmEH0bFQUn4
mPWemnF6pvk57w2KlJqvzfZ6yIGDlD/TG1RDEv0Am8FutpkQYmwesf7S+0H8bSmAUmOLy57oEQHN
KD8MfwWL7d472JcHwFsScrg6sE/TESf9qYnRSKylCqIEMzM+BYvxpYmQZZtDWeGKW4eApOdUCxs3
i46yC23kXQaipO/gRNo0hoDmDUskoU3sP6Ep6UWATOlQPOO1LnRdiDnUNameRXk80nCNxMG79XjR
I8qEsBQ4AGHFLSPS099eyzlxCWfa/4Az1+h8MLofmhFhDXNEKXkw3ChBpbNqFiEW6iNqiaGwEGQ9
OLi5GY2BxrBHaDOmUQd2ZJRx+6FYVJUoBn+fgc0bnFiX0AASUjijAQLt1SiktJDE4FVT/JuvGCyY
rfE4AmY9LammHlLGBofzjN66bvKBMeY6x3pYTtZMM9LXmuU+Uy+hvieCqt7OZOhNYgvBEGi2sX7S
FKHWIlK2A4uL9GtJurF3QqQOCG1lE71Of1RHQY1jK+MqxTzprTly5vohRcFlfga8jw5C5UKC8+o2
dx1VvNxllZxki+eQfNy8JykOQDRqLq6R3NQUhDXXqGg7k1JaFpweEo7JHWbYhsRUnwGF/BhEWb/y
59SkiiqRSytvjGcoJSyR7k7wENAAmfQFrDjmlAz+U1UwQOl2OuWT6S1YC1xyaVuh6CN3vKZxCYc+
8cGGd7JXSy92P+yHiJH5uyaBxrQ+ezBadCHRb0G6RhWeKTp/53M0DRAbY1jbxw9D3VuwLw1MMNT/
g5Y8WMWhc+TUVClKBGy7IcJqqq4QydzUZT0PKFUYrQkcb1GlRPKLzk4EdcpE+x2RdCyz4DjZbl6w
Ce63cWEvA+kFF92zQsXHRuFQ+2ySx7ScT6me/JRqz86yyG2MeRCwuBle6Z90EaNVErXZP3defqCz
D7XQgv9FnFMtojGRGZQ1sh3BbWNBJr7F3DE9Ax4fBpuDugjQC8OC5wS6JCcD2np62pkqQDsn5O06
bpZEWc3C9TbJHp/piCEzBGjYs4eKQEgIKnNUWs3edQAa0wJItFkZzwhP4fVjQ9VewWdtJCStuyiS
v2VLwG6pa46xLH1lLuCyMXPbTC3n6eWP0chTnT5frJbpoH5iwqhYFnfctcO3mPUOSXUIzby7tyw3
OmSlnpkhrXSDI/1AhE19BnHHZQrS8P6qO1wqgomakStjd7hgu1ebn7OZHTqPEwPbvCkzwvuf+5S3
vWdWwhN+wEOPom3tzSJ/NtAO7/RZcnkKvT1TtVizKcZdmavMTe3bdAIhkAMIZc9+u2KO3fuP8MnQ
O1FT7+IvsRJZfH82W18LSAHsyR4RiRGND7XcIuZC2A/+Qg4YRTAOAX+qS9iE4is8igrwYcjhgxh5
BrTmGAG6Eci0kGpG3RJexus1y9iDCEIbuPhibIIKnciGQNJlTi2dJ+ndRdYrDIE884OjKz5x/29s
mM0V3CXundncR/7Zyhg7TaUwu9ivkRu9hWcZNJBEb0Njqx/sqfc39fLzkeMIeXW3rMoaKrxCrvle
4lzOwuJVpF4AG6x/3l6hgymIEhl9EdUHRvoDlMH9fZkjAjyTXf3VQbhgkqxgieF+dWSo03dFcZ4M
9y4sKF7+74Wp1QXx7sSHbVzVNSwRbK6x8xGqVYHrV4oeb9jLz6ZuMJaLhFVnmo2cZXmc9Ajy9vIX
XIeOo0BdfYKWJjj4WckAp2nRER2ppBW7OLJTi2gzX+sQzDabotKI1e4+32d9haXKVGim+61lqPpy
AI8FEUpfAv/P2hsjJz4Ood4sbG1lLA1VPsqqKQ9KrOdXCR7onlmgHSNKwhpZVSxLCkv9IT/70baA
z9RjnJRlXq7o0VR59rELBlVi/MahrXeJLwrJ4W0Qyzq8zjx/eG+S0JqLwbAS/kZdZkiZQtl9RPze
yCDLrIgMfguMMQpzKIXJ0sPOdbQPY7/u+sGwkBxm/E+2/CGOOluDknyzYNHzFVDdDlXcnJ0ORgJJ
mw6bAPi+heJf8pf6c1TK/w4uVX5YT/vL4HvBGEfgUFtYiqcQlX5GSqEwHfIawCOqTlvIBJCsVdit
hz4VWcg5EA7hmcFZY/cfz1msvm+Lqxa/67zC26JhqPWkZs/9xRTHKixR9ocXQJNRYGw0r0+UmqFD
kXVBLhZ7jdQemRUG1Rc5GIo3teHahD/F+Df8YWlBOPL99nuOtejtUS3h09ow45N1hh0lY8/CurpL
XK50Py4Vf75jB0OmUWTiENFgN1DaG3wS5Z1Fk4A2OmQ+kaqSUMZZL9B5bi71FSVblZAqi+HJJVf1
DJ1naY6NcyhLSvgu6xQb5YA7TaLhxlgJqT9KYA9sXnPFXsV43/8gHAEe7ApJ0PB7zguqaX5xr77b
3XdAn+B7dC7rs+j7SDQOEV3PG7gkl2TywqWOksvqGN+13phwfM/fnEUtOOPQsW45yADuYolqmWM2
aK5ZWS3Yhspp0OrZEgUIlSAYccYnBT9FAswfBE8zHcuk0BcbBRRH7oxfiXUqBjwmgIfQ0fTsZM2f
+SVUE/XfJoQ81q27/6/tJdd+4DWZqX8F2mS8zlXBjcZY3F8yCe+Pp+mPnWcQcW6/NlTGcMKDecb9
17nsHpDbj1XWtRDPihPtKe57bflJ04lOpTTNh2l9UGlVrz8kxLxafz5hutGuidcVCkPmnbxdkdoU
vR6l++agu5N0jhtqx4a38i9Ba2EMwEehMklYZEM/x6qjze83lQ3zAwYSjPD5X+lrn8fqFvmjKGOt
Pdbn77aLDJHmqJOzpJfBoj/MfadO+LcJcod0aZIGtuMMr1/Q9Sh33D2/jQWlYmzq+tJO+meZN4uY
k+kVgR3zAlHRSDpQfTiWbFViTjQ2se6f0yGA8gvTq1brB9g7iAL8pqfMNElXBYorrRo/EVAs5RSd
ZkMuIilIJ0LouR1OEi0ys/t8MYxpPlEe84e6rexTGNBmVY3IUmlD6wjJUtvwncOEEo1gBMcRBn9o
Dia08WJn3EjezdGj/KGHhEM1aujTe4nmdPukcJMp97qWYuV+fsZ3jIFRMPawaD2EMGMkSQXXnOJ3
iivdzOPE7+n3DEqCtwEa/WOEroeAiOLcV5K/zpcSPViEGx/fa8LmbO0jpvW/EoahD53OVaA6fpIc
KhT9S+ln4VrCkgLQ9xWmIfHbodPSlW0q1ASftPWn4dwZBTVkYdfsIh4vDREnWMLfudDEeOcm0M9v
1EIW5g2fwFQDa9uT7odCb7xz7kn4X5F/XFjwT436RC9sg3w8RiM0tRTI2zoaMEN1Ww/BQeMAYjJf
D7gBTXtZ3LXDCUqh+ZHUJCYmV43+oR0FBV4Eg4QQkrwxY4q9FQf/X3kEo4nf566u2+b3DAsTtPSG
euajtLfcJuw2JbjL2SO2SZA+gUxBZTh784gafFzb7hAowBiYwli0+b6Tb4mk4NTOFmdfeIk0AlML
yXcnFoS0zTbJ7XP5I0yjIRzSMncYu41MbJ4C1840QmS7Iva+nMCsuQIksPRWPHC/r6ZD4uGBIFBQ
UbNY2n8t2nrVTGbY1waXBwaVKyOyGINxUUG/xDnrvH/3fGyskH+WInEkxs7dUNC3CMVeqzqpSNbd
q8MFjL++qAn91VF3rSxrOYEKfwp1YOnhEIKE8TggaInodyALr1iXzA7aV7pkKBPVWie2yDJxs4Ex
VUYeIzSnTqVZWWV667lnR9lhFuvHFK+h9zYWUZW3FBl9PReCuxC8bjiLDhMS3RLHli1K8PM0zTUk
B1yJSgnEC5r/Og1We+klKcMJG7Cy+kBW48KprhkimTF01zOI5TqZSAjxdGtizyslVqwWO/g2e0gh
sIW7aAX07LpE1sPk2p6F/Pw5wMTRRGN3vSNwsQf26+kBTFRvCWCe6ALZIpIr2OJIyjgLEW+NWqSj
Uocf3ORXxhNB/cNVxFrueKg08FcUDbuIrBhXaWLr2B3N3o4VeqHKkUwEKIQcHLJcL+eNEhkMQw4+
Bot1xT9xyQpb0Yvq2DRq6iDrJYuL5IB+j7Vhr4eJuJtRp435XbRkxJTTmdeC8B+bmTgBBK1ZnWGw
Zl3MmUwnXy7m1e9nwFnx7NSnmk/K8SC8CUwg0Ll4sOgk1dLnrx38/I8ciKoc8QTgUPULMglVvG75
5yA/z8WMlvieZQI6DGhy4I3C6Jr+iC0VSZHgkOdMpSmR/EM1zvHEFjPDSPWjwYIpPhlMQLIYdX5k
uYUMJJHw/JMme3HMCvsrOkY78sgqO4XQ/MlYB9rggeXPQ5Xlo92lsjL2h1EVqtxkplXU1bStvz/A
Nk095AZGRTysdRc63VjLyhAeeg0XDgPPfaF0pn3d5uovpsAnlTcXTu8WNXA2tZWnD0SiZtY5Eoaa
TV222d2mgQmyRPElO1FLLBDpr/d8ODg9Qm/ISi5BzhyjU8zRt5Mg1EtLTHlC4Fxyki/o46qAp9gx
51UoPFuq+aC8UZuMUv/3WCkNUZaotXgMb5ITBMy2VG3X4t/3nbL6Ygnsme8CkcOYeaVMdQEirHSJ
wof2JFdolqoTIN+bAQgvUUcgdD81JEBfrj+RqhGuL8s/TpYkMbC7ksr43xt5YVZw4DxhMPhkVdPO
J3iuJrObPviqY9lK4iqgmVb9AxjgGrbA7Tjzpm6xDhzl+pZZd8hUqURKg8LhPGAgobT3OJFYIXwn
dc3mVV9WGawn0vg8jcWOF2S2txu9NlDUYcRSdXgnA8MDLnly2RFTOC/YOnyrIFKE57HQBw68QVh9
IHoLdrmb6K2/S8+/BJjHsujQMBPCZeUzktpoGdcWM8icschPEdNud2DHKCeO1R8S/OH2MqedStvk
BWWY1+34j+Qn5yVtOhGweyTxhJgRV+L3g9My+4j+J83Lfzex67vHDzl5nWbM/X5LWbq7CY+g/xYY
qPfrzb/eIwMNQ0G5iENWbQBrAfCNjKZIxX3YSAv04u2K50bjPCuzTQCeDnjRms/xG/7DW9Fnz1z6
+EJj8PL+VcZNc0lISqymFi6PCchofDZi7LgCVR3sqbTynKOdA4wtia8kP6yjMESyr2n1Vxw9SlaD
bZLGZ9CZscqc74okEqOV0Qe8JUZd6VyF+PLYUJiYERz9LOvDGl+JWXoruKa3iyZijcO2YQvrVb/g
6ayIw9QwVTCSnG44F6NAEY1oqgNeLGAZQoUE0UJhlPuNK1Weymvx/yix5It+RyOyAoc6CwhPtzmT
D8ay04zjQ42puMtPi/NWWVzKdINaHeczY7b25oCoZyl8ShXRPBPlFwYDvr+iHAGrB3OOQXQAyvH3
7ANHfV5QicIskDbB1ZGWKVzexSzpdc44hx4uAGAgS/Eg8PSahfWRZQ48m9bAitHEsSr61ndhVhT+
Ntslvq1UORLLIbigASXE8JcwVJUYo3zmGRUbpfEcMYuzFnDhndPxfk+y65I+iHYHMuZ2mvBvMEU4
eags1jLyK8ug9W145V09zD+zUEX5fOBem1jeZOiEEx0uJUOK+KU4xI1E5ed3DhnWGgTwnY5e2FAH
zr1Sv73uBbfMRD+qGOoz7R0gAZUrr/jnIzAlQXJMQiPgVbqQSuVYplVwrSwYu6nLV4zASCJWZ3J3
jn6kulLEqFxZRZxTQrOp3D7KOgU7SClfaFjtopKBAXx2KixQ/GRbKF+1rAqfyGra0Yf00oG76LTo
s7hTl3pY0Iy4CNa5Ps95IoTU/TM/zLJXmbeh830Z33+G+1PoBIvSAs81TlwuxtnluEcb76ajxkpP
jybev55Eo0JfZhBYodXagDZcl+Acdi7SUaUXJb1++Jk11JAT6B03Ojj5S0lYZRbK9DZ3sbgrARsN
aS6aKq8Xt/LAhJn9TAReo8Fpb1vw0ZMlsCO1nOC6vV+iytWl2kpDF9WRIRmMIGiQM+IVgRIG0jOl
yZ/G9XpLkTB6WK4znogUfhkO1gKVO7kt8fLLLsiNNDu1tnlk0UWQQHR3Hi6IsOacZ92dnUf/yAAH
cMpB8gGCqnzedSfBGS40Wwob0drNpdYxf2reyGI33NtPeJ8Gae3jOy0HDzZXPH6KYCeVhKps9+Gw
kXDqRX80i9n3sLoO7Mf+ej5I4HxYu2FIMkyPkCCkcqL1Ck6yOD58vfbS+3j3gyR9LwTpY+VNeEY4
e50kH91FxLv3uQW/l35qyY8ux0PpS/eeXqT3c1ejnIj3C6kc+fn1P3RckdmUxL8VyISNtMmxhB3a
INzfNoHEC7DjL2hy3M//FTanPuvvcLEThQgKDkCgEVcRPdRAJHhQFG95PgN6Jtk67kycCqJ4hMcf
Gt9/XCVq++q7QW9lui6Grt2nFFy9NNSxXln7atQY4RBk45mGrj81alp7MRmvcmMOq2T6gij2zT9u
xhRAbwuDND0CkuiKy9usWk1hQnzHFmQ1Qljar/jyq8kLCwMd2xjfTWS005F7lAujeNG4UT3vGjZg
qPGZOwuiVx4mp3FLLbk1rL6lTbNzSo4JI3XfFgwfIN2KqCjpYGrp4N0nRExIbwbhNRBepgeVCfTF
MgjzdDnvLnpsKe4s5ZwNP/tb3OnILkCKRi+WvsJSpoKEAPPmJh7h6no0LmvWSEpAP/5MbyS4KjCk
RX2/jRIsXA7FUR3Tnm6uWQrFrlFfeGb/ecvBJiX8SGv9DGz6haHyiX6zZcsGkb8f7A4RHbk0Fhci
A+zV5S07VQsshQ93SfW8JGSNTc2r6C/R8SBnEGwWK1co3qh/JQAM0ubVkP3FH/e6MiPGyS27HvFJ
vHp9+/IXq4TJ21nL3M8wyQxdw5M+Ta2HS8RYb2O04bmQ7rQOvkUZXZZg1oTmkQceZS7YTI9oZGS+
Atcqfqdkmv9fLTzIl3W+Z3ZC+Qke6vaQkoNSwLZxEXDAN4ASl3Yk7niXs9WG00ERs73KmBmEmiQ0
PTo1IKFOPa2NNFTBiv6u5OCgG7xDu/U0Py1NsvnaJjB/5DlPDmvXM8Zk15iRIkJ+2h5nCTS4WLDO
qWW9yhCBOzfZqbsxdZW9vJVi79JcE8w00/kzZiZXgsEFNzp19m5tM5ohchgj1kWW6h/JEuOuwBW+
rQGzYg8S7m2Si6wYJKJjucu5Md43+ChOrAAxsCRf7Pi88ERIb1he1kEO+VQr25sxHiSslG98NurH
PnAEihJnTYhl4m+hgQrnGnH5jVRVz+GNzpHV/JeLWW4FpYzvv3+x7bFvebhp4FlIssNflgzkS9B1
uYdQBo4Q1KYUyzCJwqOjIUi1YOXp/rx6s02dTAwTK0Ou7l+LT+RfklKfhCIvXrkIcwDpLZ0cxiE/
a9rMpXAPt0blyyiWrvziJl3NAz8ZJFevTajKxM1xnfULDgYXTGoTQACJrWMg0verW9metUAN/ExK
r+p8hnBEbNgXBi0oXYPNyk0bBwdO69US/BDQNQOyNItdmrxSNZUbe/GWvugcFpUcg1wakzFc0fsN
naODG+oWY9h0YOO6P60Rr14uwn9UyFvh7PhNB6nTlRr1T87amWE04ObwCO+XdvAj0MfZKRylK96/
4GQFDjU/7Ldn4u2CTPJtFQtfyS0dyQvZctA15NcJhfAcqaMyvvbZyi793j254wtjjpPrYaF9U0dm
pfppgTqx2mLdTKnG8dKFyN0OVcnjLfaLEBodV4n9/SXtjVM2CQu2oJYqorC/+Sk7c33UixhI8W4m
REL95x/Y0HTEe/6gtZnPMQ9jK1I5d5UIIrZc6YLAK0UE5Xk6GPnEEsf18M16thzHdhgfwes8tPDO
v2LOy143sNbpAJdcDhvVDvzlrCdLvnKGMDOrruob5PUdT+djH0vU4Riz/ER6QDkYj3VxffTJe+rA
Gwr8d7IOe68Av13SnB9cgQgxO99namL75KR72+/yZjmP6NEIBkAp8qZQKp8FV3IUaSSZrP/qHOA6
5zBlz4YWtdBwVCpqM3XMrXCZHXYuiC8NLGZEAfLBljsaWgBnsPVMSCWDP44Yr4ksCHtgG88GMDpw
ya7VsEEKaH6DwJqeECHbc53D4NVUIR3/PH4c2V4W59hhxgdJzuqpjcxJfxIm3n/PUzXzi0tXXY9x
zyJTDGmG7/vDDU7Xu1Nv4XbO5rA1pDOMb0fV4/zLLyGN5KleiQ+KCKCapjsgoI5cSGIzympe5T1O
jA2xrXTLWzktPNzd+611DBgRmHtDb9QvcJE15KY2q3F0KBOr7n0BOBUk+TB9C4G0xj1RBGUN+pEW
QpMcVMdguzmgB9/HyrIq5xIr8c91WnGbVUmxYx7jvmCD3A5dQ/Od8MasSE/ZGP4BEcEoEXpaErtM
PdMbzH7aiMf5GRYlrhemLxf6a591M9T0JUglxgc2UO1Vuxn/BZkjiMEpzuBKIdhAY07fPazzuwgw
Z7AK2+4YAec/jctuQCbA1GxO67TcFtxBuua3s6AwwfVmrEZrBrpv/KYVzaKx/pVGsnVQoReHk/Q6
GkbUNy1AwSIOD+vQBZ8E/lhCWP1TJ9FNO60REpSwKGKtp6uF64NGZsn44T9jqAQQ9fMJOoZToKM9
LJIy1lDf5seKp1ACVhx5a+vaYdE7mpTWP8UVOpWVuDdM4v/CzydkRSAVhxlpgiixxTOG2wK2IeOI
Bc10c0NAsVoNeKFSDR1dRLgrubSOQMQANJHQf+6gLPoJctcWsNdlzqe3DTg4BrWGX9JxgzqQVvXP
IPPbAz1RuvXEDOKZsLvB57dIhjjXwYy/jlgLbleUm3lZvbEH9mAjjz1tWIFYHgCj52jSo38AebJl
jdgDBU4/zYR2kuvRS5TCGSrR47yNB3+sdOfCM/ZltpjzhRBv7Gk49RAyyp9qD8Vb1oavNVcQ2WUi
W4x1yyEhPvd+6nLEAeJXr6HkIGSH6jBdX1WAl9C4NZRGshKzieelkyN6HdrXm6L57FzypGYX7781
mCsrqy12Ja2M4s0w+ZX2etKz3trleX+MzX5RbKONCtlYBh/A3ENcpTnIvD698h2bI/6wMHl5RvvY
7Hap6heIh48OonLWSMRdiV7Jn0ZFe1fWV6SHEyNK2e5iy31XckOpQnO8GN0YLD1lN62UxDfCT6k2
Z4DwEO7YzwHHnQGw9VaMqipI8N4HCI7DC6DLdRSBLNo12rPI/v7SWIYPlmM9DX5ddTUBdMcWdkiE
MIo/lwM778rw91OPgvXejNq4Eo5w/NdDMfP96QegaSOXiq2YUaV5xF47CRjKK7vpJ71AQFPSEyjT
niPwNUaF0UKtVMtdi2JtmhKBJJ9qq2tLE8RE6xkPThxPbCsXQAkJRaqelnn7rCMwhzvYb3Thcg3G
EydFtaeXpQ/H/deI3pjZvcqXkRmhlJsfnqJOkQS7/DoHUucKtrvOxSeWX+CvFvbHkEebsXsjqfni
ekzHcXZgc7qZ0+EJCpRhwwUGG7F4r4DVn7E89xVfgco8RaORhTkY8KG/xQl+wa47cD2ntHiDipu5
9teaCpy86Mu3u0yXWoh+rAeL1fwogQIxyJwVyATxosLevNafABJFANr0WwIfXDDOOKLBWORFM7r2
2jaVb9K5uqj1h1/FjtbQkxz/6qMS8Yk0W5YX7fu/TWXIw/H04Qt9xOeRJqeiwyGzgRg6icySXHUp
AY9HbdqbdkDevwBOOsQYYeTsfVH6k5iqgplOnfho7r9TgFBhQxvPN0C9YB1XbIEi/3vyhJ6Jr4ej
Yl1yK9flAXe9/CcNihIIvSrcVam36SqggrFsuyyuS9EwZNPRNT5baOlpIRCiUHLVv8YG8z8JA3Ik
CfZrqxETUsfmqxTyJ59RpC2gAIAdPmbCT7jyKkUDyIWMBVzRZO1l4AkzU9yF2Ui8AhXpZrbwE7Zt
gngBAYA1Z+JAfoy8u7yUV70eEvQP8NH9MwiJm/LyTyTokV6ZA/uSkD/nOZ3ZakWDfzFFCQcxGmIs
nx07cQCfy55dDPcBXD6rFvvI7y85W+ZGPJfXVBCNiBMRzrxDJvd73TRjbOMDhuRaLj7Usds7OMhx
BwIk+5yOdpG0dhm/ttSjoreIiHsSGFryhVk96L2QuX8/K6+C9JEcySOFYtwN3RFakAjMKxrtnqFU
1487o2Os74IfYyv0Mr5DLSgf4Gh9QjJhVHpk7V2dkDhYy60IVsg/HcO+NmNo9FhMwYDkcsHPOyIb
pgQdpp2+Q4Y/hbx8MwXr3f9gDvM07RR8Lq3ltB1DbwtAx4j3PiwyM6GfyrzhZOqz9xPRl7Hg9xvI
fMqPa8xmGix/WigjvkSiI1eTiiguwzg4cIlfxcNqYHJ3Fx+5Ongt9GabD22TDRzkG6/um1uau6m2
0VptuKJHhvKXduizUizc6M7vv1lvvqIKU5+JhY/Nj2jD+3vwlIR1vz7+kTX99iDIfSOwM2m5ydC7
bfMzeq+YKmYHeYbsHFFel301vgqmxKmkPgYVUeGAiu2rVt00nlNyfjbb59k/7fVzq2CNmY+3A2zK
4cI9U9n9DF/l1GOByMu7ZVb5GgymoiDWWxK7amplL02ALqIxZPHcvJwI94f2Qa70tp3UTDEgOuTt
RPgIfHXq/wBEGx+EGU8xsTJvSyJdeGpGgQlTO91UW3ID/xhIXOrY1Ipjv2OVr+AWVHoumtpj9DrS
JJCkA+wBl1exu2HIchVqkBjlZFf9zOWdL4MaSl2ED7veaP7RxEv7F+oIhJHhHokCFYBmCz+j3aU1
ODGvInATpL9Cnltj5GIsK8Ly9dAgq0W2E0yn9BjLdq4a2JoEXPL27EzDT32e0aauEVHQQOcP2tWp
Dj6A+RDs/O7NkVSURx/nalhfIz/YLdZLtA6fLUJvcvCeZgdVSo8dtBy1G3JsjTZvesZ3P32HHZAU
iGqMkrhMeqzqZYd4IrAQQcEkVGShkniSDbmbbbhnDRzjbIsucpYUOWf050Y4Xi5HfS8Y/DHyEMzV
bend1Rn5Y/gt9KDGMGeuT5z2WeEe2Zg09/rT+9jJqFcZSGnECgMNEUtyCog0Ob4I58SAf0GO2+sd
RobMI7g61BeSvbqWphRdrOB2o2gk9eee8zuaPgvxueFnkkR3cGsVuxq1FJF5U/5efjmyo1T7A8S3
2837PRqQ9QgDRvEZH7PztXX3Adb3QtcBEsOaIIapLmIYUfC37jiN76y4TlH419LcN3JKJRaIoCie
n7PbX5TcLv4pusKj8NV8Y1x8X7Z5iHYH+lWp4J5aN5OwA3RZeT5pX2nEBQBMBypHWxqJNvLV7jvn
aXyNKCCkkYmKWiUgaHex9O+40KoKDyts/zcZ4aJZuq7ieZt6dfdmAzndx/eRnBU/fnxgDrxtMzgt
cs93v2i4d8jw/w6sVmwtih+5F+FLI4rpRvnnxrHzzj+8924rmNd3XJ/OEiXr0S6TeOrYyinq4xKg
urTQIdDjCX8dHdIC7zqI95t066QGTuxiTE8n+b0d4cHrZ4yB0kDfooY7WVvlymxcNVrJjAjro4ft
Cjb3OTG3NShoO5u8uPWg1EvSk+bFNyEBwc+/EYWzPNSLlWgjwyxcqIBK0mSHH3hjcO7rTTsR7EQb
2vnXydWxqSQy890ciHgiobXRdg1k4DuoBvlWtgG/3k140pJJ1kfnog9BABrmrW5VMtk+8jliGmkX
ZyOG07ZIOm398xOWmjoLg5r+BUkHOvRawVJPnXPsHjlFhI1lXd1wYnX6sNaSogEAAebvsf1eBXa8
4dmLppx/xzzDgBK8wxVbfe1n1G4gHg34sQ089LmQrc9f9BexIePaprxD45+LIiFvRpF7KPlhl33g
cdPyY8wpckAcn1Z2yul2pJyiqf1LLCT7uEAZkpDICOkLeanGGdsiV5Ix4z/QYgSNISq59iwDE0EW
RZ8nc55OM1AFxmxTgiw0GASIiN+uixQtlq5La2wWCCKTM7GnuadqzujnjRkb5mCGfFkWWkiHo53j
Ima4rYxEUjWfDSAAoG5OapO9XEuq3THDtIRME+j6RrhReTxglKUhWjm0Rt/nFysKQqjblnDEWYL9
Fx4B37gybbd9JA+n0Q9AQPZCaNeonamowE2HhVkRpKojNWnRAvHmnaNmlv9hKefh8yjqy8lpOx/S
Blr1oOfoQKXEKiyQAsKRk3S98a4TI/wpDxkPAnOO8aJc11mMcbrI2mYONB5Vujh306QRbIApvi+R
wQZQlgmlyvXee72RsetmPCk4QenZ1gA2U73eT2w2CeMextawUOSl7KBGxRwYUG7a1syJui7V9JII
A3bqLi8KWJTRfFiMTqeppuJLfiswTDShHDEP8R56X2CaZKdEA6E1FTMXJIG/20nK3fX7Na8x+Naq
rdS0MtFQYeoLvc1jC3DNLYCcK4q25D33KvvjJYs8oVA8feEFW4cGY1RIXCz+gbZk0UCnsrVOtDa9
FbZdNKFJHH7WSWUoR6hILhMV+fuIewsteXkTemzy/w0rDjhdfCddhYLq+6SLgKjdQ34vfgYnhsCp
pktEU5fKQVjOV0pVGoBU5Tje9mWH/41hevYyRUliDJTon5X3uOivjcPlK+5yHom1TarHwLyoccuA
nMx9ciOUCJwwW1cs6zToiHW/6+1k3jOMfhGvMOgFxJ9waRrmkVj04MH4K7kKYbn94hsVWwhvGVGh
cqfd0BfmyzuXKriuHaFn/nb/Lew+lkR4b4Tte0HQNsVBbguyCBIULV8RzoD/mmtuOrt7SF+BSkM9
2zvQMBS9xMMVZZfhZ3PsGH0OO+LYErmB0jvlYl6uD+3Y/DTSBLH+M+n/rGqu5NhejgKkh01YKmKK
UBXcvvosgISjMMFaAWeskjV5ZWC6Lqd/SHx6Mp/Psyt5il0tXc3JgCNBywAvY5yBGmvDOmsgNqxU
o9AcWSq1O3holT0UKmyeHvLaLN/bg4BxOt+a9izGz2FkAdEED4Acgsc80hxX2ayqS5ZUfo5UGzzh
9mxz8lUjdz8qDxdFAILvF5E7C6bZkLjAacRUupjhPFT+tks5d3Tz8vchvJ7r7csqkjoDYdqFQ/KF
STn33zbJJ5M1eSW1jcuM6OFfj367iSPMb/IShZ9MG53533KWZgAxzb44M7OakqqYDyPsGrJYEi1L
V4EGwLieLsvMfaRvm3dJ7FgRtLgd1p74VkH5uMonHhvVlVKHEzeDm2jWoykuFPTG68b4oYvrpe/Z
t3cBxznYOiyxMO+SQgMr6ecnWs63DLMMt3BT8Jm12Zn8mJbtt/d1RK8p2aEzf+eClatyH2Qj3GRj
P3vcGtIT3yc5R7uCspl8xwjxHmHvk3pfzRyL4NAXPBNT/GvkViPYV7y91rp6rYq7z6YA2VVQlqQ7
3/ynF+vD77ZqMVucEKd/0QQ5efbFMmVCwCpvVt79MXeL9wXHN3EdrJpnQ7TPqAKyvpx5F9zvQd8z
e9g79IbwT9ppDM2/LCeWHoPUwDgbgxRPNSTuNZAVoYHoAZjFecaGL8jrahoc2+3Mu/qN2FrDhUIq
31KVSbOeKdRudc/FjeDarIc5lYSRjcZ+6yT5UMgd1ixxdUqZd3klG77bFDdHuxDUohofjaxhzrPI
TLD7thtiKIVl/RuvYfO3XNXe53m9IGGDNH2WDAufrwZDr5R7YzsGcRqwAvVmNiV4h6q0A9W+p2gJ
H5bFQ4ebQoAryf9tygYN/onmOpVPl7oa4U2uhrySXZmEsRH99Ld8++nnFxZv9WBWxycn/HEFNZPd
mvRTNheuac3gOeJG+Xi8rUg78y6yb1drGsyh4o3xilysZrdd0xcgsXIb3tekrwMLere1ePSX8INN
FVaLqKVFrmBSZJTWhkSeOLSF71DE2JIuMW7zdNHdcXGni6NLVifYN1UdCtQAIbEVu18oOTghQX6o
Nqky9WXa9YYal51eAXAlsQN8NI/CvGz1AyhXBsJTQ7vVYEHurpIKxVSw58W5MEMwwYZP6vnTGfbO
UVcr1frKPElIqNkQpAS5xcv6x6oXB+iY+adGjNDUlOJBIHdOiY9XY+z7OGFGgcBgM54akvaoZl5t
y98UY5/EAjwWvGK5CNlAo+waeAsaLkxG9LuYLJMmX9Gx7G62MjxBFobyJ4lT1ZR4gkroQ8fWFNZu
5vvlDuQYK3YJenqkNOMMBds9fgkjftpVpuY5pVcoceXu4NWaUozXjM0BefhmGQ8R3mthCU41uztB
3VkNJiDd8FXgH/h0027l2tUVz2WYwtQmocV2bY33wDO4U0OT2vcUhm9/3N+EtW14lyW3kU6Bsf44
+bBKrnfRC82dRGKsBwrXlaLJUXMoELmxug3oNKJHSGmnSPd1hrl7V3418/uBGV+0jYvQAemB1DFz
/Id9fHgatMtPfptr9llz/FN4n5rnvH6948J7qvmSukKqK+rDqEPKChekyf5K7iD75sl6KbUUgVfV
qxxQxikaRwaOU1k+E0ry1Qmdso41MeOST4HpZs/zpqW+WOgOfw/pz0S2KXtiPS2EoeFeDv7b8Voi
OHNfAC9riA91EK/2AfrpiUzF05TXFxNH0mjFJkIbbgomBWzPwzuRit/fPiO/1r7l7Ea5sokZUVbz
eW4fCGwzmnQwPaswUX2WMsceF9S/wb3RazGLZiZ6Hwq748x8mML9XCXI7NDFqI/JPaTQdt9rXToW
gvGy9qRhcUgLkQCWcPfCyWwBJ4NSKIXjEvl/Zsm4ZQZMeC6ucyubXPQw/GztFqObYLzeJ5v50NFl
mdGlqPVQoQi9aqgRLVRN90vI33zZXAfKG/UcysJlVcS2FJY3ARz7+vsdF5qCNIEM3PCHt9Nra5cx
ngSjr9Q7a2DRIhWyYOxadw2UjyNNlmHrLlrJs+Jsg2ZdcbLP5K2jYEeYPhr6c2Tya5DSImofTDvM
BgeKwDGWBokRraszQhpyQsONDBpJ9H0vg/zh7Zjp3jmDYohUZG4fkAUmElxRjaWfjs0LBatDizKm
YaiMWcJ2XKXG9IPUZY4QYtLkkIIMOqugs852FJhsQKAJ/IcpamDJv9NzqbdlSe926RVI0wMdZtjN
x0L0uGpWYufS3fHRWtAEcR0QjnFt+9whJhteY5B5NQ3+3iSjJDqfOiMTGNnxwRx3toGy+O78EL/j
5xn1uttRXt2kfCdIoCtnTRvSA7NvUtfmm9uRMrWk1RidZgYbooihFBaU5nZMuTVsLb0A2e1yFv/D
0Hlv5YpbGkSr7vtaHby1/dLCFgiEhN/LEkzT4nHIhT7/Oa73Kxvyq552pLcSBgxDw1Oby3MX/LRW
F4Tg+TVewYbBsRQYsm/SFnvhh8v1nnzcBb5igdhsELcYtFCcaptyACRvtVC4oifdCHelrtihDmRT
5OE8msBLxxvr5z3RbFBwiui1ez4oHVqsKZ2+8xZ/Njd1m0mJXNW6UAIWndU4YclonclCRyRbsFS5
5GP672OdHOM93bzrXcC0r8TkF2/QgmE1l/4NxUXEdqVyMYN+fWrPqd+biKZ7qy3cT3vhqoATE4hC
m5/9hAM5GkD47L8bX3gEZk/b0/nkBdKuz9HZ4J+EhlBDCq/K5ckparo1OR6zL1R8L+twuV5xygvI
d1JJnWr4xJsAe4/9xvAPP/3AmxfCI6uDxPVso41o4updTJw6Ni0JixSqBi8qdetD0TnRi5igGakK
nKOdJ1d/l5akyzfyt+XJXVBC+08kiAh7PdUBknEvV47Fay7LcyJSoEPITrrjE2TvQLLkWw8rymyO
2N8hdH6gZuUq+CN6Pj+kQRSqYvJ/2KNmdppH4SdJgmS1ZrPYD1j0Xs8Jq+xXzVxxEG1DhiuJZ42F
mGGppjU82eC4Fif+Y6rH5BCG1UobdJyCMs7E/sLvfbZQM0jgbft+qz0tNZt7i/bw4GUn2lkZea+/
biRWPrWEj574YUcYtVsu7n1pvDPCax1XMf1eijxUxXeo47ZUpSskSD4lncv99wx0D0xjYrH8Z5WX
43speoXG3d6qe3C2Go+2krhL2RacXlD3P3OxmjSnReCdLTc1QWpxt4BzppsWmbQsMDcu6qhG3Owy
+vd9O4S9uw96NL/UxBtyMf1PnTOaX1a7IX/KCZQd6tMOz0/QcWhHmzVeczvzv1jbbPzd8cRMsYVd
DEbf8v6SJ4tHRfoENCG4/H4NJQZ9BTfyPwls+mGZXf8vX5FKFtsARMXGKWXkhZavdCEfbcGX2j0E
b7Hn15cw2k+LFIHDnSGTT/73S6Pg/D8PemEOaw2jum19rSu/yqsbddzkmnVJhTTrztQRxweHz2Ob
zBmxwsdDDM90Uh+FTozXye1gLLQsBARp8S3P5+x9vlxiQagYJLHInHkBozLw5H3RLxALjdScCexN
lYb74lRi8rP5oSUh5Slwokv61Lw5SRbdkGSQyKz7rf0235laxX5SwEaD5J8X+LJAhXBwlg55lAse
4M4F+GCOZ38XX4Ov8PTjq4XdG44DVPammnLp59pUd6cEF1x0eCUBJ2Mp5x1Wk4BkPkao9eammc1c
NOEWwJ8NkL9g+eHZ8L2GHnJsPi5Vo59rRH0Q//SsFXDc3XkxicIx7z+AGgKJM9wXkBB3yIS4jHwi
JXkBLaSOEKHNwCQ/6bhHXGU7nmWCDiU+yDxk2bvi5CPx7IXgLuxS8kuYoLhmgXt+zdZ4QXIRvf3t
75b2BCogQUqAmme///DRwqom2+IaqivI+nC8zyalgAEISKFN1shsn3breTgmNZ16BkjtTL2Fc4sx
ptgoQS77N/OfbmdFefKE60iAUMonIBoS8t/CX5HpxBOTjnL70AABPopkrVTZRci/zyL7tIwV9Jh1
guNeSD0/kxiQfVXH+Z+qnD4hpHk1PDShCXCABbiFynj/XcaZOGdEPi7xiMUb8srdXlL36om3e2ix
VxYfV2WlRvThS2HMzHhhsE6GfjlNIb38mcd+/OmzCVIZH5p3Har1JrReabd97PkHdZn7RDLI6POH
Prq0K+6h750xRRiUvcbaOhPr1uP9+JxRaLcpal3dWocRHQSSUJ+zKoCES2r57kYi6Gd4AlXc/RgO
jzICHkGUlu/t8EmIwms6bIcqXrWUeyHFAPZ8aI1k5mh/tRWbA4OK9rvj4eBmDELSQMADhAhx/ZsZ
eCj8ykQvk8gttbRkdrTJoPHll5i1iyWCH399Li0xoR/iDKSjFQ2WGKvrFR3ROnFZMc9a+D+u86tu
9zOkeSL1cSC5aiirb0pcd7Xfpqe7BS78DBsB+zWLTiJfEO+pdfsOGoD0qhAx82RDvSAyCFQ0WBLx
mDLaJJOzCJNUuRx4/8f5PQGjURpV6ENebwmte8bOUG96tutZMKpbEKShcv9uaWI3WMJqGYXiZ44F
YGYl+OHx0cJioagHXvC/rC1vG3XolwRS3TkAAZs/9zYTIxZjjK19CqJlAC3WZ3UzCWbddOCjJC6J
lzm+nxNy1SXvoTh3aX7UsJOX+Q2v1d+MwWjgOqbQUnFmDCgu95as+YOtL8u1C7YlGBsATQKZc7wW
nxeYER22UxfV9GL7uGRJrVWj+sx20KCp5DY8Tpqtc+84Xg6AA2earhsbzDzO9ar0C8hHFSyTtT8k
ivW9zA5u7jkUR5SKmU1DV+S1WrHMDRzLdnH+nUwz+t/+tDAvhjEQhGG1W4IRgUgUWgRwl82waU5g
WieLnMhsJvB/C2Fgo2Npc9ULXInl2H68MYtlfvxI3ZmNXJgBlxz1Y8WHN6BNN/djCh5Y0kdRD5je
Ko4uy+G6pCbDeMrNYs/saAs1/ov1Kw2+2ZDzmA4B1RgV5twapyM8UhODV/KN2gVEFrIHTN/sdvqZ
q815brvyqdfB5pHDD/gtvQC4BvYR7eBtyXvG6s7qwOiJb8wjhVwBiVx4nDu/q6mwK33VvxX+oTVN
qhUHZHDmRZ0DPgYwKyKexLsinQEHlpLgPL0xm59pbRQQHnSqlaV0HR1OjQQrs148mXGFe0P8hiH0
VyzHVrncLW2sjOxMD6QTire9LBmuQtTZ6NUJp5EEM/O/lLwD7Dl7vcU68UmhJTwMyxxUoliyDfPL
vga3Bcq735DWIuI74RbW1m9V9yDWFOmqK4apzlDpWT0PQ5tyxanYW5m9j/9WAqKcoydNIIQMANVf
zjVmML/Wb9n2K1qBdkNyszpc1j8lLwePphZ00ekhjKh2NCXJluE/ZpqvLq65vAMjjFfWbfS3lK5e
czrzjw36kgNBdW1nGe++DHSrqmdRgsGFCL55fNxW4DJ6MdpoJeFRqaE7dAkYpczX2+Kv7X+Y3U3F
mfe69KR91hYjWddX2sZ1mZ0JaHYj/7D1dRxl8Ejq2euBrULuHrRwZCcYK14fyp+pBFjH6k/Z6+4f
gwDxsjulP9V8i2kFGyX6i1B9u6mPCVzPZNqndu3L0j2RF9AtJJXGuv2kwHd0ncPkc39jhknWbrBu
eoEJW9NQkn1+Kj9WLY1TFgTDkMkt1O1BCQp+/RN8Bhx3+7lNe5+jXpyS/9ENxc5GViNCOvGU2zm5
LUM3vc8jB6ZcU/MnajDxwXaQrW1MXXiXlToHXDr0DITmXwrx+T7/eOf3ydd6AQy7g0WeaVGTPZAW
lscoHX1dlzZE9MBxzdKZzVXrlE7sAozj249+jpcW0eN3pysvx3eAaiJGOAkPFqYWl/Vw/lBbrV8i
5SEIfxzeGYsRSal501ahlbvIrwn7/tddpHfZVSmxdAiahRo7bxVn3JuDiE2RHVg5GYSZ0XXpEmE0
mN8YtAqCIg/yZvGGnteP8omWjodL8pXvfgZlJYkeFalZnoq8R5kY4Atsd4SawhoT8xswfRuu8Xpx
8hBWyWPHQAmBdO2h42W8k5o4ancn7OeCsOurkiJWo+7uwBPo+ILL7YTXIpia9EoHOvVxTylwOyCk
sbge1t64eROeR2DYe4ZfwtZhXGeHo7X/wlSl5lL6CBS5L/p8lMzR52L62lFXqKICwW0WbA9hpoun
cOFBUMXHo5x+JLg09/Sg6iKXGvmALsNMqF841YUSyZlZk5XTR11TvTRAF5XeddLxfsRX68rIy8iS
U7k6keZhLXB4gTPu8mgRLLkEknqXGM4kplVvPrQOX5VfzHEH7uJ6t5rw+lmwKssOLSCkDM/4r3WN
ubQR8DGAe69lSL6upib5GwDcsLciFgYcmt/FwC6UOZ1iN/dg/7MB5jYIg9Lxu6rlzbzNTCzPITh3
O37tEZe5HiELNI0EW1PDVjyem8VUBxOWa+fzPKXCDy5CYIg69JO9LlMlHzfFMc3HpDmBAPtAmIeD
DYe90SY9nxuAKtboNWkSfGyfKOmK3PNT/CBN99qo/5BaSWhwG0stUG0tcVNFgcVKbZnHDzhk8Sw6
UaxXj2DbFBOTuZzizQtYg+YXLSh/bA5FbLM43GPQGIAil0Kkh7hnZPyckNSaCLsmEr01lk0RaxZw
JUHl6h/OyPJetLXd+q+AXfNxOIHa6bG+uIrcxFUS3L39l82oo5uhuiX1FMIH+KCLoYegtZHzx/dE
hPY9tSojrxU+LUq5aXP/P1o/jI7asBOK/BiaN2hGvk3T8/G/TqxvHuUpXnx6yFx30Vu25eJcMtcU
IPm9oxvK605Sw3K5LnsN+RMO5HQKDmdcZERtsGb9huqt/+2HQTLX6CXfxH37VJv1XNiw+9nX5Ovh
tv8+yju8R/Cyw945iLrSmE1ybMgTUc4kM1C5xFzgv5ew4yoy8TZWB2MJHCmrrZrNCAiRph6poJM7
azbd8VTmPGwZz9PfR+NiCOsPjVKm5bZYCZFY8xZyuRco23VU0PsIX3UQpzLRjEbB9MbXFA+ewcLE
lLpLZautpKpPy0F3ZJCoohl/t8YfsYaAAKBUTYUt5VeNXcHGrllVAn+Fm8w1Lv4M/6lViIA8Xxf7
7jaxG5CQWmj/JXH1cAXNya4n8JsYRDUItCX9hYqTgYtVe8N8J1v/sGHWX4F8zJEHON/tY70hWeWy
fEQxKvPMf6UGzQyu3zykLE7kCI7R0FWPyfLDzx3bsF308wAopm1F3ZxKwA6Z2efhBGLYRUIqblFn
asyyNihVuMRx8h4ofI2yKr761T6XYubszgx/Datb45W3wEGKwKrLcWyRMrN5DCfV2iQ0rN2Cqk/M
y5p334Y2s/O1jXvA6FrdtVWx+raNwPjVDKIU5gZowCLeEiTXdz9yLc9eg92VLBLb1OxIPIhTN6xD
340Q4yhqw4yG8qdhsLJK99FqxmYD56BhMABMi4YJ9XX+r39YmhikmQ9pz9pR4MeExxoerLsSmaWL
R1odA08qr1paIpXqkMvuyID0GJ7ZPifF1zaQWJz39O6XurjvyecwNiLHXSmHw8H1ZmKsBdDILiop
nza6P3IlaZHuST6nQm3Jn1NF41p/pFyA11q1M5K3YCCczUha1BvwHeRNk0NkbI6/ZZMW41lj+05s
OxcMYH/DFgDVIAD4y6c4BGO2r0U9NqW0/QvCM7PQecv0AqJuGnbTrmfLv9RJdh+cniG8y+BW19hG
SQhAj5tYY557z3iy2iuH/IEXA0ycLb1OinvPzkKXEBftCajC4iaL4QIvncECoRu2KTGDFXlwYRiC
muY6pwEAFe29PhdcSTpNpsYHMWjhNhpfJTDcHnduO8+A9vv1Rx5vP6qSneJRcUyrjc8EK2dXG8U5
R6C9vt2PN3lbCC9iDVtIxVXBbdBZYFGJQ8ucjme6QVkK7A2jwpO/iKFdDTKbapwYXmLMndYiZ18T
qt4NZmMEqvCJ6TEAX9cG1YsjFfP3hxeGyCPs1T4gaVJfrPiGJQervNLGLPQZjEOJJW8ZTCDZvv6R
uT/axLqz7+CMU8kq3zyHKd91Geszt7at/MsX8BEcYBKhtWMnR2j5MX3785WGcHt4549xZdbk0Vo0
XzVdptzBx5iMggLcx0ow5tmzbkQLtkOx1K6ntakjzejvzxKTbMNFvILxEydftKMGErcHzvNSZt/6
aYcdjZEmAsOFmCHEkcKZufDmLwyo58MaTDTdHxEn2P+QFE2oXLcLxRFPFwAgGUYd0Lsdba6qQo0u
WPEopiqFrc0Pk5z8jRIWXzNjYfFbNbXl9KWtav7ldCEIW5hjfT8d9IIF5lDw+eK6rbKAJJh8cpWb
NxfEVqxBSfQkys4Idj3DQ/xfW+X2LdaE9hKPvrg/+Zpl34yy9NQKysYhWGGg5V+g1w6+2dgBBA0I
gJBRanBvs6R35LLVSJlzpif/WtGKEOi5a8uBZu7jr0s2uvU1sNJJzXXFi7/dbSKep+nwQY34wb7W
VKfHW72Ca66T9klXKFW0eqU0/AOCSHrZY5a+DRYtw5rC2isZbrnZ+oajJFz/efS7aoGhI5MJYl3F
6EwcRWBnE4VZxP0Pq6G89/gjjvRiXd8QSLoA2Si29ftLBOHHi04sWK5PsHumzKjjn0iiHSiDs8Ps
odyj24Pf3PullGqCxqi4QzZVM8Haop4CJgB4dL2CsnaTN6UAcqc5EVw8pHHNoQRnGaUwnCvX7wBz
j1ZVXdCIR85rn/p2bUxxtDDsCjliClka3ShA1mDVmW2tfQBQygJEq/YdHVO4ds3DqpQzkm2O+o12
u+x7yMdrYRVygUrlAuhAr34sbJ0sViqGssH9QiustQcMkr2P+kZXfbIQqkXLXYSeqszyYtWfguSE
a/1l0x66DYtdfeTVvTDO94A/DhartARAp9L59XMzTmMNzavlJPZHyIIFlQMNFslKVb9/2tVZzip/
kRhQRwHLp4OPRoGRYpxmcsiU89wdCKJOJjtN42gd6Nol61+MU312CIM/7NvGlDYpTqw2LUFIhas0
EJjMB4BjiDPLAqIGFmuEc+dwP8jXj96KzWiEfzzmyE6h0N2exr2gZmlkYhmQJ9rrFbWylj+qe6WT
QdqZwoNLNUj/B4m4OK/eq/683x7N+S4xy9C6HvJPU9Cw3xVnFRZBv51JNxy5hjBiY17qYWDYK9C2
N34CYfADRzDQQA4FLajcVB/nsaEUPNUwbicFwbzekplGWuhYggj6Xgmtw5ExDRrnRYBSIq85eBMV
7T7K95+65HdDTg9sghV4VI+wCcElJLiAvZJmtwlYjDP0YgS93d+HxlpHIr+xR2/yKmeiqkmpkL8a
WPmm8Hg9Da8FdyyTtPcKQoRSMFYsUfrlhvg7YkiV6OMZ7+0FwyOjMUvfyAPUF4cqH5ciY+q7VSCG
MJoIimIpyg8+IVd+IWkavMMkYEelvU/fP/5OmFPXGZsYmqyaH1NlYho6ugQrAiuzINKXMRgfSo0o
z4j6JKFNm0SlWun451b+91KKRF9CBpwEQk0sheT2mzwGOU+QXtK0iyTAkd8zLV1FA9Db022tl7va
8oTddeI3duDQokl1NVWrKC/yYQI4Vb0+Z0FJW6Acrz6AMpyaB/wa0TsH/Wp+KvhMRN0uDUAd29XG
u/jXKIqCFllXycUcV0ZpRBHdAPJS5VOeb6L0cS8YBULbq0wsRHw9RPRrAsqmglV4/BMJ3SPJrK2k
eafTNIRhA+GGz36cbh8vGI2Th6GlsGxjC/5zoNxuRJ9tq5lYZrbKaVTasb4BrzdFDwy7punLsJ3Y
FnuGuh/GskTrOr0jRJ7HuJNJPT7oyR4qbsc5EA6fwuhgOeaDndGsL+uOGlcYJisXx59y09dJuoiE
diYvcpRCsRIAYJqoJCneKCsOQ8L/vifCcPp3GCH46+V2xd88flaXUarnXFUKzPyGpUkKjQ7xDF/+
4UFvZMv69hoz8lWTZTICkxJWSUkmpFC28yelxy68OVOI5fa+PKCXgqueiNrL19pTlcEwjkeN3oey
ayqSNIzy6Ab9HT8VksH2NxA2FT0wYsu/10L2IGxmjvxwNIsV6BPBpeiPkb7u3WSi8yUiBgte81Yx
HULKyQUAmEHNThWBCGzV5r148wyLvqQeoTZNn/OAjX+pEB2kWeGQhP0vsq7RqpyoNhUkj+/TPyWa
9W5aaXIyR8FO54+DrBDPxHFyVlgtof7C1sv7IkBi7m6b8MzwuYVf6Iu4wViHrDO8/5QH/N8gXzxP
SO7oCpVYtyjLFW/NSlExzilkRjTvo4P31pFG8sgu/ahljWMXY2MckySDq1AXvoZ50fm+t2WddV64
+EfNd59R2ccEMZiybFLwVNoDM+UX+xRbc4a/sRx3f5Db1JvBZoiIp+vdU6bzLvMgSTIGGhRgS2XX
lAFc5J53QCMbnOTCzJ6UyoLvOAX3MILzwCGHP+WUErrToGBlEdH5sWX/34j52eOpjmO9t/mr40lU
7VaYXnslKqSNAo2wIXJmfoXvVOXpqOhaN6FzAlZE+3CP0/I5NocXqkvXacJLfyHHeEeEUGhhhl7g
9rerV87zQrosifNsWp2CBWvU4LIgEOtkdfmA1NpwkWxzhrA59LYVXsfHwMReigedSRrEm00Msc+a
wYD0hyI/shtI8GW1QEsLBUTeGcdmaf8DGMdvJNrUZrRNOhC2u5GXRIIqGUGwH9oxspKA8CJXi2Hr
hMHqfNgvb+mkJa2ssbKILVJ2jJuihSjWXwa5IC+rM7kwUqHvbQmMc79bVkNCtYw22/BpZMhpW2gG
48FdgiIEf4l9ADpgYseSZsUm743kppfMTBY8rKGxu9TsZ9/sHaeUkHGxFrVo+7MZjYX8rpei6GyE
HrV0aSawCsxe63jvGuWnXHh2bfD/sSGOpenRrbYiqKLt3sp2p5QUiZ0RCRSsL2Gco8fruBxn2U/3
aQGNKdLmYpc0W6KndsQjY7uLpEnYpN4xbiDx5Hj2czQi3FlRqPmivRD/oOLmjQZp3VlHpzTrjww8
fyWRmTJpGcyQbhDFP9aH/O05GwJ6GCJqXpKQ+CWZw0zcbUvGx7peQoX9kLRt4w3C135So2v0amTX
w4omPRg8gja1fkZ7Wkgb9lUaP5HVrH9ou+3S5GKni6p4plGSghs7AT9E7NDiemWtN4cdzPfparcC
GSo+9InqBFpDw9StkEt+0r47LFx88z0aIbudgN00gz69T7padE+6tKif/F1hs5ukTatptU7VynYp
uXyZRvakJw6jN9hz1FBSfAeQisfEshZ2bZwv5YG9UWzbeL3wTbVqu//HIDMB69STf6AtpF5O04f3
YiDY5tXqNxN5KuHcecM1Fp02rOucdkrQgjSgOpAlNmCYOL8DA8RXIlRiuVB80IL3Ew61Ka7GO4rE
YL1F5aRFpv11p7P3Ox3xF8t0sq/0bDJxt4f0qyMtPGHSqL/2YgF5enlq6+LQqr7RnK5q+3cw7j+b
acfTCLzA6YbssBbbR43YxGi4GAwBb00OC+BQOB54n+qVL0VKP7xgIceY9PzSXIdvl0RFdM7N6WuY
xf/rylSYuxa7ovvD1x6uR5INIHha5GJPMtrfxXCFN/l02BMetvGgFQCVb7rTh/TZ6wvagR5fceXg
nh0bn2WQaZY4ZZaX4lGB4RzUGhlwijIHotJmLNDx4+3QaJuRtlkzH70DSXcgIqDARZqiKcAEWuHW
5vO5uTcDs7rAfMcFYtDfPq7tTMiP8EChRbW5buCxRWfsu4z2ty0xH1tPcZEU+h0yyzDIYl3cymnl
69Jrl0nKRVQhupue2j0gVhyjGOefKm+9pTPff6d0cGNHVgtcyOjzdKRYvXqFishfptqu+v/efbMB
rCX85UIB++s9zkSyf/fYO1eAmS7uTvyoShOBHeoQeLGEaVvUXrku7td3FmeVUkW86MPSx5j8NAIo
6uZSmbMdPHLvlhspG+1chkZ3OxnNd+bjnl5JvEMmJ1vwXGxmSjBbgY9+PSpyLQO7QtTpls65B9Do
ZBsMaWN19aJjWti5rB4M9rBwieYaqSQssYtvfWPCfzVANKnQ68fd7OiL1OjnZul4tQLMgoKdvzjW
Mrk6b1vo7kV5J04XaKn+jKwgh5rH5YH+OyR2rSLLIjYggY4F1w6DZvUC9kAI9Q1pgGuI6xbQEfAW
686wseydeO83FbHF6iX+HqTr4R/6EaPNDWdc2qnluyzLRPe+feqlfkfYyBJ1gLg24PFt+lYhZ7FD
6zI/HibMaJkwdmDGPE1M2Nm/7VvRCdJqWul41Zq7UAQBT1h3yz/sAC9r6ldnMdmPjIxxO4hfP8Tr
AqUpuUTQuIfYxc0ynZSO+EyrS2huyLPIGhD2jAk+S7VtAHJrhUHoJ11bwyEBRGQFadHCNeTzG0a3
W+t80b2rFeijTk+TcDfC20wbAUMWjSUC95ib5DXZt2SnVg/8bshDU7Tlgmq5QpOm3XhV0YVspgwW
7ZZNCHi6tID5ZkO19oZxnJbQr2E2rhgL/beZWaP+pNYKIVvbeur8GTTM1qP8uU/+xXaW/NITPhui
uZQAlA17Iib7Hhezg13W7DAO096Dzv2mNCjdB86rVkJfvqzs0oSirRmFjq6axB2sl+0NVOLCfKBV
34h27f2azBkeigPb/ZwD+6/odP2xwP4suCc/D2Gip2GhNexq7cKeDwxVIO6lhvMDsDBAqE5+FqDw
mubyrkZqUI7CgYirknSu6RbkClqIPHBTaikPhrQcSboNALrjM7NH7dbH2yM3TUtITFdW17e0oTRD
mZ+SNLWRbu+e68/fHRw1lBWsosncJtipCvdye8kcKeTwRg9lmDfwMcidxfuolxM0MnAJZCrVBDa+
t9p6pWoADV7JVeURsLws0yWdFokFQYL7D4mSLEypAyjlyWUYRpXSYTG/Xlj3LnaxPjqyic1oWbSj
/9k90itdutHZWPYIoFy6DsEK9Khe0vFpFLh6egn2d5bQ229gvYv+78Jrvv3Qak33PIqa/p79sPFp
z6ZDGkrte9tq748M10UuJquBwAyHGNwwMWhXm/x+q7bgjk7NsREW8Oj3kV0LX2ZeS2aS1R25aBfy
5MQ/WFah8ZM/s0BVtBaArfRVMAXM1m73JJbQNZpccimuUhAgVPZzfqGy5Sg9Fl1asPCLTFUsuvDV
nOziZRbLnMBNDhl/rmlTRPgG6RO5pDeBesdZnuYFDhn8fAwNJyxU1+ALxKDcEHPV7jG9LAaChjpa
XruKj2/EymXyt6griC2DQXskfESTsDO/jSpUSTjjBblX2/UVpxFq4QEvDYuu9ZgznmMANw+12fe2
ftwCt4CLo+GLRv0TE/PWD7lhQJ5L0ZzwLcw2+9KtR2qpfNkpCwejnkMNwIujINfB0z98kHpgu+7K
SR7S9wsl7ysJK0MRYfg1uiRehW/BysRYeTS0KX8GI2YDox3dlj15nDJFsFTa4tZJ5GIfy3L6pB+J
bpGLN1cbUmUoVkZ3HaEpZKMhXYLnBRlWq/9KrRU/N+IPGY2HEiQj1tVx1w4rr/4HzDvOUGziXDTT
NhcTCXUEaU7WwkWCwtDDcKD3uqKLjIdjTyUgqQy9FXWaqhyVXw6JzDZzNlgf8qObLcO4Zex6+DAc
RERVifMnxi9U+lfm4zATVvkBlHhQQymYzy7ciM7/Y45G+HgbQF5gu04It0/Vx60WKlKHMwASGW14
uKyK2zBasQxx6aW0qfG1U6611x22wnnbjA+/l7uUDkR2YSg+bo9TiqvFQuymEx0gobUA3A8reOUk
XpsXNNEBDtsSI1YL6cXp37u8a5NM5RYfiN8crF3fy++lF6yvspUigZz5wf+/jkrELRlzWJNcyZ7A
zY4gvrB/iO3iaXpAjVW6yLM26tR+gTpPIqjmFuiOOiKN8xKC1YkUGxbd2m+kbx0C2Z67/2phMKpk
+6M0LU9n6HZ1vKkkDUFQ0Objnz15jyaFXJKouQjpEDiGaGgOe8bwzhx1MwGugQsQGHLIrDXEM7mq
voVg3Je1uQIvx8IFcxrBH5/yvz+AO00VKkcQeHKDC8Mghu9xH7cSkQiZeR369CejaqyVnw9ex21p
UHpF05ZeIOkNYH6XbxNji12+uQyrouXIms4w/yDlNjzYm0e18349NpI/yTnR/S99zxZRR0KwuftT
e083Mas5pjJGqxjdjyCO2Kx+IOyXA+RZloirxe6eYajSpl9xvsfKFqsysnoEgf5h8a66fSzigxWF
i8kZtM1cLZQJ/aTRXEtxadmj9al+7svzhRmmrWlIX4YHwsUPg+k448sHYNmDcgsj8s9xer27t7gc
kMdqlhXg3/8DPXtiV4i8AppFE260uJn8LiyOrMMiTyA7dsJImicF+MaEFD2H7ArEn5fLQju90q10
SL3zEkmuvBEVY/W9yFmI7gmPyrkL+TDxEJcP4CMBSauqhG040H0XiYv1MJdhJksjTnPT3bqDNNpV
LyGSJdALVNItV2zwPnMAm8cWyT5a4iU1LlFWOb097+3fx3Iw06GcXrKNQbDD7tnNqTUveM7h7aW+
uzRJQWRibVEfvqi1BiVAXizC+dgXzyRCkY+A0VAxmwoedVSVzCxxxNyXvF7+1DAhiuYKP7uVPvqe
bR1PFvciM01wc44gCGxV7hvyGBqaHHGKkCDFM4KxxRLpl29wa1vcbBROQMTnEpM9GW7rf3TV/SZ6
OlfZwwouiaETWUXDMT6LUjFyg0fNlToxKesTXENZujt3uKiUtv/0rztLQ59O0m2FiYOUUpJfuVqr
c0XBGiAs+sDSxw3W7vA89R7TtHS3WF2VBGLN8cjrxZyP5piE4vxK40+1auLUd/56Pj2x3MvCC4lf
31ZG1qpI1kkkhpxOKnlpHdE2SzTuEwbKEb8jbAiCMtCwAHgjpVMm1iEPVKbeDsNLYlExNCQ85X4/
LRbo/vkXW+OdqCH9F40K2LB/Cx4aK8B5GQw21Ptctbjc9FDtlEHuCbhMDR2mW+AUGYlcPnVBQ94G
MPj/jRQpsuLVIAVgV2aJ2iwTMqxCYgG31PwJJNBNupaLRqWhuk2ztzTl5Z0i211RZkTNch8DQbQf
RA5IGvs0BAP245aiYISIaw4dGT3QnJo8skJL9ORSr7B9gwkauoSkrQyg86QSGnl2anyk3Xs3XT88
u4IIOHp4DBot8iltDKy5GyAEgNjVW0iwFjQOEnQiR/YP79vyiHd30vS/9hMdiddTh7f0vw1ExmlL
MYRJBuBw9qF09pO05q2jdhW0Bh71mwznQo98DQ+qRrIVG8b0fyPJNaSQZ+yU4Bi1wr2hAiIZ8grt
pc7/eMZvd0+IMusuP18DfZL3SBBuAJ4WU39HKeBoMZ0ck+3x3RIqT3dcHYx20SIMW8AxvVmpmmJi
eLLfcItbjSGPvxiz6k0ckjZOPl4cWAFwhraSDWHriNpNsnwnR9hAaZ2GLStMy5rPTJDOY3nI5juE
v6oPQ/6u+kpUedMVeos7AMo9zWwxwRhAlIiOP9pDF82qSczACa1YaZOx+QI50aessi1vVjVN0RMk
UH9rG714eIfXNy0kgPtNUZDFJW6/OfO9Qcyl5VddwDB4SNng8FjI7k54ZtiWKqUPqVo0YI7Kigg0
FKtxQHwpMA5X65xR8hZw6Fwp+vgGDHLEWlyEyIw43ShSXWi0KhFOP/1yEkI6cV2Vtb4f+WsKaByw
GgKXG3mR2VCYzsO/beuwLv/o+PSgcEyBkDcBiQKCKc9YLhU3hUMg44LIPt0EnySqhZbFxT5w23Fe
PnDMCUihvCOViFvNDT8NDFTV8ivZ5/zPXQ/fB82EFgWIzJBsdBTdqyEOrq8oXHIboPS/Y+02mLN1
KC3vy7BWFteSyI6zxXsZtWNYOuMC0dt23VhAPBfZ4gNuyBicNnGIZEVdYYwc7dI4PP5sVtfz30ep
Tvkv5kTS0fh+BA81+rjnhHoW6EPpmxsu8CzCyZVW3A+KY1dC2S4buWVbXCQ/u1plf6nLjTPSQBP8
J5QT0J/LNk7RM0NB52+Oxm2wc59lvN+eiwJpyb1jU07D8/+cfbd2cQvBLxSKZPME7kos1uxtAf2b
B6JL0In+8jT6PQqzpLj+Bc+ZTTp+2MdaUHV+TdHQEiSPkpkuOUHQisJ29wn8S+O3HIbyG262LTB3
LSfDBS3PSa6WRJNIM40S4lXhn/CBA75zffNwGl9s69CS+obabu2iBSvr5bwcPY5tolZRjCQyu3/3
o82cZoAoOE10yghyNWuhGZ7p8ya5mPd9xs/0lKufvm/jo4L4roCPYUoWZvB8houxtTMvQI8CdWYA
/Vv40VIGaTVp1EvNAhw5itKD3FfmSGbAHSZLOqLVYUSs3h8KjRT0tSc3jx2fw96L56CdhTBtnqCP
GE84QkplkXefNCIE6daCXPTqPYyOJG4INIwSlVvV3foa47i9PCGE/YeQCwNTXIOLZtnMCSkdjt4k
GhIddRihpKJm85S5L9ayo/P0uJJDs1ZO4G7A7wNlidII1uIuOZ9sAyf1NlqqPtlMfbz6cGOLvAxb
397VrtdfSZkhcjua7bK/cgmYBzZPdUy7xN43eCsEcHLoVJqGSMtPZ4RGrDHwijBS03RLqQ860Jtp
75G9w+Z4UmBI9cH8MJZgnCYK5Q+2wUUYh/6vbs44MVIs9qgNuBqXWK25R769iBRN5K0qziPtIDGb
enuHISE4k+AUxaiUrZfL2akjlUmM3tJU4EyeEyGFMevFcSc4nQgCVm4RUgSqnAt1AAS/RJDKHe4z
TE+7Lf4Ts+NBbFDt5XJS0kg2bAxzK0iI/jtBboojPJBQ9v01/wxxVa9FrDf+D/+yEOodLs0B+9dD
oSTgVx75jUYObT1KZ1ncX8zq/X4bcyxfQ7+NgMiSdUQnjbI/J0QF5tTE+PQIjMuqCVzHSoDt+MVm
WD/S0vhsVukOpGbx2JpJSXpdbRqyQntnb76UmjjlTw5kjWPdRJXZevaDQC2vGZmCje0KUqiXrGFF
clDqCyIx+ptxrtFdzKPCkwI9ynYp0QFMiYPnOTvLQixttuvzxsRh8AQ9ow41mBkVwZpmMMdhYMj/
coyylMQbMUxwei9X788DQbgPu3RZQJZnrE8UvCnpkApdncF45ee8xY5Jw7LeYRbjvAa+UKkjXiNm
Gyx+9vH9ylWegjj3pWDalCwyeBhI0ZlM11WnhAbNzJNIg5eM3Vy2vjXrM0LOWrD3IUVPVBwkOwCm
F1/1I0D0G/4AX1ZY8YdqRT12Ar5T/AQhYQQZ+vRM1e1930w00zkqpFEhnULzvd/fWuT+8z43CxMt
c3TltG3pWTP3z6vLGWfoCUKyctIVTKy5JO7HXr3RFKMcGeYEWDm1ypWF8avodjTLutbozIRucQFx
MvpFIRnw2sEWu4gphNe9648m1miBPLbRZt+WsedWmJ84BJyMCLxcIkS9I45mMz6uf8ME/DzcYfNF
xEKmEskMnThFGNjGf+bYAVgttgFBF7HXneUN0A5OxjK40+hWJBlaQNsS7EUmhtdg8tYusx8eJ2Wr
1at4fK+W0on1OeLMCbDleBlzTPWWolaaMr20JCroQIDKxCMcgn7MwvJ18uVhFEX5K9eF9UhT6YAD
E6EhFXAZ60eUm5bjEQwkLfjDY2u0sN3Lq7EU/N1Uu9iyhwScix8yJ4YU0InPp1e44EfgEDwpFNHR
VIFpN5wfTrzJxvKK839TF86y9/jYNdUdMO77U+AZIzDb74xI5KR3J0RAobbBenlLJc7pUZdYsVwf
WyB4kaIXnDfn1Ek9MoM+RNbUIqOVVnaWb7xG5BxJjgDD6R+HQHIOiOTmonLXdiGsPi4LD3bw5F2p
6LGsPYdrGIsHKWjqfk/CgVrqEqlRWg/UbHEYd85ZpmcsfVafE0gA9t8511aeUovDYbcAhXVAF5PB
Cd/mIX6vQ2eqFOceFA6XxlPSgWVa2rg5LIwY8vbUW4BVY/oG/gRsW6JV+hgaGVT28boStwh6xgEK
4X3KKSnl5+sKa90wB1vG4natOodsGeYMO95zCB/wO0C1OSTnykPoH/ntSyA6V84gwam52zftrlCi
5B2yyl/Hn1EQYM4mmfE/HGzefRNqO59sB4Yk6pnqp5aW9P4u1roMKOUTu1C4JeuXIy52dhZ/ljt6
xViCS93JV1+tzkVUj7mdEUPYuALXHaiEzOaN8jxFRrO9ZUnAJkZIQOupSugXcN1TpQluzMzC+XTa
SVPqkZ91P3DFtdxFD0DCrS2fj45/FLatI8XBrcjfeWMTA+UKvE2bBGcTctOemvSLY8s4xly1Q/li
JYO2H37HDicc/WLAHY7SX4Pbac4tpc1rTwOVUMUawc71g0Lc3BTGLvW6w72mYWoRW8elsiCo0TW4
hvlVfa+RWBzUhYyqt4HFuRB9lK6BughQJFhy8GC8DogDDJSIONFsNkhhJguEBc9hQCjo5qSSaF1M
k/YCmHxKd4P1fqy6dlvr/pEPyYFBEOKs0loCVRLGN3a2m/8lSepgFv1fybgsnLnvaOcqJQGxUlQV
YKm5Zus07ZZjO+Lz9nbrdwSa0T2RhniRnxuVw7TEQZ8+zKiEWp2zYWoEEZar/Yegg5v1M140Dotz
6icfAjWMmRPoWDsnJnEhwyt3V4IMbKldtHSzRw8LSI7RCik4DVrBCDLgiU9zpS9EEFRu2LCltINs
GMXyb8+4Y0IkyHU7+uZT6Z3XZ9ouVP9vCZ9N/S05OCq1Z+ECeJZ8ikT14R47Rh5SIOAstpav6Oqr
ARd6G5ZW52LPCXzaWybHZMxS4nbtfDnLtCCyF9yjE2ckix/ZNrNM7B2qjMwrPtcZRW2ZP03lOWei
dAnqDYLYI9AUlY3UILtnYfeUZaoYbusXjBChEqfMoIcWSBaxXgW43FIp+ivX2F3JR8I0g27XBkEb
Xesk7ch/PnblyRkCMdO/YO/vnzOYMhXc8sP7wLNPvYpur8g35t/M/TFhnr9mehUrYuS5jXru6b7I
w/wSN180s5pXj0x9FPONe19sVf26EIHgZyYbaVndv/LHKRS5b2fuhp6EYCKCIi1m8bnCPkXUn/ss
zWysM8uvP6NjlBh9hT9Flf8RTA0/abMzcSzcWRvMS6MChK2/LiuBV6uHJnNw4oprO/bJb4Nu9G1c
9AutxyB23g6whadUD0xSY+JHPQNoDL7M/GlzITuo5SKu99omTZvPsU3kPyz/kjQwRMGWaiA7zslu
F6C8iehTuUElC136kwUiyXCuyolMSwLRMvXyc+H0+QT4bClQh/QtKZJOd8N63jFYKKsCr7HYdrBC
1n1uJxwnNb4CoeOaQjyjB0kF5fg0793sr5G0Q0XtvRCh+3RKJn/JclcKsh567HF3ZPGryPe5IvqL
+1C7G+gB9OAdREkric4tWbA6kXKR2zhExrpIxqVBn2Uyy1eyppLfQyYqrz7JUeRS8CG35UmmUHo+
EmMYlmwbAU8L+U1XIiEkaO8AgBuh8YSTX3I2Vgoe1QjQVwFL/Mug1IgkzgFSo3sGszBgnQv+6XPB
6w8sVYNhXh/E+Z6US22SZkFGp9PS+pldxmWDTxMAKB0g8xaMw5U9QidnLQoIpYDJCWHR08HngXNo
9AyT04HdWLBxhVVJpSKmLtDxcYvAcZ4SSgvW2SvQ0sPSevsQbUkuMnqZQNBdhlUCLnOv+s4i8QCc
5yfrg2MgxIVRmHdB6ITpMapX5BEJ59OP+9cUheoWJxMhwk7kY20mCpJcHCCpGGxjq2PqciIuhQ3T
aHsWczOWYa7DQW09BGFPwvLrTLp9xVhxPkVTD++Qb9GBCN7gmwv6PKFVylEOBV4XPrMB2Z7wIfS4
j+JSg/t8Du7fABJdt3XbPZx7YZNWXVFFNo1gD7usRM0zti8t+WJms1rbAYrm70qCapYkhyW6faWc
WMUw/wVyWlE2lHaEO0MwLpxvF/PSBaNZzqlxH8hURjLE3pJumVOPU9TJ729ilpOaryKdmxNajt18
/6B2CLU47w77p90EVjkhY3AMa3xX+mh7LKSUDcCn00JNhEKFIk2Tmp2lwcK4lGvg8642lo0zoAVr
B8g8RAC7XnBn+SijugbMv+iuhAI++Ns5cswEFDl6ewdVLeVugnZjYurHRIEAu7h/oigGUn8TBbhL
nzNtZSz5HxSIGnYc4Ek9hWmVUsKanhiN8VV9fszvkKcPDO1g0It7amZGKAMGT8x8mjyBCWK9osrX
aCEfJ3Wk8elWmX5sFzPIbZbrSPKAgN3590UqOrxDVArK7PdWzq+f5DRGlSzfGmv9q+61UPMIcujO
UMYENGQATs6eQ2hUwKxALCe7Wg5gk3OOpkH65e6cC8qc8NKPuD1/6ScTlJgyDGHl2LfTZ47cy2tO
yl4mh+NQO6Rhp2vNHh/rUKqWZCvOHxeTiTl66+OXFhbir0o+OvQBzYNlSURuLnlRfNWYALpfysG+
TQsXfBHWFSwePpmaeZenj5ztIVCI7WcH4h9Xk1tbyf4eMc/bN0XmKV4Nnr4JWTYOdq1K6RmCEYlM
YtoAFips3GBQUTudf9MsFfcg5Vk3DJIe8ocXi2vhkXNHb5vX9dtfz80iaFhfcIZsd6JGDr1viU/s
emrmi496kKPSIeMelih1/ak8QR/Uk2tFyulxiU9w35jUKv6XDQkVs3nWW5it1FM7kG1b01PQqkr/
oQ1ggZJc4m0tkgbMPAPKNyAXn8MD6XGUYe7mNByOt7OIpaAHlWNoE9+oHmW5AiVL5vZNQbQZx1v/
WTPhYLT+UPUm+XiA8h44hmdNrKldTfTuVoAa2OYfFjyEaVh9rUeD3O93PJXhz9zk1injff9l20w+
4Szs1JfV4pcfrztW/Q5NELtE2MzQc5qlz8OpF43oG4EsINvW1WebG2JUCFotLv3wQ47vnxWeNiEk
+OUy4t3hrl/bQyde1QyPk8ubYA2eSOIBlbFLEU1WEP7vBb6x/RFp8kc+kuVp0QiJNYQvSqNUE/k2
7AajudrBZpjC+OcA2Dc+j6P/FbZ3Vgx+G28FLe2pjjd58ygiLsN1wmvPxL0ZnlxB3HmjnMrsyG1L
YoGOPRLcd4wfcEzdQoMEdsG4/1AsihnPgu4QnsFJqguSeTom1QGSSYn94LTJWne0VJk2gHudOsUe
zgBT7a1bDocMtnSGOqda/RBULnrY57WXCIJPC3RBkdAVDNDa+nLBTi9L4u/0rdGDN0loCIYiEJKz
MswEZPb9ZekkeaMa1kogZdOxfu+hoTM/TV1jtGcvmOBAmVoFfkEScMF8xqpklG0kT8+CS0T7oUmM
i53knMDosJDaP2MVq4BAFEEEk3f1JhZ+GP9iYKPlGwJGxY26Lo+SuI7lDfXC6AeYiFQxPH+pJG9q
EiuwOIQNCvplxl8PqvGySZalD0Zgb0eoJ05zrlyBqKvKGY3gGO1g8uD26M7+uNUrnTyomlFBGw6q
iCxdKGKm2oy2pM6/ic4OiMMV/Gd50fnCTtIaQIGMjiVUjaCC3gYn5B2J0o6KHLwleQseV0stt+a4
5lw7eSuh0a1/JenKNikbMlg3OPpR0ZezxIMj0n/1YC9lqFWR1/QC8Xk6lbMJaNonJ6vyoNt8yHe9
p4r/7g2KsUVmoSv5PetfLW76rB5EOzi5g0H8Alucmo9Szgnq5sGlGzsV4FTTpDUhpR9zc54Kk1Ei
01rqNyiyreq3Hozv9bOgH2l0LSBKxscOS0p4Oqbh/08KUDUkC8bwz8dn/Vo9Mhe3/6IeQvvhK27/
wfyRRO8P/IZcKIyG21kQj87EE3zINlogNoGnZYQ6SwLt7EghZ3wFgqF2lU33JWdQ/xh0k+lihy8y
VP5/N99HDQwnypVl0SFgxA0ZdI2yR4zqqBxVIHUYjnx0yjVUF82CJUkpWenFPToH0Y9kB1LoM/HN
n3IeNdz9OVW80wPi/4TsbJanUO7UOhfSIqPmbIaUgvAhgYh13C46eKaZk+VkzKyvbw4cB5FTtUbT
ycJIofTuyGamks96QUoZ5gpsJNgPP7QQK2N+kEWmjUoVgYPBokh2p03p0847YJm3INvHV9tuah92
02vXjlp4BujNW+/46FcR2LclRFOdJ/fi7ri/9+HzThH0yYmpU22xxoktGQz6MCDm+qf0Ro074nMY
GcfHjTAW3hAG+/0XHCOj8BnrikgVF/FIAAz2M/MnlI3kMs/oRPQAueaqvNk2Ya9bd16MYppaQPcL
ubtbHBLsjCigzx1vs3wrKfiBkHO8y/ea383+MxCD1a7d0vhzsirf4eQ1H5kMlmLEo7gug9e9L/7V
B8uuYdI1vC35cS6C0XFbTrkhae18dhD9COm1Vk/buKMzYKghsiRAlvVaTkJBJxOzm1ZjTgDyP2xZ
lq7sYHCu89VnS3pzATpWFWkTp/U8zcT1w+S8otq/PmBqvVz9rSF3ycMsCLr3R6TbGKjK6ywA6yqD
mmRRGQ2kifTbkel2t4Uv8UIVgAD0clP8NedPix84TzzR+y23u9Kf6yZ+utUNeLHMUYbBiQQQi+YJ
yPrn84WYuKRcqTpa8oTbigvzxLgKJY+ry/ZUM2Cly98wi73ng0uTt8mngc5XATHapr6lbsE7uKzv
yLUPV8qgV6dfOf9h7ZRT2bzceRbFqk/pqtxZYaSjJu7kYt8OuIJzKSs5/8KD/3TCTNIj3nTiq7hO
I0qr9rFcHGxMTDyKewDPx6pOooffSCemhSGsqapl/zlBL2hZBMK1b4Rqbu416dS5YDL1mxXtfrgo
A4yAvIH86YLaFsWAVmsTKvLVvH0KKmMkpWtDR/kow1/4f5v1hfB4VFJoYc+y0DdyYw6o0Oo66bt+
VdoUXKPnw9qSwaC7DEh1C8+6IolH6sA14cPaN8ZkS/YxyB7vRermH76gJ86soQcqEb2bx4/1O5Q1
2W+29+HDilAwJK9E6mCnpgOzyBXwtIUnzjMrR44SHsrqAXbnIYZUPLX6sKJTFNW8Z9od7hY4LJ7J
1HtH+Lih5vGzM6zMcieSGyUb0ZOQEeWkXtj9Mx7q+90KAU1Jmv5BJLB8yr13aWU6QEkVtJxlmLqm
0cDU20rfoJu9NedZdZHD/NrPw/prLoNyhNZdnmbrRF+40AVQ1vbWR7WolChHqKBdjZvA9/Q3i9R2
J8xEwcKsk+vE9GxFOJ7JGsVd7Ju/hYEg8xwQvrofPdUdits/AlsRwgiNC56jBwYULv8EKgorEaIU
Bi4qXpbkZxLD0LCPksK1uv3dFz5B0kk4LYq1wgj2UPHVL7KkghR+3YQohZq4hweOJ+OGxSwHIwa+
we2v198zlLBLaEAbfJ2KCPUKI7pPOUb2dR91mB2d6yWLILHEFNofEZL/eyJxWVujUXNv6V7N3zRw
Kph7ram5Tzg7kw+1Fl3EPfHf/S/Ri+Jq/gjV8F8WFMzVlL6nOKcw3+KBbzl0x+SoXz9SI7TFieP4
OhAhD16FM/p1wMQh6HJi1Qkn/JPJYb8ZDLJqXhhoOYVCWt2yuvgAYortd9zccRG6s/U2mPHtwGOy
B39biDJcVzCtWes62hOOy5+WMp5vjYFBzvPWsLMLuMZkVQV9g1JG28tUQoM/9S3WyNpFA+WLYrhr
40StNJwM99JEywXqbFXAPjpfCCBi086LvpUYsLgMJizW8EDUwf5mDwk2vqQjZyu1L4/L0Ufwdy/t
2O4UQW49VFIdpCpN/miSeghouh/Cs1aE1BN9ZameoSAR+As4+kZddZQ5CB7FT4CeD3IDlmVGZJeb
zQG9LaRg/ex5kQcTGhPD0U5UC7NIcJ0cxVPcgdtRLjLk+z8BrN00JYh3QPx/Ja01aqnQYLk/9Ya9
cy44G3cZFqtsyV4bth156+H4YbQHq3FCIqJTKApdUhaA6E0bQRAA4yNSlXF4TiH8VMi7UufRXURi
uRhBqU5fQMjH4rCQbYIwglmUc6wPvEHDrNSCSIsfINv1aX0WdB4Qj4HpDb8LVvMcwax1hurXFs3t
5Oukd+HzSWmMS3E9Cd1T1DyNwkY9e4vWqffFLA98Lxe2xw0/Sr5F2g4XNA1tcipBZ0xYY4fC9gmE
IjHmRXihfx0I7tizxAUWCBXWUKX8M9so3UEqitIXMEoacBI1pm/i4q1e/NU8vK5Twto5QPLmFyMp
3r9r+v0cpigN500y8JIZPwzRCGvcFUiYk+cz65m/nO2hgTVJkURBTeBHnq5f281ksup0rY5ZX6KO
kyspXqjBFVS/extDFbSCAcj2AJd9m0jVbemtlBAtK7U97d8UaoHCPS/Go8e41m1/Vi4heF1rSMXB
OJKuLzST2DYGHv48dvSeLtQZSwAyCsCugR+oTxg2QCTePzn3efrwJoSkmz79WjuGl2/chWcDsK/Q
EsNadkW8sLssDNMXNBxPv1njF/WZb5CeDxOXSveYMn/TBvKu2zgAIJNcHreFYFo+x+9zfSKO2aYp
D9WoNvUXFEb0orgJuzElItnk0IKYhDABK73gEQf/1OHIK/l54TLm56F0ExZp0fBc/x5BNSOxElC7
ZwKJW6HsVwk6C7p3UN1/4Agg1OOMob7mx6o4sciSVoYgiRdaLIEJhQRhy5avqYtPUPmbKN0tMKp7
9PVorXrMyI64HhbHKVLRoF0A3ZKMBvivm278pm6K2of1Hfru4cLbn6DCTylQg5ABMgMHgo4mWd3O
usIPHI5KfmduxH/3IxcvAYByGQcn5XB4QL+yDEKSLlvtwVt4hm5MpjPyi1BuTxR1OHQmCANJWVa7
EykqQaXY+L0h4kkFy4Bbiadf1QWzb+Yx8YkmiYbPncnQ8BsTCKV4QWtqhYH2EgZFaKznXU/TpnV9
VcD5O21eeygUFpbdPw44DmlW6g+W5zx0QDXgouf5wI6Fo3TupRHskfO3E8/yP1tKSBoXIKgYPxXb
7j0ON8XoWP2uZl0BTSlmzrrdHA4mj7qk+Lht0srPl89I0X0CJS3flLi/rhGNywtj2kpco7UqOaYz
jxjIvRH2ijSohXY/EXRpNPaV8cutXH9JDRyOFFOE1pZCyat4UDeuaYngX0SgIWVgVjd9LClOwYPC
uLtYXoOWDPrrsuulB1Q1h4Xsv7HuWYyCKP1vWc4wfiqxF/dcfcwfsFV38HaFbsz+aHdfVP3Sjzqz
zQfqJKusIOBTkNS0GgLHidruB6Ut/c0xmaebaqhmdIpku+/ERZClGxyW0G3FtyUKu/lU3svLwUyj
7kV/YZlu1R8A2crSFlt1drsswWWZbHK2Rksym2PQxid38ULfpkwGdCPOReq9cRN1PWONODEuTojX
CrVsYRguZdVVHpden3jpfFicB8D1HtPVTJpWXKoiZDQuHaRciewRn6yBpEyAu3qbsghm3mcXrgV1
/1mCyoBnkq906mpQQ6T6RHyxVRxV+w4y/58YytKUo/5/+z02y9lTGFI8p8G3RJdHvg6dJtAdaGaI
eRF0aNxM1bm6NfI/Gy+43VCcB54L9NuHkIaJsCw0vsaQbZ/YJtaNyxVYu4WEXjzbiDlAiFpKQImf
31tuAjMuwBn3J9xRodME+R1OjHRXyeg2YEUDp3y97OFB8PrExm00HkmoKfwgJHCsWSjKlSO2UHhe
DQeHhenWOTpdVsgiRAqd4+PYvEriL0myQodMV5qBrUU5kQHxiqX5rfG8enBjLEna7nxMX9kBx9PA
mUqmAMD35O24gT6iRb5cgBzIrmav5w4DurB5PNRD39clYAPbsZaaX/yVUy2syklbYP9HWQ+FWz4S
Jf1RS9bgu9czBns336tqaTdlqzTo7US+vaOnfk2h3VKs/yR9Hpk5pvikDzkw73q7mCQ5RkxeT59w
XBaFu6dX7tz9ddQlVpFD+5POIlVd8Ola+rLxVL1joL1DSnYt92mRg5HWPsoDTiPljyGA3ftzL9+Y
3rIIKUsyrWvy5EYoZ30bnWg4TmQ4Ds9P7cMnLpBus2VEUq+64zn7DV0qJBGsF3lmLJCYWqZoZWF5
sMFSGCx1WScKyCh4ObfSMCV5sNeMwz7dWcsmtMp2QtO/wIQGXsR4Bi7u1RFAWWF7xy31qe/3n0K+
GKB3zZO5MRkON7lK3ErAwBJXt0XDbomHtJfC7hkOdbrU9fweJRLkzVLYELsPEx07kvAWb9Gb/UDU
pvztgMdMCzBzrHCbJtQAxJC/+G506xEPAALqAFCi9grjHSJiGdECFcH73rtjTZ0F89VdfRaUZ9kk
Ia33ZcIZut51Vuow/311K9EPKITE6b6fYWZ5P5VU9wGzBtAWHqnh/6w9eRHxTZycSgBqTUoEymdM
WJOW/MilbNSmx+tGubAskjhja1n4x3gA5xzVl2fMdKsuO6DZwPlefIYtgJHKDmIZ7bysglbTIgUF
WZdqVOzPeApvJOpiNOh285UB4EeeiVWnjxWAwYNYj82VKyYkxtytjNwJa4f9zipD1pfdTWuCiRDd
J9EG0/lsVYtEuaoYpbbqAFv7ArrYI9w40JiIA2but9R+IXJ6BgEtACv9S9dUcXCtC5DIZlqNOMLF
W6S+VgV4XwjIQdqXGB0Dqiv7iQi+Gz28neZMM0kcu/CyS5XYVkAYMBH/39JqIu8WDgRtyOIvZFEe
NFPUxNRBa0D0w/nF10DKgL3ubnynLJxCU3ymsmjZDLB0F9Ds2ZhiGI0avGMsQxjJnfEss0Lrytqt
OEM3fgDwvo46ijjf8wQBevS/lwIj1FIQD0gFj9c6E7o+OuJEYSktgG4DlqDYvDpb3cEZYJot5PMk
gkCVngbSNWELJp0g5RPmhAkDZYmMUEuRxJk2Zwev9HjJ/sfN03rGdvYKVPohiXZRTg9aM0z/+IiI
SgLDkvoHyNzXXaWz92KMUgHeIZLEQYvoU5mcSDYVRqsVB/z+tn5QUwICwx2It+COCnfltlM9FehV
7oSp2va2RfvJtZaf1owTwTSKXxOX3C+mBYGCs1zYrDuEbAUhy1m7/dOdnClikGqx40e0l4CtkAWt
4f+YTEyDY0ZMzmqnOpK2GondIhDPuUeezaJuYyUo7mzUnxaod1SVBwvrkM/5E1GyJTrtiMV2oqSc
Irfg5BoUcUsB08jhCOMadH6GUsRz8QR8SFrAe46D8t9TLDoRsioKcQ9jBLQcSiUfmhNv3wdedQiB
grq9smFRKzLn/fSLhuR0FK0SCN5a7yb+63fAMf5sPVUxNkNcfO/2dRLPt7v/hApFy3fFqxIH97ve
fbFCJe1GDzm8e67U8lWF1OG69Kv0HVVvL7RvOWEwvJRxUEBfED+m5t+2Mz+5prbzzA7GfhCEJfd9
3D0GYtMJIVf5PqHn4d6idr+tQKuXRkWu5OBs4EHOdBCwMJsIbvnLnXnXkDeVDOx2FOOS6ZVrZl74
4tn1SkkJTCH6mmvOdKG3LM6BFNjczS3hSXKKl+EPDDCPRDSbJlNmmLXfsYSvxM+Q1C9+Jx92Yuh6
AmI+qoWYQ2uABLl4USxPFl/TWdx2c3SRqc0zpX8fyHi1lXQEjJZfRMPxSY7jynjBfLYS1RZKUtky
+h/Tot/R5ZS++Ja9tQqtStGA+1hDUabVAd0CXvw1IbmItyWSwjSVTYPIOMbaDLLkpc6gjyhGM1Vb
MDmy9sYXG8eJ7IKWJkgstWFrb2QDEYgw/Q7UhwJdqzpeH4T6o+8e+CMzLZ586xmTydT16JFyoqni
+TA4uS/mrD4zlpbg9H6gVDFFiWUbeQt86qlRsiI1X65VQLpf/kzHtF9x7bKnKktAmoCYYkknNLVp
yXSP5P34aMkVydvXXKnTQlG0uJc3ecU4DA1PebBOtBOtuQeOhs9wPDPhy8bg/TmFXmiY/azTkT6G
O8zOuSE1B8lWSkko1PHvPNYzuZQaOGgdKEu1TJpUwMstrAPCth6YFs8fzwDvImc7QO0k3okPfnac
62kmmFJSG3WsKbjI/kNleTL/KI2IhAkCkPeJmPcHoYhHgFLMduwOCNHV96ABNaPFmZxIJEdGTIPI
7yaSY1uK8NSs4eyPRaLDV8icgaDQJz+rVN9qRcoIh8EVmMNrlv990sRASGZNalgjY5c8ypNyjCuY
gINCQL7jM0AJ6MlixW8UslF8kTGLrp+VsuSz7sOGFU1HWNu32+Q6eHZaLr4mwMDQnbhaLT53m4YA
HOf4uqhaC4ruiSa2o/cqHBZ/7QzFV7o2elnA1RURVKrcGH95REhTyfiNLBPGBUZg2aevfAFTzh7J
M09h+xsgUiebGty2fg+jdvv5Q+p5V1o631QmKCFf5UejFg6BgmyITsb3MM5hRy+CftOCq4/IJ7H7
a9KLIig+8sEPOjCYyarI+eUvPxBgL11dMETZyxk4k2aw6z7is7oZpwFiLfnML+LkVJiMXYRE2Wxb
8goFdp4uOpmyMgd4ubtNA9UDN7T8dI7KYMIqBXxBGG2Hyev24yX4z79aTb1/OS+QZC/7Y8FDx6Q5
bqAERCKsA3QxqlbtPj8iEiO66GSpfg+fZJ82r5he4A6oJHLmq3X0xL/lCASu6bS4HdP45U+w53OS
MkzwUwL7v5FigOfSGPf10pOBEH+Sa794LMmt/9X/6Jllas4JIVeXpQwlmPWkObHn5JmWW2PIo6VU
Xex++edgXZs/c+gozKP3j4mBOqnnI4dVwFI76vfXrYQtyVajPQicwvg0A+qoY7NpOVFRvioTwDRo
MeJKlh4cFr2OaUAwwSabG7GqTxfhpH/3nysf/UikOPAfeECFrWMQ5trxgVR+Tmaj0WVg09tirpUE
NpnlRG9XL7lyyaoP59S6gbsh489+l0iYJ5AgqIPTITHtiVudJ2HnICsJqGcUVAxcx6qfDnxTe2QI
VbmUxhs75CwsbppV0BfyCtp54A5SM5Buw1utqUqVITBLc6tNYFRq+2JTC7p1ze0kVqdhcMya/hUr
54ELJbOfmlmMODcArakrVqAEmqqQoAh06L68+ZJdlpMJ+f8NfBEkUPtvjz6bA8KNu58n4yBCcuiI
QiXgwCbeL/HCwYOmt1r/gKuLlx84Ni1MiysMNbPFJbEBF0/rmlXsU6N8SDECa438VH2s+7n3VVAR
YL1XIxmsmAYDOB7kBCw1tuKT+47TnH5oqUOgIGSXMZhmxWSLXNQs5C6hu+XTP74qGjlbNvL2vBt2
HBrL3KX61bTa9Rb75Mxm26qOXM2yeJDCO071tYw9oNkUVBBh4rg+h1JUpllfH9xKZShUCgeFWlEm
eeNvbkjf4ApdZIB/GX4CtMOdsF8UoTaotFMv3wQAMpgMG5zNNeKBy2WS0MQCWyoB8zZcMpxvZ180
w2hb+1r2V0HTvmvWehN2A/qiBBzh1BRihKcVsYaItIQh5w0sFJZnZa4BZw3kQduZ8qRGtHO0dmec
y7kFVEwCXE7C58zrwxck47t0nEAbfKjQxWOsTYi2oDZKaD1vni0vbDR+CGUC13jzhMTD5B0Bvb9Y
ItjqcRoTgP7kwtVA80ifPhOAd3vheifkAB6tZgB5w5ip4iBuf14rUeMl6s/Ru6q9uVppzExPq7EM
p5XJT3Z4AsEByeNJhbu5cvpYeK2c2iCTS2iRqWL5UFlD7tf7yxewhumiNNqboRSyUo3WpIZGbKvv
+L2MgrdEomS190wilb8+ScoONLIyPAfIhJ1I/2uDmB+I94rv+j5KpUKTx4FH5GjHba0aRR204ftg
mN83OtdEDP67npS6W1WGbzMlh5MJ8VKiZE+9m/q5pge2GPG7cwRrlaJUw/+1A6vzaei2KnZDMw/C
TzOicM5P4rgCGqyaF1dRVGkLjE/Ni4FkSV2/bsxKkSrLTAoVwiGdDLVRIQocz9PZfQ1CcEEZpjCw
c+rri//uWYCKLn7nhkNYvaAqZhte/9BgzKz0Q7IgKWrm+sxzIwWNy66RrjOZcHd1UPoBPgCoD379
Z+i6eXBVZHh/fu4qwPmCNcJP5/sOqus8HkPMZVfzqJEDBxvZoq/I99KanaP+nWbITsHHcQnw8rtE
pWFlSgzlUmUJiHy3+afCzm4I43Qk1aTDd7rL1vlKRUZUleG3UqTepH2LgPQd9MH7dgtGNAyeds1W
5j0p/vTWxNUf0WQOEstkvZpk+MmPKJUvft8EnZCIS1CT/0T+hCFvi4sAoqUtsbYXYxBhH+0tTcJ5
824YPjIpEaXs4eQoDbk4KaImzKnRZwnhc4d/Mo47KTXm1HXpJThr6pTOdW/ojK2N8ta6ijG8z3dK
J7TQlVkxBFR/A0PPM5ez+LuV+zV6HR6MzYSMDudl/iDVjrAQiduYHZO6yaHXwOjzbe53rTKvuUUJ
4uqJppZzCBcHjoGWGuC4L/52J0CDefXpGD985Aa8CMNRg5dOv6GYXX/FC/utTZwN9t3mhHILTySy
UX9/oqpgi4EDmm+6CI8haRXK7No7EusUxRVRSNGMmW2emA+b70Os9HmcmpUZx/y5XEqsbuvQLtwJ
k86tXHpelvBbzCFmqGaD8wca5M76vJuot5HfJyNI2//H89OlAOVLdGc6/4Xh4mjhq0J4oGvJHo1N
K1KBwke4Bqp+QAEKCms8r4ARD7e9B+1iyxlfTZ83DbyGIgXPFSOjxzjvgzRS7CKzC7UEoBGTyuqR
atXWAY63dFY67B1PYwDsm3U22dm84/N0qxlbvAxkWfH5yxJEUvSgmY8zwR+HWkNXke08FBcROPv1
bzoBqWNuxyxW6p6bLeCouGxn6KZF9T9kxjmSkYSkS0pSWWfUW/iYK/N7PIhmFZ+DJG8efsovImOO
p+JO4N0KttgsW8jwu8pD+RZsCKKEDdZFnOKoPzBpGjs+GHnjM0yhTJQAxRAH+ceSxNKkvcU7l5+v
E/aITfv/K/zqmoA2lWOh3RD3l5vtFtTVwtcf9YAcVkmJT3oz5kYQBbkeKtBpg4Uit/U6UCVxWIde
Go2mlCY4BavS/FSmDPaVq79Z4TkZP5UdN6ocboCzHLhqm3KI1i3m6HBs+8tSpfQugU9RLFIAM/9S
G9jpJ/Q1htXIF1NSX3nhQw100P/7HbtcTblJaQSFJFtho7zuzZIsYc7zwc4fUNQZfvAeZv76cwDy
HNOA5fzYRoBeLGWfKYmx5/KJXbFzRKDTWG1QeTpIncNAGwYwjk5CjgImOrwxqIWcPL4MtMBMa5OD
3LGE+DqG2Tvzwz8+oYAlb3DmcCAQ6zhKmLOmqktmerah+topToYj02Q/SM7+ybb4/Pm8m456BDRK
hiL7tIslS2Na28x+tNv6oboeNH0y3wNx7Etk5+5G2VIFYSN89Zgz4ETmYNMz9q/LkhhhqtU1Fzj/
I8giVzARfkOlu3ZstT/O/0sGkWRkk+dCE52oCK8DhfRNBLr+35wBH7k0LC9tO5M8QoMn8NKaWrfO
l9hf2ixq7giUPveZvOWnez+hUd2pBcblGcj3Nit2Q/Afp/8jZzC2I6Y4R1jOyQT7TuOJ/WnNc6Cd
nr6Oi7L3pqabJIO7DG6Dxs8Iw6dcsTE/I4hBzKF4HDraDns3ElWNHQ6hVl/L5Vf7cdouofmszjwE
XxVOwZVlc7NWon6j1cg4gkOvwRpXrmBEKdLr1wxUVx0cGkZG1qCZDVHMo9nWyX6iD60IjXsZW6P+
3nCtGxa7zcsV5jXZ8R99es4rEOLCH0dpzkkRC1Q2ZZ0JnM9s2tiFQc/PjBDSp4Dn5wUrEoFT7bHR
Xu9X8LcwlZoP4iOxTl8gcg3SFx3UF90ewkekivMQrG9Eo1yGJ1/GgzqLkN+SIookFcfHmLRTtnEI
iYuUS5wYExpafzEjG0mSlc579vMdIgrEpFryLyjFE101MfF3OVPJgOAS4CKGfZDPlR1cYlBTtnKU
eLlBQMlPBbJilxqRumACeW5xNPONwJcIA90c5JKFibMryX43tDR60y74D7vP5Bf3pSjulu1tNHEq
pCevHxfP/gSCwgIPGmKKPl9zN+KOYYuJJBUKccBvJDNsAki6ZvBoY2+8CJHD9fCAat8ZZOLqCf0r
7zE3am0XY5NzNavrv3sbYJRuNxS3FCV6E3VAl/iZ8IPm3LdBA392/qUsZagJCQ0AkN5Jr5eFjCKq
kCJIvZbsfLx7lggvOWfi9WMxcIehYV4Fdykm10rfYTvOcyDX7mtO5+pJLToI84MNSDC2wR7qzDGm
k0JKy6lN5WulYZ68wgn9j6MNQlgGj2FxroardzGqA6KtldohAIzxcjLPa5I2yjK9ftM8x+CWb9W8
GnX6mTfbH78DjoeqqcjCMPVshTxuYF7gUhGlHfprOk6bGvOfeXzWsQ6rIfRffVA0X05g2lkUjQ5J
Iu7urr+I4QwfBL2HqFV9cJOLXL6fTKFs85aXLYGGyxeaU5ad1vk1Geh/wkhuQsI8Uzd87qoNERie
7KrHEVDHeM/8YWeCUZsJdvPJh60nbye4uElhF1HGzWKZwQey6PTNeu5byp22EJYII9fvPMJivqMX
a7adDcKsja5dAZzJ9+eqC+F9WxYG2Pk+z4v+zyzDxp17dDgjTXIX/4VyGKpaI8KhZkisURBV0KLG
Dyv4EN1b17i1t1cUArWfA5+5lcPusda5FwGsc+Z5un/V06U+Th616hjxyVEX3TLyzeEBYelr5mQK
ACsEx0rD8D6FLviCnw+XTU3njEWAR6ckBHo3sdLnQle4rCePwUXeQDzJzhPuPQdBMiVnVOLAn0Rs
/zmUpqRHD5NXaQRfUVoDDDgIR9v8KHmWFZ5xyXq2rkx067m2FPBIm3dJY/bBdO6xa3HsyhTAyPpz
vmMaiUNeP5BDbawCFqE3M8+usGx0hjhwxbAG4cSHh6cCcp2TxZ5SYhQhzFe7UEda6teFtTcAYlyf
svNbXU5xHD9cQSTyQUgZiQqTp6ZUE/Fixo3DLDMXFXx6K0cBFIMKgHKBLYrZ1VqvYbJJvN5EbS26
f4i6L+Upy2RDHPvo7DmHH7h4Kb7I4Fn3f4YrvsBHvrpHVG/N7VpkFMbXZpAddppurrz8cBewZ4S0
auKFVRhvTvAHiaMJM+b8kIblNECIpyF82qWOv4iKplTf9/8/1zVbLO9l5zBlAfb23hh+Bb8hCdIQ
XbOlwlrWtvjhxgWlrphC78sqDxGaSxC4pp863gwAA/yKJTdxsqdzwKUKHnDRdO8p59wKHLfciE2i
gEecWhhm9GTurIRlFVljh137AGb2bKgn3K9SlMdiGR/P05ohsA31C/Eh0SL2l0CkFlQNO4wqpS/v
/ULol4egti86KA+zkBNwGGVSk3yXb3swj8HV0lknXX85mpfh3J/yDI8I1lu4koZmlAdO0KSLF3Gk
rST2jqIRA4C30XrLDDJzhL+j9UYOYDqs7VG4pKTtJqgt+RVA+4iHh86AwU4my1YGkZEEJG3wXIKd
uzbMYX0m7SajjbnGkwe/W1ERUCcSfzuBgA0AZbKXJpCfneFGlKlYCCmBO1mo+ojc4ObGMHnzcYTB
PBeVdsC0yBzEflhIDsF3dY54NWHeYEtxic0de+MktqUcLI7giawFrbBL+f95jB9y2ewdq8cRAW/4
sN+cQWmMCYme+nuIR+tpDdtmDpE3M7ffADHY/UM88DN2M2punK7OIaC6BYmfscEeVWfzqBjDFvJ1
BteioX5WAyPJo1Avujf77kgaBbxPTOvi/AvPSaCJGzD1e7Tnn/AeziTTLWeSiTuiftYaMnmq/jj6
MI52qsCY7i5V8GDyfhcNM+mHCM/mmtsNS6EE3UYJTlAG5za1lZiJFYcm0N3zVwqGgm0m8/funTy2
k5GT2JQH3lteXZp+kh0oRvgES3W/vwvgMG3F3gYTh74c8sRBv3PMgsY4zgLtw8tRI4G7GGeJJNjS
cJsfeylTgmj4KNnvxS0r/nFDn8eKWiJx+wwNWAQhx37rBEEhoBodiMGksufR+gb3uRmChLX4CTXQ
WQi78TIModDbf2Ls77fQ7O8YiBB8fRgu/f0w6pRR3wLUDLMTpXm49iBRvsPSqVPNbvgKAbYHuRMN
jXU+M4pmpXl+6lci69tzm2ESHgOeDWb3zs64BsDsKf8YjlX3X52DEvTqcDj2/8IgYBB2Pl1JR+5a
n/JLAOIJXOpVj27ZDUSuCIcbmP9XspiP2hHkMl9hBQbhBWIPeYJDoaQoFGkhNaYKPlIdZDdHJPs+
vTGVVX6XRMVq/OQjbmY/fq6ooxiiD6qflZQk8wlNX/cctjYgcc8AoXeRg2glFI02Uu32uFKG8twJ
1LHDsDowdVs8yoJMIf/0ZElTn4PgqU/MG8wqdsXGHFisQYub89lY/P/eSkTx7K3fAuIJhQJ77AnK
OaLK/W97ckogsLlqHCjUTaQLF/3mWUfe9jFxuuyA/ICj8sZQfazjkh6+ik8p1Z+xVJDg7HIbPtSS
y/zhVxzhjQmuk36wWx2QP+AYtTuJvp+ucKzHKjk7QhJ6vticUr5txjvbLGghzObTklFMSFPMzcVw
CrIuFRCPW8DIM89Ou+nfrFmkaiqmtI5UOxYa7ixkahJ0fcaKk4u+J54mMUKlLGg4wLSAQ647wy/K
gLzR9duKyK6x6MYZ3CEf9rZKn5+QJykR00MDLIiKMHz9u1p2P+XmEWIuvV/Kxo0u2RECc9LCsliH
lG4gikc3Vc3A1Z3dFXlK+hpQJD6fiHmpCKxbhq+6uq7Hdw1+t0Aj23xaYr1r/OU27d1GE7cQrYic
bM2yLagakE7GzN/bsigrYKunpUkTf0SS/mLrvtTX7SkL53gT3932DSlFg/E1OjZ0GdGmmoWi1J62
0zlPLbH0iSWW2hHVuEpXHD/olAJ+IodZ4wCwkoOiwT6iBhzCMJ1RSbd18z3Vzy67zMlH/jrdVvnn
DNrqTVQ/j1LDiUe0JWRKKdZ17XLteaBBfIWLMOFGXjryV5HlgnLJnwZecCWacIowSN5bg+q7POAU
mW+7JBf+h6p+h48A9pgu6xhRIPJXZDq/J9mI8Kda8bzlkGFKNpkuiOoRsG4SfmkQY3hcaicylaYQ
hnqaii6ayLMUlb9siHceE6AK8UG0rlcszmZcxFNVhlKbpVWE900qR+B6WULVquP+9/FSolwxVbrI
HG51UKenpxNIicibG/SlgIn1pAXUbnSHZ++JOdxVLbGSY0qTS/nRQCmFsMGgUoanKulehyINH4Wx
4MBUXGrXmoJSqAtjPKYd4qS/GBwaHtqDvPJDIT99cxpdlocbQjrvd53ybjy9N46sgHAfqUxDujv5
qGA1iObmYX6dIi2fQcWHKVEhx1h5YpaUGc2gLGMBNk5X9z+DoxcOo9eXmGbTjg18oNf+GvHclkag
E9RYqoajwo+H2YY+5ZrNfamuEm4s6t4QGHbCN9RBRGHJ1+CuPNO8q9BEG036rqM0q3fpcIDwXhp8
ko4NJookTs0lFdsP5zP+tlN1vmjJRG0X92xMLOYJ9O59MZwaDGnF9qbDyGQJk35MIqkU99jwwGsH
pMt/SqvqrBNka3wr+GblVpwW0w40JJ5dQDu3V0lM2WK8tw4/cDjSoORRcmnHI0523/durcp1lQxS
VBkX0LXU2GfvgrLgW7Aeicww6nXhduN9OwQgn010prFFHc2D+tn7zsreZjOTPGw6h+aqZtXRWBAF
ZQoQR6vW3r6gjeKdGgK0BzKfaVSNDRClW3Mr5hqIMog6q4LdUXe9sSMIrdrVWZj1mtvKy8gI7C2S
MEYE4dWXB+XNCMf8PxOOPd1sajbLI+jrrhxc81NAsZWxcbwdHc+5hQFVC1kZ00aLGZXiYZ5VBM2R
zHRb3hT8rff2rhgPY01RJ/09nuIUamrWdrnddpIK6EnH+xiMfySba2IH1qzom8N8fSWgxy7onO1j
UZ7CNqiiZILQr4SQui5XeOnK6JecBEfHC6IN+OAELbKH084crjtGVhOkBDghgD7InPRXvir200Ff
T99FyZc1iYHvePWXP8NEeO1UrIYTPIJrAGpPSteov+bS8UyFON1s+X5JXPxoQ3kplAI9rgprX6Y+
U6xFj2OE72OwUpLu4QGuMCUszVq1k90YX9TTDOvbsT/JQF/EwiO3n1p+5x2NvQFH4qMnpPd4lhpP
AlHEoI5zMLHdMT4yevedKmmIR4qxzBSJ5zBNGkPWI3p9MwXDUUJLAN4cnZTpZVKwT7X4ENT8AlWC
pwYDKE3O4LcZ7oicRZiQpcRZwsrEGg8Yrzysq7/YA/xu2QGx4DZZAo2my9vCJyf6WqO5SiYZ/Rkj
14g3ppcSFrwulTS1ZkVC3VEa5I6VNVVXJSXpYc4Mrf4mPTiOF8iM+f+cWbHrGDlEhu/RljHNwuS7
BZHJiNe6tXVL/BWvSXmyTq4K/n6nq7mgKNtsPVIqTPR67IVCTmK3UHdnGjcPQ0EyLIhIAL1Wobj8
NtYTmmceeNxS/o16sSjP8TMQtXPgf8pC1k0H6TxYvdETsVsvjZlSJk7DqzsVabn2exUYot0CHdp4
FFrAHHXJVwvtK7F8WHLXoYu7VcITIX3x1SQK/IkJ2M+v++kTRjRIJcme4sdhZPr6sO2LWe0K8l8G
qJ5JW6/q163eGwmR6YcdEayqb4LdRFIocxdr6zrjgwr2/tUYDHahCzouuwcPpunEXpuaua8W7bGt
H/jG2FY/qIdSzKv5AQSaTjcvunxcFoQvRnR7ZVSihEyhuenYJxVuyq/7BSMqw/4pulTlSTdu9Fpn
56qnUskvthGuF6ozhd2weZZkGkDdq1iWvddbb2iMc6VOdRVQo2ILQ2Edbcbxvbqc3u9y0K9QARNE
/ppR5HsXAUrPeteHcA4so//LGlHaIu0Gsuhlqqrm5TtkFRnRKlRKiiq/LhKRb49BTEJ2ViJObqvp
XydbGW25y7yulG+T6zjzePHlar7FVNgwVholi2stUNybbVHku/rvhAyxexeC9C/d8Yo8hGIrVm1i
9f/DMf6EwayxidFbEFF7OK9Qy43aDIZkjfjb67mTXNceyAHS7mvC2iMQ3yZr12SiaYET1yeunDhi
tTWi/Dx9safFbT9dzxTrFjN04YqQYlUS6F1AtrfefDJ5ewdznrWpXa8obRfFwPo0Lyn65wt+/aei
Sgu0eKhjPqiKwGmAhSYFGT+0gMJPziskIeaJldUljPd0Xnc03zT8wF4ZORnqD1R/DgzsSb2R3UvE
RtsTrNEuWrKGAfbwRY+Dwlynz3UJqX35fpNuNyiQcRoVhkFQAQzS3IByhMngHlYYnEejZvvebygs
7K5ykFHpXOk4zNVzIO+7xH+ObJqjoy+x089TM2WxSd+YDLA5C44uCmVmz949nu7wueVH7hzoS1wn
9tWOeTSG8rOnF31WOMX2sZo5Bcx7zlryvmOENu44O0S3y6uPsjWU8H2aAPGg/Fvw/IkPbpZZY68B
toX2eSCUh3lLKpcMH0nG8Tf+9l/g0Y+615lkF5jGYkJ6ldLPVED4R+ubBWyIYikVwLJF/LjRCIfn
ePbHDRJZelicf+ybY45UbrCBCxvE0ayCqKPELRxBSFfNJxLxYhDPefrd3lDrAYrxnQ20o73jyvtT
ZXRSnuFjda+gzzYM7iITnfdjGqW9sl4j8GgXj+CcAqppmYOyHBCaK+gMm/NJPUTvpbh7LD8iki8z
K1P+wCdiPGHhiJAzIobC1ulrseUQbs1DEoQzWXgxnSHqtpWVYyPoklANOzo1NtWPDuCUqvbHQRGK
byceo0+l2ToMNBwu0z4hlAd47e5UYeyCA9PidrTjIk8RsflsYVIIq5BEPgVYf/WEkdlDJRxrkAZy
H7/5EB/6k4dpMRopYB9V++IItBzzRkQ6pVaBMUvMBR+pwb39rGR7E9xBo+7QMQw5D+ScZYYzyzil
51I1SedHQv+ODhPuC/x+HrTKW3IrL5KsmddPzPx8muMYm4xPhdRpk6oteIAwIu4g3G4PurAuitww
T777g2agkkP4MKhCZPKauml4jprL1dzw4h224GndIJNCDr2qJzjn1Y6eSZlLc8l5xUpZJD94Mibi
SV5bdddjvvAV/aNpCUNOOxt/+EEtQJMtwX59s7wJKdZGHWZFJy+NIH0MELAlJlv/vAT3BKhpmzWL
sQhhd2uM8fHFs6RcJTkYPItxzJNbDX6fFk+QMJuqZEue8R7zKiYhBCVYImYIjymIUuRe1BKZ3Sv4
jZufS2AstpENcWthxNNldCnA4TG0IS/IMbw4K7IEB6QOzfHKPxzqSvfhwG6DkHesqIN3/lc69yrg
UbyH2PwT8+pUSCh+W3mSkeCTyuS7LSGPO68PO+C942xwEH5pRrnYDi3M9duHsiNjodxVuYKVTxjb
55A2vgAsf0exJQ4N3u+kNlG05XVerQYtNZ88ZEBWT78P64R6NejeXK0sGukOsSzZsL7o+kLS+9Xv
ppp1fTFKmKnGD8aVGinZv3NzYtaQ6gFtme5ZJ4qDhjRofjJb4UQuHUWpqqUJ612IeTmkhtH6wFwO
snRSdO6lbBJt92roAYzxNxM7xJSbDMEyXKp9QLztrKlBtXr7fUYKowQitp8Ptr5tg8oaJINUhaoy
OyFRSx6CxczTwubLpfPDtqGozvuQqUcaWhk6yk7YbTO/mUz19bv5Obq9hXtnJej9xPI46W7QDsIQ
VvJmG03LQN9EbV/JhQBHnD+t29Pr8bVQYSfXY8iW+gAxKlhqu7jR7x5H6cwUFoc4MgIq+374Dzkf
rZcxKbNydv9D8wTVPPy/EeFjrD7KjEpK4CXY3cPSgGu5FBFyztfmYOMWzv4tTs0gsAb/SNNJtbq4
ETg9Jh9CM7zle9a2L2DCsNHr8QZTlyyMLLf86ANcsOprtuAUiryxCUk9WAo7ZxnSBOwWeotx9Qea
0QRYCJmq6/dxmPGXugaxFtDBq8RlfoKkpg24jKPWpHLEWRJzitfQlUc76L2NlC7SwzIzn3xa5D21
Ni4ZOc1MRr03Py+Nt6jHiO0DttB134VhE2cyQ/R64KQOkEacP3mS5l1LE4VtxGhVxpP8bDW+Sild
mJrm9FHcS2PK5NJHMbinDnqbhSYSECQ17w4x4rZRKW2rAVOWk/1x30QhCQh/NVDZlaQIJnTSGKAD
/7rKjuwtERauBaOh7ld6lMNAbVqYBcXfp+CYOoc+vILFwbkfhzUq2+tgXTjqvkw8gbq38LCHPvJS
voPr/HDshyEXdett4LLIsyo9foTQGHJpqdLe6R80yAvpxYF4NInoe8rolbUGD0j9Rf5yv1VGpWsN
mf6jaUa4nfQk0cAhvyUqPnXfy0PhBIENtjwO0hEWVeBRGwaGaAo9Xw8uqDvgolLxYXgGv2mYxGzX
2tEwr04htM/3NQzghHWhgWiOoN+INyZ9icb6kS+aLB9iq0DqY7TJX+OmxlN9rjlKQvhGfH8N4976
aA//iUDo0NVmQJulLtUrhxEeKZGJANWY5WWJ8DtVkc5F3ml+UNhfygJaiw+AyJJePbBCxjsfLM3+
31t07zohiW9sBfvjpnjmt2JtlO4EYy2QGo5x2734g47uIZn/kN6lDnsikDK/3GtJnkPRZ6j8NbVj
nxP8uM/ea/bjS+4YGu2V+iYXAQc5DnNI+8FRw91XdLNs4gL5whNL92uO4m/jrHx+P1CA858IstkP
IuMO7KEsAC/Wkhl80QZqNhGJ2jsX41tQaHfltsUrdGDywu/1zXBMD6fomiRcNQ8iplipAu8aaxvb
tp5RcZgOecwOe4ebaQWJbEMliRjNERdF3j0G5l2/YxwhJ+oTVp2uREFgHD9ZNv0jvx4sGBHx+96N
PVv22UfSmE/VdQ61miUzhSt5De6WlJV3YQB3quJ2I6cSC26mOIAIDLJBkku+T2RNv1cYmdyESAWO
Xk4sSjVxAgmJv0drwt6UfDdhngy3unjqJehIrUMzDCEoGf5wyvs9ErFoWBR3S2WaRLU4aFF0d60Y
JY1g/CKle1Yp+v9yNP+7ZHdFlUFzMzfeXf1S5z16JMlPr5G9eUdDYatEuONdlxCjsy0CQ79AWk71
gGDpjZjoTu/69YaJEXw55Y/rh+fVYeeM5okjATuTJ0o7dLNtA0tn2UlxjoVlfrBOLmPWVpkN1yL+
HtX+7zVM/dqt9EfsdbF+OJRIpdolKojwCUPwwfzFEp4z9p6C8a7o9eCIZcd7Zft6MS0qfLKuboUg
saS7jLLC3dRy6JcmKwD5oxZ89Q00A3D9hvCbOiIkns2NWgjDzOyP2fizfRrWpJ7maL/03N0N0tTN
JX+mE7FLK7pSz2EhkYy/CTXz0vBsvEyJhNUpBuABbAU3PGFq5cew9NYrqYq9ICT66Wayf1PsXDWl
uIAmrcByjwbQbWKa5Bqd0ACyOcp7oh6OAPc7fF+z10URobNvoYZNsN5AgZFhO97ua6OsD19A0WFQ
RbkZ6r4sI6YXRj8TeFigeN4vNBBbdBp3+O4JHsowDV2Vx+IUW9we5GZQdsXldbjsnu3wODfTf8Af
h9yF0MmQP6LBUeuhurEGDe9ZYbtbFieCTwa/yBk/FSeF9tn1x5ntQY40HJJTMY6PifmTNPsCGzs0
woQtQssIgvGHSfdJhUEvlK5G/FVWTdWqOOY1xcU5XekSDx1BdUmOzsZ/8Hh24L7R1kj3dZ33V2tY
EqTcVO7/0P3KbYAGE/sS78ZSqTaz37WsoPKPRq70x/pAzvsTtneEOMoNsW+F2fNRo/zeuPPIBYT8
6YhwZs/dZW68pEgdzJH+WuMEM8vsereP6eFW8EoSRbCXtWQiCaSimvtuSr7gNt8Zxk9pgY78R60+
I8eTPd/qnvAEp09eTF/uD2w4pfO5dKoRxCct9YqQTOPGFRNwt7qy9zZt2jpj/ezlzMZDOKqaJ9Z2
LXfMXwtN+N/E60pz/z90LtDMasFggbGa/MPB9JMawe2kd9RcHmuNUA2QtMgYCrY62MhNf5SplWOB
SutQhPA1TxCYknE3g5KUiGMJrkoyni5KYF2sJcfy+a2ii1Cd7mPwTpbcpoo18IE+PZ6iSorXY6Uf
w+OqJxx+srQUKWCcOZfjE3UBkd9hYjMoOcb9GUQRGxHD44lgQ9SDpMkcsfp76F6UsELVURCbKmS1
/O1a5FO/b+fg3Dl6RjXGTq437cJDvSQeMRX5HWLL2/IbEAefokK97PrGFgo6DVZjfPeSMgD0YR0p
K8vh7tfs2aldZ4P4kaxlI4pfjFgxQcMaBEfbcshOSV9Gxdq5Fwn/O3VWWZ1vp711zFL0bw2kdLHt
hyjy+dPNq2Myiv5+ghBa3H8fZjCehf70h6QVtGoU+MzuzYLwGFgSJMLDWFny/siFrbqrw0SZ9opt
jMH1mQ+OfmFo1QuRs+RNQcbrOhK0Xo8SJ7AOAWC26JGMhTAn75R+3MR/Gjj15Yx30ujoVYeDqsc0
rmjTSjgWOm92S9WeShnCr7X41dO0oCKbKFNr7CclAmi8zpHINHPv7gi1NfHg+QaGVtHmbC58qBxy
cJdOWppdg2Wpx6/RG7+3iF9zrPuuhl8q3l7U71bzMz4ShFBaI+jhmJaIRlzTiXrf2aWEZQ6UVpK0
q/72CMEupINC+AxYtWVxPyXmFeLGZoxrHK4oxTaZgpl66Yy9MRm2G8t2f8yEysBGljBHI6ACygzO
fWXsuNMdzBWHc6nvzU+X4GaS+BJ4TpArRIahqWoChc3wavFvC7eiuKq7PSi5k6T/7T7FvPEfiTBO
CeZrIGu8K5XOdVY2DgwtKTF1DJ1bX/fpsHu9Xu8pniNcSQnaBWphb3Fk0BGwc9m3pDtAFEDeJzV1
2Y2jxA2Cv0cgTGvTZQkFiQEvCHZq/4OeBttITppWs9s8HesnPBaub/0c75Z14N/bmEMhw4nsCdrv
ClPUE/pVBW1/31kHCZmhcmZnC1XOFy2r3zoEl4yD+3kGt3pHaIpTzCL0YXGCB42zVpEkz0VsHAKx
zhLoCORucE09xHOxQ4HsP4yV9aza9GkkF77Hxl/8MmsqYNnzy7cKcsN94CTF4hlc6LarUZ5ek51u
qpiXYKElCLReIJXGLAO8rQ5WQj3kwiABf7vxcxR/uX4JAF+cwyE9ru2r5BH9mt7WZA4NaQZMdDB1
dJiCsDspTOKTEvWHKa1CacCpDOrnak0767zrfJTG8g63YwYgLSVKp8nqegtFfaf8uIa5QhX8nMLv
LCh5OztmwYbEOr3DqQkLoEXnL6YimyU1O7WEDAsp3T/d9YAYsQWlp2YSK1FBvUsmCn7IpNxoEtFg
VANajbPFRxRAwZSj6tEjqOoEfDBFvCJb6cpLIIcPvK70C7fayvsTvnyGKekLc7ljS50gdTzUWl5Q
MKDJCWcqSw0J17BiHFgVYI+EVOVH+u3givumVAKN8Nw6ybBA3hSrHM5vkChOuWDTv5fRpiUfSQKK
XXicM1DwbTRd6GOe/g9/XvZqFt8nkYsuTsrP2yTJURlxLlMN8bA5hReeN26cGhZhm1oS9Sn3Xz0n
+cnVmmhoV+RLbLOkvArRydG8NH26gLgf1ecyJYDQJR8DiMkP+ayCGiM02UQ9PXIpBOribYAoeBoX
McSMOSE7f0lOvLIaz8vWxMrSLChBRsQH+fnUnNkkcsvS8Z4aezTwPraRy/xuxsbCHWg8YRMEnkuQ
LCt1HR06Qw5Tg1e9Seg5rl8cxTRN4hQQVNz3hpfZxR2au/DFjOZGMD6Q+UsF1TezfNMAUVzC08Nh
MtKnWYD3uwp6owtvmmbWhmE7+noTjg4neMLIYUczQLZtlEUjVECm/dt2dK1GDt0pl+2n9S7Ijogc
suqKI0fay2YzYZtw4pCpHmim4ry5dB77XdqLlVMAlp479r1RK1bz+r7b9xSsYWeJ9UjShXg1DJcZ
NC0uw+oqWZ9iJvV+qb05ULPib4kaYUvq4rcNRVvCN3z81hfNB1cXnwmTYTBImJToUKNJTFcgd4vU
06zbym5rabDm2FJkgKcUCQU9L3uBkWvZtRym9rMh0cb6p+ZrPPiQHSfDfDCqyXqiM0bTlCjiePm5
swPiXr1frqcgbcJUQIUfMaxudoAdfgHtfdzWopeMX9Sm27OgmLlAl1cgkVHpNAPu/BdQSgFLvJd8
ful3MARZlgMxCWGl88Q8JcpZf4uJd+VqgRAWBBLj2v4a5NUjCtQdaQaYAhuxi0nAQ6NssVjgPASK
fZrmyzOvWTNU5/KOZOSxOUrr/mU94wO6LPZqsja7MhixgI5OT/4bP7XH0tORyLcM4RM/XJJW2LnP
AluVTasz8l74wIACSzJFRZCzBbNSv7K2NY8Sqb5zRD1Jd/lwbBYtpLO5n85s5M/u0AsYGbPadhk2
t++uIX/pZn//2e576LQKHPLhy8YtYknZbGp+xto6MQWLqXCuEzBnj2If1fUp+558C5yOkXqfy7fw
jzMmLPaPpUxsOQ0ZExjebwR+QF0jSeg8MHWoN67fHz4LYclO62HAIHsQot6+gFUCLr5japDZPcou
FYjUoASnDropDBUrYna+uLmcwJLg6K1SCgNU0f1nRFrLZbBuLMPLYUxmamGq43uslxVwNXJg5Haz
BwtdmgSXfj8bwO4D/Nr2cM4S8Z0RtuxtVMIvSHMa9V97blW1GI4+G5EBsof18DZ6LIZ1h188HKb4
Dz+/SqPxw4oJIA8ytS7dW0tuVDOXiZoUSXjC3z1UoYoKg85Ko68caPnp1haigPV4RHU3qivk3JTs
tQ71xVz7iMkALiFNbL0mDSQadnzt7rHtk0CctCgBC3dvcGTp7w5/D/AaN+P6tysyjyGhPS5Q2Cz8
O7f0c8erNjTSajtMjTygT7ie6Cl//rh7GVGT85uLlBjnPj7eb4Y3aLHwHL3nq7AQ5M92Ee1jMAl7
tr34Da7B4e7ZFWEZGMmheVGYN1iF0aXqKwhBmic3u5464fQ8kQfMMHHFAhcs2iNMCFUBpZUlPYPc
td+npMBTpLRNw4vqheWe7AszSDceSs5ZUQ7hMVmjC4ErrzfLviBOoKbq0kJXwjMxtwYjNAJ84LxK
x7rWC9DlEYU0zWkgm0YVpaRUSHqbMAI/W9MXkBTGW049QjE9ojNv6x+YPveXISSbEnXR5yqjaYLN
p4HxJ3GWHuC+nYhJt907yUCrv1qUswzNEZk7YNUXOPS7wRSANEp4xbEoVyI7NELMwVG9TeYocZD/
eUOJiH1JCC7g02yX5wiq2/q+ajuadrwdXHKMOBvXSv/2b3VW68VZ/ZLlRaMeeziBiN/tWAFzrF9S
QVsKg19khsvvh9ZZp7+LG+molkF5n4/2vpHGPFpmt+8glvIeM4eeMZCztYp0SCK5mph30bS9IvOh
/Ji7MeNXB5mIm0tE3E818GpbeQF32pO2FZFF209558Kin3t2r5JwXsnLy+m4T5Bf+2zjdtO8/iXv
wnwBbfleGbFol4j5A7oKjStp5CAzalKCODsWBhPOrrano9Wn2I2SRTcQGGNGgcG2aF9V3yn60TXZ
JLq7JLOIUXkaai3KaGVzBhhSrXNWISJzCuq/aR9GqAGEeliBzv4X/jSHEodDd/Faw0ycHBy16+AN
TDv1s+YEoteHpORB9PW9w15ZngtX0J+EOVnNBYMNqbg9jobWF2aZfeWj/rn+XJuvoA0uDNm5Fpzx
is62jnAfRn/BHMot9TwN6QsL4JYFb/A4k1h3U8JUZU+qwHj5uO5ZA/lkK2wnd6uKdsCrOCkusQdf
p/5j6g7czKWwoAd+szmNZ0Z42uyLQNevhbHqNryA+HNRaO6OuxmSbc64ECJQ9wkirjH/Fm2F4s1I
BiLBajm5Y026uam+63gJnB+4rECW1ckgsqdVI6N5hFhc6t/i7vpOYkyFgYbhv9lrbGYhEsXzJb4c
BTWfE4rjBe2eYF/O0oHSHdeidHeriCAzIwPSq1zEM9xy+kcN5xID7bmlb0c0TMJUSSdimLWW31ww
FA9cYfNHqmbZ8SPNmBto8KC1Dyh20HfAm1TpuiGjOPeGZTueH+EQJisVdc5EPULKt7ipP+6uQfyj
sBQKt5QBQc1O9eiYBczUcWG997OEuL45ZY8g96K9U2CtlJRaZNnZJYwJwDNVB/KAHr/tW7UxHKnB
a0tgXaaBhEd0+YaXz+i/keUxdX09AQLlxLGQU71p3pcaNkT5R0Djat5EkNZJRIgDmCkcJrMR4tob
GPMOn07swoSH//eJ7pfztliyMoSWd/Fl75oOZSRlFy+Z6aGfKSkm+ETrEwrHv7OgKcd7SKT5cImo
+wZ3M0MtMwB2TjBRS+YEZcQdQq9tNLxOiHNfmo5AJ4hbPa80p3K6Bdmu96BfCKb2Hmrfv+EQMo6S
ZLRds8vzeNftxBeHyqsK951S+koeyBUJdarsSq6AiWV6ilyJ4VW/P9R0CZDgWNjnuEMZ6Mk9l2CU
axKIiPV9blSyq1PuWq8+va7Q+Vg1z4yearv/0N4ILM5cq5p/fH+w5wZgOT6dhgkILFOyNobhaREG
kIOifk3ORAkeAKRTD/oonce+RKGZTQqj3CkI+uzCLTf6zugwzQx6MxFS6MclbQJosZupCLQ59b8O
kwOxNNTEMQPfUY6QZHpbqxFt0Sqk4ueQzAq7aCeI6kXCxn7RFkrBbyDj24OfSL9r2BkzilvP8rPN
M+3j9ZdJ2D5P95xuRv/Zj2DuXKMWUuV/rA0shpD9m2kjzowUu4Ypei5uX77OYjbixpOK4Bb9V7Im
YUyf8Dmyy6swplYL8+iG1Y7HisG+7SDaaDKfjM2Y/3W8grzpnYs1P9WPMJp5jnZxoo2L4/KlEv3u
O+CzV3wMqYS3TBswibTz6DaEa45UPTPi2aAigOrqEdYprjJcAr5pd0+0NHIX+rgYtXK6fB6ugL7B
RWioltAxnonQDspgqBhBaTkMj2io9RzjmZhKvU68mYyiNFx2F8bvP3dQc2yRuLs0UVVBsbZabW53
DgHxbq9OsGvFbk+f2/PnfRimfodIOA4ykr+fIZntMMb/VSkxxn58H4yx87HgF8Z+CnwAchxRzzXX
Mjng6G6tag7bMcfURc5EsGMbnESMrvqeaOqYE8wRMkgANIDatxPCh0jPOGQTUvDt40LxcBkxii9v
ixVj/SBZnUNtlb0PujU4LJynkVDULK+3zC9c71wadhAPQJXf8kyHb8ILYNMgvcYulHNCAF7D/lfF
0omaO1t+/vdJQTRuPQE3iuyQLDRm2aB9VILdOKhfSMikvsnkAweBmHMPnrFVolHqxXUmX2OHdseJ
3M+sT370wXiv3JuMOwslfZr9gRHntEI2k3LeNC7fXI6ZTGg6MjdyHHF0kdFertCyL0xaJMoC1OK+
YdSjbczImHLMiOfA9oJHeeA32wvhCrJKLlcf0G5/KzWno2U7U8BwMuFT6DEfBaEg1CGYV2/lGjHg
i6A7qYYMBP//hrXwloHUhDG4wRG7FJ6XzkTxfGSgQFUsWttYrlIkHulIdxMUd0fYrWyBcLj4hu21
D8gSjlTtzdeSvuN1lvUgGmtn6D7NJYAwpI3Q0RZItOQuCHoLAw7omFwRrWHfU1Z9ZCbQiMuTf3Lc
aRzAQFl1VAGOmDp4AV5eH6KiyVxqIPUNUN2DKUMfO4iU2YOL7SZXM0af1CYJzvzFxNXZPPDuqd6v
hlJYzr0J6lmdOat3Nw8Fg3q4jA46QnhqkNmJTxLWcxYoCnK+xfmzPJDd+zI5GWbNapZ7mXLtAT8M
3CLcQZvc7TTOTbbrIDker+ZOXI+NPMbkIRF/idxU3LkrsOjytali84BPyt3Mahz3ZHdPWNh+6rjS
1ooMpyMljNkPEaqoSfx9aK0rsmwlTyAqFOVGyXErQ3RyumRh3qMnVZVWox92UhN/AD//aF9a68Li
BmhEjYQoPy2Oumr1Gp82GnMYk8sNnPTd4Oh0Olffl3JlxeQO3wwz/dz1UXCKDLeVdEjXYucyOo9F
EvWe2qDZl1RBGQg10MaLGvlFEP7YUcm59W1G5FV8mkLt02Tny42VKBBRJmwr0pniEGBbCKoB8eaY
Zw8XMh+y9qPTB26ErrCtWMo5uJY7DpA8QZSFw9BD0Jh1c4nwas6YoNKc32NtQj9irMENcZxcLVT4
R/rb7F2RVV4pt5EJSWi8SKILSKTbC49OOOkmu5OcKOX930e5ElVq+PLAXWbRe4tpLPp1UrcJYO/7
3Qx5BbFqqP12l89GmX2tFo0UX2uGTXBRrpH/btIBEUS+/YU+jI/QQIQo71VX+QMPdlAbQXaafPXV
9Sf41+A9s0HrtlmHXQymmzmnrmjn/+kQjAVGMJsngDXkk0PGmDz7ElqivpKkjy49RUBF9sqaiCVJ
ivvu/GGriBCras4W95Fpmra7dxkYF2uvtw8gz6gFGmgikFw5EdSJcCxjFl4CTjl6Uf+8L13LLPbO
GKrpk8NLu1TlSQNXzFSFoDkA0AjY8mYmL6mosYHVqI7GLCX2DBSbub43dF670hdWil9SJT/CshiY
m+NoI5sg+c95Cmzu7tRm30GGllDtWG04NURRLt9w7aoYYXDMgh4GAWdGr7hf9w6r2OcnDL0QrZTx
c+zpmdxqlKsjXWijay6CWcqz9EUE9F98gkat7RhDskdEAHIJR36/q+i0ZXxcyRrcxJXVmbAiPCX+
u8DILU1MiE3H/KEK4XQACGaTGpy/pmoFXWSwPBCvFBl8W1M1GkPlGKn++g0Y+cABEzCh0uGwZbRs
CKfLzsSREptVnB7X3QEIeFFCXrruXrab6OF5fstRCDm5yarMW2aBROGNFI1jXzn8rJJnY2Gk/5sg
Z1RfUdQJc3SNv/7SgWEIyf3zmHpe0df+NjUBettbzwVThJ/8+JNUdMt7B7h4wzfQQCeLqj+ak3ue
zTOsnltOsm/D3aoKZGuQZX7MxV4TJI8PxuhNo6lFjtqupe7KrRjqIFNtuMyGzTn7GzNi06aD4QsA
tlinpAI92v23xkbxlZ292WnZ2vBpUz07fRZy++08AzH3CFRFGMicA+4fgRTMquh17QUdmhsBljXi
Tx/0XgQv1fwVTw22GodQvuDkP17Hm7xPyaDR5UjwGYu09YbP/AF8ayEEsa6c6JKDP2xlmX8s1Bg3
BjxhGLmp+MxGzalmEEIplz6EKkH1iWXxQuhtbZRN5GwPl0CqI2GU21LmoNc/lDXR0s3fmQFFrRmV
T2XHcENpgXzf/DipLCY2Y55Bh4mr4qTTNb82A17s3B1SOQOrrR3f0Nkj/eRyB1pjUZ6vwm6YX4mE
EA5y8cgO5tCYmf3am3oW8WYv0OYfoYYJO9t2RCftDx+Ec/N5KnyDlIJYfdps/hYxydSABhlPa/fS
63S2ILOyi9s1YNI0rH5Qb9nfwBugUVJ8wwNSjBuaoG5rkjSX9/VF3bb7GGv52tjomMU+rC8qFM7G
D8jxsBEkGkjzk/dFQv2sKHTZzVuPF1QsxlSanUpbI2MZGLzhXwYvH+DCKmM/QQLqbi2mgj+kRLKg
1ZsoyzKcQbumbd0rk3G1JuHtBclTOdvXX41pvDdLZz0pgeWrglnQ62bFxdu3eSLadWLTenQcBPJp
Yk72z00h215oKR7QU+EynroDeDbwaB/urdi3ZTr59z0FaVyWCX2QGK+F5VTwgZVl/+cWTRSDKXn3
J4q7sDzosQCYEMZEpkqWi3g1It6o3ALiFmK//hN+cj9Sxs7Yn286w70hsWmQLAoEGCPYj+j2H6ev
W3s0h48WHc9IQfrhxaBXtKaRumd4ZOz+nEV8h0XD4KALFpuecJy2cIO6h3RlP+UENyQxzLJaYjpk
ueBJROHnazTj+ZbqB183tmEOe4FpFJwzIhrg3gEgcZ2PaS+yI7XdOjCyx9FMcQzFmLVgJcesIW6l
jUIk0m0lyNu4KeHnSFGQbrK0C167OCj0iu7e2JmRq0N56yCd/4al/w2fYHh8MkQD1K2oy5i7rzjT
yHr5ZPT3hnOpbB2u6R1kqEPpu23SaBsayhbW2faGyWNa0qany/d1MZCXQXLaIWciDFU0Mj7C0Eci
LeA1Mw9lW0wNYZz6kf7/98P5Xo5aBWQ96e/UpidlI3Er0cWjVjUHSvcWOFlMKAipDUW4lkuqf6nu
sk8kXiJTiFmJt+FPGqO3Vrs6P5B0cdapBIzCwxFxWJY3OtAtKMjThPCFTZmZzSrqFE31G+qCVe2N
roO87OcLWWoq5iF/UwEj3D15TK7T40eKFPNQ7kqXiD4bsaelQyhOjDzOyCWDA4NOpfiQXVlanRnh
LOxS1OViukDLswbCIYH0hCCdk+znj6brkeVPJ9MIeH+2X4lPG/XfQnhV8q3QoMzynTuWcDz/iGfh
8OVfHr+pYxmYwPqpX5EGlITZLuz0Km1l3x9hAA41wz828V/E2GB2N1ho1CFsPgst0C/6QY/hRGlk
GT7k2yFAyEXXapHdbxrKwhvWYWEX4poGcyzjUeJo+4ArlCNxgZlhjjO1gP2npHvC9VcDBFdkGLZA
GKsOoQFCQASCHNho7w3XNAd0mCfWQ3wvG66L3Vgdko59ede3sVSN2J0FZEHXynqYQisGltaMSsHi
cRO8OJqqCk2ZbWqhCRFZW+97nlQ+mHVKoQeRoUe9TgAdnDLhu85BRMmZvrUFnwaV5ymxiri7hYnZ
uN4gd8vP7co5OASJMA68RKXENW0SreUVoz+KKQqdcW8VQdFkEkRIQfAI5x3ejc+lkgThRySaxRca
2vNf+vJ7sk8D7oBTWVrwxe7OeTj4h+24J13Cn2nnSr2h9scyovrBETPbnVnm+FTlgrhafFBApETq
3Z02RWZd7vqFcQ0WuJqThFFlLQtajn8zsT75i5aU6KLiIJLBbUq+TgsTA386YH/rQo/BEolfeXYd
6OtczcYcc7jfTArjNMgBlgcRiDE1/4EZUMl6Pw7KXfMirO12umWS2Ge11uMt27kztqVjBjMctvZX
RWN8i/W2qh3xu3eovk4zeX0zLE2IZwc0HL77bVREBOFE11aFza0GBaybKvs0VYZcCaIb9HcI4LFl
gj9TWSPKA/TlfCyISWBMz7WyBgOlNSAYvpqO8BtMmn1qbV5rSMzUFy2xlDy568Np2ySBtrZbpTRW
yxF1wloLRXsly5UMFcHfhLA/tAKJUrWr9gVicmrYdNqhmj3LFqPKF5Q0aTU79JDRB+aA8PBtJM+U
tVXsIjCGfCOvEzcKAbegz5WOWn9IB5TFgDTMKJUAFaIpkRaeL0h7/g2lZm1Qn8waU7tJcN8mqH4J
6vax1TNsw7fOWssdBzTX34en5kgiDFLmOJ1vnJEXiXv1tYRcIqJuUPmmTb09M7h8id7UEfZZe0Nr
NgyqUSdkaRdILhb6vuJx2qFrehOZ1uod+eTNwk121jWJff2ylsxWOTqWZHAqTAsjHUTIl1StUv3Y
4vD12lCdGPWXWuH23O39gKTGg9iuQoBdJSLX/Lozgc4bMlR0FB+WCwHl9+ZtYwecgsZyd7bzwQ9b
jTBb2vXVZJ0Szs9/GX65y+DBU+A1dlCkM2qvnaigWZeguYrtR18P0PCNqAblHHSR2daOxZ+MFIfA
RDL9tG0G5r0MthypicuweHlMdzafRAIFVPkt6S4YBlNjVT5VJQTBUg1+xpRn2nkA5VFLVAT5jpHe
vfhCo+7pUk/5zzqhMhmS2JsOyuEamx4NEzmg1OPKI9Cy6bHtg0zeAuaYMmvVDi2NsD6pI+/FaVmV
HxcPh/kdRu5ohsP4O4KuEgoIbV6/U52pnfZG9+MNY0NpL8iOApTTDna8GZdSSKbTzXes9b7aTcax
ZrIDDuhNtQxzRuo1yPvoC+LRoT0Tcja6U0sTjc/mDnwMXswfTKufnzZFi9fWn/WnC1FJ8gr/hVa3
0uifeuBSXX6bbhHqEzue0nUjOVcpzb6a5sE/cKt5kXZvKoqXBDR/S2E83LHxhTZhlAjIG5+tqBTn
5suJz3izRowi8h9NMcY3xDhvaBkGEONkv6QaTF6pG7ZyPD0xBqO7r3UWsKMLpHMSP41muquSbMJI
4Wr8z92AqL02vUO8zvjtiRWcbtHShU/Qg267jaLfD06rlDSvwCWNsng8oBNsFKkBbaYa/ezmm5+n
nYNiGhBGaJKGaSlZnLeWAISeF90tohWp6CGNFTIyI09tDVj6PeA/zlVz9+27yHo+om4UdUO7kDxy
rlHf7v08GzzspfXCCx8GY+phxQ/0jCC9+ihm8jSBOCzNwdOxezBsbZahLgu3pmJTbXvLQWsvSPer
fwNOj6FWld7f115lWcLEf4oqZnl/hGyDE6YENX9Oy2gfyn1wTJc+qG+REACs6Hh4RVS92ADfLyt6
j2Cj507zUUmHZQkd9SsMgdMXpHspQ+BcgsvRqZ088aQinYTbIQF5MVwyYKMi/hXN0XWS/3v75s2R
4+ZdYbSoIPHY7/s1pYgxCsKT+cpuJdndt5ENPwzV0KVf8MkcTC7C5Te9jlziBiNnKxLqEmcCplRV
HbfMmkVTV0o2YWSgggDOYbpmZjYsGpBh2vDXVGbrEkJpmxyjPzYyC1ubXXgKWvi0XJym3RAFO+k4
UPvvsG5T8z6VqnAYuTKSm6pgyzCNlkJO188tHm/SyRspnCLQBZEji/Z3vc4ZKF2ZhhWUb7VH/uRi
8mEUD340rLlOjK+lzPdKxl+ix+T+XTfExv3s/iqkVz2gX/JsWlwTIq3OEZ/KqzUaqTxG1KiFgOQe
iibi6zqipZpnLM4deE/3M+Jc5yBmxAQvBjT5SzywTo+nT6A2M6FenbYyq9zD1bNgmFJcg3CQ1nhH
TAs+5C+6VK0bAU6OBWDXLAU7ohrQLw1WXARgj0BTHiX0y7+j4aEWz+Q7NsiULvDfxjkOopY2WR9W
zopSUBMQ0AR/Ym5bWDZgb8tSZqZS32NzYfhA+1+1ja8vxvJd5bLYv0N4DCpBUkntb8CkZ5jLpxGe
lC8m63WvcOcUqe3Ilxt5OJ7pNVMxIXEJjOCI7XX13lnDLrK73FSi1dp/bPASaMOh0Tisb3YbfkxL
2sAdcFc4XQigGIcqtkDb2ibV/xmr0DVGe7aQ65CSfPtNe7FbOAD0duv7HbUo7aG82fpHbTIcY+nr
23zDtbOWw8xaTyFqX1dMoyofj8YBFid/D93dC4jHq8Up9Qbe3ReGV6z8jt9qvOp2M9PjCWs4rjYA
fqtkIn+4lJDvlf9YAZge41AhoxVJS9cExHzzLWQji/oOR2HsImUQu/mY0PepLwmx8jzKCH/D61xX
wimWcG/ZsSbp2xQ/ND5FBAjJVKaH5GySe84Kyc7EpiI81dEnUf0SCp2f2UIkbC9MXSrGpD6S+pDc
AAv+JVVzqPCJvVNGkhIVETKLhBHXR8tlxcqQGhCAvG8mCh4fIY+CU23T9rCllbbZqLVnVyRT/aYT
zVIqhSUCx+gVe4C7M/4/CbEzgk4WwW8mKrFCJYPuPnw7Hr2q5gLH8KeGIvD9Eb3rRP2JlWtNvlOJ
uRxcruAonItat3oLTUFppteO3bc0h8yckqCLQ26GanK4/ARgpLR6EHWt6J6GIrkxUAxq+rvqub/h
Eynqo0SC9SnXmLMzGwRdhkTC7ZgMmALQ1+enzl56mf1RjxTpNb5N71wBbD45n8bz2eEQa4g48rlk
d4cJwMGjJxMB0PnMsmrRtPjZFuB7Hu7HeAh+iSkkt6l/g8qoHenifKPOrUkj1C/90fUZj6fS/qaP
4CCdt+Ae9rKhlOVHKKQiLX/LapPUBdmlLCCtjLJHDPYdXX+uCBh+BpftRYilqz20jhDQCBgZkXqB
FbKEqVPP+XTEYLbVO19An3oeKSEtJp+mPZ4BTe0WsqeH4cMq+Yqy0BZ5G02R0K8+5MTBAPbYSl7s
NcMatFxZzMPxE4/lJpJ8MnL+sX5dFVVKLusbSgsferKNW57WsYFbnsbjzgTq+fte+uIxKjbhmBCu
ThUUUGyz8xu5E2gsc09gLAaPOZ4DxmC3J20VHk4VIUrssDZP7V6zF+r4BFIdwFQgoxzc5CSB03O2
3/Suv4LtefhnKoJwj/mg+VLMyI6pQbWqYZLUil3wD1ENRGkXDS++vSBrDsAVnWdI4IkBtRke3zaO
y11UCpeIcV+FP8TVj4XBpZxw68uSuTL90indgokuxhSsKH1Ch6NUzWNU+9vmSq7SQ6951IlFdxvB
/sZkVuzSOhUt8i72mfVN0c0vQuV9ghed56wA2s6GmQ/JQWsqbcpTMfa+j8iX3IzcT9sZ/ZL+H7vr
QC7hTJI5QZt9g5oPd+ajWDCjwywknF4I1IjmX1bvy6b+7LdkGYylW8JdgWQ4MbkJhBwUhs6lLmd4
s0FDZD5zaKpaATNrefXVEw0iG7o+1qglA6IdMvGgAaLqFpBxJ/MAu3D/0f2yS5+WCafByWK0tWsD
xFMPIrBFzcPr7kfG/PLIEy/tUrmGA69nS/+gSLCKbqJvvPM/GdDZK4S9N/KSVO2MBy9gUts4m6uU
Adf03fKNMv0ihKJVal0iKxsx2dn/AzmKy45Ph6a7mMOtWNR8nnkNb/CCL8LkS/z+iwO2noqiNGYo
F8CLNh17NmSSCRF6nQMCbnlXTsgBxLxbwmHh+T5e+8SxZ4bn+MsqvFZETzibbqp6nqpFy7+gNR8W
NIG59zix7ZXu5jXB7JFBkgnMFTTr+rowVjtqzCQnb2QvTkKzfFOTcxyU70cOcsdsUvqdkl1Xjt7Q
IivCcpMQ2S1SaylFFORMk9mzYq+kp54JulO3pwvlDdmbqze/eNbIEuBl9aHiPS9hM40CsSKbUh9a
Wq57DH84bYJQ2Wz6kfKulNdav2bw+06KIK5ZzbmCZUt3R1NJLXxSlOi4ILHiX0gTPFvw6dSe0wKT
+kgkpZWkfm7Gra+40G7jTiM8GBuKJk7i/4717BJMpHYUstTG7Ku1hWeseMCdpxkQs8mtBckUaEAn
M/qKBH/QAhmiRu45nan0vB5Vwg4p1GGa8hndre1Xek3n9FpHYhr9UH/c7iNiZXBwJk/lVVvDeRJy
hH7d8mSTQBSHrtq8J93MmUU/8ccuAcNEwksWGWYaG6XfGYYJYxiOOq8SCzgU2mAQMFLaMovOJlJd
nphB7XdCWe1BB+oP8J3iFHJK/4EBIzRoJXmVcGL5QJjQ1Hd0YmQUYqw0zpP00RsvKDRG+3ipyHJT
BaDAPpeHpq+CoQCXiuFnVYGmuHKipyiwSjfcYs63dRnurJuFX0Erne6m0lkGtiSblrsncHsqp1Mj
KvI+abRJ4OAQWUQxTG2kwl5ck6zpq55PZ9E/LbwWOPKRVZ9Dgejr9mmNFbQK/+GQByOchW8o9AFy
Exr6wP11VnZbqma80RDDkvHXw7UbEYKvMX9216O9A7uP6N5FRIiQzpWxC1IhaZMHVugd5yXJKZQT
mGQF5nlJpeL8obPki2E1Gjd9blL6Codv2m1+WiDKb4DIpE+eUI/6Qjlz/WrNlWmVGafbFB9OaSjt
Hg7Cg5NdCs3eW4lalSNtIW5rOwRqjF69KKqpR8NBFSR0NV2sLOpDST/4wtIOcpu5pFKkWSbFVemm
u+JmAHY7oO4tbqK4ZO3iWrppMFdKAHB8DTpUhpthtnqXACJvXNaTktKTiOpAFLjGH0QLXJCg0zaI
Q5BPVZjL5fObTapWie4o/6v5tId3yUMed/Sb5GuCShbXDJhPP24afM6CFcNwdv5oSTwe2Momz/J7
61Yona6MqhbvPxjR1n+UZ5955UJQ9pS+wWj9joHkn7wpqPrGH1pB/GuRbpz/53Cjp+gwY9Dd5wch
fjwLFZqhQ0rHDLQbJkO4OqxUb7J/xDSYsAkXXfGzxNx5euqY22E1N9Gx/zzsJ7JFIQG7V8XCrhv8
6isiPAcCk02fgsf7mZZtychaFB2VAFvS4wDs0qMqzKI+lWWs61DbS5R1fnb8o7RGgaP7YQ5SLrU+
1M/uH6BMFNL8/uba7Ivxw1VnCQEYEJNpFZwjoZZ7L822yYsChENo6N34Px48JzWu7om1FJjG+IFF
h6FoNPLJM7zaiSZNzOQCgyKJakFnBFS7wms+E85NH/lBrDKkbI+I9mCeVC55KrG8DIBh8tGCW/+q
IUpe8qkmrqLmueAgcoWU58RemyhY35Z2rF6R7Hs7SgGRTJuQmfzaRH1LKwaBY1drjFpmv94FdG+M
yZ3bo8q/UrwR0I8+xc3SjmWYz4COA4DjuWnLcFYdFEDGZW7vACAYxiZym3WM0JnJLdTOEC+A4q8g
3LjTNKgveRliONyLNBiMaMOirNACz77qKD2MSDhru1YEP5LrxMMfjMYAOqAqWb8h7X0tL97mGqFf
5TjCkzkSajl0MKkNhQGgPoV4jxgCVunolrM1Bw/tBWHBNBJzgjje3FsrcW7hRbZ4qdNsmTDWjsfu
XwiECnHz1xAravSalnFu+9NtzPdyK2safPRAHZckylq/wREcqwBiOlVHQ8DbDJtRUX7JEJjdBLNZ
TyN/Vim7k0LFfdEt34MW5SjACoEyvkmL30tsyzN+HjP3dYKMT4TpnHHJK2ij660gBU+9hZARznHx
SLNEyeM4e8m306enB/qHLWoS/TAMqPJ/bJGHnwZvOb61NJJxeOKaIf/HTsBWRV+kMHCiMWPJiosu
EtCPKIu4ae665bSSwx1Zeptp20mRXKekbFlmaBiiZ+STs9yoqtJF28iyu+uz5oh7ULPuKlfYqhNO
izcODUP5JoZ/QUOIZTXGAQCtbH0d+A5OnwEP7KA+IGhuWvhzj0fX+17JU0+Yk6/0Wi9rdkeqhG3Z
RSL5tXAe6os7D1aMn5ZzKrQn++17csnabi4O7Q/m8u4r2CowzRph2LPwFdGroXZv2jd2ASLhETOo
yyOKxIUYInCSqzVlvIkTHmJVBOYUsD/ot2Bg9iA35PF41KfVMkMoBtRh20YMbyZmn/SRVTapdBys
JLGN7LBDvdIFwr8mI03fyi5/KmZuUdTuEPo+jDivX/ajT5OTvi2lh8k2D/md7WClCTwozKxbgDy3
voZSrMwekLV5jp9EVGnSri4iUzPAb+JoN/J5+3yF3CcO2V1S1HFY86O3J8eLsXRNxIpgScEBB1IQ
VzJn58w8N92No3xOwSpIdIO3721ZU/C6kn2oUsXCu9GZ2utxgWAMFXEu8RYIIRW4diMt2xyCEonS
a58nYmIQovd/RWGPm9ySzklwDqTN45rKsuE2dyqjv23uYzwhrLmdo2FmNGMiz/vdSm9Ty0e2YaGD
Vfyp/YHmUJ7TljFFqvsi1eZUxk92GX9GzMirLDhGQe8pxXkxrP5LfKITorAUKb+NrNZtCsjEYOTa
aRFEIYhtuziiKXqN5GEfyshBIrgzDpJkylvc8PlpTNLVH0DJ04aZivcj+7r11Ya60LbipJpBGWv6
On7XQAP2PdNSaUXqK6SOtFGl8TmM4stdPI54lrAjJs+NwYs0fUIghLefRW2v1XJe9ILFJa/FIhc5
ykUMifym1ZPoqUi/DirFXdOqzAna9sxLN4AIhGALKcVkAtHtdOGR9KNgIt/V6qYlNDf7Nken+F3c
o8JIIyuBxA3pKIU1+jXzpAoS6O2NWgwARV0KEtWeRJIsk+a5fnCM49/imQQDeBPO0Bj02ifkmFtc
TNQg7hRYcJ1oZJHBZGpIgPF69fgwDeDYHb5Sl2TpF7rxZQ2vl+VCyi1SYWPQSvBa9ch5buG7tA+D
xoILzuXBjdbFR7+WDh5ScsBFMMtckXaz4/+ldC/m9oLwe0EC4XwslOTlc2QM3qlw3NZjgl8ctW13
F6Rwq7sjOBBHXa2lSoQZLGTUnlEebQ9Sd1/7ILQ1zKGV0o9wxwl7E/8kcjA7N44pKD3H4lxQk+u8
rCvsWvUfp7V+CqRXQeTQMYQXplqoVC4UgvjfpRNXitbGdC20rgKHP9oaMF7OhcS84hEk5XiuTpKA
bPTpk2PFfmayAziArojka6IssiitJ/zVqGcn/xtMX13oI7G1IBKJfI9Q5yko1KYM4No6Ox/ayYw5
dQ+8m/yxG6s90OJdH2K92LKLNmBs6qNpcAc0rLAd+2QI/z5bYpkzJCfDw1xkvCUxUEbLLbXfRwyW
VGZL0qtau4FWHF7X1lHSfmDbiRAgSDlCSg18HfzUJtE0cRIejIUK5GPe+u0KaXWwiPTgaA9VO6Mi
pS/wTXm+j3bdP+BTnN8Rgkma3g6sVE1eYaeodFreoTFtwRsi3IdQslJh+vKib21CbCW3YcWx2OJe
7B66GAW1mr5Cs70gpKezUNyK9gUBK7aO6pxauTpmXbvibCm+08UmYo7MFQxc4Mkq4jp8PVyWBV/Y
rowFVUSPXRV+/Bzp0dJKE4MWJBQ+8mfZfRQ0MfHiWgIIBKDTuCpoBxyXHInYflmWATUyv2uck9W0
aIPiBm7Kzkm+B0Ty7MGEhqcpT44/LAMgNCKabX9PQhBn/lC5Q0/jgUCXbQOQTGD55G+4C0825mAA
DDnflSUrxCjnSpa7wYXpJh7U+Ej7d69G2Bv/hZKmh0ZgKBn8jO3aPAGQ+DoZrW06ZSK4udrIBANu
JTf1XM+9MHYOBHSPckpwDCnrCJsTh2jEj1zM6An/eCKpeu18spsl0v2bcY9j7LpQcSfTpOII7IG3
53Z+oIp1g7sjJsyspcCiujnKeVOPjB15ActR+QfErT2TsMyotqdR5e+Lgu4owPr0tMIRvFCjJ1cM
hVlu/pZIPJ5BAOH6e8e0wLXIVaRVydYjmILFYvB9I+/232LbOKepAbRf+JsY8vxmcd9ZDQlxo4Mc
zV/adoOcJo11cj6sUjnGqLachYngZRJi6neORejiQXVR2cU+ZJgPPxJh2E35UZbhFz4i/OuVHqe8
iILaVvl3pe2RxL7tQZNyzUPucehYzwzFeXlybe0ewkLoTArLVbR5YjkNijiEMr6ceVwTdP6KQ+bA
wl9HmuVCNuQCSUBenPYiAr9INLYy4pinKXeXSZu+SVtoR59EbnHo3HBj6vEgHyaK9/hxArRWo3sK
LtuhL97xWtCgzHKkFCYdSwsqInksvTRkyOahwvVnAZDg4E5JjBGRq34S8hV2lBUplVw0v2xKvnkl
AoettDGSPCLFOQh9H+i6Ry7GQT5mcmI2mioZmNA74LIs20vWP0M53662VBdLBLuPsc895KOSqx6U
vg4ZKw6z24hO1URruoWAK1H/byOb0lygFbFtb03bSC4Mvma7QijCJ37d3UE3/qLQ2oSozqEKylxE
BEu/iqJwaaoIfEZfWRHQRRZfCGApPSM5HLbTERiabVglKCpPUl+fySo3ASkqA2ftPci8uRsV9WZj
qNC2vmz/ZECFuPMEsFxM7hpolSaw7ITrxkokc3FHDRrrqr4YF/EJ+6+r8bXELz4kF0g1rc2MP4xY
s5AvjTxK+iItzRGSfdJW/xeMjYHoHXG8gytCBvptdgY2foscHM0T8LXhOwwTM7Sv9AdgPIuImZlO
b8WpcDRmrx9E7i5MLq0buv9Vc/I9MAlrEzVB+PkvjmlNnU3Co0DIDv3+IxI96bCgiBlV+8RIivxh
LvA+9uXnYgGz9JlqNh3UOIv8oiA555ZjloEz49pICxJhTUW/yPee4u5RZT1Wks/Snw35mzjvakWg
1zvlZgW+av+y78T99MvyPIbffSvMexM4WuZzxdpJFK4GodiQmsfdOvBPSUx9pq1bdpuchqlgNgsL
MbM9RHHiRRoqqiuWmkfEqs8mYZxm/oeI2F2uQXcFYmDACWHRKvnxfRg7DpWBM9Dpx66Om8nyHoep
KdJH7hm0cixxkxcBS4o7jjHIPlfW+88SrXFaexqRBet52C9WXLW68bskYtrTaKO+lZRuGuB+n+1k
NZFmPf2FLT41lxCKDyM7INAp0kt/nhz1caHHwnJ6kKrpH4mR9iJx7cFLAnaz2KZ1yg/SnZqkv7RB
yLYaX1FuKyksN3Hh5jkIHE6goTiZW0kb8UsBiYcbnUiHbVXXGC8c5X0aD/QHpKflsKis08JKaBCJ
csWgBAfneh6aAYyYEdJN9XHyVD3/+frnbnAFWFboMr1QFdVNTNhDzmxRCRU/FWbsli3YjUZKyKIf
s8MG+JjZIv6NoixHnp78bjOP91g98uk1msopSlDAZ2o2B1MQLl/SR6hpNAsAtZM7OneaSeEzHc50
p/7s7OF+RGcx2UH5W2suXgPfd+OanYgwTfalJRI8x+oRINjMpcWMiMZRDtdqsAFL1uNMe0tC/frD
kAHRNZ7UjVQ0vg3PL5hHZaolCGS21ttIefsJqSOwMhOHlfVeC6SZBJ0hNx2a5CFsOXnOZrg5m5WW
rKSGXYpJuKxCySZcXCC5shES7SRoSclzi9h//nB6yQsipq8qPRmF/sDJYpHtIM2wdPYHXAVvZx6s
WtPJmkD82o1/MSQKYHsmK89Xzq8TxLPvc1rxIbiu294kRXVRuA9WyZ+fPUtuwSb6tQrs7UKRarbI
7DS/x4fCHkRsOqlhU/SSTRhQexZdbOxvnqEo/d4E4SzgQYCucdtOqNEXqcFZS0HUb4NUbKV0HNwp
TNnFn2fHcOoXew4S37y2ag1vf3JyiA+oHNYNVNQbBSFW0Ba/Hgnddv9lmMo5jkVe2CCatiKNA+Id
v+s2VYKw3eadxD9WX82EvRsqzLlbJhffjI6gAA+EpzcNHSoqg6U6ounvFfNB8STs8UMoWkhwaF/I
o7BD5a3lTWWLUX9DVeFHJIFhvEa9mF4MIbba6FKshMXaxPNXAaujPKgb1t3ImCk5ClvWWpeKtxLL
0VHZ1YVy5T7mJv3Bo7TOC0vWI8KXCA1JVMkItS+JyVkaSb04VqumsheWuVrRwP1ud8AuQZeauceb
AUarhImwowTSUUDgeHGzjueZzG91kG4n/bNCArnXEu1+SqSlEwsnRK/JpJPVJGtiSUVWpwkqpRwJ
0IxX206MhIrAK7GjI/dXTmzs1BQw9Ksp7kpsiH3BYMDVgy9BWN0GmsvF7tZLbbH/tK11lcn3ELaP
JBTvK6OhUTCiQMJke058bhpWfl47yIlDj/yFndJN975cDXktXP9WZls4zLh4LQsaEF2ZTd8yAy26
RQZiMGFs87YJBgvErj+pUUKAU+vK18FJKeDXpYmgQ1q0n/4qWa2btA6esacaiiH2QNBoyfGI+/9r
KYoWNlB3y443I9IwfDwQko72D+bW19gaicJkXLZ3r6QsOdt93jcrPH7sf1bl0JsHTOeYUtl/L0Yu
kndbUxR+tAgNyxXDRB4jgLHEjL2+ZXepjep7ppb8yCihPkgWBHEjSmkMoZWBcHyRMM8oVdgdWajC
09wp4a3s33Pg5P5/BXTbS7Xi4QbCjXdagH7YiIA3lb/Oi77pSKWo5HUpbjFt49O7b1Kf8B5Z4bc8
DIDTTXaIC2cc3WgqEOgSPv3a1XDLmp2A4BYo9q800aVT8WTb9TvzYuCFzjg5L0ad3YQEnvtpqLKn
60d6+quG6dwVtlVtSv7dmXgPytxdN7CmDO5WLpe5T2s5xbHXKNmmhzskEwhDC0yDps1Rpa21FYsH
YCFcTZ29iRHn/6GcZa82eKxFiu84JsktZcKm13XzbcN14H/+9FGVGgciELWCWjTL7/z+YOL7PnbF
ADPEEkjwLGN5hEcAzmzzlk8dWvrWAhkLlR9Q14GjV199MNCCaBElxi2Cagzmw/4qnYsosSxJTymb
WLni/V+Jin4d5LuBZk+e9eBp5FKvGS+PdDp5e9IrXUJWn/QWkn/6Xj5/j04HV81bLFhKhBFOCdZs
+pYNaqA1sCK85WmCMZwOaQjHmzLPTp8JXFS/ytNiabBgpstKhahDQPJK0EYjhYHHy1HswbQZ9t5j
fj7ENeuk9TIIUWV4W6jSxHxfUWuQQpLRK00ap1P4rILdNddz/t1nORLXwjgAZkCvcfafNqcWvh+F
SKbIANSA6+agr37MT6rTyDLYyaGHvSalMhJqcPefo8mhtiWq1LRQntk9HZqbz4u/wT7bOG7sZb+a
/E1/pudcETk9aIv4puNLnl+5JhbZmfFVojQcznnV6lTrpZVwhaMUBy32VEFYy9pFdvUEDlvDa9tF
6as/h5F92fxyBMh1LcLFWUuVN+OpoIMcGaaxYsSjkLDJeqjjaA20J7Sw5klRzDdnMmt045sJat0v
IWbQxmLHK0cYfK/wieifwq2NVBxDMkXPg/pUR3PZ/tFwzAQL5vnvhCtKI4n8DHsVK8nkGsHU7nfo
zmENYkRhkHQ8X5LgrJZD9wyGOk6vHa5z3+bPB6Rj1/HQKFa8o9lzBoHELM4qsRQ/s22Yi0/FI9Oa
jQm6SXOUKMdDG53/mr0CLR+P3iX0hqx6EGvMCE7HXucLvLq+nShC5ZBjGrQjnBRCCgdkiIivnUIO
VGhQIipcLNIrXMxcH1t/xZady8mYIECCkto6Jl0/1XJL2b0tKHSv5IZC91J2NxdbgErI07dbB1EK
lnMQh/6gEQ4LAxLzqBkwwRFpe1GtVaIKbNV41X/KfKSsR0aUn0wiS7fg6aLTsrY5zVPWqLvxtgwW
OYB3JibAcd3NIUn5PqMyVYB41Z6CtQF0gztZejvJXj9EEKMjfyeZS3U02roXp9DDgoXAkb26pSWZ
pBWmgAU8e/+dURyxYooZWXD9pQxkfSnYFWeQLumuyxiAfSYwghj0BMAX+Gc7ltO+rTnHS/q36sql
6ZfUmePgccgemFkRymnl3FQ7cFmL0gg3RQgq+0Nsz+K2EgkSx4aOwTx0zyoSBfaGwamMrd3lato4
X4AA5pqeYGJ4UO1hQHItHSiJAwA3iYS+rACGQ68IJ2rnJrJV34dcXKg6j+yKV4a2NzXywg+tMGlt
tPvtb81YAdDpqeslr2nsIqMczfSrD2EXb5DBHpB40UszR70eUuNyXSfnx6kPFDgi5xv7j5Xcejjp
3SqtHdr/yNl1aB4jY+Dx8kmvWX8ysRszXq2zlu7LypevZbm+liLg1IuOtqXvqzcKhcNk7SSukqxR
WwfCECUZbTQGVcLepML7ZdTtNPgGoebNkATKT2C/Y3HkFeLJGyFoAYtnkkLt8swB58HxYfYp+Gso
n7VVT7rXN35h60eHEb2eG73uZpf0Sfn4e29xXen43xPKfzUn6RHiC57VVhsKwMPbub15t3eoQEXP
dOLP1P8XoICtviu4zORFUUuKpiYh7TjWC2Kf5AcNL+bdiDWX5UB8eYMrTJvSqgdEpOjUMqEfCtaI
lP43agFz3IlFfvEqNk/AeMGWKy3cs+/8cC4XPsoXwfzByFFlMcZm1sEgJGLEYwSdQNYhEH3Tuttp
eoaAS9ZlHSLmduOaCuR6e/pPg0VrdPvTkQF+sOiQjELUyKCdHFJuel8xsV5s5hff3oI7/bUwrpXH
FmVqIU+a/Wi6TYxzuNZJwyv6Ac4x4X5/fxZusZUQxdkdFKpFwphxLePosog6pYORUL5q4yX9KTUC
HZZbTuyI3dZEvgQVBxYclrD3QRZVLnfbRnp4mJ2ITBmCYhSZo3uGpFqXygL3eClyYcEEWUSLiL5l
RZOwONyub68gmVwWYFf62/DUvEP1GWg1STg/pRL0eXgJY/HTXzAJBZGtEhMBcuHxXqk3JcGhD9p5
TfmSnk10CpipT+zc5tkUwHwCIlbWpDle86PiEFRN2ywKJQOKCB0gFpVf1E8OqKImbfYLDfa+FwhX
oU59Xsiln1X4x0oqFz76TAPMDFlVaiEe7W++b+1EGfhAXxSVJBcbsF5MI8mjHYD4MwwQ4A9Uk5Rs
UzpB8dl/vtvrIq/3Yde4Q7wwymBrTPojnEjsucJ9rAIl/br/2gQw+jhBE/4iP0lpD9wpIiqFGBtO
XgqP84OugZ5DAfqk7pWH1WlRH5nxWThDhBrIu88Bs1CVfLJr7JnaY7yibMf4RF9dvEE87kyR46JK
nmUhI4R8SwE5RIbz4zEyuS2MXR+g2/F0Rh6mrkPnNSOg+oUa8jOnYgsLV1k30HAGd1qcY6tkulCU
0zgkEnweh9koo89X+xgj46oF3t+mFclX46o2cTO34rQh2oly9tq6VxivknZlfpEWxrr6T1/GViBK
YjpKCFaF2sC61Wno1BuNspbi4J5oBEhLu0vw+aRBY6RMS2Z+/PlX3WgAx2qemaAopbbxkmkMGvWX
j/woS0hVdbkdPJFJmR+LovNW7qALfxHQHDXBIb0ilhm3etK5js7IXdQQ4/oSBKGXuc5hFvwW3Udw
0yCjE/M19VwXg0tmyWnYH+i9rz+Jgwd2YOyQYm68vBbfoDLbJTnQZRsaNq/UuP0v92Lk0AlU3WCX
cm7ofoN5mOs1I1x6giqMgnr++46WXSh/aLQQjaXXet+03zYRMJOouN0xwqJ08BWA1oDBwDrrJMRd
THrK8b91WrHfCf61tcxEd/fYN2CoQ7vwy1sjPKhgTnfzHyhYSyPh/TnhKJzoWgLQ4g7+wkPaPnuV
Y3VuzDNR0hNv3B5Iut6gKvLpcSadwfRYutiX/RBz7eYYf8Y4ZWlDCTvKDBhOzdg+Y7FrxHzc+AlL
VwprMdMz6ql37p/7Q0Y1Nod28+lCHpnM8JecRkdl1x8dwm0AZ/uiDEdB2AzvcspbAtz+OdPzOJTQ
JhKhWEUlO0aniRWgSPS0+QxULdCJd1EWH6wGMxs0ounAw81YrCo6D/Nd95xdgjprhA3M86+3APuO
b5GiF1GuwrxS80rhDO4r8+RWu7KGzw7uG+Jt0Jm+2Vvi7srMGKDbIS3t9yWI+KGYWc7ij5Pqja3P
eSzRwg1d+ls/IfwHP3uFCje/SgLv1qDdqgvOUmB4ob8qgctnx/2EpS5mtXmEBWEKPpyuFZzWhJst
EtAtv/hFecJRPcw+O/IC9BhKn6uK4lveaOtmVf6Ckd03+4lZHGR/hldyOJbMVtW/cVJR/IyO2wj4
VYFHgnXLZWivwlQstB+fccAtbarfRKaxtDDsRg2uOXibL/1X6q6hyyYfsuh/DfJVgIOFLKkizO2X
m5YLqktIjOP++CGdbIcYjNxJTOl877UMrHOu2VKoDsIi6NMtsCBfHQyrID0WpQQ5pOaKGVaZTT6C
hDPtMaN2Q/zHMi0HDUF81oezZRrdXJav9WRLLbCKT56PmVyuNRKHMoHZrqcMpxiAOfmWIvh+L71U
BotbgXMvWFHPKu4ik+wHqrtZ0AH1gLlU7K60huImnT5Ypk80IaWoxNG7QJhzW/xnC/EGpftw2PbT
loUnQ3+SeSnCk4xzHwJ4Vicz5QdtorXFH+R6YE4Y6lcuOr1doacurRJtAFEqqZHcz6Y/ko+dBkQ/
CE3qK6j50fc9Wj+qGOP2MBaEzM1MRN1c/nOyDWLJ6lal9sxhjpSmYIyjpu8c3HpvqkOg5eBbxyK2
Pn3UwzY5GiJdrKwh5+LYlRwrfmPNlclWJ9jJtniqb3I8rhYJPc5iSotEnYSx3Sh4r6rBHJpQkMKn
8lzEKboHQYjBB9dIG6tBCphvKeyA74qFrqrVVdvPgSmHMmq8U4uGgW2GArHAlfKB2RJssNdtV8fJ
/YISw5WfGI5OX4SuYYr2VrP6/MKCqLcloLQlu25SPy7L4qj3UJ74W9K3YIoXPZ3lbCbfaTrv/OWD
v7QvK7Nu2lFtEruU0KvKZws/kWOyvD/8JZJfPXYDg1hgeH5B/KJaHGILueESymiTuFiieMBMk7w7
J/Ib0CsjiLV+SOQL4z0wxb6ZgzuudaV+BGQUTmIMtzT2aI7mfG13MC1xSUm1XCk5D1YTnurbF2ls
2zdM1o3WBqGF67pXEfn9szGPrIBXHb7ce/I5MqZTCcjCkN+AqquEPgs6MJyFddhudcdtdX6L+b+E
m7HecDQeREqVNjIMFmb5Qr9SOJ7Uc7tceaLY0BpgnGonhIzAqjEAn5LoogcgKFxfVLgDrqYFg/mN
/Mmfqo6wlV66HK2RSgO3hpqJypEZ5IgnH00rCbN0oOfuH+6TKVIabkKaHb9oHMYo0I6lS/ur9o8z
rIb5jRAGqpEx8z/H1qTyNj5nbFwJoV3nJqvqQMm8rdwTVuf5/ZlxsgLdMgfjqps8d5xkMVaS3IAY
W+jfpIVM3apVLvprOCsTBbMADO3re0ta4DmHgShhWpq6W0dlKFDkdhSfFgXEzEQ44NklbqGkaoYK
xLNdxKWA2mKoDyOl2JFU0D21CSUyZ4sL21NB5CpkKL4xxKXVitMdowaneQ3ktjwKvjyRmqVWwUmX
yGpCJNYqhbkTwYGvoH5xoDLNPlwiKw7zSx7l0EGpqUc520xSOdD2hg==
`protect end_protected
