-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rsobC/KJPwYQvM39rJIjKMWX41n0C92FBsQHv69i0MXBLUdhxq/iVO53Zu6FYNCCFXmYzDly4RqH
t4JfXXZURxOQJMG44qDfjHImuZdPr8nc3tta53BJiBGP2KaP2FbgeN9iwNPsmq295gWb3/UrmETO
yxyxuHHaRRiosb+8rpzqm1r0qFqOFy4Opl4Dgl7EBQuWivVgpuQP8w6fMp9LTacnJifPR/kIkiYQ
1iZF76Sg6FqbB/1DIhVjY60qvpVuP/ZEHVyWtr8O9WZWIDKc/d5H1gBQjG0XqFCjcFTtfIIAYuHl
IyTd0KBe2pUh44r6980g3yz9zOE8m1CMocN4Fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
6E/SiyfDLdrY/zxBJrz/QIsFLaR9vIOXB5zMzqLwZBL6HorIOi5Zd6+J7oJMySEnQXE6u+jHS5Op
g629J+nFqu8geJ8IF9JsxrcEqmgpM6qE/4+rTpYf8zpNenZg3LU8KqTy3e8O/uQBVrWdLpBFe1Vh
JRbGs3sEOFr7pKmwI4kL48mSoUyUTZcm2pU5FV4jJKqRSejgXG02736yA3irEbfRNr9zWMJQ5aAT
4okSL127aoBKXhF9SgK/NsTOShp0B7pVtjsrB5odObIHptAHzICJQdloIgyPIVOb+SHTGFpl01pa
SxlYKGsCDWiDGFC+5E3k60QoMSOI+4VX7dyWtcLXfvhFGMWpU+0DG/YpnGEvF/o+w2BUI1dv4e1H
ehD1NPEgCm6r+UPrIoXRVn+P+b9f77jwxwi/yMbnx41Os/Xc/+AvdF3d5kQVErM4VZ7XRr1jfg8S
ZRpy3ZLNyupaME/AMXzEU+FxigAotHsive6x8OZRmCEhTF//Ia/b/ZWiX2jdvVTxdEbSDNVfSy7Q
oCp6SQHv1pTSLxczV4yvuqYNE4SN5iUOgPn07MIEDf6cCVZwApBLKHfU8V1UNbewdshLpDvx3r+A
hhNap9gI5FDNv5TsFJPzUDZmdZgP9OjzZ1DQ8M6MJS1QVTpM6QMZ/3cIhddORGMen4eE8/CaH/BH
xKT3YOiv7XfT1HNLlEp6jKviowLz44TdnRiRr9+tsNrDqco4a9VjT3Kg+6k62oBQ7Wh6c1KiGgap
R3rkOYrgZuWMSW0B4yQkhg+5GD/4B8fRsQvh5TsI7EmfecOZ3lEvusjdbrPbGv4i1MR7Q90S09Aa
aH0jVO85+Pf87ZgbAKEXA3BqYNGPgyQpObtOoiTBrRtkYC9XXlMY03hfRaF/n9sIoe0044c+zLFn
Z+HdyDgmlBGI8ViNguHnekhdvyVeU8RPrsXXwgWnjf+Pp8SbJCwEmTOM/1ldjDJh/93XCisFqUMM
POwef/OKu57HwHZSxwGIhe8k6aBlnBcViVoCW4q2Ruy9m/hB2rjygRvN4rYK1026dhMwayaT7kNO
TJ/9gN2VH/xYaMXoZImslbRDs3P1IsAP58cmEIKpu4LUtJUmC4h7wUYoyIHwRpVp9w9CKCBzr+BR
eRosrudLLPNhenI2/b5awBBYfXaLtm8zXsxTEkeG+9zRaGixzE4iyClGo7ZZGe9qGuIwJkjbA5ZO
FExOP2vH47ZpMS35VOXGWayqAfnRjQGaUQINozNsc996RVWacsMN0Z42VdYDG8o64fyIVOyonc35
ad5UEinIo7ragD148bQsXzx1I8EoelBo82yNxtTaPqEfyu7RXDTpKcM1nr1KNJXmovNtdYkkgyP2
B8+DBKmQWD6VH3xdRLyH+rq4fNW0u29DBkJLi+kA8pW3b6m6w6zsiSV3YDLK/blzOhu518GX6RiE
AbuGZNOnuV+m1GuWjkSa7HZfNJMp7sdR8Fnc6+PIR0HiZ1ewMtlbglBOJSBEBazF0s6HI0vY0lep
Kp4KWYJicxhc173+vqFBt/Y7HM/bDYHTqEGkINNcUH7IguyjyiuUzGXpTpCEBmXboy5Kg5DW59bB
Q7Bdqp+cBrIA9HamrtY/bX2D3wgr8qlAiVAY82mCgcd12W+i7IXqcmZwBH2oQ3nGIzdgyJKHpv6Y
BbZQUlwxbz1Qoe2CtnZkWa1hjy4Ou8uSJrpHNesFviqW7sadq6SnIk7aqRQqqo1KS4EjUnOsqLdi
9bDxcWBuOceGkfMe2Q5YfsdVouxjfzpWNGtmlVRxe+3bRf9Mtr0SR9FbODW4vT08L29i9ZM3O8V7
dFIJWAAbDbMIs0FLwb7kHS+ZWqB9STfcVR26LB11UCE8QzcJ9jIS9Nw3SVvymCzVtzEAtALu4vdh
xVYasmmihomlkd+HGsiAY7RgX5XRlcbtVDd4Bqa8PIMZKska3BtGYtCRtzGpu++++nBmZbkIMzR6
xuRf4l1i6mRq/lrXUh3wgd83GsLqjQAk8Tyb17SUNZ74HnrHtCw4JUk6VwDfcvq7OUi3w5ZghbjQ
iy/Qdqx0CTjoQWWTI8iD6ktTpOkOGAe6xWE4FAX9xqX51RmZ51CkaE0RvCOf+GIjhZGK5t7ML9Us
jSAFLC48l0Ly+qLOa3lwDXrYrw7LeWzElg2ZWKL0CWJNsC67KrJV8PWXpU4VoVPDUeylpAsHYPD0
8ZEm1GnPYuMKX+luwvthrD/634m0lWCvesCpsprVy7zXlmM2Q22mQGedz2v+3yol2dX2R+XO6nZH
bYGMbfm+o4NOBzBZZ2eZuZge5mjXzYVEFQBkD4lZF9g1on7XelOFXPzsk5GbdXumnwR4AAtwSi5r
JeylA9M6dX9MoNPQ7zIH/7LW3ZOyFKrWK6+uzvlcO3E0Kes9eInfuygzG27LhO60E1DDoSI5arIB
orEZJcvFJcwU8yZ5XDnoEnMAkvXqq3idz7h83j6MoZOzAx9KxILnycciFM/CRivJlzNK/8NvlZHZ
Qh5hgFpbZXztHLOp9i/672XxnN8nkt6W3jGveJsdKUA0Rp7euNWVGw+lrFbpj6qMApVAexgOUBwY
wCDnxsNIlGCO1pM+oSTXmPryGCwYimkfHrdOiwe0onuLK39/6TIGMCR9GIIBzoawmCjEru2cDier
NB4RYbrgbNsmghJxRK/fZ23iUYkF0sSx694DPudpqJzIXG7JluhlkNyXhEKIaR4Wg+bU9gplE+L6
OWjE22CPoF6CWwQD8x6K03nDeJpHrXnjstxB1Rv1D6CqcwTyyFL4JoUpjaG4uyJ0VbXeub5trX+B
Y0F7k6JmF2+rGBfO+5ZA5wSI4TIhyHeo+wcvZcQYP0iNFE/BJkU839qmbnf38u2wmLc1Z4FsfA/U
LNzRxdO4lllljp4UCOFEAv2hDzpLIEjIJ6DuAgPbi/kQFRt22+c9Ecj/6EyVpRKbJR0pV7vRkJln
jU55tIduAeXCTaxviQplhJub2XYx1f8rzpGBRMyicDT8+lj61Fm6a/dTF30hMp4VV5E2x8nZ9hFR
bmu2/WL/DeLnuj60JiFgJZDY7IjeijfY7csW1T22eUctibuFNlTy0nraUZLiHK4xQw3/2fkx7HbI
uriafmtQjZnj3ehb8P1v6r2JUOwhA8dH7xUxvs3deiPc2SLsRjiOenc7EY/1+a6VigdyggIEuVeN
aOd7ePB4oiPZ+I5NaB6u13btNb3eAKsluqwgh1scYAh740AiwQp/ZS04jdpg5YTNPi8nO8IklljA
X7++atHA1pBN8UNjZT5Ii3knDJSlowEynCP8Ocpn1cPbMUXBgI2n5sz2pvaqD/B+mEKyS4KjK0Zz
W/FNNZnMCSCw7kaXqa10SdkBFgZDjLHiWd5mlNS5r7yyyWvb9QzRkQgrBRwwIZZDL+PJq3lHJxaR
ykV4atbsMz+kP9m0Qjevg9FRipQ7hI4uqJQ/+YOUPz4vuTKBEaAKhLJsXdXKwJHcf+2GEwEAWmcE
6o0QnBeFZLiC5KInTfrUtCfqtv+brguey/sZ8IeIXgv9z5ftlAIjNzUTA6O9irOfs2GHoUkrp+gG
ibRN2DFpT+tQ/+05sVz/+Uo0+nB/7RYaS4mc4aoBYOWJvkJkO3xA/5D1sknuH1oUaGUsxLGxsmxo
RGHADGXiDMMwrsJA6nPmaTphiqc4ZSAv6L3b6OY9hggk62BE7jM3c8u6w53dkix6lUhJw0D7yL/W
VGIkamNllsLVdI1KpJlrkBMn6p5hv2Kfae9hZhEiS7mCQ/CYeteyhHXtB2ShBNFVMD2ExJYhCHhL
FfBTYe9oF2EyfRsPFUDrfE11fV+ojmORZpQ4mROSavxQ3HIPzXzrmb+k1NyI4BddjPXjyA3ptrGf
bKAbnyvoqmCyVP9rLmPE1JovMHX+jJhhae2qRaaOlJ1z7AQ0vUAzNxX1td55p3nR4eXgrv1E67KJ
Y/0+UG+dkJIVq5XlFA6qB81Wbo5T8J4eqw3vu17epwHOT8+AJb1zuhUsRgkNqb+pk9sSJGVy2V8s
JiDaAsfvswj/LnqlbLvO9EJQIRHXDfSLaEPXBQ6OCnAiTm4YT6+u/5bArieSlEe5Y0ERPLZf3MMu
XHrY54TUYy69CF3KQmWZzKPHumQ8mjAYT2pn3UGt0HnQEHkX7jdgwq0NgdiO9+xHgn7vvwKPA6It
s0hQQcndxFSKWgX8tupAhwkiFx2+XBWHtTsltakVq8FV/bmaakJCc/fS5irvcldJY3hUK8WhUshH
b2dvbNDml4jMbdzobPxOmU+yhcLtkhSpqX9IA6o3TtRQF+pn5dbWGfJ85YkQjv2m8Ggz+9fi2qSy
sY07uf2tbzNwto71Ikh7mAOnv0mBJfjuoD9FOKovY9qg97/PZRQeSfpeJrIRBCvuE0LF9Nt+Wz2O
Tt4S2hNL8x3xI/njwGq4S6gUQL0d13EkmHIwSfGd44aaz2TWKOEORqqJxmDhD7VAn/KkE19GhPOv
wBAKfDfxYxXtK8ZNAWA/dOZ79wBylvKT/uFH57eHRiyzCZguYOrmmj09352gUeesNiG4a/vsoOt/
y0NdJacxLItlk5ryXSBVI48GjJ9xCEbzV+4JSS0jg8oSLGDoz+hDO0scBWtkyvin5/63CmLbPdVb
73qG5yqkjJs9oLSbu8qBr2lOx9+hHBPlFYfTcw4Lcc83L5WuRQzbjd8mbFh7kMlb4GZMs0t/+NQ5
3GjP9TXCYh0ehhshkHeX9gV9sBrvkFz7B3xd6cndxiQAtBpPSmw1Vzm2xyrBJMtoieK0DSUe1j2D
YU//nbCSmUhT5QWPEVWExfmRvotQxZVgAjCieBBr1gn/2LPW/r6LxTyZGmJ6zhZa1yQr7oDVipof
u+NHuqoaOE9FtgC0/w7Y4W6mJJjXIox1UBJqNNcvttHRcb4EZO/57bhNOremCxu9SWoph+4gMhBO
dYYbMe5EXEfmXfTt/NJKZEpqTeX544nmy2v4jtwZQ2NpWG07K4uoI8TrfTVaWe8b06/vB9VIivTf
ERkyiPDNc0fYvhCihwwuFlQS/3KGwgeFjk4gP3rrAYNSZ6dSR/8lBM3UUf6G1ILp0g9b2RwyV7jV
e9b3XGJHzjeK5rGWbqHQZpaNwaoIZkzoszHYGShMcO17hopIUeCYApc1W07DdPXIGMjTfPBA86b3
gvRS9o2heOPIr2yxuKeeUhy9g2pTPuFuhmTybry2d3y82HWSkwnjsJN7ffIZrsW3kg5G5uSDefYo
e05D/EGj510LlJIqMOINct3pUisLSsWhaaoyIGn/cvSl1+FaEgdx8xCKaiOg1s6no6ZoMfA2/dUO
M2WC4eGfP/RqMXhSNItAOb0Yv4v+/aifkNnwVziOfKB+6aHq7XQfYNMQZOlYiTdDIEip03ESj3Bx
JHoeG+KwGj+QSwqPsop8ufYh5+XDIfIAcMOG0LX1RJpPLP+cMwksYbeSK+2SrRVZwxLywJMUItVz
XBxvpyTWRwEA/M1BFjVbF5OVIwJBf1S1jfER+8W2cykgZ1o2GIbCyG3wMKAD9tfe2kiPdUi3vY7g
QW1xRIlZZtUdRBfmRl5bymJewjVcVLFno20GKn4wlx/dCh12vaB9M6fWOZnVeHDZCgHJ11J8dt1P
6NwVb8gFc0E/o/Vc/pXeWT2/29RTlKzC2Nr1LQf5b8SfAd+2/ERRuNkKfkvyyhVFCbg3AxJcuBz9
ljhufbINOyzFw1Nnk6nLdxopnvUpL5oiPLXH5YW5UXkgyLk+j3jrt2gjdDRv6xPLoJDLyuAr17VQ
zMtLjAB5HOZHdULNxg6jbEKqZ/7w10J0EbDlIFL5bLdqSd15J82FaII7mk/XStXcnzekpUwT5vwo
n55zOPxzIjlZCnLGrsvS+heuh1bNEE0chKyXZdCF9ebF5BrNcK2OL8bhfI0JXcdkEiZbhtwy9L4d
GbhlLF8me/z85q+cYxnhn8CbXQMRD5vdB9duOt98i2omodOTu2nxXjG17WW98oA74kTTL/XmafWu
VdEz5ni23/9VEcv9nbel63YNA4vPybHJPAurjnHZdBCwwQ7RrtoTTtWphlq0Oyfox6xjuWtDGa69
7Eme0HyPiZDxKjhzwZ8tHwjZ43J1hABz6M6SrDMb2siRgWblRBf+fCLUg6JsSp4wVrT8tlOSfz8+
iiXuzHq4rgGKzbGQahRQkZEuXEnth9m/g42Xfuxmc9wO9sdF1sqSEZ1A9kpqqKMZzYlu/BfT/kOS
M5tsyXlMGmx2bWPlGk7ZtH+ePmiMiz4NDFC0S8srUV+eTEnZX0s61WN07Ol4d3z0Hgg5FwL3ean0
0JAlocTaSPa5h+n45Ufw5FwBBA71uSpPxh4pny3ZcFbmmzgKqhmvVdSSDrYLeG3xZxBskPK7mQSl
5rDqQv98mBipE+Z0chm7xsYLeTtqV+qu58r1oMOvUPkQATArOhY9OH5rdoDGjnIbhMDVH3SUE5UX
MsG5ObMJdSwMurzjlX90DTGo27hKh6Q0XOJcZhKq4q3+qJKVSzQRo+F7Hq9l2LxlB92akxfpWnF7
7XOZDbH7tv0r5BRJDK9r06kRKf6XhCT6+fW6PaPZ8u3PkXh9nUUtADi4+IV+clKghJjJLZkhqvLn
6NM9v16VlqFtbkjN2zl5KAlSkhcSArQDrdY+kHuwxZB1fo5Dr1rE8gp1xygSlMC9DZegn/Z0ARK3
j3jlePOeagHXoJ+HxwiVF17VHw4hyhMed37mdrhpPIX4tUQ08niC4H7OoQbM2LTFxO4FDbedB4OM
LVw0TVE0Vt+Bb4YboAN5h6DB9ge984kKJIabG4AtrM9rRAUxUq1a7iU4fStNlS4V7C38oFiJ7613
Qjg5EKjqkIQ2oACdctkCDiSy3SvH5Z3a/6J81IPenAbhqZDQV8a33fHEXbH7IOzED2Pg6B3kXSWN
Kv8Rz6CShxvpnJQbogujT3lkHHgsnfBTt8VOQnjNg1nYBBTt+vN3TTFGU59HuhDOJh/ob7m994zR
DQcXpgF26LQqJ/uUkkwTtKqyuK6Ms4a4lhPdWHej9edpuu/tMzDBlTWXS2lyJGxvANpz8pxZYeLh
SOJaitTjRiJ1E83ur7qfSWPvZpqbQSSyRbGL6k9Y8ySSmtr5VRwsanlQH/Dn12l0u/BbCaDFt932
xhDgjFjR6xp2+L18lNfHH1LyGzb7zh1umjK8+sqMQzpRfEjVRaV0tTT4RrpsRqnWtFPayX6927f1
7btsgfIrZ7/+pbSk8gEOjmBu6P3H0eG2gy2+3kB1mOY70clKZ5nuS1dNK4aSrkwF9erHnuMh6V1/
RBfZgx0sfC+tUifqMV3swy4IxTno3BkKOSyiTZuaXVPki6uPpxgb6Kvsw7y5pIdlDsdQ+rFhkb0X
PS1NDzn7cDCeEN4Xd4iZdBnQnsKQI78gRG7gaK5qo8ZDOrTKDbm5W079DeYqPdmcgSK0YUZ0p0qc
0IBLlelba4S59hNJFVHRQx9xjJmm0zH+Yy+g1rg5V8K5uA4uGQ9rNA8QeWnJwieMyUc02BvOP2Tp
hYw8au7qi8BFm1VOMnDat1jnfAE3rpFE4PaKtJFzznSxy2kbh+7G4Iewz26GvIqdXt3Gju2ZTNot
1Fuy1XrEO7rzd5476obixo3RSRkT69QRWoH9gRX7tp92NOIgbv8Sb0+QEYrHhuGiJFoMh3bZFK9P
+cssNlUwX3kDYWpPxebiQ8adm/ijH20Uj6q7awnKxCqZjl6vkLNfFc/ISaX1TZUZa3k+wvhWdUpF
kVy2baw3o5ypeAY34qoJFLgG8w1edeHQCTDGBXgB2nkPIZf+cVLsP+PFmh6MY17E4rrC4IUjh1Mt
f8AcWdoMSjg+257SkYYjFLJHWgGto4ty3FU14RmePE+yV175UmR9XqOBC6orAboxLlEF5l+HDLee
kZgd1i2enG1q/y174Vlb7uUDtnAksouQB4vDVP0Ow157LnakzubztwLqxZ7/5u7B+mzmArifPUpm
Y0pqBIykxSNoBxTulk7dp2V2oViU6OdXNzAbtitmMK+vNkIK5rhJ1yD4GjFq6/yMs509JElvJ2H9
dBb1MAmrReGabSENKTHhcrkWJ7dJImjUxlgLLcqC2v2PKW1yd70xcw/UFguBF4Gcl85Gs6IBSWVw
TEBmGQm5WF2loNCK5prtMuMtj4T5/M2uImm1V/vooXy0kEsQu+9ytbVL8dANMP9OqB5TuvCwZPvE
m9Ic6spYQoRWraJa8JrQUUqoKuGEkyd/Q/jCoGiKosYSAGxHXRFVhWy84W/VuWtQelbvVQQT6DhX
+VxsC60dE/THkjAH90xC8YCxw1GxnovAAcbHf1pIoPBLn3KMh79P1hn/1G1RT9QTfyBedN6pmJXt
RszpiWF8+Zo8SJzcsxN2wxTTUxS8CfAtJjmUeBr402MG3/ZM30RlGCJjMqW+w7NRhy/fkpDd8zKP
C5fzkH24DQp7lDf7WdVqLlfTrV92sN+Bd4wqp2A7jvEp5pYYdTiukaAtEjtQ1tpvC6SuwjOz9/TX
phSuEbWZ5+7227dbMKsP8FT/GvtL3ODIzzlvn0zyLL6ZS5BqXyN2oi5KDXOpETACQnAGcGefYlKo
4sCIjhj5a0Hs1bj0l+4vXBszZGtXKFdwgRjcIKg7F1yG9a3kXvT+H9GogujIoYR2pS1a+eMUevNY
Yx3oT3Sh3LDWDvgN5S+TQfbI61dTjTKzJehXDesBB2GV+8xmI2si4YazyFL2rEnt/oPN5zIQLUaW
pD5aTZju0wF0BQQCRk8LC+aNTQuS/Q1KHyfhmW8lWI1kFOy13OGui8OoylVuvsMCssb12YZprbWj
YnhviJEgt1JEXzJ1M2wYLZe/qBIprTPxKmc6HN56fh0jDNc7RsdC8ZzwNyerS+f7H9TNs8DuI5U3
M/JyrhX5I9ZdgHfAKWeJ63gZsgmI7iQ4crh2uE3PdftvQPExyPJyGGjhRio8SxHegQ2ep4x6RbqQ
nXlQNx9phSS7StfJKUdt9xQEriTE7fajyJrGwKEuSIx2UMubGGYDf52gbNulihLP96BulX0QRPM8
2YB8vlCvgqww2fRaGIJ8BCeMEa48rzAZHUq0MqqE0jjmtWdjXVFOpamao2hJx3IhOE9ZP5OPlSr+
opW+jXEw2IEQYPkSWZt0BIcv5g3GCyDYlsLsZUpsG3FI8/2+CZHKdHiGhpNIvDTurYDK/gJMovrq
IXHqyuG4XZPt5l8Smtz5Mv6yKkK3BiTqo8/PMb9m7ZwTwrNqKTUuSUEbBwlyLkXzoSTB6TEHiBcT
OCS3d0tOTovtAQJneirUt79rsd+uIUswbMGbYRbkSY2z54DHFhH9CnDIDmO+Nbf/HJxzPN6XXzUd
NLm0WXmLYwoLCo8Jjghsk6gLWwUe2QwNnnfL4/XUuGvSSUsidESSlHzi8vrp/X3KGaBdEDEfWrko
/pP0lXLDSWOt3s8lKWpGZ9qvJ96TDkjbBaSDtqrCW3DB6VdwZGEf0lcEPcV61acjvuxNVXnehXWb
9zt4LttTXzLB4VkhN4Qdzz+bEEY8Nmk7evxhP6v47kW9EDMXlOrYjBmEZSbJ4ogBQmY+4pjmuca0
tfugpsnOllVz17FxcjhhxnerqQSjWluGGCym/ijmzP0N5eoNl+6XAx5lWF1Eg68JcFxoPulrBhjx
JsoATlGjmFgWYdkO7pjMUlsn6MzXQbbCtQuIBTlntCa1/1zLPvNBspqpZGO3SfUEeSFCMh6ub2Dq
LRL/5EuileTnzPy+/krIPFYTDzvUUEob7+Q/flDRs4uXmlB0UJjGq8N2z9hyW8D+IoyHIsXFyWyY
7mtliZxaCRWjt3m4spIPrMBKA/yUlu1oech3F5w22uV8NNOiXjvTCkvQCEKi5Px7cVLvwf8mgk1b
ClRUlA1ygLraf/U5GfsT1okpxyhRtkuw1auKjrXgxGS1wzl/s9kTX8bAyfj9b2LpZs/ukLq6AnB6
RxJgxJp8wlkw3qBnBBJC3cRkL1exo5L35fK9If/2qPKcn2IUvu+1MuGrInF1dMsRZDGymk77C+eh
JNZFKcyANZjOwI/ngJBEQJV/Pq82vPNVUEalaMTwVbaTUbD7c6cEpemlBtN8VuhYQuAs/iu0Abpz
Ezq6wMeFIsp2+2ZEInpTCJ4XqAwpUMjcoFr9CC0AMKYfbIJjP+IBqsal+POe9z2r3K5AWZvhyAMB
Sj6vB5VX9u4x7TDvZrxKRZNYWmcxd27Bn6A61fUuHJWzzdnGzqjGQ4SRgtOtTNl/TBL6mR5sTqIt
0nlnn5SjnbPshGpg+jTn1rgi6HhWKuVE9JFhLEzmcEBvH7JLdG3MXyi/pohVYIHQAdgTsz3hkBTV
hlq8bwth57kJ/69t/zYqd4LxN02LtFNVx9kTwfWHyoRwZ8/R73H/SFRRqAY4LXk48VE2pVBZAZhe
LOZli9cL1H3ViHg1YrJHf2dBnuCNm4Reroiz/gRWycNRVaecVHwRe23YUUFu0wIdTr1aSP2XEFWO
KHf3SeIk3mcGYMFK/Rnkam6hXIPVgeECpTY+5cMKKoYIt531ZBoEBpiIB89tnoJdiH1KDsCFqOEp
ptdj/8mmQBEh0vxbV8XP8Kj3kJfCJueh2ksIbUAHgwrWU6FgzgX1tVArs+TF9tKdGmW9qJRZ5xL7
Mayq4O2lpgDZVuB6yCsSKYjQcsK+T1g6G+6bCD7aac+CBoxZHM3LHLhMqmSfboY1fHiDOb6DlRne
fDmSmi8q4MJuBrvaH0PxplL5/3MO60xcd6egiRy8Bh9ekRIJJLU0wZkOLlMwbe1x8OjP7WQYglvI
9NWstXOeWyRBoocJGSgGtegCeJUjtjSLJbjOyboXeSul55srvvXcBUOmFwzs2BTnaeYRXr0VYlPk
a/k2nGRbTbAcm8iK3RvqKg7S+ElT+3BAwWQfFfTwwN1QvSQxJoYFYwAempH3sLThHTwRZXtovPIi
2kqHBX435w6CqXCV3DN9YynXVzhhrnT/2Cp8pxhjhPnHkrpZZL7uu29GNPE2bkfnb0csMAA5JcOc
6yHIn+4CVk62WVIjDaetRWPi24pi2w/UYpqvAgy/aCKRSnf35OnQ9DAwD01rBY6/n2rqrRAEosOm
JnRIKtkEXZV7GDThxxRBVI3n7H6aW0jY8OvHDjTHV2a4QElvsDlavsaKCurI8skq35Cplw1ZKAPI
+bv+9ov4L+r2FEnQ2snNDPYzJXAUcHRw1bYn/6fP/k60FGbQGqiEiaq6mtgT/STEqvpC8xfZaV8r
zrKZOqz+8ezi7/t9WvKMIEe0TcoccmuwcLffDd1DmtGHlOaYc+7JU04mXxpjg+IhqQuIZ3d9Ca3g
G8W3EPum8L8MJcEOcILnLSL1ud7q995noJbVNO9wDzCS4hxMh4oU3PC2SoblVLUjskdPxhgXsiKx
JbJklKWI5wJDGhWMDc/v7dQqQZPCvo37V2pmreMId/oSyfxnbpUCI+8Hen9IYqQLNX6nRb/s3Tp6
JTeKxfSreJoNqDKvtQRLce01Tvzp9ChTr2T60GB622VZxJ3YYCsnMCZ4Bws/E60i7694p1WazNLH
SDdFyqJDFLBo8XiKYNi9cWULhefDzlXyBv+IOsqnnXhsKlCNBqVpS9QEEJsOG/vKxNZyjdTGfxEE
ceVLUmS19V6J8L7vIsy6oLUJMwzn3nH54F7fbsLNuLs3mS9Pmt5XFm3zbjKza6dp6QIDrt/jNS30
VZ8H2iDOmZdED/iFYarCwp7ASAnEhYvoFhv46K4MqGSoEkJP8Yl7uPgu/Ekkf8Aie2bUdCL0N8jX
8ZGPFTQOoOw4LPXhsQMB/QgodG1MY4z3rqlMKl440YxRsjpHk4+ocJ5F3Ng2+XcTmD3CJJwKlSBO
t3RyQWQR4IX0RNnLqTAhSz+bum28uc8IK+D5WxgDZoSft25563a6bpoX46k5afkI0c8WSJWr3TBu
JSVK8mT5ZpFJQvRm4O/ywkMjWBKrp0pDJaDwBB2YKHY/lqkmfl/Mrjcgh/+LlXba8lgkI5R0wObM
yejDNIW01BpmbT7Sjdf6NsFlNjGjKnqklVe1aZcsXE3Bicymw//QeoD3fg/c5qMcfmwSXfEBLIKl
LoZ1RUXDVpfaBPuJGmEcr829OgaG4sr2q3P5/PqnjLPXSa3J7B1YTu+p5IEKtKKTaQnpxQA7rFa5
vrHJvNwiFifO/01z8/dNgIJdPug3a3V96o2DB2zx/A/v0Mwx7suwxac2biEtnAm/xn933WwXNShE
oAVsy5vBl3Sn9PWHSUNbo0nj0dwJnL7huGiqavGTLksQTXpMpXQHifScMqqiTzwZ2C6jwp2XktoF
oGD9XvSAkWNT0P8q2lEVpBniGu//tXWKC/538YxC3piNrUvUPy7dDYyNQkgjatlB1TTpdhViwb6m
gDVLgJUcKng8KjY6RLPHbRSsj+EfbLjr8+KJw+foQg/XpEjYrWnRfhZhXLz+fmYWw0qsW0KQgG8w
A4fdg+tOEOUX4JLKWluDBUyUBjgdEuyq/XrLSOBBj3L2rDxZsMR21sVwKErPyAMihjtH8xXhSWic
+1RC7gtB+KO5x6j5OBln5rOQeumEnAHKvbxxpTm+nYMxtnBVJi9TAjGmCeuZnNpv+OdP+mGtM14J
zY+kSDr2AfVY2Wo3G8nnhr3+nOYhRZzbSB7H+QYCbe2DsWqU06Ja2EVVAT4Xexx2Tm80od98V2FE
e7nWUaOpgt9hlSOvCUruK7DUBXcgWjyq5hWmIPP+aoTx84+dmZTciWTGYt8n2Ju9bbhT8rsWFWPC
pzchcEedOnlflz0Rq9SwRATRu1X7RIJ0uotpvn6MDtYcOjJ/5o5uZdUFgiR3Da6gjNLtV6s78H75
MrvpSUP946TGsi5L9eFjKIufwAaOipQpBsS6Tlu0YYmM1IFX8uMr7pv27DBLnElVGpOX7JzMqjX+
oklny0UgUtg6c6OMFmpt+szrXbE8keL7fqfLZJ+tAfY59NrZlE7CbDoVIU/crJsCgVP5h2Yb6mZN
P3xV7yOZMz76MgYdKJzTQflH6sLxIHyOZYis3qk8xzMxIBR3m2RmFp5McSAtSw+avuk2hTpeCeqt
b55N/AUzsJ0RMztqzUCdkZppYivHAPaDAHmBgP+6uVa790uajaqX1KNLGWnwEWMzncgWLa+o1zag
lzDLikIENB5ftiUltyOFdheRCEiseZCT6rX492oIQ+elnNPyFRNkuW90aklY/JvKgaybe0ZyGOO0
YB1ELdH/w3YOs4ngLzOzVpXlcRUeO/7WtX6ylnFba+zyYE/D7I7p76yBax1qe3OooQmYRw/m/hTt
ttE8N+JmbQMhNuI1GG5jYMQPlrO8Bt1OisBMJnH1z9slf98g0PLvAtFUcVuze+B7BGSAvAjlk99K
SLDkh+ccpeOne8//hk0R8o7H0upACnxdggs/k4iF8xPAXRVtyizy30iaW9LntGAUCTw7OgYQx6Cd
GVGZTCfvkvn8Z4bt8q+WuCmk3PZMnSv026y/CsShdwb7S3C4Yi1aqQi6vxfGfzCNq2ffoRQhRjW2
2hIAkHPC/K5DP4TQxXHb5Tyb5HDR00JGUdvAEBOs5hk5YyBI6TftUgDp1kbkwn7toeschqTmGhdI
yqhw3d14jbqPfdtrIZUQCfrBu8LLYswNobTH4a2KU6SOocUwhXJONUkm8D/2wYyBjnf5knYrXJ/4
XOq927wxCsYc0MXk0tr81TsnGyEySZNjPVIe0DZ2YuAxPt3deO6aH7/NmXQRSknCJGbMz4lH252K
K/s3ElNzOQRMM7G0ZWZMO8g7ZuNYQoIUx1V5vDVW4d0WHdcQp6LoXQbAGuhyLRuv9ENbWsbCsSOi
/V7NJdUyxQFcdB+3CrGnif9MkxkAMKY7wkBKTilgonX2cdcscgKaNzc0hlI7OS14NeSYxxYdptKr
lso+i8aELuFQKiSgvMb/SQvbomfUC0fE9UYPSL73CjRy+fNzWI+Z9lG7px5PQ3ca8y6hi+kKUqwj
8w2nzzLOVIuvyBbsitoMVEWc9KEUgIQGT5wj3IoVllMCTt5UFieDgE0CaV0gW3YjA/nRdx5F8s/I
gZDWjhg12b1NMEQsBcnF9aulm6S3NIcTCLW8DE5kTR/gin4Df2AAr0iHZOgHupyQYggVa9numZg1
ZRZDF1hr2K6oyUQKCgVAvn4AMYD2j4uAUKqUoRRBlifki4laYcJbNo42+3EkDDL98CHP3t/iGdXy
TDc5UZ8yqeBsz2D0/pRbyAJ3KvygpPqoazX5A23+qfO2bLPkqJ6XFcQxMuJhBjRDJBHZd8Cl8icu
hYlt/Q97BIra+N/Yq9IljBwixpZconkMmMybXzHGRdFEsOYjHW/o3n2LNCoF+EbMkJ9GHGK1K41f
veCrajkicrck+7JP6VS7C03YZ4abaAdIsStd59tFIT5Tr4x4YKS6R0XTLBDyGhRI1TnBDlMQ+kmv
J5P4opSW8oxPYVVW0H3WRoMo/82RWGE57kU1zydf+ezZLOUM3G4l7Q6NxEGWPahsk/D9mMIPR4nc
IzPT3ElLa3lPr8tY07wReKkmW7rbDBVJoPFL3+IpIXpuFLNauCKylHVpiycZtmgzuItJe1XWhkY3
BYCxOBBMWdcr7GDNqLBHegOhLOoNDqSZw/VHGsejWM2u+uTYiCNmPNQH13ryBWAANyfkPu7o8zp9
TWQkOke5af13C6ci2OpE5GSSzPe9qxtc2dTpj7pzjvaA9jVNwWlsLzyOtyiRg2djo1UJb4frpNRy
vcfQrG516Qms1upsXlHouQepnFGBTDVGaa8EHcSwYEfB/eRfQsOIGhU8Tu1gbiQJ5Wxy2NDgIuHQ
uiFHqObPJBLnzpPuRtb7aSjbQAJGCnRtPCaDOQJPhYcjc4QDwaYEltkRAb/lM69zLNAkKoSm0MQ0
qgQl6brZbe8ptg0eQwXCpFcCsbeP7tM/FN8bpbF7bIujJvpGqAHlZYe/18j/DrCwatprzVWk2+7R
wcF7T31XhliJoUyPfOVnOvb6vDAFPEE8YHY67ZFMGOVLHk+nqxzVbI7e/F3KpOuSFG23kld8ocJD
eWlXIwWn2IPvBBVugFLjdgYBlumHiECSAS/H/gsEE7M6anMshE0EaVp4+uminY3WHT3h96N8Udud
I3MHAFIB+bLCLs4gwmrLdRx1HPpPvOEn9f+I01yWsxqtn4p0rxZAC/tq7VG+eol5w/UWdGAEHpYp
eEHmYDTzASaOI5f0eHd2brf8jX4ZUqel+r2EScoH6xtoagrE+V3R4BCapYegwivt93ltTU59LsAv
q7Yz+JVro9fYwP7rVkIvxt5d5HmeCjI/oOfGYVCsdPUKqYHeuvu3CJ51JOi01QUVxnFW9aqvSb1+
jX2rN1Z/ujUWCHxCHcH2kyH4jQKWBRsIzz6dtKjHPozJpjC3WLobP4jNFnOzOzjZYUFKFIqmyL+b
6ItFMFHvD46rUORcsrgCAsWfHEpC/ir1QCL86qDuM5V+S0GvJGy3RF5iOT7HfRf+Dw/MgSyKyADB
5r22wVOhKZF6yiWaoA8joXa2jCakRPaQ2AR/H+CMUgSuqB87W7NEiTGXDpnbdK+vt9sQ2eVY3ist
jZABQc9IWc7G9FngeEcGEGX7Mmr7NfJJtzdMRmuAmk2cFWvmoeWNK/YAy4+9LgaYUC3SHQJif95k
HBsEamsEW9ymJBTEVFr+snHHkvCYzusbfw7R7wWhpkOXxpvW/mMD8u2x1qN83koULKphNVmNNNQ0
HC8aq0sgTFLOq2J6Ssys9YtqW9hlrrJY7Bxre9jSCfUsdaRgKcZjcBZcA8sB6N8cC5yZR/UKN7Fe
HBhQaMh9L/OI17i2gdH7n04PfKqCNaTjOwQ48MwXlbp+n+UUWUnLG5f7SPMPHtsRJMIx7k9Bzi8i
cY25U4+tNdwC0e4KP0gO3xXnPPmDULLNeuceREtXHqs2X89WtOeEjO/K2NmI2P4gACIVbb9eaLrw
myzXc+FuKNEcP7muDNja/hHvEFyKndclPUxdvvAWhuZJX89e39MaAmjA/C8DyTQyUPKW56jED/2/
CE1QDDhn3/Avp6BfOHl23aMMgOcR2ikRQT/xOFfxmcrBZ9BtoX4BC2DZOdEtoLXaQrL72z91Ov1D
597dHS5EsSVTCqUFQ+cFndS+oR6VoVE4/+rV/SQ0zcLXTyyWV/47DR67UJG8uc9YqcANtgWKFSvM
a4OLag5efqbQwSBmkyU+wrvVPMPJkCEyWQtw/OCH2ID0GLQ3ASOZKymejY/YD6mYUMPLKwSOqZO1
6NzDTiLOh9HSGJ06B/PrhnUN3QsRJhkk1SyVZOCZRA3PoZhbtZyGj4TizoNFZMgGoOVnRjTLcL6/
aUvf+aJ/BCJV0bGXICOtqwTAVD0yWERpWUgmbrKg8/c+JpdRXHYJDV4jn1fWgW6RloJK09Gnt7iz
I/qHTBrpvnl2kiZRXVI8VgH6NbGYVRgR0EutECrNnpIA8jno4XJUCHWgRlgyFI0qDuWbeSJ9VsCW
KODu+MSZe4Q+VKSoYWhBH7PeFEwVu/SM7O56iPrUSXRtUMYGP/WLaYakYlPe+BJUFM+xfdUp+DjF
AK7EXwi4WCpK9JQc3fYz+b1c+wmOw348fK41mAQKJ/Ia8Bmsi5jq1ekmnE/EpXxjQC/jLqm7LQSs
TWGTV4cAWKjgvsDS2YkrrFiw6rei69ODOpAX8SkdChrDjDq2D4X+Yd/dK/Lx1CATTkGCdaV6blMl
qAAP2N87oJzfULn4z08jcxJN7OfmXtN2T4lFLiil6cRHzStdRybOZAPGopgjXjaaWwDa69PlbgPh
I0GUuupPaOEnV5o2UJ4QznsVBvSG30O5TUt+Uo0h+0xaapATN8LBGz56C8LHxINzfEMlS95eC9Cn
lwmsL4co7QrTP/YqQcvNADyCee5IQEK0gb5YeG1dhKMAL0BpQqidec/oTSqVkM7L+l7gBXJ3lrqr
Z9s0TgANJ1yz6cKUWTpGNkSNbpoppJIPEXxZAJn3Phnfy6X0eOkpdy5lS6G99Pp1Z5XiieNawb73
djAuVjuP/DvH203ZCNBXEesWEUqMAdwNtX8fXz3V91uoaXctJP6DyuODpudbI3DY2Dbv/FlsP0lV
4WarolEFaIJh5C95axyk3BdKa2e+4+cqcFiLMu8JICijveyRE5YjrtOCx0k/6+oLU9Ce0p5SjwzW
oGtFQYovH5vQMMazm7Kh5rPETczQBXMk79CTsWtCTRfRaE9i8nwgRZgSn4r+0Kpl2Q0sS78mo5UU
EZjLwVynzfvZf3l9kTAShzg0s52QtnyIQqG92x6VI9Nz3U1NAEq/z6jSqsuP1WlxqCji7eMef8SK
j/jNbNX0Ea+DeL+0WkAiQJmpc0qB13D5Wk/NRGM9cOPsbIiDwhS55OxBPvp/awFyGm7zHPx4z97e
YXhQgbeThkHsSeFiaNb1DIbiBpfq37TNSkrhlphVnRdWiIQzkBrz6/w+ONSwgq9rwCnX7WBhdQiW
YWpGx3zfWbmOH+92mPZfD6Vpd36c/rg14McZ/wqqoPa1X4+BEz95HwDqK8raQybErGtX/Tn0IHZO
9NF0lD6aBXsGITXn0Gkv4rwTpcvxyRgkobt3YT65HDbJRH73yySN/LAxaV0lgnHktAUzO9/j9bvJ
Gzi1iZThpISRx3WyAovHUcC9brzP/UrJU7mmfnaSEZxKqzQvYoPhklqmOfPc2K2B0VnzqvcZ9aR6
pe1FovcdVDfEgDy4nFBJbj5mqKyugef/zK8cbSQdtUoFo2TDVFeDPtapaT0PfSML+VHYE1KvjyA8
hLgCe3UeIbcZOrbpXl3S4yrV0jII32hIci6qm/Xfg3LARPS7fBV7HCEqhEoi1ZpjAoF0rRLGaPfW
/AbOXagMsuqYHhxLeIH/HMxmOVgUzuIjKwpwkv3FSISEIAvYSM4RRHJDp2SINVnDKTmh0NS6GLWg
OtyI9dvLjK85qrmyYmBMuvASofMfBKAlQHbTYa+lB23yopsDJuedKwotylt2zjeC+0/TLc3fO1pk
P1hVUag5ZiyuxjuSvwVrF4CM/eFDSLPo1qA42Cz5SDPASEGPS5432JhnMLAokJ5jxNvk5SB+a2Kp
kVsmmv061T8aZHJtfN1o1MsgkpUh399UtgV7fPa4jCsss1TWBwfXyB8StSSxUsA2918vTtABAabx
/cHe36gyAEfRn9Cg4fxyy4hM8tSo37vt4jX3nGzN/MbZQ7JjGSKb4eJ5VL2Zx+4MxqXYQ7RSFdDL
d6seBEEbVDItjnEbN7sqgEr8pyt/Bbtym39pdNMQjImokX5A9Xd5kXKnBh8DGoGxWdVMceNAvAx9
hJNvQdymLZdEawjNry1pud05AP9FPqSiz03N8LU3MBqLIVUfsuzKiwYdo+l/QkKK2mmj2fCxlcUL
5UZSWKFFamkcea40Eis16kjzf7M/bkqw78rgE6Cu/3WjJ2PCcXSfzHszn8gC3ELd6GEUd5ZwMK7f
0cnT1O+vhWnx7tX71C8cOZS9MK5ft9wqoEJYeRTKev7rcbIzgqdmG4JiOKK2rjf/X++ZiJko0mIW
mM2suaXXKd86vHZKris2RvOGvpNwdtJREmsS75prjQos+SqU9Z8S5A1u1j6svIj8C04+w2jZ3d3/
RsMmoe/uDJx9oo3M7DXHc/DZFI93SWcYdsMD1f0yQHGJoyXcV5XCauqozMWjDCKP9rK4FxsFHCA+
wlXM/K9mi5mdirajGvexa+GiVpRyD8Q/GpPgnxmKl4bVFBEKPz13JWx3iUJZzt8y6NiGgLImCzW3
8kEHlHBd6PaMSCXWHtGIbKzQtnBH+WzyMxH/gKY42SMSqlZPydGHzstgKcnI4pXTQGyrhwmXp4Nk
ZrNb6shdJEEkO2urCaJ7XppRpg6ATLih+VadM5jIr3ylQtPnC8Zp/RELYEimy779QxCODiPZ1xfq
lQ7/a1sLb2znlIVXjCC34+pF0QRgBCinCEmPMDAB35W0UeucF6NdMfmgGqGMEoPCKeWYDy1s6Tkp
jfFy5CuIDhKTwmMJVufclK97mB9Al9nnV/gYPFmCBhuuL0lrS3bqb+8MSDN1npCp07wmP1JJO3Od
qP/iJgWPPwSXMoofcNmctQKK1s/0W4wyUEMmUhCM/fwuSnLx7oDDLvHD2s/ROABLW3iB8pQ7fR2Q
WcFzHUnp6Npcl08bMsub9xundIsU+k3R0BckcpqAZndabigz1GIKF1mbQGD5wCrfNhGtcirYBeoi
FDJt2olVx69kcsPdSsD7YODtliTN9NrILnb3UfiR47jXuSx1bdoAFO3fac/7XBAvVInmSublqzV8
R59m/XmifURec48ZCvLlTBlEeeKrUmlqndOC4XACjZGG8u7a4qaw5kOO6W4hCNPqqmk2DyPNPVYg
e/e04E9kdGM4nF1EjAco57NFFdC/gbtTFsa26brJdlb2NjgmmvZSDlZWVOw2swQ+W+AvLVWd+Rdr
JR88EoqVr3V5Flkk8p6N1iEY66YDGR475mmAH0Vr4vxRJXoMbFMZ5hceJgkFy+6B/RGr+TPw5Esp
oQw/hEhAIi3xWyZ6QZ+jkw0wG268WpvhO7RBKXIcbpKjAwywI+HbKESJ/EW6OAdoveE1XIppgutY
kiEOvOcBJuaOfqCrjD1R/dbW6qjVZicYvt5dfTHQ54WNw2ursGO8U8/SLBn10WldvU7h9tAyWxQi
FN3g2TFE1MlDYCcwfv+ge3FnitJwCrGG+ul6n6MoC2dy9WgDChQMCKYxDh8A7kzI5f+1Xdb4Uib0
xddIryq0rSlCyKdoY9QPbbcprZRR8P27b6rrtXFqQGPU8fGya7IwOm67KGjWThwZ7nuA7gaCG8uY
iNTyA9A/truIYD8vgGbYLt0gY915nMWEpKMqxrwqge3WlCR9k80o9kgFB5ySP7Wk17GAOvYVgc+r
LynC+zEiQVeNNhBmvOzTCmBNToZHcMRCcv82p12uG5LJ5/UmD3UsYcSQ/aVjswyUgr+HXeuNiQ0N
LD1eoNUgmZb07Z2HUxLRLUUFSfDjTL0xsWPsjDp3uLN37bOA8mv/Invb+d5oEPKq/U1hiFMjfXQ/
v3bwuSJ7UZp9EMrYI1SpV83Z2P23Xv4YLxkTfxey2EuNE39vTMSEkG5uE8peiUoOO5sgfXyeJ+Fu
Is3p7mm1yTzrz01MM1E4+EsTWKtK+p6bYpoGRxfqz27NUTz60jJweIEph9chf51FrHrUvBO2GT4i
3VPNcVdK0NAIvYOXUkCogYwaVA400NlmQ4N9kJSAaq/FhUIvH9K1kbsfEeaxpkl6thW0B6sjFOLC
KwmgU2HAIYu4GlBpbFy+xPIdX+L9CMLvKJw/Jwo0hh41QFslmw2Gf1kCb5+MebLbKzU/JbpqX6lW
kIfrXtornZHXCJdJy//KdIGxpBWn0dlPrBo3GJ18e5EJnHzGx3niqOvfc03MsqkiIjnjdkL1fpCM
NXHXlBCKF1gTKhcsDu30N0HEf5KzPULI/xFOYKzAk1vVoOBYXoxuhn9PXRNkWRHJnT3dSnz/y26C
2MGA1nliqhC32iIDsHri56tg7pcDoGw/sLStlMMXXynosCKzivngj8yTiakwn2FOkTlxktX+2YGM
hu+26LG6E3Xqam8QRSm/DXC8EeqjtEHQMVXINywzsH9lpwxwOtHsgvar55zYDFcjmjlz/xCCLhy+
qozGSKtrhuti++bm/T78IPASpDkQ+bK/fkiOtbl7KvBJI/7+OMUPLuKTGKI9sBfZ0xie5jX8vte1
MX7aF40f++vQqKMgGOWaVJXdigB2GiR1Zzm++fV0MMCXl7FRoaj5DREebI281WQcEeDSuJ7stccC
1ausK2/rDcrhdljQGnEwuzuXeGWYEa5yWebR8GTgfvNC0Qxx1XomTUJ5DD3YumzI+dGai7a2KYPW
2+l1qj7FRWnxYtt7aJIIIfrHYb4yq5/sguefVCLA22/PkVmm6dZAA/KWIhZqnCgUz1JrZy949cOm
p71sRFgEbrA2k8XCFM6hNkYH0U08JoLcC+V6xv/eHqfRR2ZdFq0YF7Y9t/LRMeGT3s6A+jXiyxiQ
BGbA7gmGdJ+LoR13rWB/oww534YvDNuMiz1Yf+xAkajuxvTnmPz9KuaiAKZlbaHniQpdhQxjc9GM
Qo6gkD8rwmAfNrE1lV8j8HNkyPpvA1kaDbDNykuM5HUGBBjpGnPm0gAUaNuatCyccakPeAzg1r1x
xWV7z4g04iC58t4HxXt0c7DwVJy5nBGo90srbFEh5mWKaDvW0uMAC3PlTRJRCqhc8OaMMBQBW6Lu
cZPgl4G7nwz/GPsptdFYYf6nnEwqiuv9cFvpYBe3vrNuzOx/j3YnQ5iuqyarIBMBEYpi4F5Jejbt
qtmhVBs1x0q6VHj2RqFtFWJpX4PeVLhAkT+HmQ81xkrzPe8fk+0qGBucsSo2K03jJMJUjQneFcDb
ay17H1F0F3uZsZIdXlmU0Ko2zYPj1RN8DKIXOFEJBejQjc2P/39+G4oYX2N39lBPt/snCMKoi6TS
SgMgjs6OAETZRGeRurgW290Vwmf1O2xAUBqhbrvJwAPOORh7XQuNGeaT3awz76UAtJJ7z7hamRt7
o3li1CnbYbv3bHx7ug3/dFAxHbgP1K6+vYP3641+wACBuh9dBbKBRgeKm6vitmhdfbP3iJqEwBaz
iZSp6+neR43nBq4T0snrHJUf3jpPev3Hw2/8kd24/dagVBMWBup0w/IIrFJqxpi0kvmHugHNRJsI
FVkPRal3hpf24qkgou7XH8mPCudlEnxrcHmFackfGNWPhGNiGJwlhWGLjipqjBfjD9n4e+nsx+c7
De5lARlA6jqw6ScqTKgUByajntg+mxflmADnQZWrCUIBqFlZVvYU8lKbbfOsCRv5dJ6Bofzo/YzF
pPMfHd2WqbSW7qJqC+PVpaXjrGw5obUv1wOhABg8Fe3pmFlILReZZ0BqjAaXg+HpM9u0kEbCmeWX
5APeyhxGwktfqL/YKMp3NYZK3d70CDt6bXyivUMLhfMAqxiBqNqgMZAd8w+ZK8ehmEtTf9RRE8X4
IFU3PTet0Fd/W7ou5Fa0Uv5dlWY2iCFoYZ/fmCAD7IOYm/lz1hUZ1YPGO69PPhZp3Vy83Y+BWDde
ZXaHv26+SZHfZ9Mg/0MTg7n4uljlwy2nsW3XuZfIZVNvHf+60sScB5wS91O4z91WThf8fwb/09tT
eapJwWkRo308C0cnV2rcrytFzl3lMNFC6r3XhL82nSweY4unzYU+cJnkbmyhS0V0kkpfgaXhZJPJ
b7muI+i99B42VyAaIOY4TyBHg4SpBIEMAWiPhn5Gxhwdm3dmBSHP6EmAyBSOinT5vDHvqoO2P5oV
FZSuxqwmdgJHPS1NTHTBe0SAeRMwQvQ7pLSAp9ZI1d7dOwAh3/uBHMm40eFmcoL3yfo/MXdPmNfz
F8d7rOCHSGAS0oApxcejBGnE0FDAurPGNRhRNr7Nk8Dl/QSOZ7Jv83SBV2Dw2sacp+DHzy66kNFX
BA+3MLPkMbuTsExg/ux/LexTPm0DYiurBlqJVEHMnSeFVhsNaJQ9y+Ltvvu20DfrIfzuMnMprC1F
/V0aBCF1XoPBRunKvJB/Gm/C3/h/TPMICGcVsxYfmLWZjH/5PpNXiVhFvOgdUiTMsmb+zJOZiDF4
yU5sp7Bg7sy27+XODmZnk6+ngzsIAND/+c+wWjc3GpJVM1YspD4MngDGtXO0bEAbnN/erC6X+4my
4vdRSBZ31yTcLgtWPlEk6ZevAChXy+acUOY7mEu9/GAzjNSd33o9whviRR1fghk9w45BvWsiLFUX
Zbnq8oxExAG3LY12UPxLzcAfYipFr2Ae9a7y1Om7X8i92T1O2C3o8o48aHADarrJjHdLQoMZZeTx
Ia1ho3Dh6aYZ8CXuA0Km0rsshZ+CYLCClJBHff4EeKuHfgdAEMA30CxK0GpU/lkvVVy3z1qRx7C5
wSrSMxRS9JTQXYu/F3ZAOcys/Ct1ttXPyPbeq5J9XLKzY/tbkJVtqqlpcIhqSg1gr95+Zvba1plA
TvE04XAbRhVP4YtLewIaa2bw5yc8+O8K+74ytdSeXXBmQ04ASIAlqgfo18Sr0U9JCRCtG3wTBtx/
EdJHa5VbiMumtITPQUO0oK875dOO4I9ywsrCvmBmoTdzQ5O73g6iQH3Z9VQoUMBNoFY5fi78EFId
CcywM2EEexunGtCyJ529pPkokIJiRg+ZjPIlogI7lJkhXkZwwNT74/cMMhf9dkVrWFzi1Q3ONBFR
TOD9ZOqYJVQmdYDTZXjqlbleHtj5+xNciWw+BDG1QrioAoaLfVR5KgIjYFpx48jqmUxiQWyfqpoD
CcV/b3jlSr67BGBFYGDVrmqf+P/EsjctMhpAua40hVCriwFGSq6GtaZHKK5Y7XTnFSPAyVh14Qpm
734/moLERNpYYSxzcRaF2ltJSUW2kEX9PI8db0o6q5b8qbOrLezZXOkdLkJjOdLowGoBllZv595c
5Q2IUIkbfOqjtR97We4Z5EFx5ABFmDHjM2nfP7sS+OJLfi28Bnnh2bIUAD/0VXODWZVV7sp4joae
+eeYNP8ZiCDk1mzP2oiaRcDSrvX+q+sfF/mAsh/bnF24b7ALuc69fwzggw91FGGtSenvUFi+Z+fs
UHRUKRlZ2kg56BlRjldahIvMG5FKo0lPs/VsOCHqcDr6TCcTsTL+RUKr7oraaj8a+z4RpjuUl3RW
JXKZMI8KpacyqwmyEA4Byu0NyZpddKe7fMT+YNOeFpX2TdCe8Zorn1Woyv7+rzmyXRkHjq4AfkqJ
9WblktvTteNjBdfnimSAjSlNGH4ThPzzcZK6yBr1mDLtpUAS4ibn9vS2ycWAoV0ps5oraTCubjPD
UujAoWs5fZUBabMKgIERJF2uoQcSZHEiTnUHG4q20FwrzzjPxBHyW5YEjBNFMYfI/BS3p5m1vwPA
1f5Nb7A00l/c9EgklTWReFC37+X8TSsSXuoqF2WsHrFrqnHefTXmoLgxdH6lx4qagkJRde8U7j6v
BVsgHt1uQWeaucUK4a370Aj16eYeba4rtOM6DTY8YIiXiSRkzDpkZU5N3IYrXTLb/mVB9nBk4+k/
96fM5eY2YkTJhH+3n9aoISDKme69IZJocbxbTjjaKtjXd59sE88o/GTEFf84e8wWRyOQOi/3OU5J
r1f/r32Wi1MRa97zumq42ObgXDy5ryNbVePkL1Kr29mKRXiyOZayJTjUHykvvtNIPHwUh0TM7fIG
m5BbKkkXkTK7ItTBQu2I3QTl73uUJq96E2Lth/S6ROQ8Bt/axX1gEz+ieSCsYke3YK4HRo4HieUF
AC6weMa1uUk3AgIVhbG5PnN+EOuTZlUa0XilXSUQvwJDlvOqnyvPetGn3mA0T9ry5h772AQWf9Fd
tXPj5oB/usKalJqbbazusAnGqN4EennnmOupx7viCcJ5/XupcDWcMio/TvG06TBp1wrj3jM4uJbN
Af6Py7k4OdwNBl6xlWW/Ey2kZlqvW2bUbNLyYo0ndoXxjmNeBeiC+e7JzZ6O5TCbj6x6FdBExNRC
vdirVNYQwaNLfPNZv0z5JgOmccdFKv1KerTKEm7HsjrK0PAGjAYf7c7J5sTfCFaB6on5OMD+0PeS
D4YI66utyfryGgz8U7c8854ZhDL7LizwVOQNsiBa7G9yCjscK2LzoZ/Nv+j9vSkh7Cj/Xk2QGMMR
U+6SS11A6E3/8Fe7Fbb6RCYtmBbJlXlH7erMTxTOzsodv6itLZUpnpFsWAaccjFsqeFn56qysF8N
QXARnbBT2S8RoW/FEQkXZ2zabjKbSPW/Ig4KBMIWrcFwNHv4WvDA/XRQCKH92kTzSX8rVNz9Ta0W
0cMX7xmX/rjTf1sHi/PIknQTwcvrExw/SK8hpvBhWyZPkALcUFbdXIjQeo/XW2obmS+u8m3lO88j
h6I7oqdgOt5RCaofvq0YjQOPLwLWVUply4mxyxNMwpC/J70RODLi+1Md6176MOeL2sr8coiTWPXK
4zwM+DF7wx74LvSmFsGKHsjQ8MOwP2dBpSqO1igX5NMpju9aDyz8itnkD3spXDheIYFGfPM5z4yr
IzqfP5gijG2jcrpwmEl4m+hTOr3eyzCgb/o3j75SLsX/PeAUlizstb7uHynmdZIc80NzdawocysH
miT63q2BSUm9vN7Yc1kWQNacGzARFLdy1bcAE1MlbTDM4zkRYsfwQzvVEviinZTt2O2jWWJnG87x
8uaC/JKd7lzx+J5Ie+tSLsFEFBo0RZ/cSqrY+nSqAEojIxIwhgzJOgCkAQkFGsSk6RofuTrCdpOQ
LuQJvGWYvUvjUbB9/7kdmzm09gwCIvSeqmWPPumrtitKar2vvPe1Rqrwcx7I+8v7dv30FpWi1WwH
BiCVT7Em8A2RKPGH+fn5ETowQa1NKMZYCRQkYsj7di5k3LBzvNb7SfZJxotABfpr+cHwi71F/ZEc
YdOqRESvYQtf8du1JygXGw4Yx9m1rsie66Skq8ThmkoeBh0RNOFLj3ptkKGYLy4i7A00haTjztvz
4ou4YVGtef2/kmIP11eqQldyB6stP4V30Zj8SD/gfdGeFy5UVORMMI0ZHwhSKGD42Bert2mx3qIr
1BOV682kX+gH2HdfNjfxr5eLrS66FCKuv7Tvdw3M4fMD1SGITLS6zkEP2cyRqu6jEM3TusaBYBTR
qJEIFQHnt50TsXQsMqKgZoKVx/LdlRctYEMhA2jqdZuekqTqqDJNOXV4d/x+508Svt7UDfq7aYvY
XjJcQGiz2GOgZ2sIPmAoxKxktRjGg/eomjO9xaX0dV4Se82BxtkAUZJJiTrXPYjAlDsbt4QDQBRv
bIM7VjqnQ3Z1RhQtVhvmBumkYHLPBFV4O6NyCn44b96TRfoNSOTfFINp0O5VXuoufhwnqYnyZMEO
oMfpoVZo8Wbhr9fC9cFXL5xqBPuY9RYoMabto9C/LYP4U8KAcSSzmKacDWIyPprUCr0EK+R31FOY
b6GtSXK8lKxk64axdmQiRuri1vpjhjuTa+A3S+L1qtQobivcfxSGLsiwCFjsw2XgF3zXYZ31bMOf
kPrMpPT3ZV+yETctrH8xxrI3+XIcrI9ZC6kMQGgoky0xbHfHC1ACKElHm9OjUGXoDK5AhcGK4G2p
IfS8L+H7jxNf3rK08/uTxl6p73gwuFqzGToPo1olF1JZ/SypgZ2dG7ZmjsMlxLISScCahVKJxuCJ
udaPX1yJSuoTtvCRaSCVUxwyUVll/BYckonJFwoQbmC5iYJa0IlnewnjqY1trLsrY2tFDTbTcf4V
zb9TSUegUb5Dz5Fxbw4rAaqsJK/SGPVXqjf7nRyOOKrFcPlnYH45SFytI7ZxasBYYJIomIyf8vQn
TDpqUVQ8gKUsR0at2saSBLEq4k4igkFwX/Yk3+4e+W/CdIzcX65loeuFuIeM4NKy37YU6RmMSSr4
qdJ0rx2K/xc3loWiFiaLLMMqAVl/pUva2BI4Catc2duecZdY1NTJBVMk4ZgGhiVXgAgZVYrV8mUs
GOJO+vrr8ewwNiW+Hlh95HL9HxAKOE3hwxREXpYvrY+/wL71DPDP1Z5Scv1qEktHcec6c0NZW5eO
dpcPfSWyJk3LkL3zqUt6qVl3xTUO5RLoBTzpXKDfd7xy7to36iVpjou8FksMyon0eViFq0WcvfyL
c72Uq7qckIc6ILUIiPCRoSxAeXb6AA7uM2i/w6VzAAB5E65YCBhAVMVgH6mlCQYirB6VIHTfRyq2
2/k/zoeFtW7EYJfi/Yls/jvHVVnbVSWmB9QzDGiQ6tIZMxE/DCsMDWqU17F5bJcK7KvEaTPeZLHt
Vg3Sp/iV0Y1KjrZAMbiD7l/F+BPJZt0xkL+gMorYWkpnIjIRiLy2ej2rA9L71wzxYtu6V6TuJzxY
MYREdmGNbdKK7J8p7u97pf8RZDfvaFz8DnasXAm3a43skvwdngrTRpJVuspDEVZ4RYD6Bmz5JqZ0
/M+wB0gX5Eh5HwiQNDHSEFga8gs3tSkNQgXpTczPXPj5D6cSqMOMUbZHRDRujTqDDQp4AyAcsCj8
gjHqZ7jLqqUhTWCN0t4ur6v+fnTnhJg/aYPF+XSRDj8N1Uv6aPPA2mNU+hi5Q3WCut87JeTHqQ+T
ctj6OBO5FpIRXMgWg7nBGMsqcjMtm9zqN+JxWBOSulhGdj63NQIEURbm0vxvEKNCwgoaXGrPQ2Cj
ksDmzX+Bksvb3yLiTWD2Vty9Oadb8v0msG9uYb99qhIi7JQEhuK8xSWF0ZCHdPqXat3OV2IUfw7Y
m5ymu9SzMryYKtru0sZ3Bb7jwGBgVF1/I7mzf4cTcHHZL4C53VkGB1l1EOJ97hqfxxcGYXAadq+4
MG13OYtDF+ZkwqxmSjeJ73cFSZrlvF2vUKi7ws/06lbl2W4XXLMP0syXK0u8jigh6bcqeRJYVvpm
a74CVimen47pPJtBL2oTtKHp+P2pDs3qhvixKLeCfgUd46CaVFSeeEzFfALqYC7UOfIdf7gpyHpd
iTuvVrEQONaqemc7x+QD6fbw6RZPOsfyyOLebrCRovawqcKwGWK5+5ltbRZksG7bhEgenHir66c6
vHKRzepdqwT3RnEjGe22QQCGhLMXgqSF9q3+srQEqOU0qW4lAcdvQsUWeVyM2RF4kA9bNRPDB608
CqsKiYJmeYttZW6TV6FfOKjKpiA7Eu3buZs826CtI7i5EdfgSCyVZgj77BL/pdlSnHdaTt/cgUZY
LT2QYkz03xYRTH1KKpGzXGUKHNIx0yCtBAQtIQ+HpunYs6tYqxaOkRDYDtR4Ift9LuP1jHyuGoc5
infX6fkA+pv6y38BJD6keTH29v78G6GGGCUUKhhFB2eFd58H2h73jI7Y9oV2ewxmyiwYIltyuxWD
N5l9ZbV9lUn5aRK+9nnA2lanPSqSz/RATqBHPQprkjVro1xEqWJCFH+3gIEvthJ4G0dSjXhzYASt
08ShQz12PoJWQgFPvyj9E6NXGPh/fjXW8YZ36EWkjGZKlIoSQ4Fyp+cfXSkqY0eTDfqUGrfjz78m
4ZJiLdZieRpJkFQ3Ii/ARGNGmhf1Sf2Ubuxtm+i1R8X4gHzOy7It3zAq/kcMNTB/8+MEnhXh4l6F
HAjVR+iBTckvq3Sqgfr6IwxCGn0ylbMh/A2s5xHP5uVNssfTUud3Us+r+2gNUhvb7ee4H4PFCays
qsiVKZyW8uEflJoUH5Y28txcOzPx7AQoMlcNnkPNYqTg1/1TbwMFZJjg8O+6Gfo5sZzsln+aDvNy
qTDJZpA7Cg1SNxFQf0F3cE4WodONo0rjUpi5N/DMhkK6s5wo0RJ5VeHbGbIIwSjioLISiSdPrLgh
CkoJG3oXwpFTvuFGR21pLt7rP/bW0DzhjzE23VcBL5MGK3S/8Y1CoO17pOdFYfa529esxIO4NE0l
FLRGwj3JtcAp8rYaWOhipcykO3IoFE67mGgTIZiwJpXc6YbYNOSEX+AUie+Yuo+7npBPEXr3bEky
bdofojEb5VeyT9LBIPsdOlBUEWFqz2DPL0N4KVxlx850paVXJlqH8h3g5Ti6Asrvktf+55HlO1Xh
eSiJitJpKqvZJDV8F4cpHK037/LM5kdUfUO9z0NAjW0g30KCSE3386DvkbGFvEhw0MJ7OMRRlm4/
8FjrLtEKPDpWVPGXzYCyBmc9Xhvhk7BMxv5deaC/Y6yiat1raWR5rTsOf3DXCI+rejTAhuUIKQ5s
2/OPiyW51zo726yGW87raois4jpPUX+YGvJUIwtJgOzseWZZAmq7u9fWphNhoTRqs8K1Cws3ddHq
mA5TbqmU5RnhUTglSVNQBr/8eIFtNUCAftw5GRE/3o33kHtGdFcs6MAO6fP6dCdSehimUzFCco5Y
H4AJD2HLoOIVOYq1UQWxFt/RfaQLCsOy0vd/vomy4wUf03BAn1IOo0sSQt4DAI7Z6QROy1rHPyGj
VMXKjdVGGEvxfAxhJIjZ0b6Qy2ZYGiBwGLB9/VkHJCCEh08ntC8ynSeabjXDkHhT4qSYOWxh1UCH
yhb81cI65ZeEFKJ1SU83rn3qEDwJMnL+GIaoHk+60JuN/d3qHGEw/wGQ4gJaHbcSTKFF/eISlDg9
qLAAI7dXyGuS+O4nagTcNgTNeC2OX+iclEA5oayF1WDV5geynSEOb+oa5SGXq+GepS9joAmd866X
3bLPBT418m+/2/1KTFbWmcdPR5KI3Va3sW+Jyyhld0jXgQknzY1I7wpQZoYTOxKWea+oZxHZJ20Z
9wRqHUKwiMfKf9HZbpkoiI0sN440f5KT2PlWyOIVtkwB8AMAHETMR/qbBDVRqYHcjdSf+d/Kxr1S
FcN3Mubr9c30pL5Tw3qwbxMgQ57Yn6wnl7Pu5ZHKd0MCn7IqBYn/FasRlbdzwN8nNfWvLp/cGZLt
NAwrhXyi5bgjHWAo6Uw7kwAJ4U0zMpqYTwIzG72/F3mtIN4O74CxjMQmgz8mN8afAhgJP6U+S3Hl
PmFX/WTRBKYMCs7DGAyWpUxAoHI1KkuAqUhEGQb5wf5gJHl0RVcyUn2amhBEITRT/5dXmIeo4vhm
kd8eXZnoO4xSjA2bg/TlTXyalGOrAsl8iO4kvtMDzcR9eKGThAbtcux23Anoh1G+uLq9h9fnkb00
GZ+ezJn7+AOKpFJkQkmduTMBvUl8K5FhjZ3Vv0SI1r7WDNkdIDgoOzYqePP5+22fhnsO1m+DLWnb
5B7unIaMXJP9ukm4VXupOfACiu0jvqdc/Dj6TU6sYSFCp555Cgacal5ydqkt8pYTPt2fEfA66VO5
5FhbcxV0JB4jvi5L3eNPEOXPuqUI7GHCjCTf2Xz/xjo5vp5GetjdnYYZ95PxQYKkzI4F70WABUdZ
hJhkLuGJps62YdW1VGdMCogKtEHvwgxCmjAOiYx3p5lBomkt0V8RJ23EXAkXhthjWGXTodsOycLI
57lje3CJcFroHtwOF+LEk6riAR3zAWVfu+g8vaBJnvum6u/sfgiEO3Mx4x/X6BBrkwYWdlPciI1O
BrRvn+d87aTHUSjnnU9ItsrJeXUr0zGE39tGtE547wogAZwyEBdH+0n7Yb0AzpmFz+Xyn3Tjqbng
AJtLrNM7YH3Q2jMIwxjuwCS8c5t8DiS9+umph2GME4G0XVD+0bQSX4yytQtqQHIh0xFOsbTQcxER
Oyd+AH0kR6COAgXuuFqD4OxrQIcH35y4+E81sBBokO0Uf0vNxNdq/kxD8QfOJzcIt+lZPcn4IYN+
hvJFkOk0xURtZ4wJfeHK9aLWKQPhq1Mc6892e+lGu9srTFAziM28GmvTyJuec2Sb19tn8m9o9NqV
PE0KCF6R3CkaYDeTTcO9WbcMZsKL9FQScKnqe44ZLlOgamF90zKF1NxxOvRooiVPqbkfB4oxhsTu
5tSsqbLpn/RRuTZEOZNIsESJl9UIdEnJgy0NsPCVqV0GWNzjlLXYOT6dhDFAzcURe/+zExbO/ukF
RLI3WmzVFjx9y26xOt+9FWIqWpfqjKl48clCfER0/G1pNL59UkmlhjxyV/Fhah51EYhomFlPe2Uy
7sJGzWBDXw04su+Tzld1IYdbDlHASZ0nFPTaqKDSzA4fyQLg80cDt0TzCti1jH3/NnY+ePWtPQ09
O+Q/jnEG9nD7TsHAcaY3bbhv5mx/0TWPZbyiNl3mV/yJWl/ZLRrVOT11Qx0yf6xKpN5PnTy0FAlz
IvTfP9InVhof4CLRlIdtrBVZbHBwaxDzO58VG0IR8y4S8LeR144yFPq9elUhV3Fe6nKAXqNs4rh9
oElf/xywDOcNIc81G+F7baTaSEGykeodM7Ot/ANS+QggIy7x02fqIITJVBxMTM3Ju/qAtJmwY5yu
1qXNzO8+GuBmsAqu0ZdW3nvOo21YaZCQwMDhtI2ELpsLzh/G9jI3HCEpjGzmdz5E3DwUWhEybwQy
fX+khhk1Zqyvla3FUKeNvTosLNWpk9NGEZArwz86qNgkS+QCRPS+6gQX82DBSeMyG6neLUEtvyTV
FIW0W8N1bUS8YxS5W7JujQvO8jhL3lgzePAhreJYHrJr0gvC6h6Amtos/btR9A18ftMoo9rrXnV3
UoE9sEsKDaxxXSfepb7dUkvbBi4/FlbieqNMB9thCflZhzdu5T4a+8vVCvveNwRYjbe1NxNxGbo2
oA7dKOQYVbN+6CMzVSzLO+2ptcW/9N7XU3e1QNzYbvbzs9pwf7AuJwo51VbAapfx9wJODP0Dk9Ih
mK3wL+AhpFwvtAmXYBAFxUap1ItzQSmSyfYQf4lxY2+5S3hiOePmXsdRvuwghUJXyYTKN2G+Z82o
dEAP6aPlOtlNT+OZYOxpyY/e4aYlahmiEVMgx/9bUX1cKCn88KYxORdfiowWI1IiAJ7zxqF/t3AA
uLhDbd8sQ34z1u1xegiExewzxpbnVQk1CVfZnHSCelQkswEU/jGrpGnLlojaEu/J90xgi+fmv2PL
BDN0OUF2kwLnbo/2yJz1oLK/cDYcNSA7DI75gvhE6Oripzr5nYbnyR+vBqWOepmIZCUv2dyJWGqX
Od8M/XdadCNWoCDr8JbDWchrm+CK31ZOtrqTokKL+9hsrk0hSQsYBIDCh1Uk5zDTuL1P/jyIj3SQ
QE+0uy7tpW5nkvBS9b3ChTEcFv8OQbl6efbWEIaCBilT6tBb9MsQg2UkyqSTtFf+iy1yE8flXXWK
jUo43Z2fWtAmXrfsum+rre60UQ5cdrTxlJ/WxHBZOpV9NOSw2IXZ0QztzQwK3kOHqokUYSA48AtR
vd5KmOEE4u2ZCF6bNVP/bdbAaBb/XilP0o/nZRkMwpHXqAGRHyOA53XpLBLkUBipHR+tqF0YDCol
kSXjKJI0AgGb/ehccsCbFcyWYjzoWGWsyvcH3oo09teKxTglbw5MUjhKjAYn0fyaAW6PsTRWkKL4
PLvKTfRn9h2lIrz2mKP0sg1pGioCIHjppNVsBA8rZN762EE0vx5mpTY3KYS+fpFpYx+lf6kXZvB1
kV/nEzENgJf5KRX1nxfEinr/ZhytEYfkDbucRZ6DJEsNsoCf/1rRTsX+L3pls+W/uHt1cWUapZS6
5GEqE9pa8n3OJd+cnQO9OUEZdvXkOGD6csD90H24PziCg4w+O5XVmpsMNa+jOdyqYm4Ghl/fZN4A
MO7wV8zqrPW6s7gmQ563uCh150shpzc94XA+Pc7dAdH0g1DVeUWH/58GWHq2XvGxu+4VmLmEOmmt
bhzDoVn7kg0OyLfwJuzBwf7bfpTLgDGN5C+O5DHDs6MN1wHDaY98ofGgojUgOSNVPChXwh+sd5GZ
nHVIm/nhx4UCuSQdIGWd3YxS29FXA1r3jrhcCFZMI3BBTSg9SAH2oT5IyOW+m8o6867PVS/i2Lnq
ZjCwizb56Gl/bsP79G1ugIyZbZUGwNms0WgzNWo7PbEVuuwER9BlbgsZCWsKa3fQJgoX4FzvhYtt
al5haNT7uQtipdF2O9oDda8mqjvecfVAdfTgCJJdR1n8zr3BSVYST4/xxlsWjDw+3+8GeQPyBWH2
lx6GUbmkSDoXb/2oRGUUg/GtKJfMmt+wy1v7oAp92O1S98t4P7c9l/FMQOv3+UvtDeO6TmPs6u2L
s1tBZgno8sK/N21q6Y1ZrGcJjNQB24C+5133h5ah+lqNY2wE8iAPCI2q7PDaMfoN9i4gcbqm1m8p
V20v2HrEGNvXMOZO2C7i/7Oq1BSgP1CMQNLK/4RTeqlvAiWX87SG66A9w+462LNC2g35NzNtVUJ1
5EIhBrrlha+o4QlrhEVIgNPLH9OYWxufEOWWqRiOeb4cJVvDL3UF+IRU9qzgB61gyu/aa3t+/3jk
+IipKhdFSUIXyMVwQiAcu35Y9oHJThLalh/ha3W/zxwDnNgBoWUEdCwgRwYl7CCF11kR/T6pSjEw
uwhkro4qGjDyysUjqzH8Xo+JAo1rgKAI1g7RkHzCP6JNR+BvrWzuH2WQN4UPLVHflTylzsdcR34p
waHm3EMdT6tC1bTg3I9zwwzv9q1W6wopad75S5lz7eK4hFkdAobpA9cw3b1MOxw3n5vzU6fcZNdL
mWlBiz+M4kQPeTAuwkotQeBdkahIOwZ6bl+gZQzHHCP86b+YC+QgWGuIOLqc+sqe5sSevckWzLVI
cVzSNCF3HNBavyoAKhx42a77IlFYH2TrvA+3b6/RvNf7d4jFSoWeTEXfNXrkQY+MIg6ObpCqRhCs
qx5RLUG3CrJykp5KltcrJq89h1h4ZO/TdlNC8jb53Ji1fEzp08gvlKAUO14Dca6VnflQbgMzmQuP
kFK54ttqemHjUkcZ93CVdf0x1GpE6U1FvmC+zd5Q5R7QT+ReIoBqFlxDN/zUXsThlbDN/r5DIuy9
bDRZLVyXkW41Ubn4RE42c9TRCSPvT1DLLlyxrK69IL+KYZPyQ/4KwlB6lvY7a02GSCCTIox80qfa
KwT+0u5VNhpcgV2BIkjAby6LpSCoOw7s0bL/MoQeArHQDHeeZQCvuiaB6WoyR/30KZP/0YQTZ+kL
8UY29C56IVudwpuh1zX0P1Y1QSAPgrESm4xbvbceDI4Vbmopzp4uKNMWM5qxpenidyHvRWBOkMEC
I9/Wb8+ARiVrTANo72Dazn0O4qfvS+zLO47TCl6Ao81EngDPk7A+PoVp7IwwA/tC/bpYR2M6szFi
B1K3Hd5xWUYbWvF/ZjNWM0WGTnHHdQzIEVFvLvWthvnEHdiCAywqwoSyUqS9Pjk2QN070X4qKun/
bR064MHDx4CsnyIagSpfERdUffxCN4GpIvhMX3McvtENnoAsVhN0zlwYP+xzitKFWz0ZYyxMy0i1
d/YB0HkwB1uJ4As26zdgF5gkv8SOICltAejZjGC7RI53Y4S0Qj8n1ahTJZBsSYADqFVwuOPpUhsQ
43EWaQpHh21+ZpOw+vO/dH+U71pTq/MMgiWjhsofWBGVREClCJsDGvFWZmMpDDB9VSoIAgDskKeA
LiupENkemZRymi/SYdTdCtYp+Yg2J1iqEQFcrSOcAGBwtmsISX0xG9DcqX2RdWWSsXn72x/ym4ZM
hG4C6fLdY8aE77D9TX1vGIYwIkFDw9AWxHgWcSYsjnkxTTiK2YR9XkM6anlkMheyrTVjS2WuhfgV
1QKFlo3/VdVEFP+irNtktkBAUfQV6HtNCGvSNFxIHkjeSdegZTvLsEgP0MvC/XKox1+In4FQ1zTr
iI9jyIakgs4eEH8Q9PwX0mA3uYgDg6rmU4fug51SfBgwwYqlSRE+BA0a1/TqEbcXp3PXfNP4MMCx
cmNqsNcRfyKbiQOzX+qQPb37Y6OBxFJ1Mb2SBGisOtQD7wCoUkgOet1yhBj2serNW+hMWOo1LPAc
LY+8ouYEE/aU9mVYwJAz1kvmAhm3RuND02fYel0iOsf7H5JzVkP/kJSANviGu2lYFWwPnilUS5y3
8VABimI8Dv8RuwLdWjN1T8dHlEfscxSoMzCfTb5oF1saOxqS2O/g9A5MbIkYJtFzp+YoepHkbtF7
JfA43R5G8yPosvNONHJwnZQ/2ns+7BtpHWpurE1nH90i9mXtwYNZgL3Q1ymZtZm3Ph+QikI2JJRp
J8NlXu2Hih79lgZiFDaxJPyDbLAEku8L1DLRYIETGFfGLezgxjpU8OmVC4lEBEE08jUdHWka8hmr
SqOAhHDUrCyRnhWbE2p4+H78bL526jIuXjrTT4U3mzWZvS6JPmb0ZKHbjKiPTPsiHyVau6HPiwT+
GjpwwgwwGQDO9DPlMS7L4d8b8jtFhXVoB4GlvYKgA8Qhbn47xIUg/Y6cIToXsOW2wgeIfNt1np/3
P0yamgDzuONVxfrZjOEeN73k4bUF5MRUnMC1OocXrx+alZwaBDKqnCxCNFd7NII1pjDhRlW1NwTJ
X8mJf8jZeZrMxDWHJCUp/auxQQOPy0/sBCr3a1B/IUcqc3CDFll/7vXIcJh/Xv1rsYHy5bYuwMdh
qHUjh8j05Z1EBROBikGinViyphNTTolXTLSTK++x2OmbLKN4BMltmfBWRvIjmdFpWjoJQEwyD0Ov
5AM4KX27BSjx7aOEC/K4lbs4KPEaBaVRNPRxPr2nDSmAMRoC2S41HbqXnt/iKOuhjPurLjFw55EJ
vzXG11/6T//qN3HufyVC4IrQJU/fJq1kokQjInAL5GsJjYZL+DgUzg3X2MMCxkITjjOpLbaRXIDy
ZOp6NVEq2XdknWCiS1Qwqgu/LVS1o00GR9irRkFIxasf97q05BEmn6UkLj+HXAmbBDsy7jpZgoz+
Jx0JtgO+5KvZX9Xd4wO0uO4TAPHvSerNzOG6W4x8Y3rYeDTFzPaf4qwA+N7j//dFMhlLyEaIKbfe
V/Gpy38I7KRNUXEnVUJMXSX7o8z9VAeBzj8sQy0lSdJM2L1DO6xZ5EL6hjW8RPm9iHE5aiw81fuw
3uWRCZGjdYqLOJf5GCTLTTfheaBiTFExIToCd5jdZR6pr2btahDk26QLI4miHS5FhsKx9/gqulP1
cymAMyc5uesqbcpKODjPYnr1ML9etlHXj/9IxTLyfzpgXodhn0On2+RzyLnrYohhF4FI2cw1aihV
GSpO8bZKyU3ijhoysg7j3ryrshKvHDMZgxKS1PZl2lESySOSe4jejxWHGJ2PrkJtKBnC2Rg9hzRw
UapgahwyvUm+BVKmiWREXjrrKQo0zGLQK6cvcLN8TRF5ydepee750CBo7nA2ssZTI9gVHHhXWUzN
f3NI4UUUtOo2Os7j1CNDpwQCIOsPC3BlrWw2PSWVXQUxVpmu9uXblHamai60mtu+oI5Zh5Ir14uI
cwutal9qKp3PTXmFZe00OPr3uQwlD2nUjDxo5MIwmpaAwgoe42KSNv43tuwQdN6WMDxTdkLuCiOM
oT6j80BVvrZAsD+eza3tzqilPbD8PL7bqphXncQAkGimOXP7ZLHsxMz4FIPxN0Q7kQOECK0gqUga
9Uo2Uc+g2+rd+oCQ8OCanP3k8YIR0oPMQWCmyfBe4PCXx+qjhVH7XoAETwWbF9dsu0EGbkWoD4Dw
hozFNbcnJai0vEbnF1zuTSbksn4SDWVxx2kwOifivCcagenALGVDzMo9OKPfEbmeIf2jMK8mD+PZ
X05E01FyT5QJWbKrgmDO1sxcDb49othjfIrEn9Cg8onaAWNwMnjCT5W1+qjWj5eUrdbWU5BI9Xxp
b5RhwXMPHwXu22VTzUYotKfcHvs1FA+fz2RCrLrQ2RrC+WVljXdsm+geatCZZddtdl6RWKvi3qru
0oFSxJe/BnmcQVI13JmAHgc9v4W8w8IY4FhaxFS1nIEDXac1edWsf9KvbTGi5rSjPmYDgZEaAfcR
SqKk9FYUN+z/KeV0vkaMil84PZOPymg2hoRM6HhO9tt1y3bvaFBGKRmm6tfYtRZKFozProUdvNbl
jjotjdagkI8x7VghTCfFiDaGTD2v0RmyTooMJdPMLW1ROAB2EJYaxzQQrBrwmUSGPUMmjz+TTBmQ
vmKmSF00AYX43SWbX1EqRaQXSnlUo5bVhgdKPKqgqrgY5fXYsiwaxvVnYEMm+XJNhvD1I+D+7ZWv
4oD7Eh/msbmJstN1JRmjW2+ceq7+w1gmtAC3HTB5jD9jclfp9MqavtNsSoWVrPZ/XYcI6i6etm5v
LxUvIF+LfFMr+BSpst288nvmJ1JkvkTg2/mbrRBWKgjn/Hi0faLPfdDc1m7ESwy1X8Bo3dPrv+k0
bqlTPkTTLHw1Wr3yuUksWw3sWQym122ZpSK38ByJjN9OfuNnMxaHpzoKLmxJeg8GTmB2Qu1vxjpp
0on6MkFdtTtYmRbE4o49lVrdXeMnQj+TvAM/gbyWOxt8T56C98pqGY+PrDsloMMMJJN2v0PslQyo
utVvaCaHGgQFJm8biQlaBEgAzPwf7/F7Wx0jZ9z++SrVrMztoKDU66q9ELouHe0I9icigS7Uy20B
r4a80VeH1mtsqDcOnzoYBNBvj5rALNvLqXqLXkBJ0hUpnCAoxkrcc+hvKT7E738qSKkTCIUp+NOd
lIhND36X2wq1TpfE2YVtTc41t2qX7c2AS3SlHpyIMJGhgzhjFPJYlcd97IaqGQCq0TrdrOky0uCO
0grvaBVT8p0h4MyJ24swDneqYU5q2R24FSjK0XAYuVxSoIV5kveO5/vsCmrkIg8E3EGIcl6QnQfJ
hNKEaLTyxzkf635rroaThI3Zz2HS1AjGnf7lQyqepKcT3F18nn5Y76eXSxX8K73E3HveZws1yF6T
idXE8R4rJsWT7cWh8ZDn9HzHWKhxTrmFTfiU1tSn74ITPbCCEA4yhpgmqXrhkgTRb0e2ljlnzWY8
JxXsNU2WU383H0plDG3LD+NgVmJ7tZ0hqJbxnu/sMJLCorFEm4txUULV9RMSwliMzvqU6FBvutIQ
GK8KRu+rLvXuLsQmqJDs1gtD+nfVOEcTh8P4DCdI5nMom5M2gm0hZcHlQcPhHdg8m0YfqTjG0hGJ
pqyvpePO/d3NIzcFnXG67oGHWFk4z3ginNbUw+2cV1Ebeb0D/paLWd2Vww6LE3zOEUXs7dg/I3OE
ErMmw8hpvKWprZAbMbvckzUslaejoUTmoohMOFcEgUzj4k2b3ukY7XC4oBrI0J94w2wQdY0Gyqbk
k9FLBTv1AI2IZpLa/kc0jbaLOTQik5+d0KwO3Sg/WFhgwLBpDgIxeLsk30ahwljLk5+u3hRkjPY8
N8mBuRYNum/EmU5a2x1ydzGZqM1Hg3AN9rrtkSRbBFvGjhbZQqp1t+T09e9dSXw2tFHFg0f6CSyy
uEkjYhXOUQ4Smgl2dSRlbxeBsfGdMFKe+JWK/BAFZC5O5YkQZpakWVu5KoJPPyTxF3qAaiftV0uC
GLLaFgzJcDiR7+W+RWlD9BZtGzKegkghxA0v2Z4Fppzs5NDnOFagFW+VOOwNQLEA8oF3SASQtS48
B4ZkFmuDrycR8RU+02WDQtTIcJB3LQ/YsUcL4QyAqSzPDe1/M3PmcYQ9fsEozeQrVch8BnhbybAu
LRSV6Bp4do16QkNADnfmVNLLjHBlhpeMMxxAPZqzyhGbmg/UP4/dOYpDQW9nB1jHhY40LVLGDK7k
X7LLF8BciPJ9zQwQ8NG370fYq0HueLTELfTf/vE1hyymuScRjprgcNzPZN9SyCfwC6AQKcW06oj+
lDuUgf+MuXAqGaJiQP0fh9/4S7ZVf1NrkWnB17siybQ7PmtD6zNeOSXqqeY6m55idOYde2EW8Mtj
mblgn1SL781tSuuYDhm/JZ91vJ1G10w+xBMau6GrkGkpwEk6TK7vueRioEpmkWfQqWKsCffkJT+4
k7+pwKogqZlJyzDQ8zQuTNf/wM8YWMgzH5FtW4UCHYmuOq/GMogm3TKDBYuNaVDjwtcpEeGy2Dnb
+Mf+AUtK+vKDcgncLe6RRAJrxpeByMuGAWBTicCBlfYvPNNnjv+Zm27dOaZUNw6yYN/zVXZWCOP1
MBNhFPW6ffm8/cJbe7KyG8IFuSprfcy3kyZDADsm1FcnfJso+5IQGvZnj0ycmyiggrnJ8zq/mSSN
ePrObxtKyBvATj3ZZ/MX2WUxCJkDbnHs5q3oyF9XP+xD364UmhnFxvbbY7mBx3SyVSWKMCK/nqBK
ASRK99l+RxaHD0hyrg5G6QdRRUBlLoV7shEyOdTlmLFUjQJWhnvaPIKXJk+TDWFQqcLPDj99sXwM
foTuxEY0qjbuxNM8GjhAdQoB6uM17aY3kLyYLQpmn2wU/T37Lvo7ZYTl6CgR2+qKFx50WgBsH6fh
32pg1SnB+RA80AEmY+OPJgCCafq6UH7m71GHZtj63z/cx8TJrEiIR2fZvSTvOSlBuJEZvCTrkv1k
pYIqxVShpb9kYraXYGIl0Zze1GRNSWQqRIkjTyM04fiaVLU4CTfuJdM1piJxUuKoOhDique1bkF4
lXMYw+XT5Rr1CuUmUIvqAx/3dzBTLkVhyP7bXNIHZjvYtaYFp2HkTHwDY0dedrwhvDFnshtM5UHb
ZFNX1fWF7ZZyROE/lpbwMp451pZrCTYZWxYqdYYRpuO1kITInrnPHpXW9p5+pA53MvXaBztDZW9b
aFNA47Xcngq0xoWy5w/t91z2hJyUOzDpUQH+pHn9mmiBPsTUvkaGx0nL93kBDgp0SdpcjBcUX1eB
4oBWBRSSXJEEo8QJFF2HZ6XKoscpXJ/FKtc8IFb+May1PrX5j4rkEyEliVwtldjpQ/yV+eHMn2OS
XfyeT5hxPpQUjAutcElRD7wu0z2p16NC21ijIyu1sShiMI2NQLLevQDSedWIX6dYYF1T/V8DIEe5
tm3YfzsXsZsV8/CAJUuIQIIKQW8fLzwEb2S4o5Ob8WvBanFuZe85t/38ZTTh1+ajUEVrSTYc7uA6
n1FKiM3x3bIy/mWEnXsS7Jj7QKQmmYDo1ZH8pzEc5ZEo4cRmbMY4FjU2qPOEGhKaynVGTCokqGtc
vWIfgHG1SJrZnKjFcEgytcyGfNCBT78nH6YrWTkvsjuT3naENAUjrL3PXlS4GmENsEJ6+YO8K3eA
cdEmUoNs0U/FTh+jrgP2igTnBOAhvksshOP4qDwbaGHarZTrdcqhFLRAbrYpg1D5LntaCg+udR17
dpihg09sF9mRWEhOm1dShYk+p6oJfPbB6O1U2wNvTb147fh+gooJOnRJVgpnFEocNl87zdn5HG62
dgrIpVJ4HZLjMuMSYCVMQgSXOys3cyjSrA9PyOYcZnE9apy7Ya4lJeGiR8YoS9ow4DrEbPD6Ts3z
ibAPSBdeeujvXoX62OzPCOpXR4lKJTVyrDje5+2wtzSYKDZrh9YeKbVQj3+vODTgTLEd9SVvldpW
j72BXg0e6S+SzMN0kyqYBekk++1+OqIpGmJ0bxOLBtjVLFfUUazlC9zHikCLseGV3BPqQpX6qbYz
IoOKQlqVHTYjJr6I2gbxCUDmcc34G7uc2wpWlRHTdgneSy/yr0Q+WSHyzGcSudtQSbSlkKNojPXj
zQimSvH3zWDFAzuoOz56kWThErBvVRCS3R610ob5yLy4wRJkHj9dyQDq9P+zox8Z0bOSL77AjjC6
f3kBe0YrPgXE7A5wM3j7ld/GLc8qCKuWpXo+/3MhFCMLQdfQS8QilhmxdBQPdg9eYbqL3UCfChF4
zUmH6wyJR+Ps4ct2UAx7FLBupFtlfIMWZy3fvdUkxY55ow9X+gNCeQfnNcWwTCNEuSQ+Y/cNh/YF
JpSe87lrajOKhepzqmavJ7L4kYbuU4yE/RaHnirPNWYDk1gDp2oxJTFvzgLE2vdR0pKnCQYW1uq0
SGJwp7K+EWBs1klY9PPmeijQtnMy9bh1cfNEZwnEXrAXbFQHIceDx1xEWcXieq7bSssSMYVNPzlJ
0ZQzamH0cNh4zCNjMDSLhmEztE+APGwMCTj59SyIVLG8xojEEeXz42hSBIRae7qLV9eHv5vvSGkB
wju61GTCPWUEqrpt1PMasFh65+szTKqQB2y5e3pnmv0EkLDgCPsg0eeZkUtSErnHeZLBChxABOQ3
aYwo7KMgi+t27UnDlaOm/cEFgm/heEZ4+4gF9lnG5CgNWkRavZZOAayrA1aR7n0GXyJYfoHsr1I+
Y1njYQ4cTYR9J2RVHtlvDI7+7mthPL9ujwV1ZHJKOvmhzFMZ8w3wfXoIn4W5EuEk+cyhGaLXu+4r
ut1eoMhhxbI4sikB8tsTJfhx6mXLnQdH3idsNYG50Ix4VxPJGb+Dq0u2ynW9B/nPpygjx183wxQ/
wdvUFb50eVMeYU8YiITGVSsTESRsj9punqDDsMoUJS3qE4Nk5tmBRrhMmRcGuRHLqIgyjK+HaEsm
9yDRD3Oa/cH2i99VuoWx3obTw3h1n6Up0yoj7O2+AELmzzkGOhbRpnrRw+2rUGUyHESO0ufuG3qX
ZLlf39he5J0lyCJctpeAKSVB5htwbbDHxN2lrQ2XMyTN3BkwEj7AtQCC51U/f+O83wrYfCjr5zTt
kDOloKtWYp1G2G+vtW+hOnWK7NERy+Ell/b2mqK7Ml2qZRiidG1l/Bd5xbtvhC24DRNp9sYnc9tx
BhtmkqWw1APSUX6JeGHDJw7ogss9uJDsFlvzHrCyPBLEMN9SwiRABbFK+PzvF6jN6ZJJMsPXDHPR
E4eo6NciOMJ92jnLKtIz+GJOpWqBf5a11SHIl/+kj5VF/b0+2u0Tql5x21Nog3h4BUx5viIuXQWJ
iQpi+BrPiC3XT3CJ4oKxX1cuHfYViravodZ211rLe4TQq5idNy6KgY+HaCN1k1R100EcpRsAqZEW
Ke/Nl/pGKBxkkytmJbbTPpCeqq383jou0s6gtsKRDjDAYNhob5nRp/FG8Fs9i71zipoUC5oNg679
baqyTU4a5JlOk9cXrv98XlsRCqBR4VzuGYD2omcJztEGQ5fVLw/iAU3AL6JUdd1ZmJS5+HQnq2mR
zocKU7F/GBKPdvUtCpny+rI93vrTKYFwdPNh6mXictPT20s4pruDYhiD/o6r2D7kKrs14hpko6as
TiHmjnKLdbZKN7G3dyuqMZvyKTZ1eOktsXZ0OlrazoSHH3VCUpfdFR4LtEBtLTF/V/eL2CS/LBKa
lZL533YC9DEWwvTgT/3K0RJKlo1lFAysRhg3S0bqIruvr/ecrTwd2k7lM34svLZpd9rvEN9b+bT6
N4xDRjvasf/rXRkg/8MH8KmHYYHGQtZQMdhytT3xT3VuXZKXFpbY8zjhpip8euBoBgneVULd3AM5
cMspjqxp4hlNZDRJoLPUbYEWS2duQJyl0I8+apvWB/ZfZxBjzEqx6n1CjvnCdkGC+Nx//mVBUlB+
a2Isvww7nOb7Fs4tjaVcIK94u7EOmCrYpElU+9i0xM9ZZ/ueX+OS6G3C1/E9+9DRvIc6syt3gQdt
yG4GmFuyIQo6f75uwLluTAFRcAL3FJqoZKr3kXDpm7rUpNjK2VCpuD7QF/bNIWQCAuwuc7Jl+MlY
3SNQqWGpm9T7hRWMmVY6lx6EUDX08r5+B2Nq643N9dr3u6dr3FLE6fv13VxVYQeD5CPLGtkuhM5s
UKzqdRr3Lgf4/pb+L2aP5Xh2zK/A0DHsjAOu1M+4nz/VSGeuUSnT90CyBmTAuppkB+b3mjCyHXyz
Q6AMQZnq+BjCW6RvTOyF5Ahz3qaIKSwCdD6BApZA6y/08wvJIkT/IbfF2bc4O6VkCIPhzeD5sBV+
ajElrGbFQk5qcClmah/U3BqpjcJm4aR+Fc6lWpNBdlWwLQCgUZCzHXyA7vF3EJcnneCu3InM8V2Z
jf1i1lmQwpIsA6GVrJ+GVGl90xE//Yi3o5VbmllbuEYDLioByw2dOVKyZiFp4TliO9//dSn8EVIn
ZBwDHNOC6+DFTag7o4V83LBJOhJZENgV9rloIwxUZDRz+dzGnXGurhMB4ZXFJnw9vCNONhxuVujs
Ilcz4S7AYTIG4HTQzA48k1lkK4qrGMTBYM38WAxyEOaE6GKkqvXSuNk1LYRoKR8u/OQeywP1/lpo
9zs1cDmak3NpXyQgGkCJVgA9AHlLOfFFlBVpydZDy726NmQIKWCdHgYHY0d+53aGwetF+bYiEAUL
UnPAOH0PSL+DEvPqmcItlRDYdi8klRCM1anG4imoJcYxrdlC8JeXqTSyF1GqojZ0YTADwwAZHn6R
mSLCNt853MVNc9ZNrsjQrk6B/TyBOU7VPlyNUZWIDXKd6wyWbQwplHx97+RBDdO/7uMAMr5nhF1V
kPzfUiF/DxaKlB0Te8+okVFg1ddu0fap3rAHJKRBHPGxj+Va9URUF7FTU1G3vp+5Y/8GNtf53rtV
W3PiHeg1BCPC7/9gpodwVk5bt6LC8tXUqf/Gx1R8goEZhT1kaHLi8FfaV2+4onnfRJuRpAbRcuUd
RFJjSB8OFmR1po+dCGxtiUfmAGhkrncfYFMA/Sumf7GaiQOVvVPlI6jtwoC9/cmB19dhSXjqB773
T6kwivi8fZ1puaghrgeOAtzF5w/KKcPBlZ093SMdyPqJcyaFxKUsyrvzCWIp7B0+wp5iXzh5S1Ek
7lEFZ3PhcR/AcT6kcvCEqQjRzAYgiKvdBD3S6bG6cOzrSmmdeGGxLgq19mf64I0Ci3ZbKBUJ8wv8
8BC//U5aJg94Ep2N/vKLrjdlrL7VbSjXA7SvaO9vm+Qj7pyDCPEqRBmvOWX4YfU2g426CmDOkMAO
mwwpjzCwf+wB0rc/uxnoHNjYOzyaKRRo6XFiSL/T83cu6jOkIGuGX0zI6fGJ9PTCZam/MMHBAPi3
XWkP0WkJHD+1znathcY9dGWpW2xEAfKMl2rEjXbQhj1w05MpFAP2L2acAd15yEGmXq2a5G5l98dv
om+q6EhM0orGdwcdy1Kh7dfOcLF+lisUPiNGaXxF5qQnES+M2RC/QNculucpTOGfbvs35/LZSwlg
btcTGntE9CS3o/FijxPnz855A2nJxbVs3Abn97JbqFdW4Tdcxl+h81GWKgHbwbNJueEyX1K4G+K6
mdekAQykntZ7pkGKWkV865T7TxqgMwKwtPdBgj7l1xFmiLFWXMJWN1KKhI6EopkkMDkjizo/emd1
e72vlPjXlABL5hYM5TPcj9wKeSaHcZAQWUBtj69fkfztQzeFRrmNjxIdKtJ1B21bXZzJFF2KKC+x
YQh5n7wX3TXkFWhfODAmfplqTsKXA/4Zx/eq9jIYjmFrBEyEWlytVZtFV6bS8hIxOUWJQRekOfrM
GNYpB7jDqcUR/zzyz6BNt+VtpYofaNgeZ0YG0QSAykb9HvHFRV5fQVbsTjakIfw+OMDoNrLWvXTH
tTSiJseYW9kFnaDNBL1eZ5AwmzFEhh57XzrZTjbiRZ0cySCfboq+4UtovBCnlQcUD4gn3Th3SYdX
WIgNfRLnXxIFSRy73QvzdFk1q8YdTkrNnFz95y9LW0z7kxVGaiatnN6Kwl/Cec85JJNy2pVDXXYq
K10lrMpnd1Fs/HJUy1AG2GPPtczV8yIDbrUUb2x1iQySrG6GoTlJCc8s5Ix3qXmGBdP0X/cQ03zq
qJ/6il+wK/AmFlIOEUkoVyE+SBlvyWuqEZRWJXoT4INPUTOJ/J+63VdYa8IzUJGJ00NqyUtRQLCs
Cpqw7CgDkCBIyUyFUJRoTWPDciDyt6bQTxwHYLNLOYIGRJ+OJ54kL7bb9rGKeivtWkijXDw9j4gk
kG9WHrGmuN9g5n6Q6Bud97njD54MVcEBkRAd0dzF0Iy3VKvcdpKMDMJUzESuwtccQ6p16DEk7W86
Qjket3EWMPDcLtgzXxvOSUlt/Z6uF5HbcWByh6vDmpU4PorPdrNFsqjsxsyIAp5MvC9m/1U6VL91
jAbRLvPGuIUpuiJkM0SYcv0a+C2rQHA4VtyU/kVelBqGTBNOGFNA0cxdJi+a/sKPpXDp2Wi4jOFh
KZitJRPQ+Pb5v6CDwZn6CPL1+Dvl1BW7jKaD8Pg9FsA8QpCWb3+mapNWu2Qptl5I5PvKlrlp37Cv
732kBotuuatyf0kyi8gC9E59YxqaQ/SohagfI3IAUPJ4BpTmvcRj0VYDVyM40xenOJmWjIRJXsxQ
nEWXlW6Lx2y7LjTGHmacYeHQ3GcOsnHcH2UOjfZcIREox9A6E+mY/e6b5LKTvsaHoqrhTLJxGRLj
sdDkGqa7gxiMNQ4LfN7JCustE5MoI/s+107ewdftSpjUhT6ke8J/ttlIaQxCMsl+blWoAVzHLCEX
7YemAHcLZU3Oz09Y9pntprBWggav8oZaxZTXYWq3sNMnsdiM0TyY0XhDBontJbppa38JHRWWYogh
K8Lsi2E2Cu6V3+VzocBWZm6RYZsOtoruvZe9Z4s2MNEx5Z1J0EDPyikETHuwfNv4JRajtqzUKiKK
5tSRJL/PlN61gttuofDmYllIXQIkQLxBTrNwpp74upK8jSfhLfdo4FG2iSk1Pw67GHfiSxUarNI0
qzobRy/MzV3Zzl6nnfVGb0wTV33lNUYIAVRH7YkN6PK9EGe7uNpqAGU5PqWXmfq1IqE9gsQ1wpup
Lbms3Hh0cMRlKPigMf2vszR1djm0YedwFqk+JQWwLlzhJQWgPYqvD7tPjt2PkFaMb/H8GeQoYe2s
X25eH3Cc8IhaBx62AMz8yk6N6MSyOWtHIfxas0G7DUmbZkEE0nIlVvOotN69XffDd2Eny/d17Cra
piDp5ZTgl86Wt6Vg6EmhcSHwsNdf8dt4dcCCbWNfowxyJrkazVS8pvbEd8PhafOQhWg/VBtMNUso
DHmkUA8RFvgCYWlP3jgUkCp7085eERSn6DwpgsodRcLlIOGmXYYYAfHSZZC59RIbNHOmOXgh8D3h
2JU+5p2qUsBEj8DNdbzEK+m1NyzRQgV3wQ4+TLlkPlPsnxGtBiqaUJjWnCEQ1Cv3WEpq6WJPy20k
RXZfcLUuwBus1ZUsQFzdrGV9BaTprNSIZIEZlEoRcJUGhh+eFyOt2KWwzZ5vVLuuevP91tJMA39O
A7n4Gla2UmlhC8u9D1NBlNJ3kXTTkLCBAjKGZhtlLE2NrZH3q8CoCUrl94eWoEsyGNvWgneBEQ6S
pGa8LhmrEudJG9sdPnQTbN8Dbg9CJJ7txsB8WpKBCqKPKiib19b8hdNCoh2+2mEw4UP2LmmLLGU9
Ob2/M5VFQrVZviqkYYgNG5Ce/c4phMA4IH6XGsEGXRA4StteKUwZhEBubtG65B/6dH+KeADWHvvt
bs/3frX4R614pPyMSV7sxi9bleMJmlaWTg5Mqi0CbSCYqIKfs1A91ZVV+iV8IZ3/jEZJbSMsAUGg
YJ2EdaVncma9P3Dmy0BCoLXYR6hSPTzrLRE6SGbWWkQKmMnI52kYavAsO9DBChs4lsCA9se1jU9l
lIzSH+eu3O2ubj1H998y53ygYINUjRO54vCZiEtXnDmX4Sn4kk2YxT7LqeWdfHXhTqAJFxG1ko89
jzHXOpXhRBOj392ioa8qZXQqr1Q37u+UGynhmx0Ner1vpD9tC15agPYPjGIdi/EIVokATlzSMP5U
DOO/oXnbeOG75Bbkn7/s15Ue2gYseZAdk3jBWqcFrHWbn+iNQb+DHioMbjlFqbHdCWN+t9UxMa7K
iC3JQC02aI4SAnBEocIJQw9U27ZYeGhDR/3e4E5SSqBlsAip7x7RP3tL5sJRh2ycpYreGMA+Ja/L
S2dE6DCgd+w96VJgqnaCdllFu9lpoZj3WuH4fUjUNVz8hIsre9ds76v72jLONmMbQJKi4ypBc2sv
oO+cZ338PyFqqpKC0IHZdhTkyFDl2sBA70LBwkrOVhL64/jpr+P4rtwuV6qZ6b/kLJCmccb5bXQl
dAM1dD3+ca/iMxbL14WiN0xZlEgbc9BibdmmZ4wH5kQrIIj3psEbN/pceY7sXLkJUPmRu73BvIbB
awYlORGut1VHMCq7xYuFsgXwmuT1eQTNklvKP5WJ9fEF//9hi0ysXLV8O0XdajFuBdZfsm3CRxN2
zar+DQYd4tIfyxShiUSKlokaVNxDiFXCccR7A3Sz8iOF+qyq83u6NdLuDC3NQ6qoR76rVv7xBGlC
6ZJssulrEIsN5aKTbmi1enYZjTNq/GgJ0U3zT0BGqfA9hbr9yijLlr+VeLldvsItpu2IRYJ9rEG4
rFBOOg0ARnmPp7BRKpuvhZk2o0y84h6JPt+mA+itNETbj/fkGHtQWmc4u2HI/rkCA6itqKGwubyF
11cvC1bPq1KoBZjmmVwFjrRIbHMVLjPsFmPTzWxhk1zOOr8OseMujZ6b3QLNJSPXTSBc3ZKQ9+OI
5Dz/plS4GKcejMTyou2zUMSqSrqZ9nNE4JGtGt/tsgp/LArj5cBXtmSiJWq6qHZ/kBG8dcPo0qY6
RLLWF9a920X4U5yuRFussGJ5rgjpbqEsvD76wrRusv/j3399R3PWZM+FcspswNZMDOkfs6gdjDEI
E8GmmrFw6bl0FCxywp6Yr2FntucDo7OBBY1CgFtgkvAf2vEhLQ9XcS7r9oVwUOdX734Xm5D5CWn6
HU7nDjR2nTIw0rv6Llp3njPaSj343/bx3/TFJSBR4Vu6OkkkWplPhdb7pEN1YLaRatq44RGFjiLY
kZdC4KsRygcqEyR0UJu5kBOrZ6m8whK0Iv71j8+XSAcGrAArdXMlNdgdujAc0DmqZ+4fHPfYmBAH
Cds2eNG4u6szbzwrlea5TGzN99jno6VzS1EsV9X9+MOUGXWRv2Y5KeYbdibR0kUfg/f4KD1b90/9
C9Q0j0C5G9eD0WFt73w11gCJfxuvwoXuVesEtr4xebqE8ql+EYY/L4GMnLwtyKfnPKqFlZfAHABv
6Sx5XNpVafyZ8LATDlT1IDN2M1LP8tZyAYY3n2KxJZWCA+xj/hD10JioVG200513TDrep+5B2HMn
/t01FPeWY45+dRJLQ1Iifq8LmfGCtif4Pvu6qZ6abDU+kuNWwe2y4zHqK1kvLiFLrbIq6l3eBNYh
/v39flwK8L/FLX/1UTp/wwtKarZJQ0xRnlPded22p4l2ant6DK6s/1CwR5DX4VNlXWLGse6hq4bb
jk4ZKliBJ+1MSIQzSvzlwEHvfL6CjTUtZDE2f0ySQ5nu8BZbKQG2KLMke9+hxwInHBUaj6ldSHf/
3o+kN75xyGyPlyvQIxB2dUqLIdyI4G+48Fzo/c6wuNF9ceekZNbUZrmKIAiRp7Ae/gkaKXUpQjF1
WOYn7PE6ii9cjQ56bga4O+WfGSy7ql795AEHQys0bZrqs8rOg9rr7GbMf7vRz3gTG3l3oAomgfND
6CR0r8JYcFlkVBZz+T9fOLBv8w1cTguoWzTr9rKajJDpZhKpLRuGLvU8x8LfbXgicNpMaKDH/ALO
nIFDSojiW1QqYOCLL1otyHzVmbttVJJ73ViPMDfEdpNA3KJlJXFcyzNliw3Yl8ZpbfBNBp432Vy7
Ilv/e6txPldMo2XCxSbTGMhL7c+G5EZfyPw/w9aN/FtLSavEpkttK4A32g3YTZNxFicogOLc7TnJ
A+FB6d1jIAy708u5Bt1psWHlkJOT9eTE5qxPtXu0x/5vNqFJSsiF63P0vNykYuZhtT2P6nw6dzFz
pmIALKUQQPwk6v7tbBj/vgrJXHmeHPwGRnKk/1QmO3FE6YbKGOJc8UQuXHuRqE0O8/iA1/S7uAI6
32PTaMT4bhTgtJKef7ZqzmGgCLOpaPpwK8SjYTQ4Cjb/WooZqF+uxAeBJej9a0hN9M/DFPxbqBV4
E4guVQthgOKLVRohNNscAcw9i9pF7Rb8QdJ9/EZFstVUvvC5J1vm9XB/iFiIng3WX8v7dEKpkxKR
mqeyGyZ26vtOwHHIl3zErWm44gZ65SVTUl9eSAf1cD9hyIaysif0hbkAd1PNZ6zLNobYus4jWEhR
p5uDHGLQdiCJzrM3rljoGNsCWyWGbrrKwBl//ZNd2SW9EqTQrHdHL/pvobf2wfIzgvzWH6CPSSQZ
W0+9xfba6+pQoBksk1Wy3Ifwb4csi+K1AO9EQxpWlOiKinF19EtqprmlJ3AW0CPJGzXZh4nl+4Tb
XdMbQr7axKpu0+yWJ88ltORW5VtRlUD6omfzU6EGkXeV6YSuLFywGJue7xz84pFm0eN1ZLNURLJm
/RAQHNrXaJj6rJ5hofz0aLxGZKKlUDzuhm9vrIZgEKc4BkVsivUSey4kCCL1wmZovcaTV4xX1Lkk
fOMKDXVay91SquC3McNkRodSwwTHVyXJ9v9RoVkwCby24S9tHmetrZMwlYJYv9I9Hyc0RFSVSRVI
bdovuEOuTGvv9hRoCvqW/+NwPajCHRKFKcc4uERAoesFVbk/mXEeXwTyC+Ta+PyK8yqe//Yrplo6
706hmmZS0HFCZaZ8w0Mx5IfYF9XuP/e9NdBom85f41t9FPrchSTqkgW6ckmaYs+RJE3vIRGKvFy1
MUYxEr7lxpfncc0FB1J+/z14/ac9Ww06bCjr/NCn5JYeitFYY7N8CVvke2K/D7yvz0N+Xc/o/ZIT
W3eAwCdCPVKo3laTE2v4q5BQVoNA3fUZ7bPw0llfOjYC4wMKlTAVZyzcAwhI+uB36oO2vHL3CpK0
tX/kuH1UVTmkmDSFe/naTXnlCdz0HqQankDE8Hjoo8yDi7ePbzRIa1k/w7PwJvgKcrEG+9toiUTz
7C4Glk8VVFvBpuMYByBWoI7naLGIZiAEePoCdE+hDU0LADEzTNQ7SgAZ9St+vkXFk7piP//o2Skq
m0GvYr4teJ4/+d4PCsNCWBL7+g7S5/QdbJKqC6Quu/fqEsaOeKL5VPJx2XQUheN4ogpcnMPbeZlB
xHLRjkslr/o908NjMRhUEEE5YO4j9B4Lp7fuSWHWpidAUAyDiEJCe2vtSAthBUCZ9WDvf0XEQP4/
QRxYjbXzfJXT5Frv+36XqOU1VXVB59fcqFCnceyrRnGu8RQWG1j+CEy06xx2+eiwdKUxTjuzaMw/
PHbdyJc9BzoR6VKH3dryEWXE4ySqWR3AEpk/XwiysRXKQN+sZA6Ds9zyMFZ0m9K0Oc9Tmw9YVCPZ
oDt+n7UtBrfmZDMl65N7hUei+00HS7LlOyx2Okajl76/IABa96K51HmcEGSBSLh1w/ynBXB2GalR
9G8/K280FBqBgFVKc/C7+nAh03IvrONHn/VJJSyX4vbMJDuTytBFdaT6hdfbe3h/Bmg+MCIDoa0p
HCoKU1O7XJ3L7VCWWjZfNYdBpRcfFBeODUBQlgevpttXSRcUsIbOEK/T3cdpERGduIlxKNqIzxAn
pI8+dIjr9na7SgLN+rSNm4UC/CHnqwxlQDsi1NHqy8b7P/DFh4fwLfHHD3IvPGjCwo1a1Jf+ryFC
BaIYtinSkNooc0TpwwMrLX2NDiGdOnSQc/3pXqN3yBkVROvmAD8h3WlhodnC2DhyrWscFoMMIHMl
Nqlz7yzhsmx4SaBWD7EZ3tuSdumXar8MuX80SG1ItsHUoHE7cVHVgUxu4Pnl4r+gKORws0Yl7JWQ
i5y/KnahofJgq74ezYKvrdmwAXj3z2YVMGmzDrwN4io0xOj4gmvDKg1aGrQjSly3CuxZruO4ZKiR
u+Y2x43lL+6GFCjuagfvRDL43RY6nMfM9Bbp2E2kqs2qzuQDUwIbUC9VTz+EnBA8lHh1LBS3b9XC
94N/t1rE2DZZ6R2XIWy0OBXd7blN1qR2PhhxLrkLi5QMnjQyMuObv80m18IFgpLzOR8FuLWI6KVq
pu7Py5GhgMFnQxM6WOJJ/xVq/82mlNBACqwjjQtzq+yznG7FtYdxaEn4ka3VFVoYAJ4cRRqM6WUw
DTFlAf8053MRc11YNYxw6mSA2+9aUcNffiLqY4+Z2nKvPNqGwWO/oPPog3SQ1sXWrKJSOCP5CblK
G4IF6OkiTwOiqKQ5aZt7MLFvzWQT7ehWJB3PLTgC+mkIHdJROj0YdnqStfYuQUI8ezmTnKdupdkk
t2c2eFPlG6ifV1pkfN0FTtmzYzcsx6QZRTyrCgXLGbtysXALuSwsr40Hdb3W3st/uUPnTIJQfA5p
rjZqAMyCzYmIZuu+ylOE1GCBcx3G1m2hNTLpAJGvKbLRRix9Jg6WEfK1XY34SXGk7+yOk+JijmKB
X2ORuzDuOQ6vRFM1O+YDYNc1mhw3EqsxuMexqWlPSoT8Lm/XOy6zv36KJf8T/zoiFh/XI/LFNJS8
hxUw6tGGwfH4HTwTef7CawKuiy2cxjlsEOfXyaLZjjNG/V3LLqnEVIa1Gr5cnXXIaGIzTKn+VN/6
mpHXm1n5QZMlWvLzgpHtgRFzqlEDXqDgn65YLxEYL14zaxOV1S0/+Z6wFcASmTGO/pvNU5J5y5xw
AxQl/QYCtvHJg8JlE+y3XMlTn4kXBcssqx1kFC3RR7FtibC5F1B5lmOFxiFAp+wEjFgPwkngd3rB
akFhLNAUxFs8G3NIqrAFtAkEGgocSlTMTGGPLnfkYsvMHRirllOdQbGSCcs2OkNQq4iJIazbGtlg
Rcfu45tx5d6j0NnH++fCRsbFTqI6+fh+WXFNJUJKWEnjgfoWxSyjAAJiQfolLvtMSD05opQbBZVz
1oNvNv9cJEesP8nZHuXsvyLW+AlFdegmIBdQwlr7wIJ3UvtkEnBDR4BChUj66p1Ki137tFRSG4Lu
Lx83Y8f9sPhvRqzGnBLJJzoWnjd+YtGiCIVuFa18I9D/yMUVUdEbSxS1RTOoC5oXqHjqsFoIvicf
hKozRdaTHxRLysnPfUsoHZFJWzbcvTF1ffkZJiDkC4vMBDMP+xi8Cye3HWZLgKyNi8lqiJcpuNfe
wqSkYwPtZzHxHK8gZTMUWotn0Pyw0UIaDh44mqki7PozaLGGZEZLyx+unQIasPUz27Fx6XV8xkmP
3YoQa4TK1OHE+04j1WWsMx0Wh3vqjuwz34XhFpYwQDQUETLBU3TJfRJJ9UbDgZ+lIzV2qamCK7IB
xxsPBeWOEKHAUpzT+iCHYy70mD39vgR6yhWqtnfUSqulk/rS2pU5TNd9FxsD+WPwGDTtKWfwAsEJ
qfGvnKileK5QkRkZ0BYWMsFgaUkxJohmoC3hKl0bVlJbxzMeUhnT/C25bDgRBSmi7XsICdHGJb3Y
V0PgRRUt8FA0/PkdQatqjnHEzQoWooIx054uCHFKdHobwTtyYeWihqHl43NHTqnb5m8nG5i78JmV
cxKspYL8f4TuBNSFD8i4Dx/uNxSKbR1/iizosaS5Nq9yLnqIn367LfwR9q6AnQxiaXRIB+4RxEXm
838ZVVETZUofCbMd3nBaUVWP4zTDJrmlj1kf2UNR0CFRUpE/8psHT+LwL69fcCg0dBPYMd3+2S8G
FCKgZlbc9NAzBHc+kDf5Ep3Tl9EUIPIyQBFKgDMl9Zx3t2M/fPrIwENW5u3+QNPdFJDqEdgJAp/L
S3qoyAgMCoTdRs+fnObxsJPa+5kJbZdvU5DEqWyBpUW9d3vKb1+iyfis014LSZoksIYlYUFBX8YI
O7c9/TkUxjkcVO8s34PgiLQfLEcC5XIS/JZkoFsiWJ0aS/pX/YbNo2LiuaqtxFVszAXGgiUvBJXo
alEokODn3Xp4rm121d4cpzygg2s2Yyo3Q13vz2c5o5yopWuu4GDQtAHRCop2lWVceL20AiY9Zk4Y
QymnrPyyQ9cqz111STPJK6l9dysDfJKej4WvdbKWsjKKMuf5yjTvMOy1znjJBsP7oVT4T55CWZx+
/tzw/hICaueww3F8Fn3rpkoR09kwoAzd7YldfKiAiX74OEiFXm1Lm0N4u8HKPueQIDY5btgwu2Di
4iAl6N3RKW+ye9lKOAa0rmiJIDAqUoqSKlsSXPZD9Yun5KloRhf9wuRkdrSCLi8MTETPeVm+CI/R
9hId6x7qvIAzncbI6wpljcCD71+b2Pa67skHOm7SzT911xO6VQfWmFsvPS9dNx5IPOk2o23J7W4T
tAojGAbxbSAyc3/pQYANHYSI/zcqCbkYMKGxdQOkthyZ4M0Db4cBW0kcCcT/W95oVUvLfzC0dwS1
zL0GV4K099u//GmLrG4cjyDeT5KyyWBQoGaPnz3sJNh3FcaMtTCJ6HH+1TGFOJSf0uzt8/jFsxOQ
4plStben2wTgeP5+2Xtbfwn3askAbGbAMb6WOZPP7sW6Tqg1ER0ujposzTqj1J6Dgg6Ixd6Hf1J2
aO3kH1RzZFo7jZeaZll8Z3cI+U02Z+4zvpov1U6wSkgYuxOmp9QZvdoAoRMqB4mQ1YjpE17ndKa+
smXqWwF3vine7c/BnnGwVaGgBUcYN9gCZiGiKgmkR4wsqz1RTDUGJQlqttCJrP2RpCY29JB0VLWV
0ydMnYvjZiUcmI73Na/9tSu000JM2NBzMOC7lmfZtbs9sirUehsplKtBlMKQHiypmkDl8FXHXLEn
TcW9bxdTlRtP2C0FJt0yH6hfkcepA/Jqm2rRQtx+VCrlzh5El95469GJqY4MJzPAhzvbeqD9wrLq
aA490xQMxXueoJjT45z5O8iiZYRD7sOZ4q2QmgRXWdxnivUCK8DsFvV4DIXhDt+MGaYCRIiE5Wzx
wBJUstlRhnSNFGuya6End0cT0Z6y0wnY46H2d4Ev48tP7JgCReLoIONbmGcRh5x+fmso6c7KIcKJ
Hgd0ldlcsZ5FO9cQZcJdYyzp1nNZbjtUbH6Ee5f5nstCBWeQIieAYyFvsOlQTm8OIsB3UymTmARt
EIGFWKysuPrtVS0EfmfF+kMwuAunUDVZHhiKB9vM1qZoGfJqBbi0FWETIFTJD5oYuOBYtjvelv82
tttfDW8k6lZ0I3FNaofasnLWzZxEsxsRd7jb1Pu6YLBEexsp0sewYlftFsqkvSOLVNwmj6/zPTF7
DGQyM6+KC2HR3qspz4mQdYyWzF/53dy32OMyCqXSZYiRL5clBfkjr66sTEPib9WaXQeYZrWzULyS
eYpQsZR3E9ZwMej8VVoUEM0psnCICRfk0ikhpYD4riUr6oObqW+SoyBNEolEhEqu3kVB0io/CxE2
SiNC97VLB20B2Trf2Rfekuw974/+56ZBKJ/bAMf3q25CnNEYc0z4rI6flB7aljYXAtXA/pbvS9ro
Rp+dsM8knjOq8Jeswb/SkQIUdOyyq+yg8m/Gd/pAgpDqEOIZ1vLHZdfWpVusUVSPT2tmiy1gbOfN
v769F1RKZW2Z553hGdo4Z6G8DrI4yTfxk8TzzDtWA+IYKQLpYURNo4YPjJ6/CteNgCVpnSLaaBWK
SHYnZdwxfHxR/W7W90udkVoErNj2XigqqITgOo/ICE0Oosk0PU/36Qr/abHUi04AaqQv7/+IA775
VFckNwwdHx/lBwXpj/lwwB+/wG3xQShNA+XUt0n7pAIM8dLO77KPPotZLt9/moYP9d+HFdCIR62v
PW8C9Fz7mkC6JDOzo2eBV7AKQwZiAYRxzoa6nmAYXSAbaKVbuVQuxiPpy83Bno+4cMAtGT/WLCMw
m+qPIpwqvUD8jupUfQYYEX3oH22gu1toKli6qcwb8hCwD4pr9BLJ3Sp0mdOu8CHNYWDBS5tyCAN6
MaRbSiL6jp2VhE4AiIzn5oAuZxi7/oQCAQ9aYAbhEydY/LXFH/XNxz5yvNcN8CtQwc1ZF207VNoU
LbjMADGr/SQsQ+Mz9OGVV8wGoIMN3/w6BXjRSOhoyFfXOy/bYkLbLO1LuBLdHAIwQi49YFumfkbq
Fv9Cfrphx0cWD16clStdiflALEtSCpeRXoCcoKKVScijULZ+qvkXjl9OSCi6TL+U5J6cxi7LAtmb
lZm0VTU7LJHiWqBi07lDqhLhRVNKWvyGAfZOFEDXF7o5cG8jIHv8SQuVp+klNVQmO+TmdR2T4ywn
5jJG9S8vgFyhNBoAM3/PABPuT/VG7MgWHBy1dvlXxdfsAcVhVPOflvMnyyNkt/gNikvzUb8abTyD
/ZIiAkam62ru5KQFZpWi9DBzVXc2324+TbMk6vhoNQzk3R1uLuyqQcmwIT1texJqAVC9qtQLeWUU
yA9fkMR3YNfnZiZBs3A50Rboa/uLx13TnZiolg8NsYPVD3d99fPdKFQfE6+/OvKTlgOp3BT2LyUk
Tk86Xfp91c25zaHj0uwEiEESA6uELa8kj0BxToX8Y09rU9WoYp2pInd2kUQpQGZfpndItJG7kk2c
h93U07UC6kYosE01eohyg3tHduSXqe3oQ7xyLQ8gS+vB+oHgU9mOatHmHLmp6i5nrJ5priHjhBQN
IFVD7lI0VYTl57N8heYKVBHGptTjiMfM+H3VGGwbW5YcoH4O1VUtm467NPV8UpTzwJiUk0EO1F2W
7B4cogelL6443muQiSTbkIg/i6keNDhLcE9RvdMNy87OaocFvKsYrnBYw+PZYHuDeGVO50aUILRG
Y+KFrVTiiiyTUYfxDWIJFjzNQFaCr01Q1JRQeOAw5V4Owdx0s4lA+nX9P/T1UbBp9FOK21/9ho+p
jUbxXhwKHiU8h18mf1+rCL3O0z4E3g8YmrHaCGxf58b+IP/911TBmRMuM9Z5bGhycbQkHsftxeql
3Hyt+/YSCcto75p3HgrOPrFy41GK1aU+d7fRlW8Ybep2ADjR8o4gG/o16qNtoNV8WF4AAwNNrAdt
Ymfou4KezxtEP3rUh4VgKwUjOhTdJKBERlrWpyObbXjYXheJKFYS67Fx/AoX/8JSJS+RVgyhh9+l
NYGjx+G2MCBz8iCD3wlElU/CLQaqma3eucz8Wo+499AvuEwTVWTwNS+j4isuVp2NFpOaBTxtYdJB
VDRltpznVxQwjUc89gMbyj63ptX3OfIPnhRnM21TzHcr+mHpHtkTUDp6Xdsqv5I5CIi0l2aYdVgI
uJ9slYJW7aaZ/Kl0nZRaenbUTYY5f3CK0qPujYsq0Zg8E8Mb28jDkjPmMisbTuuXY7DPOZZNit2u
QrL8O2G1O6qbyNCMODME+mBD1keZe50I5UgjQ9ve1yoabct+vELCgaeQ40LphiTcQg9eRuRgd/kw
YUzvFQLDzftwbqiX+nxp/pojXRhLXPDRIoqVrKBHGjtYiH77IE+ETMlLXpaL/3EOpg6SW1eWohNV
C8jBKMMtCgpCFN5aKHAR/ogzS6m/zYQh4kFJaQYJJgqiTiNdiDrN65/F4VJRpRomr/HBzWj3futA
8WTpnAZ/SbLsX5o/kb6zMuFwLyCpMZvyFAtptkezKKpS8BJCMSevptDPAfLlaQV02dcchO//Rd5W
c+N51duDicUhOp9jlMn5NukySelymSoZnVAnVhNyWa7QmgRpW0TvoSxAhIw9wnRVC01j+DFI4r5e
CJpHKh0Fk+RddjjsiFzOWcWILsy7TSAScFoy0WMDjnMYXwnrYL4a7NxZ7s0Zld5Y+O3PCprNapaU
BfzfJKALUMvWYTJG7EtSP0vqkVd4w2H6mg8aS9Ckcl2nLtCSsfP1u4CXHHJY74Zde77IWJsimY7+
TwyIH/dAYv3tuZE7ZS5ndxMjrN8uKVZfnGrWklUqlNGm0AJGnkUXsvtxQ3eGgQZsCkr6J4QQvshj
08Bl/4B5Vboc3RTJJeVpKDHXNkrHLKZxgMQEb/j/fXV41MCRdEHtn9YlXU3gwrZ5tDebq9lDXc00
GDCfAm/gRab5WlWv6hU3RnovW28Kwk1nTunHoPr03WFITN0ObJGnBcjcW7cG7JriTsvttkJrv/pH
rkoXWJdyIJfV6mw3wJH3jdKJam1A+xAdEhjU4BpBD+hMw7A5f0GdYWoPA7sc30Ukfn0wOV/2RgxX
rBmsfZNkHWyA6XSX4UzYSc/ZBI6WtJBJllXPNHgIiat8gwwFZBI1uGEkvY3U0GG8n+0IkUApm1GE
/nVviDAxbaUU0fEV2fs3kjYAfOWuOOKIlsqCxskVJkGCsdLhMWsJJOAA/O2Gl3AzFYx6Ho1bPjxN
wyD26kDQG0L3Z05QV9TTGnGXPmpdTWWRVuD2D1QSzP2CMj6PzYhALQNm6QkZ8tRsK3SfcGSqiJOX
lvFXequLzzy0DC5xj+5obkykQ+2b0Go0TYcDiOgQwvNDQpH1ZCitAjaplx0FIgZhBHffPvEeLo7q
z1NySMyeWggUkpCQuvcD5MDXFJNEdU8WfGnA/VCE4dAMIGMoEGmOcMr6kV4UAV6tfGIhvdpoVoT5
0XJKsd0zNmqpzxGi0hOtIBQKGd9lks9Tlzmdb28xsTNpHKNi6m4YBTk5mDLaf55jBOO4CqwvxnY1
2QnYAGf+MzzXaaGE5WAT8fnozlih4IDjr7/FVOh1zReVy3L6ytPIFXOX2Bc57Yj92sWwkPGEfI1m
KP5tpHdNJfi2PWnU+RGvlP1CvdRXXEmL7SGvFvmrHnVf6o2bFP7ZHiAP/RcyaJn6Q7V72VxPxZut
kP8J4N7+kMlOCOGe++f1RiSuIS9b8cAXbKrruBU0gny44hDC+YLW2Ar1aQNfL8JnoS4VTOD0lbyS
lEDjT/6/1yLYfmuenVTVPjDvuFhFZNoBwL9j6JfkDXkbiMbetASDVbbrkZk88+lk00B1EXj3yYor
bo+0RpYoFfSQxSMtVML7BepAA/F5o8xmt4TTrVh/jSKpVFfM3xOlqesZrbiixz6da+aVl0Vgk7hB
2+kpKImHL6hfOFZtkDARlucfsRsIwQrTtpndvByY1I9Fj3OsZR1Q1dNw5MKOPm6MCkKZm3JY6AjU
E7x21doEUloj9uobJNFGj4Ah5CZUXcYhdSvrf7UXLvwydvS5FwiwLbipDlWNH2a4902HsigCBS62
pFIRYr0mU2s5sNk+rEXEZu8/vRWQrQmVkMJRDZQFewYu1vsRZrqQtZ4wgqA2rUCFpO5Ute42Ub5I
XFpe5+NV+5T8RSZ38ZSKgM2ysLzf3hphRSBTuN+nqMwAqoKC1JhK1o/+oWCy2x+dfE6nMU4k0FGw
IqYj/ED0wAziV6WpPvojR+VPXSvCXBGfPEH7+/u3erRSRc6gLsrPc3XmpohOscm6/EPVoagybfJd
NUbHKKce9kMlVGB6o2mdcFTnettgrbW1oYn7GamKe+NQbRvbTPVnGPpSuDYLkSagEE268LAp2pSp
HtOO8FCeSuMGPTQFvBXtwZwTZtmp5/2NQ3dB6iIaT6kKRiwbnVRdi9dcIkWaBJLcrTLqWcflC7uD
TNAw8kdrXCFqm1UUACmmgxrrMDYglN7355VWqbp5uwHaOpasz1oan/hXqvSmBL+H9r/3L9k4aZ1g
2PxN/0EymIOuKJgal5wySwu8yB3xydXZLiYrpAbZ/D5N3GCLPDSvSae6+4bhG++42d4frF8AIY39
wvUNvWnPtRKdxZP/hbphoB6i3EGQs43EHUXDhQpqDVEYVH79cX2c1n028NoFtkJZl6E88Lehp0d5
PzUFTJwtzt6b1sJ1D0v/tWD8a86re6ZRfrtxMWCSfuz+VvL0AdLf/joeyV3TiQSGDRIZq8Zca6oX
3r6fk7qrQO0ngLCAfYwCfW418/kL6yO2x+m60euY2Jtu3DjUPl7/AEaMAyh1Xa7LawcDGQin2FMX
DPoCVctKqn4kP2umwfRosY7SEVG8UU812koHfYutJlLOAngYVj0P/w9xFQQkZNROzv0dQuJFTYfE
yRH/TAEbJOmlxjNGkvE7ahUZl6H2Fn2RtmjvNg/h1jVmoBO1QMuj5WTmlyyWZQPcIT4lMAIWraG6
c2X7vTP38GjXu8+mHGiomzBO3OEajQAQjhyycnDqwRlOEtdKE2pe6oXx7DBJL8CzT+hJuB4JUByv
9qaZxLso8fNw2itIgFndH/uI36m16383QfPQoaNAFZUKTbdOMRxfQKuD9a3BCM+KeIExUddV38L6
A2oFWmUg9JjDDrBBcY/nFOUIvNBPSyfzwGjyCz0Mt9Uo6JQtUUoY03ZTVJy7xmCCCFUZH2lwW2aQ
L4TCzO8eBCWkPnEG4oK73bG/mbFPsyHk0K9D3FxsRUslEZ0KRI3MnaNrYuZEZDTSvBjsncpk/9vt
S1UA061cn/6TCLirgkyLjDDprUewwK5eohCWIrHb/uGUumvqJN6M/0500nRQ4ul13VMT4/cTeFBv
F9FCMeTv2dTOrhZymXvlz/gaZs0VIkLk1nnqK8w2CSj0KhSypY4axEriFnZ9fC0icHOYn2oG+UIh
TGeC+XTK9QaSLbRz/8HxV4YmNc5aDF3Tq6VuImSclBQz04zW5FvP8uvYsmzcpuDm7otWqq8G5SZA
FbO0aNO15z75neOmYls1vPXO5SOBqmSoMwLYgwjVBKQt9maGuIwESGDnHswvIiyu9C/NMB/EXJRs
CXsDVu5u+Bg+p7CrweHtC5YlJWjaurRuAzbXICbbewlstQDeYwYAqQGLx+1d9412oTDUXhiLrBGg
bwn6ayeQPdSv/8QAdv7Hw4dRpdlkObzZaXh4qfbpmupm1oxHLTQ3JcvMPUjMyeqjTvSiYyEcx5UC
ICvDY65HR028S/yQYYzGtOn9CGCLGzhCNxB0t1pWVYzL/Q41XNBkQdVn3K+hbiMsNtqWHt+v5YZn
ZIW0X4J6YTnIOLIc3rKrjlQIRdAylSnJ0oflu165SUh3pgNbTe6cbaQN+gowEacfqQHllGouvoY5
mBs5/Qpx5fjltnufxLdFu8Sqfz7saA71pkEi7KUgw1Mfs4q0siM/gqyjsO6A/S3Md6BihvreAYrE
PSV0dcRB1owmhipRzuGKoX/wscWrotc11t7bwt+dKhCl1a6CH+eojsEw648gb5A2lVUTOXcZkpFO
o4WEMkrHrJSsGDRbZzb7nU2yB2o2qLscwm304l1XBBzPVnaxSsysWLn6rKZqEeSMl0/awBahvgPZ
CDqLXKoM5nmYm7WsXnjy1dTzP+1ZU3D44p8R16dWC6mLM6GNhY9OGRijdpDmfApOR+9bmZHJDkXP
lTCquisNETQ7NKL69khzSFuo1WOmyfgYYtrqGv3sfnbJ9R0tWFcAGnJfJgtleIrZAHw2tHGw0/hy
wiYg5ej5BOSTO4e0S1RVF7XyBNFFoiXh2k+Dh6Wvh/YAWkfNe4ZA91JwLGSvA5ziMMkFCYPTSdnw
9NcSc4wcX6/PobBHlQIs4O3rcr8bV2dNaCErMe4fiJgVKiHZ1ti5B33z0IUJton8nb9NuNt4y3f8
grdy3SprsOpm1zNOThbfwdJylxjMFoAPiCy6EDIzUFTLnd7jC5Yrc3di/4EzFxRZ8EBXWuQ/Ttjz
uxMXYZffNfWUqjl064dEd1CGHitBJg+PwUYm2QhBV/TQEQV13Cp1j4Iefc+BWR4g+wpsVWazcxti
R+931Opu6bH6KGwVKk+vgTfNobvw2xNxmCmuGOFOeoUMV0mKeCQPnrRYhe6OjfOF6AEOyR1NpTY+
Duf4bisv8rRHW1qQYaRQOZ9qad16GnCAT6AuiloROpwdFyDlHr1HvctsWKd2+aebPud2ALk66M2F
rlCKsRJdzIvNUUwIRx6C7Y+fJ2yVSBF8U7+iw+IG1wyTf1C5ZmPRlUSV2O+/7LrekTlHvv7f3Zit
3mhPGTh8SSLgYcDQUNXBGU55Dcg0MZEmikxzB6XmtQKaFpHrIAB3kl6vZ6d9ho6NaZMfyP4ZSHHZ
bhmrCBIxNrtbE+TR0Or33K76lDHqZAbGXX90U0yTD2XLlmSYGfRleoqAqMzYMOIohuS4XfEa4mu0
/1NHm7Ggo+ylXyKRDP7dRol06biE0o+6Uu2fUNIW5rzoulfsX/OqW08JF3xVYfTsaDv5lSU7h7be
VQ0TPoN5UOpbg7OPfH7/U7vPzVyWlatKZgGCwIt68JOgD+6EDVzL4X4nzvO1iQpuEnHb+VfZP9FJ
YAw6LSOkPxbxkkWbSkO/tlo7cYV6tYNvBxnUdqucVLUPjt/YTstx5CcYSfQfWHA7JdrhfCrTVD0c
vWMybrErgsqhkTmtm52rcBUcKMTwjMwPqQ+RBhRQx1sAs3JcymyiRlj/Ck28mYTE5m5mvwaS9vfK
u+y7FYtvFua4jRJrMX+qdD7jIQIsHRWhupp2W8CI8Z4k73guCzWBlQAUfiE6ihRR7dRHco3XP6jR
W6cjfr6koRNYBIlXgxA2nqB5pgJFB4o5N2lz0wEzJLyRKacKOAiaXf4hG7ibVeAUbh3dwmGFrx4T
ELMTv8mB2bM4K2E2zEU/fZ8Yzqug8fpqW9FDtdBLlmY2DdYFR6A2HUfK2QCzGLPt0A6taSCpvKAg
JphcdIIciJb4dItjhOGwJtSdM7FO0etlBalsvqAsmOf0KMAsOEhHWwLvG2ugAemaDYHvg0eCLRZs
Jco3qBaqmvN0+6WFFO1KG+hvOXoUlorSDdkxLVxstzQsEYvggMkJUpURZaLvOKAeehLnLZ+60CjM
mS19VCVgvUYmuYiJ9NKLACy3cc2L0Nc+jDcSr2v1pjbEdP9wI11nDXf64bvzTTk1i4e36usD6yYW
zIdKPAUeIpXStgcUMoNYwPodDCjMPa+U9tGZp1fhYnYk5k4rJxaktgYXj/0vJdrGLbzS6ozI85Oa
mSTp6jzjBW2WXEdWswVNKktyPJ+vcnR8cXgfBkXvgMsHKGTu+wW1D8CK7WYwDz5l0dTm/vXfEHCb
bzwj4dAruruvaMKEjYxvSi3lfdO89NM+rIjSTOvfFFFIHs/A2sjdCYeHJmS/miZYM+FIAs5wg+9z
rcSuAz15vWTQdu+F3G7dPNpsTeCDF+V3Jqgd6nkF6+604Er2n1PXLtlBwCbMFYXnCKTzr56Qz8QA
0vI8hW81hyBV0cSl3o1cpVo3cyc7wu/zqcpZCU2ITOShHso0LvTZdscCHDgOzWBY+3xYREo2SpJB
12e//A9zO+cAjMLqxvL36WBG9gUXzwQ1B+cL5TjWeBhjeGLHXarpoXzVhQdGLGzqWm4htK7tQhAq
RTqD6Wv61iw8d+vLbnDOCtAUrFSUgaQmtXx+rIVPm1F8bbMr6Oi1s5X9PzuNXAL+aQEND/SV5pyF
Wutne43EKEKj3GbcQtvzf09KXcFUwr1geTVLbqdUKVT2yu889ajlEdZgoQF4ejILlwxp1UMWVrMN
crUDHUDnBezeglygiIvatm1UF9i5GRsW9AyRySeAOgS2cVKjMLPQD8YEx2GAVKH4/eQCwygvk/Ji
QxQETHYzRxDqenn25svq7UfCYhJHJ43JvfmGNgM3opCbhxOahy9n31F3oGXa4PwF+zIyF3GQ10h/
/+VaFbMVNF2mAyIMEVjEe68HFoKLG8Q/NqQAuPY9kS7dOgHBbbVo0igGEQgNeuQN9+Nf03gGFZmw
UHt654w7XZrbc6WAeJT1PzPMr/Hikkz4KgEQR84HV1Pdxw4Ab1BjXF46AguussTiGIS+S0g4AFqx
EJDG3q+6Onjg5yhNnvd2ATpz16Yq17w2/Xj5p9agmP1QVBEAqyYgjcS8Th6V7/folwBRcX8zR1EI
aip/UTt06iR37LBOa9004ij87UzwZQK0ebUsh1v+XSuPHG9qqGQoASZwXFHphB8gHRPMrZqKpoUU
SG8ZRl0ROAK7WKPe8Eb5VeQJrKVZ9riyBDGI5XnAUCtHoISqpWe9LrTcIJCrIVv3nOx/qUJ/ePXD
kPht1xJ+Akk9V0MCMsTG83gxSlfnp3qZ26X09yzuiUTdAraS6ZrZZNTjwbf4/9LUeVDDngKlJe4U
AvcOEPSyQRNRwpHLvCyib3NA7qTQeethQEpof0DPhquNAZFD4nw54QzxoqkEeHkfvx2q3NBfSrHv
HpQYjHgHE4c+4uP9Rzb09V/VknyjHeEccggkw7wDbZ15ZJ8zqWVXwEffYyFKRCHc+9fCswQ9uPdn
Os2f6xsDvR637AWez2nkMHjampb/C4o8OoxcVxHubUwCrl0DPAoMu2sBCVuT9cXfw3q0Tx1MOJRc
NNC/wFZeygzbttimkOTPXXjXp4nyam+mrj4XQ7r49sgkiN2UDKN0ivAPlAa+6d/rd9pueue8FGL0
vfqi9CzU+1v3GF8Yl5Sm4GhWRhLOyYdNeq5gWH1HS/ExUbVpMmpFvK2QWumYE3OFf5bcDSvpOEMq
6EL4vb+WL3aJcd21vK8EyZa1p+Dm0uoXlHK6lH4b3a5b9pWc6UM5MNX9+V5JqJnozm3SytMJDx9y
WzI0kdyf7jG5EAJ5BYHfrOKl/zK1Ih09zpJgdOL/vE0D3aH6Mp27ZX/gNUvhyoSQv8EZd4z3QmCM
1HA1wst1lSIgL5ep1C+9CgxaR4xXp0VX8J+Lxi4VvOwPqf1tC+j8dUNiKgAxefAOxjhW5xPdTAEX
RVqVzP88o8A7wa9N2yz9ZGjIpNp63PCRPW/FsxWUwtIYXyK1bQu/7IdW6G7Db6aKLRcqje7Kyb+1
XdbMLXmZcq/ef/hdHJcGeyWTcj7GBhOrNqRM1AWyA5S3ASUj53KCMQgUsN+6591d3KmZTyUrWoOQ
fphSVgT+xiwWdBEuBHg6xqxNggnqem/O8u4errR55117GuGti+/LL+H81WoORiq7KYghoWx+5b4T
uYweMKuWEWajsH8JUiwrqz5EY2GGKIWF3daawZMOAyu0CetBbuMxOBvExX5Eb6a8fcpl7PwIwqUp
AdlSxMZh/npDrBmmdWQwV5fLsV2wHWWFQGjeZpe6YexgiMYiTpE4wjKzVFsZKyrl9DheFkOgTfDR
IloFYwrtfZI5f1eMXjoqe5xP525oHXbf2VKXkJp7W9ShmqQd08AKc7X9CHkGAs4Q+Eb9Pd7nwJfJ
DubIn2H0CDfc0Bq+GdJy6QIqAvQTslGnDMZ1adfgCCXxyjiozDVRV+Y+WygpAT6/TY/dPomBd6lB
MxX69/DWc93zs4hhIHsTnGCKY5RQOMdTtyy3ZrbiV4E7Lx7dEZ9RvORqaysH/tXV83N2YXr8FV7d
ZH/GbtOM+HFQF99D/Tvc+P6ds1leQEWFj9TbipU9mIiGJkmgvCNRMdFGnaCZYJRskJLamoEJh8WQ
UpkB4m+AKPYnL4B1zlnGYLDPmk1ayIU6c5OUJB+y6X7TX7N0N/Edet42nPX+XeXqxiQJfo4O+cTR
JcOKIoTPRbmmug/vtCCeZLjJwu1LfXs9F7I9GC0vbbhZLvE+sQ8em+Ihsr9XBl2KgY0C+ptjIa9/
ncAPn+JgLtb3GlxjLoeAPR0nIivd7mZr3RZGD2UjBJXjOegM17DwSnJmXGvWX2IBptDAcYZx68T1
cFhE4e9yQy2IYTyUUt15c6J96m5OqvLn0jUgQT3J8NmExpOBxiAHeSrAI3kwGybYWnBt0OJqA7j0
g5NOJw7io0mdLy6SCqlhX8MQiguYo2cw9WRKdO/V9eQ6kaZmw3Yub99TcKjJ2LcvlIEkxvCFe1JZ
IVVc3WkJOl170bScSmUJMtT1737nCoea0YiHbvh+Qv1ojE+xPFwoZZOZg5XoRrYPfDswIASkDodW
ni4ykghl/eyMttBiZBURsOmkept2zI0T7clB3osmbRWW4Ygyp1wEFWuSEsxuwWcDz7u5p8oIn2M2
x3Tmqn3oUP3l26s4Ev5XTWPqVBh8oZr5w7GvTy6W/AVtYsQMowbqO+rwdTXxMIUHAybOurmauoZt
UnkE8JG+lO3iGxRPcqplBnpHG/NcoH8fCz6dJk3zh87hV427skFYsAHrnFqKM0qTjSUgL6KiZCKV
6663Gsq6tJ9tYZMIn7hLmVdC72kyexhIe2f54tHhXZ8hTzlF9UKm2JBCta491hc+JpmUuuNL/6FK
3yncpBuJeiyA3JaG5vRIMLTpsrSccOMxiuQsdfHmL1mVFBbI1zz3uWgsI/0OeraDx+sI+pk09KlO
U8xxMYLiLYioGA1kja7uV0aHbqT2xBTWQrf4TCIhe6wAtN8yZGtpd/Dd98+H8J6UvQ/vAS1nDJPb
fJUZ1qq6RUCPD9uPlQ4PvwZTWWGb+7QHw7moa7bGBbHjIbC0pgLkGS0JEkbk7Cr7VzRpsnqYuTEt
vn0ggVu+7iXS3rgohVFu/yU8MglT9cZYm2pG1aSu0swy2CXrXcHmA/AuWnlblIJ9rhAigU72E0sl
taIQyyJEw9YiuRIQJ5kT3agup40QqJE2VMPepICIfq7KbsmNdz1oDzVT6y1klikPTzEGQsRQr3aY
FH/mzfkWEuPY7Qh4jmS8Lxl9pfelVrHMZkzbLJcTkEwyxKlPQP9Yw8JL+syRfadp/6Q72EKDyJTk
3sEmZaWpFuceROLFoI9o8yo7QS9stNmvuViMLvlAh7Il5zDP9WYhTn+gKbI2Yx0AfMO8F4nGvwzg
RUIzgBgEvQdS/67S/VIiPJK1PfILhl/U3usZYJvsBA2QBfH5BdMA553+Cfbe6C/rgUeDNRGb7X0v
6WKZw05V+8PUPcf45Qjksq/FozK+HXuJj6+lMvYKcMEz4BARoY+D7UcI7UUvNMOYYExp4sanguLA
oSN8xYig+gdHqEZ0ZZ/JzIhZgvaxssIDAW8KuCZN+SdbjrUG/VLOcd0jqAQyNpiS82tvmMCeNQdR
2NsWSPfg0jrPB/JnzRvR9j7LiRP2aaezYmSyIELNK8ueqkqwOKjP3XJZo97/axCcOBh26qYfyflX
kpGvMsWlFuXgwj5UyesmA19HW3Ss5cMK+4GoMo2AhYhsq+XJIUhPILeyve8P9cZqX6bES9ggw+IR
EKH+RSRit1hdofcya9UZdMw1PmO6rh+dcVBMGV9qUDRR8a70udZEw57sNPh6K/BaYO9lmNqbLbUS
3LKyNSMLGm8vF/5jKmWizkVWA/lJo51iU4VZ8Jq1guYLnOaAyDz8TNfj9EGbs98wjiysUtEa44T8
984IXA/9FlgHimUY2XyyqU2drt69he9Ko1R7DwhzhBE/Fq9XIlw3ufNlbJRQjXgevHbPOCN/WB1k
DNnlwPq/AJrez70xM5kQryLabx5ezJxu0aKUzR8EcmRMEmhAA771WSCRdfAxaz0xx66VYR/KrPrt
ym4b+PlDGOps4E9rrnLhg9TgJT2rpQrE9epMNH2r0HaZzRtisgEP1iJEfvxPVnodd/3azL4WUT4R
hxANbjf25e16jdcEaKm8TE4EXa6SmDH4xEY8ZBf4OSClJvKI4YxwZJHqhnoib3ddi1azDDO/r2O2
KBq+1livSroUY+kv7/yuzDgVNkWqHtff36QB3IXOCWuqi/sGKv82EsO5DT0I3sC1MveHQC7QCDIH
eWpWoZzxEBRJpi6GAwaosWeOz8e+G/DxiUvn/eBB1UcgqHnRLDCeur2fcmCdtdBaDzJ8hPoSbri/
rzn/0XWRJOxNV4BsHAso8o02/weqfRAPSziqUnoCgj/sHmESuIg1ERvAd6Y1wFGtbbnM0QD73UI0
UmnsNfdRhnNLu1iHWJd6kdq5LxHnqs1BPkrYmXT0qaCYxnqFs+fyhRRsDPYOsOvC8rrsitwLpiL5
KTfRbAtchO3Om24jKSSsY4yf1GnIHwDxyfFv8G5wwb9Eyd51w30zvUN6Er4oPFa1pZ3wc3McFWd5
LAlKiY4RwEKSFWBhBR/YkISL953i+lPsTBSRr7iNfDp6dg8zqclEA19rTJpvQcbDKGV6qQI89jxG
/YPjXFyQ9YnIOAAgkt056r6Xq8Hp+p++AAR5DcYMB0OpZDEOWF0yTQdv1F3WtbwCoZpvYMUrUoXc
c+sXdr4NJZdY4iDEfIHwgZbQ64lew/3WQUcoBC0Stc7shxC4jyBYm2+Mz40tNkPrRmf+P3hwkSYG
qJFBJ7/OW3BMfJo07lzOxWjA6tT41QhBY+w7MYqbyk8Bur60/wMdpXvoKS9Iy1nLuhG9kY+OGrzE
A1taChllxwFqn52IZbktOUy4rde87A4hFEcDBcuG5gEJ+p0q54JAvlSy2dZZwXpE7BIKfTcy1mGU
fpSJQc+OH4DmOcemPF2uRhxr8vIWEhsDWhDKWssS141bJ7zNdgSncW7JVBaN7JWPBX9VGcv0hKzr
Ip1o6dOd3FpTXBcH94DkpALIAOsBti5iE8V3frW9fh0DoIANpOgiAsU2EPuql2B7jBcse+SR6BXS
i/m1oPlmtveGg2QCAmupIInv77XN3PuU43F4J0ky+TJRIyhl/o2QSIoLpTMjzckI+A1Wy+VadCu2
/DxijnOxKIfxbgspFSJut4IW7+DRzcV0ntxzbCvVDW6bl333bADaFMja3J7KnHngZR3ParnL1CL0
sZVY5fo+u0tVBXr0dcbIIh3DdFV00bWyrfv4Jufx2tksmUl9h3mvMuseiZ65A2mfTAxwL3l5MYQi
G5X+WpSsKV85Gcrh1Jw4E8n58Mov54axiKHRIb19cOOnASsFoVmFl4DKTz38Sq9UUbhBSf9WdgrT
7u805A/Xy32FBFzgwNt+eA4NNOwxbMG68oGbFZClJQGUWS/gTYM3FPhlD4Il4KMg2kVYyijOwEuu
m1NC0F9B+w2pNLjwuO+Vw4VOCgIfK1/tv/BbUoU3LEL0GYclp5sXdKykpOMPLB+890vnjjZMZiyI
VGOw8S5UwX8dAyXgg5rhPqZfCLqjoct+5B6T1JSN+sU6OZakiYQuoTJC9PeKnEN40XWaBo5sGcF1
na6BgpUeeu9zb2OSIe0WVXd+ejslgM+X8jmNbYGC0IV0tFQi7Xr5gpDWcde2p09S75VOn/JnyxRo
nRmD1RNEqooAY0+lJro7ad1sAxBLH9aaPs5ibTNA80Q28thAqIE42zDu7G6PFjGHSGqWFImMih74
K7fKnoQ702J1F4cJHFrImTt+X1gO9ul9FULrzqOx1kTPbmIqzP6LufZXeXATH/SQ/IL8RSQyz0eY
HbyudHb39bNYLN7/+v/EVMZKWg6Feceh6UJ9URMYzc1u49x1WlFDhfm6nV/WOTJiKSeCeG6+D2SZ
nLasV5fYcevy26by2i1YtlEUQbhgFgi5emA+Jov/2Fkne6JG0MOYp8cedQi+jWI/sYU4Ln1PD5Qz
9q4zyQ/FXXtcBvTSL2Q//RCIAZBO50KD6M9noAZeC7wOQxMWBR892IaYfpKq9oZMA06K3aHWrztu
q3nN1c5Qn2XkDIj5SwUzeN1arv3DuVklrMbi5Ifxxj7s04BLqe6s8Hb6dQFa9SOCmYkwNOP05RBU
4b0EFVUHqffy+7OrwvGFPqDXuZ9lqzdbMxKUWcUwD31t/Kvou/JTWN5ki2VnUZ7LqizlAzIAuMGt
3bZ6mDxR1rBCWKw7hm6x09BrsfMZE5hJaslxuPy+uhrt1yA56Ed16JzhJnGHhJq9EWKl8u/5oUNG
MaszMT6ci1DzYyXFGuPdJiHa3xxtxFLHWwFLqcnTn3YaoSfuzb3rMZ7e57FhyOGsPqF1ObIDPqvO
Fow4yWbXFS3C1DKNssTkR/dOxGprbdZ8QTgfxbcTNf2/JNnva/pY+X/RLwPea0g3bubqeJYELIix
TuWxuJSdZUqb2+T8d2Q20FeB1uJU7hE1+Vwi37b6yQITSDwXmWuLPPwTwJOB/i7sq/lKvhYlXEZ8
1msN/UHVRid5rASG1cmTYBQCd9f40vpathLM1rQnhwnXD50DdOG/346dsbsbpXg2tUUwOXt+19O/
LducYh9gSFAeOrz5r5rH1ksN/3p+sdtoMkgNP78UVZxGCr/FC9iyxfPXuElg7zODpFQdo6OPzExW
uoc8BrSK1mOqhYp4yI6W/IrKgnUd2PtyZTibUMI1Wd5+MK/m+kq2GIHSePq31LOgYCIf0Fc3Kx3K
Wm8k3R4MY+DwTVX2CnLhIWklJRwMSy165JorhQEuNTLOyR/oGlNQ82EX2uornZU+LosYf54RIPWk
Ot3/RybxR3qIKvcZ8sVYxbFu9YdmXNZh4j6C1WAeAeSNYKuehRwO+7EhiUYRNGPF+dTRfgVKrvFY
omn7F+mnwpFPNz3sudomrZPz8ZIYQ6yVlSA/dCz5MLSbcJvp6ybGUWwd6F871eaXLo8XAAQmOad/
4KvuWKMslRqTD5KzMrwTGXyjP/r8Fdm8DecDjc4yU8zREOHSTi7jSg581X7zsjyerWmAQtZxGbTB
E/kUEIy/xhVq1VqPgAwL5UJxGKTFCm8nT+0cxwggbflY5Vmv3gIjUCecWjKE8ZyxQtftbIYL6WIY
hbKtR01reqqCGQ21fb798rlw5uReEh+jwr0PbbenYYlozHQj8ZVmrhUuQQuVlboFE8mkptsmoK53
1vALMWazakG1T/SoXe5Bi4ZQ4ppVDFoVaORbgQBl824xa55Hjh3agIMj+O40GUUbjYA/wacsi2zc
UNC+paS+s5vTUPINvBWLmhsl/jthLP0YrCfG7wXVAB6tg+I4o5pxjtZ0jtRmjiZDpFSrcP13ixdw
Xh+NkRPb+cmFkjuVikt+76D6amX52/UO1/3GmeZB6HmDrTmg0NSnod/pTY8NVH6lM/gNi3nj8Zus
dT9PirusMpaZmaW5qr3AP3/gpsJeK/SydnW5F3+gL0rinPeysNpW1FhrD5VVkpWXS6AX1gx7awd/
kkDL3drESYiuydEine+7FLMYq49Bn2WaJu5t7SzVhASkRredx0b88y2Y8//Fbvo/yhUDTJrnJdXl
lRyKYuzpCqSYJnXk6a6U5ElSoTbAYuTVqdtcoQaNCMN7A9b0zNeHSfaLJbEhLtZhIlGRDmrXY5Si
xe1Sj8t95PsH5Et1VFLk/nhVaRvxzWkc473QOE5jDXEzhWSAudTLObFk8E2PIY9eS7QU1XJO6EmY
PgA0/W2+TUoVx3ojzSSPKI1hlINgFU3JvVA45MsuVnheV+so9CeJYfP5X1win+gbgesCc5myhq8M
CZcPZLYQdnpuvaAoL7sA5bfcY/AlFbuu1STCsq+LJ/N1ESF6xVYE4xD9MZwfDI8PVIFiw/G5EDav
XiwkeQLks1cH94tqyCtBiNgj2ddiGd77E6KGu2+C7VYQGIRs5rRiJjeEUCN5dwnxABTYv5QYA6s2
YPbAPjoMIhDmWFuqfUgYWLJsncwD0ejlvDX8Jgj4ivJzS6/11lFkCj9SzmRuSv+kxP1ng2C1YdE1
BekI4f7ShwTwkXDkKurWlnvH83tMJ1YmstLxYM2tl0I79Kwi2kiqc+z65H83TKQzEEUgKPvGcQ5t
hV3gMGWkHZxvefB9rp5zn6iCxb+2S+U00GBpfbPBRgGbsWGNWuapwBt6yL0kXoJdG5UkWj4gZfxV
Epy15nYK3tOxZpX+KxhCU7RleGL5lItlQ8H+ebPciKUL3Ig2Yq9tIWonkLpr+eQ96pR1npd/bfC3
KdtbD137deS1yRay3J22VLldc+CJy/Dc6Nq3bpbs1/nZDr93dWds8VEPZGHo/Y7K+4QgUSRhLE+k
99d2Mvsw++HIlsnK3nE8txJJAlIvVY60Xidvc2y5j7VwFtoB2LY3bjwSMsQAFYekOVD6NyIDz+J0
GAeosZW7sW0VzowngKLEP6FIMlyG31qIkF11/uHpaZvcibT6IoJYz0NesVKKsX6QhzAEXtRzOCpg
PLbuNv1QeCwF9a7b0TNRS1/ohpiPAkhTwiqLdv8BxrJV9hDAAypHYuIXpa02/WNZTZgq7aOEnFzS
9vCs2K0MpDDE8gGXvCskOwLKA9DnfY2MDxCeAUFLUUvtIP4dHdwpwNvrepwDVRE0wV5fuHlawHvM
n8Meuz9BxPa2azCeBK7k7rzninfC5Hcvfc8rrr1qAHXdiNK2y2HvQnTCeGvFu3GekvJ0FlbfBbmq
WKVC5+Q9cm1auLmlduDh/6bb74e42ub6VBfyEFrZPxO9ga+rNUkNgG+aicoR117ScLeDgnp23CqY
V9jR2QVWPzxrfOjjhXzRpPukopozHcyQeSINWu6VBIMiL3+fiPRT0BK6jcGvV88f30DypWlbZrjj
qR+ZD3AKL6FieKeeruBQU5xpfnhTBIXzUR0X96rnDdMkO5nnRzJ79xIqQ4po92ryCfIsn/TvYmf8
R6MYlxTx6lXm545NCYBq4odKbtO02SPoBsixlIjfLdS9n/ZMNYlQMQiaO4LynXU+B491MMMm2ehB
z69uoyLbIq38Vxzb3a3N3FR4F5v1URnSXJLhU5i/k6mVdijFsdUdzuvT9O+gPj9MjYM+wgcM8MzD
sa/QzbNd43XqXcdd0A16Pjwtnq/3+7zzj6sYCeZTVM4fb/0lrN9Eel+ZLC8qNsiczBgoFG8amaQY
i0FsiYrTQyuhuhNXLwBxOQL7eLoCfJmNleFLboBrLhzCpD7G4qJO8vQEIc84JgW1huSpA8RbKmy5
Tii1b/MyQIm4hQ5/rpdZFuING/mWY8QOacSDJnZVT62QLcyM80Gyoz5PA7qoaPi/KJrB9VJOzZYa
dVVtMAyhdQNd6NcnSP2P6fCrS/Cqv95ATAqfmOOPFMbE0Tzg4KfneF7KhGE/tfdA5e8srhg0Kmru
oKbKIM0cmbwcYXcJy8P9WRSx0jwYAVMlR09lEoUXTsJgqCZKIrXbIpzxWTSvxRBhh7367OhsHWQW
T+8UkyvNNuHC9gn9qW0WpEhIJH+Gf3d98FruJhnXQ2LuOMsys+6ycCjFzYAANhA1pAKt0lfZegDN
Nbm9fiVbp0xTuhVBrellH9zhzxwOGTThRdCg5GO/TKXs06zZ2V1gVG0ZVeLyql77CK0Uk2YxfoSk
jsvb8uSBbRljBiIksYJBncctuajAHpy7OglFXcz3n/cVcxoq3HsDWPaFAwuiZAgbIJ/N2daNnHOk
R+qlfUf1aTbgfYcLax0JBKOaTANfez2tVJmutEij/6m/P1baWhzU2GBqe4EG/MRPFsGbAkuy7KUY
FfNxcq3NaBhrU1ZHk40hkdVSqSSS9Vo5JokxBPFdsn7U1+N/N88//COzwEg5mt5Pgb47+hgT+1+a
/9qct1Gh2cUbCfuDUt4ubkyg3pf3too0Cub0rlaehoLZW9Bxp2CCQH/2TqxUCGaCO95NXNWXVTzf
omQMFz3FzZRhpYV5+UzASDFJcUBfHkFJWeo1laf5wd/t2ZfF+eS8nHR5MLYtwmLpTcwmVFAAPUhp
3gvmA7Uu9smcvUG4o/4Bz5y8l6Lw3t2PaetJVlvnGQn0oVnYqRTTPkM8FtsqTLhizC4buH5Dirqq
SKWAqJXRy0VU1XpEx/l/A008PRd6tXcweNJFpZwocChVkcmEJ2nr3hboG2Kd36w4rBLpgyJyNX9X
aVkZxtVl9L61WOKXCkK1HCilzaGT5UgMTNIV971FgENZlUWvTFMLDE8bSaZ/NmDLJ4d5LP02sNVo
Mb7wQuXYlCXUa0ALuqarI6q7e/0um5JD0jllq0Mkdl1PDT/a+Ule+rgi5aFkwkuTDKLesQfmUi6r
0OzGNYIIM8tFzg5zwD/elJyJG1fgpaezwf5t/Z0795k4ggzs3ArnTWSLB4LQ7RTn+jpZNnWfQRcy
UmMyf5BNdu96JQ+iKt8wICDwLVTfvG3PEcB6FQeab3B3QFg5zen/JFedQIqkOqQOx3mMElm31+29
qS74x/AOk4ERce2llJcP5+U3+NXz7ape0qUvAq7ZZ7Wtt6Lx4wmfKbGW8m/QB+lWtMiSBIGEwgdm
7x6gy91tEuFBSgTyByKqURxUdc/CmHKTfsiSrSyONiARnaMFsjUsR63oLx+BJqC/ERWfkUGJEX0K
UVLMuJdtE0LqAgBLna0YHR+3Pht6uEejwfewvbFfYo+rrm1ZSxVAtMj/SSAY++/R9eD4MxDZ7NYb
rBi1yigr+mrgp1Okd29qkgPxxJnvLIEcIAeSKjAFVZphtImF2thwO2dC1VmLoVni1STiOXZ56XK7
yfkx895wgF7s4GYOWrNUg2LNHP0HPTRJJJkJy3jpQSqKHxRlbE+Q0mSAjCCbas7N/FL1lMkM57BO
hz0c7UV/Ic7gWhWQ5dP6AmB2YRkiUREjiOz+oB0dOECgJy/6ypUd4HAcg5x4I0TiYCDMxg/swrJu
XDnL3tw64TUFz9lhM9hqFchgcF6ydvfZf0xetYNHYAEH5q5qKXIbV9ENCcbm0eAZqJ8xwOIC8W7y
thf2Da3U3pF5LL47cY/SG8anx1sUtn0DPZyVpsEVLd6pwD5Zp6G0aZCgMWKbwUFh1uCpdP+4TmT2
oh9DiWwDh89XqVWW/VfbMapP7b147WqLovbddr8hH+uRJg8VwDCSDFknD12DUbD1LDQeSsNGgTBG
VNupw44QfDCi0NgxWOFrPAEvkUoWIFW7QFNfm93S49KB7tglqhj8uR6DZ8ZrSXm6lPMX0JmKggrT
qVZKH080fL7+lAO/s0+JynSgKZjKnpiVNsitk/Xwkn8LBOlD+mXt+5uAqmYbo8sisFGY4rm0A42l
CcRnXWAj3Ev6Q5zX/NU1ApEp63fJ7o5tY3ARnEWe3v9IFWqc6pwQVfNLfSA+/LG/VWv4/Cx1U3X4
azc7kMUMvjGPmRJpAXcaQ108/aC1Dgcz2EFfIKANl4+rroK3I8mHRZVdm6GRU5d14+u2jWfSCCRh
BLf5UwGuxAoUtOvD0Ce/UyUfi35gnnyM8BUNXtZkbA2uxmHeizhqcmsu4sGyQ9/ujB7LB8nQQENl
5jLJDZSQMQIuIKUTj1IYq0tQV9euVJEoYJ9sIXt6+RhXApkq8dq8pKee/vosj7sq3JNTqNeYp5Rl
20XnqpE9BOVlYhCRKtBJ/57uVZwxPdTTXALcZNf6DJEtVWleUmkPrf05rbjLD5+aizBGLSZA+Cfo
lhpkaJow9LEwTWJk2wCGHeyCuAjBKlsmr8LvtW6sVWPG1aqkIlbrAyy8vXzPfaLs5K0aKVOfsNcL
gKNTuQdePpHeEQCP3DRLuM48tCTnM6UOiMytWADvpsRRMXkvPwIfgkGpryHa7ortr9sdleM+7OyQ
yBsyjUL2K9BRXeUtBeUcND9Z+ZRMz4mpPphR1bdvF2zdGjyunpK1MzVHza7tMRXAk/eNX+ewxZcx
1sP0qEeIE9OexlvM06+8BYBmQKXg6Db46rEaQFUUVrSitf3gl3XBiCO0KGqymGDYtqayvunVIOQh
tHxzsh8v8MBJd6Or/PWVPIdlJq1lIlPJ/0Ku8Wn9TtNm/iBeQDTOpOIwQTG7YTyKUYL0s4SJZz5a
jPoaWZQVPMI/XxtKeKyMoEZMPrUpczWQBlypY2auP1rOoTFVuzVGZZF1xmCNpdMb4fk/ev6tW3Rq
REivdVketbKT17khPciN13GD6HIszNyDNJzNSKw6+aVW1F/o2PUWJ9o1U6AewFbMFbZo0fWODqHy
wtVxfrcwm+T5qYJxY2zollPK7fpA3nTHxjJ5ah6s+jwVaPyek3OQ/LXRX5WfemZDQcI525AtT15x
zCqWDeeGmUo44Yv2Nu0MXL2kbII7Pk8CfoSs95rvOjh/TIsnkCjmB+dhrvcUUEFRYZ/4szTEjsQE
LeMRe9yJ+PYr7xBCYdGyF3WIIVdr8RBB3T5uVFaf2botKzYemg3lqADV4ijYeq1GSFs9EiGZ0MRs
mjZeiD682SBlL4Buo718ETF58vHBhTOOL4uQz8sIU6TEHJ+oHihExSD+EwVn87WEdHcCxjQp921T
CHx/gVzSbbUNwejISpyXCva6Dbi+s2mCmf66rZlD+vsC7U06QwoNuUfGMaK3H/HBnVKjWsGeDqKY
2zjXhmkT4zIKelh/JCNgEAtt5FNKJoZOA7d+9WwI7iBc12JMKYZluTFPsR0FYMiLq8S21HghsYMw
ehx4ejLnA6/G/QnuJ7W0fn3m6XQaAlMucGrP/eN08XtCJYC8zm5y4ItN4gOuawFlyzKjeJFPyBhA
p9o0mXMq2ORFk9GHkgaKhml+F2onr+QPwiMAJBkCOau8eSaIxgbL9waizElPP7T9n1SV5L9hVJmq
F05RWMfreeHJtVX9wfl7I8Iw3mmsMjzM2FhkENtgnR4VJZM0C58EbNdlPBhWXvxqXnqQ2Du3+Fih
4tvbkNve7pXI95Feq3xUZ4ovv/oyaw7+GcTJnDlnaO0OrVN9KO/7zvCvGi/83IWIyKH+NCOZkgLI
W3Q5NdvWTamQR5kJyD2XAFoWzv8lLZC6tDVnrd42RypvXwUJYaNi6nNzzxB2t4ZkWDlhMqcykP90
0BtZ5eyM22nj8eImXZHwxbsr+3G0+6Efl0aGHcKM/dlZgPbXyO1ahGD8KAAdc+5OMbFLlFRzGwIJ
iOSomy51PekIVlppeA2QHg7cNdObUgXIOC0HmEooGSmfHqWmB0nhahrUaduPxnik5MDnKudZeCLh
v9XVSan1TANuukGySsB8R4av+Z9Q8vfyhfntUrkT/s/q+0DRQiUf5Zgu5TJSI/j00ScQ66z8a8hY
5Kubs9YsxkW6PQ4uGsYEIM7bxidBc1xMRuXE1UYZi2N7bvV527K7i9Ow/LWNlRpDDE8Mewv34PeO
ZKlqVZ3nkEeAP5n5Z/5DMswLfB94IQuw4Esb5GANlEVDsiG6VKZw/c5drD36lRxPRi8FqWl39kTp
pB8eQDgFsg0GFeVV73uSc7IXe1D0GNjD+PyEPyvLEGKi4ltBNPLu7HbdzI4Yv784oZhDaPh+oO/R
LQEYilXrwa1Sv8mZU57jK3v3NxHYKcKyKEOaWEpsztCW+Bi8OOyqBn7YLXq4IorfiUknd7RMW5WY
I1AIDg+86OVxW17tYP7g8pvDDYvGisO1n9DLp8V9OYyic3JGuMwovaMnMHbjMDqOvUOhycbG5Lpq
3a41yX808ktWK7ASfLGkdYcPtP9qLoZ0ifkLJpIo6DiLs/s4xevUmBVdGTahmyQQ3jQRjQu0HEx1
J6IPNEObmyC+CF8SYYzM5wxre+9z/MV/lYqUNl/hlLcLcSRCv0Dem4t+3ahpPoaVwvRzkws8ZqeW
3tSVmGNQ2FciNCjWrJDqpyntz8oG+jmKDFqPb4Mbw1r1L3qQcwbmDH74QAcGhuqNZ09bDB/cYjYS
2C/YMZ9JIDwyDDtjYlTMJyTXwcR52iXsn3uzoM28c+CI+gK3XBiSXReTfLhiEQoFUfXIIvvWjZ1J
0fvrbaGM1mFCE40RpZzD8Iy2CCAU+d1FnI1wUirJG/RofV8EnwiPWGWtvkTLNwDusBTg2Wm2Y6HT
+kD2nnBEC9nSJoi8jGBr8hijYZs/mFQHW+x8/Nho/Xyx08eitJTBd7RBYFDfSudi/xoGI2H9SI/P
g/zVbdIQpz3gtC5VLZBKxWPK9O4r6FwRj/VcLDQM9/upZHryiVX5VYlGfIBR1L4UgXctZp9pFawM
j6iMWREr4dYgro+Eu+vVlt8Beq9sXH5OiEcEIOlORnv7KhwYzSRaKGN3TY7VS9ADRlPKH7sGQeKl
abYWyUwziUD1/65fLTQP1guv7iVuESl4/fQEP9LIc/W0WI19XEkFf9/PEZXkZjy76mfQAdoB5XBx
BRhIq+VSWNTgeIp1xXjFHKBUz+BLzRiZrrOgk4lZDAO7i/ZzM7/PfJKx86WCY/DhcYQ8DuoT2Ibc
EdWZ3caHAlUg/kQIDkQWA5HhHkhx0Loe2lWQaTNXavP92iIYkqI0u0V+3iUDWrxVRwU607fPBBoY
OZ1NZUx88tX64GSTQBWDmxHDoUdkvJVW3kgksz5DlxKUEhlZBFQSMTtczA4dQoXhqZFnXar4Wf47
vrPPvsirRI2xjVdEv/NBEIcTZVNH6d9MDOh/LRrbVHAmV4r4yiX6vCrHURzc7KEnt4mkimcDe5Kk
Fc8yMm8TvLHRGnYnEbfMGJU0oGIcnOtRMcjbR221AbUxSB4/4pNsaOhYn1wChM7f3BLFGKiSy3qn
BgI49MkFd3anogV7kmGbXWAJBEQB5FjtK++g6frygLYOLPCMqXvel1Mp1xupT9LVMvx9tG1qliCl
9vhI2W5AKBUL2Zl+dxUaXnkndQhFke5A3fzfKArH1G2gWuSRj0yKbC3rQ/ZChXnX+T3GTl5uDseh
IsLXSILjzYeFdVllFqoQUmRO/2QPOOZ9GOVX7wJyZ9D3bb1dC83bcpJ+WAUSt33x3dVnWHCvFSZr
Q8chFlTaNlH/hlaZRU/PW6EaSSK6qTm0BL8xrXC8dFLzUTwlWK4nBjBFqmvsTybbhpSENMnL6uFy
GhTl2DlyVqPxExTNQ4oyfSRLpSPFE+GklwcIHvBdG9tkKyZ49bnTzw+zE7nFyEGYfM3NOi+v0IGN
qV2O6cAdr3ahignA6VJWUfIg/Xt18OpGHygv12nqIZ7uGs8Yo7Qay9MU59k029FGWLc0f9o1t64K
6hB30uhub9YolgED5XxA7jGw/53z5wTfLDAbsD8nnL7Kx0iAmpThc/5RUi/oxl1DJMlmV/E37nxm
bpl/FZKd7tJsIDp8tJk2QaW5RjitW9bEVz7Lb1F+e2W+9aiLTMYPh8HX14x985zaYURdlDexsV76
cSU4FQW1QTSnktJvaBq7al7kN63CvxPHIhnSnHnpq9DxWCAVnnHdDTPJA+LA5aGeuzhU26KoRLBc
9VYhEujbTrrAtq8uv2xKUSxbU9o4Knf1FX17W+pF+ZFHlfR3sb5syCkjzBQI8seuVCjK/GMr9htm
iv84V/skQt4Yxgc3cglEDoK+N5da+yc/SGEBCvnkehllqcQqmVRtr5uUnabhYpZavxZKHNgv1ND1
91MEf5ugE3nXVIV/9D5VC41KEe+i3jR5F3wnrBYR1b+oAuqnVJ9LcWeKXSxKLIuxa3bT8Kt6x95z
N9MUmkYCJB7zPhZfFlXqOir4VR5+stvwcMjMTzUHno53Lb1UM27lIpprs6U+iYc9NrRwcOQZmAte
CSHnz3Gp9AXkTVRGbhZTYX6ZrdAP4PY8RLgNCW5ePp+gXvtyntXEERewxhX/JAhpHlSFLz7tW1sS
vN8dHPQM13c4Y37pHI+rbEQD+JElflCt+wktx2sGqtrSFTN8tv9wvNt3i+opogZGGfONhBD2uaRa
2XC79TOcJuc20jdy8rOrIgAFgK4D1XdYobqIdQsVTQxWSr44FjCYShZ2l4l4uko1hl1k9z3vTMQT
gaMjrTaTnw3hU+u1iG0494+0VIpQFPgbDKEh6MkbynIWXTnUkKS5HzngP4Gof9F1EkQbBFgnqZIi
4plpzQbwD5HdTko9vjrgend0xk009F5kV+yx7Y8qz+i5FPYANS5NMyuHz/0mg/Jj7U2SlViNEbv4
NJXD/hi8QIBFsV8bx6tzcLDKo/vJCOcScHIqJhgDhR1CI3lJVL6Sp5Tm/6lAsu29G4wZjlJ5co+M
u8OvPXdWr8mRwrQugE0bQmm8i7RBKEnbyDJAyNNg4awtE/DUOpa6x5zpdrF0oDVsHgpsO07IYXpi
ARUMk0Y+aVBSXKJOqgoA7JyqOkC62AAHD+jt0TyALmjDqexuotn1hQGTSACFeWzA+mgi2FFLhRop
TjyBDjZ8Pqa9eeasiAejXDXwv5uMY5vtuPx12dfFnN4F0qDG8XfuNWRAuoUcAyY93ApBqTptjctY
Sq6/GHwKvYM7pmX9m5Gm9ZLGgd2ybg/AsGKhe0sK/5vj6zGF7GruUs9ZayV18BzZnNTdXthUZA1x
4Lo6D7A5Il0iefhCSeW+3Aj8dLr2irjeFefYFnn5RY7QPHwDSx23mq5+vf+w7+ABWVlsFm2fH+XD
1NQ8dtUe2XkFgsgWv9WDCCMQwXiOD16m2Y7aXnZQ1kGHV//KcjbCmF8nSoUaqKuyLG3NomLq5oQl
juhHRVluNGNG5YbYKsIqQVksEV3kumBr6mRHbc7X/QGzkAX5hNMoRW9WicMJkfaqfilI3kAO/ncg
/7BiYmYWrhmT+cuAMDZhiwZ5e+rjwU9mf3tpFOGQ6a8bqyeBvwmPR/faX/YxcLMV/fhYmLDjAOlw
n2Izbni8fNeGlUb6D/b2siGrUTN4YT3LT4jzj/5WQMb31lEIYDaXGpR0WxTqYaittSAvpszvNDXX
DU6Mq6CXLt2hP2xK9LqDHO8BUqAVfyMd63Ua1N2xB0qz79sx54TgoCsJ7SOdzUtOISfIMV3oSU3J
JN+CmK+lk5Ktk7/lFsVXh+yxkJJtVvL9LGTUortSbfgqSHuWaSiFtY0kZwZoKpAhBEUPwIjtrIhD
guj8dxLP3uXFC9IIFHPgrnb/J9IAsh5JrGt1e+H2cfUFZY73kTxTbJPTdZEmbAY+pQbbBGX3F7Cc
0DDBsFiyHGuj1KdPGbd4wzJkF7lqUCoY97wfJh2a5td2jUACMNyy0EXWqfeIWG2kOftB+o3Vf9JW
4JjSnMyDLCYXfCmmplFGpPfcFHFI10c9yMT2pRjp5FkF9LY+wZ6HyzxNToBBYgv9/jBeaTYbWveZ
SIEMKdQ7RqMHGqz1OWLW6isS/WUE7BUq4r91xNYIovJWJ5ZC0wyNwq0sNV89exheOUTeXJqu6VqS
EyBaNvcbx2dsL1s2I6XSgRjeAicytk8TzqN4XMTRBRLAxpsrNGw4RQ0S3a2dihuKfbb4WkOBlDUr
azaYXwp0xuuExx+hRAiTMAzy4h+6vCFHqUAzsqC/FQwCpaQolIb0LlQDScjBaZ6EePfgdrKGSKE8
aAxueuq+O+jpuAU6p2EDhNma0CY9XY9uT+s++AuRRH8YaXxj9AtQWIuBsBqbLD9vTOmuT1XenQmd
oKoQ96UsjI8q0lyAQr5wy9Cax0xhrn4xc1h/gKLX0cI/9nNgC3lIjD5v5JRuC1X3JDUbR5z6h4lA
ezeNVunVMCkMDRBoYAsMF7ZiIkxwQNMasOU0kJLU7CtIS92NiKMmf1bbyDeZAJDyI65RHNhzkICm
Ljy1U4ONzG08D0tlqN01xxVGWhhMAPmVCAs27UmWi6FS5i+TBURKqQZ+Z5Y0VXCtplszF4p8Kcmx
TgBkCuG1PFSNO68FY7HQ+xU95+FtZpT/obqi/RXjTYadX+KLyf1shQpYv3Ec8Zd+KvPigN0M51Oi
2ZKLCKz+o3SpATuyT2sovBSQ2DC2xAg8t+FLby145K2u8Vp+1r1BX2Xn3cINZkAGPvPUVct/HjRJ
rtUZoBnmn6UX+q7rUQmAc0rAwS0/Z9c5p4Ak2KDVOK+6kurE7gNuQswjq+E7mjgPnqIqr7v46Heb
2TGl9zYy6Zt8Bl1Du5FzEAkhZYsWAI+gYXt1mt5JzvgItHg+tQhxBJe6mB5m56F3121drDcndqby
V71QigKR7YLirqbmLhjFEVn7ku6yujlRW8Jb5DZSc6DAZBpg6JBj+dWRpw9zyydsHOMorREF3hIp
/JWRoKW50WI+jIUlZaqCIBOR+7dVg4kDTiJyW4mGBdta2+47wBZSi+LPVYfKq/RxX4MS2bg0E7rP
ep8T+Q9qYwhDNBlto9SO6fAAeKDitmxPnbE39430yb6c2uy9UPYkOVqflPvizjuTnpWEWeKchUeq
A118WGDwVN5dzVLxUJ3YvU6v8qkDc2BY/ujHyMbjJq4gT1eiBIUxU0hvdCuVGpO4iIDUDYLV64F4
7s7nkrELeTG9O5RYLZ4eXzaFWHtGv1olEbiHr6FfxIHRqVBhL35gQMPcfJwp0PEH1gdwv+smIHzs
i/wxADKcNdqbCR8TB3hZVR5nOcVhiRyJytsS0JG5hNeIWBIv76sS0o8LyGC7fgNXktYLGXZ845zu
Ep1zO7etAuTH0Ivs4DqXIMZ3CfyIxMRPZ9L4hYfu+1Oc2001kraH0FVGFMB7McYFJc20JDL1d8ah
Ef4J1FBl2NLHFYjnitaEebYdrmwgODQeHjM5l752ccmIJHOWFQkOS7Ko5xuMbUBcY8D3+RziMpUk
DZ5c7bZaEuohtjx3vlqKmu4TfMj//E5c1CXBugYQ35DaDoO/ipIiYoqMtX1A6LuoivHcxF6R39px
4Px+IBz0JxoB5Eyh7tWYDjcEIiyg+Zpfo7pr3nT90GMzuqLznDxfo3oSnttkshrQyPF9FZmvuX9n
BgJte55r9UM+Pb6EkqeSkht1b49cB5gmu7oZZqzXY13TV3e1PjwAOiCsInL83IIMuvHVAiHKUlrT
MIW1PPnLMGKSEye8y6ftno+Bu/zS3bY/+7J0kDFDLe98zuoU9YFarEw3QtVmsJj/+uVP5Rc6LqYL
xtgZ7sqdzmwIZoUa/cRscue4tY2sBxlgMtWf4/xLYn38Ged2fWjG2gyAa89oJ5SSPoZA+xsiZPHZ
PHBTl+kaR5nYTihTT3rPrxHjmWrI1Ej6hUz5p+ybd/Nc9DaSE68/1Vpy9BycaMo6lTLqdc01NLKv
oiSDoTBd/rxNERnrlqNEmauD5u2uyiDixtsblg4gdtAaMy1ba61i2a6IgvCakq9bnz6c9AUoN6ml
k49hySyL2NuGKsEI+zuRw5W7zKz+4A8kL64CMakAFcQQAxfzQ3jzwS1h2Lhr7WxOp8gL/ekQTSyO
QRQWdcGPyirvmXZH6FCmDoCelQNNjwfAIujZ8SUhyNq7xSqSPbuIIhyinnQl5JF0THmFXk027ONC
pzqAeytTscfo5Ak1YYgNYYMDmmqBslfV8xJGzK7HEPivSOiQDd2ygGkXM3QKabSwx6KNMZ79NBno
Ub21Yt/1bPqJJ5/qzEg2Gtd+r2UA9PazCLUH9WmyCPbvSX1gTWwDhChfMf1taM8OK8xAb4ZN4s6G
rGUlz2g9pSj12xdW8U0ZxRZVTO6YeulDiTlpI2A9ozsFkBM6x3jQtIVIMyvrB8aurYahp/iy/ayt
3AqPghdGFs62g08wDn8uWtgtcXwdAAyNyVKVGT8pmmVGH6KKBT+HKoPYCmV3RVfTVzoQNxa0HC1x
f0Xr7+WBGumxzF/KqPiiDPnoAGe+I3+BJHLXff8gxGA383UBTqwdAgMNbhhioRYABFfSekQtRpKe
75L8SW7Jhs/JpUN8Y+0mabMYfSm6B/k0++a9T8/ZjXSy0hBdOJhJwsOlYHPQ80tdfFoOLx7yDH/u
ybfJ8A4ajFo7YUsyKeMavi7cx744zt9hrKkh6VjQ8eN06se1rJLb4/gXNBuBj5J8xYM90fziuNOY
Bx3G1348KUEG1tjmfKpni7twZ2O6gIoPr/LIVB0RMyzmEYfONAO95CPrrxuk7vJZi/VOdiQfPxp+
68v4aLH8/Qe+ygcgVtqPjm1At8PeJeKO1RFZFdSfgFMl0z3/AMBZv9rnl2GhmD96DgP7HFKyMz11
PU7bnS1zCcMNOALshsPJiPZ904n172M/PfeIlOaNTw1aYZ01NvpDvZxrNnRr5H/B95wdfXExI9PK
xTNVjfAbnXoM4W0DXSN89PopadQdO9bMnQHROtkmRbhpA0BD6U9K4mpVaaSudnsuHPr4+mjpCoM0
jolyKA+SA2sb1spGBjYO8JrbmGopXTikPmVewkLH7hz6HPxpr9q7rU/a6joN8xzaxSZqILl7veHL
csWFYsrD4eSRjjDv5ZPDRJDlBWfYrYJ5aPEMMEdPGGZGxS30VEzEdf3V4g5be3VOsNbJ6jdD0ll7
XL+bGuBJT0LZOSC7nJwRIKMa8RCq+rZeIjMBpGZb3RggpPMwNaFKrOSEMxBUiPSvRfOb65dElj1W
PJyDOded5vdKsl2lvv2LS4FwGfZbUco1pzzlWHcY+eJR9IF2vBRacssoMVgCYFGKucDJxCZen6oU
avqoAUxlmS4IbQH5PbGMoWtfr9KMN26uK6Cwhwrn2BpViMIOva2j3688w6MaUf7g7r+3mgqJI7GV
6rFmWv1kwQFvXc7rlXaFv9u6BBzXugPocrvIuaqTcR/8TPjZmck3SGqaW+iNchl6Uk1g9N8wsQRy
cxU9eLVT+r5i1GHv6SSHucILMbUgO8R+9NFI59uNdZfUtSwel6+c+9gVN0FosAy5DYuc4cXJouwn
MqlQ8XktdqO0c02qj/pvkO0zw7TaOnZHcKfBnSGAtlD0Hm1fxZ+3DfGIpwa0H+KHDkyqT3iNYk7s
w1uSTLgTy+Xe3ulsW0aeiHa2t2fHUYfchnBwWioYYg/UbJDeJwFADeCSK04EwhkLKmCFC55tXktV
/M8/GoDSLFa5uHgCyOqN7CMxKA3WzreRQWFQN5stZzjYmGwUdJWSr5HkM8Orfk6ySdxFjBogVgMo
TQo+of6ZaRdJa5KBGZBR6fXqqXBDlH8UeyG/ArC1GGEo+YowtUNqniGC37h15wPvdmKIrAHaBMt3
WGiP7oTmedkDBkjswJqDAe8vskMoqglh3tYZSNZltMnzSsEy22k1RgApFWekcyXeWj13H1dchwmM
fCxyfN/fvCldfdgA8tWh9NM33UMcXRUPD1AkC6nH5HT2zVfFxHv7Wwaub7shNluRX/qkZmD15U7/
1IEQMxQ7BIDs+gzQBLNINcaR/vje5gUQZoN4Y4tH3aLljJoeG4s/yT0hb5f9x5XnLODOPdKe0Cv0
lbwKOlqcclBx7tD1LDR2mV0ap0UZ87NX6GMgQeboLFUixSsrcUyRpGLDQ15CgEYRRms/Ekh/+p04
7EdeR8t007xEA+F44V9S0N2WdAYmCXwSer3mSbjrtZF8HMIdS8feMIc3e9JbPyhuKwxThsVjxWYh
FfPZHNfSZnx0KhWI7lOUpTF12SHmX8DRuwouO5i0/VockfAfNaWG3KlAqA78KMX8rAa3rOZFTocN
XBPqh/n5uG1srZfrjENCsjltdKBNkgt4qiTFXqMbkg1x2JBXdymhzGwlV0jVGZf4ZkOqgtFe1o9I
KIbxmgLi6H2AyeeTjKMQlxdwKjz8UG3vKhQ7cJE2QOXx4cfJkd5UXNQERNue2c7zikHgQYMrw3o0
6qLNDWlW4grVC2ap+um9VQF/yxkyxYO4yKahH10cwu9H1bMk61YhcLHsEGXAsMmbltGzS3vAZ55g
gHB54PpqBED/HLnA2VnWScnz10wfusmmdpAiIsN22Nv7oP1UNWa72yMZkBmODefdH5SNODdk0afM
YIP/bABpyTELUXmiGIngVc47SlZpyM50DzGFjcfAMDkYJ1jBKQf3CM9YtZRF973fy7eLiAXcnoih
yf2voSlHXdgsAt02ka0OX1OO03GCsQsDl6p7hFND5wvzZYBBP3G/7ZmS42vYrPfDJrDXHVVnojNI
/4nZObFWl5bvlJDfq0zywlfkAXf2XHAOoA1V2nDKBtoZ2iUPKwEQ/zBy4CmvkgrYa1eCIkUWghqa
JFzWc3uwzjmLIke/ISSav2Qsrzo7yKE0+tqOQ3d+izorzjzDv27Tzum5fRrDFZrHNgOl8dWn6bIL
wz0Seyhb8Dd0sZ7+DC95XcsS2TxbQJD4Ije1PMgDpwfx+6G3KZo+DfTFq7fiTvMXFc8fl9NB5f0W
TH0VpWKGvX4qK1WmMi9oaiunCNKk5CdvrEIhE04BnehIpHf4+5leVRsHukZ8ydhePQihujoIyl6O
KyaNEb7dgcxdsYpZYVKMo9+C1KcUyZYUiNi49SwmaP+N8CqkFat1vuGHyZoDog9j6VypEGIQIr4z
qAIvWHF6A9RYCQ6pr7yXni4eT2e6bC/t6kXgmCv7Do3foeJrMPfKlA/PHKmJ5AZb5eUcWQcmf0WJ
skITL8VmhfzSZxIHk/6hqf45TIznhQHJ/ahJpQAnCxDHh563iAo3ADZ05DqToWsaW1ugJywY2BQ2
LsBmbm/BOFSbTr+0JzAZHzklcJqPz7cApLdiCdVkgVPp+syQ4RasF1yFmxiTmrn/tDYEJrqmcTdl
dF82Z8iZEpllozNa9BFIE7lfVDh0lnGbuVLkBrN9IGYug5nUghspC8CM2AImAYkWmxYglo0LN0YP
QqV2QiR0UDkI+uOxEFGJoSXIGtP8AbquoQWE29zxJHFQB8FC6ofFJ16TF7ub3BdOFXWLjbsrPdGr
27wYDzOMve7QW1CAzfmfxUt73TykXkqJ5a6y4ALaxjtikol+upG20LI90b0g1xa9bWxY6kF5iWPS
1Yt2kK7Pvn96sr+T23FAFF11Vm6PBukoQWDsvZ80MWw4EaSIRswxABfsXPRg6xfoCStz96iZvC7V
WdONdjjyRasTkK6QGyRuVAcnT6F6145w4puHswGWcSHiIyCZ6EteoBVE0Ylo3bt6BRDrgns7z1TO
LYpmw4ifqNvtA6tINlAhcAsHWP6wP5fqoKCPwwi7XR90Vk3V8DnOCFShKKgJoCrDKETIy4Xv79md
5fKERausp/L5UPsPCYEwEjo9I1O7YgQGxMC7Qn/u0XnUSnO/YpsCZEpsbk1SLyGDYBDGXFCL0EEp
xCocdUizjuG1gAUiu4IZdIIEvObxxrAfVhdgVLHbSpmKNbHtLqyWE2e59kohKPAUVADOgxKeUVWJ
a2G9YJaZ5BSfL8WXvSrueKSr4Pd4PskpN/QVMvMg5SSBlfQDXJsMuMP+CQp+ogGBsS2fvWsQGRqd
bAdXwW6R7MZz3woPYsAhGszH4D+zbX85hfQdI/ZZWZ83E9hzFhBnHq+JBawd4yWKijFQb2k+kIQA
heVijUR6LULhX5q5/VD5eLspBFXyVfl21pyH0GzR8ashxqwA+42z5KoHFQa6Nz2SjugVszUR3iv9
nWEjOLHmpfK8gYoXc7aWmk6CqgzzzmSMTjczpfyrFzdL8fkLJl0teIe/o0oa3NkmO3hBy4VDNM3u
88m6wN6AWXoebGHScG3XrUZoXkJqTXaICMalywkqf1cSexgKLxYiEhCO9nJKRQetOL9SXkt0lvQu
RLAu/Jl5TA0ZxuZJdMA8WRXn2gd8o24QHVWRVe6R+kuNONrKyO44M8VMvmutvwtkw2isBThxNuAN
TVLqEoMm+fcTMEnfqCDuLYb/A3tmkoseE2QIY59W0JuzAZv224Zy5vyzhdv/XHVpuyqBSA1hO3yu
AGW5I3LSXiV5jtPI0CsAQkCNcuLhp4N4xVT1toxUOQWUmZoTrVFhOIdnycTXiLUIc4QJ9YTIxtJJ
DMHhVCjnq77mAgznHMp/VzfgFoGiej/n4+Mapqo/3Cu7DlERrMkQXtXY7BmswXmoUlOAu4H3vHD7
V60gY+kJXQMzWy07h7G7IBkXMhghSmIpIgtrKBi4VDMnkQeRjVGc+5skc5C30vPg9zFOBgugnOqv
XlqUHigG6NKs2SBqLQILreTIZAbEKBupqqEUzN+FYZf0Wk6Thk8keZ1/ysiPMWSxKXvFq6dF/O9t
kF5yMPe8hrzNXbp2RwJNwGmSgnZP0B45s0v54/ZDp4lbbqizgfEO+EC7TcYyGt2WXZOIlQsKr1Qx
bOWQjKOAi/Z/YANgVYlfZexdrlBj+2D2PvdL7ya/koZ4PPYAJSA55zX3DBzYfy8VGJEtlTv6896M
C/eThy+btb4di/YoY316LNrDdNVV6N3HoXqaYN1yGWLeQl9ZZ/x8LnGhfX+fcm3cye+RRk+brwm1
qdPQjrXXAzsZDMYbeqA6oCTxrRuo03cws54t+/h3GI7EZz0e2sxVTOppTJ1pDGZ6X/ps+8GlW9P/
uCw044chbadWn3QbCpHt/BhnjnkPPh2aVaVSH0sqFBAkMyBR+Vg0sD8fJvaifFKtpOwJTodLI/HZ
3lzA3+JY4lHSS2TpdDIGWL/qD7bWjmNVzsUEGFhX+IplG9yc+8ndEfWs06dC/SWoLZOjNpvQ9FBz
1OZpfbSF1DUywX4iSsK8bTWTidPrgwLH/deN6PkAe75SVWMRPbqZNQbxLcb56n4efpXPrMIw9erd
JHeWJbOkLKOtL5jG6l+G8xON8Baxontead/MXHy1N+Ykzu84oZv/5GROMT05kn2lM3G0ALRf1Dqw
l3Nn3aLw2wX1xCmZAK2G+4Q1IMXx5jzys3e4bx4y/2IIbLepHRpyT/nP7P4xDu5y5KT9mYmLk9fR
zCQnhmvTas5FkICGV357UcofWTKSU5sJk6sQ9WfBE3huTgXicxDic5AGqd0J38ALC2EVN3USIqFU
BNeVyfK7kdsoFAMk9fD1zZDJaW37gGgYdHNje40KPgigvgd/byFveXtJUhWTByfFe2wLKTWc+Zsc
kObN2vrnNUo3O95CJWkoH0mt1ipJFh7TRlXF8vHUZ3WyMQ4viX9UQTNIZJLi4HvJRArRuLujRKAr
dJqVeqCESu+DDAlPw5rLLT2GxsHZv+cTe2/+DCEJaHtHYhQFgVbAEQLnyK1KE2MWUqG9yFfAyVd3
FKwwySmtWgmAm+/NQk97pk62PwoiZqWVuYKhTDm1X4aZPU4nJ7Xd/QcE8m/d4rciK/8PsF0j1NQM
g9VWFhH1qHJXzYuAbZp+E1FlqIpYqN4V+s1eVxa5NKh70FlQNvuyJy+y3V6PbYQceftbhthD2tB5
+911/BqI8EsOHcRK+w/pbo015uxfYqPKr1BIX3o/9uvf4qr3zu4n2tfGprhDIWxGM5S+8ewdiQBP
ajYztKKGpIdaR/B3xNxZi5C2hUiX9ByQoVZLv3f6e/hFGof7rLcKtsQ3UCGa79/JtxCbJFNjh247
VJH08thB7u2L3Flp8/6173w51LuhFKHu/8BQL7jOZFEId7QQ+jvOWTkmiqbL//cIK/MouEL+TodQ
uN2W0yvwtb6XIJWE7CdnxUhveTGtyH2S+OKSkI+ToJM1qt8mfB/3y0yqOvC+HYV4wAT6Q9EKdoHq
rnOpL5U19+aYjLlkYfz4cHNIhku0qelvdfQbnAmOAERVXGO/9Hp/ZkOEIpWAO7YT4pVllT50rTgD
SmHxQwPYQeqiAsVy4dtel3W2nsdlNq4EokCWWhcDEx+ju9DctLLosbbt+11Q5Vb1qs5jbmAHPPHR
p+146IXjiu8FeQwOkRw+K2Tbz7yCGrKOL9o60P50ixomqTloV1Iyrfy9udQ3zsErJSfjTqnxZ1vw
iHhD/1hA1SZNQ1/T17PiMbndM6jNtRAyOKJu+4LGpQ75qyr2TodWSdM/ZnPjJkpZlIFmitGH5XXp
2fH3bXyX8f4x8J/haNThMHtkoLpnVwwvUH8qx+w7pDMVQ+MA0Mw3GJjuEqkritoyWtUcDZS9SDVo
96FRZ2HweRRiFMGXXzJTl7YvRpRP6SoDBLG4T0t3aYlHYrFqhQ+5QzertRl0UGSQcsSbOoWX8j/N
4EfG9BJSljRofIYUVEHvH95xKmgeL0Ug/xW6ztM3dWAQP3JxwuM5+Z0XBx7A1q87EqNHLXNh6tzv
Mj4Y8kgZqZ+276v4CUr+FTrK9fFOViU/VbT9AH1mx65pckC5KXTOG60EmNMhberEHvKS33L2Y3Cu
umpZ+cqP1/7nwSGy8lzYUfZBRLHINtn0qLqPQl28VzB7Y8uOzY09ziL9eCcUt3yZ+5KMobIDTC6X
G4uN0qwhH+7rW+CcPSEbRmLjFRN1xLaPb61fK3uBAdxkjt7eAfKVFb0zoQBo41RV5Qqy467eI6FX
iFClKJq7khMuqqOuqmA8Zp7w6JQvo8Xw47n9+1wNSG7HFAgBQsNlQFKuQ1abtz1KdIGx230eUZsS
5e7czzooP5aFkNwMfB9Py8FFyhwqAGfUKxeOv8kjPe0jIKpoA3qBik3L+sh54MyqknnbvEpv/qkN
QffsdjEGxrrWRymEyjsuWwa5vG5/jvHWIkWevEAAJWUh11X6C17NNrmXhqeg8Vr2Fhiq/0ujGmJb
B1NB9d/fQotu4iH1ui7BQDSa1bd94UgojGDalruPhbTM1s/jOYy3tMhKkyyDTtAD9ewR2h1fQL4X
S3WzRY25yMhhMp6bbrcldwAb6cjUgOVLzxW4J4LRtvwcO1ov1PPCPDlzOKjzDc/rQ2Hdf2WQ9UUp
tTDieJlDLj4yGrBjqQQZludk9qFItUtOaCz6hVM4xodtl3XxV1ChM67TGTGKAyJN9pZ9Ji/Nomr9
mrtjYXGi60hlge3X3f9fyyLE1VgVB7XhOd6Gstv+XPHJxZeG44RA6XfgXX7KhpNyPyYkyiCtUwWR
CN+CAtN2TKJfbxXMMA339QxiC4BV8A2lMB4jpu5n557acJ+HVKDYn6C3UYHyvdYw/OIl6haUhdGS
ypSM+Ho70lA++ML4uucfn9Ad2154maPezErQqZsyBtcCwH+UMNZ+1lvv/MHB2rYEvFeMtfmGaUK4
WgTPWkdvTbhrVwmsdCC0IOAd1btP6IAceHuoerdG0ATWE/GZs+1cuEtRt6FSu+wL5PpcRo5DV5nq
Z4wEqlpNgO5UAKeMD941ix6GQGRIz1WxSj4Pa1J6HmMMh3cTN3zdGXQ7DR7rJgmUODQr49l8x2fo
mxta7Bxw7UW8wBAkzLsL0/j48dfpAWDCZ7VJfHq1JuYec6bv/vsh0jPSFHboGfaJy9JQR+QfIk3o
+lE8XB9I5Xf4BsetvokqSstcf0hTCTrk2DXhErzplVBXmnDKpR5F8l+1hEKjvClE6a7simvCkI76
Cq78Aewi1m306F7iUP//IDe0tOgEwoxbHLNQrCg/vLMQzQy7c52gbBS2XvpZXWKdszv/2mUE8cit
HlidsWdE/ZlMZGwcxhw/ct1KPcSvr0UF7TdkwBS6BFyxHy4Rnqtt2HF25wAAnNWrKjinaj1fFHLG
J72ymS4f95N4gsVCIaMslEZa2RNSD23xyyfz3Z1fnD5Fx7wbfJOqO9fhh7KJOtBRpZPw/C/AYkZI
jS2tHbKfb2/6pHJIH0tSB7fAxjJLg7kHvqxKGFaltGg/2G6fEYXx5VYykAppgLx12lCT9WP6s3Rt
FL2ciVrrN2L7PrEsHzj6tXOOXBByG5Q0+rQH1tr/F60MyZAla8hUFnzrQRslIETvv4bng7zMTA8W
QrOTWOix3i9dfslK+urclL4O3LIzy+C0iuyxwMqPcRlh3seEVgE7bh/swyW5N9DsQ+sOAArMRizh
FBRjxL/FZlIK5Z9vuTfZU3qoaOCUYWTpuv8I7UuBvXezIK25J+uICgoThx+eVvMRcM9WoGx4UmIE
/ObCK5xsF0glSp9WI1cGTtL9Sf48DuS6LOOH1EOtfYtjyzYYiaAqyvQuPPsmtOT2MlbWC+EbKMvS
1kliz5s7UUvSH/mxJrGUlr/5iD787IGz+ylF9pSR+W1Ice/TvbhnGTZ3AN5ZdJybbBFDmHDbtMSZ
zaZRcj4Ls4+ODqUVQK+Y2WH3lQ068Ghcgqp9kML9hYcW4OzvFjt3MnNpUOhroDL83vyQx9EEKsel
WyEHzBe7InPhXIyeZf3EqO/yOP3JnolusRx81m+fkTRR+AZEpVenAMY4FRkT1MgaknEjrgGnGln+
OcF72+Qbzki5c3rTIIcXd8b1HI/hsgtZnhlrGshvw3OCLijfEUIdijlMms2H6gcVD5SvUcL9rJ+2
iUbCooMV//NwP1CynH13sZUkPU00xUM9vgAj2YujCz0hg3YPxebjQOtuUnzyG3ojtEBkqw+/pVxa
C6bnodAWoirppK7J4lbBHX+rqN1ZWg0WAvjQP7bG1exX5pPDxC5PUM5SSk5JudW5CQaa098pBMMD
AtVLttSev8pDmmjQkDCXU9HMcZaIks+jV8bOa3OHGwL4uaBTuDXKFtv0Qio/hTU221pPaEIFU1GS
T7U+tpYsFDFSy9ZP4tOJTQ9KilrZd76mVRbO77SQ0vcQ+xGgLRy3qX8EacFiKB8/0HkMMbQ4a61r
Fcas98A5y7SFAksxtBYg80C0+c2YhvPG5iMmbRiWd63lUvewsOdbZqJOupMXl4IAjKJ/VJU21Ltc
bYXLFHuVsGyRXCWnPaUg+yvL/cV5g9CUiweUFn/ql2FZDeQQPCBZwr87VgXO71m4gJKXrRP3LCYH
6LKtDl1iEnvWkQFx0UMEc4cni4ZOt1EOzdP5ZY/0nHUEWU77LppejUb9NF9h7gmDHPfeonkiaPGD
wqBvQ6Oo08Svyj8KCyCzkWFzRKmXA84FtoJ2etOQjF6uhLjd92kSKYkpop7NUSCDDRVhpiOPOkFe
UoZfw7HyUdlDrIRzHo3PFAdqfyiuWRSPYAPnP1SPyqBD3TiXiQ3GYT0hLjOhQZsjkONIwnUs2WDM
YxE4yL8IB1LeMi0EvkithT6SRla1VAyO1VCVe8d7yC3LCSMFiIOf6Bla47nvulfDS/0Ktemmm87D
xUpbSqkaJipwOxTITU3ULsK7RaUzTn++gwwrvT4OC+7JeJNlm3Hd9imQhOG6hBPuG10WidJYQWJN
gSQ/Z42PYxrVdrvxZgClSHU3NX1yifSxqaLsEbrp2vcd9SVHuZKAi7eQFNrkcHpw3Y6OOpuXfoyi
k5+QiY1ry1GE5qu19fK/5LUEYg91pNNTVdbdO0cyNug9qeQpjoiVqmY8Gsh72TVCXLZ7H8iejtg6
LzTB+6HZpDKoCREXy7TvoqUaI1kxfJ7XrGg2YJlUnbeH2rQRyMwrYjVFe/IZEqkWxJO2uV6b44fC
FdpYARX1e2CtEL0sP3hB6M59OWOI7sX71OZdGQ75LCjSrFIJjlshVh6PoERPuZZ7ZjhPm0ZUL6tT
v99PdcNEnR7v2BuiNoB0NNI0K04TnUihtvcO9Nb4AUdEOiTpyA0uYc1OEicRTbd+wYEisuYz1YEB
kiIyIBTya6h8+/fczTe4Nshl1QuylWIRhfEshz56o+nGdh5DScp0R4Jn/c4a/u1kZ+Y3yySFRDCM
OCOztAB1E297yrA5yGXnWcPlHUrUuDV2yB/lMQ/pinuAxhgMqYfRdlyeOAjrTd2qX1XJWOdNLNeH
nsk29twu4oAfPlPgK2Ghc4e+x63LG/l1aYDU4ip19vVPmOvt0xeNB/4JTGHwbygrn8WxLN8B0lag
F2JcZeSwtXZTtf1hdQIiCNLctn7Co12vSyZ9KahS3Lv40kouli3N+ctr7MLP7/gH0uubTC6+gFmt
97yVugb42IeK8js+1fCmZhsZYpyICCp4RXvq3wPpl3l6n78uGPJ4iErTuKYY2Y5/5uhWqZ46YjB8
0C7NiXa9dHF90f44M/0bn70YhqB9plPGg/sJ/P85UGMRh4/weyfo0USmIs5fLHKThiIdUckwezHj
4Kn3lRD0NynXvodExx/2lSH8l2x7g1IzvhzuCZSuO9mXXxOcY+P31JO9avMeYgfbxaPD/tuDJZIJ
rx90SiqqbTUEFUdemdCB7oG3R0cP7yOKBlwX4aT0DnCczYLdp9Lf+d6nTg0M7i1mA6oI1pPXyNnn
7zvLmJhXRNIeV1aZ39Mx9wDuZoJNOlkCIT5/d9EQuxINamkGwcwdAxezKn+Bx22J5ZhrJ80rbAHA
ueGQ6bwqooB0IafiG+I/eNiEswtLrvbnFRiKiKVQkjvazmq9LG8LkmdOTxnSDMKngvIQ2Im6oliQ
PCFJlDNOyJ8e6H7RxKNFe+u3Zj85ywzqjy9CmHl+QhwYsKNLiJGzoJcUuUGPCLTW3g2nJOF0QPxy
ikOVkjfXWcul8MBb/sVLpKPKQOZck8th9px2c43DrJ10iGxZzZK7nykrx3Y0q8gZuOoM0WlACxqj
IxyrapR8vRBZPE6YcoLCb2X9lKfgGYXc+vWIZfMKsayp6dYuFPbucDtbnF5jKOAiJ//enTX8x8yo
sLBf2iiipw0MA4Kr4pZryfKM8L8mT6wfLv6BjHK0YBFLDL8imwveCqRYw+iq3wUpJcQeTPMnnPXd
gKIxkZ39AWP+ogPYofEvvQFXH3uDg1ILBbgOq6tgxq2rY5iFHWMedTHIYT107AsIHkKaCUC7KOEz
iJS7xx5HYYvIrSGMgInaUZDEWOE9GFlDqZffdhBnYRzZghaeEmdrNYiXOSPJJ+KIRnDyPlRhrTS2
lJDsyPL9xS6gCZnV+xxRxE2mPjI52e5/poUbI5qqC7qN7gtZDLL8CfP3G2/Go+ddakczz0ZNUzZI
wZXfXhbdUcF2TKON38MxVZ/3KE9XIFVhS/gy3kf5ChggWVhLeo3m9Wz6NATz4nAIh+L6ofXSWi+E
cxqy6HqQuzFMJydOv8ndfQtTb6l8JGa5g5Q9iW5LIDVpewsQ8Jskm9ZFfw+3hL33Ro0u9RlAL0J2
CexEII+dzYCfSKgonaGn2dwccIn9s0dl1gC+bwBP/+u1BgSGkPgmhe0NmmIN+CaMbSeorZvSw2iK
GgytOyYONyVqo6nWBiQrkscMvc/XVJFUJIJKu2ylvnZPsTqOk4d/MYc3B/cfSSBeBecFSQUmh8i+
pk9Tsi735ZPdzEcYooD4q21z756Tx7QtSwNUIQzYgOPwtInsK44iBLwpGc5LDesFU2GHl7v3Zgp3
M4IIE2IG3odrB7Cv1IZR7hSSN1bnlXYfUWZJIA+A0oLipb9lbA1toLlJXtXi2B7izvmpO7AJy9ml
2tztVwy7xNvoRsXqkHvlml8yIvm3KYvK+SnOh6WPPIvXIPhNyAOoCp+2an/RS60hBTDRWQp5lcOW
uLv1ChtblgxjP0GgRixAxO2vKY/J5HwOLMaogCnQkR1gddd+O46ASMgKEFuegfWtk8ymj3GOMbur
AUg4kXgZ3y1V03TYYN8H/IPMgjJpn7Tsb7dRELe16cgfUMkt2PYl374UCOuQ3Om1RSwgt24JwUNK
CJALB2r69ZS2wqJHb08UIyg4/13eig6aiRC8jPWl7UR4bGfUYMV1vLxZFZY6k0W8EDXuwPD0f1km
yfIUtrJQvrmhKFIE3YKtEVC7yRaPD1KvWxwi7uJb00bq9zfw1V7AWelj1JZil+6//fGbzLVQ/DLb
DqmpN/j0xrJEQ6cg9hF4McokvxCunD2Qvyvapftfj7ddkQtpzLBsKZLdZgoI2jCUaUue97AcMfvJ
FQY1ticUfLL1iKHWCkBqZlAgjLyUuXWXKgPdNbKu8/IbFzU2RPz+8aVsptfHsMKMtZjiYE4z5R7e
3tTOu8hQBK+vwfpeiDJ2SNATqxC7J+0KMVOysYqut7yddnKfeAH7UldVLC61qpL/N0BSw3CVj1bz
Xk6qH/RuiTTZRjroifdcVY/hDglhVnKe8m+hwuRKFj153lKt5G5+/8wjFJ9UWTvDtcGhwOANgqC2
rhNIcUjpUd0LwOfFAjkT5kxW9oR0JHainvl4Gp4u15KzWAHODQa1ubLBE8IxgC4qmJ3S7TCha9Qf
GcQI9xg6oX8MvZGkIlaVb7HEcPNKj8MCwxqEylVL/fz2zgSHnV9bzaimfkYwuNxvonmRt28B7fwn
315ZjemydhFpUS4ECY2Ew7fuqwwV1+jnFDCLjTlGU0D7xVqFvq8CfkSelbi0AlcAO3NkMee/CBn/
aBTgZGt9dtrAIbo2YC0obLzFTEy6Huuj7ZKwWHHtRpmCCa5EMWwKWGunM2LZXwZU1LPK7rUwC5IJ
cHuVMzCMOS1LUHKhXbVTd5tZUF0gwRXXVqEND57v0c3dj8PJUL8IyfVK4b+16fJhToygL1VBYowS
s33+PjLZjQ/5uJgdoUvGCb5gsALuRl9XH/cZ9/wsSV778PODJVj4COVxwdLHQpxDaljxeOO0Bn/6
E+Lkmxatj2IFo5OQIlvUy8/QcCqTJDOwPt/ovagdZ7Y4OgDutngCR9jEB1iNzWHdU2LBD94Xdrdz
zhfyMnztUD1djNE2wHPSzHtpD9c6opfAPNWp5KG6n1E/B3xE8+bGsBonrNWE9yc1X5nBWlD0C01N
vB2ooYQqwLsS5pDOfK0oJymSdDHezz9M9FaRlhRmbcq5hYZ2D6EJRwlOFZ05/wyWRJK+xxL6VX5/
FKCmXmXZfgOrRmoUmAU6KRRmYUq9COjgxo8u8AGgMkBVdo01dfXv/F7uR98rr8qKQasnid2DAoeC
4pZKMFY1oGA/6tdw4R7AYIyoBobL0YPDgI9JsYDn7+5hFMJTWrJd742xLuCM9QlZGok5H4x03sp6
IDBgfRRZyAg8VRnnSeAI2JRED5zMvRJNnjb0RXuGhuPJ9TZwEpfgW+6x6K2NZ9eZU8sgI/ljWUlz
qGOT8KLPJqRQpAX2lxw6oWisYHh1MCbpxn3FlN6YGz7DfiwgeFJylYhVEiz+CPzyXpQC9NqCYKof
zkHYnOxlmaMeZdoFI144VwtHpCZ27LPpqGZtkWhHaOVwbVj+R97WuCYlmLjF0SbSlRANO3B+uabO
fb6O0Ke5KIFIH8LMIF5tfviyX8BMzZkIhMf1PQPfqAGTQo+4LMvOBhV3MS4AJUgCRJ3vUPzxtAEI
3Wo6SEoTPxx9/j3ZCbVMIzyQsTTV+Jntzx76GRWvFv6E+4Wf4eW9s9NZiYNSxtx86WeqUSJUsAIK
4sfedfO/j6Sz1ep8r1f890EVbKm1lija1HhAYsYGU/RE4F2e3Po6fzQ6CS+n/kiZ9i//5j5K/lDF
CfW9D6kPTD9XRCtwce5s4/YAnDyEhYkE8lb0gx9EDkG6dp0RC8Seh0mSscG75bShhHcT0aCTIEmc
Dv6Sy++BkzXgZ1RdFW7Sjls/NGueG0tYB/bSkLBmvJmryxJrveLdOEdK7VCI6Li0wZMWfSMxMqho
2/e1IMMahB0ov8tpjREXY91mZCj0Ok8y8WWc9fN5GQ/gbmVuz768UMwes/mebtozmCz6edgcHTiq
CVsC9VWOnXGVtYnpLMOWaEqnZd58i+XT59FsRBBf3MqK+KwLEFnejjEPD2ZfbpNAHDqJlnKfnZiH
W1FsVO1GEEiXHaMFxMru1y0ZnVJbTSP0/dtM7V6dN3ynh1vWzOX1QJAOdu5+t+ZrCrkUqlyks0PQ
aaf8xbcXA/Zg55uHenOHjnbNpQDBEZzx4AT2rpjhpwvJ+jRwFRtm3n88xSmNsIctpw9c8HmLsFC8
Yh7u2PmCabP3i54cVDVmCOFE3R2Ostk4+kmqyE9tJmeexC21uSLmuBgAzsfG6/Ah2KgRxMw2ofus
ZnyznZiFwOHl6lsMD7zYmkElEfHr3pg1EzA5uwEdbMwDSTIgaTXJULVjNi9WT5AYznisfqkcGXHi
k0C2Atn/HGEjlTGqOaXLOR0WamFVdOg+s9YcFSwHC3iogOoDVMa7ih+O3Cp20c7H4W63quG1O5vI
Ox5V9sge23zDreBzoTP4QTE9x1aXVtOBUrPNlGPUnmKojRi1xKxqZAexTEKLu1whgt/KmwnDA3dS
JfbpxMacB/sKvDj5svhtak4rPhRYtVdi8yk+TXhGJV0vP4eCMjo68hCLR2ZV4GdtDSuLtXnrKvxp
D5rBIG9wbpCkgLEHixemMaoSNA0eav/OVv/lih05Gs9aVHNdX+x/ORCkjYRCpjghmrNDovsXHfQD
RjgMibyrjxdrVJSP2rIN3Hl38zAs1DiId8cRdUbfhPMkpKTIimM5hK6rWbDU2KsU+yprNOgvnfqE
SDecJSRdNEMJ+PBjLrdrzMEr5PHrs0vbjbjNySmho5fPJ8dl0yCEZhOBc00XG0MPPQK6yblpgcOT
eTdEcvHngl6ZCsVEmq1aPgJYQF1LX7nPy0aglCNEdWbqa5ikQguzNgy2WkuEUOwzNhJw5RQ9C0Xt
YPCUf1teeakx/3e9+3vrJN0Cu101oivvNgUQrzSqdm3D+JERLVVxaE+uVacRBH38L3C1x+OovYSA
V3LV0y8K/yq2VosihoNUeHiiM7yrDTqPPjL5VWxV5oItz9Yx1Q0rHwns8lcrfrqYPeL++bCJra5P
mF6UfyD4H1W3lcal8yy4t+CTYlob26rV5Qmpw4uCQepkTyiZtptHWJ8554+Y9UTTxYQ5oa5ZSIIN
NHTVS98ZZMGpyYJHM8ABlVwyaVA5YboV37KgtSKnBjEmvuq/vonTPcwRo2iROSk/R6ZJv5/gJ0oU
b7LnQbz1GhbDT5kXHWniU5fka2rhzZowV89IQ5HNRnVVFCV2wzCd+PobYlcTVOosa8M54QGh/URM
BG/LahtAYmhKXWzIIubdMgegyXcXncz4KE4YVmyaqlo0A2/7DzEp3XlRbyLmxKWgaislOerDqJrh
GnqXmDYRSwgrRhwSOTvojJyioYW3oMjtnjGhtsvjOgqtEbOqBCQAc210eY+v0ocGfA+PjHMba0EG
1On4an5brkGl3AcaykQtEGfx/FzoqukXU3SFKGm228Z8j9rR1yfVjY7TrSP83BAhJa5f1b6NW3YO
puojT6hWNHpAp04zGo7z645VS9LEAxzpu0nRVq/+qk0W1FilBazp/BCY6SkDeZUUfw5DUFaKwcNn
I07HnsLBMUINs553OAmeuif8rCTKV7YN0DQnV2eKO2HpczPozTAJsAWBrusbL+Xj40PHZh3YR1kO
tBZA8ZjGmh7vvJ4e/Q2HZ26uiW2TKUwRA4a+GFu+wnS+ahYbPQmR+bDRfVPIDQ1JLYFywNg5rDiX
6Q7k8VyDiBV1r27WrSSxjhf0c2DELBs5CGx6XgegzitoNGFIRHUDTziQlhq4NST6GOn+16FghgLR
3v56QIxopcLTtUL3mkTqu+I9UctOVW/SHqEXDYJcaRBFdTA3P/c/u1TVmZI2Mh6JPYhxDpLKzpyD
f4nXRCDX05M+BkMDurDbjk7J9QKNqZo4h+AgWoRPQlNQS3IWGbEYVypTz7dBwabAe6bu0R01lVYZ
a3raXTvDbtSiaEOs/qZaQrDzy0miRZRguPq7MfB/lB1qbeZsIFFLim1Ge/5C4iG3g0Z5h4CXIaZr
Sro4KDXXm4Zi3ZcG/i9+4Zagznml+AcPB9/ySMba+2DR3fLcbBVDxLmKjMUGu81x/ilp77iD/KzX
E8Qqiq/vHN4KDGqv0LFP07fjGbTblG0sFzwvTh0cts48YdzcCWsq6CsS7f5qJddEvWh0gESP6bCy
swN3KlanOn4AKcjr+yboZmkZcLBMaIFFAf7zkBSqIn1OH7aBzvC9xAMipxf5TpnhoOj7IWuoaSEk
m4Ifkm1vqBPCF+bPymB6rmFbXE0yfOuRGfRcR5+xb1F1ByqjqLAS6Sv7YAMVBuoKwgaVbBWYrrOH
FBsx9EP3HRQHTM416s+Idz+EbqWIBf/7K6f/EdTkTPaBcB7VgEopjuftJsasORoP1qTn5a41EgbA
X6oMYiJMTPYbxxJklI4c099URae2hbYyZBsah/zVrB3el0WvP667cgRKH0V3tBeE4kmZhUIBO4XR
g4m2qniFBx1pwJ5E5oHVEFyn8DuAg8T/vaQBG9Aus4Y1LwDEErXJqQw5JK7jIpxiwdsv56nIRpOI
UAOP19sq2+tE452ftXf9YUAul/qljGgZY5dvNDnVCVT34wOineoOzrcNZ6kk8LEod+RyAXlrgSMu
3XkQkJQzfo6pznbasNBG3T846TmsW7zIWpoetHjt6Op/nu19i59rDGV5eDcMKSx/NX43qxpWD3x2
41BQdqZDMt0qujmxHJGVoU02OTr9pSSVfburw7bYA7SiLmL2jNC4VXrbTIUjl9Mj84GNaMM+ydFP
fgM/XcSqfxGTg7ALBj477wGj0QEVTaN85RiqppRLHWQ9MXfWORC2GqfuQuCLEI0xhhDhqJSY1mHq
U3GfghOcEUiM4uzxCd2e+mK8NjgWC44MmZ+zRiazJRWRYEOJadGxhr/QCe2K5cavGUl6HMp0fxVD
UvyasfD4BOn6+RsuEtny5M1GBEFlHnZe1rahU9tr5MJFjLY01AllBS4gViIFNa+drRwUh9m8OXeP
L8HypmABaAsOt99HpGYA+Q7U86E9TeOmcj+Nbt/JgCFuev5SmeRTeMeTpiG/NvERjXAhVAn1S6td
IGsxw4nWRz/Ly6UTZ+Nco5wY3tDXw8s0587qN4/r/N9THXeqFxE45MRDsBT1/vZRtawkZcftMKSb
1Iz7TpMrK9hE46STtsVTpb8jWJsEvfzD0mt2PJxH64Fikn4kYsJ0q6GmW/SqjrgRlAdlvDZhXyMY
GRAm0SpEf4qpkJDJaZhyWQysyuuVcEfe461eG0McyjYJGddRMWwqXIXznqRMbrjcS1JuF4s6bLJW
/vVsqBhR3SWBZGmbeJskn0YbQmuREivUZFbfE/jZ7vfu1rtIs7t7NWfbtgbx6N5fnJEsie7BtenP
oR0oJ6Vv4zncDmnOzLol1ZsIbYDBFl7qsJhgm9cd4mSkl0KOE6h2z59vo766U7QCSYr/kP3AKjp7
yuGCqmRCjMT+OJfRCv/O2aoBj4q2HK0Q7dr1CgWK4vAUPfJZIJ+ZTIwyDEq7UPx2oBJZOcDko6i6
zlvih4ZYZEXMm9yPV/PwR+vneZMGfwNguOKFvDmos6511xAvznchi8dA5O0Ty5gnxSSlTGtKUbDt
jDA7hUJMBctaGaKQHXc252vjdjVLSyWDp36wP2W+Rd3rI30cWmpETgnolipAGI3g2Oi+AnH9liH9
PnQ72BsxBMuUbB2+6UxHDAPBBMj5Imuwzrv4FfCo33CwHrL/itVFYxrYQ6SQ1W1Xw7CjBJ7H3ojR
GdlcVVaYbbb6FbwHfWCp5zFvKbChsNkMYp99aXluOueaujFlT137sTCjoIuaQT39WDy6MQt2nMfB
YYu8RrkcZ1F2nNHWaiz0ketAb8dq5dq02VCX1gHgZGXFyq/3NbI9VI9gFJVG9dsjb+oeigo18OlW
QhI034fcBWaHMfJfpDOUnm44bWOoB0s0xthoZaxHvigpDI67TglS18GP0Y065zV32oynpUoWkwNm
UDD6qksJauvwyRmED54yYUFINbvAPic4bfIPpisfakC467BcO7CZZkaJiw1JUPLQM6rQFWndNC1g
okiF4iwhlQNEmF3QHzj+0hSSFYzM6jwZdOzxJKNbQ3C5JpweGXdK+OWnVTDRq7kVKZmmkcDysWR9
0+/sneMFs6WQWIhu0g6XNkWWF5zQuZrf+zAMtMHu5kT8WsTVRkYnga13yjFBYLblnDNr0Im523pg
9xJuXQu7oRaE+eOpF81I2petJuWMIx2W3B6LuMkID2VP5PBDLLb2qdB2p118VYdiyU7hx48oengz
KX2BTCU74yMMGv4BEti+Gw4tl4QaFPV1F3jLuVWmVxrSqK1M1WGss31N0jsU12bgPE5Iy1K2/M8I
zrZGvdXVhcfPF3XIhpcI04HI4nsEGFisuK5Fk6K4tIadiej9P/L2BwZU6yILR9nRtbhxii2N4lAn
AC45tpg1BiijVJqOA1x1t8UESCTIEumx3j3i2sqOiw2DyBbw9KkmqDq9vVfWBszSqftC29/DMh8U
ZK1GH6vf6R07nRapOLPv0nFSoK77x/2NWI9xgOL8r2FUtKdSF55TEjeulxtgUzEbLdEStaTnJUQT
zB4hvsb8ieJDwLC0CqcKyRMOEW9ZJnV1nyO578atSyx0yLH5T3lbQgv2bSrbxzEeFH4HqtkCQUeS
k7oainDYx7IKvPOEW+sn+OrEmtokMTPqXSG2pXb3XZ0HDGf9os/+65DLfLq6QoYJT00kaCKVoPbG
sGiFS7LChsRrpQz+i/sBWRubW2QX7zhgQD3ARf2X0RlOtsbNEdFwQY0HyKVP/PPDI638rfP8tupf
Ttw1FLwtFfpi+hz50Pjuzh00PI3Mpui7+6zJOcRgVKkwsU5FOGa86S+mI+0WD8Y1cZsp30e1yeE2
P+McPWp1qft03cSOXfZYXh7C9os9BwKBlV3uWO8FRPJ8zrhcmjR/4MN2LHMbcuqp9j260Nt+beTM
zvRtLodMMIi1w607X6uQpy15xaHydsrtt9OA9H5Yo566AqjbMhr9FmsxXQJy6gmlvfppY1sZ9/mJ
+P0Ud9m3iW8stHPqVTUT0QDDstxknZ0TmYz7T4vA1I1USdHkO1iW/NfZmGK0v0HwigIG68irgtVP
Dn8c6EpxgYjwnq09zrT0j8ZGQOTfjYqG5Pnb1koS/YZLn2LlGpTZxEEp5pUCx++32Mfw6935EOzB
b4Xj6bdGpcRYaBl3EJ3/lL3oQj+mCDPj90ek1kiSC6UXJQt4El5wqKt220zKE5tuCo+iRhmnPU0d
PdfeUVKwrGaEgQpbZOGBcdBgKXMT3AdOkj5jBf/F8jfuw3cjcHGuaxYz4DZRVF0oEKNRXMyGoYEN
hctimTO3lCD0zmRsKl8tYCFlJGMUPvYPam7wFLkRWVCOCKcleeofBS745pLbKRmwTMEdsBdSOx9h
KJQSkzhRL6pgrt0JnYcuB9+XpwrWRl1PUNfWaLPHfaeLGF2Z8+7thd7cL5h26UdC1Qg1XDGPSG46
oLfxQ0Vsi1YDQ2wyxj/YFzPfLL03uvYBeEyBGmBtPwjqcJIY8rhpFr0FMUgp6XvpZpGD+kgDwtnS
Et+RF38jB6Z1Z7kqK+cK1J9Rvxotsp3dzl3Rsju6CgC5tgPMeoGtoo8QYPta1olCZP8A0o7Y/Tza
x2PDVuK4Ca89wBMGHDtIRz8arEfbsEUVN5YaISFKDl4xtqq3L/3mEOfIWsn/hKs/UnGrKPHOYUeZ
e/jckvBi9FMwh6BezzwohX7AnsbQYo4uBbiryxQmFD2W5DhMbq1xzVDPpgUmAJnqeI5a+2Er0oSh
evls5H0HD32GzsAotM+v0u4+B+0lRdC6hjwhwBAeT9v0hGxKXXqRabtSyR3ISA+B7/soB1Fmsl+9
fxXvPbrN0YgtLTiUzmLDmYm24ghnBDEBfQF2xvuqixZ7cxAYVx8Tnnw3YBODmExxWKZ1akMViyGJ
DYswibkt3jWS44kOojTnPJep6wiFfLqkWw095wM2UuFUQdzjtejd3cGQHxBNO8ljeXUxaawz//z1
2YTsnvYSAa99dg6wWq+VIfH6Xq0VPcA6oxmy2ShNiOancyBseNucvEF2+XW+PPAOjfJfY/mcz+LZ
5TQ0pjTmIOkIkRrp+z/R9LgGBVXsvSta2qhFdm2B7MFN+Tn2RryTwn+9gZRntOF4Pu/Oaw+75hfp
0U/aaz2jDI8SPi3AGIfZClTcymJdSUKMqcs+7g71ef8dTApRf9BQEHmQiSNDrAn3zjuyK8nJqcuR
wJLzy/7AlkE/ZOnH3VZdHygLytQ5ISXCnyCVdnpS/BnNQW4kqMFbPI/Tqjff7tz/jHsirFm7CWfa
QsxPHdEQjbSMa51ud1CfvjgghkJUxFJa2iZx+lUGweVkK0m4+rH8SsaKYXaN8zK8U/hp5yJuL6w4
N6WgeUu7XgWLymhQnUSwC4iC0eEz2PVhXGkLyo8d7bHW0okIYok05antwGZcZNKyvvv2lXEnRYQn
jGfMxV66c7vKp1BcF8X+Bjxt9N8Jn3XExuyLCwK0XitWwb26XXl/WClvftedZL/udQ8RsA41RRK3
MralDqjTqnAduH9Kwg8jWFi37hZzTx5lzCo+Z2dQLseayvX2OFsR4FZQjiiOxva/BApz2FsPM9Cd
s81wghhtuoP92iXcsFvbrm/iYq75c68RFH3mBgMt5VEn2hSLFdUz7MlzEh9pE5lGENDzR00J7qiB
yTyQB+01hWZ5fUhKbvutYqhTTTV4AswLbA0Vd8rvdvNgfdkW4oDgPTaMvnlSl7X2nX89tYRQldV4
Da1MXkgyRyGGVlWPBhymB3hWUkgPFDPc391efBDzkrrjvIqQrw+RTP1V1KohVCpzMcLOhFysXxJk
GrNNmm3BpIWOSHK6pbg5pT0BWu89n4eS6JxhEHtg3ZNG7LyYry1c90+LloXcIGEdRUjYVqFDfjwk
gDtiomYzv1GGnKZY3+lBnMyIX0OM9eSM6G2fwWLxbkaeqMCeBZgd0XWZ2jpd5m4r0Iuqlqr1MN9N
lFhD6a+tdzTFHTtVapN/xyqBOZi4dAFBT/yxQL6znNR5Bqdt6dyks1nfMVnu2fgQxwBs8yAySGhJ
0+Rdtd5V3zddCYrknRyQnSJLEEXPdoitgUu9QOwkW6URlXam5gRY/m8O5Y2fFwI+IrahPCZ8vq2O
dTuqskvJPvgUn/x9/ZRagYycUvKuqFEv0YTjf+cE66aMl/SAbt4EkM973ReRdLu7BJUvIjhQTtjN
WneTx8xQ3UwCVzb6LEunUDQQaMqcPaWMkpd0H6sOOZqTyfCT7LdpMVOdjb89+Y2sPmarcW+D1zi/
OxewBqH1I1UVVKfOAQG1DtxHD+NtMUi++zl4R+aRbEyRrtIDkyS8IhoeDjCHpgCKEzwrgJTAITp/
KoB0XhWM8VJfE9ANbXzRYWE9aG7uUN58fa1YY/ixmsqAlQIZrFPtr7KaWZHgkoPNhs8RUIO/ZuYE
+TuhjKiL7F/H/MGB0nu1XwD5jnRcOFTKpiCxGn+8ljlR3j3AICG4YgnnjNPdJoXhJyWCFcsmneA5
R0ucVJIEaZLBGry4FGVSbKAOYaXx9nJf6ra8W3pO4ou4j09ia3M/ZrTqfPGu9KuYkOnES5g2rn5q
fVzw6UvMMNTt4p2JRYmVka0xjqS/qomE0AC6r6UyWjdzbXqrvaC/EGM6SjDpBLT66TERISNuleUC
btB1KFv1sh16tktEdF5bLyaa9gzT3mMxDFHCEHqrJUAL4oFbT8a6ENHLL4l9gpvMR75JpZ8osXxb
u7zouuu3nl1WCjAGsz1NV+K0upbxUYyHw8JVm9yf73ng0N2lJc445yvXCbg3XdoTujeLrwXvcIO+
8gRZHmUrqlITmnelTY4HNIFaNM0tfzu70ZThO2W0VjEeFW2IoFvbj2q6AV6E0QsAG3LuITLyzsgR
ViW+xlZWdDuf24AWHmWvvI/zan5DeAtcIhCpHU5gDu9NUY0mAeSTm5kKpJUdvpBbZOCOGOLd/Bq2
I14r/f35RGeRogjcStu1RTtbTcPVwx6mgGMUWPfqDTEYT391yIfC4GMT/jua/a59v2Wi5DHTVz5G
8yOLYY/zUCAvOLDt9srbMkYFsNQs1ZHyHoo91YrmFtf+6vZcVeMKl9AJm19Z6eo+AeLvNLRu9f4E
Q/0UgFtYa94pjyYpPY04rvQy8m8/JWqIaGZBMfXdRGPWh4aTrNdw5VLvxRQ8ONx+SXDD30a7qsOq
FXpqIhTrdgNVNxCwIz83wxcGj1i6GrakuySkCbCtRpvPyCM9Dkw6j8lJEvzldWJwOzLIkB/zXoSA
CjnNFH5pXdvGUMyQGoZ5vApwOrRnOW499yhGnz5MekUoZ5SeTlSxdo41ndKYGsVW9LDu1d+cZcaf
ghzqD/ch1L+Ilb8BjAv9ib5KgU4tMvA8deV6k91hWYujnvT/ns0oeQOGMDS7G5VbkS3DQ0nBw1ZH
cTQO2rHqcFw30huFCqkeQFLaj6lLJBdVuTxDFFZ9DKqj8u6BcqFYThepQJd5uXkvLQAFj5f2cftB
K58e91f4XSzhFfLMZMyP+rvj+dVvvEWLf5JnVkCf9WobeHcxl7yvkh9h2Pq1an7E4f2n1BR9IrmP
bV9COEKwQklywAyWTLGcOXnDZOHmP/1mRmxoAzZzvVY5p10lOGBArZgo132fmwVYsb9W14PRcUlT
EYzc2tzvW7YxunL3G7MabtFDfJe65Pqzgm/34MvPEARPf2s5XYKwCjF/tFkiaKorg5xYhwJqA0Yr
Cjhooi+Br60hht/Ih8FsjIxuMuz1JTW2Tqv2sDOFEBPbOYVo6d0D7yOeSjtk/aQ2D41Rdp1DWHhY
UNWRK9BAFOYoN8VirXk3jHXDI6pzbMf0POMEjx+sPko6RGsg3yWL2ZdIQkuPPQNcVZ3iaKDvJBFC
bAjCDE/c4y7DzPPrg5ibb35Pf7TFCElIwSrJRGkMnxlkxhLStnC3LL8/viPpDYM1NAVBt8FRyqYK
C6hUPEnyL6Irh7lv8Uxo1BG7ThjIQtWeNxD+l1SoJD5sBKwOaIcbpamV2USWci9kX7lKjwP98ixm
Eh9yhwsLG5Si/1HTyoytWOaPO/0KTHIH9U/8AlteX+fcd7S1UssorQIwlcv2Rq+CCfZY38Ilsb75
NWKFc+MrKzbaXSXJ0R+uSn7F/lWxksrOfw0JPTITXlxxcKxHcUHmuGUAOP1q3PhtN/oilBllTLMX
1IgZxJXoZzZgpzdFHN14h35fcb4J1/CJcYwzHnyec2ts4JO7/AMHcc7n2KBKRMZ+hxc2eMlw+saC
l7bcBnLoqLADLCYCLiXlmsEdBEz+imitYdEQXRPnnjotYMTStKwBLq3OhFm10lZ2WsH/8nARfU4G
TirDpdoAf/AfBdWFBwnutoawqtH/ZuhYqAZRoduPI5Sf5St5s7i0yhVbVUO1kN7xM389AT0n6kuB
SQHB9K8ZtYxf5YTjSH+8LuNqlkOFodXAjf2MjHPoHNUW1ymCsufD9uSif0gQlEtq30/unrXdqpGb
Rl4KJfRsPY7q5hDGOZhHrrN9PhF93MFyew3eE+pK4W1mbdtVZtUeTGEOFRvAxcDvdQ0wxqn+qVhn
0HScB2e852D1xyeEx5SMq+xhdi+QCITsAWreS6CggIrvBkkTFJQ9kOkLFkli2ef02zhpFGRh3pqs
2v3Jur/1Xc21yKCHznw7YCEp4JExqN8qWL6+cYdTy2B7czOL7AERZjN5WHzc6vNz99PGlVPU4KK4
0kVat/BhSPA2kjEO8zwGGxSY8ioEegc/GcWaiWplbr3WEItdqbOagGpxvh351jwEkeJviouX37wc
Zzk9UhthcwMbAt/3iOM/xkRiyDBOPkv8UjCVwQiLHJemOIIT4z+L+YzFrjmEbpdinXhGB8yhOYgf
G2OrJ37TcqbwkZgbTOh6jDa7rqiOuDaweWtLgCv6tSo56zeW5Js5X0qKtwCqt6J0+88nxSjlY5TV
YMkqB4OJYxl463qkTqin7gtlbegNPO6lC+IazbwVyvnUW3IBMCo4skk1me66L5DQxcpxwnCa4esU
19SqQruy9BGeSN/WeqIbhRbD+bUXtZ6OIyixM9OIZr+aNCjQ/THPKIuaTd1k2pHrB+wLJGOoHU9Z
+60aYD4Awq1eTEhVedbnZOOq00Mnn0ODnSzhTbdZ7WBwhll9EoTfkp4hYreFkA05eWPsIv3dDmQr
eK06IWJhYIJ//JXLOGlZNTE9C6zrEYlb+pvLXz5C8BVY/Ev6P9lvenzn0xGBirLn0F9IB2bd7KCG
WEB5LJquUKMuqRSYDKaOTtHSnjj0FFh/nF//AOpvuBTY09DzlYh6ARyLt6oVlcgWo8wD0/OBRl2H
mUqMY8UMd76kbMgHDIAq6/1jd07Vm+2Dzm1RpdQZl/Ri0HIo+ocyOE0UrOouvhuzG0GULUpN2E0F
j65IDM7NpcLuVyEIb0RAbvTwYN4csjELwsq6a34QFastxN5XebiZftwoAke4fwIdoiVhg2UI87xF
alWNzKApammnk0T5jjBfnu2d0f7mjHssvb7+uL03y6eCKR7ZXhz+4T3Waz69YzVbkTykItoo4ds4
TKkKraCpqmYse+9xZp383dJdlLwxEZA4JG7QKTefiTr7spX9F/Q348+xLV5feEPli5SZgJw+zF6Q
GomtBkuuxFdsKZ3eM+UYN5v1OX9u56l9PkM0LGg7TaDy/aiUD5N+NWNY+2OCIMVAWaXsdIqyvvwK
/5RfHrn8HY+yxiT+Ym0V3IihRIXNMMGPTf8nPPVEoB2u4/OxZtQMwPxMxRwiS7NU7wO0Kzvwb9bL
XkuZVZr9V8lWxcOcHtljXUnrarD3fDx3OU9N7ZcwMEtzqC6IgYK5JDwcWfHClOLaFobV4asRLdQt
lmp07eEEdZVwvWmkfjaxyLtm9Vj/Yl8kJcANQiTIU7VuIYuTHtdREWmlENVDBSXROLlE+XdHBfgx
PCt8ocYE212157UAqUAaOdPgnHMCWRC1qtIqtCiTqHKt7P2ZAKKlq+S1NlHTqCdgculPmQYtf82I
IXU2mVR8HrBAg/pQjI4UjJpYRVeRgJkYjsSf6d+SoWWDwZEYCO1tLKNAj3vF+7Lz4ugQnTuSrAQ3
YGIYNi5dsUoVOlmSkB66VWfHxVmMVvazV8xqQ3lFGspSYoQdyVkSd48mJGOjpiLz5magrY+Gc7MO
Gb9gIojHnSz/wwRrUE7qCod1aihG635smee5L/sDU+6fjRTR4USYJySIiEPrY48iDjt9KnNQw9kW
t4JqAS9b1TY8NUioM0ryZJXY3uFRj6LLT5WCuvzF1vDLLmtNvNOA63BvQ4Ad8oBsWL+sa79mT0pK
E+kg6k8vUB528wJcCW6A3Q8jfGthJtrlDRaq/xwDZsWPieIvBVc7Q94qi0HGNbC7Kk6e5zvhhKS9
ajzSwfCDbEq28OnKhMsQdH/wCNkF0J3vyeDS4xOI1nDLwN+PMQkugTwDWwxyVDSZX8YySC6y2Xml
BUbn8QBduHToCtd6naK2TKgE+Kq54mKdhMbp9HxyLzn7JcueC8vpb9Ge3gWtpW9w1NZ7fKR/O86b
Sd6Fs37QI9wzGCEDm2r1f5XWX+JFbGsj93IT9PMCodA16kREs7KAz5nPEb6FzDnBs09hl6Fpmy2n
gxWGeSCYFAKSiSn7BFM4j4ug7dxike3VtcwfjBeH5iAt/BgvDDTAxLsfYONJiO/+CwR8MOgYWJ5B
QAbVMfj6UXKR5zY5OHIWoNO8VWVJ04MZV5AlrSKPTg3hsKS8ORArUd1JUycbC/to6YcRy2WXQAuQ
1v1ARLJ7UBZQNf/KXOlWzc97m1Lg4/zoUehXZw9xrNN1uYuAbISA/RMCynYuvpDJlRW8x4ze3mbM
o4qI+5dQw7UpaqSqY1/of2PaZP3hqpYDMQWbcMJRhxA3Ae/uV3yKHzpl+k19COmIpuz5DUjAhuI5
rsJNCL2jFiULH24apojurG7LGuPRTi2oc31BLhVmzdT5N604kwN0dypGiQjnnwkfnYzCGStLKpgY
7l0PsAl6yMPl1qDlfsyFG24cT+7wdo17JqYco9cc2eoMdQqMMEjmhebD99O4avHSO/qcSuopcS2x
7HWJ1XpFJBShkRAoXB6drllyKsuxIdB4YB0EQiwaGZHUCLL/oWELQO6jHV3MHzxiVp6wxsOrlJHR
8mS+Drn2zpMT8FWd/L/iflaethaMsS3kvQsIwHAdMXv75lBIKZrrWd6QsO45QfFzrD5RObRhKMK8
kdCIKiHNVyu0+RREZtgw2f4BqLrwFCH4UYDICsBYD9AMhHMODSGCDon5VEr088tI8GIhdA0sTNyf
yqC8NfypDWdPVXiYNckSI2ApuesJPw/t26dgw7GTx8bsHrrjneqg75Gr0kE0DZoZhHhZGC8TOZFj
rJVjV6j6pgwaXL4hw3IccfGaydB56PBktiiVtrukIuwxOJbd95+P7i2zHMruSAb0Tlxty47APj3T
YCw/k/ZVTQLEVyDqrUN4MHi6j37hX5MPd3Ow9Cla/KhxsSeKfJ7TC4G86+FfrgkM5g4ZXUNZVeDp
AJCpYgIAe6dO3GMXrZ9aurcjJsydJb5wVUZ2PNPcKWWsvCQmMOmjuc2HT8nioKwJpnrOaPODB3i8
gQ56WYfV+z6OtYZcJWxWbToHoC5SJq/RwmC+RPs0LdvDy4gmBOGTadCJbVUbKntea6P+/RKqv0kA
h2EZzsOO+PqE1wC3YR+LkYGuH0vJ3odwgYkhMP+CLpFDE00jzCGOkTuQGx9ZZSiicPiS3e1X017y
9gFoP86XRG7vusdAl+N9ti6rbd7VwWaQmas7KNA0Yumrq23pdFvkTZS+xfd5wZwOduryauf33lAi
MUCwGpcQ4hCFDDsYkbAVA/B7qyOsYz69hgRgi7rIaOirZPdnllYCP0gv5QaxKD5ce3aqyEioed5b
yJzSiN5tmQI/StnAB7LJ11Od3fIIyBvPBUKon800u+U3LTTsIRqfCugS+BISv5dqvBZxJQm2DViE
XmIZR6xIABk6rpkDVKqgA9JpWffCnoWroKSDFyHZZvq+FBESImzMCkbcSD/FYhkBdOzfZib1Wt9f
zRtFlJ++64jJ7oC9sje0IUmD7qVxN5gnnQUma+FvjMnl4KgcJdessfqF5LQeQdbBocXyARM1XYcU
Z0ck6xeLrl8KAelB1hYFTCKAtU1pQnhecfVFdLyeTty7Qb7ukf7dih6izSjOkKLb/jN20P1vTxxe
YMIl862YMqnFrwG4liKgEdNq+Xh0c5HcUrGW/kDRJV6iyr7i0ljvdWRgfIIhRyR4/6y3hw9H5lrA
kOb3Ir2/xp7anoK93AngkRs4OaD0Jy+N0bItwVviFHXVhhUhTJ+Ko4bBe6SyeCFyu/38qpUxUkT3
90WetL48p4u5pcdq1hwsxID6kiXsZwGWdwPbsrmub48v6G3qaAeWXiGfeAxV2J0sRoCY4e2i9x0p
15OlI/T6VEcq2fow9IDH1l5E4mLtIHfx54AcUf7cSvwIpZdUQy7fPhwZ7jJGb9xov0VIXe+GzqbO
RKv2i7JlnZQn4FRBsu7fGGN/hOZtz62tUezxHqSws73Ow8v1+udZMG0iP7lmu29iLzPGhRekPF6d
EKCNP//bRzlef+MGHptCkNowtSjobLQT6m4Xe5d0rGkVSCYiJoNXFEsZi08clmVemHqvizCWHJ3O
WlocrDMlQ2hKf6lo/s1zaw6ehsoT4KHEyQwwS3flCHEXKfUuDM82PCMFeyuUCa3MfDOtN6rOaCE2
hy2LOW213mGO7SQiLp7mA2PEhCgrn0JUVWXs3FIrdnJ0gKSS5W4w77UMJqn3ierTwg0lMLf0Ekll
AKgitF7iXRmueBnD2j1WC96bm+F5OvQ8T4HhUibGQhJyHkEi5IYs9UUqXFFdFeuR9jQj0DLqj/6Z
9SjCQnKVYpPt82rUiMYncB0I/uQRrD615M+ylD5w8jJ9yqdqjFqJtjNBzoSvedrWGe+1GXu2QMRl
khSuYCwKRjs662oegnc+uwcWpZEURmrt+wtbKiuHRHljf5AAL8QX8KQ3W+MsoK/C/8yYYEEZ4IBL
u0Huf8sqQFOijLNiLy7Exu1LiX3I7/faBxrx0XlN0pDVSZq25CedjTC1KiF2G2GM9dF5CLqP810Z
whueR+cwkU2Gu5azyloPPb5ak0HipeHll4fjNevvG2YKHbJV8ncDTgi/T6h7K1jQDKHe81KxTMSA
htW3QSKOvlh2//YtQ+znAa8PNOs4wEtn4MSphKRpD9i11u3vxGWbKyieD9O4fVy6Cc3cx1dIRgbl
WRfwpkgQkQ3NCF8c9ZlI5rp4OmepmpAhbNehr9lp8zTpOX8adTIIcxTTTBGUMWVVIUcndjv8dvXw
J8lNJ979fIrAmyYbrXsSgsLGxk8f8GQ6P25ktHbCOMO1qJdHqcFVzw4V1ZEmhDWtlBVXvH6HwKEl
rh2PX7IPfemanE74XFBHxWY0WOZOuqjJg31HyQg2ztmobHRH0/rMxv9AIofMOwOP2SOGOqtprv9j
koZcpbmbZ4SQX+IjkxP4kj94hvdl+TCLb4k8PU7AWhWAjWsJvss6Ci8CMaqP3m3galC0Ef1LEAdH
A60/6hcHRR0PmSEbEPyK0CMMrky5Fv7BaewtMjwlvylivyqPDX2RnOa4M7n0fQWB/Z11/UxuFJhD
N0X+akfoK17+8xiMOuohfrs01ge39uKM8zLqRLk0kDa6oRBzTEXvj/PPQSDpvSXjxF7olXb5P5E1
y4GWGke79wIc0J9769EG+a2Z2yXiBnWiNaGoDSe7YhPVH5/mL+tgj7Cgn/jNTS7rtNUJzy1PXgaf
BaiJ6Uf98XaGMt8QiyHkiNX2YCuZU/q0js3l3x3l19DOJa9eOajVtCO/FONGdrsaW0OwmKMLFJQ6
fkWUDwoaB/AdewAHK36ZLSKqDOfAZoMy7HNWFPJkHWouMQFbUew+Sc/afg1B3aDMfiwS/QIQYcJE
U3+qT87A0kt6hl05iZFCodUo9yfLK2cVYY9CbNsryDFeulFVhr6ZxqHBVaimcO+9Qx609uOvBYZW
WU09tzlb6SFXIcXxT7XgqQswYbhKpYAuXgeZJZVeyw+Sp1laBbEZ6tFI0kU/w5+9HH3mLrtrN3Sw
0Gr0wNfjSqy5VFEOMI5Ftyqe44URNNlt7I7ZoDGj54fjdgVrslZCfdVo3l3UDx24XJmoA16pkQcM
TGI4bxlfP155PzsB/C8siu8zPltvx0AgEzfsvZdoAX+KMBKhJbFst2mtiK7nLyPPLwK7F7Y4t4ct
mVfXPYVmv4Fpe12hSIFhFK9ve5TLw8GQlpMbXkSekMF336h1czcCEnaDWuGer5tCyHbBpV7U4kTg
QiXnJIrdPVbBTfSluo5VSBom37bKJKQcR+J5KiouYZWZ1mfQx6hkSW1g3gbvl98p7SLJwV0vlrcm
famgunLoHwhs7TQrKS1h9LfL52VLFScsipJ8GoS1pMlzxHBY8IxBGuhf+HFTbL9YIh1Qp1XDUmDm
OsjdrWg7RoSQJgRXAs8LX2+osqOK/tzGu1iHjuHDJunE/BjFXA4AVdeUsm9lp8HYW+G/ZLIfbAKD
OvDmXSMBUlhRMC4J6CKx7dm4x5r6T0rdoZprQw5GJh8nGxWV/d6bfL6AVZa1RlpKRINXx9K6KuLO
QNc8WFnPiGBf6WR9zKQZPa9M+jyeVSqsNeKPM1oL4uBJieU99G17ID0ancY3sceyF0CYc4pkU62/
ihjiybdU/W+NjNi6BOKlUydJxJcT43SDMTKOLiM2HeYgG1tkNAi3x2vuF2tIwok+yz1QrfvvqQxl
r7gkNeBe5OUWAfDf4Q9NQ183LagemIiscyheJkh77RJJ1kuiwKbUfaH8TP16XcsS/ElUX1JM02+p
l8IG0960q95eRmWHTPDZwUel9/jp8rdjbSnGiiNFrLW4w6NNBAKvKWKZUj6A9hhgH0sy/GysiFrT
arF618g+0qvww0Y9MX1u417bjJMGE1Kn/s2XGd1w7MlPiguk63TaZV4tSA7L/H48HXSVpdfYTN3z
o3awZzSRpZw1JUqs2DceviEMb+FKcKqVe5sSrsdmYoVEgKJcSenTA4QEZSdEVPZb7497Ea7KkHia
hVhrSiIQiqKF5bNRFbQ5PuyYkXzvsipo7qMstc0pVaPZL1nvo/II1SZ5zuNLuKPam9NXt7lwHOu4
0FFU7BcUz8ky7Wvd9fC8U4Fejwi7dK38o2TOY4mQcM1aC/drVb1xlWcY3ccNR91QphSyBvvWNH5R
F8VhY3ZizPvSi0AchUC4uIt2uqq/G1Z1mdwKaLz6eGQJ9W3883SfZP8b/lqc/8DFl7FiACDomkBL
3DOvNoqCBiuFX2ih4OyPdxFc6ss5Jk3JKsd+PxUwT24WCDhMt2swkji8q3NYbMcnMliGNN4STh49
Iyh4uzP9z1aKSQ6NLltPKPHpxi08jGGHjaDZTqAfenH32kiXsX9Cp/c76wDpJyq+qhJsNLMv3hbr
8fZcHYHTW1TMPZA9L2Uy6xNM7ov17ARu5hjALBDxS6yqoisPrIdVKidlPvCJKz0a9mjtf3fDd8Jk
aLYJvdni2NR8lOplxjLrDwE1wq/JiugdWa6dF8aVheSSharOO/cb/llPZufmj21wcxRG0QKyillC
SPbRzXJshNY/mrIqZhB+I7jjqh4c9zrZunUm2V9mWFu1I9jFRYDy/JjO+/nyIBV7VqHAOHrcFiQ7
2soCHnrVn827S8CLO86LsIgpxTd77hmtqLv5kSHeDCP304vtsC9RZn3N6341S7co7hcqEZ09plPA
VD3L6XVT01+cDn+b6LFSmFYQ55CO/8ekl11NUBTRGjV2eqmbWQFXCxDl+63tQYF1JKt1dxP9w42U
fvQ7fUoo2x/KpDyzM7Pu0O+70+yRXcLOqTBev/OchD3FR4hPd5nob8FAyVYdJj40QH2S6ERVkOQK
lvYTXfdsDklZ/mF8/yMeCkjj6ZTs/VbY907r0R3+Px/YipWZ0X0z3WpdPpuz4xDk8R9C3FctJeef
prWThdmZhTW83pHt0iF5qDVVC4aWDwQt2tl0rBTC/6pb1DFlW5zM/APbyo1AKjZw8CQLW25XuUVx
PPyuGN5ImRUJwD7Er78iWNevdBktvE4Pq2ORvJCHtneZQejwaDnIG4uP+WjjL4dIAzlgMqsZbc8B
tfGA3tXQomR1MH+CgTOZ3vcMO0IVVC7ysZk6R2kcZr2XwF4EAA1xuzcB13wx/D2gCMIpH1NuZbt2
a8Oi8koLxtrpVlrEwWbE1oKBgE+bBVlEnZ5hKR6SbdOFyXJseEvUPAgt5SY8feqlyajjwgW1fpzb
n42+ODqLn+LbMnkhP1F2l7t0L3LQo9TFsbxefyf4pfXQj+chpu+BvYaZqYhPhizpCZ/T56inkmJj
Hi+s95IaHCHU6oSh0mdPw3HxqrbtHPuIiqLqWSZRZMivBhH9KgiPrPAmKGG83u/wXoW8sUCChYPn
V7bH/BsIY26tw7iAi6xnOUTb1mwEqYrvfnIxcwoIFwKKsuUyhoshGssT+azD88tPcK0yQZ0RbgcM
0P8Rq32/g0CRxN3pjRx0wpnsvnRlTXIK4UUA6ZKjcuVwfoqJ9VrJILxXceDgeYPYlp4FrgfwE5S3
L4u/xCuKKbnY8ywJFFnsFkul1nHr8HsGroJtSCD4zlomCUkp8hIRO6X7Y9n5CorNa17rCIe1cgwj
7+dIxTUMKm/RkMIDn6EO4m5JVTU26M8PES5DC2HJY7oZ9PlChNzcnQTtVfxmbf7JQRcQfFxqthso
t+jHhOhXUeu+XVoXLqSRmgr+ICUKywXsRlzlZAuYWWl1NEYBEOsPgyatr9ioq8ATuf3wF2uxlHaC
Mxf3lHw+X2e+k6nZW26z8Otw0w9MJrosVxitiEC+i91jTOwn8/FjQVZ2fNgTnTwmxjg+AxV6NXh1
PjGVgyTN8OiNXNk1Xds4eVxQYCyJCSnl8v60a7UpotX8fVi73FzjwjrvvltokxpsgFHb5qrFhMmz
enqhn/v1pxozepVGHaPUh3PDVbfZnWL9BPWyZaeF9YkYURG77jF+/DZYagX5EKYgz9H0dbL+E8Qb
LQOqhJ23W59i4JXV9DTlimhpk3UiiMtkuqZ0qYwZkLXbMMUwqAo+Nq4I1tevA9xO5kL9QQQdP7MI
jvYcLFK6sUc/YgSl5REiMcMRcuoVaJZdDmpBRKujp5UUV4bRJHLrmE7rSLj1MAzBb3zg5+RmF4Dx
QZTZQEtZjFl3AI0UEP/f+Y2loLOfkBJYelu1g32HshjeJBnyBLNEG28OO41VuxfY8K4BdEDjFFqe
MTz0IFmxAOYgAKce9MYT2Z5HTStTVhSMUg5w2j2Sc/IOGXFBim7bP/hz06cfOXGU3CC/qq3dCI+U
BLnDJINwN6hcQ16qwkZyd7JmU4tzMSNlhnxvIp58edFkbeL0eAyS5PsELUu3Uc8ZpnN+rgfjhWlZ
bM9aGidgvWatD80cqNSOwfe1VLQP5F1iUhJK40FPCj9QTAMPS1G84el9/gV01fi9dUl/9SlmCN7I
1a4+fayUgcO4nAVBaE+B4+jO0zGSZoGP2D3XNnN5quw+vx3/aExuZh0PF/iaERBA4tK07FVsijOV
TGzV6O8gUEAdxFnphHUEdmLVI4yQ8GN7R54rDumqwtU/n/0QGdhorW9OpRenp4oGnPRaBrg0EvEi
qZE5/POvg5UyLS0h1Hk8bZNPNxIWSN5iGZjx0jGrVLkjAeiiZVmPxu0liKvt+/kp/bEZxgty5ZcH
ExkQP7esr1HEXBgVV83SpZ/oJKT5W/mm4ebyJO573TTUloOXzZ1SM3iAOtrFEa8gvIx9CWdzVtOd
wI+pBSQ8QqHUpi+DdS7uEZQ0E7HMQYTJppRDeX05Tc4eDN5AgZYvmb+b3Rsd+JaSDkVHOvhBqbCS
6rb+nnr+FiTvVT1X8r2ZfEuKrcomkt5VQfbHDmM/kal75uRFJFId56WjOTCWdSru0FGeRC62qc+t
L3J28LXmDytEav2dPN+1d2WTecs6Uscr1WsiMvkbrcpuOdckT6N7kq3oc1ngikS9Co2gxuLvX6VI
nQddZ/HMJFtxIgQek2kQ2vHgx/vQ1ikLvSAZiFK1HSd+3ktbJQ+DLrwtcXwn+DTGAGOQO3kkh0K6
a2PH1Rokp8J6ZBx7yNh7V+fj2mLWk0jrYoT9j/1ZZNgWZxE2iTmviycXvs0DhnM+vqN9FdmX/vrv
5m7vEIrZ7VS7Ej7ocd9LKSyAdeqavkxnLM/uXrb6mwXzcX3iPvWZI6D5J1/ytlYFolQIMDuXQCDw
1dvYKB1K9wSoRRDN/HFcpiw64a7uUw/auj6tvRSqbrfpIK5pcjsLLyG8Ec7SWbPs/gjUNAcrCCgC
byQUDx3OK/TEiD9SJbeegW2i6g75yR0s417gd4kI3tr4JfmmMyAATXyl13K3XFLcjfvdH+Q5yUYo
+MB9hP3BwxTAMiVq7i2iR1Qn8V/64oJrCZ7xkSbG0jkONO5oewQnaWhl1miGdSVtnxplLYii9gAH
mWuS080RueYsx3YtvIv+h8EhCADmGKXAotKGuRFnRs45gQmPhm7vUUvLiEjwBg5Q8Fupx1NJll9W
k/NGyV4bhebbQ+LsKEYQrvsJ3rVJABKVavUVdu92kAZVL72l84WXoXdwj9KRPf+KA5VbpSHNM8BE
aIPCf+YqfMgb9bK4HCAYz/MGbfUtnPELkMz2Yrny4jJwT3ZMlT8t1FBrbig5w+19394hFnD9AtEU
NUTdfr2gD/Q6rjw8+EeU+1vbdR2WWrgmD2aE3r4V7Vi+tpgIB/sY4KUavuEwCrFX8Mr8fZiyPi3Z
xDPfpivpQqY6hZPtWIvvQcdXa92w4+fdkpIa0LZ1quNZxzpPXwmgZ7Ak79UKUjCe8liDe1WTgD1P
EQ/hMgXq1KB0F44q2+Mfg6ZWrPDWkZPtLIqrReFYvG2+8pTQxcBVj+NyQ5EwDiyl5w9DSlAhJ26n
ZygkWE3qeMz1DZzu2HKp0cts4TXxwb5USDHnAf/klrJ6Wz5keclagwQeRAcpWp0493kPAInxnm2G
3/sHpcam6a23P0yfI4trgrCtDdQhLIbKLMspeYfOvpDCJ/OXrUSrKLtShnXZhUVxfuCCYk2gSdOZ
KA+ZEdv8oevso01Kqoi/UIr5HheFDs7JK/GN0frAtZonP06VmBpXtCknH1w1EGzAQcq4bwBkH8y5
fEwQADIrfS96YtBWjgz9UeBnWVE2HdBlFSdND9zoTvKjjVDHKR8JqXWA77mvfFvr/G6zFVtSngMv
ZBGhPpRegCMgjtDpJi1a7vqqGCYhSkahqEglK+LWI2pWjoUncij0DD3mp6f6zm86td/rlg0F65Hq
SXnvDhitAIadnqGp/CBfAeShbfbwjsOPJzPzJ3FzVYooVeYZoa3cKr0t2IXjg8mm8roVGXZrTXRY
8G1WRHBkPz1vmh2dPQ6iG91mu70WrBfgdDXkBBv9Dr5bzNwe1zzIDlnEQh9+RuTuHvySwTElxg6P
CrHlrFGef/bbNiFPfIqNrM0u+m1tSVUMJG6sGNubv3v/GoZBHCoAUAIDs8f2GXWgTb8T5cE7PVbP
/hLxMGvPbhjkd/yTlcp6LwBRFO79Xijf8C461PgXYb4BW4iTwWscceU9BwPk2fT4AWDsGob8tCCU
7V8GnGbvu4IA1mmuqyodT0imEkDbMTSnwCBXyN1E5DKExoSFa+R4DfQs7P0ydf2DkOiWuiFDlcyT
uQ2HaOJP332NwTFTQ4NAc879FVRgheYfdI9eD3nmhpvUHUvuDVKBNm5gXvcBvIo9lA5eGnK9P4+J
/KhTxW8so4HO/8sipXSX4L9PC2mLBRbULLFn/PPWQTW/KBTiwruFd4LzW1ekVdATZRvSo2NIciwQ
x065syVYq6LgMe2IMdfm2DdZaTAlnNHO1M9RVleq/T4sUZmjmB4gzU9ZplMljMrg2QhHxXRYagsm
uofSwVrOzKQ3pbU6yCXajmGoUXmN5Tr1zVWZ3AZb5kZryOtHch5dmsThIx8qCeGqiccZ2mGJc1tQ
R2XtoTESUVKwawDPb5/SKg5aMvHqRJydBRS1uWdF5h3nG/5CAXDc+LjuOq8Lz3QpIzsZ0mVp3bPN
LMRAXyUlqNR7mPpRivu1C06reyvVKgEv4uYIZGLJ070IpMYILYP+JArl3bJIM0dPdF1VCNkIIpna
QQGI4vwnBIBQllGecPknq5MHtNfSENq7Ri/Rkck8WTWSas1DuEPQhNXzleCkOmzCA35greBsqUm0
ZDR47oD4U72ixklEJG9HPEVozjK3gf4Lala9DFg2CX+DFSCx1+76O26M+VwItLIKK+AqAa83YWKb
56zOUPZTD6ykEkDUancTtjjC93AnkNeXdtzP2TymdRabM+zGr/ZHw+J3btlT5OC6BJVvNUkkVWwG
FSxFBmTRl2E+FnaAvH8fDL6Y4kG6zqnFMDdViqnMkd2Isf6C0b0Cu0jhIjtI4RGmFE/hlGwQ0GpI
Ih7uhaQYtC5zCS2GA+2uDRpPkCpjfizGyKTQY0zow+JnfVJEDg3FfHGgyEwsGBZk2iDu8yJhs89R
Pup2A3Z86ZPuJlShzjK8PEpD3b0PC61sYGSuJLfI5YsjApOZrVSjILoDCm+eXhCRGvxAj5SRbpbH
cWltcUMUhOng9AQ0JWo4tk9fesOgEcu8nbi5QGyVQaJUeFdht2B91sIb2gwnSksxr6u7u1VCcpAl
dfKPOzKuCVTPURnKkIf/4iZ9JlGR1rcYRm8BxyZqyCQdFrzcLIquGl1M5AxOZYtPbkHOcAyHnQNG
y2lAqUbsb5gztBIpxzw8uT+qqb6s+mBNBx//bChdROzZ5yqUw6BjXGawwzpiK1gZ/+UxmPoNFYnH
77ZZu1QszgKWXLDJm9GOGm8raWsWohq1Jb5G2F/s4uN+rnqPLTOiv2C+mA5uZfqvSjcP5rw2NCtU
0SponVVG+U+iJ67rSUa9oH8LUglDWVVAYpqCiteDMf4etAYUL0tX/VS0+Od5kEiMemK/mKT5fMY0
lCBE1t4ylEyBVgnXt4CrT8bwzNjeWVjm5vVHSQ4ADIVH3UcrahpqKWM0RuONK6whB+eVKlHkwYW4
mZCmI3wXsDBIxYDJYEGOlLh0XjOXJcKi3r1o0ACBSv9iUnAaUcgG/2KLVTs579oLPobDup4de6q3
4VWkRlQz3uYKSKLGM9TJtDQb/r/rmQF6HBcIWactUVnfeFw06Hb7u/6sDY89kX3Jrb3BB90a3veA
YSrQeYOS3i/68ZQ55b8suvD/JVAZoPzsc/gl+dNUU+ds0NJ5eydb3Wg+HA1+WZNvnstlWkhIJly8
igiU9TpfBdelRTJ53t5OG5OHAW76nJE6Ck8srbG0dE8F+WvLe47Py+d3YWL5KP3GeKtioLTxfyD0
m4ZwR6nR+dt46E6cdDixMAf+w7hYPPOJ2fCKuh1Cs65ZznVYsB8wk2SbmTm+MkLIdXHeV9NG6vpW
td8zF/qJugmXLtM+ZMQZJKBBwucOszdbWOyUeNdtvF69yfRdZEOu4PUZl88AW74U947kleU+6eYm
5ckQuLFVylhPGClS1BuASgaUgfNtHeUK2qc5teUsM+hmKMNFTXPKeDvTy0MrEtAmyuQBRYdA21zG
7CuUxUhJZkRZzwmnjS8nO/54IsMwqN6OkOAOxmXPTtCO9FR6fgA8abLd/ov2lfbnDVId470O6FEv
DKCEoeXCDJp8Pdj5j1He3i5sCOW1OlRItJFA4yRD4hQB9IhleHH8x4QpK3zRupnMXkg93dRTjG0c
a2iDNqpgYOWY1Zx0Cx7RKQQWkWYYdFEeFMl/fEnqHMhh6hh9ZpcpV2Uvy9FqmVZ0yMKhQIVpgfx6
IW+oipqFrpwa7w1toF9n5PTIwhK1gttSyfuLiqy37RaqAR1M/DWuk1g3/xFD/h0MX++ssIodfmES
F1I/1v/ebwdQMuLeqwYrzFm225WupnwYauU5Njjr6BTTd0m/qdQKkpiGfkEUkb/7IP3ja/tRakZ9
pfBF5OytMQN8mXAOrfjFXXc2iBZBWRANJQBumgAIuYuYfeH4OPGkf2HiwWCIzIrxsbF19AWl/w7j
7XJrsnZKVmGcKoFOYiJzU+s+1bp2b0QTsMqjiZZvvCGlFc+KdXfqu6Hmk9be8wNF2FzJv7sGT5L9
hzUSNOzsQIX1WioMU0qMRpy53c3LZXay2PsKlsqkDaUWP4nRvqUkqbiY4Uuv6eF3LAAG+2WWzP/i
i0murSTYfddB80Ihk8LzmUqwqpqDGI0S5Qm6QNdLKOR1Nc8o3foyuqAza/Ar6R8pRVRdEC3BC3SH
MyOQ5mMUp5EY8hRSop3DlJD3OXPdnT5ClYELVldYisBg2d2poFuf9QuezpcreENP/yLdh9JBNXxo
6KlDJeX35B44hPjF6n9k9XtLVSkM/vjig8FtLJe/omGMoqnZJVd/RGJ0UE/BuTZS+3iOLKezdlMR
PLSO2HUgG79RY8HY5iBAnJqs1ovu08NRfmHlGMaD2Slc2R/aOreD3JDN6BelIWpN40uX7l5EAT8T
yCWxqVobwYfhK0KV6X1+ttaUr/vPMAVO72wh4hpKffSxCcPOAr7Djpd/qKpIC7SV7usgekbgW2NC
pRYUU08aMKZj5xQ5bIYi7zdQr/wQ+0GZ/3JwNDf58Q3AmShAleUOlfKaxkabxuSepsSC91C0KLmK
CdOdpTBfI+SEMlXmpPZlxzXxv6wE5ZaptYRYAtdslCyhbzpg4dlP8aKdyqAVZ917O/EepDud3Vr9
S/btz73JDSTREsBF5gay4nbODQtC0aYXJy6GUq0vLuln/bU3l5lTynYPrYnsjFhBIgELbZGDn7QL
InfGw2GI10qqgcJrAtSkKr6juYMNhZ1nGrFQOBeRTbNany/yBURv26MJBb5ubK5Fg4WpQ2AYpwH/
J1iDnVgqY3JGHDkp9ETJMHwnC5CUFPMGsnPBfc93oPiNL9NBoJTLnV1ZlNxEfo5pkXACsJyQsdSs
RihRCSNqkAGW4Xs68bA2L3WbB0eNorSkf8ecMmcxmI0Xtg/wV1xZZjh9xuycyu01GtbEldvLmUAA
cVFiL3lSbYT0BpPMzsuXLb60o2KkNydoJHkK8BI+FO3zYfFn5ioYtmG+skfZ7g5NzRB4MzwZXrNc
gsCI8hvQZO1uaKRe7bzlrN2dGbsEkSyhZjS5Djke2IqOdbq8S7FMUxSIY4PZsYxMeM1AFI+1sNwn
H4Y4WyqpJSH39xl05EwiMoRmwcLlCP77svNFf/DuoIKpdVffojbChFCSiDztEU8sAdHEQXUwgvkS
gHA5+42KYaiXTo22JfbMHN0TgRa0+TYOGRJgnSsuGQMZqgUVo2bmPnUCKwXzydLEnmW/XI05KCfo
Pj/bZvnMxoLiRtpx09aRlCTpQuvfGWerJc+04pwimFHYdFtb2CduetkLvg+Qr9eGUbKuLAn322cR
g84LomSJhyQjD8IsixhhaBNlscZBAYQxf6pRSIV40D8PIpWeLzYgCkB1bkgxvy77L8uEK/VJb4aD
Vvshmu4+ryZYEUlhIhrlT2NtQyYntQTL5Dvhoq2EpqLX6V9g8mZLzfR1asvUK8QLtBOMsIHcxd5O
O8DoTRZmxAdaeurVK/S6Y12IcnFOfbeB46OsFzLX0fcnFzHFWT3KYaTsKE2m0yRnhwY8aepMavNz
i9kP2A6wAiTxRPVFDHjCI/oONLMV4MbKyiOUTIiiARsV9G3jKAfLCrDML2KjV8GQuomCEg/EhSD9
PDeLsxKl/J61+7xdwVEKP3GjkRnw0o4APZqeqXCrXTQwT/FBT+xUMEE1j2AZ4mUV8z2sXMtQ203G
UFsyWqpMIdSyAUw/GwX0fdj/Bu11wOfO4J3npiSFfMFoSZxN6LHgkf4GKmO+wXt3W3tKf8fkfeYQ
5uk//Y4uY4taIMpR0eBgMl72Yk+GOgJYulaYjKZn2TTEBMe3h+LngZ28py+sl9kwvyOTgY6+dvUm
lnLbbmpVED10ckNgBqRFu7UqN74rzKhdl1paIed1C+a5oM593RvEv+QaxIaHXjKn9+aukXYCgh0y
6XvL+rr8TCPHaQMCXfb0pfWrDefvz8bOF3XWSRjLs2eX2NF2T+97kV5OK0sPgdwB8Lc2RZUtoBYQ
QXpl2ZPiDXatIvEPxj1GS/LTjJpbAY0Uf1C0tDbqa5ztGRLH5/GLVru8L6fh2k+nCNQHArjWjSr7
zzXkm5u+iGRFG2qrRryPw1fG5s959lISBk4v6Y6XLNAcCPCwQf8P+84IPVfG8bp1NcLZn+mUz8zw
34Inudn+15+vgpp0n0KrtujIeah+lRrcS4tTeAhRqPlWBwndZ6hEW6uZir8kDgwuQLMxtas65Jl9
zVUUkCPkKtTeVx9SyLu5YpYBB77U9h4mT0P2cUvUFnJFz17fnDenoMKYGIWrrOgjTVYi7M0uHGoM
q03/qvWBAcNVBMIE6ax7H+461ylkPs8gmXa6j19RBui2IL6ylfc5vHyhkYcyyxKFzNPNwFCcMk8i
L8xEdjY7klBpRrsVgDWPrBrt8CCFBxJU03YNz9pLQtZ6it5Sbns0zy+iQtLHB/hJeyAD7eSoOcxr
xVsoZUFvEugKq+GATOPwRzeV5Rz/hV1cTPIsuSMkcxQ6cI8byfmjcYQXAoGukwh/3FIdUgy+1FsW
FvpmXzQmivLxh5DsdvMo7SYoYJltnnFxxyS8CPQlueN+qNkfKhBE/dlr1FtYz53xUAPvCj+UgmZx
nVfBywNJgLXgrpPH+gPzsgDau/6jMpYZUWBR8uaQjqjXaZAkaI/wBV/vebLwQZMknfdjxQN5oLp+
KFvJVAVrj4Gu6fNZt2nu3IcWPbGWeWvshN94qsIiBly1esNg6a+zxohmbBkDpNO4+eH9UbGQcM6m
Rgsgb3xX65oypXK1hFn/EnfWwsTCo65biV1b4AOL+1lPZ7cEhu0yiCgpDWnjnyE0w4gNkmpDLIIy
zDncQ3OreJkBIqmamav8k3z9PFycSkUUreRSenGnauPKS+RIbZ9btabIKRbwHxQdvFvi9Cbsrbhg
C5zjoz0WBi/8/MV9tYPUmHjQpsv7AjQkJmSlMEFk61J8p6WXOyC89de2Mjr8yHW7P9sbGsVfdF5T
IwKNhpQ2zk5/wu60Wkm0XSQ8bUbocd4HCvDXY0c9/veqTolefmzwMLpO2MEB+MXL6QPrru4W1UQK
R0gfmyXYeEdsDuW6tlOCgTemrpnF3t6yybx4QVu2n6mwHEGvViFuxc5u4VxH2BuL8uXBdDPrHFEq
2E/R5H4BRrUNVoUszi+l2oAqTOFhnrfouaEMSUvtt33FcMr1D2qjaGEnsfy5R5EN9WbsrJJuFcYm
OkOqpfxKFmBSkL339hkUl4qG441a/7JZUsj3hghfK8BHLuXH8XEveRba25Suh4qFUKTdYIE5MN8t
J7n9TDynWbgPbF1sXqDcUrQsRPitTnjR3+iyToWXWuN48I1ElnQG8XVbSerqgPCWU3tbTbxoa7Dt
QkL9chHWLtPdhdzu+kme42BDUAWWbXx+D580pVFsfHZ+ZhdOG5nlIVaE1eh82s9Waxm9pgMBQAI2
w7TP6lFX3qWWua/mWjPJnc4kh8qjR5XH39UYQn87l+iHB5ZadHtfRPRDiyHewRkeVwEv1e6VrtHV
1BRSdttq3Kp2ELQbsfKzza8pVXqHyPI+RRWJUqfDVwVUa825qwrqZ09xfDM2PHTigQqYi0GikQYV
mnz+O7CNtd6p+tjWmcSzLHwGRvBnWAYb0jltmfp500KketrMPgaQAVy0cfWboPVH4MrYsbSohHQw
nkbKcmFKTlCYTakCNjDv61OrvQP67ut1niFzPlotqy6oFk3UGyyOl92Qxmn7oOUmj4jvZfDxQ5l2
yMhIVTSSN3gGL2UMNB+0pMiCT8z/jD1jT+WOC8k+ReXtASxg08apBDxdVK9qdNpcnVI4w4BhcXPx
mPjDFeosVMqlnkae70/hZiPLiASP+1wH/D6PlleQopnO0oeIQIrzuSfun56nLXeO/WevOvrltYtZ
z0R6197IHyCXujOVadb3oW2s8zoRKcHz1R1LIFpHedWSs4ijHnW1Z1sm+Tp1FtDPJFcvotFzWP1T
rv7vgL7aTMETpe+KL74QW7pyANxkLqIMhL7YT6q/wcUOSWfMSL8zwH8QjkkPwQQgarI3yeq9l6Ys
Dwe5zKzoeu6D1zDcLgJXWypnWneMVjTpSlLFemVFk5nX+DQhnUhck35eTt8TJfhPBaiA+wz7WfMW
D0T3O3h1uXv4QsFVQ1eX+KSVTNEOd/f/4qr8ToNT6f/tztVexnEdmGYdzb1G3Z9+qNheqvu/xn5F
ddvoLHKPsnDOfyaWgW6gbwtddukRtQqDXPG7AbCKouUBgp5+63steKUknsmbWOHr6Jjp9WShTPqf
Klbc6S5uBTHwqkTewglNQ3QRZM4j6qhOKQgpobhx9cDEnm4JWTNLCOMtOVt9Hw4VVB4Ge4ilh1Ue
iFhc2RND9EY1bG8Pehj0HFGoGBf5tGHKb599yjxC5Sy2WvxVxHFNujo1ynoHBwOG290NPWjknwTQ
4GKWXeHEgP5rzVx4XAT5AmvhRepIhotLleZpUje8U7FJnE5KqfverwLw5sQGWi8UZKmL8lb5XsWL
gBjvLX63iY0jEzjCelcqyF7W7C2GLbHsWMu/wda2GWwCQ4XDiOEE83Scy+8WSe7tJpuq2QIt2ckw
Ayd0zczKMGy0ISYIWtNBrDJw9hwx5iwJzswNgoHcuh1TKBRwURi+33E+qxRN1Qgzi8zB8R+3xshI
5gBIGAaRpd6OFZ0WGvgqNUdgkWjX+jbj0WLs7f6h+SqLl+QzvHBcXT3+ly43bMv5MHGMsGDjPOLI
JrJrI68L2V84Y8A9OglMa4L71diw5qExANMTVt8DhwObc+jBy/7EjCq2WNj0ij0MV6ERJFIYuBB6
7aj6NaSO4RkR8YwpGvscuVs2oJ2JDG/O18amqJrV7gC4c3Rkqao3sN1OBIuitG5tZvZll1nbz80P
u3qnnc1rGXoPtlCamNz9VaRQ2Gujg8SyyPCoNLV0+dgO27M5ZZZmJk4vuqulsTdqPGLwcdAkUFc7
EKn/NEiBxt1C8zczmbUtxYvgStfi4955/8StNYBYV8La4zmFiQFo52G1uTFAn5NtGt2Tmondymi9
tI3EWcjEdgReU0hKD0ZBTUHwfLQDKuJW+VnwVg7bVc3U1xcZu9GtO0DnsCVkibWP4N69iZmIz4Dx
XPxq49ev3SiW4AOT2nSKi1EkD3vGrmbqEtYStiNQWuSkV6dU0+s3+wNPjRyIXSwQqfISJK+vQsAc
T50A7n4MCRyW//q3SzWxLVXSaY4rzk3hhccVEqIW8WRk5bloUS5Zpwk7+Sel2QErem33TGQgj1lL
5PEhh5Z4iV5BXEfTA9cwgUr/M5ooJ/f8xMVeLKiG6cwtC/SSuC39sYtsC04wAulMiMYzAzbN8tPM
FN13+b2Mc96Bhw5c6s21j88cbyoFmqt4Vmgxb9u7RQiFLDGDDpwy0D16TtB01JP7GCF27Yx23ZXQ
bCVZM268smgSRoNiC/Rer7s9ftouPkfZJuqgntavgLgqtC0QyENKywd49IyLg+exj+qRWwPo+xfC
2nxQMoKqWYDA4UHq4xZKCvqAMjQRg/PPWTLeJMnVzPmLIKLd28vJjDSGetXoOfgtqe950IFDYlUP
k81Um8tYKn0Hdb6P/GLe/xM8oYU1oDUiGrUzaoj2ulK9Uf1KJATO49guWY1eHHZhsQZ4tEC1YCL2
hTfyhQ4MqRc7iUYuet7d27M/ndryxzK3XJ4zBD20MRVu4GcmI3vW2IQFF++Yk6zq8A0sbSnyqB/0
SzKATHi9+R84v31jPSPHNBZq2XqQ4s26FpXG1SXUOuelqUnxjhZydhGrizKJ2DZq4c3MyDqmEJSe
dUMZ3fA8G5P9jeiGqEA9A3rhzZPpKUlfuuEdXhL6Qmi5EnSyvLFuD+OtCelXN88nDrGjBeQqlJVX
VUl6KOD+ub0FyHnvyNpBITbtcC10PFsqkU8MBeMd2bIKv2JLzEiFm7kXDGjGiBr/bbruaPPT2kmG
ZB7ysBAbk20eZ63t6zI9R4yr4CSwYppZmkazaVZjNJB6nxma/EFsSfxKSiS2JevfJ04aS+egOaLi
R5skO0kGwACzekVXpfLlgueBtBZNXdIcQsv3EhT6dzScfNUcf5MZrSXJsQzwMVum46EPY/18Kjas
xh6mouFDuOhjRT5BcyOtPrOexw4HqDRw2mG9wrlQVcZUYyROYGNIXe4MASB2TwGRyoThWH25yI1+
yNQDWzE/BAv6Fju8cnsLFJz2vMWnHrSMp/p9t72Yy6Xut1tac+tQs28VaTQSsOFQ+knPNHOyYZ71
caOu3u5eBP+DmA3OwXHQAk0kNBYNYbveDuDELB68aAijDd4LbJRBNYlZojaQNgd94mXYSiF3DjL5
6fBXMTWWnVMuIPtvyP59hNDMNY4dPDbOwa4Sh2nz0qrqv69+x9uU1ogxyLgpTEqhNxrGcB6O7O1j
NUnYoSJsrvBTtlrBSGajyBQuA2mlbDh6e7NsHHw6YGDc65a5+5taYJR5UqjG4Bu1JVKHlslDal3o
ZLU2R41L+ccfjiMVaVUQ2PEkH2D6hU81uB5SSAI/3CCJIEzTBTpeoy4neCW0WzAuHq+JlFfMBhbn
Gd6uagr/2TMSo1/9GQdRYWkqL40oxP2zReuZ1sPclK0rM8O9vYP1ENHxFmdQagCe09VQcew71sCS
Z4OCyA3r7NMpuhR+DvX+/HTeck9tSh//FyBj7FJz1rd/C1kQMzG8XsClB4bHZWabrYQSN5jA91JL
9dvObTUZQQT+AhwSR3Dr3TKZuihpmZhHmnCQa/tSaHahglYBhfIuiVF4KDCgsr/BIgfZgIwC2QYt
XNbTYk5h6sF61ONtAUkB3B0Pr+t4P7AujrzgADQdmI3olNRyPogU6OgTsyPQeaBJhSuqOn2HQ2hc
+KT2uSqWT0LMkKxFEK3Ar2Veukp2rptQ43p+0Tcd0cFag/GZSdklRtcojqZ11Ef+d4gF8YLf8/eD
UR6r1NSTluB5rj5wrxzOmiEkVsvZf1jtXgvI/SOLt+mHM+o/wHPpcKyhZ6+dnadEeJ2YCHZqhBpE
EBJd5nd+ZeJAzCsKk1beQ1mHXnUZWL/NVaqyv2os1EJfipylGZ5fW1w9dmj7qbIUaWrOQrM8iqkc
HCTTjLcbp7MpTBwerP6L9S3C0ZSuRprkmnHMCEWmMC2VCyH4LzCztz3MMISBIdTaWDb6SPjr3r9k
NHVnNVMI7TnQlJiFIC77/fI8qtQunIEEbW2eFsnE8vDd2roLsIvKyha7IpTP2LolOpgf4SQqwCOr
D0x74UkKbXcRulviVXmxZdmtHhpVaGIHbNv3xBaXTjeiTVKmPp46dFGSyR912QRtPNWu94oFJPID
aEdJdDD7CqBOManUqyYLewKm5IWAgiScHHnutIMXPuOGJkFAcNNd5VrJwDCXCz5HJ3dDefNZ4l4O
pMFPKvN3WYtKWQa8gDmjD3lS8BNlz4/airyAygqYinqKBJKUa6bZ1gTqWDuEeYESlu7DGoB7ssda
wNLkAZH/yrVYpaA+hvA0TSCGOE1t/RZQjS3asAjccfYpqqiIK/q0S50QlMOeROssvh3C5ZRIMRit
hI/GrNWolRzki8t9Zn3Znm1RXiGKK8W74BrRLK7RS79zbZTG6i7FbU/O1g2Yw2VWIA2HuY3jPrxg
rj13lBihoI/+jLvaV6YdDEzXBKvloOkevk8VWX9oZZ2xR9/q9FE8XYbkctBOe9tXE5eNkcPaZidg
3DAAr/bGRA+aLeCk9CfS2Zr1e9wE+pJrFkS3G48ap2RjmK3/spYCqK4oLmwrPHJ6rAzmuAHnH2Nz
rd9D0Zo3h9VrTAugFzZf2YnEKowIqxaT1Ha3a9VFPKQadHUmrBggCpb2IA0GXwUrc4+yb0EfyVQ1
UMLPINvNVVZy/UKb8WqtSaPqiGFnkkbNkkqXDxUOED8kqBfkNW/LfigvOQaEY4n1ILjHqIc+zlua
nFWpIkb558Mn1NMCpHw0rvuK6MQwjwov3SU07CSJmQ8aKYU/lF1lsZJetHFh9Lh+Jw8fmcbVo4T2
aUx2YWDu4qEQdMlGCk3WwePxmUv2LC65Jq8e29lJhXApFclkPP+cWOo+XXNY0HxGjKBo37d+RynN
gnc1X7PNCMhCbi14SmIDcw9x14LrV4hj+VhSpHTbqA6DDfBJM2qGK23fKoJa54WCzak3eKnENE9q
/y/pkYv1UTxU4f/YV1zjWQXZMVeq4FyIfdZUXoFQpqg9FfjQP8E97jwPtqacM6jnwPrad71ybHVw
T/UQYXnCzsjXZ2gulOvrYSfxj+JdRJPv1X4TFyc6qcYhKsgcRtlL4yjFETE9MD1J81KFjJg4D0f/
RHU25NuMIP+D5n/MUj4mnlgi/f8Nm5ED45Dcy6VrDdqdB7KxN9xmK5As/1rNVH/ayKYorD8CsQ6/
yix+b7fXnrz+QVE+UUKd+Mm/15zTeeSOUFs9dMeXd8MtAxvqfwcOsMZ1cmfxk+h4Y9ujiczmip+s
K1jv3ooKMVODUG3Ana/kOa8HqCKTSwGAyDl9KhRnaBahA4wAlcHplz1WLvUtpzpkgKBjRqfJHoIC
Hu25DF6zWrJXTOZmxhlw/RqleoyY7TKtCl14rSdTj3NIeOL8jJA4VXA7AwsEdVjv5CAq0Es87E3i
cppuLGG7cLJ4UrhByoCBFaboqHmJtRis4MgEnhvvqIbVhQP+bJs+JeVQZP7f7aIZbw2NO3az4HS7
wcyYtpxm1tXiCloNLO8IM7jbcxGjAMmaCoSIQPKjxVbb2eKmQ5NXZ0/i+PC0LagxfsjT2hxweJlI
f9sdYbptag+iK+tp9CF9/eXTqYp0MljvifV0jZvCG3BCgxHq9kNoq21hgE379mUaciw3CmMXWuJc
mrFnJQJPnsQcDFsiaUzyUvbT/qis7J05f6bnAaj4XbjBc50bmiNm6YArWwbjAQskmlAGwJInVnDI
W70pOk2RCRx4qYD0HIMBVtzh+4e3e0dccklRScv9JQLgKdfSYmsqfquqXqbk/XYwcp81JVk9L+d1
XeGRFTCoR3fgbX7bZcnh9008bZD+dLj84hirVyWbcFvb0nyzehGpU6xaLU9tnzeSoY5CoDi3pzAo
5JUMkizmldNu0JO5Lzzen717wHdC1jqaUnDEI4cET8zhCgh5xabrrZJvygsLkjbEVudwkUCE/imG
JG1H5lo8UytNCa9o6gYaxf/iIDmkeHuIf3zoWbaPJGhbyD5Xnz+oA/NPXZPCpOtXpkr2tjJMVMbI
O1x07xWccl8SaLfIt+c179kRJxTNb2SZ/he7WH32tDXctCiByRqmV+l2d3vsjCqh+npRdsP+q28y
RZJpezQ1XngzAI8aHGnLYiWkBlr+xPmFC2deIgbGP6DLPjjmpDiIaMOlrsyQL0XL5+ZcOjYGKzls
6zojfQ1DWFJkE5Ka8g2iQVp/bJCf7OdEXEvLCsfzpt1XvrggLSaDsE9V7HHx7VwJrKVK5Mq5a6yC
GGkLngrKnQKOvUCqhAWE7lFMAPf2Cml3APA+UhITpOYhWcEkW08KB5PNn0iTEb4La4yaEpPaStt1
O3m4JlJulrHlVQBhFn16EIKiB6jZxWVqoliHvZsZyfYQUtb0aBWk8J9Ax/Gt99+MvjqaKnedG38I
TVGXzBrFWOw0TgsiXkRuYGGDXqqrS1XAoEbmbIlF8HmerHQmFAhgb+JZw3tg01+7bzoPqAnesqFD
JCtpiUccoX/mqNct4+KDIVPB49OCtpZ/x8PUrDjz0NYllp1BgihMY2BzzZrFpVEgBySg2vUud+fI
Wb+ThaZWFXqVOyVYPVZLEOoIclMPQMYkPE+I2iKVJX+qhuUN/aqdVOl9RSE0iFO5eLlwPYPGOAb5
oH7uVPoA1vkrxocH4n+MpwffmarEJ7vw3gCBxforhfshUiaNRXw6/V/O0tTLGChF/+jIRpnk2bYj
M+oC/iT7ANIt2CppFqPoe9umOoU/xYDfuwGmPlASFuCbCe4iwwFqkoszIgZl+j8fDtE+4xrEMJ6e
2H9DJZXSzhzovwlMwRlbY1rPojY8t7boRC5ohKNxqvFnRKoL63xQ0bLiIr7PPCyuhBNw2KrXWiNB
cUcStBwsPJM7YzOs8PmMK/JWoJ9mOpVACEtRFjmdqQl0lkdLNjkaFQ2Q95zOdGseR8kokMn8eRiF
Zkbiua40A29jFsDuQBcwYR3BscWf3dNjAY+uV2/h8wgvg6bdOwYdASzWgSx9YHW+RMlVXJvN6Nno
1h+qsbd0xr8A7QEHx2hfZGQ/OH20qn6KQBEWcRcG88uIUsquMhMWmblR2A6mExi8S7aSWVrgKE64
jGfKXlDch5by+aDsJzrTNZvC5baTRUqKyU2hb1bt3bJ7gyrIUz78rq3Yv+RK6PdaKXEoCzRxtdvr
wYPY4jfOID27QsU14KXnxLb9wVz/WVZg3yOkXDNOUvw1gHzGgmYFBWUj5qrJAFXezNqByt5i2RAL
QlGm9lnJ7S4iNX/+TIwHUi11yI66y8PS77B2DhZMEQ3s/29ZPdR9kqA+gLUvFDHmrFnu33LZphBj
jS8EoeJqb+apUzGSOKZ5wV57WxkOM2Zabk7intsDngebezWup1amQ2WdwqcdWdwKXOcRkhrDI6EB
D5NiXXDc+SmkPWitFzYQBBkREwtjHywI4Tvx2CbRp33b9+s6kLpEWvldNUQ8TaLSGO7OyiyyikE0
+HjVc4IuWY1j7B9ylw4YT3fFHsGQnDf0k0Rul//JJ5imL5JPKkmQ366cKpSdqr2XtY4pKb8VPfnE
RZCpXJCqsnd4RAz/s+1jQOETXj4Id68Z4uzmSgnlEQryhhabRkQTrWUqyAZSnEPWpo3VvkU0pYoS
9N9I0/yqJBM58VcWG8BWfTF7tKrJpIH8v5aLOYR8CznPZGStBlBzRlVS99Hs0kZK+cOD2pBJ+MVI
AfHRp61uLBYq1N1KJP2XqkgIg9UfC2AkJXzA+p4+rz7WG7MmpPYXVT5yZd2SLwGClUlBz2hf3bgV
ZXbW+MGZNW1WHMkqyRsc1Txm4DouNS2PovjVH5RYyPM5BMbn2cIoyzNLExo97EDEbS2gykeBt46A
afyKVkaQTDsgpfc0MncvtWcufLwxLUlZgBsL1nHq2AA0PPgaPg2wQvB9FXLwl/HPyXuDZIcUREOj
24Ru722f3BDTo0jNg8AizHqJYFuImhbX1mvnUHWvDLv2yBQGIPFpkWKAZBOWadJSSwtM8GwH2azq
11ou4QgOE1o2spPpYaSWEVRm6BlLzxYZo7Zybm+vl0RZJxh8QQSR/LuJVoSqu2IlcyCXSnS3ZREw
PB8CxzpKFpYV+OTt0/RNoB8iCq4MazUeYzQ9p1vhgAWSMTqIzQ1Y1ZXPwZRNlbsqsa4nRGnVYyNW
YndwVBuM+cOLAF1lQgWBdxhQ7RoOvJ11GDQppy7parQa/5DDnqhtYLgeCKA+u4HnLHojqpR0sGoz
+PY4Rm5V8UtIruNdKzBg10U/RClOFl/C2bCYS/i9qIfZdNu9TFjA5YDQRxNlB18n0zdwSrVb7zs6
pTvcI20hYxsPEHLG8IsWpgQnmZY4XFOX7RpZ0f5MnlbPVlxeRjOuRVy253RNFW3GKsmxNsAToQMr
MYauDwLiNB2jbaauWEohLbdRonlq8Y16FdeUNUdkH2U3RCxC5djKZ2FpbHyHTRvEDsA3ivn2gVqV
I3TFF96qY+Fn15WqAegtNKLgFsgw3G9lvr23aVXMY0qMHJZepSbFAqUP4v9ApDSxDToRyLi5LyCh
Fvzg2bv/dg0jcInRjZ+yfd2/6FDjFQY0aOwBRHsWfE4zx1I4Xo+7LhciLjIJqx09LdfpmfEkAE2O
iRtvv3UmoDl23uvfV97QHKcN8waDuMToIRnrAoJzGaWWH8IxPHyQPOlla/AuAWjk0vHZSLH2Qdv2
Lk2Ai4rBO2IkJOdTLqrpgtxiQFYDZ53+qIifVOHcWfT7YsJb48fFC1NUngalcliDMc5fSUWuGLAI
+1jjSjQJoJA3A3BtOEZfU53db6aNANIlJ8Wr+DsCW49bnZRK2rUBvEACCSE3B7XnT6dD14jnQ2SA
Xmu+dMINTvqXTWU0X4dqdzv5MgFoYbWGh1FMRxEppqf5p7mJTs/Fp8UCwauvD0gG/ms4FMSq5CMt
5VDKVUK0P4q/vx21z1T5q3GGJjWO/7iR2qwuBueJk2nmtPoWoG9wSGZyjLcf4+BgX/DJBGxXEYVL
UJ3nBd2vEV+qnF+ouSuCeuOKfwpZZU9KPxGUvFA288JfW6h3HOeCotLe+d8BMHLM5KDbspalUToZ
LSlKS9XZFAa+/5voIAEDI/qTvqekvZ0wYPw39FMjCCep0IiiOJ9N2Ac9ahXGsJPm+oCs31rQyQj3
IvYCgBzxjD+wV5up50MII+/1UMmihqSkrEBHyD+e6rjVyKXb7yYVz00ybqc+M6kGyCVOUvusiXjc
1seKhI/lFZoEXUSACwX9k26rkNe5UeW3y1d9aXE9U4kV6Wg8abF/gAAmwq3+PkvT2+qunbzBix2H
4jTNMJ3NDV510cHAa+fXvC+P+LldQiAvHeSTzJg+M4d0OkD5Vxsukwax1mrBeN4rHXJKyXGjQ93y
JVm/06V9p0f4NX0v2wiBFCxi095BSfJEnlRyGJGHmHGrproOlzt09zzpR5UiC5GmHgL+cRsTSQB7
0obLfOJxbPPNT53zOs+UKO2BAWoBTvy3mKYbBobBtXHj6GSbgaUxnf8dFoKD8I3956zL6tmyqNL4
Cw60IyubzOavubdiPPvGL8k4z5wDFj6bAvDCvyF/ok5Lkm2vnPXySpl4796XWmzYN6bkw0jzfUpo
ityziy4uGd82cvb7KxPPlrR99sapVrRqlKe47m3QFrAyKi0lDgCNNh17R2P0EYsECSLCn/TR86Ib
Rz8LeUPOrYYTvcfLjQPAbzTqAb8KdOLoQydoKc4dHmlm9hflFIhmDidl4yk8gk2DIYPpCVFLAg8K
bnRcy4LU/Jcix+qwgY8PDCpvzTL5meHtQWUdCSnY0gNknTlCGuKK3zs4hu7wlUaAilSm50OCtBYd
Rr/ZDiwa6mETHsKJSNKGehXkA0KbUqXrcQWEO1kiJO8iwY/XdFfb1zE80udw3/imo2D2qMrus9IH
6cLepn570rlOnv+a6f3sfGywrO35hbuSIfoCAFICGJ6glFym9/vVc1cAhhW2VDL6nvScra2kes/l
4qhtPosZWKG+zAkyYUs+kzXUNYagK7+r4iNRS3CBLJFSnwpq2tPvZ+94pDGWWsCSSIZAJ40VavdB
NYkWHntTscWL/6mz0+PhRwz2ZrW+FxMpitlfl3z9B0BJ1NSnjwD2iFVi8yGn6noA5DOtvQd5jkYU
35wtvHKYYnc+HboP5NTOAVQz4S1xf4yg70Gmi+m4SjyIZ/IqCCVq/zVf1FdiwRtaTmobBbojp/gy
DddFHDpkY3kQCxQvmZIOnBMyvjBNEopcmO7N3rTJ1J3bsIdfp0rfVmVh7njvW967wvhGlIlWhG4u
JtOYtDCRqY1LVQjgw+1XZR6212YH7N+8usncWaGQBdnM0ij/V59w4unvBMdMwsNT4CyzThxuRZWd
bkxHobCv94wRsPNDq9Ju+RdBFp/ofi0v3AM+LyAVxFz8h37hAgATnSXtLX5Fex3iBGcDWgT4y/kw
tTpYAPwDmOucI6+FmdZsp7Zs+EmVIvd1pveXYOcfYQ0pa17qyqJAoqA3A96EiLcCiZh4mMyeHdqJ
svV0x1aDlDR8FU5ubXmRzhgPWRpruzPOvrkXk82t5k519Ume26ElyzHKFkmg8NP0x0NrDn84ZA2F
XgACH4BWvggdOIJl2QpO1FLglhIVInCsjHv98r7FOnDXZTaC9TR8RrYCgWiohD1WFxewZR/s7MfR
TxXB5Yf9ac+0qxBY4B1pwG3OorBs8YV07MaiBQPtEfIhx7pDFZUPCu6KPyAnHVb/Mm7GAUU5bQje
r8+OUwZ9SdhRSFLOUHOhfXHr8QGzFAQ0cxxBR49w6vW9pZCfX3ZG9M+abFoQPMbkAJ10rsThVXcb
g+6cz7wt4aDbq8UPjzny3uIOh/kDZ9B6aX4RJdva6F2ie68NNv6sjBAB6nVv+agMr/qR2z9hrMys
PMr3Nls77+LTbb5Rt440CRzQ46AGy5LiYGpcuUz4X5GFKcoTh9IINNB36GIoLjn3+5/2PRFi2317
9PUZX785wjKrsRIqK+hfivEqCRAdWHYDJ/6EpN9xN6uod5j5UNl8Is0gHKjvPv184gtFVF9pxpdb
H2yvAxfii/zijSWMZ9k/gB2/1zkXxA/JUgnqZ8FxJgnWWdYe0Fput5r7GcxpfDnkaZVaKtU6wLHE
VMXDjDSTZxuIQleKewMuhM3Qx/bLoM9rr1YnRMBiHdKKCVtLnEx58wLRKoaDZEnuvGTcBZDTanxQ
lE0pjghkgcZcT7P6zv4nQz1Y05FBRUdibLTpKx7OpJ9A+K5eS2eb3DLoi9GePMQNVMV9yC9+mskn
DQQUFs+KugH9u4FsteW/3ky3vKzbeci8c1xU4GwdPZ3vZE8aVab7VCv+cNMh9nUxZQUWTe0f+M0o
mLdxwZtpJRSXoFP2jm5Cax6GjPg2Ue9d08dZUtX2Xq6kz48h7suRfTvDKIfhfhFy+XWWaXmzsF2z
jJPFlOj2oWVnJQAGON60IbgDoV907HGCGspRxLOvKpcfCyf7Cm+Vuu61wlfCSTuh+mXUIuWK9PcN
mG3lqRFYavf2ODxrgZP60dSaTq2YgX0KxxN8X0jodEpjEyJvl8rwiZ+y+EXY0S6abKCwC1F17W9N
FCckXMFM2BQT43TuYfUwRpg+Kzv0DByJrjUdG6/diauiacLHKa7RkJb9qH1OCUcoLe/ciFiGGNNe
/Y9ifjT8lienV7+7wrucaVICIpcQg894ht1Zmi+/y5yRD0uepTNbNBUzwmzrfZRuvb+39LcgmTQc
mxJc/EJ4+28x/gAj9cAH5tMN/PVU6xU4HJSakI1wFYth6uneZYasC3sLGe9xKvwvgBhX0GBkg9oF
aw6efWQjTmO/NXc6UtyJrR4hASWNUZUSxCMIImg/q+ynG1k6BPyuTFDBtNfgcRM0tsHuNYOPPI5A
xRNB3FVeEHjelxijRumXWwx17P1PD+llhbUjb9MZidTDWekj13TsF3yp4CzXkbLUEi4J+CyC8yAt
GQWbEMCsnYw2fpgIPPWUeENmQ6ZhaVMkgtNyCwxbUEMVxQSkoIV+GXHVH1BXDx/sWWNgTcLf2jrj
86T/vSOw4w+4nfA9/M04IdzzpFMbCJ9TmMAdFu86mZBPJNo9pCNykuIID9xskBPAsVNvSgGepPsy
+BSHROmh0XgOf5ojc/zJZhULVVbxZrsfav7nDnF30Kps/vmbcqUkESY3uCW5VcDSBUGAXkj33wmd
mHfBhtdz+S6fNtha2CyL68I0uPRHamccbF/qYTaS+PzNUyihCD6BUIvDsQMd2hg7/lX2ZaHCQIYo
Fmn4lFbEq9MJvb/jpMLYywzy30cY5iPLlof6W7ycYYwxRuS/2+OuYMVlyO+uus8hl6CdaIiCXSy9
NIQ9LYC7RZ+XnC6jezbJN0/MKK5dfv7I6kuxB7RqdZJBPmsGQZ9rx7AbkgMYLs4nxkU7Q8BY8ZS6
rH/VDAvn0m8puWjKGKQHkPejZT2Zd6bzaA97oAiUOOGzd/7Q2mAerhJGO6dgq6+KpXIpC3e/B/ca
BUeb79o8DMHdqaRNTfHXAuQmAVSB6L/vZ2vdCHdIAdzRnT9gIjgJPS1XCSkhVs1+jLb9ZO5EthfH
HafetK0x97BcefsIz/rkRnUEp0FLSyPZgymUzE8ht29rZknELxxhuQkJjreOUEDqt6Q+MNg2skwk
6KK9TUinY+o0poI0Rlbuxzzj5OSSDfaVF88ZrLUjYoSTo7V4FI6vPca0FdxiLvI9263GHLvUXA7m
XJNkgcy95vGt3YUmcdCwPZiieMUCx2r9bSxexVdR4rnykdzlFZ7GjP0JcDuPTb3ucdeVxF3Tr8v7
R1ybVKjFryr+EdbW/yLqC74bd7Z4NXVfoTrp0kbh8pns72L+IxDqFNsb6dcrSbrf8mrtnTddL1Y1
8fsJEilgHuMNS/TPm5yoau3okTAS5ntXjP8KVBw17Y6cAKsEkg932DAEpfNJBwM9waQm+iOO9jcQ
UG6IMGLg7briHOlCVD1bXQjgy0YYXtks4WG3gRRjyteuJjXDhdKYb358z/7rxx4cghdN+5ypObQI
Sh1tuvHy74eizpahGOOmKPXG9ASZD237IH62dV/T1DIUo0uDaJwa3ub9ANdBnVt1VUidVf4jnGJ0
dlarDsQk/bhV8/15r/wv5MWvKe+6kqWFZA9wf3jpjsPrmqdbrTaXEurBOvIC2DJxNNJsBQ+D4/ZM
GxpN2C/zwILybMpfguogxQNIcJStBcHYc6U44Geck2ZwCze1taCgymrNUzbKZMbiNf64ipXV4eAD
xDxj9bzQ9TJ/uv1FBvbEXbyKxwmsu0PfLSTramzvsHYjNsZBgOicqLCYFAN4XA5jCPwrCTxnfWWh
8TVybFkGcskFaSCeCrhM1tGon+tZIXFPkR7aGEiq+pPdi2jWvVZ4EjGVF2+pLPVv81C9iaTc4CCV
NxSqEoi53fUzlz4I4oP+p8H54wH+dyWRAEfyn5JuqBrTK04+/kv+ASAgoDnEM4CWVBL0EUF46YuM
gZwPQn4yEBM7pE+oRKaJ9p3vhtqOVs5nCVykMEOCGOMXN7rjNDfa5oX2chYBWYgVVZHozj/1wYN+
w20CAzu5vkruBmjIAi6ux/Z0JxOa1rqo/hGvy6O5cTE8AxkyN4JQZ9oW/XyADWV83JDE3fetvzTj
QM3q2s89SYA7qKNC6Gp8ItBCOxQN9fULCaniO/4WiUKG9n39zMtQp6/9VCw5VCf5vaIjWQMViV26
baFSy0iHikc+iGvCbTrU+cnmHdeZTJtmu22Hf1bOy5sS3xmaXdhMrM3rMVGYWXg9c3Y5abfVoVLa
acEPwtU0+tFTzYDaBLoAzua3upTL+AneUwJjwqAVCs68+5BEoGL4PIAc/Em3PnOgzYn+1Yvfxgrd
CgBpiraZH+IED0/QJSLYE3grijhQIG2itwXR0Tb1Jm4IPYvpN6s5x+pNzZFQjmwuZEas1RUieXVY
B2qO+O3o4jKqTwAyX76F2fgI93U2OLTukNYyecT4YSHmbXcyahowVQDh8+2rtalnu7XGZIjBLA0A
0n77SxXglznEciCBh/1TBwV53fcboNzeJ9RjTg8VGZfd3duQgx/ggA8sKuMYGvFPN/KjD5Tpzau0
GSLm5F4shM1GYWNmrY2nI5PVk/lcVm06uns0CkFP0GKSf4WyiOxjgU8HjvSNO5fA1NXPWyOfKKKP
/GkVL69yCt65+IPlIm0Z4pLmdZCR5QOtUAbFqGDPRGcPz+qxsAUvV5u5z6iqmbN2rTZUU+ZfBkJ3
KRA7L33y1L2MSYVM0a2VWWChEir8fxMWpX43948HG5WAmoxENWcnu6q6WzVn0Q6TSQ6EvO3YksVD
AgRxweqK+SY8i2Ln/a+qDQQAgHXqBfqnGhNHtO116jbaIriyANnQgHyjFhqpnskm66kSoOmJQrR5
1iJkN012N08TWJeQcHupYihFJFcx7/YGWVuOLz3rd6WwagvYUEDemGt8f3IESRahg/g10hZ0fT/h
I7YXiucHs23Sjrzj7v+cJ9O++QOSxo5KjPuSfZSGrtY9i1jQsd5PsRPMiuTm9rJP1mcKm0Dio5tf
Um86FRCDtGKsT+ljRS7oz6Yq719egI+hTVTCaJtE2j8/W+hOTVDRqV060rN8NipMJiSy2HOhxodE
VsNfzx0LqjBkJrqzMavaxDADjo50fZwaRJEJK47Q+rcp5l35BRQuPAsuP0Tvu7hU6cqUhSKUuOCu
l9rJGRQaZbJXEZ7FNLvfXZO/LYiBscvFHqntY5lapulw8/jmuTE5rHJdWkbe9wndpathusddCkao
lcqoK8qcJIyotDU3wpyh5FdPW8r4njdYLvxn/hPWFUyJQ4otJjxvVQeujgbidisHc7SvYuvenlvx
ssc8cTzgZ8/iJdZlEFay4s/aguQwjokjv0O5yQ4T5GS1CeVX2+04YUueHuldwZ1rWpH93ivfU+Cg
Kf4W2tB72w8RcG+wKQKYJ//Ln8pvuLBbywXW0nDjBRn1AkifvNmk5CO2Tdz/kbiZsxzRXt0vHbVa
Nuzn9Ha8QEOjuy8bUqiYjPKK4gHfZbxjTBEjrkENjNKgYxtOtUFfj6KNjwYOB/THMhEKi8jbA8Xy
UnlYuQ9lxcFRS/vk6A2jnjnZdd1jlb1AAJXlfLzSR66FUPznlQSrNQSyY3QWClpV1J0/Mk8x0YEi
qoK3yH/LTwNsiGuwIkaemzYpBBpVVqLro95635Hmj8t1YX8rsIshYm11hsBVwvkysQ7r5VUW0sFj
i3j2GqIIWC34URIuGKUSJW75iJCNdHMEtHQSnnC72TOyjFzcBxlfBT4F5LC/M+YPpH+38Da8BWfQ
Nzcns5PIHygnxL4ONWw9WJ3Y2s21tX3yhm2r10kEMvg+s/thXY0UrGBzovtahMcuSgfhlvQg7cdP
GD6GLCwchCj2nUMbQ//sz7dsjzMWnrh27qm2VVMoOuOPRwSG3uecszttgaWEH8eLyV6M7FN7T6or
zdWRsrZ3wT+mivUYgGpX1kbdvFOu803JiWfv9g4XW3GJXUVXIZPuyFlyOsKeCd1LSkKwAHuwqE7j
hGczDwlu4pum4H3g
`protect end_protected
