��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�:6�E^�F4���T����G$ɢ6�iO|}�:U�x�ct�O�,��(�阊˒���#Zf*�V��wD����ק�V�|D�×�+���x��;�;nX&���'E�amY����%�#�&nh�H�|�%�J���$M7�q�@F0g�﹎_؉4<�3����a�>�/Z���J�t�r���2���+ۥ��(���C)�D��ep�;rz�m�Åg��P�30b��g~�g���fr�ƇKoI/��c���X���-�p��hL��V����w��wQg�x�犱�_-1�<�r�D�r���헪���'*���8xl (�xb�\2�}��U�����ʯ����_�u�;e�.�6��C��݇J��&U7�=T�?嶻���Yc-G���
\����$�M���Y@��������&���~+ �+��'G�d���?a��]�wŷڑ[b�u�p}���|������(��;������ʸyL$�����E��n�-��߮أ@Y�{ņ�g ��~�oc�޴��H߆r��<H/;�Ux��(D5�T�31ax�·_Z�?FRL���I�� {I��f�	΃]�2o��e�1�� �X2�$�4����>�_����_��e����8�q�bw�~}��_f����uT�x�{8G���7�Xc�����uo2�,:1���v�����h ��5�Z��ps�C�"�hgk��~zf
[j�)�L���>{~J�d��_~��Ix�f�ns/}kn~�����'8�&��S:�7�7�`��P�g��w�Pnv$�gP"�r�L��4@��>c|s0��Ƞ�U�)��� ���T�\9���m���p�L)�m���V4>���V�]9r�RGr?J� P��P�T�B�X�8{���r׋��0�r�l�*�.�w2A%�pT���YlΛ�\�����9���I
��T��]{b���)Mp�5�D�����</{*��#˙4�a��Ln���ERL~����J�ya?';������z=�VWE�۬�u��p��v���� ��*x\�-��l@���m�KJ�l�vc��v��=S�J-2�d~fQ���x�1N�Ku�:�I���\�{�sF�o�6�j=7`��}!� |R����È6��N�y��x1Ϛ"7�J�FD{L�D��,�TJ�,ޛ�!�X�c�Y����L��O=�:w�4PIM�סWQ��ٸv4�x2[��(:�����)�qo�>��`��W��R\�7��Q;akZ�vn�hBJ^�,t�,^�t
1���$r�C01I��V��e�j�kS�;G#_��.[��	�Wg��\}|����U�pIπ"�ǥ�����[]\iұd���nl�	�U�I�����i��M��$�����9�4�]�י$��|�w�����.�x��\&>�r�����\��h�%�MZ� (����Y1��CU�EJ>���qL&B�^�Ͳ��o|VvA�u-�����g�f*"O�Հ��qA�sҜ�������B( B����	 �$dsCy����)o�A؄y؍Ao��y͉�Z��N�s*��b��H��L�z\v��=�Q�P���p�yoZ�q�ƞ© �C}_��U�5t���M@�m�`ؕ�'�e.�iD=j�筄�� ��C���t��9�#_[	�x3f�m;�o�q7�V�� yY��s�-���19�bC��R�%�Jhs�_�ci�{�����'+��9��mI%�9��b������񳴩�w�H!�x!�%Us�֡A��HLJ���y�F��oZ΋g)�,��9K<4j�d�KpJbJ��\��_+7�z��HP��+E���!�鉳�n����M�y!>@*�L�:	�Tq\�1���}�+@F,���T��0�U��	��JTe8����&�����H�CQ�1�R�otɔ����v��	zc~��o��eީb���R$�AW�q��a�׍eN�O@�ŬU��.�?|��t��JSƃ�]�ҡ_>��*ԟS��Wϻ��=O5{:�$n�p�Qhi`�T����
ni��=5�O�������QӦ6�ܳEq$(��k��u�t
kyXK'�^ɢ%�Rۉ�n��.����Z�K�7�Ǥ��>Qsp�&���ov�$�'P�Xߓ�����QZV7d��O��f���#j!���ٺ�?;�����K��)ERI�a��^���>�Q>1<ڝ��Ҵz��5a����7��&n,8@���&v� �����P�K��z�w�)ޅ��?O�}��նҪ;�0��g������N,�[��e�=�J�y@�n%�&��Ǔ}��DQ�X[�����XDj�,��X�G>mO9��sM�ݙ���(��ֵl��Pf܅�J��6�����)�cH�T#Ҏj�SJyAȜ�e�*�z��rW�Ћ-����4sj��%�����x����0&���GÌ�E�U����I�&��k��Ԍ�l���-:�� ��-�����)C`5��<�-�?4Ob�6�e��I~��j��4�ƹ.����M�R�&wr�0
xx�vt�"�s��o���T���,�nG��y�h?���SIdzw��h�&nUC4�Y\�f�խX�(����~c� E�F�q
ȉ���m@��''�I��uN]��a z�r=\!�ěZ8���(����y�����Kq��l��l������skfX�w���6`�]�����&�c��.|����G�!���P��&�
�G@ �_���EYyO�<YҌ���Hd�{_?Fjz�oj�'��>o_��U7r�q<."�{P뗆0�$�]D��Λ�a������:	�Z۹�ĀNw�l�c����Yb��#|���x^-+w��ɲ!E��е����_�v*
f+]�uc"h68f02�[@� :t81�oO�,�����`J��x|d����R�|����@>��|�Ƿ����-��eh'X��Srv8M�U)]���8zRC�����-z�E2��)��d��Y�J'�곉��K���呈�-�� xI�O�]�����6��j/�,,�`ac�S!������)��Zl���%Ջ9��R%�Nӻ�Ϝ�l7��.xj�|9@"��ۻ��g����"��� ��>]~����o�ẃ�S�@_�t/���6]g�K#�@d�
���?��-�f��U~}pHL��������Y0(�,;�e��f"-����ߴ��UDT������u=GF;�W��Y*�u�uƱq�B��_G^��Y#b�7���_ƈG�@�}Uf/��/ͪ�D����U
��(����eq%H�#�GǮm�)d�u�*#��$���׀,y���X�y��w��S����Z��F��B�c
/�W��M�ê#Ib�=8'��u��ٛ5i�Ã���Mupc��S��Ll��@��9��a��1s���E���-��f�K��h�aI�ٲ��GR������2ȧH����bA���h���=�c����;�w0p.��)�;Q[�I��̈́���{���ː������N��<��"ߵ��ݫ?�U�3h0_��S��͏��&$G���0�~�Y#�r�ɦ]�B����W��a�7h�J��j�rM1:+Ms��tc5�8�Y�W�H�f�5H�Ĳy�����mv2> ����(���/R�ŹF���/�5�<@�	�����{x��<k��U��"������mY�$q���%��c�풡����<�
�.i�$���2=�}��2�r�{.�^G�Yj@��Z�����e����x�/�"��.��#�'�ǝu؊������m4�4\;��Y�;3e�IЂi#�w��|�� K�k1��B�0D,��9l]�iV6}�\"����������&�gWq;Q�_,�8U��p�5T��C�(�V%�8�ړ gY���*�l�l�4��nCp,�KP�VJU��!�\M�K�h��ܜ�Pq��]o�ѷ�?�F����s�<Xțo�R0���*��Ψ�!��/|����m����[ç��߀�g����W���Q����p?�Xp��,����(����=���4�cP�=��[�@Z���|o�rG�D����2���W;МR�����3�(e��	�6�A|a6ц����n��%3y����[���ؕ�z.��a��	��b��Pl�����IH;@��.�sؿ[^�P�}�"��7�Ss�fa"�T��6\vL�ɵ_�X�8����kA��"���q��]�A�C�p��>��=�g�B�H�� V�������	-�'Gr�i��*x
o%0}�,��>8��+Yp����j��h!
�m�k3�]�
ध 1���G�T��_t�)�o<'��X��=� �P�����
��WH����p��藐L���-�A�L�kV!�.,-�A��a�^�Hٺ�蟊W�u�[i+�'�_�Ul{��0���c6pbyՌ�k�#ĉ�ba�#��)|8@��n*L�N�	,�(w�-�i��f�dUs{����XE㑲'T܃U�骹��<���CSAPC�vO��;c�>u��,��-�/i*m��QFS��L5��y[�"=W��o��|u0�q�n�~E����;'g�E����}�5"��r�-u�#i�_Rܼ+�'���X 2�0�
�7	�Q2�#t7M�K�p��{�:A�D��)�C�k���N$y��/��������DLҭ�V��JJv¾Ib�'RC��Ϫ������<Ծ�(��k^<�����fQ8���P}��3"�ˢ_��Jh��S�� !�&�nјa���(��,��Z��̀�fb�|C�T�~�]��;���|U�%k��N|���~��^)oa���\�[� �ے׷j���*Ճ��g��n=�$�'ج�����t�^��y��gw�*>�U'zDk��O�5r�����%ĴP�������� �iu��AsFv���Է1P;Rjڐ��'�$�Q5�9b�?N%9'4����2��^4�B��*��,HY�SL�?�zSzC���#:���{MB!Z�T5.�zB��f��x�
�;���fk5���4E��ɔ���.��9N�s�1��HoIlzޢIm�Z1�Pe�NvMj�Tx+T�
���ȟ�dOi1��\p��,����L�����m��O�
E��6t|̿�� R�zG���5�E�p�g|�ioH^{���}�kי�'�%�����!�$�K�������p��$�Ͱn�}������<͟�HQ:����=QD��/�Ԧ,O��i��o�o+��{ V�?_Ao�-oH˵U�����uPQv��P:#/�1���ɫ�K{���S�\�b���C��v��v��_@�>�R��2v���|��_/'}�?#����
mB��<�N�G��5O���<���i$D�
��x�g���6ÏH4-�㇓/[j��B9ޟ/^�I�����q$$V��6]T*ąA=�>C�5�"=kĨ�7X��E_jӘ�.X]%�Ȓ�CVks�(]�A�Zs!њ!�4�C!W�p��S6��f�Vsh��f��?e�W5�\��L���Q����h�OR,5�W��|�cb!X&%���O�'�>�o�W��5c��ęC���i�aN�"���"�&�W��Vx���n �V��ў�O�;^=��`�O_FA6]L`����x.R�&�]ᙿ�K-���Z�?��9��}�5znf%5� ��ψF�>q�K�S0Qsջ���P �S�	̙'���w $��.�4�{9k��\Ĳ��Y��Š�H�����B=as����>/�t����g��"Χ����k�����P��d�ݗ���<�΅J?ӂ ���r�3NG<��'���ȵA������M�G�g�V(����/�:ϧ3��QlE���.����S���ΌYK%�s��y��u���@��l)U��Ғ/�Ę� Ҵi^��*߳��=�<�Y�M�Ƞ��.�8�Ht��A�.��{
�2�X�#�k>h.f_�4US\o<�)��*X� ������e�|M�_Q��T��(o���=D��4���ރ�*o)�$������t6��]y�T�`��q��&9qz��4�� �9�,�5(ն(+�
{x�e�|C,���?|5B:R��*��I|�����~i���7���NP p|�Rt���3���i�K"���	G��l�d$������Zj6���T��D��d����i�yyyx�5�g?y�Qͥ=p��i���yˏ�m�a��5�k�~��ߘyR�B�~�0�����>�EW:0�o��Bl�4��0�)�ԁ�g� �0x�����Q��̉�l�eS<�r���AaT��9J���9���_��x�3򀬮0��ߗ׮ �TQc�y	�VX�&��XhРDt��;�;f�X�L�i����/KbI��S�;���U��&��i`���������
Ӯ���S��PF�iEВ3����LVo㇃pr�d>P��:�J�`��ۚBO��:�hIQ���c�>�Ҏ�l��-|1&N�]g��ۂM�un1��M�A#�!��%�Z
#���a� �d
-aI� W
�R>�mC,�MgB��5�����I���|�_��j����Z�7�nwB\��JR%��;z�+,�E��ʃ),)�5�1a�#���2I�4\6���P{�(U�!�&{x��5y�]N��`������܎�G�n�������K�+���\Q�����^�&EpV�-�{pkH)�^k�[k�����_3(_�fe�󉙇L��76�(�,R��Kkh�c�tr@~�(1���JG�9qe,��YܧK������Ä_�x��@[�7f�;.���!�g��m���e���E*!��T/��/ڵ�9�k=;�MӐO�\�< 8�U��>Ï��:��􂖢��B��1#����:�o�Gj����I�jc�� �\} Q���g@�H!+-	����S���f�١ �
� �0�'�hZHT$,���@/��if��
4G��G���**q���;��y�x�lb)��CU�0��߁��3�L��Ɵ��+72��b(H�s�����#���Љ���ʫˀ[ڧ�ۃ
���l��U�!��-s���^¾�ik��X�@i���$X���[	FZxq6v|�*�{���0�@�F�ZwQ�49�BF��,��8�V�����q�b��roPs����&�ot���뭟�g��Ϭz�]����*�q  ' n�<��#�)�f��P�R�� �
�qՇ�o����g� ҃pb�ϗPL�Z��"n�-K�`�wnE����&�iV-���9,��I�pű��Nh�X�k����0e2~B��|ѻ��W(�V��D��X�l�yX�t���O�����0�)(Gʬ�N�͙�#���sTLe�j��p��
Y컯����?�׹x:���'+��B�����*5���{���Od_��~k]�U��Ep�ǳ�e#uP��ԺR9y.�$�xy�#-,]R�,�S��%�&����mš���JEy�Yd�D"r�]E����5����b?�{?�;�����	����|�A��{���������@k��`���=��w�	Fk�R1f�+@^Q��E����0��R���ٴї����އ[���!B���5Vo��jmP�_��K�C�7_�w6���u.y}%���Gd�)��5���ai]&Fl�7[�K� ~���å�v����ee�/o�g��~I��.��e�D�T���a{�{3��m�Z����oK�D.��-�L���٘�l�ǊT���������L$Ю2��?O�U.!�/���x&|��+�vm9A����l��c��&ϓ� J`��Z��02������P�����yH=}Q6�Dc�q�a4���nB�׆�l!c6(4h���#�S��t�`W�K�������ͬ�R�����v�C�J�E��x�:�U�����&�����hehn��1�*D=Q��z���σJ���nΛW�)7G���e)��/s3��G����s�h�B׻���ߥλ6HF����Kp���?J8�bZRr1+0���z�Gܯw�$w���r�0,g�bͺ�jY{��#���fO��	�j?=��{��3-���!đIv��+ǝ�B0��R/��<��@�	<�NJ�t(z�%4W���$��[�/�r��qږ\x'��\6����̆ڜED�=�xD_��PtQ�Q6!!U��~t;͵�T��'S��(�K�y�[��[�!ɴxh)�/�i}�4h=]g;�AK�J��{Ȅ��9U���p�3f���E�;�r�>�.6��=B�]�9��slj�u!R�~R55���և�c('���� ����v�uP���������۴>��|�;E���[���Â�
�ő�c��4P%��w��l�^+j�h"�'�i�8m;�`���@0�]�=}�Z�#��2�T�)����<�G8VT�m ��s=5��C�;Q�!G>YXC_��t;�/͞��8��L}H���V�,a��L9���H��� ��	q|F����蛩�co�O��RY��;����Kr�w���9�W%�{\�MG_��� �@�'��ƚ�Ø/����Y0�0�j�Ks�-�k�7��I�ܨА��K���/�IV���
W����0~�(	�p=��� Ώ:͏�g��"ʵɈY�x�`�N���\�l'HP���{\����6�S�P����̕���ZZ&{�tu��n[�ИJl���0-|�,�U���qqME�Vvig�h��{��u�GQ˴��/?i�Rnn��?)�O�_b�L�X�����)�����Ԗn��i���,F:�T�
z0�od�Dt�{r�Ky��z�O�Bj�j����͙ǹ�{�4�H���[�.5yEͨ���Q8ď�"u,�F�v��p�H�����O�؊�Opm�ͻ��0�B�5�j ��4q�l�8d����e�4N&����!��@c��prA
+�7��;�W��mی.FN����q$c�]�)g,/t��L��"�L啯���Z��`���x|���ؼ��r�fD���F�Ơ�z���=MV
��,��$F1.���������S��}�g<��a���+�P �#41Fn�r���;E�]�ԣ��I�8�FT�wjӗEp2� _��Km`�@\�V�O�X�
v�@��q��aq΍&%��Ϫ�O��0��ƝI� ��	��J�l�����4}/��q�$؍�C��x���^b�q:z�$�K�xiO򁥢�ʛ3Rz2&������mH�x\N�C��8*���b�m���9�+�CHt*R%ԗ�ڀy
��ȅ���K2����?��a�{���x��OC�	�T�g�IC��hs+[��/�}@1����ǜM���}b�ФE$�dz{�G�c!��!��G��'H�]<&�MЕk�)I����#x��"��������v��'y�1w�����H!��\�i:܈��>0�-�����~� �v&�G���,<�
�(���h���٭�3t]N�Ŷ�5B�c@K|w��o���gݗg��ġ'�A~����)y곶�Hk~����utr��A�!�R=�j���l��-ݼ��w1Mv�+��-/�#eZ}x�6��d��� Jo|��A���4�]���İ�FOQYk��e�����h,尷P�='�6�b1�Y
���1q"��:�s�)%{V��I��T�$�R���5�+oc�7�
綌��V=S��k������^/�.R[��:i�w��^��{8Q���]U�����e`�ML���T�����=��Tg��Y���vȫQ���s����dC����y��xc;<)C/�Z�A�]=��_G�@z�������dڟ��|\#���[J솹=���[�����g�����o:�[��پ��'�a}��
�N+Se�=��2iC���0n�H�Q	�����-�,��6�����|��3v�$�[j�a8Q�h�(�i�{��Tx�[R�6����4���뭜>H���c�vUq�h�V�n�c��e���	.����E�Hq����cAPY����C0�|�O��"�>�;k`�*X��˸�KϨ��C���8��Z`���,�<:�����vo�b�(���D��8���bn�nZ�����hwa�}��#g+���7r�7�銧md_�2���'����V�A �M���_���,n�9�]U�Q��3ܟ8z>�L� �{Ϡ6�UqZ�ݸQV���yx�r�pH�l
,�:��<�*� �H%{t#K�Oe6B0n	U(�'Im��_���d�BpK"����$�њ/׾:E|+A����0 =�L�&>�3�������K��_ƪ�x吠9�<���!��5�*Z4��#aIO��S�`T�k��CSg<��j-�06�*�����.Ƹ��O�� �;o-V��W��N��w�lŹ�%`a��-,��n���D/�/ƽ��l����0��YJ��Ỹ�U�a{��^Q"��n;��� ��Bϱ��}��@V:xT���E��&W7��!��w~�6�~�Ȝ��/W�q�i��擜wP��4E�s�����(#W:�h�77���T6[d������i��M���t�WT�.w���/h&{_��J�x��v��Öu�u�y�%�?cÈڇP�7�&�ڿXҪ����1짛�PbY({����`��K:���B�D
L�q���t��ΞF�p�ߋ]�Q�����p��b��a�Ht�Z�����T/�
Oؐ�c�n�������?%ě�1AơB�&��2��iȎ=�ǪB0z���]iuS�cN��\�&�V��� Rj�+i�r�x�Ǫ�V�|\��Z��:n3�!Jǐ�22W&Dw�zٵ�فԙ{��wtfh�M�簀aJ��eN&��'L�\oTF6�q;���n� �s��1�_��/Ls�RH����hG9Y�����Ԋl?	��$�?+XB�i
e	���b�$�����ňԆ��?��IS83��$����ޱ��a�BZl���4=1�$�H��/ ���0�JtULܗOLi�b�U��HV��")��4�6�����Z�׉�������:t#u^�J�-;s']c�n���slx��&\WA��piD�c�?r���6A|K{�B�\7�(["`�1�(���lm�4��&� $|����9�V����"�Gڍ��<����`��EP��ئ/�y�!��]"�w)�|��}�x�:-J��@�+ц��^ёE�v����	0X��F.�=+������~ݲ�D�l��<g�x@4*��y�$���EM^!7�i~��-�*^Y&[<��i^D	l�X��3�K�İ��Xh%'U���M`j���0歺%�iړ��:���T��jІ��KY�~��Z�[�U��H3j?5��ç��DD����@-<�T�.	ی��� ��@׫Bp�q�D$��+e�l�[g��$��&B��Gz:S}�Ѐ�t7E�>KS�����'�����t�51����K��J���}��>aC�Yk�ɵ=F�
.ַ�6�q�|ד�ɵ�yã8
-�ğ��0|�7؇؇U�!��{֓ �?� ��Rr�]i��L��M�:�Q��u�6k���]�7�����8ݡҷ�Z����%�%1���dD����a�n,���HvWM1J����o`���u�|\��Ǎ#{��P;�a��2Q��{���n��NG�������Mwʴʷ��18�_>��u��(��k)�+ی��a����b���R�cc�;����.�4��TG}3E�.�"'Q�rFq��;e��={]p���w� � �i�[-c��5�DD��w���z��G�seC]�����T?��N�̘�MR�k�	��{~�9�x�����^BS+Q_�����2�嬥V~���ƌ<�����٢���o/��4=^#Ќ͓�cQ��%�rkM7(��X3~��$R����$z`�x�ēV�3���?�5��������KI!ak7���آdyN��4=*�y����?ogu���NGO
��)�f��X'i�"��	H5Ȍ3l~�
u3P����ا-��N�8�5
^p�����!JN�����
WP!���}��]��V�@o*W�L�kz�s�B�5U�/���🸕^�w�n�0��P̞꺂�ku�u�|aO#��?�%hB#���l2A��MEn�_�C�e��;���?�\l��Q[�
Bp9.?�焖?T�P5L�+�\
 ��q�N,���'g��y1L?|�X�f�A5Wu)��u1ɡ� ���9��	(�:�'��A��&4�0H�Pj1�*��Ⰳ{�^�g��y�A�(b�z]$��p�T:^�H������[޳�\QuV4���O�Զ����1j��=�'�7��Xh,�z�R7���R�Σ�ap0�(��Mn�*�����̙1�{�����D��B�GV��K�l�:�5v;�D��9_���-L��ֱTe�g��0��S@���Yz�>6uX[zs����SI�S਱��[�(6�E�)I�7w3�^��H�)Cgn���t�d=���jH�V�VI��{���s� ��qV��K9pG��j�	&2@0;�_b��y)#Ӽ��h��\bS%LO��Ո�yζ�e����X����1�Xt�G��?�C�$��m��w&�u�z}M���%2{g�W$�%�$ҧ�����TuJ��k+!�ZQ��=@�!��0|l�$�>5u>��047���i�U��D���E:2�G*�m ��}Cr	ă�G�+�h�[�ud	��
�/tq���`4�L�J�����������(a����O�K�+N��jV�6{&׽�,]��oV��~�Ikp�^�����9Vݞ!P�T�&��[5^H��ͅ�(���fb�0�D���U�bc��r������1��9��/Ho�R�
/�����5�7��� �e���!�,��C��?*qz�h��%�H:D��!��g�Dhqׯ�g���S,OA̕�����i�Z��M4�pڲ�?�u �lzyѤ�+R��B�Dޅϝ	Fa�;t�3/�=E�B���1�-1P2�ےaKUl����/;�*j�, ���d�ջ��|Rkϱ��{d�w۬0��E�F��W�߅������3��&j���xઋ�K���Ϟ���]����}K/����=��r3��m�)��Y��ǨO���D/>�׽n�o��<tb~j�X��.����c~�2��x8�py��^H�оjn'�b�Ρ�I���I�>b�L��v���KS�����eR�H/
�W톛,�2�o�� h��B�ߕ���=��܉�e|P;�?&xR̝�Xv�v�?��D�8�>k�M1wǰ�?���?�1�Ez��\b��3�l����a�H�"�0yX/�G�sb�X�伙�^��
��Mk�N�勵�\+?�8x��,�Lfv��R�&ۥ�������ݵ�g����_�u�?u䲶b>�iM�\R�"��c�<�>ē�X!4�xG"��D��o3��.���0���uZ�s��baT�#kx���k�'ӳW�	��i������� �om!��`� 4Ϫ+���tsC����97�Y���9����?)���tD[Y�N�`��w�$?����:���`��%t7�j�%����<�-I�:����h*3Y�Y��'��?9�������78��^,��-��'�xG���"����&�ih��4,�����$��Y��,��V���D�d�BݦG,v���5'��KWڥP��P� :��y7s���Qk�#v;�W�!,�n����-`!W@���c�Lj����� nLH7?��W17T�7�+�
Y&a��cZ#U��3_c��x;S�����۔$K�����!����=ύo���t4CCm���MZ0C,Y��<Ӓ�U��Qe���Kf��a� �X�1�L�����U����y��ׯc��U;�?��V�a�������lT��!ҹq�/ʨ[]*�6��Vd4�{���i�ݧ�L�L�Z��9�����B����h�eƃ�[�o���?�����,��.nHs8҅��	�u �1OVM�� t��E���[ӃY=))���9��,fj��{����{�|�SJ��g���h9�h=}���ӑ2-���9�?i�O/4�ö3^�Q���k�ԗNrm�?�M಺eFaM�F2-�wt�<����R�`{`J��ӥa��/-�C��l)�$Иor8��"�9,<��s�k��&�	�~H�j��{�FK�,���A���K��ګ?�-�� ��7��dp4����2rm+T��y �.�	,9�p�p�
���\�3��b���zh́e��[�N�ʁ$�2��,�&��6#1��
�@	X/0�D����"�N`�+U-M�v��~�F�60���aPy� q餏�O�F�.St���{�c��lA3h�D��u@$Y�jEi���K\�h��ް+x��]Bb��.���F�`Jr/����r��GIP���)��}KF���>�/VLΣ�޻}d+� �Q�&����H�o�^7 z� �T4[��F��h�CGE�Q|�$z��t_?���D��e�(@�</�� dgnn����ZyײkbP��<PŇ�e|� #���-�_4�Y�
h���!� �yv&�ʑ�=�v���n��a�p�][��n���ޝ����}'L�0c+ԛ��޽���}#8��95� D}$�$�553��j<��~�P����j��5+�X+������[~UP6��1�83� !N�;j���T�ce�����#g�>�+�5z6J)Y۹P�bbjc��,��ͥP��\#M��h��Ud=��Bez�ſ_�?�(t�,)yXVn��;�6I�=�w��i�bǤ�'A����i��F�Z��7pP��n-�8RI$������(���*�1e퟈���g�#��r��i^k��BXO.\�u�4ٻUǹ�t�sO��ޢ�
Hl��i��>7є^K	y4�򠬍ٙ�VagJ'���"����.G��Ӡ�9�����9Q��;����>��ZI� �=d��8��=/eZ���*�R�N��`9{�l^���T��ͪH�+�����9�CP[g/
;a&�&^;�v�=X�EB�I���y�ÕPόB����!�D=��Xb4"4�f��",�hV�)�/��z:�@PA�9�
��E@	�t��a��Uա���`��>!g���\�l5�8����\;��>	�S�ʧ�s�"�G�����Iy��"�8=ZQ��f�iV`67�sg�\� qM��$��ܐ �u�4��.�$���N?y��e�����n�c��M#^��L�� EY_SSkd�?��?�qT��~F���=rI�w,V��y��׳�f��^v��By�=fV�/L���`���K�yAm�m0�Ra���:u��{��J�}���?eZ��8KX�(��gT
�'�v�B8���*֞�-��X����<VZ��w�X����]����ƞv�M�E�зlڰ�Di-B�}�A�T1�)5u�c�(�#��H�?a���s6�N�8hg6fԛ�/{�Z�����׭n�@�§I���d��P}41��TC�%E��k����75�k[��0<���L16�ϩi�a�sR��7O"�\fV�#��.�� �%+H-��\����8�y�����r�0��Ӡ�z���N�1=9��/MV�j�܍�����1#��_f��2d��������_������ʅW�`���9����^���b�SY�i��:$к0�C�7��i��!���pr�|]J3o���Ϧ��/sK�`^^�R�ӪɃ�q��A��w�4fSzt(�1�X��\�qKS'���0�^C�LF�f��)Ί0R���B38Y�ȍg�r]8�0���w�/�,N��t��5&'��F0=ӗ�s`J�.���3��ǩ4�%�ׅH
�pzDѓ�`Ս�� j3%�}GؖZ�6Vb�/lX����xa;L��R�0w���cv������nv�]��v�,���;y��&�@N�}��C�f*�Rת��~9���M�9-������%u�^�Dw�y���X��_	<�q�H���3!���$�4 ҲQ���9�ֈ6_��b�G�6��.�;C��F����`L����Y��ͯ���⟰����~3�W�oR��.�����>�boD(���A�ff��a�2��MJ�lC�SaCM@���|/[�y俈>����W����˗��`��k�H�,6��O!�O`���j#�)+���:��'��DP��]*�E�Q!0�������	�֏o��T��]Rr~����&���WZ����}�X��:�p��&�7���q�$�W�ힽ��Kx`�9ٍ-@��??:H�ޓ[�	@Wj.�ֲ����$?�}f�7�{s�=���Mz����,r>N��D�J~�j�4�y9�{��z`6�N�aقA�m���%���<g%��q��	�(L����;�� gK�6,m��IÕ�6K%�oR�kQdE��if>f0�Y�umŎG0�A�4rY%�w���[#G���-��Y`�p��M �[vq�=S��b]~�/a�����ͫ�~��ƅ@��Jw{��Y��?�+_O$/"�:=�|she�q*G�`�V���բ��(����"V�DZ���~\w,}�s~�����M�3��s���.��_�!�3��v+Y�;��j��'�-�0 =d���*8>�{�X�k�R��ұۘ��R�dWxT���{q���ic%��=%@�6�/��i
9�t�j�6
?�К1
ܖz���JbǨ���1G�����Bǎ�N� &�Dt���6��¤m���QP}����_hŹ����`)q}�3Ρ�n�:�9n��L;���郩儺r�q�Q~l�_Q�lz#�E�O��<�����=r"��Og�Y7�4�d�mf�`��R�įA��
�Gv��D�ՃRh����GT���zTZu¦��WPno��+-h���k��t��2��{ޝ|�@�U[��LL�R���5јoK����Á�t��'[{��J�g�;"�l��/\ f��2���T"g�0�;A<�!��5��П�7;]���R��@�ԅ*�%w-��1�a2�����(sf���X?�4%	\9����j������ơg�s���ɑ�Č��k]��4G���� �k܃ ^���"5(���k����CP}m�{��r�(��
�D�l�#�v	˰A{W)+b-�$\��IO�I���Xi���ɠ~ݕ���Btҥ]�~�3�[��	�����#߅�wCv]�7�@�K�d:r4��~VFy��X���>*ǥ�ӥ�)}����N����C2JA�������J��2�ǟ����O܀࢈�	�}#�����5y��D�-C�R�KpK?�%�l�o�)%,#����j5������O+�o��r��=�ޚl��<0��w&aI��[�CK*�UG��;�X�B<x�j�x/��1H�>v���cs�oT� ���m.����vt��Z���,
�XW����5�kiǃ���C�0�\��O�c�ler��@OA�!�T��i�?G�L4|ӵGF�2��D��>����.��zvu��t��d���Xn�"�9ǅ��/���Lӟ�I�,E=�W�u��se���
_���
�!��^��?����ԥ-[�z�DS�5�.�h	vyI���S���v|P�h�������{������x��5��FL~1�����D[l~�
\�0RX[&��Z-b� @X�P������7�����&r�wLp��L+�/"'������W5���u	0���|�s�$�b
�I����� ą�i#_��[�Fcފ ۸7�X�7��䣤�(V2�!-�2�Ai��?<��8���G@$c���:���O�F�#S��N�GCƤ!�c�O�n;6F�������Y#f8!/�O;�a:L�n/�9=����jVLǨ#ռ�����E3�n]�|r�(Fbt������̤H2��B�gF�!3����n��<hr��H�ޖ���S/@�zB�#��6k����*�Ep0	p��j�3�9kg�~o�n��l��� �-#bh��4s/�^�"q��~��O��65�������^�W�N�s���"����)���0H�����mOvp�����*�E�*aҲb��Ъ$Ї{oW(!�Kpf�)�"�^_?���_T,25� �7�o¶}6��0���}�������`GR�:��g���{�6�v5�
ȌA��-{աc�I�C�YOj��R=m����u^�1F��X���c̉�G��1M?��s�]�9Z���bi��ί��r�'�r���a�	�=V�����y�!�$�ݽ��u������,B�~P�Y�I�k5�{�uz�S��fa�B}j�M�	?�u���E��9և��u��*�*���{	V�we'B�xo7!'d���z�{r�81���(�<EL*!_�𛹹��V�30u)�=�4��B{�Q3�sfg�}�

��������	�`aR�|��75�2{������2��M�ԗm�:LlG4P�9�,��T=={�e� ��1��T��<���4�'Ť�΍�8I�o}ЬY]�JJ�����)m�Jz� N��A�.��Ɔ�H5V7�m�%=�[��"��d@_c���H/ ��yM�$Ӆ�V�6���:㳕u�_ ӱ�/��������J^kE��l��M��)��e��=�}6�}{�C�*4��h�����q��әu�t�Z���3h��g?����Jl1Tk��n=�l}����)��k���B]|0K*�o3�.Ɨ��Z!����~�oW����1P;J^]���f����qKP��Н���i+����J�U��g�C�0����e�<�'����!Dx(�8m��0��@f�����֝N,�8��	���͇�vb�M�?��a���QW�AS-�ؽ�ȏԂ��Q��њ�E�1����?�VU�ewf��ԆVe�5o�{t�X�F��
��N̔����Gў����<�NK��ӿNf��T��g�i�췐Z��VfBrh�e��ƪdX#���G���-�z�-�)Q��9:E�U�"���1�}��?�g�zHMvۀvW��`��\vK�R2�2J�
�YҴ�>A�Ĉ{�����KI����a�*�[��9�3�'4�!ᕵ�f+!>��ً��z!p��${.�̐��:������Ӿި���@�l�Hf��a���+�u&(I��荍hb����=#�R0CL��SQ�5*g�:��
����g���J�I��GY,�XGFH��Ee1����3�	�E�=��I6e�=����^���DZ<>DW��-����z��dN��p}��g3��=Q0�V<�;\5��_���X�mW�L�9^"ͩ9H�g�:YaЯ����[�qM�#n����*�{�9��$\d�r�
�\��_�r������/(w����U����ye�/
���*�m|`�Y�S0�*��c�|�������N��P��IR_����9ov�Y	�jȈ)�$l:�W��mm���&k�c?�a`�y�=0�)���,��_� �d���T,�/u����6�{ک� Μ���1����1�8�ȞW�@�&�X;q�6Z�T���kA��c��������D.Y�E�p|�[T��;d�e9x�;]��%O��n����֝�ζ}X�Ө�倿WБ.��i��*>�Mn.�pW�>q����6�fOF�u��`�(&5^H�0�K5���F��a�
�gu�`�?Q����ys�#��Fs���5z�-_���1������S��Ϟ��/�dV�'U�B!#�߈6� �%�X�\J���pFo�L(<zǒq�9�J��C��{ �#<�ZcȈ�Oyo?5%�Qo�T4*��i���Ke���r�7-��/o�Qk�&��m������@�Q�
��Mom���F�%�d̺�4J�EY��˿��jW�&b�;�W6�c��A �����U����/�㗬��\`V������k��w�M�A��
�̿y0:������ԓ
H.��&U��Д�N��+vP�r^��V{�9��h�~IW���|RX��$�j�8�`�iVu\��՚$���ҏ�?}LB��桀9O��- ��		xR�
=�S(\>����!sx�����Rg�-��Q�Ѣ9�*1@��(���0�QPB��`j��(���ϳ���F벒e��Q3��@ �c���O��s��~���jq�,�f������?�J �;Y��F�bm����� ќX��)]�UB�����PFi-̹%���6�΍:�r!�l�	ORln^���=��Iї&��RF8����=5�,�4��T8�����ǝ��{�ꮥ�ГJІ�+���V�mfOA�Uv�����~F�us3ໟ>��>�8��
��+�[\E�T-����|g!�hi�f��W�g����}��|[x���ie��>��P�Rۓ��`hW���ݼ��3Z>�[������%�3�ʹ�3���*Ey��(�����k<e�]+��7-�c$��k���w�u�Z�ȇ�r���jd��MQ�VkOL<HF�}��=�bs�è�X`��K�_
�|��﯐J,a��_��g���G:P�C2L	��s2���)�v�1 (ґm_�>���>[p^�U(�p8g�ucI�Y�̞��=��f��M)<�,2+Qӵ�"~��.����M�N��81v��	6���tj	w�ֺ-Q�k�@�@��p_�\�A�W���21Hc�,��#I ������FY{�h������?���,��p���hc�!k�c\"U��`�\��7�9�d����t�>�q��ꈇ�t������2:�
�NRNu�n���N�T�t��Y�Eͦ�ك4����ۊ��#��{�s@�4�����e?d��O$�6{\$9�_��I5�Eh[ż6sg@�3-��?����p�f#Cs��GK4�]�����ǘ\?�n\LD$Ez��{�բg�ў����cI5K��� i��t�v��뵎�&BĽ2��c*꯵+���
CB[cU���cCA�d�ʔ��9�x�I�q����'���-pcā�v1?
I6�p^���]-Lf<�!'���d%��qU �l�d�#O*k9��al����';��� -���2�M#K��E6�: �d<h_5+��gFڛ[*X�QC��j)�^K��;�)Q�k��<��c�]4�	u�Pq҂�.����	(z�=�t�9@f���5��������K��"�^��L������5��FfKjt,�?�R��߻[WA��%��d��?b�m�P�=�*�{�Z�V�oi@<s�A��� q�4��nF��a�<|�cq�f����ZG���>1�>�+p�Xv!�j�B)iIʱ,(���7=s�>򷨠s�(�^�s1���^�jQ����X���Q�����X.�c�^�i��i
!�k�}DmV�obc�qҋ����-Īz�� dl�G� �/�=0"E=$k�o�j�G!�ғ/c�܁vZ�S�+�J�v�з���<�,��x<4��s圼7�9g���մ�%�Hq���L��ߢ)�[}�І1�u�V��j�RDj������O�e�eI ��������)�@Gn����LS� :E$���~��tS�=M\#��}�j�C�^��H���IWz	����Q��v�(�!W�-���|���D�����W ��&Շ���	������:cq�h��Վ\��-���p�H�&�l�5������%-J��-y�À�~d9�{�	k%dd�C2{�ttj�ږD��oD�بQC�$�c���>���*��`v��������x�R�-�cx�j@q��!��W���4R� U�FP��A��K��¸}���(��"�(��x�gF��k����J�@@��U=<���;��תWq� ��]����ϚqVE2L���ƱםG  �Q餼��p]@��`|��͵�I��p(�[U�
ir�X�>-��D�+r�L}twVyv"J.����w�G��v�&#ƿ���잋M�����/����p�ы�x0�F!��d���`kD�.\1~�䓠c2�P��y��O�?�hDC�P�Ƅ@8�#~��t��w^j��R��?��]/�\h���g{�`��I��)��咾�I���{n1y+��ny�6K#�|t���lT/;�t�(=~���7�lF��ݙr��%�G6AX]ο�����.��%I{�tT��gϪ�r&o3�������Ч��<h0ys�%2��RcNc�O[�%(��g�KJ�Ӱ�.ydh��|��,�����ђ���=e�i��ԱE����%���0ZV�
W��hҧcsr�K�i(�x���p��q��BG�: �����8����V,P�@D1���2���4�п��$C��?�������K��H�l}�~y��ģ׀mL��!���)ZD̜m���U�����OJ�XP���P�+�<{;^p���iHY�{o����ǐ/,۽�����P�$&+W=��j
�-Ea1��5a��5�+�B:>�:4��C'�Sy0��d��b���=`�����o�5����o  ��Y���& �6����HCX�����ԋ�!8�]�_��Y�]V@����㻩�&υ����MWV�dP% �ģ�Tp��b�����N�z<���-�&��X�:�Bi�h�����>�߉\��u�Nf���0��%B/��#�+2W���50�/Yг��8�����������]A�*>�	�W���*f�v�x�����޸��m�L�u�\ ����}�o��)����&öL@8�_R	�!���4 AB��!��_p{N዇��&/�>���GK#P�<7���'Q��eC��G�(}�w_����^�������^�?n>�����(���%�S�ݾz-W��0C��G�}(^H5
qL���T�_}��G%#$�j��5��7�Fw&]�2��BhD�v}I�Jz���W��r%�n|$�h�,4av�Ø��t;�eTL��{ǀ��7n0O�d9a���;^d���]��w��/����s�r;{���/��~@'�7���H8�6}����l���||���2��r�ufj���?
6�J#������,&�0&������l;�I�����Ӡm/N
ʣ@;:��H�|EpƢ�o�
�jȕ#ǵ�T������u� �6�LRAz�sq�ۍ�6��Ȣ(n�cl�Cg�kL'�Rbv�U��@N��tnƢ78}� 37�z��BD�p�ALh��b�uV4�V�$���(�C#*+��l��h�JR�z�Pa��~}��sF��ɣ5J�s;3���uЯ���<��(Q�x��+R�G� ��"L��5=�B[y��\Ɔz�Z���2Z�v���]�.m��VI�]{D+��j���v�&��>K�w��?��!����E�Q��`%�͆R�<��E���K#s�vA�̀:-íeC�O�`�,U�E���U�b���Q��ɝ���[J��s��8��G��\sVn� ب-`��#�KI&�a�u�?x�0O9�(�,�I�5\�6�m�R<B+Ҵ�7����c�>��ɯʣ��ڰol0���S�I�#lR`�MȃZ�͸ʕ�`�0)�măD���%�h���0��Agb�|KigX�OÜU�*!+"�lU������5ʇ�K^qم��M�<*H�T��9�����?N�x�`�	�hg��'�J w�#�GU�q }V9b��7�D��j2Rъ�)q8s�F���u���WBE�L�e9S#	�M���HC���1���d��R��ڙN�1Tǚ�p����[�5��#�� ���x�[4{#'���&�0�+H����)�~�K���\���0;�߳6��d\̾�QG�*������ϲ���C6k����h� ]{�����A���×0r
O�����b��)��:����QR$9�[�~�?���nT{bM���P��`8B^Йd������f���e�}K�I@M���Y�Ww��I�-�U�*�+�6i������Kg��k��!�k��nN|wh	�����?	"rx���bPЙ��9\���a	L�fȤQĞ-ۦOH�3�s:�8Lp2�K�:��\4t��t�,����4q���q��GI��>sl>��yH�_�"#�+�3��Z��@�R�F�8SX(�P+Ku�z��>�-��+0ާ�7?NJ������Cn��J<��@
ƅ_|�Fԩ&�1o(�TF������C	���XFXȱ���6w/��_?��I��N�S���Z�]<�2e�&��vs&e���Qq7z�5�j�?��L1[Be6�P�+N�<v�͛	6[k̸<_9w�֩�Fi�O��D_�s	?�#�����H�A�EX��m��з.u�Dk�.ml��:�8e�;�Q[J�k�[d��[w%ރQC[�[n�I~4�$��ע���T�v� �[p8��*6��磎ƭq��9��%7ěX�Ӄ+q|���y�a��lF_E�	�(�g�p���qQwd���YBte!�R��v�Dq��7%��p	��y�bo��X�7��d�E�{I,���'�t�$Z�lt\悓�"3WR����z�ʻ)�ē�a���1�Z[N'��� �g1V���X:H�a)�^O���kgk�F׳��vR)�n	�1ھ�!�t��c��ʅ>�3,��6��!!�5��
9�j�T���w����Y�� �e�SS<���K��z�䲋�)���tr�����s�ƃ�T�g	��H�æ�P���16��_a5��L��~��jX�G�����'�D��s���"�#�S���2�![GB��z�/��I�8I�E�3�'cl+ZӉ��NY�:"ͩ�|W�$�dY]+��|�2�¡�16?�Ƕ˪�0��-����e"�r�+�x�����3r"K�W؇�U'�}l���jN�����I�{�:��ӊD��I�����o<P�f���x$�V�Uȷt�Y�;��Q"Cc��J�@��c�i�)��5,ƿ3�Ih���9������ka[�%�AG�3Xjk�Œ^*�\��*���uE
�Λ���*B��*�h�o�*LwMrdgu����Ӛ&���
����N�HȔ{>j�z�:UT�!�6s'::�
|E�ei�k�﷒M֝���Lk�o�x�x�����!��))6��%t���/�<f4UI�4/�M���,H|�O�=����/M2�T��\�'���]�j�'�H�}�;t����0�"Ӡw$1��4�K�Fv��"C�_Wf�-��C�y�%�zm�&�����z蝗�S�V�[V.��@�h C�+�4厑�����x��r��KdPF>�c���	59ee7l!��󸆏ldD�2�x*��[M����%����M��<�T����дY�G��l��L�Lş�,�}�N� ~ �x�����i�����i�O��m�0t5g�u$��r�X6�혖�kBUBRu��j4H�<^{�|x����]��U��X�b+¦�`�2q��	�{�S%���V��*�n�̱���\�YB���EĦJ�T��(��{l��>�湘��������Dh�?���Mp�T��e2D�D�<ʖ��	�t*����58�����K�ք�Ԝ�a�C�"6�,�μ��Vɠ�Ƴ�22ꑗ�'��pXI�I��p�y�$�y�.��4c)#^���΂��Ѣ���+'�uLo���hL=3�L�j' z���z����t~���Pg}�����gRK-s� �y�e��Y(��ry�� ��%~�6�8^}�U�x8���m)=�����/%���E�a
�_�n�?�敮H��{��y]@a8/h�o�Ӛ�0L���8̧��d.��Ob�Eb6�$!$&�ꢉĈ2���!3�f�WM2f��k�8�Q��f��>^�w�Ft����6��H�JL��s�u̫ѳ���� ��8Ec ��I�p�c�ܾ��B%h��W�k�bO.t�򕳗\-k���3��O��KyT�������9rO�*�g���"pQv���Aj��Se��5[�;�}�+0|�Z�9�7d������y�����c���e�Su���~x���oE%�����ea�[����T.�k�"��E�;��9��v���5k� �d�\����L�[\c���+�Aʼ	�I��W��j�=�%��k8����|:Ul�s�]��o
�,�å����J�{CB
7�c|����<D=�W;t*���w(��¥	"WaD��J[\��k��٬z>y�T&��<��Y�o���4�,���Uq|�~���BB����k����]���?�D\�ů�	����_�gE�I���*y�d�����e�9�s��e�R�8�dM�ݺVA��oS?�\^+�D�,��{!m��>��d���m~���b�n�(�]e=g/�T�aV� &�@I
���x�j�goy=l*�N��l�%n�����YouIOZݟ��b�am���c�����zXN�t��#�_lbh�
r���A^�������x�k��G4����S���Dgg"�O4w=���M�$��e �����R��sg�y�:�[ԩ���m���M�P�����6����B9��q�@ߚن���e(�A��1��w�����Ƌ�Fp*��ww�C�o����c���	l�mr���$�-$��4====��U怗�{���E�Q�J�cG,�k�_r��(����j���m�}���DV�v��m�b�#�R"���q2˩��hV����K���Ԧ��-W+/&��h|C��K/Io��_��'��a"{g����^I�� s�����֊��%O��bd˱8�ےR�B4J:ĩT�ٳ""|z�0%�x����ʘ��F`?��ac��'�[d���dCPf��"T�x�� "�;�.���ڲT�D�nv��D���'(pE#��4u^�]���,�*�ፐx�Ԋ̧"y�tE�2�H�NY͒��ON�\Ȱ�u!����A{Ƭ��"I�-z�ݛR눮[`�a�{Yڢ���Tꈄ�JJ�&/!�x� �넺�X�����3�G���߶7��y4���&w�nK��ַ��E꾅������*43_I|�~b��Pُ�d�t�.Z�W' �O1�9���6��k���O�k�r���EGN8�hf���ޤ���)��U��ݔp(%QNP�.j|�d4r��$��%*��+c1�G rNvʥ������$�nЗҺ���� ��O��ZL�}���Lm�0�i0�w[��/"ӋUP�|�s�Hqm��ס.ar?N����B��BnF�iC�|��d&�-<	�3�5�Gl�&�p[Z�ǌ�����}�ѷw��G��!�Z^e��U�Ek�.@�t��P��ʊ
���$~A�7��
FAC|�_���E��`��k.�,/R[�W�>k����Wd�#����3|��)��@�H=�:��%<�P�5�tS���`�0�=�gqG �C��Wbxmji�zV�ߠ��:=��Y
B�����M�*u~��� ��uL�K��	O� ���]Hh8���2F���^h��,,
���D��;���<MT;� N�C��2 `v.Y%��C��d�ǅ`ݡ�P\F���"�r�?Ub���#�̯���(�r)pI��2�I+�.L/�a�����M/�^_�N�t�1����Q�T��]ATt������u��� �A�]:��&��y�h�0�1�&5a$��H�]1enwtP�Ȯ��<ҍ�(
k���e6��G3�̓W2Y�E�T�uÑ{�.���:���屾1��CKR3Y��Ke�խAٗ]��$�v{�P�|	�H���>��&��ͨj�:��gD�e����2+q�84r��+�ӿ�hb�B���	�[",W�jº�i|$��+H�?���	��<c�1t���n�f�F� ^�̰(��F_F��W6=�c�|P t��뙢H̎��#��)�:Z��*�c�\'�fk]h�nF���Bn특�F�������136�Wʑ�
W���0�	M�/o�GS���g$H���L���QXA[Hȷ&�o~�T�'	l�(�c[@�)'#]	)֤�C������o��>��-���0t]��z���,�&��v����02���S͂c+ pÎ�
�'xv�����C�}fwv�x�|�8j�����)IČ�^Q3T������Rn5x(\��R j0j��mx�<��h8'����z��lW�j�	�'W٦��{�m��!b4.�"�_���R���{�Έ;,�6@tq,+�����1�s�W
}��0OG̐p�%G\��F! %�Q�l7;j���d-�P���`3O��(X��#z��lt#��P?���%�
��Zug�HsY�v�^�f��zeɆ�r6��'�Z�v�h�{:x���+P�E��.��J�%\f#Y\��+t��R�*����L���r�I�S�DO����T�|�Ns��P�Q��7���{���*��q�.���1e,rf�46!� ���~�^���!�K_wR5��{6��#�,�(��:8����\&/���Ah��n��>k"�<V�Mx �"��{�$N�b�7��d�&�7������!s���p ���$7��è9�4�t'vgߐ����4����oi��nI����R#���*�E'z!��\ԁ䶋���݄8�}�h$��Ԗ�r���:�O�ل#�D�tA��E�Y��Ĉ����eH//J���"K�C��v�I��陙. }��&P��r"�&d`n4<����R(Ƚ�Ύ�L�����+~���SF�����E�s�s�%Q�Ya�ʥ���B�E�m��n�~<��UV�?��l�!�'�����E�?VN�o��N���kG�#�CԒ;m���<�V`<����f=�'�=(Sˆ����Ru��ֲ�W�� �m�j�}l�(�:�C.F��"��i@�c�K���Σ����C2�����yF�Fk2gň�΍�\��ΑYz����(}w���C��a���?���Z���Zv'�e@M��!+�"�a ���Z��!*4��{F���i�V�LN�?{��S�`�߉�y���nTX7���Ş��̗�?��g�u��݉���H��.��Z�W�R][{� �=0p�49opg�Ӻ��]���ca��v�~Xzܗ�[ǠQ�Ƀ��)�FUl೥�Ka�A��~�Ps=�E'cy	���o	!�L4%A���:���-���#�7��(*Y�}���p�޻^�Zp���|)&���S��]�� ��^ؘB�z7(�'��"� ���-*�I!�{��+4J�n���'��G���d��&-9���DP�0��0�����u��J<���#m���I����*�8�k�q�񶄇�-$*�(�� �-���u��ﺮ��NQpu����ZQa�I�����(Z��a$xv>�ƈ	Q��Ġ��e��7�5���U @�Z�H٫�"�{Ӷ��#@�-v�~��b��]L���m'������Q1,&�3��C(��5�$1��K}��5̸êU�H�����V�kH��}���J�Ź?͔��B��{ޏǄ���Ќ���D����y�LX=B�䏂E���`��e1T1 g�Ӊ&��A��T�>ߩ#x��Sx�F��D���{٧ &��mr\�b�a F��1��7or�������:I�zn�<�&˹ͼ�OߏJ�����5В�ߑ��-���22�����]2��6i�O�6N
g�R�32���<�R�� i����*��3����9���Ө��#�B2�*���M~�U�랼���dF��aڿ� �UeO�&�p,б,�q���r���䟵^�p1�Ga��	���{���|��Q���\)V	G-���R��lF��M'ZT�3�
2uڀ)KE�B�R]�0�pY�@a���"����*
#���t� �V=ʃ0�Y��j�7W�W�DG��^`f"���U��'��������I����XoW[�N!s>�ŀ�e�ڭj��L���>9h�PK5�J�w��)X��h���"��p���<DA�Ī)�{~��@W��Lj����V�PX���.�Bouu��e0��@���lC�0B"����ᶤ%�~n�I *�E�������O}Y�/��*z�Z��쏚:-���[�ι]7YZCx{�d��C�hZg�F�T�Cӟ���}/�J�F��窻q���t�+m��QFIX�D��+��{]�4����r2ZL��S���}�Qd�H�uPt�k�tw��7%�oR��}@
���f'�����Xv<��g彭��)�m����N��1܎5⥈`*�-�"�	Kw"�E�B 	K&����F>OH����|e�w�?�-�
�J�"��:?�h�}�ő:%V�i^F~��ZhN�U�Q��+���!`����nxE
���>K5�蓴;S���c6��+�E;i�_L\H��?Pi����l7�5���yz��B�¨�#� �	�?l�5z�Y0l�,єG'�	� 86��5�V	�r��`��FCO���p��))��{{^7�'��?�z�q2�j���k&�����p���=p\M�׷��Ѣ�N%�	9 up��rHيgϪm���΅Qd�k�U�R���JxˀFA�)�g�Z"�C:�XAW�P�|Bk��S8��BVK'��Bn,��2AI*s����:D���H8��?��J���)� U2r�:֏m��G,�o�uhЍ��&�8p�T>��u�����ʀ�:�SQ[z�+��~T�G�ω�4�9%���o��&:S�u�0��Z�F?�V�K~	�<:�Y�������,�Z�ZԻxIR�%>����dny�G˨���5
����#g=�G_ m撚K�?��O����ʴ2���kmM��=`p[�i7�|�Vh�PcF���U3���8Ƭ�����BM���|p&��V�T�B/x�,p�	y*���8G;�Dz�x]a�Sb�8�W.����\)ݗ-�7���eC� �S���هm�c$J�89��V��9�DN7���h�؂f=�E�e�+��s����� ��P�0���>�,��
���-zښ�����=̈�E��(l�9���:�c8���0@$��擸ex� �����84!��NVL�H�3�1�v?u!���*]�`�t�%�Q�>�XhH	J���0/fRd�L�u�����f៓@@�otZ���v��va"������1����t�*X G��vֈ����x�u��m�&;-?aG�"[��}Ax�s���(^���_Cs/����l�X��&9M,�%���!��>Q�%z'`�bz9�YK�ӓe���	v�����8`4�6�z�s����aZl��NRk��t�Rue���g̈��MQ�����`��	e��J���B� ճ�-,����Ǳ�poj
Z�e�˔��Z>o{���� ��IZ'v��S�D��|�(�ِH��K;��cr��Ms���In&V(k�����87!%���D�o[�_7PP��G�!x�F��Ӓ�<�\�*~�ñD�`� �����hct$�Ĥ����4��,0s;�VwP�����~�3��Y��[Z	c�OY����c��SG|J���)0�Y� �իe3��IS�d�!��#r-���p�Xp�gʳ�2!�S�`��f�;)�x�fB,p�+ �ߺq$�`n�D���T��=HM�pfS���x��+�����/�� ��Yʦ���<�iq~y����Jt 9Qe\�J��_v��[�1�9���DHE�fz��O�%�|o�v�1�`��5A{��q�H@�£���]�][}��ٽɵ/2��<��$�v>-��pP{�w��Ӎ��Ө�HDt�A��E���Wa���0�}҇\���a���N����O^> N[���σp����V�[����I���u��D�����:Q���ʩc����ȹAÕ�*U������J�6v��%��1
ǩW�?XPH�<�ao��dt'��G��wd�&;*l���l�/�������F�<�ڻ�[�:"��ڳ4�87ۋ[���(Y�u>�`_5�W9����d&���dr�K�اt�ॽE�dh��'��.c�y�����'��jy/�����Wn���:H�9#8�ܥ�3�=�"B���q��}����A��g�Z�0I;$�̾;�*�r����]���{%�MFm����h�CԳ+�rW�U�s*GQ��Y���9?�QFve�;Ee��!��?J���;V�{d7�����MİU����Pׅ4�)