��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	u������뽞4=u~��l��v2'��0yb�%���n�ot�c9f�na>"Y�~N'�Pzר
܂X�B
����v��y蓈��ү{�>�U�z��g7���%��z�.��$E9b�As*N���lσT��*��1�x�b�B�_����s�Qk���E�: +�v�	R�@v�1�+�^��f?���v���!|6Ԗ��[8
�I�p6y�h�Ҡ�<�Qz��,���]xC�^Y�g1]�T����5=j]+}o�N����Y��,��K �&�8PZ��:�k�Z�Z2n�&��]�"??�u�� �m���HJ����c�t5���|�f [�)!m��l>;b��ɭ�Q�Y��LQ�n�7�ј�;7J˽�ٺ�m�Pޖ{�P���� �R�w5��6ߐ��\^Vlu�t�Mi�[���%D��7�C�AT]��o�s���*̟���7"9<����X��_H9[�A����~����.d6��%!3>��/[�2��e����(���D���G��A+1�YH �7�߭J�n�� �[�Q�[�"KX����'9�'�f�p��)A��S��(l�P�w 5�9@����}Pf᳧��X���b]��������:׈��Ev�����P�:��}����a7�X	�c���wR�Lu3��!�^ �	CJ��v���0�S�ɦV�z>�hGNゼ�ۖu�%���p(�x�@�R�]I�v����dFs�/[���l���a���2ɣ9��5��H��㕏���:<��������� ����@��"����Y+R�@��q�=RX�	�w��˥(d��v�g(�49N�N��^�* V_���^_�/{�r�葐��J��%��~��+��g��T�@_cƠ�ֽ�+B��@�=z�b��y�Q�I�\�[b�`_�v��
&��"��P�>�����Ԗ�D�hH�����2�J�C]�KA��[��F:�E��+_�;�+���+�)�.eAh@/F"���"@����<��1Ar��M)Z�����~a�I�MG}��l�T,�*�QHny�4��6z-�2��3�g�ܧq��@y�#<(S1B7�;� �x0��zϟٯ.A�f��"V�K��"�Ru�@j��])����D��DBF�� Ȕ�G�l$��]z-��\�iU��gXMV�5�lu��+^�q��#t����@3�)K���P������P�@��s:�5�R$�L��� �5�3���]*g��_ ;40.�WbG+Aq��q9y>[j��*iL�jU�B���c�5��J~WW��/6OVq,!��P�Ӊ@V�����X���X�n���w��U�N�}o��}a�3J@� ;�S�y�`�X�$G������ �E�p��;��X�b��6�$�\+�lA`�l�34qu�~"�p��vx����mE��WS=+�Ӳ���kF���k�^�9L�w;���?�KyZ�7�n��e���� w���Ȅ�M�L�<
ل��-B'gM)ߜy��E���\&��}?���5X�k�hi�g�����di>Յ�k��~�ܰ<�n e��%�?����T�o!3]
� @��Ȥ^��i7cC���K�A��<���Q��,U��Ee��yq���H+�.{��ޢ0UOYT6��J���
'D��==ўɬ�Z��v.-���>��^�6n�lN`�dy
s�U�����DE��}<�Q�f�{�\þ�k&{��(��}"^����v>m����,�B�n]m����}�^�U�az��Z}���Bbq<�m��^���k�DWm�ʋ�B��~��ӕ؜gi��s��95|���D�:1l{Ar2(U���𧆄�1��V�7��e��j��n'q��+G\�䞲sV��_ �Z!*;���)N��<���M�׀+v�`xql(M��wfP� ��G(�vO����\4��ދ�'�Oo������c ���LZR�blꎿ���(fy%a�d,aT���� 5{z_���W�Rԩ=v*��~��2�av��JN����V�q�G6ǿ6���\������s��Y���B��N��X���z�l�g��VAjմ��~�g����K  ���������Ǥ��l�ڮ�����=܂,>��Ɂc�z���n	8`�_��|A蕬�]ߋ�=Qz�ou��2_�Z��;T��y� %�S�����o0�I�B{T��)���Dp���t݉uE9�gh�� ��Ikꐸ������qk¢�[9d�_���[ŕ]_Fu�`mt�Ы[n���1���V�ŭ�*�[����H	��`Q�4�D(� j*!�0�-6S���0��d+H�9T+$?}OKĔz9�m�W����]����8曵బa&����"|8�Ux���a��Ioa6��~�i<2�P��*)��6�����_�J�h5)��y������G�y*%�(9z�f�b�B�SJ����v�Q}�sX�hF���1��� ���*�	��W՛σ��O�-A��;TK�H���"��D'�zH������%F�$R�8][��},�!v��A���oV�L�i­g�(7��mu�OL�]}�G%q��-�6�������Q^h�<32o��,\u,BIV�t{`�K���ت��?�(K|�jkaǪ,�[��V�n���U��d�'6��yhC*rhQ�+	�?���D���5��e���J���y�7t�ɬ�K�Ͼѝ@�iwyMͭ��rOV]��F6#����p���>��EJ���@�l��K�=a�OOq�f��{v��Y��@�@5�9�*�*�
�wx��[�������3��T� �B�G�{�2.�@�϶�X�?.d9.�G���4�N3���΂����G��1����i���AE�E��ڧ�fu����=	�K��۫��+�:NK��	Zn֔���#��2,P��I<� �"�ϑb�넒��q
��t��[�S:�g��>�2IVH��_�^���Q�k�<��l�"�##͍�%���鯱�=����9�m�gc���X��Z�x.�b-](���b<�k_��X�f܉ǚ����5_�j��c0����X�emY���b��[*v�,l@�ή,Y��IFe�u#}�͗�Yҝ�^��'�e�d4�~ȓZ�x��ң�4��X��Ւ�v�;7��w�N���%\i+)SKL���h��D��]9�"�V-{`��O(�{,��5��U���:�L�D�i�L�g�{u�.|�͔�Y�5ڤO�f��\��.�#Gߐ$4���R2������aHr���LU!H��b�i7����<�Q�J4{��_�ޥ�]�9�O�H����F*{����Jq�Փ����Ԩ��E����~Ў�7-�.l3@q<آ��c�Ԫ�%o��h�Ff7��?sk6�H|��t�|N�������-5H���o#���JKў�3�4�~\V�8'���{9QP�����Ϧ� oM������4n�4֏)���B�X�#s�}l���B�O�c,��f�%���Ԫ��KBNǇ=��N���f�{/M%G�~�0��{���(`��������d]����iB��,�ϊo?u��<w=�vY\Ҭ�j���i:�� ��w]�i���U4"�H);/��Ij���+�0@g�^�T�ܡ ��Qm=ubCu����pU6DTB�"-K0��(��n�Fp���d(�=��W�O�g[����moJ�j(���r�B�.J"W�)�$m�+�+��;T�X�9�v�t�0_V�W���l!b�K,a�h\��NYݡyo5��U�KMp����J��?8�ߢG����oe��2�=��fA{���<�Z�5�-����_D��X�t^Ґ!m��͜�:�yt���~�eʜ$ܟn���&툸���.�6&,��21���p�V,�y�v�%*|>l�tV������o��Ʈ?�| �*~�d�e/Q����ƕoI�ՁXF�]G�������ģq��5mtf�~�an==^�����)õ��6��~�D�T���)�5z�s6���K����p3e[����|��O6�y �&��1�A@b	���?R���po�*=���q�-;�૧�,S�~�C��M�-�w�l����e���H���arf��矾��V@�8`��z���6�L�ZCk@��#;�Eh�1O5�D���F4�m��X�v�jVn-���.1����+[{�eB�_by�K�?'A#�s�ʃ|o�_��ﾷ�l�I!�Z	?rd ����	8�@��İ|���nWF	��1P���
j��b�.�I�(�|����.���8����˰е�}���+xQ�����<'���Z� B/�4ki��uɣ������l�)�7*����-͏4�ޚ�LB5�d���Ԩ׬� �K����eI�Y�t��ͻڮ�U�M����Д�8[�^��;��JF�6?����)�e�6�v�ͫǁ_"��D��w������D��XS���<il���)u�������Eo<8�K�� 3zG�S�s�2, ��^���[�]���6Z���3"F���$U��7�Rt���n&�Q�_1�"����U[Fy�o��!s���B�|5� �ϻI" �c=G�l5�T�"�Z.m,}$Ry�Mb�+��`������� ����W~c�-9�c��.�MJ����@l�}��L�GO`eZ%Pɰ��4*Ľ����Y��^7*[��-���5q�I��U�<j@���q��3���xz�[�=�1L��D�j)-���E�E�RM�ɺYW2`��w����k�t"�8���mn������-z`��/��lrެ�5�B}�J����1S��}��Y���9�5��-Pa/7�h�gm�YeL'h��l�veȔ�M��9�D�5͵�kl�UK^�|_�qr�y���A�{rw%}����[{	I�5��!���ƅ�:�y:�;ب��Az/p�&Q���-nM�R��\u%k��~VP�n#��%��� Y=kC@���y�*Sy�ґ�DB��t�Gsg���Vp��1�����z~�� �}n⣧o'�7���}�Z#<W���C��#ۤJ����fG��ڰ,>g�����X�8�Qq��f�YjJ$t�Ӳ�
������k����V��e)f9XL�^8=lѠZ���:�v�*�$&e]t�ƭ�}��=#�IL�|��ܕ�'h��`�c�IP�����)�^ط}����&}���JS.�������*ܮ��s�:*��j�v������-�����:e�
���h7�,���v�Et��a|���%�A���X��Sr�1r�S����śu'�J�e�?�������y��0�-��<���)�A�6.9;�=��5��?Gz��Й���� �����h�?�x�Q��h3��4���K�;�~������Z��������ڝf7DJ�.�u{�@('���x-C@J?���>s�e�����q� 8��������kZ�B���(!�ȏ0v��a�X�Cl0�=��S��E�;�����a`6(�
�BLhU�e�${C��f\�5��$�@s0f�����+W��e��	6Tƀ�g�������M��Ic���f�d����]Hq@�1ڱ���٦�=4��/��x*����8���rO<�e|vR��`�x�w��͆~��Y]Yȏ�����%Ԝ�V�ɔƺ�R�ēR��#UL�v=�� g(lJ�I4.@��c�l�RR���lo7na�7�h��-����CĶf=Tu�>L�U�+kg�����I���כ�3%s�Ϧ�[}�����N���C������j$( d���{�R�Iz e����xb�]�v"���2:]+x��m��o"[?拧�