��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl�Y�
_-�E�V�R�]�� �V�]!�A�z��5�)jx�NA��g���i�U�a��P��
�d��x��/X�*�]ഩ�-��s����]����_Ÿ���#�/<��:?D�J�|��2��&Hėm��m�6���H��81���Q��1�y��o��@x�Ѣ��< C�f��4z���!hi�Q+�U�NȘ����2N�OKy�xH�v���3�y��%ĸ�T�Ι��:��2�y��Y�"��p�w����ڨykZ]�R7e��k�窪@�A����`5e�T��Z��{h�6��~+��B$���a�:�����A�>�A^��q��.&�w㰉�^�"�i��h��q17܎'{=�t��U�U'xk-�^}B����2���uCkX��C(,Nea��2�28q����Wn�{.�C5&@p�����zq��q��f,*�+���Z<�%-9�;��~u$n�/��9#�V(�wC| o�X�~w>�g_�?�aUs�ؐ*����n ����0����Ơ<��8-he�FrZ�K�V�ӹ&\S2��(�y`����>~-3��C�\+P�;j�+L���%�9�c��S ͭ1�(	��4{���*���OQ1�5DU�+���_t��[;�	�,Y�F�|�8� �;k:����@��.,�+G�nm>}N|�(���=�O�t����E)��f���g=�[��v��K8��W�b~9�JC�|�N���5Ǻ�uZ��׺��K(4��PX_�T�[��_����5R���q�H��WB�J�x�E��q���6>��fр�pJI�HկN!�$�*!�M�t���䟪@�A���(n��9����C�2��0:����<���px�/nIP�1��V�pIY�o�*l��L%���0|_N+��r�.��M��5�m�W/hn�A��1ہ�������|�.��	G�]�ʸYP�҄��,�ȾoU5���&��;�W)]���$��ϔ���;��M��H�T�Ë��t�����l�?ga��5d�fZ!�d��Z/�ը�RZ�]���Xr��i��7y2�hw���V��yk׍�.����2�<%����IQ����3F���N �p8<�A��������i��v��R��3��?� >�Q��_��B�Xnxt���:�4�"m=>4'2�9�
A.�K�|�.�O��DPe���/���4�o�Ȝ��<���|W�f�ޜ�U6�o�B7j��;	x&\�A�N����E�U6y&q���'��O�� ���T�b5եĊ�6�9j.9���/T
��BƷ�w�P�[�cq��PK�`fQ׷��Q��� ��{���|�}�t�Na�)���!h,��.��!�j}~b�\R�$��Ɠ��Մ�̅J�U5����qPU}8q$����$z��EsF�Z*�G:A��j��ft����.�_�������G�i}������$)N�2�A@7ud��uO!چ���(!�u"
!f�֨,�~?w9��\�5�[z��9_�����4�$��a�RsuHyւ�@��}%6��x����k�Q����<�B��{�S�)������|n�5��]ev�5I����Bݴ8)][�\I~�3�k(��*V��(\��,x�]a��Ik�U�O�����#�j=BRi2���+�	L��(���v�?m��}vd��<0_j����b9�$@cN!��a�xFd�;����Oc�m����ttA�^(e�F���D�u�{������,���U,���ߓ����f�x�m���=h��gZ͔��%}�8s��=m�~�&�<�S�È:��a�;֣��� ��C/��0ؗWdVZ�O������npæ���j�z~���{�����4�>�(����o��"͒e	�����5W��+����+m{q���ȅ)Z�,@��য়U&L$�玼�`H�>�F�M ��qk�\CAf��G&me�ě����P��/�c��L�yף����k���z� [�;�Mʣfgo�Qf��-�3	��FONGhf�����Ţ�{L̳����h��p(=,*%�"����hT3CHg�yC��,���Z�9ۄQ]�Iu7Dvw9f�18���F|������V��^�]�1.��r�Qf���X.�@����W��<�Je����>��b���a�����fS�~ɣ��l/VA���z��.K��2Z+��׈��͈�ʋ)�||�,~�.�o:���������W�&���jIa<ۆ/���vz��mǘ3�A��Ԡ���Y\1���=H�Yc�����V����K"��旓��P�@#�����0�u�5��mMj������BP� ҵUE({���ב�[Q4�v��Y�J$^��A	��dI�-�N�4�hI����q	n���\
��P����{Z�j"@� ϓ)(�\��J2�H_7n��;S�{O���cv�]���� �&���؇ �S���*� �_/,N��M_�� [�u�/xn�r��W(h��Hh�c�&���oN���ٹ!�R�����䮂��m�&�$A�([fl��!�p!��	�Z��y���*�O���v���&ϫ/����	g�+�y���H���|�12
�
��n[��]�c�N�ǂzX��r�ǯY�u�H�����+1��\�
�f�%!����rn�H�^�������{0Vc�C�ɘ�<q��~M�/5���&%���v�dd��A09�R�%��GZ�"���"l�P�`@� LE�i(�<����;|�7����d�e�h�������K_K����I���\����c�ZL#��B�$0�.���iD�c\���9�%MzSY����n�X���xhAc�ݪIU���,�k1��T6�?]=J*�;o�0��Ǡ�]��S�Z���}�KD~�Y�F����x��R��?r�]�id����e\I���Y�9�mЉi�9u��ӽ^��f6�Мވ��2��l-6	�j��l�_U���qL=�7N�9<¥����.%��>�6�(O"eK�E��a"�����C7���]�2�)0���Y?����7���a0�Wq7W�ff���o�ٟ���������Y"_�Dsv;Pt���H�F%w3.��.;�Ֆ+�X`���ո��M�pA;C�G5��؁��«	(Ͻ`�e0�wL��J��)퓼��	��5:mV\D�&c~����/~�e 4��K,��@���s�	1,��Ն�t��Y9�����b�Q��m��&'�F^���
�&V��P	�ǎ�����L�k�oRpI�����h:~Î������JW�ƹ����܅:��5�pM8���HN��@F�J`&Mh�̨�����,|�0B �ސZBǊ���p���a��w��G"?�L\�L����M%���M�۳���V�m�������Պ��̙�p$$���u�0�4�B����ι!5�����)�0����Oҳ?V-,{��<�@�2-���d�l�~��ڇ����=30�7p���1ϛ}[M��r3=��m��P����@�)��xR�ʪ#h�����eU6���С���NNh�R�XI������-��0�40E�Op��z�W��-�N�fst�sk���������&Fy U. ���E�wob 31]MϑqEgJ��+<�Hj��PW�
s���o����z.;��5�X:�&*����Y;�B��%�Wx�NnG��#nԍ�`�=(@��x��v-e8֒c4}Oւ��o���i:�f��������y����a���`5�� ������KZ�^HV���\"aИ��]C����k�&O�sS�1,��Q.��)+�SK˂�9/�R;\û.]�ZA_��I���sF{9P�2�Ǟ�� X�+�wM�e �j���i	����*{�-�&���)E���`��
�8U�� {�I%�������k��ޒ�k���\��zؒAy	�oE���2�V� �u����'�$�^�%�,O�G%�c>ni:&�����ݦ���'.��	w���Lhr�γ#�Dyof���tj�{�J��Rܣ:���`C�1.�A���@���)�C�o(�	H�����H���:�1�tU�>b+���:^�����R��oUxӂ i� �sX�@�/;uS_B]��7wa[���A+-0d{�S⫽��GI)Y\���R�t8�.0~�������f����y2�*�Hy����b0��ԩL��f-���c��;��XinY��zD��cc�1d��z����jCK����]hL�孂}yS�_�Q�ZI�kR�����K��<sbF�lߦ�1��R�G }��K^�_�Dn��h�R'`�`����S�/�F�~==�s�;_"�~%j���#��Ǖ:��i���Xc+j�P���,l��
U�F�&#q>ć�S���?�s1G4 �slʋ�g����Յ�v5�u��+I����NV6�=>�{6q>ϗ�C��uyk団�8x)v
])���gw�Ak�+���/�f�?�b@Ź�w"�f�	*-��Φ�A�%�r<(g���ǹRDnHNm��@�طI��t��C�/�ޠi�Jk٧����
4y�<��܊y�(e_+Atc~�C�Th�����M�ج{|�dg��� vzd���g�O0i��B�;v�`ca�m�u�<��l�$T+�|Iqo�Y��?c�>���Ў�z͎vF���Y\���Yp@2rh�a��w,�e��R�
C*X;��Ժ��R�����p��7��	-�/��:
o���������r������m�.��7�Z�w�:���n|y���`��
��iF�[�6l��wdan)�A�!�ή2Bf���Ő}��F���~`y�x�ۗ���̡�)�*�mb�	A4��Z��X����uU��(j�x�ɰ�=�z����R h���џ�.��ܭ(�T�Ǥ.�G���D�&ν/$��s�#��Mk8aL�4ǔ!i�
_�Wy��\f^���#������א!m��+v�u���D�c���I����O���<���9���8�7c(�h���l)Ns �n�F���C������Gm�D"*��/���tK��?�]��8�k��\<��ɌK9���_�O�����m�"(Q�ַhF�K��P���M"Z��Ց����W��F�C]#vN���dɏ9FV��s1�W��x:"�fT�9<�%�WMa�kA��?6y�i;��,�!�G��j���1��iL��Fj�ȓ�H�%�B�l��}PxK�w&�:s��AqN��,��i`�'���4Q�gn�|`�_U�׈m�TY�m�Ջ��{��<�~ܸ$ǔ�et��I0���j�V��h�g.?�>=�i�Gv�?��5#̧����܊��xe�:��xQ�Vg�'�$����K�#��Ӹ�[�9�R��2��s`WuRM1>n+��v�y�,	 �2�|�,�֍ɛ�������]�	���]�u�P�P*���GA��x�E]��[������$��ezIu�'�ث��U�l�{�j�H~�b�,p-�>7�e�%U�&J�tC�c
o�U:��d�	b8���(�W5*�"R�+�Db��S�*>[��P�{z�S��¿Hc�}�����ބy���t���q�>nw���^Z���/�0c�U��̏���2�ד�oE�vBt�5�������u��mv��E�N�I�je�L�'��p����s� �Tc�yRR7�PX�6�ԓ�� n�N�GIh�*nX�\d�D+�W�E��K��Ǯ ��U	�*uK0�/���o�f�gR�����XU���Ƨ�����>��Q��Q����ƈ+�*���r�RU+��;��r6�Ն�!�=���!�8:��EQ/D�%5+ǌ�`����W�����lA	�^u�y����������,D��c��Z�i����ue��-��q��+�a�Cy�F^��z�W�Jn�Z5�; ɬ'��
�b�&��ޒ/#*��Ds�gD9ȇ�Z0q�E7�����Qi�#����� ���LTt�{HT�g��4��ѷ*������[Y�x�N����y/we�!�)(�|n���|�:�r8�-�v��5�t�-*�q�^v{;�x	�֬��)��m`Ϫ$ɐ�i-�4�&"@f�����k�lG駀|)RP�ZP�5�D��p� ��(�7�{�����ۖ3��M�@j�/uU����,�4׹k�� `<�	��<�I!�͇�G�0�BF!���T��2���Z*�?�h��#��=<�`�M3`
�dj�̈t }U�7f����`�KO�;=�*.���u�C�B\q�f�|��	�σH�Y��e�}�!Bk���`���� �&�]��)?^ڵ�<w�\������.4�Ƭ��
|m�l%o���ٍ�>�-�`)���K��Ԝ��z�Rd+).�f�0M�0ґ�=4a`����#,@�1.mGP��@�9;vS��=3�&4.�H�U�d�[KhUt�}*8nr��I����P��t尻���b^�r�y�Wf�Ŕ��������\J�����^$g��ꂐ�XᅿG"6��2���3o��$@�sĿGa��u9��V�Q�������N��4y�,DF��V4r O��!<>b��ݣ��jt�9��m���zr7-wQ.���6��9_Т0�i���S�s}	Dx�zF�r=�G�4�Li��~�~ιJ͘Z�a ��~H�"�A�����֋�9*@~5�!|�����-�A��O�̨i��f���{0]�q�xn�w����=��FQc�]�׈����S5��?�WӺFK�hB^�E�N�B�M&E_����{�#1�XO~�Y� ��^Tg*��>|�ʂ����|Duk�Q�1˗ꀠ~�NT
��8U,ڋ����Ȇq!`���a�f�����?��yA ���� ���y���)ǩAY�!EK~�D��T��f������1/Lɵ�۳�J�$�����=�!Y�9�^F������Ǒ%ߔ�R���.�(F�;`��S��C��*���������P�da6��rvh�c�������H�I+"�Ӊh4��|w$�ھ��|������W�"��D�HP���	q�#u������B��0}�M�{��t.�9�ljǵl3����B�!�=W.�g��ъSlBθ��{?��qS�ۨ*�]4�N7< ��C�Q
e����x�I���@0���u��n*�gI�LQ��V��K����/�m��D=]Ϻ�t�%�@T�(�S?3s����sĘ&24�_p�_��a*c$��)|]kGFB�鏭u`2���.�i]](,�PP��k�[{ڜ��}j�nA,6��{��D��/7�1ɇ��)�d{,b���
_v�>��g��X�0-bn��АAe ��������f ��+��$#cR~�a@� dAl�O�-�\��`�Z����vQh��ndk�R�����k��%7�B|ŏ�p�+K�T��T�_�D,N�_�eG0
cJ�d>xb��R��w���D��$���o���e�\�FcO>?
�S�q�gX�ݦ�����Y8�h�5��Q��ϻRIց�ۛ�j�v����>D*
��KB�����8�������#b�w6���H��l�-xG��t�mI�A/lK�׉����.����ET&���G�e�)�E�Ks�hj0��I�-=�
��A��/(���Z;Q�@�Z SKB�BpHKBO�_{Q�Qub�=���_�ԭ"H�P�l�=H/�{��4:PC�f�Y��Y�,s	<����>y ���m?$e*Z��O��Y�U��o���>ni,�|jJBA�Ѽ? �^<�����収�mRn<��B]��s��36�>���W��̅�o�`�V��p�n]u���f�<0��r������+���@�����RO�s�Lŵ\OS{����N�+6Ȑ(�6|.��deŒ�Wu��Z� ��HE!��K��;�(�l�t����B�;�H'lͼ�Ao��M[V�d�؈�\@���"�A/A�Yhd��L��B��^�1%;�1���5��`�얷u�f�=� Ġ�T�kԅ~���q�h�Qg�M������摹��o��/���¼�ȶ(5²6�ΦG� l:T�SH
�I��p�����G��O7�<cdva.ԥ�[�A(5�	�Y}�#����2�C���[��;�ɍ�;�W\��u�F��A`��$($�oxY��qB(Ơ3W�ď�&=>�0ҝ����~�6-�@�z���z�A�:��YpQ�u�ҷz�e]+�cS�b�ϱ�<��u}����n$�,����s/7R���m;��(��g3YC��~�2Q�Y$���[o|P<&�4�5�^�;y�~�yE�(�e9!oĞ��C�s�(3n��t�#u��f�p�~���z���H�X%�ryI����-`W��S4�!�}7�P>��������g����h��^X񀄵��{�������޾+�QP?5��D6�+�a�@HS��(���.����Pb��Nؒ��y/w�Q�L-�����$^�K�XS���'�3����6��h���K�T��5��Ԅ��|j������U�IU�қU��]elJ�n�k.ye�(�X-��
Q�K��K�k����'�Hz[�<e �(ڂߐd|�Z�B��J�r����(sE��$3̙�	���)9��X9C���Tw�� �zoE8��b�/"l��8w��(;�y�T�^= �{� �C@[�{ϔ�a��XN�3pbz��t���c!�C����v�u�3���jt��y �IG-l/��?H�0�vE�\���c���q5%W�אb�9�i���W��i`��X!G���H[Ra51����ͅ����2�d�D̢p��!.2��J
<�Q�'UT��WԦ"I"3q{+��T��)|�:h>�T*�8>�k'���7ݱ�c�����������<4ɖ��/�Zy�h��	v*��qy.<nyM��f���wf��z���� R�1|��5,ު�S��*	�H�D��<��x��s��	�ݢ�W`ڋ4~@w�+��wm��l�<)�FY��<�;F�,n5�ό4%�dnȯB�Jp',�	��/���}�"��i���*��pN�Rδ�v�Mu9K:�?�d�B�y�V��x�5�v��1�\M]�ڛ%�>�(�n^_/�q��ф�91�.@̲�@��ߍX<�.u�,�ݒ���Tz^}.s�JP*��#��Z]JyN�W���E�v$A}?YQZ������c���m�e|fa����E�RL#�N����ͫw���Q&��
�F+�'�vݫ��/W+���� -��g�G��6���"ѷ��_�B�~�K��Q�`0����r��AG>�fv�@�]���ޡ9������=�fǾ�DY���{�O�{
q����-����f�e���`Er��ː��~s]�tv�B`$������vON�.�-�&��Hy2pc.Pp�|����R3��8]l΢>	�gU :���*-F���˭!��lu�B�cཆΏ�glLv2�r�H
s���%���e�A?�!���{=q"��:�ϟf[ȯX�#Kл��b�=���<v����N»v����S=r�N�c�qi)�@7�)��������������(0,�����!f��b	5tK��H�"
Ĩ`�k��,������~ƛ�!��F���b_e8:v�V�K�Jd)�p�V���&X<'�����E��eUR7	�������Tp�g_5�jf���0�y��MH(�e����?����(ŝ���O�C�׎ ���H�[4���L���g.�Ӛ���	CC���-���+޿�_�X"~6{��p�s;�R΁���-�9I��dS#��LH��?�ث����"�� ����d�$�`�c�)���-�`HcjS��%D�Wv�������� �`��7��5N˘4�P(��V>�i�a�רd��iّ���li�*\���G`�_��H��-+��@��K����ɐK�̋�X�L�,/>:޼I���R���֪G�D��p+@�\����/�,	#\��7�6��~ƶ��舑��b:�H�Ó�q������Ӄc� Y�G��K���H���X�of�7���'#T{�fT`3��� �)�H"���4��-�&��{�<<�����*.�Ǵ���5�[O$���P=��M���?��o��7����j�-��k ���Xx!�������cY���o\Ձ��*6Hp|l����X�r�E��MYYH|M�x�͡1��a��4�R*��������� �e���:=H��z͝�Ƴ	T�m��J8�:<=��;2���pO`���j��r���(<=�� �6��F0��Y�қ�=��sھA�C��&��b����L�Ke竿k?\ԩBd�x���p���Z�_{$7���VV��ȁ��90��6π�nr� �H$b��0�$���/�D�K6�ͼ�<;ܖ��z	�@a(t���E]H>��;���XmI>x2,�_���&��!=����I��d�:!+V�	�x7��|\*F3�?�}�������:�ٲ��L�{����O��� ��G!H���v���b�Ӭ�>�nxNdرr{��Hy��}g�����ƛIr�aU
�b�Dq�4̚ʩ[Ā��gD�1I����ߪ���� K`�C��Ϊ��g�& X\����G�w&��6.n٦�o*�ڇ���b7#��2�i����{����E�:C[�.5^�@W|�]��8�6��|eE��*j�$�P����\S�����s���Z�g�5�Ʉ�h�O�M'�in�'T�f� h�B���������!V-����� ��N/��\7���p���Tkܑ�{�����BW\W*U��j��Mc�x������s]�\��ҥ������6RiyHy��v��u�
������f��9F��k����]�&�S,�HQ@-Ba�8Q���,�JF0[в�.5���]�#e9�T� ���Ĩ�.�	ƒJjt͡⬭A��J��M�m�2F�[>	ry"�nlv}5$&^W�{+������P6��ㄏ1Y�3)��m*��(x|������
.
 rr��k�بsD&�S	D�0&1�y��� �����|d�j�bO�Vt�כ��[�1$�R/� ��A�28�(H�UON9+��C��
���jD�^�>y��z�$bC�;ьYpO�,���>K1�.�
�pP���:,�<`M6\r�r��W�LX��D 2�t?�P�H_��7R���T�������R]�p�*��MH=��\ZH����9R�Me�l}H�')4P�y��Vs:uj�s���ߺ]�	��9�"9�2�HB4��`i��'�1G�671W̹���yWikyCI��� �ۓ�0�7���qK�g�*D����J���.��*x�ǃ4u�z�#��q���ltiK[��ؔ�EU�!K�
=R�MKrX�i��+���M.a<J�:�j�6t`�$���Dm&�;I39Gg��~��%Ca��I^7:��2=-GO_E��_,�d�ގ����M�
�>և#��N�R>��ؤ�Ʋv)0ʵ�~h��g�x�&l[.~�P�:^�qHu�\��<�S^ՔTC]ہ�֦�A!��hCo��_n�bVݶ��$���7y휓���r[�>�>p��{��P�C`�+^y;*���T�j걨�y�pf��u���� �������ͩ���1��@A1ƾ�IG~,/w�n��<w�Q��:����zs���i���O �'��%�[k�|�Z��?�?��`7/'��M 8Z�+<�Z6і�'Pg�Y��9R{�����U}�F&#T�`��<<��l���Lo�޽w'=�7f�!]:wi"H�ٛ�ra���^�#�؏���-Vz�( �k�M^xF�;��������&(��A�x�e���W�ΙJ\?2#¯wP�����,9ѧ��F���f���2I2&Y��>.R#<�q�7��W�2J����m��N�ș�?�4f��Y�k%��2*�ukU�	��o�|?��<�g��zd�OS�#��y���[J)��1E��b��eѧ��P\�f9:z����a{�G�)���O����w%Sg��)j���޽��w���sQ7��[7c7f��w'^��+ꥭ5���ʛ�Ä��S�:s��I؀�z�),s�H�ڻ��]�emK)�a���¦'�?�$KȑQ�Z�e�p����6E����9��̌��QD�S�\�o�P�{L+]�ջ{��3Z���*Ӄ��P�)�°w,
�,�����1�>�����# �[����G^�����O=�pW|D�ؕ�#=J��ˮ+�x9�n����'	J,@�Q[�"EѠ���Ҷ��3�d�;R���ֻ����⺰�Y��q��;	[�Ol�Ara�������Y(��'DX�o��퉎��b�������z��Q"�?�u�.��C�:�?��Bv9�a�۝�DKz��mΝvK����닺�~��uB��lN?�U�s�U�����'/a>3a��5�W$�ͫ�86�G��$���Q���t]�mNs�:���Qs&�Sɞ����W�5�=��A oB&9 _G� e SNs��'�����'�HO��Z��F�80N��sm߲|k,�q�m�y8f¢n�7�ah���2����f��f�=�b
����%H�ND�r#om�v& [kb�p�.��	V��p���у����j�6�!�����vJ���pto^���B��5 �0"�����3����v�FJ߻g��q���~�Z���G��n�Hd�T�ɓM��t'�z�Y�$
y��?w��[F��5F/��t���O�Y2�����^�1N�J�!mk��>�*���9%���\O8[�m^���2�4��d����$����7�H��4�	�v���PZ�T�kQ����/�����i�-��B8s��|�h��|��t�GP��$�d�O?H��w��3�g�G]Q`|���nWu(h��op��ܯWy@�Mv�*�u�}�˾�����*�͇����K$`4�ڻ��:�R��_�c�{��RT������d֣BL�+/����}r����m���'�J�dJ�`���e�s*�;�(ˮ�>�@>�8l�`&�7�'�c���N��ɵf��b��<�%�"�+��M�4��l�P>\}:�����8'���ofDN}^��ރ�tt�+Jχ�ߺ]$���d94�q�q'�'�[��a�iv��ߜR����`;�9�|��X�9������f<���F�齖��n��. ��dcP��4U#@,��j�H[�M����;W�zZ��$���%j3,�M����Rs!�Y���@	�٪�6W���y^Q�����F_17H�`>�)5�:B
���R7缯�7[?�r,oԮ1%�٨+��o�_�S��!��4�I�N9��;7�q=i��I>ʑ-^�}jO��l��ޛ���i�e�iM�m�V�8��|+�9��RS\�+5I�io��h8����l��'�t?�:�7�X������.Qj|�g)?x�T�H��qX�9m`f��DB�
�Y�J4�D!����h��D[������,�����cQK��U/F1�w�ʸѾ�H`
�̝��k(R�5�֓�ɠt���\��ļ���r/@Y8�,�;����1���w�����d��ш��A�ned��8]�
����GP�H,T�[%ąײ�� *v6��?������Ky����?�.��攖+�@b��F���mh�`ړD��\ɘ1�c[��KG��� ��oL��˅,���d�20㤷���('�>�jmM�NB�J�}�|������7�i�=@�W󏩅?�<��cFan"k2}�D�+^V���ϐ��S�z���܆���@�J�T����ri�d����@����M�J���X�V�K�����A�g�'"l�ボ�o����Ad�rE�<�$������}!܆��k��_�:;�>������� 5��2��c��]U����$���EK�Nh�*_���4%�/A�>��8H���Q���(��NF��T���'.��ٿ���Sމ�]Z���g!�A��׃����B��������D8QL�X�8�z����H�fẛ�j3���N������kAp��V��7 R[xέ�N[rɥ❹+��Y0�~k7�]��U�s���ūd��3��_~v���?��4��~� �'��O� C�H�*��DI�jpk�L.�����'ł��{�Z�B� �}�c�,͸Rb|Z�x
����Z�X�`k��=n��>2�mB�,�<�=K��F>�qW������$ ��܄]�%]��$x�3�Y����Z3�t��b���Z?|�Ů�3mDKQ�YH�6!t�\E�
�Ls���7_�ֈ������n�(M|?PX&F�N��W�7�l��!~6���\+�珤��޼J�n�M�P�	����)Ǩ�O�m��(WHI v;3P�pd}�K,�N>0ݗ����
ݞA��i��{g[�Ǵf/�;�qu�֗9OL�������������R]��p�{�Q��4�R
�g��b�
��Ap�����UhQ����(����bA�,&E����� O�U
�Լ�o�s���0>oy�����t�:���q���� ��I*+�����\��c�KI5�`% Խ{�ladѹ�Z���@;s���W�6fND��6��h⭣���م`����.��h@���
<K����8�;�~�hY��:��)b���ٴ�LJ�V�ׂL���$R"7�v�fnG��QR*>��߽�I���>[;�Gn�3Cۣ�5/��Q��l��m�E��L���߂A	��m`W�FE�,1U�b�\n�)��=|2tƵ���D�d��� ��+�j^��K��1�@��B#M�Û�+��*
�7��'�󬉖qS�$�����Ѷ��7qX�ch��F��h���wY+�/�@ =\M�G�ŏF�R��z}ΒW&1�z���~W��y���uV�����/Nj�g�eJ��P����4��T5V�^rP�ʝ%��t�f�?���� F[�s��I�inQ�N��f�M=³x�ZB�p�3��܆1�O���2�o��R�� �����u��nJ�X�E�q��]��"��G�������0ך�ʠT��Z^x��[{����0+��a1&����?�F�ם�����
�b^�_֋m�,z���CC��&e�j�+����F�%�S �խ5����� "+.���rN��:N{�2�<O���w��D����>i+R��.~�M��U;��_Ի�FP2-㣴KV�-��{�_*b���: ���n(�w��;VS`�;�~�L�Hz/�Q� �F#	G���_��`�Չ`���.�а�gr��%*זp`��xj4�D����T��F������P�-���-jc�i�&�J{#�+뺗������x���<����h]�t����A�/��D4
�� H(�6�l��B�ZOr����9��v5�\�ehPY�����ښ�����R���rB�Gqq��6ා��uka�#	&��'B�C3i.о��y��ǷҒc���a�Q��(�Z:Ja�uh�:�O7�ܼw���� n���y�k�U݁�Rg��ӗ�/�C''u:���D�}3Ў&�E�T��8�f\L�/�Ҳ�^s�	�RW"���ӽ�Wt�����P��O8c/�H�܊�^i��-��F��.����Ú��<8�Q���)
��瓴��Ba3��⫾���!� 	Sso�4^�2vF������E���T�.FU=+�e}���|b"�V��a#w��I</V�l��T�b��v,�H���=b��#z��-9w��J�2��/�=�O�AډXe|-wm��ws��e��\�8�~`�ư(P{i{,$l��Z����z��+^zi����FW_$'Ń��pu��	��/�d��d;G����`���3���Tz��
Ո`����]�޲�~O�QK+���ߩH�2K��XuL����=�/�ռ��Ty�g�Z�����6X`�G��������
���"�ߚ��fȦ�hq���:�����<ʇ���o�f�c��0D�/�%5��K���h��I&O��ma0�&B��b�y�Q���M�3<�s&�݋��:V��>���W�\P1W�'���&���Κ������:Y���Vz����jIH��SN���^�R{ܖ,�n% ���Qlm�!�}�R�g�c���<�]��U�0�F>2x�D� �SQP��n⿂/V��Q��l�˸�e��M<�@SS����Ū�ee��C:	���w�.� Ye��S���̴�UOD	����i�pX��a��.3Ĥwf_f�|�*!!�C��A�W|�AcO��$����^�A(���C��R���4RVD���ү��N�f%���f>�EQ�^�(�R׹���.��7Z����v�K7S�)2;��G�y<��츰� �Y�/�o65�&ArO]P�3^��$M�n��'�ă^��Mk����ɏ�4���ʊ		���/j�j�hnE>9G����$q�EhQZ*�Ny�S�~�w�������p�q�P�~vCSQ5�i�3%�EY��u!*����N�U�XGE��f}����A��I�=�LϦ��.u��̢3���0 ������c�<�2S�anq�fO�N���cܘ9��V�J��Om��l�^�xs���D�kF��&�]��|4`+e��A��MK�|��b�>�1���67 ~7Z7"�S
ӝ�|�Z[�7D��4��ڋ���O�6o|ߎ������!ng4!�ra�<aJ����ƃ�QK}J� }!`۸ʜ�E��V6��^�洇�������	��C��r�(Vs�C�:#�s�z�L��_G��۶���K�T��A��h�HA���^"��٫D�������,D����0~�־X�G�k��P�X�z�gzg���)̈�̞�-q��XE��|��eyP#�;��Qѱ>E����Dl����>T�"�~S/�OG�������҂�	8>"�v��^i�J_�2_��<b\�P���g�Q=��[[�Y������|���xd�|G�m'��^CX
wh���,1������W'�O	��k��P�WSj��T���<��:�6@�v?�CM׃Z�H�kj�6�Xj�W��)�o^��v	N��,��r��w竈x�)��8�wj�I�$�7���Dɧp�5�GO����r����)t�N�I:���6�K�',��wY^���X�q�[�T�*&�d/����E�8�UR���ǰ:��� }�<G���"���^P\<5�~}�(�V�K��q���f�M�.��e�y��B݌�0^�A���?Cy!?��d��j��Py��ԜQ�u�ȩ<�;��.q��ɴ��x��O�����8J���ߎ[A�g-�s2�n�*�C�߲�(�ͭLS;]�HX��qdVW��x��g7|N�M	J�V{���ٗ��Įw�W_=����9H��V���K���B��*xgDnl�ӿ�9��O����W��W���s�u���<�˹DH�p���P�;�֎��}��ײ1ᙐY�%�3���G3��)o���f��51Nrڠ�9o䮁l�dΡ�%7AJ��/��f�O�٘����.�+e��3*£x=pV-�|�Ǽ$�m�{(�e�w��5�������+�΋����N�K;��t,��
�ﱎ��HP��&��6!~���g;i�R&�#O��tL�{k�O�;���� &T�<W��F$T���(!��hV���W��P�O�����A�yڊ�8�ŬR@�ܬQ�FG��h��=A�L }�J��j�Y�8۲�Q4&L:�����(�a��#����
�1�%|_��^�Wo��v0ǧP�X�=q� �j3ÑI�Hs_3�A8��#�=���E+�r�C�l��Ӡ<�Ȁa;	���y��?E���F�����1��zJ�,��TNfpz��0�^��T�����O����Ǭ��c�DDB,�k�:u���q�Y7XB�I�x�PPu�Ɉ�NK�A?d7��3@�� �_�z�鴪I4}��cv���|m�0�{A8���3�6����`NWF�
Q��ζ��^ʢ�Z����WWT�Q1ͺ4Wx�*r��_���������A�y?�>�ig�4H?~��o	>���N��s�4�n�� ��l����Q	�s�R�"����fK&U홺�N7wL-n)�O%M@�{��l�P�w�U_�4��I����pP�n���I~�a�A4ݿ��=L���� ��a��Ԏ���6ā�"N������i�#���88L�w�iht�rdtG@��':J)�m[J���~M��֧��V�9�'�D3a8|�	F?z�P�ꠣ9�EqQ�֜۸eS�-V\S�u�&�s�ʺ' ����i����Ǭ"�N�<Y�F�,�E�}��-y�ץ��h�Cc�����x�[LH�f���ai��t)��w�
w���#��!��4��nI�D��8�����7���R�Z_�ƅg�
S�	�	���0`5X��HD*�0�����ԯ��IX%�u���8���E_~N�"N�㌰��6�z7E4��p-l��\j��<���Џ���~*'w���?�:K�^f�$�T��}^Y	y"�-����MCI��t����o�6�$0�k�a,�Z樄ZX�� `ZQ��܀�����k�e��=/��Y�т�	A��r�?u�&J� ����gl���'�L��GBZR�8�Y�sŻf�H��
�ۏo�8j;��D��n�����C�u���.Z%��*���&No�Ոש���򄜙��qzyP�e%|_�;J�$�+[�8���^���Q�.�3D�o�	U t+kw��X�"{�jXHl��|Kw{����5c]�7��g�0���&`���������vXH�B�6��rR9��&�9�+������u��I���|Dֹ��J��0��^!�C�#�/ݕ{~����N���N�
��EJ��|��v$�Q�!���?<��U8����]��i�0ht*��@���b�}F �x�����3eU�Q��QQ&���l�)� ��E銦�d����!����BQ&���ww����U"�j����K��I��կ��OD��Y�YP����Q1��$�Y�*�}�������8a�F����C���-� �������z��=45@d����M�zdy��n��Ekɔo7F,����B(i��8	�"]1�d�����B���z�\��;�F�'Q�}�0�w��i�a�q��o��Y��m%�ꇸ��U"�.u� :x��a�8z��ԍ!�2�eϸ�9wb%%S�b-�S��c���\<����I����^����aś⇕&sj�KA��}S_��L0ZZ@x .��iH��Mn�<� 2an*wbQ����*�E�GO��'M-�q�ѽ��_�
�$�t�D����"��|܅J��^���i�-4��+
[g+���݁}�1�3�:�o���8?����(�g�
�+���M���/89g��pc;�'�C�h�7�n#�� ��H�ӈ��8𵰩,N��1d��C)O����IO�j����a�*�\�n�$�yJ}*�*5�W�S���8����3P]d�
?�4���4�@�=Q} >��_�4�ֵ������{n�>����]Z�\�%�5�8���*���LE8�R�^.�6�����J+9s�7T�6�xX��P6�t=!j��c�bX�Q��,��G�b��g��y���\�C}X �حE��G�L��F�L����`���'�R��ۯ�3%���dHN��M��z��OA�ٓ.=�����T��m�_q��gW<��Gh0~m$yv���w�A]҆�	q��'�!K�>h����c馾���K<��dE��q���jC9[9Ҵ�?�>}����`f#t�$엢;o�.�Aq�< ^eh2� 
�QA��	���YKy;R;�,>�=��.Kw�5�0� PrC�y62��{�b�u\�qW��f�T�"Fd*҉���ʶz��&<��o4�f��S`^�'�H:�-�PغC@�tq�MH�_͛������sH��s	<�#%D�>����0��4{��}���x2W���]Ԧ�r��`���e��}���9��&
�Ѱ�s���㟁m�H�;��7�M�zD�գ!��E=v�χ1�7�nxOM]$�i�ƥG����6���kκ�����	���@����^�8� l�Y�I��TNv����3��ĂeH��5���i=
��}�����"^B]:�ӄT��8;F���I�q`���>�7�.�,�C,��ȋV�@R�L�~	#����0a~[Rdc�0�XB�½�r�$%'�q4�-����ȍCǀfD�y�:��F ���1wI�ϲ'f�eYޜ~�ܯ�xڽ�K��g�6�1"Q>�s�_����'�K��l�z��R(���e��\�� vBb�fe��i%[q1'�3PݧT�&&��Z��n�Q�C�3z��j�6�kǒcPe��I����2�']Y�;���'��Hpժ�q��u�g�W�q��#����Ʉ*�}sv�Kn�
�{�Yբ=d�T(ԭ̖�ո����**6sx�N�r�5Se�,O^����Z��Dh����T�B��.�;��,`�*)r�%�}Z�M?�L�F܏8�_�ͳ�Bc�7 ���T(���lE���v95G����g�Ѥ92�2H^N8�*����ivD��Q�`�G_h)wAXҶ#��h$��a�sdNH@Hn�@	S��O='۾`�#3[������.�+!h�������nfK6|o�%�1r�8T�KcNb-p��	�9���M�nO�N7e8W�+��1�~��-R�_�E<�mÙ���,��3{-%@P�O���m,I��<^m���i��޼2��۝��J��m��e�q�`k�eM!hK�`�C*��+P�̐^�1[x�R��]�ҏJNÏ�5aw�Y5��z��S�W<M�,}}�q9E�*�xb�c�A�ؽu����J�+��C��O/`8m���]>�2h�7�	��G-�R��u���Dp`�#�T��~��(�����>p��ֆ�r<���d�D�-�%P��ç���(_8��0#>��8ŏ�	����b�|��I��:��x�.��L�*:�^W���A����,�/s���(���lr��U*�	l=p.-z1NI�/���e&�܅mӇyw(�Ŵ#Y���S�%�[��]$@P��$~�1��#H��ώU�t6�@W/���:Ӓ�4S�!С�N�������%�M����\�p���ͥ�D�� �|�>������Ѻ]K��-�]��*E�̙<���kpz�]%Z�T�N ]�M0.��~�#U����sw|pf\e��������Oh�]ށ2(Y{Ni�{j�t�'	��s 	^�FO�d�NM@�3�R��P�K�Ա^ڇ1(���m7�# }�&�~��\Њ�^h���w��[.ܳ�Gj���"���D�^݆$��>Л���9d����5�^9��Ԅ-�M������D�1�<Ǜ�i=���]ԐH�k`�6��'��=��i��L�qM������DfX�酋��]���c�s@tb�v����/l���Gx,	S��v��È�W"^Ck5>�ه7��^�3�G@�;��t���~��A|x!��Vx�c!�\���	oX�"�#牯擬s[�&�(��1_������L��mz5͠x�6�MU7�}��K�C��:0/�J_�w`�O�v������Q���s |�yB]6?C4����cC4�t��5�͏����,�˗���,�V{ˈ��F6�л�@�(I�E4���Cy�	�h�C���$��h1)E� ��_��ݗe�c��2s�EF۹���aFDm`'���;�I�ڮ�y����/�C8��.��+���i�h4Z< P)�vM<�+�H!��ŀ���}ܹ�Z��F��>�/A���L�KI���=0�Y_C�����ԙ�<Q��<��0�(�L1����/��ص�rb����/>0vv�}���3n����׌Zr����c ��A��L9^O�ӆ*��'��:+J��qf�o�~g�����u�l-e�4Dv	�_��)[�E�xwJk�y����;D<�k�r��p?�ᶼ����8׋m��N �:�	�a>D8��Mϼ�]G �f���?'���9I��`h�!�f�W��N��`礩)��.��N%qW��G�3�H�s=3�&�&��u��ևn�f�p������I�BS�*�GN&Ԃn�l���'��ř$�����{�Eš�Cl+�#9�X�S��@.����,���� ���Z��˙_���:��d49�<a��%e�����J���N��[�In������/&,�.�Sm)U|���~%�G�
�U�n��ˊ�Tywֵ� 
�(�J^0ǽ�-��	2���o�8�����RT��_2#�����o�~�k���8z�{"So�n��󺷊>�&p���i��I!ƾ���
��oe9�4��s𔝒�����onV?;�������r!G�w`"�c+�sqς�{zHCX�M��k"�B��K���PJԱŭ?֙��HU�!�ˠ5��s`
�2d&��jqeq���>!�D q�4�q���\Ž���+���` ��*��`�>9�+�d�}I=�\PbY����D�%��܀�*ؔ=-�9z!:P���Ʀ�����,Y��[@�|��e����T$@q��܌��=J��.��2���,q����^{�V�vs������ ���w=!�c���kT�~}���U�2��$_�UF�{���|M%�q���#(�iٚ��vOU�2@�~��Y����jݾ�v|J��!�����
��D�+X��U��	��jB��}>*���ɗr!��{��2mv�ͱ�:�� ��*(�ǯ�l���;�L��p��x@fǷ|ǍcJ��aU�^R8�@��줍�t旅����0 �Ԡ�%� O�=��4)����:��z>t4�����A��V�f}�"�?K����ˎ���T m�2��X���M�"U	;�RNK���%j�;���@yg�ҡ#�z/�w��\f���w~��J��D(d��dH�;����\0�H�蟈K���Z��q�e����r��f3ZT�t��|����2�z�_>^h8�A����3)֐FBC>X'k
�y��Uj�`>�A�:��h��l��s΅_<�fhc�1�_OҮ;	gۊ�_�'�����: ~\�>�<xm�\}S��R�� ���b2z��4��o�|M��7EZv��]�^� ��;^�W��WO�}��dq�n�k<��l��Ǆ�w^ϩ���XKBa����a�b�qp�m��њ)�����m��N2���2UOV$o����/�Sp窡}P 2���J^�(66U����H��x��/�ȅIC���3����Ϧ��1��[ze��?�I�c�Ǳ�����R�tt�i5��p��MM��=� ��O~����i�_V�3�v�;�%ge*7Sߡe��B���PhdS�vH��(�� xm6F�;��E�z�"Ĳ���@�`��M�ԥ�u�i�7���c�5Nl�*"%m|ojM��4�頻�V��mw{��v�Ю)!(�����&ɲfi/	��1G�&����m���oZ����*	I`�w��7H����[y�V�ν��]2�DQe�#!9T7�~���j��S�NfHٺ���V� ��p�W�ī�ػ	޲dv�$�z�4dqE
G%�Sp$�[n>�M�D/3Oy�ee��jϢ(�<'2͢7}w$�s*|�4��7�"��^O�~�R���
JI���=8�I�2�k�Ѕ�bg�w�P���,�<���ta�i����X ���{Z^s���+q'1����7��`2.6R_i+����!E���i��'�0C���K���0Y{�m5����E�9Q�E¬=X&���\!�t���$�N�ˆ:�SqϠ��K�q�IC�uiB�!�Ԁy�~]�vC<��Lb�%����3�=�ټd!��*C�����Fo���B�c���ų���Ǫ��{O+f���¬g����pf�0ƅC�Jh��Ă'y?���@���T�?��-�<.�E�x�\��U�Т� ��њ"��t�L��^�|cnUDf��"���.4�lm �;$�c���!��`���J�\�a����7�\G��s�{���m?f��_��a���8T`���>P%�x:�ȓ'�6v�~^Nő|66����m��f8dz��`V"_�W�7�衟U�=���w����E}]����2�XL��sO���͞���.�{����.*�g񭲿�E�z<=��tȕEKG����tq'R���f��T��+9U��z�(%��W`����q�ղ���'<>^@�$���sc��^P&�<6<�j�*��b;`��0]�_�Y���?HV>��T������ŏ�P�HUL�ڣ�s�	��RI���h*��Ui�����F�I��]ش ��yQ����zt�i�ߦr ]h �����ˌ�j	OCu�Q�z�C�����O��wlm�'�wW�Rl$��m'�)^��̵  �w)�<i����7�:GiHm���Z�4/��.�V �.��}�2�8����KF\���m��*�ل-����-��b����8DWBP������)B6�����!u`��u��O�z�a�6I|S?��(|����~��QWC]�Y�����3>rdѼU*aq�"�|ɹ�f�T���|헃���!sW�h]����*ra5MGZ�߆�o:�!�FC�y���0�H��c�M���G�d�]��7�<R�{P)b��U9�U
D�Њ�P?�����j�B�r�n_�u�V��Ӎ|ƴ��@##0��Ù���(�n�gY�Q�ZRaH~���vc
;�-rK�ٕ���^�c+��7lJ���͍�'_q�;A�8���,�'Kt�w+���޻�MC�l?�*)I�C:wW�5�j�%ӓ�( �ZxNI�=�1�(����o�
<�HA�K����s�	�D�+��3�Spf��q[�ǵ92TM����֑'k���r��I2�;m+������0����7Q�-�;o�Zk�A~V�ZN��ڃ�͞��Ƒh�uQ���U���/{��G3�m��n����$��g�.�5ЙQ�t{B_A�J*��0�-> �<M��k��щ���$�����_G�,$��MtӼ�1&��f>��.F_T^���=J�BJ�q1B/%�u徶����}��ࡈZ9��f����"�N�ޞ��j���{/iU7B�ݡT�vj`��A.�¯�е������#qs�&��[�S�"'b|S��c�~z�y�����m�7"�c�O�;�E �/���#d�	2W9	��X���7���4B�}!A0==Bv]EI���9 ��ӏ��Ců� �Zf�V�	��Y�Q�!)��d/>��ʻ�2܇�z.�d��,S.~��g��oǥ�r(�HyX+͛��"���9�Y��ꫤ"Ģ�a	T+(��w70�5	���"�K��_�Jsb�K��"���FN�QNRR��7���j�-�p���;kg�i����P�@�f̀>��ǽ�hц���Ҥ�=3�Y7�����Nwl��|��!��h�6�����s�ؘv(pt�F79��$s���F^9�4�ktʧ��?E���=,�gx48�~��{���
	��2*�
���7WYt7��c������f���s2�D׮�CRgW˫N���/��0F��Dj�����.��2"nI�vP6�K !1Ҟf}LM�/��S�[��(Utk�A9�`q7���^�i�"*���Gb]�R��ϻ!;��⠌%w��t��A5j�P�Kr�����	������y�U����
���a���ws7pC}~����kz�X������_ՁT�*���Q�2�Wn��}W�D�a���9�������[(t���L�TE��l
�BOd�y�p�[�#dnW�!M����ݡ�#k.4��Բ��!I5�[E����<�0�V������#��BB�;ɾ]��<͵2��l����xP愯�iv��)$�)d	;ج&1�f��M�V٣"B��p���g��K��X�{��%!�хO��/����d��̉yw��-A� C���˘& /�%���=�q_(�+�An2옂�f,�gMhqӣX<�K���ݥ�]D_�����`����t0��l�S�Qٸ�)C+��:��R�2�?T5e4�C�:�0q+f�cxz�v�"��aU'kt��{��C#�U<�r����P���tQ��V���YA������A�3Q���ma�,���	gy4 ��=�8Fz-Q�r4�L���=�V�O�
I�Fa,3]-ژ,�]7�)^@����N�-i7��%3Q���:� ���D��[5�5��Pd��F>&���P=�X���f�*�H=J~�Ϣ��c��n�nF.�I/�������>�=E-`쵘������X�&*�<�u��Ʈ,_�<Έ����y(�wl22�@s.y�^�y�5G�E�}�RI��mY*�0���]T��b�����7i
Lۼ�`>Yu7!��p��X��X'�U�t�e��Z�LEU����B� Z\�N���� �+��8����y؃R�3�A@�(Sp���W#Zl���a���7����_B4����hJ���tЧ�������X�ܶ�35��n5W�J!��N���l����Ǩ8��
O�#H�Ψ�z/��}s�j�u��S��-�٥�%��W@�a!h��2_r�uv>�������F<\���UƟ�[�%����M�N[��DVF-U��m��n�ʀ,���z}H�'��h�P穥D�4Ź����P���y���ϊ�%�Q�Kb�]F�Z�`�dL���GC���Aؒ�$_'rW�*�ߢ�6�D:�Į�Ƙ�����uހ��by��V���\j;�����ca���٬��U]U��1 ʸ���\����t�;s����[��\Ґ��48cg��H!��<��,W��F���⅍�R{>�%f�M�w��H��?^�rY,Qq�x�4��G&�k����!���V�b��%I'�\o��޿��
���}��0"~�k�7�v��5���޼e�7�uR]�	S�qG	��$3w�KDg�u��>��N�D�y����(p N�G�£ZR{���'>ܗKϔQ�@M#T��S����ԩrMa���nބ�Rs?�?_f#��|=�\��آ,k{��=%�N��`1���?�I��3���E��3��S�43��#`���MQ�H{�8������裞��H�::��\Pt�rN����_"��(`A�h?�-@J��mF�I�KW��,IA���8�Ϯ[���-���~�X$���:�gEa��yN�<����㖅�@�Q���݅�j����'i(�U�iN�=$�ޜ��˘����#a8FVyn ��15y�\,�K��+��wl�m[��S�� 4�z��p���w��;iʻZQ����X���b�K�(c���b�m�QZ����$?zo6#�C��#4�[M��"o���w֝��h�,�Q�$(�/[���KWl\R�@���.\����4ԋ#+/�S{۳)�����ʢ<�v��T��f�N
��t(��||���c�����=����#�VE�����@�Y����``��vJ�IǏLw��Ţp��_X_���*/x�#֕�=g�n�5`�K|I�Ǌ�#v:1K�&(�S��h[�#�� �O�i�Y���-"���"��S�Z�-+L����e@# ���y]X"���������"me"�1���)i�+���H��uo|<VĠ�����pg��	&�l�w��(UFH��WA��t���N�I��Q��"ڊ��W�2�`�W3V$���#gN�E=��ahQ&r;*��#��LB�[w��S�>%����](��ϋ���Qh�Z��4�W����ۛ����L}&�un�"�y7��s7Y�&��tQ3�W�͏���Ph2� �Mn	|r����aO�*��>)�.j~�Wk�>�zx�]���7�c
	G��Uj�W��TH&�F�l��Iȇu�V=�0�*�5����N��9V�P�q�	�4�'�� �uT�I�����Ј�}f�'��=!��P���7����Q���yA��)ˍ���MT��k�#Uŭ��2��G�I86��� c���"&7�7>o������3�z��(�7!�D,��(	�c���|���G�5bxqEfC"|H� �� 2T�m<�H�wQ`x�}�l�����i�*_����.�f�/;\�Ď�����X��$����^�yy����]����F9���)�Y��|ldAwOC��R<h����F�,�KK/�e�>u}?���Zt�q=4�k�Ss�˵�=}/*R��}!N|��稿��m��~#O��z���	ށ����cI�c൱�`dVM95���Ō���M�q=:���i��+_o荙�����L��P��h�+�� Њ�h5��� .%�ҎG}����M�u	���x�f��N_��sp%Yt�r�h�Cfߨ�z�����3"�k�2x��^��EQ��#\��K�J��yׄl�CL�T��:�s$�6�v�"IK�Y�E�Hۋ�C�A��?,P����S)��;ѵ�Ȯ�N#[�FW��aW����KTXd�8a�|Q�3��lg $����#y��ʒ��F �;����N:,��-��m�QG�2�}��j�T���+�ㇼRNr��H�i"�Dg^o��߁�����6�YbU��Q�X���]C��.�]���}���R�q��L��Uփ�=��^�9I��%5O��)�%9eC������6/����-G!��3:���pN'�_V=euN(_I��9:�����[���s�D������S��H�N��v2-g&����\��`V#�_�^��l8�-�f�� " �f��	��x�@l�O�g�XF?��Q��S�A��;`%�#�K��BȽ��E��燳Z�*�X7�������"FJ�mR�Mf��bmm+qI�ǙIv���<��+.�У��I�cS�ɀס	_A�A1�\�É��x]��G��8C�W1�*�sa�����(�Pث��3�����m���>Xd��%Mc�,���>i�z�UELc6:�q6.��G�NDM�T�L��o}�|:,�=^����?B�7K����'Ce ��9i�/�	r�ͣ�`�W��@ⶩy��Y��`l�g�MӦ�O�X6�~>�Mby����:ńq���O��j��Dp#a�L��Dz�ţ+	F��fN 8���*��d4�=7�+f���|4���l31#eJJ5��0X��s�',�DLZ��6.�QUo���jJ��髗7;t�	/0I�. 4ĸ�����G�<B,d��у��"'���9
6���t0�)�:*��$X�i�
=���N��6I�/�Zh�X1��@Y쇏���B�&,:��>v�%y�|��=j����Z��+x>��W�־c	{��z'�ڦ\�~e��`1�M�~"�:�ݒP!��١�{����t�3�?�f?�y��p����fx����O������w���b+�f���]�E%9K��
p�����Ș6;=�M߽0|�o���׋��N��n�	�0S'v{�	8�򙐲�d`�'�s!lHX�=5�BMQ��MN��5)�2Ĕ�j��A	�P��".�H�r�A�>{�/�o0�����DdJ�[����A�sC��1��f_��x�2�$Ýc%Z?��i�d����ݶ�s�9UYceh�íC�L�^��މ�_~O)���ȻK�����I�9�N5�o���w�0����_�I?lbfp�v�M@������D�,�����	�;��s�\ȃ�rRTF_jي٢^����׏�eeb<�-����b���J���t��ߟ(��@3e�e�ޢ�pH���bt�U=�^�>m�e3:q�G��q���|��ن��=�b�Iq�DU
D'l8Y��v���д��\�Y��]�]#�2l/3�����ZM�7���~�kf���P��|A[rY������.�HtH	��R���o`t-��	�'ӹK�.q���2��r��㶕��f����(����N���Y�I�M�k��Tԣ�-[����X�1ih*<z�%��ש�}��ln���<��?�i4��r�x6n>�vN�3k�iCt�=��o	�qe��0�aV�F�է����	ٳ�����3e7����Uhk @��§39�ŷ�R��} ���\��}>/ٷ������ZB7vӓ��f]��r�b�.0h�����B}�a i�T�q*������Gշ?V�C�� 7Zn�э��Ÿ�,�nt�t'�{<�/3
%w�/o�~�P��]h/k%�J�����	�	�����n����μ=�Z2r�;��I�a
t��0B�vr�*b���U��m����m&+I�n��CT�������_�tٲ}��+�]L7�1�g��[��5ߌb!8��-��K���u� ޘ�0=͂�]�P��רy}�ӥ���,1*{G��i�@�9��r3��<�ʭ��J�b� f��W_.�*��Q�G��t,�c�wӻ ���^>������if��~��Y�TlI1O����o���\��d���}��s������\RR5�m�͏�c*�/ʣQ���W���9�9PW@1�r���m�|:���_� f�R���qz ��}�&e����Ap2q�a�s���b�lO���[��@�쓈���F�|O���>���*�0������릭�?�$�AS(��4o��=%8,"lٽi�Q��'���k�^nʆ1Y����_�N��8����]3���;����$.ɴ��цE5Q��do2.B~x�'߰1�z��'@�^V�M�E`�$Z.׊@�� �O�H�����JN^M	��छx$�E��Ĳ��jPu$`�����~�F�9�A��c�-��� �
���a
�������9P-O:��Rg1Z3�P�O5G�� �u��C����`^��ҫ��U+�
9�~0��X=t��?��cP<6���&� ����8���!���e' z�����nK(�̧j��_�Q'+J���<�}����1�����<�K~�_�s��f�����{�v-�Zo�ް��_d�	׾���23�T��ݬ�Pn[��M�zrw�D=�9�s��
>��m/n�����ׅ����Є
��i����B��`覅iMbH�w���M����w��0�g�������������Z��-.Ӡ��":�I{3�K@(�t��3�w��l������^� ����V�VM�����e=�gS�yh�p>�U�,�/*C�K�i�����7���_7���B#��p����꫕H|5jݏlu���K������^�FA�	Ni:Q�lTp��l����/�mұVb��(a�֜�<���@8�=���m�{�x'��y�U�Ќt0��B���c���`��e3�(j̃����2��������~���OG�)v���DO������-n��Y��rJ��Oqq���9y�q+�ǡ�^�
RT��&Q%Fv���ϗs���I.@cz'�F�m�(�'pcĦ׈f�'��Fɢ����n�7������)�*�`����R�0eK+\L�c5M���-bfo�%��Dm�;��II4����o�f�@�9i��n���ˤȼ���ջǠ���奡�8����S:u�s�b��d��r$��)0/.��K���:���>� ��
9�SH���	��1s��L��D@y�b����}o:��t���U�Hv�F�$v�Q�/	&��I�?�PlF�E�*��m	o�˂���u:ǱY%qR��n�(�rr|˸��o�%z\���y<��n�R����DY��h����Ƌ*���Z�M��prU/��-��\�5�^,�.���H�s�D��ص�Ób"�Y������@`�����9]ų4�-<�dU�br^׷�M2�8N��Dx�x�*���%���	�B<2Պѡ#�&�PjX�%� ~O�b���[r�;Jy2��٢��`��gVT!D�ѿ��w_�%\��R�i��M8�Ý���/�Pa޹�śb��V`�u�{ࡌGc��Ky��ece�wS@i�Ax�c����%a �t�	s��y����4������ h���v��Iڝ�n��O�	��Y�S���pr��c�|��b�Q�!nnE%fr>ͲH���x>��
��y�5@�K�=�9�h��Ra�i¨��5(?j���;��ZnȒH���.���$2�R�	k$Kfo��6�ez�dHb�@=����<�f�E<�C�y��Mk�C�	�{���u��!���7/���@�ppS�,+�QY�8����Q���S����?����8�3�[�Ռ��@���������|�<�i�\>���*2����Kӽy���×K��M)z2�Վ(���9c>pg�U�I^x�-����$�4SE�����*;C ��@F:�*��$�'P�v%��8̢�~�s���&�\Mk{1"��k�oL=)�e���W�>_=BX
b��R	����ud[��o2a�EN4�(ہ�����@#OA�Zx�,�d��J�|�Hd�lzQ�!��8�aW�3]����5���������>mL�T���o�.(�Fǲ46& �Q�g��A���./�qoW'p]�H�h�-��?s���z�M��8/�A���oD=�4Xc2(#�tA�פ(��PK���(x>�K�jųe}G&��!W�ιeY�ڧNŒF�����P��r��4��"\q��.
����CK��w.�m�@6
�ѡ"�Y4���Q��t�}݃��V�����~I`�,+1�>��L�4�ا��W�.+���*�9�I�����CU!f��m_�Y��P_AU�@K��{���W��TB�d|�T֋��&\^s8o5���P�z}�{�9P`_F�Wr0�Lz�6���6h�m1md� E������@��U�v�{��W����7$���Y�Z:�]�OG1� �Bk[ݭ��o�A�׼�lp��¾[�el[�#T4ʽM���`3Z�	,���q8�T2���X�S�X�@G~
���A���n斑��MW��n�g����m.o��bI`���KNs��(&�m����L��6�B*l(�E��~��Zew��l� ��������0Caa�$�8�'�r�&Ʈ���|��i�3����D��������.hlJ(�1�]a�ꌐ��e��~�D�*��fu���ϑX�	��F�HK�I6KcnP�P��2�h(�7�~�2r�(y��?c|�B�F�om-���U
!lȇ;�To��׾"i��]�f9z�Q�*Gw*m����2Ȃ��S)dJA��y�w����\��y�qV[�A�âU#A�=�s�hc&]�k�Rz��9��9�G;�c�R����r�Vx�Tb�(���O~8��/�����^��ƥ�mCȯ.�CWEǯ��7� �Y�9�p3�����ST4CP�ΦPh�"�?��dF�-���X
��ߎ��+�Ddh%'B\ߎO���l�C2$&)SS1�8zMQ�����-�'L�#Uh��1���7]��`ү���C��n(�E�xY��	���,@�>X5���NKj�@��d~*/�&��D�8�/�<��j�O#�?�Ʈ�������Z�L��,�v��9��������|
;4x�l��&�M�@�d�P��D�g-�Bx���_%���mdg�DL,�z������2;FʍF�	�hrv��r������V̡}�\��^�V�z�G��:ŧ�y?��߻���B�S'2!?yd����LSiI�Ƣ	G�����2�Oy��@����B�Q����Z9��|�8�K�U:��x�I@>u����^�a���Q��T7VHM�.���q|��z<	���l3'��,�r�`QǊ���mx>I�g+W�R�h~\<��j]h���������&�kK��1���v�c9�֕e�h�An.�[�&�?)@ޗ���Wu��{�	�҈34e��ϝH$�b=I3ԙ�{*��`ĺ�A����g���f���y�}nՋ(&.��S���=�]B��Ŭ�k�p��S�������� v\��� �'	nE
�W���u<_������ȝ߮�C�ߡ�O���2�&��Uq3���u��ƺ<������H�Au谼bK�9�d�f�mm��O���o*"��w�C�r#��bG{�J��<�Gh�s�w֞dY-�\S��!|�L�#�_2���_��V�ٱvifgU��J��w��k��rȕ�ԑ���uPl%�����0�F�$t�b�QJi��,�h��7�vae+J�{��� �p��o:���r��A���)h����n�	tv�j��}d]&m�<N�~�uŌ�.`��Q��i1ρ}c3`՚+5�muv*Ȫ�H�L�ϖ+&�G�6�L�!g�F�R$�X�m[8]U���}m�>S{^���F������k*�C	�uA3�]`}��,�	�W ��A\9��1�7Y��.��S�Hґ�M_k�oK��*��+@;B�*+��Щc�{��-$��/PZ�Sk]F�\�O-'�BaD9a���N�3*��g�;�:�����06n���
b����W7����ݍ����7"�������������
�!��K���+��f�tx��a|U�|���K/]��K���s��
��_U�-�*���y���f�X��.��6o�V_,�r���^��}����D�����+ˎjr�4e�2��]ё�� 6'�il�+{���Xf�H⾎ځ�E�����H��\d��e� ���-����#"��C�uyF�_���w�����@NT,�`Bk�Ej�Ѩ%��ȝ�cJ��.����9!�}��ݥ�bH�-�*�<�8� �����g����7������RAO�:����)k+bc�u:��st-�����E�?��
Zoӵ�6�{6�ts���}��I�<��`8	&_ϟ���Ѷ�[����	�b�v@5)e"e�N.�k��ؠ��F�3��;΄���w|�h��I�!�x���CY�p����U}��@���^H����\6�4n��z����q�-L����jY�d���+��n�Pd��~e�~m�rT�OLL��/�� �$�"��*�sPg�jBeH���a�T�##NGB���uc��^���x��	�\!j�g�s�`čj�"S�������Q�)�|)�\��vn ��ϭ�#G@]��#ܺp��D��U�Yq{I����������c�kR�,0��>���Ϳ���2v6�%���&����?�f�4���2
8['\{,e}�yK�(ʲ��A�~����ҩ�l��-Q�X��%��w���7X�o8u�_�E�A�kZX�{X\������G:���ްi�+Z������
�l��r�M*M&��xI;}�-�y��7sZ'}��Wa?�h:�;*����M��e
�Jهizח����&�����)�$�q��&B�5(���,h�����^���@�B�S's�>1[Z�5���Z
�6p��a��N��g������z]�x��}�-1�j�����H1cG�$4%��̃��\���c�#S�W%�!���ӝ�@�v8^�-&������\)r�1%��H0~N�g���
)�C(����>j�Ϳt��@)�w@����@���c6{f�zI�v+>�{��� ]�e.�������ҽw+��(�ۢnj;.����փ��,�ZdDȹJ�~�n,-0ǖ�������t�k���|�����b=4��b"�?��|W��!�}���"�G�A�/����L�M�����K��p���!�iY�,�MO��ӵ�����zx\߽o���_z����*�2sWa����c�HVE�fbA��~I�\�/z��gy��-L���ЉW�M�j�8��c�~��/
L�͔���ہ��9�8�r���CZ<"�h<ܓ��G0�V}'��z:ך#F"��8��Ͻ�����0�q`= �G��S>ÞF�d$�i�GJ��.I6шIB�;|���F���6�ʣ�n���'��計�;/3G:�,_� 8��$�k�eE��a\;#�ظ�BlP��v^+��Ń�|��w�'�r����k���h]�X�Oʲ2ݳ�zRB�L�k����S�f��o%i�Ыy����O�O�fNݱ�����e��4�6��6��U���|�K�(a��E�ב�~�G���U���AjnY�y�^�+�;\��mK�"Wq|dͦ�ekX�`X���I�^ugM���v�Ϗ�_�*�F
T\Rk�2:m��I�@r�Zd�'��Գ��
]P��e���h)�Dy1C&�s��$�V��x�>΍�c��s������A�k|l��T��ZaT��9����� !g�藘��E�kjN��-���+*������n�ؖ��R�r�����\Z���P,��Z~�F�}��f���O͗]0����� �f�g�V䅛�?��Uq��z0la�
K��grw-�h��qN��r8�߸��=�ܔم�1�b	!��3���W
`���/������x�Q�rv��e��'�X��Z}���B`b`�u�ʯ���)aFT JB����_��R{��4�Ҷ��UmZ����L�<zKL�N%��
�x>yے��(�T'N%�PD9�˽bBw�J���b��'��P6P5iص!c�8�i��j���	Ѵ�/���� &b�P#�]����C����-��s�p�R�v�Ŀ��)4yd��AK�\��=j��y�K�F��姭�
�Xk���-8䆢v͋�v�����s}��s1�$&�2�,�n�����a-F��7q]m���r{���Ca���=��OϘ�fD���2-[9�?�X(`���hP�%�K�pEî4��u/Q����޵Iū/�uJ<R���v�����{#V�D�D����RT��s�;�'+RhpYX��K���"[���s(׹�F�GҔDͧuh/0u5�7sx]��&>�8G�'GJ�d�c���|>k�FU��l@g��e*��I"y[V���ϙy.��Cb�h�������͕"�0���j�l�7e�9 $�2����LO�q��}z�#Ft�F5�bJBH���6�Cjb��z1��P��ԫm9��;�4ؚ��<�{$w��v��&��uzl�� �������7�v�� ��'������Q����}�s��ߚ�c�,@Bx�V�;��lZc�����VW���ۇYG���CbW�nTS6���#'��I0B���*e�)�pJb���qQ>��)Ƿ��(*iOftwJLY���7|V�����7�_��:i�߅�z���mY4y��%��G��^�Ŧ���G���9�Ǻ������:�-�F����潗��t�;M`����wd����(�qτ��~��_�������q��@�w��^�[�p/��4qH��cf�a�v�>���y���8|&5�}$��MT�Or;&� �(i��+���:��b�*�͹�P���/�+�oA�'�����-�>��Ҧrf��-�*�4�9�VI%*��E�`�o�$�wA�sҮ��@1ЪΏj���%~�'�eqU���إ\Sp?לJ�b �W�ߨ��������'J����H�-T�`pP
� O����Qu�Ww�i�!�����ꭒ�uw��tL�U�5��up i5����RF�����T�� 	��"3s�uE��r1c��E��3ż�f���j�Mgқ���#!��+�')�W��r�a]h�?��9=��Nl��C�F��
|B�6���gaE���wE�G�r]�/�G�|���^cБ�X|u�)k���inz��� b�sqfH�!�M��p�0i�)rcI���m-�u8�&���'U�SW�3��6N��H�ż�,B�����#)�tnӐ�?��.�H!8���	f�=��Hw�O�\��z>�֍{�d �V20��m�e��
���}OH�h���a�I���'��<�!�
��ko�����
vN�@�|{�PD�L�+�hW�"������㹳�u�Ac!K�]���Ccc"�J�40G{��Q=�)ɛs����)Ky�k��d�YMe�=��-���/�fLB��Ti�$H�����u��pމn����c.��h���oPU����[��UiFXx�mG�A��!��me���L &єq"�at6��HU4�s}�x���%/��O��R��r�nysJ���G�<���	�'/@I��<8��u�ND���L�g����q<�㾿g�4|���O׮�5(���CZ��iG�寷,�`~�����W��v���z�h��&���o���[$���s�b:i�D�N�y���>�=Ɵ�eLV�(E��H>t8*r��<o%A3	�"w�hgK�UA+±}���m���R����;W��z*iͬ�'��V& +H/�
٨d�Q�-��a�&�}�_�_@�$b=��-�V���g4c��=����"ɨa�Ƴ�S����*�Vը9a,�9������Wj��TeY2�#7Z;#������'�s�RuӨj20���&�����H>�r��KMԖ?� 2�h���Є�/�5����� g��/�vV��`���Q2�f��5�s�>�[��ݸ���e�˥�:�}�y�t�SP${��RN'9p�a�
+|��f]T��`@�� �z���Hm<SP��1��t��׆(��z��M����[�ZH`Ca<]�?G�W��`�-�yd���h���_������fעn�.�	�݄�
�2jFq�fz*��{H��Z+�g*��c6H2��tL�RuݍW?GۻQ0=�[s&���Ff�w�����f���^�P)v������!��o�>n����=)uл�����k^��Nx������]����&�f۶t�R�q�f�[B�����j�uF=�����v�4.o��[5�:/�D�/
%��ٚ���!�L���68_-R�6�n� ��yE'<W����Y1�5�F��ۣ�);ArWj(B�H�ٷR%彂��z��.�!�܂���ES�jcH�'�6N�٬�M�|�הV��%��� �7 2�3�0pv=���o��Q�/��!T�,�itz��#X'����e��ί��="��I=�)�ݵV!���c{#a�ly���C[�?j��,���_q��y�2~�r<�:�{Z"�O�n�	�
�}P��V"�d�"��!8J/(�E�L�X����y��%���B�M�8����l[��!z��]�Z@$��<P}���#ju��|�{9v�;?��/>�(A��Η�a�lI��t<��À�K�J
3 ��M�
�Ѫ�� 5�׷�p�-������#��T�����x���z�J����_����=T��u1t������N�|w���!m'" �K�V)��G�1�yv�c�
��i�o.l�ڹM���CD����8��kb�]��ݗ-�<c�(Gc�Y�6�F>`Ҭ���M�
�&�N� jhx8W�`T])�����>o�Q�+������a��Q;]�o�q��������M����?J�=_�ϕAyo��+�l1ٜg�K ���]~��#5U�`)��V��e���@2����P�[��Tᎃy-^q6�d��\��M�S^�/��v/������5��J%����HcAE���!Yz
�h&����'QA:�g	w��~�='bj$ ^Aqԛ�y��4V��+���Z	��aI�9�C�[R)a�XƲɌ��S���ٍoЌ��k5d�j!�A�3��q�p@�lwP5ǩCu&&���Z�uk�[�\ro�ފ�׊�b�0
��lCj�Gx�=���O4X�pd��d��z��@��f��Rd��� 6�ں�_W(�@uT-�N���[0l�`u'�W׸m>M��^+(ߵ�Ϗ]9��]���.R�|дe�&8O�w�\���-�p;���=�c� �/�3��Iqe�٫`��u��jV�Mo�����~$�۴�a@��)�C����U��va�����K��P����%���q��k�ZY�/�N�[��Ȇf��O�%�;`�^C��5�w/�E�֏��v|��|Z=���9���$y�E����(#�q*�R�w� ��*=~&�y��H?B�*wy:,�sNJ��,��]Z���I�҉�Do��d��K����N	��Pץ�L�͇�����a̡�'r9W��(WcŻJ���WE�+S?4�����QX�<�"��� �o;3�>��"
h����Ȣ��,��P�)��df��[ꎊv�n�̘
=�f��q�J�>h�"^���)A�Ec�ؗ+���+�v����1d��������e5ii��-O>'�=)x�t��׀����KV������Y\�c���~�yޮ��=�v�X����K�E
d�ʆF��"��ı�6p���ǎ09����|���H�� +��A�c41O-�<�l�m�#)��h�E����-�b�O�k��ɴ��5*�!t��D�	k'�:_��{�b��U #9���/�KI�="4���8���Q�9"�=1�p�r���A�aGڜ:3�D�eK����6�QW����X��&:o�}l|;b̥�<U�eV���~ű��R?L��lǢ�+���)(@�SG��eT6`�X]_BkX��mMO�V^�Y*pS��D�����ܲD�k�m���hTj�%���<�K3���o����3��>4��<C��z|5U�ႅcJ����ӭ�*pj��5�+��XfW�o%�����k���A���c�-�4ݦ��������1�������8҅v(IS�hf.�*މ�oa�Nƞ�G�Gş��#�eqy��N�ڞ�*����ǉ/֢���@�Szk��P�"�����\��E�M��le�>%�!0|Q8XE*'?+���|u��R&���Co��)�3�=z��,�6�}6���Z�-�@q{&
��KF� A�zu�Qq����!��Cڶ�{�)�W�@�!�0���rj���
�ޑ�a;����b}s��AѪJl�V���2y7f�A��ٟNc��O��t���G4�e�4Q\���B ['�~�+v�p-t"�o�<��;���d	Y�n�G�ƫ�D���A���S
S^���W$i��w���q�^��WT�4[.� �I,�u�U� ������R[� 3���@�º���ӭ�_P���#�F@rTSҲrY�y4+_"o�2y`��Y-��I`�!��cg�YL�S�A�P�7��l+�Xq��Am��Y��0�s���DR<Siw4��8�KEv<Lv�4��,��:�twR��r� �6`�D��`��;��6�H ]���un�;�Ҝ�ͼ�>�G��:P�����l�[V�:EA��أ�y��t�ܵ��k�/*�߶���	�L�b(������3�XE�o��u#��I{����~��n)��i$�t."�*������Q��j�vR3���nTZ�1���a����ɧ�}ӷ�#&ۊ��k/�m�V}B�q��o�̬ǎ8<&�[�J���Cm���O�" �1Q���K���������e��r�A�z�;J�����R�b��h�w�Q�.�3eR���̲���u���9'�y6`��I���Yp&�'�mș���z�����t�Y`�'J��w�� r����1+�8o���� �8ב$�K���c�G�T��{7����o���������l�S��j����? ���7���]��A�U(N.W9̜|���5Kf�&agQ�R,>��7�2A6
�7�6bdK���Ψ��O�	�A��mf��t?Ɣ]��qw�L'���2G�k9�n��H���n؁=�(�����$ތt�pߗ�L����o�r�i��ȵ��D|��&i5�v~�	��8�M=�%@��B0=�����lO
��3nC�qd� ��j�q���,��٘mmw~����ǂT�&��g��l��^�kk*�(�j�᥇=�����ꉠ|�H�GI~���x(���E��[��T�a��{���<��,�tY4^�a��.�$��
���l�*�!�����<�o���+��$s�\^�^2����剖p�f�x@­Q����6\�ʳ�G���u'���L�"u���Ͽ��r9�kJ�g���j�L�Qc�9}Z�~��=�ia�ڡ���"oO;�a�����P����Q�S�"�l�'�>),V�̌I�qOG��V��4,e,Q���]^��\,��[.Q[���ۥb��m����kL� =��[�8���}h�{���I3��u��F�MoVfp��-7s=P6�,Zg9��XU]E)J/%�Kb��`)���U��������ͭ�Ӧ�u�S��n���b�$��
�D����?���E�M���B6���O�
�����F�=��O��t����.��{|}
75c�n����*�6ޜB�h�,ҵrW������]Bb*m5���0�o�[C����<mũ ����:�	��
Ox�N���t0d�^������b����$��(H�_&�@��a���k�� a(������`����3���ڛU��Q+s_"D+����c��@L���:iA}�����;�T!�����-�%<Y���`�+NG���W0�`��&���g��m?4^�����ގ�� ���c~��mon(��a��' V�n��/��7G�B�W��7�)�Qa�e�.�����Y9��,�Q�����fN��V��j/��޸��g���)�/X����B脅V{��� ���Z�tNI[�&�%�,������&�D��߃��w�F�f� �|�G Z'��/�A�G�� ����e;���^Q`C�;�?[��#���摥"9��<��"x}�K�p"�q�[3df��Q�l�`'��8��ձ~��Pzb����2�C*/��p!.\&�������W3�d҇��L5�FFK>C󷃅n/GO,Yk,S��v�9T�3L��z0������U!E���sO��;�c��a�Խb^�����1�$�R��]	�	8�Og%�Ϯm�k ��}38��RZ*�ү@7���O�ǹ�V�Q��st�X԰���=�oi݈?7͢�����K����GC� ���L�.��.��ײ(���{�B&�֐p�"���#so+Fr&���d�zi©��b��mbÜ��i��b��t��98ϴ�u��li�ب|���$/2"�io�3�
S�m�c2�5�l�����e3�+[\�IG�O+��g� 0��$�>O��U��ĸN]��K�&����uĝ�1|Ex-H+�/V.��(,����g>���6?�w�5������SnzV�R^ ���n�@��*f�D�^�e�j?�,|k�k+�j�)�l�JVX.[�Xt��xL�M"6R��;�NiZHw�-�h
�>\��-�uC�אr��f5Ϻ���%��h�~�<�K};Vq�J��"����Wlh�sV�xΊ�?����Hp��: -�b�b2X��Ty`I�����.w7>����La���X�4�~Y"���1t����@���2��
�֌8\՞�Á�G�^F�P���	�&z�ܧ`�guӗ-�a-�L ����K�ȃsz�%;d��ԩ�߱
��I��A�JoǏ͂c�� ���[_�,Q������]M�)kk�������O~s�/W*j���O���e]���m��!����]��@]7��Y��K-��D0I�7�S��+��2�L(�y�Yt$/m����X�����Q8�*��	u5�>�	�C[��?���n�B�X@��
��((�y������	C���O���J&A��N�z/��e�2�!��^+Ň�N��P�&Ɇ��#̛��s�an�P ��Z7�}��w�>��%@H.�i�����y��2����-uZ5��B؟Nɒ=(�0՟E�d7]+�bROM��?C��x�f�炕�O�w�W��.��t�Y8�u��"�A1�u8�Ζ�u��Z��9�M�U��:�u}����z#tX��0rI��"��n�(��<8l:H�5�n��g�8ZH�d
�_�N7H�;)x=K����%��N04;���&5��~�7^U��k�X��QB���l��+2�B� o	�fB��r��3rqN���U��#]��7e�;u�([b�J Gō��S><\z4�n���Oa��/poΣSl�*�DuB�k����+���q��	��5q�����E7�0#4''��9.e���O�smՌ��J�)�"'���y�v^�+��LK����V�\ ��U~��&3��b:mt�G�F�('�Mwt��\nؑl�y�WԘ�wك���2�i�#��d!�)rpv*���S|=��s+�X�e�xFq����+��w@rd��Gѡ��sG��=�qA*_C�+��W�ql[ ��J���Ò�6��{�'F�y����� w|���I��E"��6r7Z�ƭ�)OL��M-ٵC��DK�/n	��(ԇ�4s�~�U��v裂����a�rx%�V�An�K[���(��XpW<U�'��;:����5��D���{J<^!�J�ӿ�a�B?uJ��K��<�INy�e:
���C�[�f,�Ι'�E;H@�p�5��R_T���D� ��}�c�h�G��]�P��x��I��"g��2i�o�\���R�!.v��쬑?��c�|pM�H�q�v��Òs$]�����>@�����W>w��v2��W���Ë���[�/?�/+���@���IU .+��R�#F�px���WC�������F��W�c��t[����	��j� XyZ(��l`�����ZE8T�l1�"dA�HjH��P��d<{�7AZ��� Y8��S��DG��+N����}�b��W���1�g�غ.�_G>�	�H�i]��Y��5O�H{�,��
U�%#��;%����]����U6J���Vz�$V��<���.�l���Vi	�?3@�j��t�U�7'`��G�i]o�͔�@�>�ž���S�!�����%6��	0Ǭ���^QW����s)}D�����"�T�c_a��nb����ɥ��p�\wBN�"���d���Q-�PNq�����J�T�)�i��k-�ѕ���,��%���
��\Ǭ[�ʹq�R@��?�t�d�ZU̪HbTGn	L`�e�'���=���"��ue�-`�u�H���[$�KK�檛�:��5�)��.�Ԩ=�
;�#7�b��i����-�R$M�o�<ʐ��Cy9���6����?7��8\G���	�	�%�[Z^{�O��s�k�P�cŭ�hL�� R�a��MdJ
d�tm��K�W,��%X� V��"�zg!��`��������d�Q�"]\Ő<J�:�	����J-W�k�|��V�_a��dz����|7۳m.�F�zzh�y�ߩ�`�ё���h=i�{ӣ4����w��p�m��3���s��v|���=��ۇc<�="d�~#?5s(���z����C�����;���D�Nq�\n��ѓ��/����F�a6��I�9	b>R�F��B�z�yt<C�������m�-�	lab�i��ti.G���x�P�����V���%�lP��ኡ�9�˝�w`����ˎ�.��O�R��_� �b&�?B�$v8�b�*��[9�Rz쀷�)�W	t�ֻh�(�w�)��S^Q��B�Qһ�d���"��J�%���a�����\m�e�@�2��Y�
��$��J�~�Lo�w��z]��0I,��z���;B�,ƞ��g��@�i"J��l�6��d�̓�3�"�SO�M����7���JJC�z(�3������NK�q[�	ܕ'%�(H��y �7)-Q�h��[��ߜ�I�G��Uc�_�23�p�g��}�QY�ҺIy�W1��h�^i�� Fu�|���D�`d��I ��C��YV�'
|��H���~ѩC�=O�`FHB:����ta������.>�)�^��%ب�����NH����МFð��b�R�XJ���A��$��)G8��O��t�ˤ5�ܮ�{�$�_	]b�$����aF!v�^�Pũg[���;ʉ�Ε�_T9��qt��	V�`W�?�)��?�ٮei���a4{�i�>g7.�r�S6��}��W��-tp�e=0��b�ЫR4��yJ�w��d��y�Օde��puTjxO��z@\p�6k�j?�G>/A�'��f�� E�6�p<��!�`H�1h�=��p=!�3���Tc9�Ga��@�_����/�O�o$����D�^�Dl��F�L�>&���"����3��71OhE��z�a�q�Ѫ�ʗ��+����J�H�]d=�G�b*ߌ ۇD��7�
%��G�y ����d�>\b��O�u[=ێ�����1}�Ȳ�[[ �/�9�45\D�V�f��R� �mI#L^0T�@Dd��v#�"\�y�o�ȡB$�Pw��4�9{�,�͆9�f��|�I-l��M[|�4��LQ��W��DU��Z�w��E�<�V㒪�/��I��^�N�*���f{���b�i1ozz��Z�*� D�̐29n��-z���ԑlzY<�y����~7�;�kǠ���>e��B�3n��{۹"�87�R~TSU�:,�v#�sO����X]KgQ��u�`U`
b♟9���z�1.�=��c?Q2.��!�r�� 37&�a�<���<�[G؇츾	��#������Q!KP���M/	h-�NQ���\�p'J�B1�9{��c|(�l�������������& ^�$'�r�TY0թq+5�d�Z�L��9K��]�SB|��~e���Z1/)|�q��J{�:�6ƣK'Ε��� ���<ۺ[�5�I������=���k��d ������A�5�կ��D�|J`	Ĩ��;eL���f�=��kAy�q�SFt!$@�`�D-OS�t���}u�IT8���P��IoL��6�.���C��/Vܚ-;;����QB��7ʒP����O#����e~ȅOG9�oQ�l��QI�Q{gK�Y���<�*&�&�R�B�B���>!J����X8��hN�������є�d
������#��k
+0b,��0�8�.�D틐�,7�_����%2������m%��)B_oiUv�F��U��5Kj)����{�gͥW��l/%9Ns$Y��x"�-�W$�N���0e@'��>�+����|�
��on�n{�F��_������M�v��. ���x����B�ٗ�ר�zfz1�@���F����;��p�~�d'*ː��r�c�������(.Ŋ��������}�V
Y?�=�ֆc�THc��8Q�_,��Lϴ@���x��{�+�@�c�5�P��c�u*�$�K� <�[p�� V��\����N&H��r�y���Hz"�0}���C;��l��m]e���_o��FqIok��b ��搄�½�8��"��*ˬk�p{�:r��
��Oe�%�	�+��� ���(��&a���2]$��}k��)J��^7�E����S�L�(&l&s\=�4"sA�����}� �[�kwvn"
���.6�ό:�(j���a_�WZ�,y� �&"P�E0�+�Wj��G��@��SH6E�9���Y߳�T��r�e��$�##[�a$qM��Ow^n1]!-���A1��/�$Z�<��z;�*�`�������I
�#�nHX�a�ޡ,F�,��<�mA7�]@>��h�)MƬ��-��W�}h7��sp��ܭ`u����n	�QW�\h��)0�Ֆ�=CM}�����ub��AD� ���MW�6r�&g�}U; */w�կ�d�6�@�c;���X\�4��o�&T������dl5DFX�o��.����������-0�W�2�up-&�N�}�L��m�ր�P��V��W����A�,�ip���@mK3�d���K!�E}��#6L~���`�_*��Wk;�p�R���C�#+0���pl�}�D*����}��&D�-C7�N�A^+�����r������u�2�Ц�׎N5�|ڸ�<G��6��DO�Ġ��O�$v�����W5\��9�#>x�s��t���K��+�ә=IEW�I����wS�>sN�e��O��nҞ8u�g0�<�1I�C���S�+�������3����--]z.�Rx��Ѧ���\�Yΐ���؋<�ŗO˿��vt���B�1��������<7���β(�.�Y�J��<u�A����K�(`��J��q��i,���2���̢���|�0�)D���B�yn�5�B|p\�l���2��]��� �ө�Б{%*�6�
��B����t	�.Ʊ�q����u���O���ի�b���Ȍ�Cmg,fnHs���U̳�+�xSzd1�倐D��%�U�,�zfSҘ��5v�h���X�"̖�3C-��h�W�{�h����uZ�0��Bd�VZ�{:�MkF|��/���/O�=%�_7�҃����k�A��$�~ڎ����=���(���"a��*�B����Auh���\KMyL��t��LĺG�$��a)��~�P�b�G�<U7+�j�p�!b���!~��~ǂ;�tI�PȈ\*�cZ_��:��&=�|��U^�ƭ�n���l���5��VH�2��6�l�4����&ߖzK�wh<v6惉E��t,�8<h���bLd���q<�՞I��D�ۉ�]+���[�-��:e�e���"������W��v��r;��X>gM{4�j�^�?v͙�j�jq�r�w-}kn�=��u���>P^�eEQ����Zd�K��m��� ����@������*��_�8�h�L�l�았:	�L��V�=��sb�MU��{�f�;T��c�.�臞��@�e"�p��59�V�%��L�OڎS�{F�P	�	uwv�1Ht|џ����M��
p���Z�ׯ���[³�y�k:��Aq����̃|�M�·��:�U%R@G^������o�G�d�~qI�܃E�B8��;F�s�+�c�wQ�t�P�CT��B�m �\�����lָ<|J���=��(�y�(+ˤ?�iNaLj%%� �7�D�!_���������N��+�}�6���ߤ)�aW���)|�/���E�jA�Ӹ*N��N�2S��ur]���=�D�HC��qRFg�mo�A��(n5En��u�*�x-�����mݬ&=산���i;�{d5IU'��xڙ�&��.��?�Ȝ�7������u��}�����f�o���59�51E���3O�wK䆽��u)�H�T@>�>X	�Z���z�����e��
_��� f���A���^�ԉn8Z�_X.5�0nשpM�z�����B�P��Xs��I�'	�׮NZ�X�v:Fiw�����~*��F|���fF��a��L0ҟ�Q����o�7��[^+K� ����g�O �3lm��wzzE��/'�&�����:ൄq�)����dO8����s�.L&�C=�[[5f�>ǀ������-�1��v�R�.�L�'�ylS1{�O�AJk��qI����a�U�:����l����F��J_��c�o�[XIe����X��~�'��Pu�b�sD��������{� �l_��X��'�������?/S~�Ʌb]�����_�k�XH�ec�Mw��E�����0����t�v&���V�P�2������X4�*���<k`Skc���{�,h��MmѤ��% =Y�^��s'E�R�QU(��pK�O�c�j�г����^�è��-4�)����<�ƭ\_2?J�S��[�z$�F�,s�1y݈R�/�����>�@=� ��N��P�pM&�I(��~�@s�Z��D��l��<P���S�qB�B~�\�z�>����k�U�Km�O.������Z�}�vuF�P��Ø)��a���c�2��.J7< {��Y���UO���riP@h.��9Ƽ���2������i�"�F�=��~���jCD��d>��U���@��C�SB��4~�ɖ���vg�;F�Ɩs�/0��7���@�I\n$>��%�4),q��5;h��@�S��2�zd!6*(��3}��f�ݶO��oIî��-���| �����@�I��p�`or�M(���M��3�_���T���,Թf�̈́<9��d�N%�Zd8�3�Z��\[�׬L�b|����4��g�V�Mq�Ӕ#�1��K�k��V9���`L��56^�lg|^��{9 C���P7?��Rd$�-�)2�]0U+6�;v�`}v�^�da���0}�5���_�⢚�㠘����Q��5�[[�o��L��;+����qS��5����ȉ�|˹_
ri��X�V�Q����E4e� O�V7j)2$�N��z�np�W�u5��/[�?���t,����hi�&rD�4�8�8���#��Yo�|w[s��7�:He��m�����l��_n�kMU�<[:8�mX�R�D��<iDRf#]�Н��
q&��7�c��e]Ò��ٲC0���Z��t��YkTc#�$}{b�@1a����=��9U,U����2tF哩C&�����]N��`�c�j���r�O@��-�
Q>ݸ��������M�Q��c�[�������n퍆AF崷�q�u�p��eIxV�����X�uG�VyUq1�{���n���f����� �;h�06s�ཕ����q��Ҁ�wO|�յ�o"��N��EO��ο�o��8���72��PY[#�a�=����X_��~|��6)y��a �):�����gP��!�[`��X�.7m��>�l`%�Y�68�ڏ�ZK�7��)~\{��i��p���M��lP�������_P�8�qW��L��ᳯ��+��@/���G�Moo�<r#��n´	a�f����b`%(�8�`V*����Lf� '_O��jh	��2k,�,�$�7��⑉�3��WW�"u�]�=�V��N��ps���<e�HM��R�x�^h=�>����l��1��?��� ��Q��:jeʗ�j�a:���Ga��RY�S�Y��q��'6J��K�b4�">�AX3Ǩ�I=&a���4?'ȰD�7�P�i6v�K�'F�����Mh�{��d���f1�s� ,9-
B����<��M�Э��?e4n񮭿�]h}�sI���m񏶜�B׷.��6�,,"����{���
��iv+�u_�&Q�fN��W��C9nC7��G�=��t��[R[�RyM7��2�-��
0��������^��l�eSkޠ�d�^�H����ڎ��p&������(L�C���LP�3v��Aq���:�^J>,v�KXq���e�R�>j���Ӎ�)�19�/%�"�-���;�|!u%xB�zV�9��,y#�N`_�I���B�<� ����c�� b[ֵ��3B��65Z����2B��>�%c޾ʧ�=4=r�����3��tZ��ݗ}��6&��r�\��q���͕�]� �ڝ�� ���"��$��g@��¼��GB?1�E2u�K��o0Fo�`n�W�ey�F��+������'�v�5�=��o�sT�mRe�^Pt�l��c�Z'�G,����91�Aaw�fz�������?ct\��@M#�D���	�x��m�YѦk���$�kd��LlVbx�~;L��n���TL,�97�72��qa��	k��c�,���cc�FnM/�q~���jd�G�C���ً�E���b@���9	iY�xjE����=�[�(���f���%&����c�_��P��{�T�uw�}Pb7j�i%)�5�'�B�A��x��ꚋ��X�߁=���v5ބ!�Q�����^(�;2g���@�?}%$IП�ӝp���5�S�y���W��7�T���{�}��J�{�Q�1�����A��j�][��^��u���~��~)*۵��9l��\���(� ¬e������tq�����9��媺��GH
\/fs�k��%dX�U�o
�zs-Ð�m���n�X௎0�ɼ�u��7HAF�

΂��!h��3����>>�@�lG�@�Z�jr2�!S�y����������&�6�K�\��?��vA�ҹ������]���g4��*P��\e��^��Rc1eF.ԑ���Cf���z�˳�2K���
G�T�l�Ђ%ˀ�6����XL�QK+*�Y�	�i�� �э�g5�>K�	��w���YuG�|J�ı'
 +����R$�l�y���������T�Od$6������J�T_)�R�I�COg�i�]�cي7���_���A����隧w�ݚ��|ٱ��.�&�}r{�]�aN��W8�ߴ�uٻ�su���$������(�1�~��ʐP��g�ԩ�L #�� 	٤$�)ߍ�'t�t�Ww��④G^�+��bb�򌕠�C��@Z�[r�K^��>�P��ߴ�<�9V9E���\�6�6���*���QG�����F�4^X6�T��V�����:Ҭ%�����4�_,��qk����H����q*$��L|��@�֍��������`�uUzŧcc��%���0�Ss�Z��ZeUD@�����v��C��|YL����:��^�� h�'p�[	|�AX1B��:�����4��O�r����~�)״�>/�޽���ryEg�/R�3a��%��F�zs�~W�R���S²�N;���O�4�Zp��j�ۈ�����a7a���ˡe�+vHQ,g�P���v�ؖ/_��C�X��l�:UP�jJ��o��xH��c+a�[�����K�� +����=fT�gq�x�Ք���4��L\?/r�ܨ�z1$��{�&��d�a�zp�ˁ�Se�f�k}���<0Q��@�M�����^�k�=���b *���TOԓĂ�ۖy���˰�o��x�0���Z$��~���\�
^�qa�F]��z� ��.	��Ȫ��v�b����,�[�3����7�����'�*uB�3��(:uG�� Ώ����xDq�{j`��>���#B+2 �<К����H��0���58�i�.�7�4Y�����Lԧg���WC�/07A�ztn0��Kpђj��u�?�l�^����D!p�P�.M���r�<s�$����%���V��FD_��,�գ)C��k��w��.4��>t(~��zE<�^�����)D�|�ʇ"WL�����Z[��Vآ��x؃��r���?t��0��6B�X�e`�~��`$X	��wڝ��!N��x2:"����<t�?���"BAizHf��G)[�ˮ�'��7��P���*9g+F�m3�7�hHE~Q�{|`�-!)g���@���4����4$ڻa�� L�rӰa����'�LO%�dZ�
���\�1�����p�R�5�%^���;�Ơ��E�BѬ�g�H&r�G�O�f>7�e{�w료13��Ƿ!�P�¢$��mNS�8�@��L�7���~�����t������&�ӣ�6�K���.i��Ae�s`"��$�M�\�؈d��]�:|KRQ}�̖bL�	�gGck7������-ߣ��4g�`�|��<��/��|JE�����%͔�#JL�V�e9��� �l��Bݺ���CtO�s��{@K>*���W�lZ�=B��nH�V��{5ڒ��)W�?�vT�e�s7ۀ�� ��W�O��`�ʴ�~�a�F/�/�K��"6��2�G�1���Z�<Eü�Y��Q@g3��Fp8��_�6�$sSZBѤ.�������T�DضDbK3ےr/̹�Lax����A�����Ԏ�#�����b�򄒄��P�(���B�n��y�d@�z�R7�#{V����RX;AY%K<����޹&+�������bd`�Q]�-�2�?עmP+�h~�Y�D;��F���� ��"!�[�g��i������!np9���S�ڕj�R��hL�Hrb��ݨ�u���߾�&E��8���r�|(��^�2�l�>�jM�G�F������Q m��@2��r�r�iM��(��y���R	ۉB��>�r��k�UcTK�33i`�)7j<�Q����mI��k��Z�/��Ϙ��A\�
w�iX�eo܍�_d�A�:�_��2h<�h��=�s\p��E����ܥ�� �Gt^�q���������IV�֤��\�A�	r��9��?������獘\BF- `�t������iP��ܠ:�>n�)H�&��&�<N��Iqx?�<� �sb����@Π	�΁1���鋽7?���퇂!�;w�"/�eEL�hs֮QT�y~�.��{�>�<pY\Mp.!�[��[��8�����̓ �۵�ߏ�[{�-����z�N:e;D5P7����J��R�H����<U]��($�ӈ�1ޮeF�E���J�i���GR◎�r�h�*����U�9���Sq`�e��u��82`���p����l_���ä�~�m����F��D�~A��.��Ξ\)�rv�qa��9���4%Ûxm���f�m�r�߳x�ғ���'w@M�:U��V�[����b�8� �hm�lV҄}jkq�\P��\���v�h���V�)�L��ǌ	X���3���"l	D`SS�y�J���� :����Р��&��v6<�m�db��#-杚Mm������p1hVp� m���c��!�'a���/2Xm�[��M���!��t��vJJ^m�-,cl�Y���n>�٢���Ʀ�O�~q�Xҳ�Jc]	I�O��;��������gq0S!�u�^K5m��TM3A�V9�Q�	�\[�ޝ����&��ȧ�2!T+�2k�at��hZ/�3�ؚɰ��2Q�\:������94�p��x���8����g�"R���D���,k�����Ejr���H̔B�%g�D)�r3�E��!���>l���D2�a�^�����j
���I"M�G���(52+�u���~@$�b�gv�OƎB=���奋o@����NC���\\�'��Z� ��7�*�U�g�K"��y�]Ơ�qYBȘ��	��=�"F'(�ģٸ����Q���>�?���&�9��Z�v�k���ۍ�~K�u�{K�؇����/��2�@�3���l8^�\W�� �Î`è�6ts���Z���B�v�5	�+���/�J���B�d@�4���N����l)�G�tٳtj���y��4��i#e�<���I?�%%#�I�Aq!ζ�D�o�F�IB���c� �QaP:���N*�o:R�� ן������:��I
�q����i��!�Z� ��U��'a����W�@[:N��1�9�n�˨�`G٠Y+��q�?�~Ω�z6ނ���#a��Y��j#4�~���TGX3������><`�U/m_�����gM�WҀ"���V QE��O�V��1���'G�;2`�Vփ*w��nln�z'��n��-����+�]�S_/�����$��-h�[s|X�tI����;DE]�s����3�g,��(.�����)�ů�ks��])v���v�C�j��a�� ���ވV��
�;gJ��?���<�W�&sa��{E�������,7R`U'�4e�[v��ܼI�S����q�m�]�EY�i%tԔ}��v�����y���g=ajF���(��t�?�=��F�{�\f������9+�Y�o��^��Z�a����9V5֌�l�'q��(c�妐�Ƶ筟:���/����_+a�]�:7Mx��2&}���,��T�A�JW� �bJk�F�=2���f���&g�e����>}bJ_95���r;F�ň� 3���>m�6���%����4�����#��N�`�O:������$y��]�fQ���l��pF�͌�ˍ&8���yP8�GT#��ӟ�ƭ5r�^C�3*< �Y�2պ��D1I*T9Y� �������z��%Q���~�~)q�ɧ~U�<=����E��y���~��݊�T�H!5�~m�،k�Uw����+��yV�Aw>��]WE��P�U�w�_��/�9���溜i~\g@����Y��5Q������=X�6��hY��R�[���+	�J3���jT��(��D�8��KG���:9��3ӡqG�e��WIC�
�ek*�{���2�x
A����C=%��~c�2���Xe<�o;��v����"˗����@O�mp���=�_�tփU�%��?��n�*�����	C�;�)��k�JbK��x.kO 7��c��g`�S�z�Ut����>6Ob�B����:����yX����V��:A�6���m�>b��Q��t��>\A�����G�L�-tґ�]�g�� E���/���k�=N^i4�	����{���Ȑ���'5�Q!:����K݇���M�A
�P�_�4�_P��T;�#�F���1��8!j&� �G�Us7�XP��1�*�6�81B�'lI���k�W%�����
�m[���uWq%r�K՗͍!dsz���gڊ-���N�֯�(l�v6	|��B�$�d����.5I�U-ſ��-����g�9���ֳ/7^���u�YS�Q#c�Ȉ�G��@�F?�)0mq�
�!Uf���WӛЊ��ۄ7�#�T�,Dh�,^��r ���"-��{�h2j�/��Q��ݩ����/= =��d����u�:J��OIW.��
�E'�;'|��À�f��s�3�$��5O�{�?h\@!��{�[ݼ�_T:T��g�b9��u@�Mz�8���q�� =,�Ô��?��Cs�O�Iv��m�\�?�ޓ���o"�I�Mb�`�	�"��l��4�����
�%&L�Ii��P.Y�yxi-��)Y�z��xst7��9݃z����m��"�Ρ�M$�}�V�� �x����o��`=������T��Q	
�0Z�@.j���C{_}�ؔ����E��$�f0�D�7ka6�#LD��>J_�h�1m"���[��Ui��D��ms���S�<	W�I�ꏁ�kOW��v�R��G@�����v�t��	MB��Ԗ"'�Ms�"ƾSr)���)%=A~R,J� ��i��)�(���,X��_�8�I�s!����kֵ4E�_a�3,��gJ�(��l��U��<�F�����/��2c�m��6�p�)"b�n�'Nz�:��P�Zi�d����/=:�/׶
��3���Rn�ʡG��ȷ�o�W���r_��e11fN�)%����!x)��.Vz0Ч�EHa��P�*�t��s��M��[��%��F�\p�n�V�B�=�a��]}p`���99�4\�=[i�@?�.�)[<�����?���.lсh��ԉ2�i�9+\v^d=�%�A�VD�P�U?����	�>��/9��@�E��-5���'���-b0����CT���_�����x}�db3�6��r�G����z'=���+Yhs��z$2��U��LV_#�%�v�qy�f�T
�F��ރ5���~c$M��ڇ}�D��w�g�"{������0!P��_����.�L����� |Q�W��-uܜ�-�v���Jy��B�7�0�~q3C���)~��T<��d�¿��>�9F�����U'���݅A� oj*�ulZ=���_.�O �즐i�IeK���kڊ��Rړ�T6ꡆ�������O���K�A�ILF�.N�9�ͮ��~�y���I��pVF9^�G����N1�t��vd��,C�E� pL'����+8I�I(��rWZm�����;��K*��1�P]^�"G`��L��I�\a��F�x�PZW+�'�42W���Սa�p�w��tN���2���l�Fe?���ϔS�`��+�����®@�@`��8T��Y���^Ѣ���H�q�cf}w�Q�~n�Xvb:Ln�>����9��vGM΋G��6�m�>�ܤ�d(��\5.����K�j�"	����Դ���^z�(��/#O���w1���:�����J������N�@w�.�h���휩��w���7*�Hӷׇ�A�g\dіթ���\^�a`Ӯ�=]���!���^g��hŰHb��	)���,W����GfE�t`�"i�-��-.w���O�7�����|v/�6�4v�l���t�yg� �*��"�B"_OqXfn�+bE���78殙�!gv8�������ި�J#�!q�Y��!b�'>�S��,���hr�V7$/1��Eh7�+�7A����
�����B~|����FUd;�wf��#	����
�a��p���? sE��q°�*�g)&m6QO�0��M'�wࢼ�S�v�[`}1O3�dC�A(�Hڪ�vƲ5�g�mo3�3���T��9��IӃ>�^�����D�x}w�
��n��J:��*(�&�����ܘD���N���]w���V��0��PM�C
KC��;�NfB�2�)��C���O���?���h�����,�	� g݅"���V_l4�x~b���N�n�g^KU>�o��~�*��k��Tr�I�X@f��-e�-<�����^o���c*ѥؽ�u8�l���}�v'&>��@bO��w)�T@?r���ǺB7��uC�V�@�Z*��q�)�97�7��^�	X�Ǣ��{m|��d��M�S��*��։���ރg���Ċ�F�ت�����W��������eY{޼͡Yȶ����;qt�����.<��}�w���o��mwA�[�`������YO�Z�L^7��o�@Z��tlf(��Y�������MI^�WV��]�F#\�k�m�Z����a�
Ɛ������n��bN��U�m�z
�2��9�a`�ƨ��K��j����F�g��R�qXOK�ب�b��ĺ�36��������kW�XQ족N�I׀}� �̿��d,��w�ƥ1��!����@�����..?߷_�Q�H���ec2�w-��J\vR3����XVg�a�`� ��df1�������os#(��/4��t���y�\�`�
�gm����[��b�"���!`G��r���eI�#�&������|�&�)�7Ğ�<�d�"�z�[E�0 ݿ��1��}�%�o
����)S�}@�F^�Z7��YZ���C�h�=;��TI]�\9
�t:/?xp�a�����y"gu�t���w?Z�ص�Ob8�����+V6�,Fp�����\�����lȋv'{��3/ ��&�����-�#�n�B��j��P���^АB8�B"�%�̊���
ܠH�����ÿ�	�6X|���r�ïfY��0��i�s����t#�&�lU�����w�衰�C�]_�Bt؃0��~�Lt��{E���0�AX%�+ho�F�c��� ��pN`���M-���l���z��7Y�+@\�b��$�l�G,٦<�E<���0��²"&��+9����^0�^��J��Kg}���a^��Kf#�6%>ɆȆ89��\_�Z`��>�P2�^�Ғ�_)�A�l�M0Y��ұS�����~�q L	�p@��I����L|J*�U���t)����ꀴռ��A�xe����z���kdM�������qCL����M��v�)Hھ;Ȟ���9�㬅����L�<8�;>£�P�%f
N!pf���O�"������!�n��'֐k3^D�'L�AAo���DCG_�}E8���Y�,����e��j������V���Df,��d���h �GA9�~����_A�qVo�j���C�����2b�V��q�����ػJ̘�S�5�B���4X�8�����<�Ax���Q>W������6�E�y�J�����/�5��Z�f}�;� �|�ڕ�V$2\�wfƫ:�=7�J'S�)ik�~� q��j�}/��6��1��a\YRg3m�؄����CSQwf�pӞm��:)�X�%�Ɣ#J)�O�-LqX�ũ����b��ޥ���t��S��#rdrs��*zvI���ud�?Ú�'.{�\��S'��a7��4M/4�Գ9o*��6<nAQ����R�U�twJ>rk�8@�H��~�rrs[b�1�>V������?��_�`9>;޹$���R>�˦m�!�)�UT�d��k �+Ʋ����h����̀g�t�f����֗G�7�_�̫���R�g���L�������3\���73w�w=��]�~�Lo:���W� ׭���ڳ�O&Whx�t<�AJ�������k������k���Y9�-Rs�f�_`�|S�M��ǚ=˰��@`�F�	Fh�9]��7��
�0Y��r���rӑ�����'�֢O/�'�5�ԅ�&r�g=\�X:�­� �{�Zj���+6X�>HLA}1P�!a��x7�`��j��j'��}؋r�A�w�?�Y0��K�����-&"Ze��_I�'܅��ϒybf3]���X�! K�n�:�H��*��G���w�FP�{j�( �g	��t[��E'�+|����ч�)�F�3���&�T���rB�@eХŘ�|�4f�I+GNhː��� ����7�GIoK��"E�@��{�[��Z�A���+l<*���d?D�e�_j����:j�gUoIQ:&�>��}��|�!T�{v파M��jjN�B.�q�)�)岛����	3��t��^%���m�GV��9��E&���e��/��w�n��ԏ��lԅ�ܽ;�2��a;	���j��4�O�T�MW�)��FD6�\K�������r�	��~��C��U+�r�NJ��;�Ѳ�2�I�1`��S�(��,�`�L{sL1��]�VSn��hx��^��b� �)fҸ޽���;�Jt"��Ҟ����!�-�lZ 2�g�j���#�A�u���+Q��O����t�*;�(���#@�������@R
����`|��k�&�(�Dci�f	޷I�������=S��T5Q7��f��]�Uε�I�f����6��q<��?8:j<A�d{�](K���3��h�j��R � ��c��l�� �.ۡ��^�t����fI���F������Gڹ��7�m���H��/mɈS�ۉ#o���]V�C�"���ɥ���MD	��Y���xs�%/}�q�&7���~k꯫N�Fa�-I{��S7�?��s��Ը�&L�#��m\GQ�{:߰�4�!Z�:m#,���V2&�;����EJ�p�.���wI��}Rt1V��w�z,����Ae��h\{�]F�+T�&����uvb��4�&3
��m��~� ��c&�|B�1?B0EV����F�ө58o6���:�����ƀW��p�3T���ۆet�$���N��u�9�JNA�g3���[r
��5��[�I�C�xs0�F��X���f�� �|v�`ѣ���Mb�>z�S��9)�ɾ��a����Ϻ��
5�˸`y7�	�'���U�`$���Wc�Yz�B0ٻ4�#\�]���b.��'�Gn]���C��O�$A4.�1��]-���ac��]p�^މuo�^����Y��t��H2�Cܫa�7d}��`ے7BB/ػ��e!z��Q_Km���r�7�dK(iصp`X�I���,�B�6k���C���c�y M=���e%�`^���C�V�����&�c磣�d��,#v�ve��e�O��޽���c�Α��quk�3+䵶�*��d� m �fμ3�/JHh�ZN�X�{qx���|r�!(�!����>#J��{�`TYG��
�"��� 2I��>)Ju�yc�Yd{W�������H��w�v�"�i�d�����턓��&��lU�^��L�
��?����PI����5�.�%Ujl�B�M�#E�'5g��.C���`i#��Ŕ��!I;���P��>���%n*/9}h��޷� 9�S���38�b������xb1f;<
���UU�O��eŐC91�v�f83�<�)d���V�n���H��>�0�g���G�{}���:}�K[;��ɚ��C����1C�	�^qhr7,�z�(	'�������|���jO���9�[��G�)P���A��s�Q�eV=��i)(Ng��ɽ�¿��[[��C��(|�FV�Y!���_}�>$0x�)b#����<��s��_��d��}�5��䌈f��f:Ŷ�X�P�%�Nv��X�:��O�Y��mǲE�x�������(&v�eZ�ֺ�y�L($^G��f���+o�C �ŷ��}�V���6�T3p1S�/ߌ�ѭ�i[w C���Pd½��y�j���/�֛�s�	���Xh��[&~kD�4���\�������ҧ�}�i9@�X���G&ii�����kBl�~w��C]�����-?�|�eLZ8���z:�T�FϨPoM
2��l�Gx�ڎoZ�/��e�D>:p[�(1��7�����oUvm-�0�/צʸ"ª`���W1�]��f��:���C[�)0튪�y!��6���.D 0�*[o|�:x�]/"���8�O�t�'ʊZ�z�j���{p
�7mJ�\A��4&�#��Gg�����b�����$qPio[���2����F�fM�@�3Hl�:?��ۺ�@G��������T=��Xj�X M�:^Ir|]�*v�~t%��8��OAt���\�W�z!�R�}����	9#?��q�.� ���LWv���Y�Pʲ���f˫	��Z���o��xk(������)�����2�Ԅ�!EDX;_� 9m"՚���0%��L���ߏ��@���e���?��׽��Tu���^M-�ϧd�8}rZ;k�ڬ�v��s�K�U�
Ȁ�5�32�\��Uʍ�
N��Օ͚䃻Y���>��"��3�*�O# �I�,=����\>�?(b6w��s��#V
�A7|ǟ.�j�:]�ӕ������0Q�����/^m�,�{� ͖�'��Mc��j���xu�`�Kp���d��@R^ E!m+\��fQv�9�[�e���ٿ^d�	*<�=��r�F[�9(�;.�/�7A���۾�2*�}(��!ج��7�O�n��-h�#$ԅ�c?�~�V�]����gm�k8!Y]�ټ���#������.&�o(H�Ӛ�ӧ�w��K0�Y�>��!n�f�.�p��)�tLyO�_-���ޢŁ���_z%��0�|ͻf�F[D���veh �F�jA��VE"S�� � �f�����u���H.��i&����d�i�o��^�%����h�H����}��~�G!��ԕ�!jC"�aG������Z�)`��E�����r��p�aM%�߂�P�w��=|��@�6zN���x�P��rP�'px���x��~#1�HM�5`e�7?_KR��O��� ��S-�P�qj{�z�\,�3{�ɹ�nꅞ�ɚ�@0��Cf*=�)o��H�B�����e�6l�~J�_������?C��L��R��(oN���h����W�����]��]���Y(ѹ�mO%����?ώ8LbU�����K�k퀵����!F���&���~R��za=ǰ`cO�1^�^����	Z����C#X�`�g���"y��v�'�az��Ⱚ�w���KlhW�Y��V}nb���TGodT��uꆱ�8s�d����aPB%����X�YI�
3�����ةwD'G�ս�`�nV'��&2�[|�q��0
n
b$���R��vn�o�{��H�xe�'>�M��74o"���'�3}%�j���h�f@��`�|��6[����<�� J�t[�ׇ]h�������Q�ވzF�	^#���B/��s30(�⼢J½�:g�3� ���7^k��m����d�׶�ce	����DmQ�lL���.D�z�?>�K� ˗���@a�X�m*��i7x˖x�>���#b�o��`�ƀe(��2>��I`��R�BeBtqm��7�.=K��,Kesh�	уj�4?E}j��W�U���<�уIt5���j�A��y:8�ڹ�_bU�Ks�8�E&ŭ��}���z#GJ����yk�����.��|�^P�]SN�;��"O� �7e7��56�F\�y`�W��%�_e��&ǻ�C~��I]̓�F����X^��	ssΚ4�D�ޑ�K9��T/�ᄃ�T�}l�N.�L����1*/;�!���G:��s�(�	V��\�J��ԫ��Z8���W8G`Q���A�M\�yq5{-VM�Owɛ��{C�P(9����f�P�TAj�����7�2��EU �5�Y*�YFqx2�3�_H(0z^��-�3K��]��6 �k+�@�!н�#Ҷ]Ϙ j��f�z���Ͻei��87��yb��%d���w`Ps��V�S0�^��}�Ҙ�Eg7[oſ¤��i��
rX9���"d�e��A��4�J��6� F7n~��	�a���_n�qZ�~��ӂ3�,|!��H�|�tY6P�:K���<��1�O�f.NP�NU��A~��\���G��h��ݤ5�,�:e����h�PACQL�1�����={y��$�,�Q���M�5�
"�({��"���.EQ*�+ �`b,���<�#V�n s�@kmX �d�<�҅� X�I����1f����6�xx{��,]�k���싼G�$�P��:�Ok�F9�<��q80���410��e�+Zx�+�2�)��u��㴉(�sO�*�Un��O�Y
�D��q��xG�r
EU�,z��<_ۃI"��&(�x���T��V�C`��h�Ў�����oKi����pƣ�F>:���[�ZԿ[Ϫ���Q�0Q�\-0��v$��ޛ�#���(���h�95��_ޮe��׎M*�ؖ����,���TT�ٖQba������*NF0��#HŰ岎�L1G�8PA�<�Em�W�X��7d�V�1�Ճ�â�U����x�z�
�#��<a����1
��(G
�K�{�GB{����K��[�lʚ�J"���QƂ:b����B�j##T�l����q>�LiuIB1]��$|��(i9b��s+#h4G�Zz���)�>ܰY�UU
=��u��ኹ��)���[�P�.Qd�����VY�׬���������S$�� ��3��ϖ���(�w�IMކ��r���F�Yz[x����Y,������H�߲�3غ(Τ6�9Prv
{����%���B������LB���$����P�n[�j
b7x<u�{Y�S��]#���::��"����#2`�@��د�m�8����[����&�N�I�T�S�� ��B�aIg1 �S�ІVqT�*�� X3�Z���蘓j�ձY�Qp��瓕�hQ��-�-��z�yn��Di"}0��o�&�+��2��y���G���j�'�j����쓫���%���P�Nj-�c�jC��p!#��g^ĭi���fB|�j��E�u&�z$D�^��ʟ��7]���D<Qǩ�2�Y�m�+q�n4=M����I"�[�~�x8��7)�'Ռh�h��L��)<u�w��ܹ�4m �F�"��J�L+,,n*�Z�>juL��"3u�'�~�.��ǆ�����5�~I�-W땲ՙ{�;׏Kޚ����t/�R���]�������Ǹ��
���'4��6�t/Tȷh&�����i"jg�	�t�3t�3WQ��	�;���fbP��ט7$jmd�5��&�nk?������0���n��?��a;l�tp��m¨ڎ�͜����,sUJl�ÞγLU��:-����?_7b!���%�������]�����/��R�%�ͩ��&#s� g����|qv�#���RU�>>[�ڠ=�+b��2�����o���!T�b�*�О�ۧ\d�[uQ���P� ��e�dfe!������p�f
N��(΢=�Q��Ch��SP2�&Q��
ե�-��O��Y����Ê�GP�Z�{G�`2�����b^X�q1�E�@n
�5��8�H����$y�Z�0XZ��v�[�eO\U�@W�"/�$%��6�~ D<��U�Lǡ���䮌9������%i�Y�^-����b0�H���h��^B*=�,F]9z�n������Oq���p�m��/�#n>���������B��n$�v�+��T,�^�|��{����3�*��$r�fs��f'��L�"��D��%j0����{��=V��2Gq��7W�F�ᗿ�b[�jc+�̐j~�F��_.?0�*��[��UK_�?`Wr:�v�`i��q^�Ar�Ȑ��Sݵ&�6U��M`!��ӣ��ԚN�p�ʳ��J�
��=$<��[�4y��䒰菃�f���yڵ�1Z���#S�"��xqaV��OC�ઍ�ļA$EZ��b(0��z�O� 𠯂�ZɆ��G$�E�ק�;���3�y�aϘ�k� �L��U��ϒH��]i|�n�b�<cO���BS�_Gm���W*�.}Ox����V�Ħ��b�Q;zؔ��82&'2���7��}xom���f����i4cs\��ڴ��˦���d�몷j�JοI=k���ĐZhGߨU����N�@���u�E͖t�ą�W>�u�q}	Y�����v���0P�;]�`�ˮ1I��n�h���8��f]u�]�\`��M<��I!-�����V�I�ړ脃��4l��m�n�٠�
+�k#֚u���}4�rw�"l�ȅ;F��(j�Z�C �hыG-*m�NqǮۀ�e:�mS(�.�S��*��I�T�O}�$c-��P��>���R��O&��ڒ��>�o�g�����A�ԓˍ/��A`��Ļk�X���68��l�z�3�9P6��Oذ�U�=&��葰ْ9�~n1�~	���,�6��U��]x�;s�]������~)f:RN�N>)r���,�Է�F��{	�7
ld.j�GrP��Y��nܣ��-OJ�?�@[P�#�m��֞��2=��|a���̮^U���)���AQUˣ���l���2#�eY���6��/|�t���� d��{S�}��K�e?��^K�0,�Bq�3���3��q��vEϾ�ʹe���ƾ�8lޗ��n����m�����m"�b� -��]�h�f,�$)o��o�O��ґ��d�����,0�y�D�BU�A�����r�,g��*b�D������K���6�SL���\R�|���e����������JP�$1��@nB�ٛz��?wSM��K�\�1Cc񏑦���g���=]Jz�U�U�xO��v$���K�1U;�ۓ2IЯ"839��>xk��1�b�Kq���u<�pH�C'_����$~h��O�[��	������Yc��
?y��GnpOyw���Lو,b���y��t6j�-!�|ٻe_?��k ��,t�ȨZ;��N�.�W)�o�U�+�<>i�����7�]��x'o�7}���*��k-���MO!����:���Y[G��.�6tQM��%Ý4.O@7�����
���Wڼ�\��݅h� ƚ�Ii�q ���l��5�{zk��,�k_ў�u�S.�@�1�F@[}FԧT�F�������C�(3>CM��������Hb.�ww[
_ԔC|(] m�k���_@��=��+��h�y}0��C���D`,������ ����DY=�UC��SM�%��%f�Hm��Ҁ[�&��c�f��}�pͣj��~:a�25�J�du�nu��� �iD�*Y�����n]wd�g�Q�cJa��^V:��
�/�+w��T+�]"f�o��ݶ͋E��UuLd����$z+xy��c�%:���+y�SUߞ*o�<za���aa���aЙ��Ei����;��'.T�B]m�ꥁ��K�¤FP�/���&h9�qK�����S�5"��RG��엙֛��H�+pX����$]�֠nGB���H��rf3 3-� ��a�UpZY����.��$������aʦ�U-��F���$�;�Op�̵���PQ�F���N�a���E">��'� �?:ۂ��[m����������)
)�wi_^�*���Y�@���I
9���=o�2��5�����[�a)���=AO[�/ir���]!9����!�L��6f��݂���~N�@���$+�g澙nc'3N��K�& ��ȁ{�"�Z~�a��칿?ŌNz�G� 2HSP��Z��R·��eY$/:۸�;{%Z7̪`��e�): V3���N7�u�<rM.\�W�K ��1�!��=Az<��G��X�P*���s��Ty2bj�c4�G��g�@{�� �S���,{��k��������񾐕TȕY��J���z�ܻ��av	޺xiM���u�I�F(D�	���Am���ʵNك�r�X���Y'�yL�?)��v�/�!5����ޣ���e'HW2П�Z�6Z0,�Q�����Ֆ��/;�@�0�^_�x>���0O#��ˑ���s��8��.đ�'CX���A.�Ī~�A���!���=��ѳ��9�����q(�g^��q�b�ы�~�ޕ�\��m
��R�6E�'dd攙6M-Q��t�����I��xq��Kh%ˡ�LS*'&V�G���v��7�m�WS��!r���r�o�ǿ��k%�}�(pt���nQ猸�(�{҅`���3 R�7�$:��i�"EF��:�F��
I]���c6F�3�'����?�M��%�Hyr1{u�<�,8�b�҈��s�;�.�G@�m:�YE㄄�~����Z�05�7|��<3t&S�i%�@����z.s^ػ@蛫^�|��}?A4���c���G��_���!潻Q�͹����܃>0�Vwa���X�y7L�Fs��z�̳�%�8?�8ES�����)�s����k�K�Nx�3Ky���3��x�|{p�1
�!?1M�m�4�w�����/��?�� �8a�v�f@��N�����s��Ρp�E�%5�e^Qi ��o�JW���G9ٻB?Zy`�_�A	~_zlM�B�&h���g6�/�1���������FJ�J�ʍ�S��4��� ���aK����H \��b����T4����m	P����F�w��hH�å>Q��a�|�J~H.��zs� �k����n`���G����~�يg!/TzT���S*Q���	�ά�Ġ���R禇v&���p5�H^T�UN4�n*}��>����ʲ��r�V�����bom=
�F_;9ؽ��n���MuVEѰsށ��@�kI4�B���� �����͛x	j���14�݉b�sXw��ET������VI�UҒ�[��/�_�C�2Έ�b; 1�gA���|�r����x¯4��t� ��v1F.j�d%Ř��_!�FO�6_����w/!A����`�Oz����e�y����1�P� K��g��e噢}�Y���u�5�.{��Ⱎ�����o�t�sd��=���,�iHX�s�lPI��U��H�q��B�c���cC��05�nָV� #.�*�"Fe���96BrΝ5�NQP��"���3��(�	R�'蜎�O����b�FcZ����8�/
�M��&t��ʷ����Ϊ�Vq&�T���;z92_��0f��x�� 3{|�ġ�J��ƓD�Ah����B�}�m"E�2k���!ѿ��#Z��`F}؄�3YBn�1�>&�*��K	��t~����r��Τ�S�X�N�;h=��0��{кf1n&��.���⤪$#��?�5��3r�xv���Z�׶���6�������S�� ��e����]�t��Y�Py�(��4����ᩃ��t����=Z�h�R�����up�o�V��l�}_䕦w�N�`��s!���v�`eE�"�E�y)����.�~М1A��	�K�K�ӏ�ԣt����0�20��I����@ssړ�D����w���k_��͟�2�B�O�[��ੁ��޸Iz�w�\������������`Ե����O��T�5*ʠ����+�)5 �炔��4|a~��p�!^P��~��Z;ఝ�g���"v}��,���L���uz3f���6�6�2w� �������V��|S��'�u^֭O��� 3��G�p�r�b�^�R�Ip�(��|�|߾j�F�<��'��Zw��Q��m�&�oŦY#��;�� �V��2u��W���hLMb*�(.���HF��O:�$8���T�\�:�3��-����G�� 5!��{,��]�Z��Dad ����ͯ��P�h��gC�\4�o��f�z�EX�$��D �"����^�b|�W�tpX��$^J�M�������<��lG�CC�W�H�W�e�0�Yخ=�C/����ОO��w���U�&"/B��74�q�\�Hu�̘0��rV
�6��m�5�c"j��DIcY�i? ~��i��+����-���<d6���
����{s��cȮm��ag�����8�K'wĳ|Ȧ��M��lR<p�qY������"} ��Evq�9ۚaP|�?)�
�!�N3%�4�D�z��F,�������Ph�thJr�.��;�.�O�����0�yO$=!�
�{q�?��	�M�1y\H;��*e�/m�g�KH<���4�{�Ʀ�9֥^�Vf�{e�FsP��*�g�
 �}!�Q��ʭ/�֨��F�G.6���B��(���U��fo9O�$S�y@�_�@�L�`X�#�-f�8�|�k�9E�C���m)3�_E��5�ÓZ��ưv��0�*���*����q�G�ʹge\Y����>+�,c.k��5���p�ұn3��o+ӈK�)6�U샀���
W��_�ר˷l2��!��o��Z�ԇA�?mZe[��s�&�p�V*\C����[�	 �l�¼��-'�>������Vz걗�� s�4\����#Ot�5�=,���:%"bI���U'δ�\����*��U��E�G�hHG�u�i��[i������.����L�z	Iԫ�nK��۱,��P���f�BC
9��KM���)U�4l̝/���B^]��w8�F���4}�V�����ί�f�zϴ?"-5�r�h����A��,�+b�H%䨞�#����~"��2����l���3J(���(˸\p����Z�Dv�h���p���B|C:,��{BڷV佧�o�}mlbZbi�p&�9IFtr,�+���ˣ����9�Ky���@��4�I��V�"�vs�1Fl&P��o1+�ŕ����W�R/�3&��U��z�U(������u����\B�ĳL��R=!-��:��q3���t��Jlb?��^�N�,��.P/>���щQ#>c�D��=�帣��Г�#�gm:H�j��ӳ�Qwsfpa����J�Iq�/$��r:����e��E�dM�o����YC$��-N{d�m���P�\�����{��5C��~�w)(��)z��q'L�h�Z�z&�\RY�HA��������Z��j@8���������:���F�b�? �Im��2n�D1#���ߨ��K6������@U�����eJr�2�ƃ^�^��08�5<yǡ���|3��ado`c}�lIƳ�CEw�M izX�A5bs0h#A�E˖�5;w�%��m>�	��FF�P�D�%��A���}b�/b��δ�̇��5P5F��g�ׯ�X�տ)�'��������K������ݪ�N��ZM���H�aX�τ�r�exv��#��-Z��\dy��/6sN_0a��i#�����DM���m���0(O�ȡ�Xf�U]!��Fݤ2�.���G��#W�|=h�	WN�ү�J��}�V7��@�7�� �����9(�l�V,������ ��}��f9f�J�<�\��+5��HU�:I1�S�K.b_\b,�^�|���4��`�Eo}��y�c�* ꆖ��z�㹆�͸�z��@�����?h�Юg,"��D��܎�C�m��g"�����՘R�L�H�?;�Ɛ����j)W��r��!���Z�?�5Ƒ�Z`,�s�>X;�m��4� Wf�b+#���meF��r ��d
=�CZ���h�(�L)�8B�-a@}�~����Cr����u��E�2EE���b �*3�c��9ۍ��m��)�3p�ycx�9��k�z�ܰF��|�aE1 ���Ǫ@ �Qi2K4�`@D����
w��$�jQx;�~��Hb�z�A�I�P����! {l���S�4 ��kL$�G�LĔ�Z�>Y>�ې�g�ۂh2�X�Ww��ȥ�آr�~M�փ3�Hq�e0@`�:J{��ѹ�Z��c���Ke4��(+����+p��A���g3Q�5�>�G���t"���,�$��V��Ұ*��(Vn��]f����`�!0r��yqͅ�D�9��.:�R?a	��m� �����,�_�9o�|�{g/�J,O���chm���S�x9���vu����iǔ5f8�Za��*D}�X���G3qq7ä8�����I��bO�:��X�$t% Ŏ�[�"N��}L~*Jσ�T˅�����P�B��0*-��P�|�IL�B篟7�-~�ܜ��Į���\�XȚ#Ueئz��pd��Ʈ�����?�	���H£ԝb����\G�bM��&�յ�QZSg$JW���7��/E���	�����n���;#�;ѳ�qa%�a>��ݚ�<�MRr�����ZY�X���'Mh� ����0a�ucH�Bd�/�P��z�L���U:�}��d����(�{8�Iw�^�t���X����z$�W1����j��k����*=�q�R��K�à��w����ze/�(�P��&�����K�E1g����բ�)=^ܙ�

D(�2�~��f�!�k�=��G2y�r+���֗^}警+"@R��@v��[��{� �3���낂�Hw�3��?���`]ƚ�ꃃ4�Ҿ�-|j�s��Fic�����.�� ��)�O\��2���c���=9 �߾7�'��_�,���
x���]摿m�3\:�Z\<�B�=OX[�HM�h�5�uW�f��v�^�&���d +���'w�(�ԽP@�f���ɪS�Ed(��X�J�@�=��E9���PV���>Ll�Ks��D|��2T�0t�*����5;�Q�=���F�1J��#;�"��P��Be��j����^5��[�@ą�j���X�j|�V��Q�BH�]ٻ����%r6�q�h|���4p_c=ڟS+V�Ͷ�l�Ď�
U�P�z	g=�w%�u�p�.�`�@��0 �uj�f��d��M���i���B2���9x�/�ř �L�JG&�� w��������Kͽ���w]�'0�S{�!�5d^�X���wJ6\}n�M�H��Ûy�~�D�u��-�c�/U�&��N�gU
��Q�b󀊾��*I!�Z����"4�T%�#��2s7d��Ep����# 	:�n�	.�e� �)�EQ��ț�+fs�k

x�Is�����Tf�?aId$'�eaLj<\K���F��|���:���8�?E�k�	�|�쐮���,�ר֐�跐x�p\c\c<,jY���=ô�� ڍ!$16����0��w��l��A*�_�-�
톿��
����sd�6M�Pq!�r�Cίɹ���D��8��yʀ��]�&cE��`�
i���8��L���~�/A�%0m���T�G��p��CGޮͼt��qY5<6�+e%�a!���:�_��Y7PКB��p�Z�3�꡿m	�I�;gM�gI���d 6鱲q�D�Z�i4 ���HV��v�o�oaGdg�+��F:�GCڽ!(��ҒG
��1���D ���:�Ǻ��x���}XHp�����I�2#�����;���.���7�>���Q8�~`O<pm$Bt~ҹ�@(�U�����NӘA�&篏ʏ�f��g�ض�Ql��1��/�]W�{X��K�����M1�T���Ёyb�^S�JAC�}�r���0��/wk�&��˿~iK�@�X�K$U�w�`m2)F��/�g\���ԙ�JY$N����������; uǾ	��v$_����9��(��� �Z09�/{=�l�q���ty�Dr���Do�ET�p
[��P�uS�X2�2^��4���V��9}J��㺲ۛm��pjh��C�v�ů��^I4Y��LA�,ո�[n���Y_@;�Z����h����&��䧇<����=Ҷ����������p-��b�zP:����̶p^=8f��ZkUTc��B�M\޵����;:8���J��r����I��ki�G���Iά�ߜ�����I&��i�B�viI|or$�Y�����B+z�kH\s7��7-��$F�J����M�ܠ�yD,�6�":�C���J�K�\���UO Q�̗Ӱ �gH٠v�\C\'q��e<>QD��Ǉ�6E�E8*�x���1�+u}O1�m��t������|����G�V�zp|�4Ǳ�ϑ���v_5el8��~��K 5˹�P+�恕bMd���uE�����+P9L�Ja�JG.ԃ@�5����ӳZ.N�5�p���0��9_��`h��98H�SJ a����Bq�"|j�m"q�V���j�\�:P������L7|���%)�h�
��zu�­��"s1xA)�)���<�`���r{\T�:�o>�F���+�8�QWLB~\���&�fϕJ6����#�F9�	�Z��7�
y��Pf�ޠ�!�!��|��CE��9�P�V�G��n�&�Js��4�@�ö�>"�l����K�ז	8�&X�,����:���{k� �:�2�w
al({��6%Q���\���Oϒ�2����������R�f��'m���&�G#�n��(C�Y�fJ7&�a�`�#�gzСc�D����zŔ�77~�b�QEu�
���?�qΙ!u	��s��16�}������gѵ�J6k�i=Ғ���t�+�L��!-q�ZZ����G�/2@*	>6�_��N���J2���H�a�6�jV��a�p�4�[�Q�.�r:�qЊT�;�'��{�&"�������zЉ�jM�"�}�<�oH���qv�:@ɍ\h����H�u!5�#��oBaᐾ�W��&Ro���E|����/�h�E�֡��
7��TQt,c�� 0�&�Jz�A��kE&�[�w�.m�=/]&�5�=���HR�n�Vp��Mt��i<�8�����Ǯ|󐌕��r�\!�f-��(����?)��l?���ޕK�Q���!�<��P����0Y�?�a8e
J�5X��kgu�ܴ�D��ć�yh�r._
$��)a�<�����p>��jm�W��raޙ��uV�%-[�L�0=
[\�����܊��9W�y4A.2|��l�m��d��3y��/�0��1����;%5�7���ZzX�Q��;��"zV(���ȷ&vT�j��x�c�>�nRF���%]y�����\�S�*�ܕ �%d�N���J�1��%5���@��]X�͞�p��!���UEFC(m�!��士�ԣYQ䣚�����;�"���ٍ����K��
����{~^�XN�����!���}|�e.�]Z������P��(i��8=�����q�V{�%�ᯧ:J[�7֜&lR=��ѻd���o�uCvዄ�,�9|noL�%_nП�]8
�P�v :�\ǣx�ݬ.�D�t&����4�	�Z#��Fmm�d��D�>� ]�rr$"3�	��9>H3#���v�A�<�I��)��7�����R�.��i��0x+�/C��\��}��#NR���:mR�~��n�aB��ST뀗5am�R�ܯ�+���o����}�	d�~`�R��`f��u�'_U��f�0�U��[��O��߿|	e0bG=�)��˧i����/v���P5g�v>3��7��V�-vI���8����5�A�"���"Cw��h��Љqp*|j����B�.���Ox�� p����U	.iY��v̞9�PlzC�m�;�{�f��j2��G���*���%���6/Qn#P��/��Y����.=߬����0���lo	/�*#$�����>!]��@4s��"���H�1C7B!Vt�6u"Hpz>����7�vD��AB�>Ԫ`<�]�\z~�F�����p�Y�A�UD,������j�xP���ݍ��G��d:�`?d� Ե�I��ُ�����_J?���.z:�.F�^8I�E
 �X����"�1�tˋ��a&���%����9v($���wu�ɢ%��b��"��AU�C��U���v��à�s���]��q�hw�&�d���DFD2W�2U��8�H���l)�E�Iy������P7�Dݪ*�=؆d�Np������P����B�R��8�]�#����1�  �Qf��5�%�&�KC<kԗ;�Ğ��֒��i.�R�/l<{,��2�R�@���C+2�n@�{j#�v�A+N"�R���o~ձ������p���ֽ��J�e�/�.v�H�#)n��Y��O|�`�4&�@a�:��[!�Y�,��p����
�~B���߫��ђ��?��?��v#��:����˥����Uݥ�$�a�|���S/h�kQ
��}�K*��ZWt�3�-�p�v4����q�V�J�ɴ�I��xm�"�����LI��5�H�	n�[�+�P ���]�<�W��9�kI�6���V�H�ƊyE�W@�~[#�)�$h�c�'���a���2n;o8Sz��U��@g�KiT�.s�}S���3�[�%I�x�B��ݐ�����;غ�.��xkh�Ql l�$�8~ww�S� I.�c�Kq	�۴3׫�J�E�-jnԆͩ`�Oy4���\��9��<�9�D;Da;�9���mJ�n5��gª!k64�IEA�D���k�\x�VK�ߡXP��� �P��)aٽv��5�>r��_ܾG� dy�L¢Ѐ4n�� q%s�K,�?f4R*�AΊ>>�h�$���ʜ����$���"~n�	�~� ��M��p-m+c��~����D�z5 lI��;�x��&���s����bK�o��=I�0֬��Ҟ�ʁ֪�m���	�	�b�.]^
�	x��aڋ5�N�xͻ*��ͦ�[�yێd|\�4%�꼼��w�#��%�����L�Y$�8�aD���h��8��������������zA��έFb�긟���4�
�ˏe�7	G �}��n����j��\�ˏ�H��SǙ�YY�A��Q�
8KYz�7(�n���=�j���L��.l�ݨ.N�����*P�E�Yx�z��7��+x+r���7���@4g�jtP<?�?PT8��P�@��G����Q��7M؏zl�M)�v�������;06B�nT|C�G`#�-��6�o�f�H9�מÏ����n&���9r��^_�)';������3�u��SgർR�6�/IR������	:%�����=���̌ ������H�z����N�S��26r.���]�U"�S�v^��R��W5�q0y#3�0��К�p�.��b�:��te�7�K���^f�=�L}Qti`T87��0��	'
L74�WI 8<��A�?���\&������O��*�*;X��2��V�>C��gl�2��k>���o�+�z�U�9u��>��p���x���jnZ��*���R.;�X*#���!��C^YC��w�Ml��Q@��9�_'	��cl��{��=���*�÷ Ɲdĸ�3=�;%���8a	��p��i�#�\�i?�4�so��_��R��|����[�q��x�o���_4$��Y.|>�t�X=��j���������/DEF���E�y�7ֆۢl
`^��B�׌�a�sUO ���..hQt̉9�OY���y�����{G�GYCgL�{L	���8�-A"��<(͚�(�%��S�.�Œ!�A��$��`:f`4_ ��"�=��>�9�#0&�ߩq�?����|�JeP�}�C�m5e.��fIV�Q�%kRo��6�q_�,5}�#�Jp�nn��q~�w%_�tUwx
K�n��v4C#���W��H�>&�(�<�Υ'T�o�i����6�qV'<o����ta�ҐfBu�*���./�5��=�������@�DE΢3�Ǉ��nui��a�$C�-�K󡿷���uc?�X܄	 �ן�+3����L��{W_�Y���e�Y�Ͽ�m�����	���G�b�UXر�]Ao(����Yր ����E���n=�H/²	��\@X��͌�a]�a���<�$�Y�@@w�2xxC�E����G���\��C�m�jP��#��H��o�Md��"�-�5���ؙ� Z:B�p�U�Ѕ�~j�u��P���;a{�^7��g��4葽5�]��1���ԕ �ؠ1�]�T�#�)��I!IF��d��"Փ� w;�gV��?���ĳ�v�P��8M�tR�;��p���>' ����v��R�1ԂB��d(q�b�#|N6�8�M~���^����#!O�TD�p ~�;�\4��������w�:��N*��3~�,C��i��(xkw�����]�K�H�ԁ���Y��}�Xd�ʥ~�&����f���Ϩ��@��.�szsYJ���$�N��-VW�Kf��H�
j�_4L��M����K�{�S@��FL4L>�Gɮ����_�Jg�mY!�d�k���V��<���"�=ow� �-��`�nd���%�?t��; ��܇� >@��}��s�Xt���x�#q��i�8񓡭=ą�D?�Y���h��@=J(A�s3�ԩb��N6��4���i~x��*�;���߮�_a��<C�;��u�SU�C�5�z��9�u��`�!K����0�bOq�o�eK���mX��b�W�X �F�`�g'ނV�-��E�Um�R"]UW��|z`NK��SE��w:�+�x8��ҵ�j:��w͞juB��c8�,%>�F����"[�ҏ)���p�͵E'	�Zw3 �Z!�����"�՝��$�f�M{C@���>��XJc�A�ک�⎑g���x�0�x�Ց���Q���{3�?��V�n�9tY�q«2'�޾�������Б�?��D0-!L� o��II�U�O�a^3p�����9���෾��.Da�z��:����B�� m�)�BY5��rbq�a���`��5�b&2Y�6�Rw�4R>�8[/�Ms,J5鹐�����`e몧f����Z��mq������u%��[�p�u)-*�m֒�S�[>�)���{R���lE��oZ�T��WX��/���,3<@� Ja%%ax,���:*H���R���i�$���^7���y�s��S���l�%hY;�������/�vn�#. �I�4�y�pWե�f�1�g���G�Y{YQƸ�.n�R�Z.�t�~���nci�$��f
w���V���>�J����F%Q +���O$"��U��2�~�vm�|E�H
S��	X���%[hjm�2/c�1*��[ͅHl4��gZ��7��@b!|.�n"u�I�cH7�$�m/��r,?�G�Y-w�%mb\*�S�� t���`y�ځ�W��nl��F��l��X���)�Y��:`��`XL��t8M�dQ���ֻ%6��:�'q'�΅X�[�@R��h64#���((���1[þY���?�e}�3�|?V����;�.y2�9j4r�E�����C� �d#�W��)}��RJ�?J�6���"��w�{#�W-��� {-4�I���e�[��$�P.S	Xe�;���;�TU+����(QT#Le�Rz�<�7��*Q��n;��o��y�U�x�켝g��-<��hv�g�� ��=�i�������x�*T��nN(��V��tM��ޥj�{�&߅�nB[�W���	��ì����a�����!�G��IA�;�sL��6˲JC�G��������m�s�Z��w�$�nYv��d0^T�(
��|�.�k)|婅�Х���{�6�//�ec&Ќ����%9eab��s^�GI}"�*��Bl�9_����H횙��o����#6�*���	���������H�Q�&��1�)?��8:�t��(�շ��&W�
�@(�|��qt	�+=����=[�lL�!�ߨ��+��9������ gӪ0�dR9mWi��Y�#��Ef�c�zÿ`�Rr!ިs��R�F���ƫ ���P���!9م�=e$��5�ZYv>��6��M�����pЗD�#)���v�q+˿P��E����ɇ�����Vt�Qru,ު�Z�&L�J����9�j����{�e��o6��Q�p-	y�Υ�ަ]B���TH��������zg�~���{���k�vBA�e)A��'_�8��פY`��+�����8	zG��lt05sn�,9:������'G�t�*�9h�}���|�
Ǡ�KҊ�)u{�oˉ��
��66U<_���HH��!�>�5���i��/� <����S~�L݅)��4m����'Q��A��K!�@މn�H���sD�����N|`�F�O�2���Ĵ�V�"�5� \l,M�W���i9����W2&/D��_( ��CD;�I,RJ'm���s����N,�МYM��l�i񅷒+����-cX�� rf�0�r��%N��F�����:)��y��0o*i���~~
�/ ��wCRJ_�-̔��2W��:YyM��=:����y�����}a�}�� �N?H�Γ:���f�!�Z!o���'D�^����Y~-���"�B�\�������H��7~;�+z{��=J��H�%X2���0w	�9�ٲ���P���.��HCĶ�$mm���oR�7S��/�i|��5#��yB����5N9�&Q�r-��n��wIu��rb��s*�3���(�����ks\�!Pnh� �\�4��+��-�):��MM⓽�����m��h��]�S2F��{���R)�r̡�c�1�i� �Ie)����N3�	�����ۖ����A����on.C��NF��ݴݬ����wF��w���o�]bB_�ѯ+@���T�,n��)%�[��P_���L�'�ա�_O87R+m�}h`%�!���%"�J]��ko<�R�k��7 NƒW��t$<gqnQeG�4*��K{1ǄD˄�$iT�{l�eiz�Og�̱S�D��ʲ���M)&*B@)��[��CTr��U��=�e��	��G%!�i�>���,<v�;%�[Қo�),LP�����ݒ�S����AwtYڐ��C�t67�Y��3Y�ą�c'�w�ɛ����߭��G>��I��`0�l�-�ף��H?�^Q��@Y��*��Z��iWhl�z%߄k��@��	a@�mO��E�2ik��՟�WL���I1 ��g��B����{�\�(�0*��嘴S�4 e9׫�� S�˥�i�a���?"̱�!��S���0��Fn�?����-liK,(api=�U��R�ڦ��H�7��a�ֳ~W��wL3ݑ��t��y��E`�5ط���|r>�r�7z�|Kk.�vF�7�y��t�5�������j��ݛ��HO[�x� �蔈x�,l"�n���H ���Dt��NmX̒lw��qw�G��~s�$)���e�&s�D͸�ilJL<�R:ǯ1� ���h�qq�U��u	)��6!f�Chʃc��ȯ���H�c����1�^̖>��?�G�#=�B,`o���4j ~J��L��1)q>%��4ٿ��	��oW2���"�$Ú�-���Ҁ ��9	�T���6.<һ�,�n�_��>]�ڂ%W�D�-$���$d��BS�Xө~S6��tCE�.�Ba ���A˄�1����"�0)R"��20 _t��;�4���(��K�`��������4����[>��6�(޷���T����C���N+��?m���|b4<�Rum�����L�\K*P!|�N���21����S�k���OI���Hj+ALt[D;i��M���LH��/�l�˙�j��{�)�ù����ڌ$c��R�/��}C�Ý��u��h�^��I[����C\�}��Il�`؈���W��/%M��X�����&l1hjzT-,<���I���3�x���qm��A|���1�q��/���őQ-l�eC���1]�)^g���𞭌��>͍��� +A������Pa�]8Gq�m*;��3
d�ޠ������d��`:���3x=ʹg���al�{pDqH�S�:5*��>�x��6���V:������N3M
o/�#�)�vg�7D�����mq��^	T-ډ3�Q�׮ᓃ�Z�t'O'I5���w�+w�c�Z٪R�HL�ɚt�O�h�GhX��="�G3���T��\n��
3�x
F�w߼�h���0+��fji�&=�.p݊�gZ�W*��{B��Z9<�(�����R�>,�D@�G0�����I�$�N�U*��nm�`��9>���{N�[m:@e���|�t�®�nG"̌g����(Y�oB��1�1]���߁e�6��!���m���]^i-@�;�}rqK��":(�c��x%�z�|��t�p{'0���m��7��$B�t�L��mT�/�S�ׁ.���l�U<�5��
�dK��캴#0�t
..��/d���'�
�'c��1l6��.z��ď�e��%X���\1���̀پ��mvѴ�����{̪���`;�)�$щ����唱�x�b��L��f;�� zc~h�C��H�77ׯg~q��2�{`B�#$a6�����<m��Je~�����:Kz����a�ǘ�f����$�(" F/����S�%�B����sU��S��v%�8R�������M���(�=ZŃ�@��A��2�?U���H+�m#�>p�"����Z��Q@�-�PN��s��x�f we �t8�F_�v*��&���d��P��Ư~w��O��,�`�J�x,��:��V�KmZ:br�}����Z�Umh3-�� j�P�yi��V��Ղ]��9����KY��PƖ�Q�Ї��}�(��_��'���o7���C(���y}�����g���ZQx�F���v퐶�1��h|���错�L���#����&�D
�G�[]u�m�-�p0����]�1��*
/�Q��g�`^z?�|J4����K�5�]|xQ�[����H!7Л��^�6�l��-I/s��̭�{n'ӿ�֧b�%7���%p%�>�=R<'i)��.�,��)�H �C��rnX́�_�KZ��7\$S�p��R�<�K�<&���h���d�ɛ�u����j���z��Qb;~5���,í1��p�u� 9���`#�I�ҙ��0���q���;�?er+�x�^@>Bb��#~D��'PV��3ē�h��EZ^f��"5n�(�<��om[���*�U5�N��?$��P���N��.b���������E7R�@	)��	���dw����˯�HXs5�O7 �->"3��|N
�s��ϖg��܏�Ѭ#	n��֎/��o���Of� Y9�����#�0��H�}�C�=�a�Şzio�^g�@�7�p[�"������JqG�;�^����������M:6����<-���ze�A)E�o%���yN�D��⌨�O�&P,K*ʘ��8k�����X�c�#݋̈y	�j1�^�����I���z���1�	���)=s�I#��}�N�O@����Iv��Y��?�NX�R��J���<6�� q�[{��Z����'?�f�1.c��(�}���Y�=S	��˷��PK���낪��:��4�"	Dv�}����\)H~Bb3k�Pn�jV OE���>������/����KVɂ�a4�jP����x��Iu3]5]�F��G)u�"2ӱg�<؃�yLg ����gx���{��[u���[R1�"�2,��O��s�rx����2`keD�`wb��0�;g�~>�P;�?����X1	�-[��7vNH�'�5���۵�0�_�qZ�H����^�x0�yֻ^^���vo��w�t�><����ўw�ny��t�ex��mxm�o~�N�MwkBx����5a�`n��	�첮�X�N�տ���C飢>��-S9
�e*��8������MW�;HL;Yw?�'3w�k��>BQ���&%� �
C�E WD�Uڡ�Ѿ�����R̳U~��I�+�%�/)�{�bD�p֏�E\��X5㜞r��������\=��ũ� �>�Y+�(d.�B��?η	0&�J�?��������,��PU���u�u7f�B�]������\����H�	�O`����	f6
��4����>��|_7Áx�6���/7���=�3�W1<��of��ɰx%�4ŅQ����k�.1Rל��t;�e�,g?, ����qz��Ԍ��͛})�네e��3�����#b�=�U�"���	�32��q�U�7�{�V�B>[�E�g�B�UK�<�4�¾��#z�ٽL�����mN� ��-C��36�>��MH���U���OIӵ�8�+�<�7�����3?@��/���Ȩׂ��t��7g*��;{5�
��q�j�زڌ�'Z/t��	�|�(��c�S��-��}��۩"t�b�'���%Uï�꿤mt{��]��N,�e��Ѩ~��w90rѢ���\g�'�3���b1]�j�����U�:��s����a>���O��]����o(�e�K�3_؃��