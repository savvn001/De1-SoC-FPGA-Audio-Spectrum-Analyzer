-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fRbn9CdYR9pRg7KguWm9F0o9Tgbr4iuR4528fy01eAa0B+Z3EqMuJiMseyQNZ+EnmlNqRYtScS3V
+YvjwfpZfhT0SlBRWs8rzh1o+8uEJOP12LkuaRzAG9PSGYbM6CQTaaV+Oe/DLQvThFltU181sJA7
UpVjiAz62UsVYcs+hhYw8bBUPXm3Y7PNASUnPaY2rf8NHtWaSV8AZjvE/I+BEnJ3Syw8oEkHSgbb
2UPfw5ripZKW19H/VCUWUEkboW6uNF4AalinjBqVn3MBucU3L4adaau5y/Io6EnMr39GD0+sRfZN
1yR4lAieLGdq2EoelxMK6J5ixW+M7g2NxnqVag==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
VYkiJiWr4nVgbXQJrPaRBPOJe5aYj2PDH2WQpe1lR+yXDi86vJP6j6tn0lYk2irs0xHLee3Fmva3
n0Buvy9YrQH3RPynb0gASKgPkfMbUDn6GTn0DzLt1Q5f55/jPLifFmoRJBOJzfoIqVKf23AwAcQ2
q0uwazJmLPyG711uqntXze2DKSgBVFCb+UbgoTym5L+5D8do4fn7W0rxXx4dBVHSRmuSqcAzqlLZ
iXQbbn4JTG4w50zsPp78eONQR7eSE7UsjVpfP4EYb224yNHghujZSEe0ljJ3hATInl6BRXdrS1Ko
0PuphAxMiA6WKF/gEBxS06OowoJaaGCadfV8/8TKvstNh3LNPCUNVW7DFHT6N26TYcrpzEomqzc9
LwTHfxoIVh61THF4JOAmFNzf1YdJoh1/lzKAELn3s/aqtk2XOYM9nB8KOh9XI4VZrtlFANjMPFWQ
KvSZsp49hoFcwuNBT3ZEnpb5gLjtc79eGi/IpU2aaDcP1JpTYTyUvGWuL9lsfGGVlOWWS+wHwguY
ctG42qAjKLQRI/ImVRyTmcQARaMdY8QzqYC4S/hAwHriTpDqJR2xko/ba9W9kwpNA3m/7+qIFtQi
wPKgkl9T6zkcYb+fNwM654Ru/wNBXuoLwrPIfFiHA2bKg9PAmp7BCHDnuSQTwHqExm2SVDa0RMcK
0V+d3tNfMmWNveynwpekvpJxv26yFR8PH1lJWfw3Vy+An19AEWwYu7wkZ9Q/OiKFU3EZ2FXIWeFw
gSLN8JnOk9x4l1+hN/zXDZRx7O65OYByD/dMqe0Esj+b1R2Ewh/NVkSoX6UCH6+7/FJFDrZMSkLd
hDl3Iiy2Oa8+RqxMawtoJuVgHEaDH8CXarr60G/yFTGDOqFzCQ4z/vkPTfdF7OILXRBsLL49262m
OOsX2ywviFRiLX8lloN2gB/KAo5oZLai4LgeCQTNQ23LbfQHmg06shmARBkqdw37QCA4fFTE4Vih
+i8igEeyQQka2nluh9E+aislltWD3wSTl3nOANcmu/z8lIzCp6SmhiJFzdAszH8glITWX7aU0Mth
zwLLSrXPcGeSkr0/kEPk+l70+Jbh+6EeLzlcphNz7stnA8ExWACosfxb44yq/geTCr+/ceWUD8rY
XkpV45gl8uqMsELPSZ84k8RlKpCuLFrWAi8HgmuLu5FbB/egeZWhyRXK2GTGYw3g2pGwugROeTR+
tn9GlarhTlWAchEKWP2XJfd9q+uGIBU3NIY+1Q/M+lTC4vj9gYVDxaBOOQbp+Q76tShHDsiQaSYX
TzZ1BbckrjmvFBYyfZNC1HKTmTz1o84uRtNWGJTng+Neig0E+9go+kjagbQ0G2s6qaKEmhk0KEzl
3+mQyqt6fBAJlWChijHHZHMiQGNQNa3S4KmOQYBy16hlyCTJekcgvHZbHa2TgUsMNPkLAhZUIwMP
fc+DRI6ghXfplU1ov7jVBxDtRJ3DOl32RkXfxRPCsm6T0ZiCRfCjez9Ns45ytqQHXRWbnhi7q3XP
+qER4toikSgVYZZaXI8TVVPQ1TLuKIbOaMhTyCQ04Xb5VrLu3YVbsWPlIaA00ipwaWJmGWkqFZGT
TagUeYoUonMkVTzVb+lWxCVombVjFSYemvKGXMihOtMz747si7pLzCT+0nxTpvFOq1nZnWPcM7T3
471twmjyjKQUBxcwaiLg9+D0X8V/PDH7fRZUmGLAZU7OlK2xtVdQfscE/0VMOcLcd5K9OWzmbvji
dVz0j9UI1gdIWb8TjZw+aY4HTKxAIMy+u5j8YI235Aruzh++WriI+0z6lkjp41rzuW8NEuz50D96
Rna+SnUrdh7YDErgKFPndstILWxO4KUJ09qEY+JwvFF5nnPT7t6twJapf9xosGTRR6ocOLuznniP
yMC3aXbcwWGYqCAu75P6unRKpJO4Hg0J1PL4nZEQznRawyXxdkagjx3RN3/SNsiZIxW6tqJ7n4w/
ZMMHePCIQk2Z7bim/eLL3jUVxG1kHy1U4bV0rlZghHNReEyoiaMrYGZWROBC7ZDlEuEsoOnHFJGK
tzvyunkQerjBvbHBT5ZHNGfVHGB1niI++7/ksOcxlBfX3B4dhpaaxB/C6mKLLRgCAkk4dvJgo8eU
Kj3B/+9KhsAvHqKyyyEU2k3kNDhgLpxv4WL2zu8W36RZK2x3+NkZhHF7JPg+rJJ/2+7zaufgszf6
5g3Iu6/t2ZpKIPzJbBSBFte3ID8BEsuSfqW2jhtD20qZOvs2KskXkkio83t9PxjyXSHORGq+ElsI
4rDRkgZa/wthF/wzlra9sJfx6LEps0f06XQQiLhcRJtXWWBJR27ZVfJCeKzpW7GN6OMaxmYJ7NwZ
TD3Cr133J+UZbsEGS4eweI8yBiAbD1WccAdeMHc8UHT0kjlr+C+i4xtd62fiF3o4X+1G+0mMlEzh
pIdwvybaIsrvQiE2/n08IgdmyG2rIeRuoo8tXMoHizNQeKCj+yzGs63rGXpEaP74o6QtLAMRleyc
4lnJE98JZPRkvzjX4eDe7X4txb5Kq/c2D6SM0F1UrpSwvKAt5htgRc8N47+UJmo9vh7vPnZtSnFX
yUO4B76O+TldghI4E4f6vCrAfMGuRwcJn/4aJWiIgSlw9EJCxUbq7LZwc9fK/qwpw6WRuD0plZWe
ntWX6uAQ/DBsgm4Hgbl2Bo+D/oHoTSZc7R6fXEYMJZl/3GotchfTwrpIkqBNEUh5XCx/wzY0H50j
VXyHLTBWH01Ne4mDgXncXiB5t6geDbtdNkaYuSf5lplSKSYVSnxQWrsZJlssnSAdWpljt2v7mu3b
5rof3TaWLIQn9d46fm2yA346ZURr3co8KdHxrxmCPRFgoabYZ44IQSRg/1gJDrT+SZQmb7ttjgM0
3dCjXaCh1xi/tfXOfD9Eo54Oi63sBsf0LnjDkNPupHfYWQcQhwMdaz+xll3rTvegQGXV3bMyV1v0
6xWSu9oJ+hiL+MzTX+k530m8tEhdiZekiIqVmu+CLhWj2wph1UW53h1wNWlaxcI7R3pHzSMwmLLD
s12bGR0IKGAC5DZg2hlBT9K6I9xDaX1NbHoPmd5Y3Jj6uJ9W2susdnUm9pscEPT96xoHWbkW+oSC
QLv8ua9KqcDu7TlnfaN4MDsdXC7KxBHn+F7urpVCpeJi+90/Y/RO/zsmhG5mg+Ms6ZmUx6lhv8dE
NePbra7690XHkBKY9JBjQ/mQGCXg32FnVxDgR6GiEI28BsQCK62J4mKguuUMkjWQs3dx7DqZ1it+
e/+BCzM54Y91osCDoKSMijzsbdTi6HZPaNbPvu1EfDYM9TwI1J4LArdtIGvLcm60Rmb8/bAbdC6f
ELdk0SWCQ+PR3JbJsU+ZCPaDEBWd5WzI3Ut3V1WUwjpFHpjlEC9H7V2dR0Nwf2q/sMR2XYIifLhw
BTpkrLabcgOeSk88KlSwybEgecZsZ4eEw5kOu6biffdTRzz8eoSXkRxEs67tWQjHHKUR6xRNd0vR
YlwP8M738BUgx+PF3NWJCJayaI53Z/CCeiPVf/hrNJPB0uLS/9Gl02av81mdjt/i2Xo9ag2xe0Iy
IfeaR86zzOZm1K9z5p6/4pjHCzyDgz1YOJvYjwSKsyZkIWoo3+MOWFCplo4zcRN59wCMVWRs/Xi7
mVYQijfXIuNUu5qiZU2LdU4C2Z9JcPICDuPNvOuM8TcYCZIWFdLYaXV88chPRWQhA8rLM1jYOAL6
Dgm4cF/ucfdbW4N/p6TDIr/aXfX5RdNfCtODgfThNO2bMiwWWTe8uWtGfIJ24xx2MKMO9jamR/y9
t+1ZldVsEz2eKeibEomE7Dc0QsEmUEYrpqPcfb6J/ixsXKjAv81yv/Bkzsr9un25MZrqpNjopCuY
JL4X3ADnaRsm+hEE5VsoKxp+j16p4P+/EmnYzkvRqIMXgAZmKWcRs/fPPvFMEVFA2F159qpp/fse
zFzq8VsKmZubw/rWvH3TbF1g5Y7Zu2DKG6JIsOvumVdm7457Dmljh8WixtEv98DKTWCTmYkN05SO
Ldk8G6mGAE8cbD3l21kFqczcr+LzoIzMkXxBL1/xH3QpaEBjL0GAoJ9k0kCRuehi9aKJflyeYZDb
4pFCmI2bzCAOYuDhbM252u/N2stofcVK9QEFh2dsk1CgL61Upyr2xAQLT3bB8WGrdbkpcOXKkvt0
vLjw7QHKpUtcYqISk5Rs859lRGWLowVCPb5r0IiTS77aFKXoLjSxgWWU8d2FAOXBLFncLIzMIa1V
8Pi+KCM7hvOf2+s/hc2oJmkYwsyFhZp3UwttS3vArBepHylCN3IYKGKd5zbm8nuyoYAYueQ79tQk
3cypZljOtiRR7nqXO9KStbKPDHFs6pwNVXuIbByAWDaUxV97WUIPqq2T6Ex/5Gaf/Yy9B4oUwNZ3
1st3Y4lEU2s9zAadcMjrkY/RFz9Pykd4h2pV8roeBEf1Lm0axq5akY03VaNbmNcfN1dO6/CuRHCH
cIa6ys6KoRaLTgyHe7xMGL4Zx2oednuQ34ESpjfHcIgt/pVBCRirKrLoO0vzhIqudgUyvp9p+9U+
/TOQ6lRlYBpHlQgY2hbrSxcq16Mj5gLWqp0FETHI71gcnjUvVC48m/aq9Xk5wE3zYpAuLJBK59w9
m0rYoB2Jl/67KG+6Crh0f/rOfNGh6l8CQmwZcb6xLdqg8fchvrnDWoFIqS7IsiHLtGX+6o3TNG50
fs4BZ9KjB3UxhRx7zTcQ2w7UJG9xAAzxg6H4iI6TxQ44b394Mul7XOcB4iqa0hQwdP9ucx5cuPqJ
BidTEbADNoYFBXCRRDQkCWzvfet62EgLtv69+YnWxoxT+h5HqrAyLa85/4FvNvU9YzTFs56r7grX
/0NtZX/oBeJXr70PJCDDj4jQa1WwH/gfH6fG4vIRuY9MuWTrvWyA1JygyMyFs/f6kAqgmeOcRiVj
xeK/Cx3qJ/Wk+siFqpWtv9VocYOmKnKF9ilZTpX8NmTpSO+WfjumizFrleDIq3t+eFYPv350Gx9K
w3O0HgMglxCMiaSZF5eDixaGYBNJUr/nbSoWn1ildTZZwlJ7855hGcTQNvblHiJZbgmuF5AR+3Qs
hFljDvl6ZlStmQ8iVGVqbusOFQVP5Pd7Qpife+iyuWsZWtcmyGsPlMB9rb+eF9OzaWljqDJAgppg
fsE1SvPfCowe4xYupeR30aH4HdYZloDPsFq/msWw0LxIPYLAZwlEV89TDXaRGneyk3we4cRYCvI+
6PbAZpW3zVV2FEZmIq2DxN+36ekejGNYKLRILJTRroXP/0tbkFlwCpCnOC6HJjIrKQS0eDFgJfNj
6IhDQ0x00zbCJvEYOZsPZF/9D42fgtXNdL4gZTfMTe44nYQYy+99r4iJIOGqhl49BpvlGTiLxZGi
MGdds7xFHs8Tf9v+8z+YBCabefJKJbYqHHsU2JGtIczjAz85pXqZtbABqgdUNq9LLkG5T1hiY1l4
DXRxjAz3t1IBR+e1ierVaeWT61Iv/433oGWpYl9r52Ul+YpDtOz2lDVnXRKwcGiQ1TygXtY/Tm1i
kNh5btAvl+htaPTGVChgl26A2vzoy9BQleVW77zCPDnljwR7+oCYedXc2nC2vU857yXjvqMRTGDe
kKPOGlyvdVLf1135aIjm2yy5m7HxoQbLl6Cbmqg26eV5bREj0K1PWiZqJ2EWRzLiQ0ezXkvWBR2L
ZXf2ifThuyIpPse0pP32MDCyiwvXrmbHiWduhKjylgPoJiGvX8EzX2QEiSjWcPJgaICKnG7TyJVx
sjI9f0ydtZXb/OPOiSHV+gvNgTWhzfRvljAYBV705pE9ED5tO3eENn3LbhzOweppiXQ5ZLJcFGU/
FkVuSZcmwFzP9KRY1VEokTjS8JXh93GtPRuzlEw5vQQWl3wkficF8ttT0BjIMiE2iFhSsMlyYI+i
fEJN12hO7TbzLP1xuKdH8gS1OL6nXNzDV9EOoKXHzzfqIj7dk7YhkDb8LRimu3dJPUpuznx/fC+E
WJGNvlkQ0g3mYguO/JH8k2wFkgZj1HbxdkUWaNmM6LvhDtn0bW+UtqwT2ENYIwMXlK6qwSkxF81F
cq9PH9+7lcKVCLid0UUfYjqdoigxl7Rt4TuUfmTRGQMMUE2C2kPI2Kr/E8IraWd9AfaBtSpXfCU7
sSo+n3wMltJKGZSmmiX6VpTfUt/jjrHmfFZsgJqPTXKs9IzBiapZKePcj8ObamQffK5eFOVo3G82
BOQ4uCh4QL8Qjk7RenCoU43LQYHW9tUFkRbB0aCVkzohvZZ5HS/mAYxpeI3GwlWmJz2YKt5dUls0
rBaT2ROSxDlFSfeQ9VhFpa/qzn2zkdznwusKYH0V+y7zXy16moUC+XYYmHsBHwGOrCEuxlfgun4t
L70nsh1oKs3ndPLEA+jRqm7WWKhQxaF0GBbh+Z08p/aGg6nJCInMkN4fJmOw9TyHVf9yKMmRMTXO
wCyrxnpSuuv4SuDohCqBQtAaURooFHQAeQ8LCfbTiKoLk7qzvRE+6jQO6rbyEdmSWGiC50URt0OC
LoxSPFqXAua0G1eTbFxXp/aZKDuIWvvrAjRhX4/DO6MFG+72678nlIUPy7UlKHtVVXuRka1t4xDM
qzPvJnc3spR8jaPfgJ1fTlldzOgLEm+i2qg6I8/xgZKMFFVxvc3QV1Ouj21SHIy4OSP6+cjMRzYT
tJnfghiEmM1FWSHPR0exEWHEUoXoMuuVlmSal+iR7+dfqLlOxwTT//dYqfYb0c6mCUCGHtmKmCpm
BFp5zeGpXKCP3jCmA05/fsUIpfvv0r52I0ZEQqP/unUnsikLzpnA2uKvmQQq07hHzc9xrCfJB/Uv
c7jzbK2Ei+7dt1NsJV4gWyDFef1VfbKK2gn3+hEQ2cMCyGOmtkmr+7MwNFXcOWxxwV4pjwzrsOi9
B5rFZ+5Q3r6gSnC1qrtpQi7A1qu1OjZxoDes02AQGDIxRcWsbw91cxu6X14uK0SKSM+vjppHVsjL
mouLxglHq/nu0hRnh/VdXdfoYNKC8/3a3v6m+TfomlvnUlEkrwY63vTiZKCePzcaT7WFzeAaEGAR
nUehrw8a6m3JzfoW1/GzvcbFP2R8j8N+WvStVd8rE6uAC1nTjvv+d93DRd9H83Xm5WSg+vk/jwOk
tZenIo/l4lG8AcpwNtUl8uRBksH0Z4AMIU8KkMpuTQ2sg9rhF6rhmJINBGMfFqenBZxH6oLqMpTE
DP1nn/+0lcBe+D8qryW1lxuVrngiXqY2mDStK8j9dqX/YsTofgeHUIGCX79pLfm4/phwIPjFFba5
cci1Tno2SzZDHdkyCFu5jg11JO9bNsMCqEIB1ejk9cb/sC4+BVs2hKopxgh/6nlyE87OfN8x2WHI
JeS2pmSgJ/gWuC28Z8Hox9FYjy6V7rPsH9xNte+l6V8GMSDW9fA9GYuGy1044HOtk04V4HDK+puT
OITaVJvcW3oj/OUmwmyXoez+dlHuTJtm6LUY56mhkdaoPIUShpvV0OgjmzKCCN+QSXWQg6yua+s5
cpXivw2D9D+P6u87bv8Baek6Rwg29B2qo3rhcBMEaA6zZi5gVwiQMjzCrC+cm693lwna0cpdQq7H
L2RlWcluTpW4J/ahKG38VlU2dsWsJxCO+9ZZeIwJ9MB7Qb9J2KerPyFugm8U1h6cPeNOOzKA6K2d
+s16zwR2pMX58m3MD7CP1DoN8+SM6JA3lmH3WZF676rhljlAM2a/trlEOt6HoIGAK7aeUYS15BAE
NLZcT+dX8RvmkVYI8IA/MTsva+gwT/PRZgO6RQrc812NNQSDKj59LLqe6P0nEx/r+hNcEfgTDoAq
T0db7p/vRG5fWHkD3TZ4PKjz+Ma47PLn5rVD6H7IfpAYk7BBUl/l7QRAhJiVoZ2t8zgmlh477EqA
munSqFHmrc+Zj0ZDZ62Duj0kxEPOzjQ5XvPTYHms2N2oMO1Eu6ZYXLqkuT1BDQ9xILzRzVuuoq3Z
FWANsQ5OtiW6KZKATg9c7BGYIKDLc1WEDidzhWhqETV5TC1docRTyG7utgIAoCdfcFfG6bR9zo7s
1lVqGlQKis5Ku6cvLH+5L50M781Hn+Mhd/ppVs6oXf8o0ccguHzyBk/e1MYS95yv8YLFSSeQA059
M/tE1UKYLU64K6B7SHbmc0G5x0Hv37uWpyAlJ3MqzxIYqUx7jbWUS4yG0R2Ojo68w5IvjuE0hBUD
MOQCKE8La38VvV4bPzNA1FvRhdk3g8bYMrTopCnixKfdn4y9gLl5GgNlvbO/wnI+nNFsPtFMME53
ooLF++LqVhzKmX4Db6PL2dSm8f5EsDeNwrCL63PCnKJ9kpD2MsDyQB4x2JfgvY5u2fXL2Q/T+MDG
RUgo7S5rdOP7TgEfieVGajLypsikHcKZQQoFKpGUp1hZkanqRYFdNVMOKEUAY1/Dg+R0V7lugPaX
9/NBcHjjdy2WJwJ904Ugdkw2LzI74ZzePBGFr6R8yNdT0nD74lQ6ofkqmO6v8is0PohFNJq6e6cN
YuTEkobfYWgNZ6WNlA7OKb4bLO4oZQl65043oiAgHjf4TO+rP9MyKHVuoiQBmXZloGvab8+FgYmu
WyVAcwXsJwf/VXFKbFvONBjDN32XvEggcXS8rfdZBS+iCHzspiazowYx10JcXEe2QbXy4t4fXC8l
9f7u/aqAJ59B8G6wTK5v+By3P/96UCYfSFZ8A+mPJD40wTYpx2g1djf4T6rKuQ650RVsLaBKZMAA
+0RhimPB5vnVrYTks5LxU8J+zNz5QWEF6zr77rSzKl/vDAPHAaBwtF7omgpQTvEE6BIsj6qd5vmy
XgPXH5vUKHjAYDLRd9EqMwSG0yPpS+cjvnigwOeEb66soe6WVa2CImT/CLp0LwwMgSJXT5n9xuuf
fu2AevrgyiOLJ5aQGevi40cw0OgtyTkdIj8xM+3KW0Q8P4QIS86lD1cfBGGiEmJbShbk6Hwg7Z6W
uLhzx8hSj9i548XayaTNNV26QaGzkiPWXSawu+YCT2ZR9PqGX4ZEzOJpFoZYrGDEjyBRgX6HYPs0
G7shxspWxZa0C4NfW6quo/VQ2S0/Y5fBTwfUkz2bYieLmk1BGhk/RWPSnWbELyYi4CA4c3VBiIvi
VU+eyXuAL0C6Mag8rfnyJfERZo81XvH8LOKa+OJFJUXdsAf95Bp0M3bBTxoyXToUkA3dpX6Pz8OS
eyKcue9XybOnVXzk9FMl2y1qVMZKEi39mhYNWBylCNbKKTPh0NIvxGSEXW2RjeRAyolLTi78v9qK
f2KO1IHwT+ZpnB4LCN+Zj3IvuDvDhLoIlujl/36a9hVTsX6sDP1ESk90n1Fb0MBWuvHydFZRllv0
p0eqPceuXTN1T8RT5jVOOMvYGgr1zjTK3PCT7ts9OdLPLE7m1sMWYp7k+K/lEt9lvcBZgifJlayX
5WFsoGOrsRkuKwnoJ+0SKVJwDLcbTtq+bpEjdE2D1K4Bew080KR/8tdkBC3++ksXNQyBQFQp2xkd
n1nGTwwt9cz15Xs3rEeIuPDo2JDRj19sMK0VQIQ+YFT7iQJ/N1RrQkHPCwpscSQgDsOUbK6X+7gq
uFEA3SbZ4g4VLwkwY26X0Qr3+yU5g5kXOKvB7qeD3tTqhenZYqEwszDdwTDT91G0/bBiN5G7ya7q
K5OUfCVOiyU/9PwBHBtfSS9rRdcDD99LCihqkfuAG4UIwXZ4V50I81KJoydmRL2hFKysgGdC5kDk
HZaxig2pfhSwSG3Xe0W7j1bbhpBCvxbarsq5Av2Wo7QW0lxQN4+/k9k8eBu/Kn97E0YYNpFnfUXK
SoToJHJz4fEsIgDvQqxV7lJcpkSIMosE0ySFm4lTm6MTEImzOLjPjPOmNl9b2+Yk23spUmXU55oX
tUKI+BL9IHfk5lugEKOBeuBC8CQMYILkLhlSvk1x+qQe883PqU4aSAKmatvpWvzpwIyNEr7dqkaQ
QN8tR1o5mpZZKPQAFx67D4moI4VhWLZyXTuybgyfnU/BH7hZRs/3MovIL/8rXgJFMcTO5jjrDw5g
7BGlCE7zUU0sj0hI7YRzLMwdETJ6p233+Z/mRIM3TLecdNlh3pVpG7iNKKSQZaTdM6DZNYSrWsGJ
lptB0LXAkf+KUSUbXlI4/kzAmjkcd1hpB25jAtKbPIm/8feHLFp6ba8KQZfkoVxdrOju7tp68N/m
OjGVFsty6lF9wrwWmmXwY9ZzE9IImj7IvG73M+mDmgxahJOFPDW1HPiOEu1Spzv2JWvr+QNEWl25
UQ0eK1p/s+D8qKETjEelyOprgjX++Hjem7o3ru866SD1DwcvQXqkHmbDBU6EK/8fh4A6BlpefOdU
cxqcukWT2UbDPE9u0qQPLua10NDaYNDi3EFKcVi8hIgHMFv/C8vC1CZ6fsaVSVcHN7+E7FKvqz0b
78v62BkCuZjs2t7luvjQMwv7NNy/NbVUJuDwyid6bS3167nu3nAvS+58C/nopMDNX1U8OYdrZpza
6oYfPvvXYkN9sUtZRvWXHDE7n8bbdZqqoHv8HwLOK/3QH2avoxonMZIQi40arK8V21/4HUg/6ItN
HiJWChKeczVbso8puXB8pE0aM3LjqtHj8mvcR2bV6+iik4AK6q84m1Pkp1kdG7SpEQa+IIdGWooB
noNoUPMLaWELtjdZwwXNdO3mLZfJlMZzUWuB2Kbt407XBc88WIlXT71DTE4d7yXw3aML1DPrcLeH
SgBi4oQ01H5D+J2HnP3/+e/AVwQl/4BgZgQgpS+aog13AAe6LanHDIYYV85A4T3W0WwbxamXMTUQ
pWJncIOyjRD4X7Er1UayzjxJxQKOFlP1NGvfBzkUivKU5s8xOT/j49iWmErOAhbzhH2HjkT2RwEQ
F3QVT3pyLt2MkCJmTdH9wHYHbLm24blooKPIdJ0kKreJ+DKRNQrWSFOl5Huy09djkGvrUH0tLjsR
7n3TJmdTu9ikkcXfShGsx9bcEX8GDGbMu7GE98j2phN92JAxV2vjGe3dqOGAZnN7RIq+nqBmR4oO
d6PMkATCHXkG9AtBApO5hb/SKwy8etMMWwKHdMZaqvJItZeN99dDFDjTdFQzn0iQjh+xNK9M+K47
DRxJ27s+kgysj7uYI7vyNhJTpi2VK+THuuIa6E2hghHV+s1bNC3JdWZ5gAKzzN69z++KFHBUl7nw
imn23fVrrwCs7pHFtVbE52sw2iodwS0OB21HlFLQWX1vHJ4OG7qj5OaZ9rzFTMiNLIrUU+b09kvC
VVdHILBnG+JIEs4mt/7TZanBKE6z1Mx80sjBIYSnSBiFDXHi0zYvlTp6DRcj93kQegjAUsC/hiEX
FA3YurQWaNQioKpp/nHdrLowHNSnapixE/Pnab8QjNT09CKG7RZru3c0VYimszK71aNBWk58/XE3
71wIINAFdcxWch9N7wB0Nug0q4JhIethpkjJ/FyDxGnAjCuEB4ae4TpFtc6oJXDeozjJa8bkd+xU
yDMzSfHEhjy0dBMNVE+hV5QS0LiZkfkVnXgG+5mkZVIp7Gr34iIIE8SNsERLDdCWxfhMX/dGtB9v
9LQTr94/RLpcKyVZc8qyIamEyWCmfsE08bRDZGBEAuogw+hgfk9xRtIvIejZxiHRcxmbfLv+MTp9
/CEExg02w8bweJ5ZUQY+O+HfZpZzFbnjNAYdfg06COi6FgJgnLP+Qvnha4vEsZiP1qFncUJnQGU3
hKto+5TeGS1Ln70n4rDiUwO4nKcfDPQjmTMWMeXJuYHNkx9x2etpAAF1UkSDbV2xdc3XMQlKMdyt
7xH1tX6qijmAria8S0m+lw6y1nzULT2fRYxM7O7Kg0MQ7dpYoeNNuHXnwfcS4qZtKtYS83FEfj/R
eyr0StMIBqWPJ3vuKKWOhESnXvsHtzhyAM9MYXidlc+KteWiqqqYTnPVjp7RwVbLf6deZvnTESs3
Ubs9ZJheWGFxVrZWrtqkxyDpOCozO3DCTe9/zVahPgsAxbCQ55pNtFikavb60NF/KFAnqFMwvuuD
Y53AYOlxd0BOk+/ozDa7AJDZr/ZwesNDjI+g6o37hB1AjpMDUndahRPyXFAbj0RT1csQaGuUSiI6
cA8JzaSINLNmD88uVnfMTSEUgaMMAcVLmkHxLZ6OHNUhFbrP8fovZfl8qxEm3x6GXpLBeU1J1QKI
0LJRtiDA5mRAa0K8nvqaA9OSUl0yzXZsIaZ4eM9gJjDywzqjkJsxi6MZD0x2hUFplH0vP4j+rxpU
c8WJb3r/6GjSLzVtiWb5K5zczbKW5NMy+Zy7Zt8OztbIPVajWdpzq22yAje/wvNExrHJA0Edyv+w
WYePG8yZE2Jehrlrr6rnsXI954RPv2r8xxwccbadPx9yjVVnsNIHIt0dhAbqhLg9op5CHrJiidky
6a7VBO1UzStOtEGvoDPvd4ojMcg5bL7XeVf982L4ncC1spXpKnF90Oy8L6Tlqsvh2eEex6oWbDSC
ukbjth6ReA/k0b9qaCuK5cgoBwXeb73ZH0KTbdS5wubeiIAS0JwWfuWK7CKwfP9k6s9o8H4tWn9V
pmJWq+Kl6jC32jLqUKwLq+iL+TfFP08jNS8c4x+w4Pmf8dtnQxNWepB8EAs+ZP8ADqfJgHrRr1hp
YnzQWSppkseZo1rMhL1oFFZvyIyVTZWhRfXSOMyKax2qMk+UfDlSXWh0eD229Ld77bjTLnX6w8ou
BymsHv8H/AITyE5ItfQ+PWYqN9gSbA+uibZw678qm8abYzfPq1MHrZUqOHKxoQPqwmHsPoU9gXCF
vZStkhDVWY49cpRPFk38cpcL9JmekSWzrldjxhTxhGsff7TV8fmXpwHgwbRf+ANySJqgcIAk+5hc
eY3MZvjoHnAxmbqcHt5+zH66Njtbhv21ZbCysBlLIyi+mSA5ZLUEgQ6UfYSe0RaRLrrDAptpVWGi
YEnc2DoqoHd9msTilr6mvLpGG0YZ4cKmNfjrbBzkTjIK4uhwnmqJn+u762+hXAoNSwVy4CSKa6A/
j0XgtLhb1k7ZuysexCKb1bcJOWgmvuCAjsFq0S0d+kNXCfbumWwCwIxl/neGiangFHNwZzh2yE+y
qb/2A7l2aL+ebO5aNEjnhePuP763ZdQyPGqw46zL5bvYLGXV1IPo4/uMNxwY+BZvT+50fZ9W8g5A
YgPnPB9/jKZdDEfZGQ9TZ2/XNIicG94yRaNbgvIhCZNYFgM/vVaQcTnnnWPHGI0gDXln4Ftb7xMX
bxAX9RSNQs7/wV/8kmUmUcxVT0Sx7pB1H1nz5WblAZ0Wv+ySHGrVObQRwCZvdSDugwyX62mf8Cfi
JYi4qoxTpjGGLueSW98YTUu45D+CV8ZF5wonQewB9K3lPGU7LHe420qSri3gQjlmOGxLmX+8uxob
T3QfuQSei5EyUE3Ni4CjBwNhWaSPZaSNDIfawmBbRo1Ts5QJdvvMjVSeXr1ySQigDnvNpWmLmDxI
vU3gCPb6BdMmt6ypkeuqUKM5myFR1f/8j1AiSHtQikKbfGPuE03GzOgV83ZPBLCOMQ7iMa0E3HEu
yAAs8nWoW9xvQqQAYpWhVJMlvxMgfDe0yhWPDq6ZKSDz6lyP9saWpwYd1qcnWw7yWid3hnmi88+8
GYayRdrCfK0pAM4oOOpnTlsK95lwyKTX82xCYVIolo71i2Gy+RaemhyYQf9lOsWG7O62YpUKcqp4
l+Izn5EYrs7LoZ5qOHvS3I+8t9pKw5blzyMt9qYYIi6VH4LPrP61Lc3524knfNwiLriFXA7vQiUF
k2DlnwzpGHN8NLMyXgCDX4rr3836ic9aNqPiZa4da/cccJVedBRyrtnZxUoBQCGKqMIiz1ieep52
1euZWP5/L4gij/lO30Yvg7fXFe2h5vb5O5MgdayDL2RtBYPaCfHTvWDkcXN+HTT/jGE+Cxol5EYv
+H7JkFMgOuVfERmNo4TxOo3Qs4RWar2eZzUtrd4ZV1a5ru74oG6dbIlvIeFtRpvnsH0mtq5HcXTQ
ve2cVd8K/HX7GiwT1SWy4DjtBhAa9O2Aw48qK2WAr2Dexc13uvVPOOrdilTB07KFkhUf/f2cbWy5
AxxiVdCkHx0u9GQFwlRFlJ8rezvNkZbnWn6+zsGjA3+DdGkNVF5dcnfnaMglp+BWZTHPdh2BtROw
MVkYdLTYC7gvj3IhYJH9srtudJ3g0FfUvuxu0Dh4RG2TvJ874kKOCuWNLyULaFZikPoprIbWm+nu
6sAdGnM9e8y6uE1NpJ+rYC++CJdftqhWZNRowentSI7N/x/N5h2Uwbs9KPO6HKXPS2eoYamrSmqd
nj+c6TA7mG3h53qysJF6B7Hqs517THPsqtGe2vSdZYDQprE1xoCkgct99nBA/HxGLvPiZflDbGct
xE14mQDpGRopVdySrzu3bpXNzF9iMDoLZlm3r59ypNrAiMbmjwoGXjm4emV1lG+CgghBl7GzpAqH
0QYq/FXDYTIbaRIuEdCKxMoBARoM4UVcnADZ6gqhr6o5aD1J5tOga6HCNWH93lMyPhVHIrKkRp0h
m0UuWJtAn5L+PJR20MAOEnKCzMa2bvmSDYm3X4OLUqfv//SzssWqwOlE/vGkxQfh9GO7/3hXiDx9
6bzJvjFy9WyQvn8m1lfHtemdxe659MgLdOkDq0GgPueUgKTj2R9So/++FK55+v9qWiegwO60uV5i
XIYXzC4CF04dlbbdwouk7Jlm+aW8E1I4fGXhqL9FrjygMJt0BmWkDhMZUfsoQJTlCa3E0dhQUNEW
WI4faoix1lwOdjDHa1Ku7mocqfxSzEwTpvZQR2StNcWbCBhkIpBh1ap8WCWtQek7xYtNW+kPxR43
PZTE+mfzh9GhbGSWwGcYCqQ1WvnW20LN5ZQREkX/10qQwSZuMtv5pYAr3iZ2KUWH3CrR7qwPx8rT
aNY66rOn3exRK3lRewRVL1SRMSobWF17KRIgdGSj8kjYu6P+5y+so8KdqF97VQALvykjhwKkR3Qf
1AHOxlB3RHtUQNB68eafSVPv8hVdt1ccW97ZhiTKNaA605t3iVta+bv1M0DEfqyoagQYdf29tXcd
RZ7Z2BoOv+0d0Mea92q56BprD26AqHsvQYsZQJP7wJznw9GHBeGKzAZiY2uCwcoJnzVNkv/ZRRGF
ckvLi/wMUQ/N9aV7Dd6yvxBui80rzCsc0VkSE2Pf9w71iEarjZlbtD/LqOMFKyyaks1Evo4yS+O7
wk+G/neUHTG6ccDlOBNEgzmDyaX6F3YUQxaFhZwuxuds3lk3PUzBO2+memFiVIjZTwyqkbiU2mQx
m2Jo8lkUJ1+LG3j6wDl4hvgpY0WdxgOGxADSdokAoM83xeW3nGgZK3XUNqwBmhx40raGVidmEsF+
So6IhLH0fAZFekFJFXpGMKN1r35fdQy0z6zdgMTXvxa5cU7fbQ84rsqmQWVQwGcC/5DseWxps8Q+
EsXiWY/CwYwl2N2PnBnkMjGea2vgW6U6gMiP/HudCtAei6HZ7fYbRfHLhHr92BbvMsPdNeeQUxeW
EOCEDy89M4fnAgzmTntmdBfeqCYnJT8l4uWdSQeXhKNH80TRhlbxExOLicC5t+vgJFtuN67/+eAD
YeHCs93Akln/xn43d+Ts1nbyb+DL0Zn5nJJWih5ltKcEpt2SJnegeEc/fP7cXfRfu+GIGj3XKipi
trf5p12FEJZNeqB5LkSnSsptZUw11ci1Kkdrnf1mJERiE2qs+Fp5WJ1Qu+TtohqiNcGD3kSVxpWj
O/0dvizX3mP3cXk0unaAJouXfaMuLVHjrfcIU5XHeszVVYUsL8DJ2M4b2BnvnJW2iU/FeLiYhMpY
HyihzQs32cBpneUWtQEaqGO5Rm+P5xaS+FHRP9aVTJ48pSO7tZNpNPXbCYi6RHaUjHALefObj16E
v85ja7o5zAtH9367H2tfL1+9OXuR/4V/D4eK1T0+9Zzi67CNMgD9fXQMxJq0YVENz8fww+jHhnTh
EzRZ11k/iEgkNVmTlB2Q6nstGXtQBRHO9wtJ2F94bKDFsMdsac8W7wKDQFxvUx+oOHANk+7fkmys
D68zAxTv6Oc3/7r/yu9/F9SGudRH/HbRd0HSSLCx7wZZyy4ew5dvgtMQRyLmBQGjS0d2EeWHw++4
RHWfcFgtOk0paijXTOL7tR8BpcopwCh4Ns0LsVXnqFj/0C367cq6r1esEKuyV/NBSlZ29Mj6rG7e
HJDTNIoju4tMMCmkNrQzmFXk/fK69PJJkUKg4lairZxGw1q66vRGALKskOZa7cZbdhuUb8g0oxhZ
jHKoeDiE2NL5oCQdtLpMmJAvtUjSm19nTh7l4o9GupBowyTgrYcWYeMN69fJ0OiND92LrYiwi4kN
hYn4m+JX0+SnVOagS4ILBK1lVcl1MlLEdnmOEY7pdTSntI/S7rZYSeNWef+qtGpoN1mt0kzvDdUm
cG8sSqtgcoGtZrJ3sn6tUrQBZUqNhFhS+3xVv0kdWMK9oKBm6ORKbjy9GepP1WlZUyJpjXC2fj81
I9QtLW2ybfj4hljRDqPMw1gOwPAs4xWwtXOyl5kQlM6Ln5EgzLnUivgsN/1Fvf5SAoCuF8S6rMHl
bI1oHjClIovjJHaDvSrih3aN89k+zb9Nfp/9EQYscDPcC4cxM/m+kk0kka+/r9+s2+E3d68PxinP
l0WEIW1jW0Kvd1L7AheVfqAb5ZvrnzCcmZzBqw6XTBuoe7V9YpAceAaRw/PU4tNLGDjta7UKf7Bb
3fuBqq5gwKjdOyPutDAleeubAO/Ac+0yA5pYbtde1ieYdAf+xWrLgFcxBm4ExkSM4sFIDmKHH+ir
m/uBlJr4Q1pAqWsQdLk3c+ycp9Jmo5anfGy5p8mVsXHt7T+XwtnRUCw9z3MB4zh4yUCM3bLrZ1CI
LQXxm63OFj9oMyf2Fpr7Nit/5U4Efl+GBHschvWsZp1raLIedVB4xxGCVb9o+u2Z97MAdGnVvEvY
kkN0BCweLQDAyYpWgAHNK2IKiyhaTY2PTFI3l2YIq+Jyo20CjkN6yoobtraRzOc7g7QUfhHFk1MB
39k4iKtE0tme9ubzXuOkeYI0VVJLv+d/+PXen+g8HQEtkfsODUVHKqTgWOCeLu+oYW2t+kft36eW
7ULUdhEJ1Ys4NDWy/JOi9s75b0Z9XQx7mx2WeVeLJX1ZgOTmHw9WlRvLiZgiQHQgElDT400Hmrpt
bgZLarN1RDU1CWIvdnnADcGpQE82gIA9fDotBYdhh6jtVprUtRa2mot6Jr4fp8IpngHNKGCVPXea
Uo/UrtYo14ouDZYaTyVAou2ryTrjZuKLz6J90HT/0CK5uNvSCm0xkptv1bYt7tjDp/gA1VA4hfN8
RdPrgbjdvm1s6TEk0B/jydISX6gmuTZ7MVUsIrkpc+bODuAK75AszPPXqXM8c1q9wLl+ZG9+di7X
AJiL46KyaMXxfkOypqAGzLPeqreyZ4KZEWnyiki+jHwczS08SJpy8X7ywAy4UGByoM/Xc2t/sIa7
O9D46ecDP3FjYsiD46JhMohGPOD3Swr8Yko1/0u+WkKiP7vWLfy8ePlZFmxzFr9hhgaNzSGsVtn6
KCY9SeSkGr+BiHlK2cDSNh0J/dQ9+kmqvEQmwjcFB+v92U3muIyOyC7ohHFRDjB4zDoZ+fRrK65S
2YthsZgKvWBEzsMmkYEd+KeTyAybJdDUern/t+7B3sURqEOPVAW/h8ewbsF1pksqyDFyY8hYRRQA
mtxCMhSZhbts9PUhF5QHIHUhvEQJXzFf7Ql9rt77SEL3oxocaosWSsBzmnDgBN1yKsThBix8EHH6
dN8vB1QXdj8aQDF/dOLcBcoYgW2pISPppt4mjeTvUsoK+OYhRfkfFXonYpsvQAyoHBxeI3QNesdn
oXaOcgurDFFj2WZy+MuVq/axnkDF5PLC44AeI3oTVEzyrLAjoZS6vlvsc0qadjRKSgc6iifXtDXY
hm7tZOiNzEfP9e/+LEHP99jX0aKpHGh0jD1RpRS8xuvpS1TXBjC5POeqIYsPkLX66dMRbwLdOkgZ
SYHoUlx2XCJImYmIiCbQ9SFEdzFFp3F/q+thGlmPrpJoX1f3qz9rQZPjmd+Ksz1PvMME7Afv970U
IcBB9es4b0z5lRQqbFqIR77E9TxoNClEf8ber/ODrdJBCc4lBQ2pw+NWoduD/YFiF2uHayWY9ncP
jmjAA+C1QVOo79xozKTNasnVj40RQO6fMLarLKxMh494S0bhCEYJw/eE/mnEx/Gmntwa5ri0Qwe1
BWthMMJC6GWG+gpT4mLCrOEu4SUoTUGSGDYhE4AlG/DuEoFJr87NSIMfOoYhc7kj0B7B/x5EUIKy
fyf2mihXbok13zgTzqGYzi39w/eHBd32IGLvY0I5qOAnZKyKHXZPz8povOwCJ1uNpjjUGDe+oyoT
apHLGeYQwegTeOGER7PKkL1+bvh7zNPwVJ5QCM1QJOY6llqJsYrq5MW94eXPjWXU98sMxksZGxE6
wyxaxzWgsMgAcdnNpBlf5GlJdeDiGN8+oFxXqBhRwYkInC4dMZ57EQHIYBamLWFclALcSOMvkxu8
rkvKwdJGD+pN7Pfv1nVg1CoV1kgLNbQtjAVEnTaRGULeOGX6LMYX/fgjfkgfLn14wzQAUfHVfxdK
fQTJd9d25Qm3AlSNJGDs3GdUn8IALU0OYFG8bU9N/mnXsCe/1w55BNjC54c+NXoNFrbqXAn7QbUW
Z7D7S2K3MhpXQ7o0rRY7R8B5tNm8GPrWKQecwHXaKE/hnoRKA11qTYtVdUqe5XYv1/SU+X6OGjog
g6VopRAqo41yJx9vgT3RWa5UzAPC+hC5FFAYAlkELbc1pALzRf4SvP2VgfcTK1HxpH8P+iN5Vj/J
iwbygcN/kLeyJ9/YXN4xJeiNR4cxL6NXHT49OQ4AQ0r/3bhbYC9SdBZjuFEfNNzs2J5gyU88tGH+
0G6e3a3NrHxfdhrPpy9szjuMbNYH5FbmMjH2nOF5ToK0g9Om2UQXptAAqx7og5fPTOziw2sYj0ZP
0vrhm72WOfKYRzJM3XLbNUYxsxfcl85+HfeEBoHV8jr/QioJ8HN81wPDv1+8AXhRueFr2lR6PA8e
hYwO3lMwRbxRmWXOIxEgMIE4wflvg8e5wyCW7YexhM0NaLlLf+S6FfZJOAKWj6eCTU6sfoWOj8N8
fwhYCo2LzTlYMb8SnvM46dFoSfGyyBjlkNxyrzMOzGEfuLOej5toE/Tva6MHhYeZ/BNtMeAOGVQY
le/i2P2tDanABxil8uB9esxYVC5Xrqy9jz+qsxxlNz7yfQwEco07iT2xGB+CTCCisFyG/lyw5rxo
vYIWTpV6kVFP9FP2EpffG+jY/iIbNEzHSqwvGU33Q/GLyrFi0MkEFNFaL8Fw30mlNCg3EasNm8M7
hxtazLiAnvgXc512DsR7AlrfFf178BVnaN+H2+dAkM+yHmQPTwoAaAGaKKcwGdfpNt/TzTWFJ2Jc
b34+lcwgydL6ltRR2rKBUofw9lQYSqjK8wh6R229hSr/nOVlcVvLAd/GtwMYJTAoW5RDwb2IOz8F
q6SNxXmXFU2nbGLUI9H5G4rxYox470B4iNtS9kzXHjul5uUJVpMmPOpDR4q/H8j2qw54M6Keil68
onanGSSEOFdLeY4YjZfOpsMzJuRR+lYvKrLfUic1BZQ5d2R6S1EkNAVg85lzcNesv3t9b3TGNQJZ
i3FGi3xmqpaqwLHJetPcHAxONuyqMwEokLZXVbypYS3YKh4tUVuHDlZDxRKWrh+RXdSjxOLx+kdz
Qcg2NDZIYMCEjffBtoPevsAA1NGvywkfHTodn3IyRiRpG3TOOvIZfL/sOAK9fKx0auKcQw8Ulf7w
ViaHvAxlpHeWr/eN4tg6iS6p93VM2eAzsx3QhGkH3DNuNK7nBMgK1fiN8DbZnwyNHIGjlkyqClFT
aQn/6gBb2C5s1Tp9lXfEp8fiWwGvxpEZ0UrEoRCS2F4tXSEuKA3P/kLMpC4wojb5FUd1HGh7JIpu
JA38QiwpVwmiW9vwC41u2WC9BPCG8JTeUhGQAjwbpm3g7mBx/R4AF4ya+KXS0D2UEVNOC7Ef7Cy/
2BlSID9iv/K1FH3lU0WyfBCIKN2mvLF1rBBcXgZw0b9Uj+xDH+miPic7FfDRwFyfnlvuqvN+kpn5
TqUaTQK8hNGQaA9xGsBNt2CMugTeNo6Aoo1Fu8vjU513pXPZBYM3zThutFYxOhZOje/h6Znfvoer
lK2Xu6xxFBDSTO5HAlCWiBAHwTwq7ckCJXb6DE1ANy0mK8EA/3D+IFfqFbSwy1DRvtqntkuJLK/1
Hq06IzLEfIPDNFC5DlrQy1A9tFQ599tFIhbDMg05qiOwMRuDEbvoqoy+iX7kEaXnqFMSSBi8Ec+p
whsoYuil876yAq04kEb6e+Pk4YVPMvrFmlFf30yYbO25vxhnWxMlzbqgfVwGW5Kvk8JK1WDloYk8
dpgl+Tuo3CRWp/h98cxaQHfQsrThxF6V8c/rpt5RdRpNtSrfOpIx+Em6M0S7v0o+kXMBtNvqZUGQ
RG1OpKjT57lMi/fzKg7bmDAADa3Wj7eiJJM6s5J/gU/WZtLo74vzp7qWdh8abPmA6v7oPRCSq7mi
KJY2H4vWZEXQfgPoQQjdSQKhw61jt5K/j1GI2EveDBQ2i+G2Bw9UK/4zVBz+snO3+Tde8uita3fl
VyG+6Q8tGBfGKrvVWxb7BIjnH+WYzrKLBT3+TFTh7w4+fp/OkFa6bLL/JCo0VpKWs76Y9UOVT/Ng
uTX6iYRTUdr+9VbivFFKrz6WY3Qjz6WxJVI6kUgI4drOLK0jERIhdS3JHxML1Aj6ISU/eErcRmsa
8ztaVpH5+RR/gSCX4w3KuW2uDyv+m5A69nfjitmjU/C7o4FKCwkAaZ5jeOECOMwJvXfB7bS1NMCJ
ic9nLf2dhaDB6jEa5QymbwkB72wGwux2i4vXlfXvCLoPJssaJ2w3H7Yr9RoZV/hVy9M5D6VDjuRA
MDi1S+wYonsu+7+fnbB6uh4BjO//Lj/pvj88evKchFWgN59kNlYL5KzP65kylryyr4y5y5jRE/BX
IdY98/awt7oDmGDyOtbXL+y0p9+x84YXnMUm6MaGSRRMJxNx0FRzQ+sT3zbXdqXj8Np8wpyspIBG
p8egJEHSIfZOM/qxFInGikOvNOt1Z6HeaQ7zeCegd86x3Alg0ASMhozWP4Ox+5/Azl8mfQzTG6lf
X8ueddSxEEXAEqIP0bMT+109fpe4NciyNeu1rpgsggEndbSgB47TE8hW7lhzas2YrCJU7cW3Wb2j
oYayczKiIQliqD2kUw5Knl//ndXk18ix5vELjrhzsoGfWuGiU2srib3Kx8wijzgOSOqutoNDe/Uz
VW4wB9+sOLCNWSAXvtezBkbfNPQuMPTL3a1vV2gXVSQplBqE2TBZXHnqMpVb+OvuvYH8coCxtyAv
5ujZIiZMX7/43V4Zniu+e77hJKJkzzAUDRn3uWVMlIOBQtaF3Vq5cV0FxpV+8Y8PnoyQqKCEQoG2
PClOo3DORMHcrcH1oY4DV9VtEubneCTbeqFN7oA7bHSdvICSCNyDqSNaBLaHys2Tf0ZagKQ8iPGy
9z073ElR5R+wN9dUicu67svbchj1m/WLC0lCX1G+rNRH8LfoWTgqs4KzvACfmEXokAh5e1f/WS2y
dnYhxPoRfzjyLKYbokB3NpL3FK6ULqVJo8ex8RQh75Zp2QSTE6Dr1TV84lM6nVu/1H95vf8mHTow
1pBv5TghuoJmtcaejXnvFYXji4fyon6kKdyBcIr4r2aFXUDzsxi6mmSMFwkVmjG2S6NJ6czeOJBU
h1NTdcl1CurUpA4JUUfg0iAMp10FW3zI6aE6Dex/IuwduDyomT+mokLbayljOXiFZJboMMAoQbfi
0jYDtqTNWNd5TT2Jv3Y2d0f/+8kDnlIjQ4WJ5t5YLtKkic/nlebyEoTUWSnJKkTcaN1T5eGvC2au
cMiB1eHMrVEGYBsPbb+2rgNHvbW+hn8JgVkRG4zTYVlz0q1k9TBAfnU59rPaaovg31gr8QcOgBD+
vnPQf2IRubr/6Z+qrYGZ19CSywNB+LaCpCyVhuDG2CpRUgz8GY9EbMBJbbL7yRuy4JBCujTA3OmU
2IJzx5hPxsKZ3ZlJ488Z2Cd2JJH/JKzVxztkc78dBXEr9wni+T2TtdHXSX5lpXhNwqDSmZtzh8yM
y0KxVXNmbJx9IO4QNbuQlK7F45n45Kv9zDFCDjeGLsgY1RL3SbFhyojYx2Utb20AJUhCedKZ3NOE
NLeDo5sz/LCiO8lySNqSawFt1sp94IGN53kUOvnOvBQDfKuSytjRWRV7MjXItviO9f7shNzFnP1U
Cz6pa7K+ryE/v8qiZrFxN8eYpIO1LmzppCyfqT9491a0sYjNej3IzuRExAwua6np3JAX5OfrAubv
5G60TRLjshtEKZzPQ9VNZXjQtURzU5/Q3hcsfl8utfFBMXfE9Mj1DYpMGDlibp8govftxX/C7Xt3
9GR6I/3gzEroQZyRv6jKqFfZK4+Ra4uVre9IxR8C719bE4q3iGGPCDCg+5IiDSyfRStqjcOR51iG
1yGD1YTTW9xJzuv43ZcMwB2dGD4rETeNZwIICB8Qpy6rUt1e+55D67sDwOkiXThjMctmNo+Ks8Ay
LJZTvK37wrShOWXcE60Z3eFcnZ5ItKd59dqWHfZc6c1WSB50a05ufs4VphdvPNQiLplKUyib3s8o
zkfK3YFtwpgvJqJyaa7VwJRuoIIhfAIw69zY42ZJKCGUzdge9c8w3lV0GPXgu8n2YRPfhIbv1e0f
SO6CllGHaSyzmikVlWkAEDb60MSuOaOclHNxzV4BV5K/l38WJxy2cwR/CJbT2nTxmp+PI2OBxPYz
IrbbUbvAvYl81m1K87iaZmi1j2kmstwaJfRCc6AnRKUR29yVceWPbMCOBYm7vIkfpKXei/Ck0AkA
OfW0NNBio8VTV7sEhJ53umph++pUbnPCAaPFBdlNgoWfPcj78Sa18M+k/GzCY9+8ZkORWulpZTfv
SAJ1/evW1nTp7WzQbD5M57xyWgaJ2gWk6nEsJSIoQp0OPB1NZdThPjoJDk/X5ExYiE5E/4WGw+SW
53YUMLPQtP4abafHt/zFzXyuwge5npg75W/lhcDClDUh+kLNBZks/Wlonz501xP357fWSyoD9k5m
FFf5XTSF6sdyAyVfFK2ktvo62gYdxSHg/PxvOjIsXWaN4rsW8AfI6j36klM7uu3d/9l7yjhcT8WR
KaTiw2c81oNBtS4jYMJHgIhXabhD4ZKlf1mZIEbCqZStrC4vfaQlOtXRl7XwFdDCeCeLB0rEoNze
j12qHb0VodcQwYzTCtC6yqLbRkda3rI/KMZ71GnRBsaYcWHHHAXywY4Z002nz7+aGZuIF6brhIzO
MVqtTEPkDBKwx96t86SzlMfXHJNto//21Crt+Fcx4lwLCX2f29672NjqjNKNaBC8DGB962sgRrVp
0cMhs5ES0ywbpmuu72hfe+gtgvZjNHo8ci18A5yCsAAIiPK9kskh2SmW8wBneCzGQtxRgyw6Eb52
Jb+BKWfsiMTVDRYxQvrBVleLrn0Lwa+vadwXYjvWs8eQFwUgnKB+q3vO0/282MgCkO8EYw4hNYZ8
Qheuoj4wrYFE8m811qv0Nb7nMwMsW/vAhnoBI4oJ0J3QUNI5AUdRVQPx9+9kTiZESA3P8ukVdZXk
BciAwOjw66rGd6oaVnnnqG2NEjSbH6SiN1PVYmxM95lp3beyEwLHx1ovmpjDvquoqOyJAZmewOjc
ly3ms+lg6jHN9BfcL+coagW4ek50kL5yG0+qByP4VyRykLe7xWXeRKnGpgkMH3l4IFoXKVtlypjw
jym2oCEOSwlIg9yG6rTOsX7KX+X3e0CdbgP3NYcvDwUUC7eHlnvjuKIbldJ2eTFEI6Nc+8/wHCFY
54bg+ub6OFCs2hpXKaWUSzvm0YCyNQAWuNP4YDsaf+Y2uBd0EpWgolM8tm+pvH3E1ic9FogENFPw
y2rYRNGomZNABhT6m4odjrLqfChNbBtYkscFRM7n3gN5N4QZPAOFgZM6+QurLyfqXYFXsWWk1n00
jH7XJ3LZQOAk0/vhWsebf6jrqG6CmhqfWXFEBEYEMqFk2dJk5rLDBUZizVppNV+gfnyAD4uNIpjn
afKDiHe3gHXPtvKyaotMBfHceiyB0C6u3CE+GDtj/VEZxnLTukJnW57GKQBmh5lzRD3wmBre7A7u
sr/Al8YN2woKaORs94pYUqDF5cM7STJ5pLOjyjH52ojnaaqOMNahhn5KaRXGV0EUnZ8KRL2YJG7H
xf1vVs8CBx0f1T1nYXivUPGnixfryDOz+QXXvnTM7IC8tcsm2MlhHoXNI3OVvhKnWtIl/BtJY6lB
+QiYV1leOCN30oyCao5in03wFXT73fLoJ8JbcXtOiF9ZwXID3QriKkKZsMD+rSM1rMSSeE0QQFU5
O7Y7CeDhFJaH3riL2Weze1sy28Bx+yHpYkxzHZDo9VCz0EZMLlll9uvcHoDzyUWOO8BCYyPfi3Rw
9Mj154MtYov1NdSCvIxSRZc7rlTJ0IMnvYxruvQKT+VFFP5gAlCt0/4h/Cl3RTPxPKOq7QMU71M0
SaRUVp+fb37alVRijZBPzcAaQuQb10u8hxvyXEi6Pfs5LFC4vlOKuGa7w0Myf0TB4qW3fZZvD/C3
OOLdEDsqRC/TAVI2m4GMhs806hjCheSwgq2pKLUYEVr3Hq2Ng+hebi/6zIkEzkuLgGvWvrJRVxTt
lpFvKmsiwIedpkUKyXmzltABgYca/0NxazRC8FJ/WI0NHIW7uAtBK0nmDBzNjgiH+L4yB3r/K6pb
vnx23OHdcqp1i/5YcEF7Vc45I4yBpwoj7fuhLfYJCnLPXUhQOEBFUdHjRUvC05cUTTv2ZOV0Nr7O
g63MaR/b48uv6q5YdSE+FkX3mU2kkBppdY36fdGkf33aLc6Dt0abbPuFNI2Xzr45UQ+K3KIpLHJx
rg8ZFHq7a+8KufiJNEsaZZguBsnt1UAf+dnC/SX84t0bprFxDmyIFPbYdUzYMv6WzjCJFhJpLgey
yXR0PLtE9IqMPV61bKJPScxDwimQzOQoJ4s6khQkvck0QJiOkzGHPZLLsz5t5wc599NPaED/lm91
6j851Vwl59/+HZB6SRlwipr6UmFGzRv9ck0J9Z+ukayjhcRLJXK5YIZtgc12znLMJsjCYwkcvOT5
AWMxW6/c0fG3/1DR4VsJ+ARSyJf8YEoHYix6owpJRjGgXqMCdbp0sphhPDi//32FSM8Q5wpV9eUW
Cu+NHBjUcnpjWFbRw/vt92+szl0ItR9mUo8PlaYpIUshKJTnsn5dk3ThmfGT0bXtqpr1xnOxJcnX
533MrcYxBgfyD6KeM0cX0+3160g9LPdwcYPtao7/AlxAy14voW/UJGxVj3OeGh1RVTBOgsZR3hjy
S3hP75wOcMH56EoFvSUrh8835Vxu5LiaDZJ3+S/OBvSeZsuNW35N1l5hc+1qVhPE1wIFtD6ez/IV
wLdlOSBl1H8S9WK+tYDEoZalycR5WQUPGjZ6/1qdTOLJYxn2ZwCHMHf7Jy0zmRaYKo9utT47XjpJ
BW16UtHqmb2gIt8F0IRmiVxwgh/g+EepJBABpcyfD7nnzZhARp6sAMSbVAorVdjKtuZeqh/385Oq
IV1vS2uLpvWIGhgb48wBjZ6a6BfPVvVBe5boBaf1bdii3kPkPrLcOHri7WI4XLOztmHRO+nbIPvv
h98vvkt34szA27f6qcMj/2MZFbBS73EjOGWd247wbLuS2pwu80LLlkTXlt7KbRTZ0Y4aLVcwv40R
k7bjXq7CZz42wCTdCrE13KvJ40LRs35kkjBh764jERzOa1oURjhm+XoG/fyN7tA5r8ZO7OTNNSL8
7h5lpjDsYSycpihQojj8faqB5xxUpIBqeUZbIYML3Dw/YjjmNsHQyJCLNWXmeabFhhzaD7SszeH7
a+HDfKTVxXEa2sAN9l0COoujet4+clkJRruLDNNqM+XlyeiNJEQ5o3qq89zkqmPi2PPlmWDlvXrZ
MvCZ5iIfCvxiWFqpWMJCDpdWm5bcSfueGDI0MLdlo7wvjsHWHfQglwrnXzyEFJc7cEP5enSfbNrN
DXVNpBjm9SNo4ecVg4WX/+K36qNW/S8oEkr3B95knQN7S0jUUSCgGjNu/QNjo8OXyrAfXx0qctrA
irvVYv6CaB7Ck29tfjWRZ6qcdXeYnyTIAv6WFuFKwB8J0MUntNXYSP6kgkd05yQ2d5dnlhpJlDZH
pefsdhXAHplqzeLpevQi0FNKNJZdOJ3HzzhCR3hCPVeVZBHAlqWVLuAhAIW2BbibChMIA25Q5t1a
bAYqGTRoi8c/0QR0N7MVg7Wj8/11Ljo9oYTR2BJjG0KdI+IELQ7I3G0pRh+TCxqfS0HCqwWqmtxC
2Wsf2wkvPyAbQZSWR32YNw1dTVtvLYQhcfafp6zNIpLGrG9GIinDxnDae2JY5OWxJiuMQP8jilMJ
jtMN+LYLBFgOoxlZEdHfWQrBSFibcbk5Plkuyno9087iB2RMZNnRJcdfSZ/3QXdAzMtAPXBQARJR
0JsoCdcRVeMJoStyv0rJfhSJQacnPXq8oayzAqrlmVUGfUQFTf6wrcUGqWwxI7NtVQVt6Sp93I93
+IsQ7S6QTSVBXbFZj7damax3Xv2j8MAoZLH/6PbRsScQ56AKW+HPFmNUxkb6IrUkvyMnLmQYAC9A
85t94QF4PHUqJHR3anvDvyAQ+uapKdcHp+UHJpgj1LQTAOMBN8w/yroRUwUCau2xuK5W9Yr3B2VS
kwFmJ/o8kLnG+DBa/c14lpwYL7SbUx0lKUcBpie0ovu+pGzkaRe/qYzXEEV4CKZ/HpWp0qxUodze
jC9mEFIAQetveBeXeiJXKQ45YyUApasm/M759SPuYp/fkYOYqeP47tUnjM8fwSRXxhBs7NTBASoN
GxFnL6/5mRBORxzLGPBiyTeBXNMjpHe5y8yUxYboiXRRmC1lniVDpJgqtyXAJLwzqeSfcXYwzDj1
nAc8s3k79boSX2iWydPQtkphQL/PcyEEuknHaJLRevSphqAoT89WbYe0zfNtnXuZ2vCWGxfqlJWp
qn8siM72GBZH2jKSgfbaVOG8mQIj1Xxf56f4WUmY0eJ7L0U9GM6HA0RdaV50umKvxNBFOhxstUCc
ZHi1dfRTHqeAGhhmxAvZGo7s2Wualkib4ebRLsNbS6OonNQAUidhTo3qyc8rCJqoj9ezNfTc2RDu
0/84PwkSKL49jO5y7tGnUP1+76yQPlzfSe5eLX90VUCdCQ2Aueae4+uR4P/5S1xIn14HQrU+Vx8T
fw3lBibT3Ae6geRzhTf5OwuSGqWhXkiNgWhNQH2s2MhFzac+GxcqjT0FIz426KviVdUqtfVPBiHj
yLVEtS2jfm353U4qciJA76bucEE/EqQekzViU5KD6aYsHnYF6gXh65maYA4kIPRDC6mwLflsZ90/
wxRn5hZbGJ2DSaw6+PZ92oZa4rO6VwhUsvYOUbP+TJRKsfguqsrS05b4+vjeyYwrCfqSPNM78VVL
8eH1xa0YC2mWbs1hvGqJDGpF76ANo969jfwSTG0uiQPQ2lPYo0G79Xfx4BpaT2xTEZZyd9bxdDL4
yC0717qW7/EETUETftMtgOSxLzr9rL37zZr/s6jHswIvD0Eta1ECqYJEoeYV6hxVWpeAjimg5Rvg
abo7ypmdfHhq8jZOXdtwkEhFf/KtZX8uIbtIcKKAQDhsHdQd0bpnBheW1EKOSUauxtqkR9Aa8FOD
dMvHaGptdXDxjPbWGumPQkyFf7NfV0uxM+tKhsB7ORGmrKAHsXlUAtzpKexXN9b401bRPR2osLfC
0IvuALlTbNWQks/qH7ndMjgOPTnro2zlwRgkGlDcvo9I3lWD3aU8cZeCElTbT0uJ07YD+ee5zX2H
iYE+4yVymgUTfPQDKfd/lA7gNmK5lnG1z1OtQy+IQYcoIHw/X/cIUsTVfR8hDJSfn5EdymM1NB2D
rQJEofV6Jd2UBRcAjCyzCvnNOVdn0T5dBS64/5pd1G/MAhvaJ3ceLxTdFpuA4ynO6EJaPcTIh5uz
aiWO9LKYvXIuft4ZJLaoljw64xG/OC4jrwStdRsuGlRiJk9w9vo4k38EHBoJDwDHo+ITtuM1Lh1b
fGS+S9IYixNmMNrwpoJijx0N8tgfHNqhtY22bcps/Mi+QUTrOL8o023xuKVCcht+DcpUAZS8ijTN
EeG6Jd+KmZHUIDe8k7dS1taC2xVpbqs450Oei0SnLEDNkDUA9BQfcNRPesF1muqUCbtb44SpC7QF
Z/s6FAqFTZ2SEoxC0oI3YTvxwnXoH7kMpk1T1x2GZ15bGvU/G7XaArMVTUYy9ByTU92982WJYSgE
zRuh5QKxQWaOWO8CfPtTIsp/XyOMfl7dUQNvb6t4RDVU7BhWEIi5SurfSm1gdpE/orrNiCOjYNCk
DEK1bZUXOzQJxXaLMPNUKrmBBf58q4lw0N7IeH073Q6jIVRwXAGxxnBSiRAK6TEeUbXyKGx2vB2h
cz73XR488T4P/g+t9g3rLTiNQBey7h/RCMLgGGzMRe3alqAKCx5EkvSyXWb3wzvceoW9lL0C6TjY
MSiUUjPU+0Y0CCu8eGLbmj+GjcCt9lwlRxlSrWC4uL+VyuQiMyngeL7YzseH6Ro9RBt9xKJIiFkZ
xdNFFAQf6N07ccH/YWibhWcR3pvgQ+O71dQzfF5LES+0+8nOowgsiztj2Vq8VCOM0p4+dVcc13nK
sxRsv03myebMk98c/XZZ58cCjfBBStjrS4rZM/OwJaxdmjnzCO5xO+XftoeqZ5HchwvjGchmXWFi
7qAsd9TUEs6QppjlU3KvcxbiMtEG28w+F7WTzOd6fMbSX1PRpHDU6Z+2bgbHon/hxcGtfz11Srv4
JvyJ9wGtLjz7GAv/1TebnC3D42NvZt1eT8EauhjQ1F1YKRJ0vKUN6AHKil9gwP7kK2eHiwnBGE7J
ou+LQnWJ0EA90bK5358fnFSDPmuNkAQuH8XHWOMY7qvMJg3YwI74cxVBdxu0J81CjCmyPCsJz+IZ
fanxc1GokWbpfOZDIMvtUq9YffHzwrFGO08uAuVdPArI6naN3tkdV/Yl5BYH3fkdh2f8M2kJZer5
+UAT7cfOLZfwIEmPuyid0bst60H6fcJpnkqvp4/uEddEStK+GHSRy34zlOvtPKbXipuDni3+3dnO
Aj9jZ5+w9Q4ojvFVTBNDreCOrcIBxwHKqOffwjdN/NuXgpAGyCq4s/TCGoneXpDtI0pQRThs4gLB
Ny6Bd0ABh3bEupN8jWcfdM5gZyVJLAH9AK5LDVdqxkWNdKwOi4OuFBjVr6StPc5dTbEIJzXk1NdR
BEsIgdpjlPsNtORO5Ubc8UgpV5ZAeFVT7fTQAyfydJRYTxlCYGcw2z2rgxUqI+fJBb6V938Xewrx
CSbyGzbASGl3D0vGyxdz4cHETQHdlZjzOljMqjLdim2yPNN3IpCje/H/hbjczrXNzrMjQC8uOKaY
b05ebvtriBKau5pY5tH1fHo0P4+KqAw0Cfi0HOyg3trq+/iD0mYVSPqn5vi9X/qWHPXgN/3olIL/
Na46i6+2o+x/Y+FwtoY1BtLp7VS4o/hUd/Sl8DJAy/8hcDvAMuWqUGxfRCvnMU00SIaH7bQib5lQ
Q2U9leGEsrlhm0z79YiHrrRhLelLQG4+4wQCyjjXQjuK+HCZd2eWj+/zkVSq5j94gEbxPbpd7vq+
38VYVr4SPJxdtsLdf43ayZWSRNdFOSLVcEAmvIEODdYom3BSgGEGB12Tl8wODWEmAH97/mRnqnHB
PziSpZfHhNTfGmlcAe4tV9WSi1irJc75Pemrx52yIE3mOqUOXn2Ee28ud2+7/jdhTew2IM1mvH7L
LMXLsZ5eHQ3rjouXKySGpcLARVfvz6xIX4/4jht7HwhSCNl4Nmjnk43wDmwFIu/4wGPqGmqGNgYp
PzPvsvNZ8V2YroctLegbcJGoyMllWuISrjy+UG06EuI9Ks/hXns6ZzF33QDJYAEiaCIYl4kyfKpQ
kZk9rMeflD0a7Yegtbj4Ej9zkpCIxXtJF/3Jhv7TglEunTd3eULy5fgwVMI3c+UCAPFMVe5xIl1K
9PdI8iZy4WrPzupe761lLcGUzfRfHvmXdl/1n9N/bhh/ErfZUJduBU5lKYUAoz0HK0pbbdeyeu8d
qUkmRTj3/g0JyNcPQWUIfg08wkbCLx3gV/CH6+McBmC0rbYwf8iz/vAsvacdCQSQ5jbZ+1wQ4MNY
tQoazdNdTH9ZV7U4CES1kDBZ7bpZDTZqdhWQ/fSpnHZXb9udLubBl9BEzHgKxWaKLQlaPZXpYDGj
JVmkcXVWU48eo5nBQVnOXIv/EaV7hGEW64pnaNF5UUwJF3TqP5my4X0ZfqcV3fqiF+ObHDpOPWS/
Z+Pi0hbZv567f2p3ihNUMbSpx99ZZ7AkteYMutErF3OvB8yNBq7usgqvFG5mkSgSB/X4RO41KmNG
PxQrnYjvbtTb5fZsoQi32IPGL9oUoilxelghYylTV2jfVIfMkQVyDvOmwRUbrQ7rHBTDhPeLcjKp
wsXXoEp82trLWJW9KMQv1tTUlkUXMm7w9W/Q6RulXQKs2lct1bqfoa1zVppDdnlYoSjmMZpRMWFv
dctRlrGd6yeY2/XxTi68JYP+3l6+6crYWOo1FyOHHfhdBgssFG11CUjcrRv3msjP1q/66uI+AuRF
AfMpSOA9bA+a21ryVQKfmvBu2iS1Vn509dz3ztXbDwmQo++ZIyV+69BLJ9zhy8dbpzzRY1NKvZ7k
/QEivG5bW82At5WJLjNLgQAu7uGfwHnoR9PpktThjWSN/SAWkXpuGNnRZLGuHg0t5qG6pvV5+KoL
Z6QXSRYS6qN45UUFtz9mMbnSqwhLHyVo05v7DzzRgm0GllyYEOO/6qYe5hL9ru8hAGEa11jYVnEl
LY4qqSEdhhfcZsUM8OVZRnL3U7mhAqLgU+p4ggnQoJSkZVXjl/ABOZoTLlA/c6iGg5gYrQXgOFqY
n5uVFETtZUcmubpTHFW+CvmEx/ZyYrSY4F8xf7KetXFWbyzNBx4Z6y/2+Dw+uCHhcRqxa/2BX3B9
tKdLfYPwJdtsEkw/VVuNcV4ze3CP/Emj2qWGTyIrqRsaf3SF1ih2Rt+WkxQUEDI9KG/r3lBkU/g8
GuyGx32z2PxIYB7zNdrksnl9DIXXhHrAKpgDaWleu4wQ6oaEeK1hpQd/esQi9IuEJt8HPmrD0drA
8AkHLxqdwIEEV6mkIjLJILzbgo6CR5sxzM9FfXBXP8vnk9BJVxoM+tnvzZ/lyDxKwQx5XpZxzira
cYxWTdlyJBZL5OwGS6sZknXj+kZ166O6RraDmTsT6l7EEYhwKpfPDUEL5+MZwaS+OspACP1U+gya
YU//WMsFKls2JL03EHRXoZtnaDVhBBV+eA4XxaZAnEtqAB6dUoHIm5mJ1fClxFSzdvgyF722qd2x
9VAKWwohmcek4drgeoXXyZcmCJGWGB2JajoEPQLAbZ/WJpkeJsjitFXI/kI3JNXJRI32es3aE3Gk
tyXrv1TKkC+hbf8e+Hp56KKiWLMcFXUwMoxQWJWIxXqEf4lwPMMg1sp0nV38mqf/WMsU6PKnBRq/
+NTwGt8RVi4qAj380q7l8XvPXAxvnVN8utwyOR76d9FysINORMYDRvv3DfhzxB9EKykDW83FcaT2
0/9MtO01EgJMtPna7p7tSwr13EV2PCrv+feADXV+TGbtRgoa6xBmTdCEpe5A3WiYBB28G00AoKSj
oDlarXencZu8ZEIF2ItwhzIGOyCuJ2VlsTZErKYrR9mZzh41YD8cWQBhwI7XC+lSYg2sYarQolIV
k4w9CFd4meQjhai9UEgavqEv148KsYMrTIaApllDy4PMqjvMpX5W+tetFV23AhQb8WOf2OVXv83J
xyFAaC0ZD5WexJ5l5OPYnTn6Ws1GwsajVaNWxDqlEwO1HR2oHRD852ioqoLKiMo9KFjiE5+nqVnW
NgQT6F588TXu9Ss/jHR75Q3avdJ/Lr/DpEy+tu1X7aFiovDEqDqRGuIUJi9O695XvbSVhSBdOWkV
94o6dhzM8OM9C49cCs9Fen1re0etC5JmMJfkJRqPgeuvL4TTGGlDEL0SDlUWuBwLeaUy2QMBENIU
mQsZQuT6uRPjZFBC3r/85zk6q5IWHosMpgXD39R3KPHBuYfyuHrd+7B9IUF+JOINg3GwRfsM55Fg
SGPcf8mNz667h3UKb3vYUJt20u1Ka6CfZqOLHCUhwgec6xmkdkPwKvniDFpCINVpw41L0tUS9JPy
5SZ2BfPN0R56j/aNRw/N43QpxNvQORnfGkaC42jZ9cBrV0fqjRseVfviP37x6kG2930hVb28SbAs
xFMDTa77lsqHzlyxT1JfjGIZYOiZxT1yp2zFSCl5RZTscctaN1nlPdXyTfIApHi8HbhNNxy/3nQR
zFZmogYrmGk8qBEvirzoxnJ0z9olpHx6WNlaAv+1BzsCuL8R3Z0YPcIYOFMyZlGyvubesK+q6Xe5
r0w3R8lvAw0F3JOqE7RvqQiPcAiJf9qWiH1N4GUNqh+pHzlheT6+ggVk6E21xOqdoz6K+RCciEoW
GVxMhkdUtMzVpWatQp2yqUTU3F+Qf6OYo3oYfw9wJKofAvRcpT2BSyDWThXRqPmIxiRIbeaqTdB4
zTcbktuMKU4D7hNmbMGXL1QW74pSfrX0wkwWTCpu26c0l7rZBz1Z1ZQBkuoq0N1OmflN6rniv0IE
kD1d65YYrJcV/fiVRG5fvmRO3R2pwNG/+3tNjccu+hUKSVm7hd6IjgrEBt3C2o9YJHaayJdEdMFf
2ym1Sfs9kudqQn7XhdApkHSvmH59ZSm+EZUTIaS7Y/Jqny4sFckjk6ZWdA/Qonu7yib2EXJMdnmD
xGy0Srulv/XYGVtw7xKTNySqOjrDNP4dPmNwSrV5IjirDz4KCFiQEj66KbQ2hICetUR+f64U6uIG
ArC0do3oif2+yjDl3KUdfJQydL8YeEmXOD52bDSrHRlshaRNez9WfdWSAH2MhnjaPMEDLRACAEHh
/CnrksMdC6BBjrO3TBZHg1MUjcOimiAO/IUsWzWVMu6BxHn77i+JuKnnK5vG0iNvYAqj3sGMo/Kj
ZXoGcLhfzQvBqJ9bx8OZiJpKUH8KvgI3vRN8QEyuOvDZ0YN63wJb0gdToXKxF59vyE2jZWAjJEdO
hCHfibOZ6wSSAHjbgCpCnPTys1/2ZwcTGeP5DUfbziD3+iQfY9UbehDybcQbD9TDUwhJAVqvECrK
pxUguW9gLWS/6Z1lY6+AETyxaRvkCn7ZtsT9jOrMbTHseOf4H6YhpYhc2/s4VzSMMcu8U54qtunC
geE1xfbijNImtesNQ7h6pCirl49ymuDwhJzd5gUGtmSPxskNybE6j5WT1W3QTXPLwSdGceSUKrU7
6dtYfdDSppnTjLotUJ2hCDpwDCB09eCIlcvejzp3pa18EyLRjJNRfaMcHyUdXzK1Syq8GpL2aHKL
/79q7RhpLYKC3x9eYi7/g2zo/lULAVI5oB53kJtKLuf16cucP2umxsV93rtQrfG+YaoKCkLKapA8
O8siTiVHboOlcVSLdaCR98JzgxErlt1/ti0bp62YTXh6iZ16QUWH2+sTJZWQBdv9x8wamqbC0t7p
+bY28qJyiBLZlnKeZMT2qhrpavVmp6/NL/ltcQzbCnBq3MOPhxsr6/1sCX1qtmAhEAF8PnKlyyOt
l5SZa8+uLTuQ6xnmuIuP31GtKuKrA1xssnGvKR8XnL/wg/w1Jef/Sgal1IrlpWvne/b4E+OoOvT1
J9UKvlDPBEJPM13rFJ0HfHH+I5tOgntMK+J/J4/1z5usFFlPLHpeYFAtyC8u0A9wQ5jRCNaOXFy6
U0OVjNpuPzsups0cxGCnk6twfBfEX1immLkUj9gGeeW1JcXt2W6UTjCsa6rjS+1K2p4F04UPWLyq
LF4QT2rQezokTqTJ2SYzvEZWvB3FcEJh0425lBefwtlCtFFDWcb5yjx4cxcj8ccdnLD+vYvAhD7/
IY/8htveqezLm1M1ABu1kmZEQWBJAfOO18oYD1FkA99TmfR4YO4vCpuyWXoev2/i6j9WS+LhO2Yg
HC91k6PCGRrHpxc/0ZJ7Qx2TiHfG8fr1xtHPh7tAn84HpE1oSnIlK1M88EHr4Krd7fD9mbHktc42
rm7S8ZnVCQR4S2gJhOJdXr3jduI6MSTAFr2Rw3se+TrdVG/UoT7rZU2fqh/9wS2lxYGp5iihel03
Tk/ZLPjkKY7aUzEQ9XzirCpkzB9+bUzIXc3pISwv7s0W1iUUrty0l2pZ4vYXmG1NiAVcypcYvguM
hW22F/9RKUAg7fKeUzY2WMx3lO4/RYfEpAhqAYH7vVKeWI0Ptz3KQJ68Y9JBgeYn0G3Zjqpm3rx3
zgmof0xG1Xvc/Cqx50ekowXZ3mumejM3VXPLp/BazMtPKa2NRCzM3EI8EXy8YjyFhrGVx6i8x3EV
aUN0XxL5QrYX/Mat+ugEnFOtK0wiFAOChvB56TWHAf16gv+ykMRIVReHJ24o0zTrI71VgNIl8enM
TPdg5V6Y8GuVu921MeWcIhhn0s+yuHVviwaPYAJQjoiHBlhKTdIRNdE7RRPvcLN4d5qf7BxHEiLp
Y5HQ2kBuQk83LYEQzLkr9uJugQdFbqznxwhtnU5DwbRIZmsKmI8hewsQAbjWwoEsfSdb4anR6P2b
bagJpc0fR/gBU1KmHCTy33rbi+Q+9cwF5CUewvjVuavK+vkvyAcDgDaiuNffB4eS4l/SgT1K7rqR
hvkEe/NKnvNgsQ6wrFSE5V1n2er0GyIlyut+TSK1BrFfjMjtk4Ec2Co3fuKrf9qxqPgg9c444Jxz
X7vvPgQ4jJVd3YWvsOerbS6xPzGYrlhvfAoLg7ixbDhBdwIL7rS5tXhZ9z4C27mATOOXfyibXV1x
FCsZeCb2dv89+cgAhBtv18EXoB0sgDHzdRra9Q4VZwv6lvxzwwNyemAqvdxClXLWeqbCoMDu5NcJ
LQYjJEp0YRcqTlGGCSM0AZq9IIAVZ6QiraZYJF5HaAqizcxoUNLS54eIr4XZskTFxozU8QzMBKnR
yqGa69FUZoY/CCCKiL/xWWz7WsP2G0ZviaBABmEGjCx23CRPWefPyNJcVL/kJwZFw5zMIAxPK+i0
077lqg8knjKFlsRLJhnMqVkFsSDzpjECQixcDmyXvLPStPqn/OaFfspZ8+Gg4maKCk5ZDiIpl0Lp
w2RDi8O73tPDVk6S7T0QZVKlmOUxzEU7uwBA+Nb61PVznpTjUDZKdAbZTlzFATPSMl5WptrJDIgK
a0249zTonQudgBhZ1tbepgRC2RexBIIhwCHmApb7dAZMls+6nbZ9G5KZeqYf5/f21FgRPQfUIzfG
Nxz6ZroTHCsRzb3URpZBjcXAR2qcflqPAh81LWnv8UByo6NwRu8hoymeIbJgShhRv+5V5zUeTHj2
B6J4j+Y1Bo5RagKbJVNacdVzpQHFP8WwNVQ5t7VOlP2t1ZLF6mWShSDJ7Jq6lAIDyMKY3JKAYSzn
QMX6a3m+YOl1dJiNKGbh0/yLxu0vQh0ywKvg4qm66ZAIqmrKwk7UocrjrUn2mgb8jnbZM4W7ISRv
bFQrPeFa1552h0MbwArB/PNQidGalX+MaWDxGE1vVzLSNEyAA7f4mugWpb0iigVyrfbRLhQb04FX
j/Yf9lmzYUnqmNHBbHW0sNwMkZqOVISBiG6QPBCEsGp8iQUZT/j02t/xETldaAE9hsb+we4Al2cA
qSe77O6hSPjLFkuRrrxi6lUBu/8WDPptG9Ny9b6APcIoWfGuHIsgQ9eBH+YRjmqg71V6h47lEQSG
KfFqRP5fjsEBinu0LE3R2GhadfgMaBqmy2wpsqjF+UQIjXeouYVqBW2p/LhkkP7I30sN9kDbhaY8
/av7Z8hePKU7lPANA/N3Q3iMHW06NmA8lD5k3ZXgkqTcTe3jKrcdJl2H43jyuByGgkcMC39bAeSo
c0o26ylq3sl3ihdBt6ANn0ZgSZ3504riLrlZn7bZNj6bCIYM5NOZ5AFRW8E7uf/MCtCKY6Y3IIOP
qR3dbwFFpnm0DEbQNoE6z1h2JC1bUeCAmooq5QpVwpCHRhLTMxhfab3A0JanBOBCRISnsrveADul
857E81v8QWsGakOc/obZu/lZ9MU50AvLVcILgw7ad53kqGX2Yjh6JCVr+X8TPyE6MgQSl+ZIkPF1
fP5SZNef5AHM4Np1Qsq63k+A71RqFVJfHjVwl9niWDdjauK/sxZxyqtYWM6m36zwdy+2C5ufkbA2
8RQ58SjeJLG07V8Mg9LZBIp0ySV9BnKm11Ce6HmesDRijYy7T5T8ryiCavQRgFeKLSOq0yMKBlpY
MvB5hH7miDOj1GVr5jbIa18TsGzu43tvtFnswPJNj5ULsE3oHwlt+G8wEjAJgAgarakYas6cxwR6
iQtbcXgwUkgxY3eXcMa//rYue1vurUqfNocJXYobqViuxZYgJCkiMqbnBx3bbuifjcelGJEA9CxA
6Qj/+hCvoGTQRXHXCmtHy1WquKyG58uBqTONYd70l5dzl7zbq44r4N+n0EHIuAXzfhwu1bJ7Wac2
4eVEvKl+6ewms4h75hks66ipXAExFg0S5cX99XcQKtbkjNCB0t5Qnp2Qml0iMBbSBSfcuK+KtfE7
pXKNrmAs3Ii2ZwFMGysRDm0gF0+VD3CBstlcWthvF8l4+jrw7thO2ewn3u1BB4SBoDKRmcmQtXs5
WO3vKepY41htJnhrscHA4jn78q2P+EO6y6mF6+n0NSeAPH1qv/OZKFfUexulLsvBhBg1N8NvhXd8
bYGOlMNJJwNV+yoc7FSxQj46qfhA8S4jPYXU3Le9kA+XiCgV1YCC0xSjlKxBilHwlTMhaHfWkYiR
Cdckbl3iAla3dATAPmEpfqgc1MdMV/G5/pCEEDg2oAHR9UgaIeJaAL3ms63H+KACJ32IKyYhaX3n
VNkiISFWRHXmCiji58yoYKcJstgqoOltDygQw6U5cVj10QnrmEKwdEnPlGUIyMHEOIugv7Uyd0pu
ChMiDWdFXwpvEQ+XcaDg6djtY1q+vSqH+dEr9RQhEBGp5+kSqOGNp/1GcW8MlfDqP32acnLbG1A8
eSVNQ/Bf10XfI631I1a/Gok3IobvFVI5eDYoa5fzZ7kSApvf7vU61LA/t47EvrSEre7Gi2PGwvFI
0sFEtHmrypCcC3zlSuEYmwCSB/1zqv5WVSZQFVIfGbFudsaQy8Pv29lb75TZTaHUu1xDTha/lP7a
VK2SDbUUYm2zcYbM3jjnyqbw7ZsF1d4B076p9HRc/AE9uJ/pNtTmuqqAmIvlsTSsU3PsflmcD/FY
pdhNGEkFKnP9DxsZWDuMyO00y3/lIzgmQJKmOQESeMZQaFGL7m6B6WWu6db76uXlmb4G1qg1va1q
AUlSSvjwkPLkodDRISoj6L2ABAv+qZ25Gz6GXQg1ZFMC0mMux5ZinrN+2EEsLP3bjX7SC1gxSsIO
XmiGFNJ43VkkFk6NeEW6dnITPq2dax0xiHXcE5754533JM1Irvf86fMjvNR3hTpqLxcj3SI379aD
vqImvOz0ZwYNwBZLxOdEcqf8BXjQrXfAMnKC6N6Z3iqNidMzubx7p462r6fFUmzD5331dNrdZx1N
qLfTj6wyrRNWG9FSU5bHT3z0QFUe8IiEBwNrdICr41+lxExsQtXrseHoaW5UyFXvy55hlHziBaTx
8Ume4QF1KbqixNfXvqVhImBC7QX/v48bTCUpfxfrBDmljnAzwGFIu4KQ+Gxr7jhF9tCSSNptog2U
5U85sXf14oWf1wQPDgVNK40FdQpHjBlSPzW+NzyZGoJO3I7nd0rWX9EayWqcpVQ3gy587o8+b3p3
EAQ4DxGUk+pJEBoX0AXvlwvAOdtXmUvIg7iVsZyYjRJ2aMevz+Xz15nFT3/LISSluRhEznWl4Cum
AocFGiXGSuLzKQY8F2kHCL9vAgI8kkzUT0bZb7ErBkr/8V+EWEH27URfG0MxrEyPSQKG01E8XqKT
udP/IWCfneFyK3Wn+NgrWqL/A2WgulyBKNEISjB3qbois6XwLvz806tAeNheaBHFqV4j+n2RTFmW
A9caLG2q0VDxiGXp4hHlaA3V7bllxiyYtaON9R1DjqjTicN6WAwZJ6h3xC3q+LcNPcgckc0u/v+D
6nQqqi8JGRmPYvGJs52Jt1sfQTw9vOxfJuf2UnRCgbFBWcTyUpA4eKvrTADoXTthzX5YUArZVBkM
NN40pvCSiugmt+5b2lMmFG6zDKNmL1uMMsuua8wGp/KIIuvadllSUM+rzyKXM9lliB+I8Ffpokpk
sn+zcgX+SrMsepqymLLDeC+wyrD1VYTSahtu0jAAgKcdIx0FA30JBOZrAe6WJgnWpLNcUHa9QTRg
8VTABzJIWIg9kc1a1l8gTa/WA+rFWY9bCHFv0qKdaIgfFO5DR2Qq7Gn3TAycQBq4InVROaXZYz8n
cWdorAgcI/k5LuazZozq242JGERI+MmeBBeBDNHMJiuIvSt1hND48BArN+JY546ynwYvjDA8nTVs
h6z5T1Tdpq3LOg5BYDcIguj/ylJ/QzOLaO2VlQRJC65QI9XhtWkuQUrtIG9qTMJCu1FJrRZIfnLw
317uY/J5qJ4TuuyPdHucFG3Iv1gX4z4i7+ldaxIC0sy6KihO+pXg09dMKZnR/F6ScpbINH1ZwBwZ
8mh+a2r0guGNGTd1o88dybJ4SOdjwqIahHkoSgJesprRll0ssaVq074+xT6l7RUpRXHR58B8I7QS
0GtS1DUD97NdQgf2eVtKluLMcwnhy/bgx0dehEsbxera/1w58KEbD4ofZN73ywBvE9bWGVvDbQ6N
p0dw2vpgLzFfWVbNm7uX8qzWCrUEQDJueSYLkzRFk++YzoGhqPlUPacvk0UBvMRFZmaDpOoBUYDN
djvOeuRYg77w/swX+Yoe8ooEuvikUVsT4Vk+UXm+UeNeSCslwVFM+QiaZe9o6KNmwSTciZ8/olCS
l/ig6JA8Ib7YB4Hf0p9NOtaJm6OtCpMiTCP3cCHrbUxlh5OnxJgecajERqrcsgOQQHsuKrQWh5RG
kqO6I2smh/luY61+Q+yX5g4TR2ZPIpWhoxNSs1ZQTkGEfsT6RnClpflsZ6pMsgZA4BOJRdoagSzX
EImyH5cPU0mOE+57MwVO0nbB5IyR6lrZJZ6INabzpUbYQ6gq9fHP83IPgyexQ9K8z1/Nw5xla2sZ
LJjFA4w9NZdrJ129Ur7vTQmGwWFlKu1XmTo/VQUkuEUjcIPbQGHLJWKKrhkslXAgkKlvJO/MMjEH
I8vo2k0mpZC6zuoI0ycMvMo3joTXBD/39zt5wk5E06cfpDZqG9Qg7r1G+Pd2j1TznqkSAcky4iX1
VDMnrjZgY8o+4sI/1ahDMfs0rdAFnArOfokwIPYHj2zeBLXJslknlfMRqAav1OSX/AIAyI1ABpnM
1peBIxBEnKZdhKTDPxXqWXpPIMVkzIN86fOqLCGO5jJ8Ilm8sAO7KldP6kwtGN9YzEvpMu07HR40
xtI9CQYDqKT6uQYGbDlrvinqHwot4jWEFHOFJMw9rbBJQndm8GyxyBI5VJBV7F1fdeB+q/qn6efb
luv/EI+w/u5U73j9++RRZkZqVOjnZsJ8RhVRZbm13oEuNdE2kik3qtQw1Bp1w+JQoirvB8q170tM
oO/7cLwWl+gXfO5R0WtZkOmfNfXhQ7bbbMyiutY3pYp7XhhwrRLgc3Z/sMMBIcRY5BGzqCDrbcLw
sxfqGV0XFulo23gcKlK3X+xREFAPTGq+qV0qIAWX4o0d9XvUHmXcJpzrbXPU5ywqCsITfK4JSn1c
VRJEUF+quYLi/kxOKKWFR5FitQoLTIDnFVhyB5+JYCaCO3NlliufeOCded+Tp9iog0ZFyv/+OScV
KYqFQXiRmv218Z9WNs60b1oeOlHhHhgFeN+GZY1RljjMqDjcOM0ZufYBjXQuVgxfmlGKdJDLKCJk
8EkvnUOJJSr+O5gcJf/W/LEgnhs1NbESQhZHWKJPmcUsQy1zJy1aExEA6ELYJ+n0JMhfuMCpw82q
7pxsMGt7iDMM4ViGc5d6OedlqAa3E7IZGEsOGUISCyFmi49Fzjl7p6iwfwiBuAu4/ZhfgfHHkl34
GHKEtkcZo1J1gskqHuk4vAkMhQRLE+ZWo8/QSH8fdVDuH7aLvOgFT1WTzTWRTd4Fep/wFchjTGSI
50JFCBqZu7D2d80AZcn+Y4Ge4uMEQ/OZ+CPXetWpieVFiqgt89XfILXzmVTTMXNj/7BnLcsUYB9w
zHU9eWeuGH8jHXsER69ycwornYrXcSvi/+IOuEgYgYGxaBvnGUgPnHL1rEZFi/Y6+j3aavcCoju+
XWlMu89kkS4OgYATEAG8UIUv+9ohv2aorjv+LIPfNdZZy18Lly5XdHmh75LVGlImgyQtPcl0n6bk
ozBcK45LNpve5bomBmCFyMSuCTXuyjXEq0tqakzi9ka2aTaZjDrH5r3l+1LQkaFpbxQPTIO0vcvD
JN0A6YZ7Rc+aVb4kym6GGLsBJJd9eP52slEH28U50nCIXCbuMi7WgmKTZkEL+AjuLSr/oveW+AW7
34XupzuxC6fXbQNhGztfAn5sfpbIAwM0ncvbitiOvwl3GMKMF/2vp9ObUNXKPe7fzctRH9vRk3MZ
7+2Yiyik7kVz/mUxf+z8Y2PparRFquJ2LFYzKO3PC2E6glnIYemvukMqktK30kTTuchjKAQkcwqg
HrQjk0DPTTcCKAoYD7WpCTAqgHFuIH99IGL3v5oagqVAsry4Nm6CBwkgV//juXl7EpSJz34Djxw1
NeWUzXdQv9IryJRDVQS/Dq4DoH81T/eOOxJXKrLla9P5pJ532GNSJ9/Y48p+A7G3XpvoFzTLqDWH
1i4pACrnmeuq3nphmE/o0Pp+gUclWXWpQa2xo5jhaAtH3j+auOf4xd66dScTuvAmb6E8CRlTeujU
X/fOZFzTZnSpVcT3welsXAs/v53MAh4p99eyjE6HntsgAgC5NXX1Wd6gIO0pYKME9NZcxtyeZwbK
tTdw0tGq7PpoDUG65zi8EsqswrzHOojYytPWgZoq8ANvZj3mc3FGL2THg1UW2OronlPAO9SGpl7e
wwg/sk5B8G/Tl7UHK2UZFrq0CmSt5/Wzr1yJQ1yayhbzgQRfP+7LYgFVhD/JpRglSWnPtcFqZB2B
qsgBpl+GvrJKOYp/eR0cyWfRAdBHxjiGsJcwiBGmTfb2DxWkj7Menw1cNyc3fqP3P1WoFX4Ncfw/
3heVDNlIFkWtnZ1wb9CguDbBr4Z8MRwqBBqch3c5biHeDTILGd6kccaUeuRet7Wn9t4cvAWIJOdT
0xXdHCBfOlj4m8hpZO+hX0G0ttlGp+ic/DqrIZCMdR6N3vRW2xtAkk+dEszLSS7DNgMQ76p2tQna
qj3OL/uUBHqG2stvCtultTch6JQHQVSudyD35FImW2OgwmGccSqdTTnx+rb0ZW6u97CO3KgwCwoP
FUyuYKpR0C6w94xHJonOy3SC/HTLqoJPvZySaJtss4iwGR2UUbCUdE0vxitVxSQuloMxRP/2yQN2
m8ZIuSEBWmyaq0gxIgD4E8DvMeyg1qRyOfbnnvuEpKi5K1U8s6QLyoy/fGg86j8eWda6el1Vfb3t
h8S4t08RM9NL0vjbvMpLtC0DMX8H3BOQD1pOPINh6T0C9wuZ+KAFRuse9Q35RkQhFzCflfYaP8At
1ErZbaGnvxnW1bcvsiWc+o3w0W2p45balrwb684XqemJBVqMUFg8AIiUK2EC2m/OUsXaCh+KKZ2Q
S2rJH3vWWd1BqvuKaXjzKax9TwVtcapMRSHq1Q1VK9RWiSoz6q3bq4Rd0829cF5R22Ge7oO2Hona
vMQp5UjH/ULVxlKgNaS8O5U9G9dc+9zrNZ5iPaDRUv1xUIlCcFl6uXiWyZEgpmThnENM34mFlMzo
f7hDrUSyfrjLjqw9kjRYuUKuI0D3/dX/dPaMuhzUmvsjhBSxtkrZgvzKvdDkYCTKKZtIDTt8EPtP
8axAuJD42XrZTzduR9ZYiOXQwPhH4DZ5PpxfhqFjhhUf0YTu4eR75avii9NW8xNkSQ6va5ebPmLr
VAodB4OSf/gjI0J7kBMA9QtA67z14tAZFdjVU2VgKb9HL3RhBfA31zabZREe0iCMzAkGGA6kqmMF
v54bmbKkqkIPwA7o1Z/6eAYkI68jUEuPRoMR9wi66mT8QzzZaqtUGiMhF3NkrGO1mcIJwCu3i2HJ
hluBfwkgid+lwJA0loOriX/Ts2Y19E++rCNEzkjpPZzNyh7Zhak19EgIIS2OEV5dQFNUmm6XjArg
488czpzM69ZUgeBJgjadUz9bnO2kiDl40hsW4JWrlIBAgcIEoC59opJpfBNIgHnP4y23ofXKO+kq
MQvvTjdQJ058LNu25IqhuMNPE+JZpNguq6XW8MCm9d5a1IfQDVGOzKPRM8pw6nGtd8tDP3hsZhfB
UXiUE9Yq2TaOmEW6GfPGIfKZi0bqD9sdhz3zH2wdbSmhMWrdxO/TnNZaC7pGWZdNFrMk/NCDBXuT
zJ/dzyPV+VGS4ouj9FWFA6WQDFvTP9c8qIdlIWa85kzwRo0QP6GoMLiNpIPD7gGXD0YVloekoRG2
ybJjQa8/PC5MLTLfCuLP5XwStKBj6fkaqzbwfPVMae7ZPK8pTyXsOed9Pu0+QNyswnc2updh0PNj
4QZW7OEO47CqLfXBtRUrJtGqOm1flb32hdAlstDHhD+c660gvr+JsRaDksZB/7XrE/fHUcBuNcqb
pNFO7Oz6ktz3zsqeHImIuDWRoEK4hRVj6Q1ycsfTrHjNTJ50FxUGb+SJo7TdCGgaesoTaRZlqVRA
rz63gAinLTN+9rqtwWYPDOM+ijmBi7OGgc0+VI7BEggLVUNSl5T899qijuTjqC1MBuGxnIcO1PWc
mDSlTui9S3KmVvak+It+6LzAlMklC+KTJnl/mw6V93zcS0luOuzxFps6VPJANfdLL9UG4fRKErHv
s9hE1j8aO1o6av6RpNzq0mF9l/Vs1JyUJkBGovmTSpRQzGXZFs4Mws0AMmzsF6JBtoEpbgq9+e73
Yie4AdJq2L7pA24WABhtl/d5N0aCwVmMok3S6AG9mEDdNQ2qabgTlYH+Zlo2UVmRRu7ryelTZZjR
q35NsXoSGLQzOKTsoMnICCcCPJ+LfBOHWbMcyNUjRNI3w3uKLEVYyv8MWLH7VyCEbLzfLmDAWu3R
lt14CichWlRsN2aBCEIYTC4tkHyc00ybuCEnZJ6ezIYEYBt8atqDuaXpNfFrg226vPOgvQBwjU/7
dUhN698CahCfieJwdi5/Af3dCaxxrs1XJd+9EoLe38DznSFo3aDg1BPUdd7IBOu2Dxo0L6KTP0L8
aZ5ttnHI+lSz3ec9Hh+lIwqpDlsGe+L2ib5YPwWhgIRpMLp3k1XAtd8Sa5H+bYXWcPSPkgwfwRFW
s7oUegL1ojz58ne8650sq3B29l/htyGxlsFrSeOOsq7huNK6dN6vp72oSFbR3cNVDigbQtV/u2DH
B4MkVhe8HgoE0A1P9XbLi+yvg/4STY3lLb6hKz/FC9I1v+DAtl+5FyWziOG4r8guVj42qEG9RIF0
ZhQl5c+8CJTgj4cT8IWn4Uwyq4tyUQNbuhbybOl24GOBLz4NBnsNkZnJxohwsg7U6pdao2qj3DY6
gSnAnzawHc9TIiG6Ui4I+5PEHs8TVz2H1DkZowUnwostrO+TN9tYaXeeiVBRhPFAtN/OfjHmUx9y
8apw7qsJXTgZYXSTFOP9PrBk7CTFw1ngjeV18p0R926cqaLCizpE4yiCuLw9DS1eczI/mrEllaFJ
zt1DPmiVSxNf2wASVq2Ign1r7xAGZCzNil3k/43uHwCBd8hoeubvSypS6T5oS45k8OH0W2ecaLoD
0CFxNx33AhOJfJOs4qGHJKxofd5vmo31xNuwXw+dJ/BaWVs8RlLtUXBBNWJbwOxetSOu2kNT0+X0
sQoMsocykMIcPVnEipoqo2PdpXxc/7efUBNT19pvrQf5UPIJFGuEOECALMbx6M0CJL6uWkvbvbmZ
DwZBI5TsrQokAaD+TVF7aurnb22Hd3xnoJkSkzJp/vhO2AvoUroqOeBxCb+Seaerfpzh0CD7aOQY
T6KvYNGIjLnU8XsoFaIrQEMCxyh2qMAFA14hSrAaIdh77XxKBN8HDeXdOOFH/WDVYwfAzs/BHohY
sIR7tRi6aUiiI8PUYo+ByByAc6MPgftqoTcsJRmE5hu3TsKacXZXpFsJ4oTkZQP3u3gLfZgH4bM/
AzbG4JPRWfeuLX4Ey1kvZnaPzJhQPbGQt4c4oMwaZu/Rnmt1Zsd4gp5bJvG+1IwE/EBlg3aCpS9B
aRGUEwlNKGHOCIEE/W2mITOv/zhsirs1mNcL1lcPZUYJTX5i9wTzGpjl7fPfO0mi1/rp6ebEqnSO
fHDE5QFNVwbr8IKV/2qAZd4wfboCkW1XEVBYxu5E+Opu/9eVklXOIKsDqmLY/L33YTvAlW+101Bl
A+UkodtqVpMVQUnAHdltC3K6myFI75I1BKliy3SU4CrwN/LIUSYf967zGWdYBtBIkcgFCeBl2I8t
ukKVSudVficY6ustyDrRsu/avOIST4sJ0c7oKygeDwLPEodeH+pyCW1RW1WhJ4AsDmjPZjnmwiTA
7O4ZhJJwKz42bNbV2XlaXYH0jvMg7osr6rhiidM0LLM0QXNKSrwWXTOR3NcpE7Mf2VGtpnJDysLd
oU+kLH/3LdnJKTkOSjpY3I59dr12WlGbI+wAfML5xABGDe/CB8FAzhcDmGhthhn3oSUmVG/fDisk
0kc6jBwWaUErCbyqiSv7Y6sEa+Qsq4p7gMKomiLGPW0OEy+WmNctVH77cZfE4g1C7Txvuf/Xy7Ox
szcnwBVlHm5vlbRt/AYX//nl3vZ8A3CLlkVPUH0CAA1utGRG9tYWpP/ZOdijOUVBmN3x4GflsrjH
GzPRC6bwxW6ZDjoEaaJg312VSbsEfGyCfQlfyQf358Dr163+DOdSvNsPBu3hShkjJiH2BhaQA3n6
ffuGNg2s/qYYHjqf8+aANf8O9rkrRbcJI1g52a27fMk3/EnMLq/iF+2MiiESEFRWzUa9hPcnwq9b
lHmDv1dtYqxJOdkZMhSwAY0xrZ8x5RMczdgxsrLJ1jOxei5skWptrhJIgvrUBj7FQdfFJsRtQlVj
q9loyfGsG7LlJhfc3+WeM/MF84oJL7QrZy8awQzetkDzGSngK2Z57XOgnI3uDteuNHwp+5g+8HCx
QNMmPaDnsV0T6TF/f/S+PuZizj3f9GY9I7f22GO9mIiwEfS5Bg02yxlIgYlgKgdlzZDYAXlbJfQ7
2/qb3E2S2Lc2I2nY+tJcCH8ydx89cnjOsw8ZxJEO/LREsYiXqOfRZIJTmtDXHyXpQeA+BDLxYjI4
FEdROXhS55FeEv3XwNYLdfYEBRJk5pgH4ZyWLRzCLCRLEsZq3xgDxbkNzrUtNT4QGSsZuhugMR8R
jnr2CLfb+2iDb3mH/kFhqq19ADXrcRAI1b3moeH9rv9ll8IhCnh94qXyFxmg1xKr8QgbRVfLZ132
9N1E7CScJ1Cyzic9OwTJRLEvyMDq3YfFfR/q76XgLUhU7ZwRD+Z1FEHrUoOigsJ1hZz8+mTrNkZV
46pPn3sj4yOEMjyVOWXGu2pmWWMBIgo0TOt/8zwSr74LLxzUMwW515a79/bVwEQehAAAnsSmYRAx
61AFNgWdPXLuMrOAFgs/RzEIBMJFi4oJtA6jb6xayaq9Lc5rwaALQZ+Xlh/VsOISVhJJ7JkqWZBU
PEBzxkEo/087UdeV05TMSKOGEZC5Fm91XT+t5vSLvNtvLGMFZXDvepi7p/VfQg+52xmb3XLCohUk
VMoTN1YEOZGMvTDW27wTdU57adIgMfHniGG7hP9bWfj2TgWBqABUkGEmQXxC2KTnfmaZ+8BDjmjq
M6X0I7VJ4JxIZuHKLfctLsP/hzWLErWSoTPMErjVPpI3E49nAFXgoGUfotTVDelRO9jIHkDsQR+B
MpzctTUasUHw+1QcEFOVcFhT6XidvNrSYBRvzKa5vqoWpYc96wv9VCzVQGEceKSTmVHKeHyXKHbN
dd1/JUoyfThztNvX9NteR0xFn+pwqCq8EaXqnuvYOhDknln6AD+0IpwySq8l5HCSTOoWRJTxbgEF
aERwOmCiGPt9CZlP8KEHnnF+XlKrsRwbfA9c7HEaKS8sYRqpkZw2PyLIZooHCa62myaoZBbl6iqm
X+jWvbKtbhe+asVdtD7aTYN24QUGfLCx5O0C0EdtG3qWLBocKjCG5dytzkLnNABS6Gm0Qmt+eEQA
lTyuvaryusQT4SB4uFjU6Hhrj27hBRzNa3ZhExfCZKak6Uv5CDJdI4xDh0K6hxMK+ITs93AV0JXq
vrXSeoJ/ugQxsN6vJk/Cj9WiXOjrvoz0lPRT7ptkDDCABwzVPUdEWh/fYKlEA12gj3PU8bRI87j2
RPWU6VLur2vihHIWd/+gA4I5wPRwH2hMjzNYUUf3JkDDv6Fz7oUw9i6mUhR9+3a2AFssrcJW0VYS
iLtKBE9WP4iXQ+mGgnynG0STRmuNUgCbZLa8BIUNH3Xm4ljg0bWB1MdKFVqLyAMd7fxkiaNxDBXC
tg4JZkRvOSKocZQEUY36uKCD8NbMpkZwhBS0GHWWDpmCGvuqbFoWaJtLmturjUkkj9ESLZcKmqkI
C/2YNN13twyH1Ymz6s1JDyyeGLdXbBDMVfBT0Cg6HF4z1QOsGFOkddn31QF9Z9G85Xj2wmGq3Brc
mmVcbXgaeUPgCaCxgU7r0OEH9Z7VKetSlvWrGTSY4eYTPJJeOb3OEjKscR06ikTLjygdTsoSowgZ
uUZEBoxjfFV2k6ScCBMtUYPzG3ub03XizJtZuQpAnnMWcIcNLzOWz34/1v5LdpmRhNj1o/JRqkCX
YKIuWCDBVEWrVKFbMG3h7sRXvFlChOBA4xDya8QlAJVqHanhxfZY+GYmZPCe6yZJJnT1tt3Cor7T
/ZCEYKc02WjB97Te5B0kcRhYrHXKLNAGTLoFN8ueIkpra6HXS+F4H5rWU3ODd63930a7D4nti89l
GeZDsUlaOBMvyS+un01g7G7FDkCpfR4H1uXbWihqB8v1A1RwoyaomToFmnEn0DRVOurAcawZMdEz
JsIrEEUJFEDt+QErm8F7vDacisEaxHr9Rv3SVZNF01hF71ekzlFshz3xpE1n2ATbvyq0ngOALKc5
cQNTZXACZfZddvb9uAWJVKFmysLCsVN6l4OK5Mn1ROna3WLeCjax/1DVnyBoV51zHIHyWIOXaBkE
fNly6cK72NhRCyXON4dVpOAFt5/iXDYI2QGs/Je062CYyxafJ1JfuP/KzaTGJfwPWUgZuwdHmdo5
xvoHYzAijAf8fHFv1bapNJvb0M8U+yEyUYRhRcQ5qJh9RW8oqhmKPMvxJwEo6d42fW/I2ju7tdfz
Y5HzEegxYTv5H/QlSgK6I0fZE4jWpwPnB9LCnHD0d1uhQHTRppixfsa+nnMrIX5rOhJMDrbv97af
8cdW3OnIXl1Piu0AxKzgsXQLT+770C+Ayzdz8VnNSqHg3t8n7Bkdvs/Svlvmh/Lt0kejL9gNvJW/
Fz+Z4emxOfXmeIjMNK7p/kSoJhCqlbn9gg74wy7uNZCGV/Cr1fp12gsxFKdJtI/sn/W20GSsTNKG
h14FzPfAcKIt8BHOGXwxRZjqkff5XzLQ0tamyXwNtIyPVMfdJs4k1HZTY305gaFutVIyowhH5xuT
PfNGtNWw4yoJ6/LJVgwzL7uwGWOfPSiRLgrglmL0vweyAKsdpOxi9NOGJw/og8lw8UyH1hVmHFX/
qNh/pVf3SjqDF6+XZBBS3U0rZ+svifTPL7boo+7CDD3gvFhpBBvuBYdo6B0JwcuUT5yGyYX1vqcE
IVS1izAsFD5EPbHZntJhMAkFuFBWkewNI6FBw8ZIgFlBtM8wYO2M8D+s9rgRGTOpA7QccnTEz/e5
JdAV2Sec9idQxgrcN0muKdL9zumS58o1A7pz5u8sUFjV4NkoyWTCj8gG4ldq/t9g8SKk719wTks4
jQj47Lhpc/rE5VX99v/poYodfgkMvmH9TpT4yf4DRw0ZaBperfrtDa0tErPUKkpAQUr/XV+slHXk
YfaRs90dMgsZ7JPgsorxugBsuCsfHvmx/RkSg+lZzoViUE2NsC5i6av5qS481CS82CUPdMujXq4e
YTcmfoL4kf0FGrvJXicRfij0Rb/azBdGdgR1zxOqdfMnW6AEjVaoDJu1VRzjIS6ulSqX5OS5gsZz
11Fj8NjjRt+nx0q8Mz52qSL/0vlJ7ZxcvkpG7rcDCRkkLg85wz9Xb3uphFeENfB6AZrWyELkoJ3H
2Rls7nM7whmd1WXcpOpEZc9Zg4ue6aJoXAthL47q6wvhv7BTJBW5S2LqJlPAcsqIL52HW3QbX2UJ
5zc7/GUCzLD2sXrmNIQQotQYpBQS1hR8HEfOlCQ8Y4NhFAhfR4yLU6O8DORhhJeWBgDRBIzM3BKM
vVHtyN/bSRh7p32gBpcxLCtTwPPbG6xSPrDLfGR59xjEUyiGT2RgLZ/yL/HBZ7E4GGOB+cw7VYdW
9nAWMF/FFRukQ6FVIc7VdnwfRKt71EJtHu7kQVsUJJZxKwHeQEUABtQW29kR0u8N3tnT2ig8acVE
LZ3jKm4XimG+6Ggm1tEw/hkVkhRSwROza2WAZmPe8icPXLdK4OlA0tfymZ9mwPpBAiWjUil2xObD
xYX+FXR7MJuFxX2PyiadAdyixIjsqbLYYhdmOMrI0RJcgqaeV5bsAlleT+rR5Rsp/OsH2bvmgWVF
4mS1NxWd7VV/c022F4LpGedFasCgxbNgbEbiZ38qz2SOMpp9mF7zYhBBoLU0EaH9I5YErRLcWWpT
2CFLqaXW4Drgz3TNoTmxA2AXCH72XObQ1bipd+1dpwpfhWAbl00f8DGywhnNOOCisdeUmNFLLjLb
PxCCSVE5euu2qYvnrAasbpT0/H82u1k8R0XYuGaxgeEL3Kz28CIxhS0Sg5AHYvuYtoT4BIJ+w22z
2TZ1hUFDMOkD6gxZxcXJtB8QYPAA9c8ErRvLnJ402gweqmfYU8+oktUB/enePiMxVwKJ5VbHm42V
ILh1A4xl0l89Z+L/vUD37qTFX6tcxX0FgboTiVcc+fG9VCX7Y8RUG9j0DQ8e9DPssySwPE9W56Oo
/hisaxEUuOyLwvbQnNx0mH5me3Ot7GcdFgwbgcwkONUHrirdpb3li5CQzlDhdfK/0bhVSutoUf8t
DLHULVyL5ecH/lknYut+cKWPIsOVJGrdJP5Ya29JjjA1jfwUAULOmo+j6kuoueJ2u/TdSGmednfH
/o9iGYHIcTj3UQiVX72H66iZBsxY6834zRWJCrxegdq88UVRYkLREQekhvhNMi7qbjtOyDa1izNt
Z5hnZABapY1su3IC4p5vpqyU2R46+VfD7x+UWLXMF59Yb4zWgkVTdP3tqcm1GjZIlVbUEwCTcd/x
SypsoGY+QLypJxt+/lkaa9h4cu1V6RE1xqa08KO04gxN8Q6B1bZFFTTKjg+rgv5o78ZtM5Rn6L0s
n59g+mHbYqqOoy8fDiLhWMzXLcrZJ+ZR+PEXkLr5YpHJ1h3zTjapEEDErJZXmv1daV5QWokyvV55
e/Az5mRN3Rtn+eukpFhzSayHJclo42p/APZJFdn1kf5QWv1khBG9NaAvUDB3Ez7Qw0uoYcJ46vru
b16/rslaf2PcFuKzWhvmAiOhunKPF061r9uzmyhHO8Y4wwKAhUnbILbbI8n346CtVnyhFHdJv09P
oFWl3S/I+miypb8E4hUqA7b4CDK5pu0gfQw5QA83Cuq37VoyAvUDfxyD/QQMZMVT2JcEg762phUu
RuHJF+TjvwusFRrff6+baUuPKtY9
`protect end_protected
