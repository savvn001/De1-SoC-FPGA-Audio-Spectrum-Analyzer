��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjH��mR�L�J8���`	774���%�<���/�0+�XP��1?��=b�>�V�z��k3��� h���'{H�ؿ4&MT���ɺ�Ǳxo��4�c�C��N#�R��fH��޶E9'�� G逘��Y�Z�X�d?[�5��p#U��(�ά��4�1��ܮ�Lֿ��r"�{�8�ǈ�ةLd�V�tW?�Bfj�If_<��ը�}2��o�)ǣ���#fBÄ�T�.jI���ĶB�5;c��B�.PX�ٚȢv==O�M����n�Z�����O�պx3��jSx��tl�z��	��O����ϩh�W�kD����jv�6�ysB{h��g��=�!���V��wu�2��Z����K�&="�Wھ(�Nmp�5�Ӷ�{�6p|7e���j��	Q�\�	���Z�^9�isY���$g#�8��q������\����0b��D����F��'�^-��Pv�iT�4�n|���w@t����.+qz��,�R6�SrrJ�;���ϧ���D��D;�ōTlh�;�\��A�y@���D�;!	�x��}�D��Wx��hdeH�IP:�S�:Y�kO����	�0Z�U������E�T3!8e�$fVm١��ϻ+�	�'���Vq�l7@��Mr��/+鼪�*E��LT�R�?��t���Z2p��hCv��8�-�I�=�+�f�7���
��9��ť���貰څ��\����p��s� ��RP��P�����lz�j����7�2�mK�	������58��������[2��(;	]�Z| �0ų�$*^µ�h���?Qq3��D]�9o�c�=2n��STG��%��mv.�ᄠf�o)�3C.H�G 6QZ�ۄ�ќi&�E�8����rj)��������Q���wu�I�|��c�j�
�7w�<���몂�<g��ρ+ϥ�����[�)G�� q:�#��@�e��Tqp�k���a��E��,ö�5W�_��r�i�<A�W��q�O���D��2_o��i7E� :�L��k���Z	̦�܉��J�N+z�i���xX1�+�C��Ҕ3���rO	��@*Q���<��2�8�Q�ˍ�Fb�xZ����-
P�:�6���W8D�鮚O��S�@uѢ���/1]��TS�s�%|���[{�[֞�&��Ys{r]	�����#��|OBҮRO��b���r���8c0��A��	��s�NG���y���/�s<vX-o��U
�������`<�iQ�r�ݠF�s5���H�L�|oJ�W3�${��5���o{��G����p���|��R�n��X`��5�F�q~��2�� ��m���s�m�	o�w�w�g �|WS��TD��Xx��"%�G|wl��.�Ӣ�P�������VJ���\
\C�4D�
�B�<�5����f��� �����9�v%�[��h�;w�Ŕk�f����=���E��1���n����h3*_;�Ɨc�߈�7��2m�ݓ����F�*8������vM�k�`��Z���&A&N`�Q���+D�/ք�>�}�[ܪ��RY.##$��3:^�u�lL��Q}G��g�a��?(��~��JF��&�"���Ԙ�8���4� �fl��-Q�ͯy�z?�Eb*��	>�'���$<�<UT���C���\B��z1�\Z�ݜ�C�?z!�9/p�'��i:�0�1ўdO�`n��z�!���{u'oN��P?V��u.Fhp�׋��DK^��r+�����G'�D��t�z�`�
�cW2�������^�S�Tg�wn+'�{yR���h���UW�<��ABm�8_w�������b%k6h�R��Ǭ�����Ŭa�֍�0��{S� �g |����{l���u�Ը�e���ܰ�������CI�o�g�l��
��<�C�΁&��O%5��6�R���#$����c���{0]�-�Ju�ʠ+��|q[SO�	*�D��0�L^0]�s\^�����vj�2q6ݭz[�ˡ��j�ڃ�YZ����@l�6y�=����q��S�0A	���X��/��-1sճ!�_[w��V�v�m2R�� }�B��28����C�Sb(S�FS .��V��<��Nfή>8��w�q{	���N����䒾�5Bu�Y�LK���}�}�A#"�ɽ2(��slIr�e��k�]���SP�����Ud皑��q/�W��u!LY�-/B�pw>Oq��p�v�UtQ��R�̑��<=����4�B3*� �/X�B��W��W�9D��epW�V�DM�6&>���j�x�ȉ��Dg������ڋ\|Bm�����c�9��r���Đ��c[9Ҧ����;�nT�Cz��X�d����rC\}�9^|���w� �Wf�q��	�����=��`UF�.+�����P-("ZA�����٤��WZר��,�D�1�`��#І�tپ��ޚӿOt��ɇe��='� ̶��򼹌f3��C���_�9kr�gi��ܸG�-�wMӡ`��Z^�eD*���Tq�t3�Z�J/�}�ϔ�խE��k�����<$�r�t-J���ʲ�'M��GH�7���(�p�JUl2)�%eU�b|͐���S��}?_jj�x�)^e���[ǆ����=����
�����ib�Ї�M�$��_v&F��X
��������^�)��o����Y+�*��C�V��;&�β:N��)�9�H�i�^�������¸��p���cL���ȝ���TM�[�f_,N��Vx����<�|+=s�����ﱬe3~g�Xus6�}-WM�ޏȃF�6�q���C>�rg,n�?��d�Ӵ�NC8��u���)kE�L���L���S ��s�Sv��#�[y=�E7�a#�,jK:_ p=?C���u���QR�螹��b�S�V��pQ�U�X���q;U$PG8e�#�6�ܝ֧��r�vџë��炩CO@Ϳ���%X�`�R��n��X�� �ٷ�� s��6��8�$��֨��Ia�;�.;����۹>�eUZz��m#�$��-ҏ��OJ6�K<��Y���	V1�����]�������ֹ�B���x~#�Q"E�:����쇖�/�Y��$�d��b#��%z�!K������|��p+����0%���I��`��S�o����!�1���H_"31C)�;�޷�1J�a<���M����V�tɇ�C�V�}���_�H.�^�#�{�b��˹�����h�̙2��֧b]-��sY3��_S���K���)R<+|�f���q��Z.Q`�+��c��)������4^�^ �]�ۦ��ML�U	7UŲq�X�C�˓/d��ʩ~eK�,r.y���P!~@���S����k��0#W�a�I�
�(V�l���3S��ܖI�.��kĴ�Wz����ӛ��ⱡ(�rҗ���s��n97\L�M?���:�'��1�j�-k�r���-b~?4��D��51�Y�$����w��6$p6{�E����S~�,�n�7�N�Em�)m�����N�-z�&���ܚ���Q���
��������Y'�	� ��26���_z��AM�U󻢲����=Ǭp�D2�0��顠#8P\3k���ѝ`��\6d�*�� �ƺv����a|����"�Y$�����T�uj9r�Č�Qm�j��p� ����Y�qY̆7��ϳ�QO%��O��W�IK$��H	M�F�ឃr蚖�xM�qj,��/�{���j�ZM(!g��f�@���ļ"����xn�,M�r X�'�UJ1������xM״��@V}��oN�!��v�YG�hT� ��[�H�ɋC����S��x$-iARy+f������o�*uJ�4���G7���]��n{ݹ)[���M��bEb�#�X��
8������.[�k��=?���}�0�=69k]�A8G��8)���Xv]�K�<q�Y/��j��ϻF�\h)�O�.TŊ�"��{�$�����Ɯ �hq��?�l�0K�>I�=���w�]�h[BH~}���ƍ�0Lə�ޝޜ'���ǳBϟ�]�@5EA%v ��e��u@<����81��K���ay���y�KR�^YB74�mC�|��Υ�s0�/�Ҩ�<7BP�0���鈏� �cP�i�hŘ��М��ky�mk}�? ZuU�hiB9��&����X����7�%8h���u�S���d������l��q��}�t����.���^8�V���k�M�
5�Jl���<�F�S>�mK�P��,�,St��O�ޯ5��!���,����G�z���z�;���=��s^��X�h�j���S� �Ԯ`4�7D���?#�Q��#�<l?q\��Z�����E��o"�|[W�.��Ut�����T���Ǻ��P�(�_�j�.��7�E)'��O%zʍ�t�5�n�A-������p�O�^�w�<����kG��8D�*Hyo�M�?���e�u�����#g��@_Yz�4����ަ������vi�P~�C]_ :��dU�ߋ~4�c��C8S���=�>��f{�/l�X�=���|8+�ޡ�t���R��L��{��6 ��iL�ET�P�E%>V1����taH-l|����1=¸��.U�x��E��Q �-oy��'�w���P��W~����5�}���PU���[e���=�řބ�:�P�
l��`��ERo	ꨈ�<~x@��W��d���n�_2�L�#�w��t������U]�l��T��OaF�>L� �VKo��#～�m�E?UJ��z��3=E8��ſª^lIM26"]�CǹR��A-�<����t0�W?B�TT�ϼ�SuuK�Qj��>0�ز�:�3�T\GQ|S���A�9E���]��r�@�M����O?�ϒ�h�ڮkh�`�jΗ�ڬ��O~ckZ��(�}�Q@iC2fK.RB��BTعb��;�Nr$�����^��F͐�W��}��R�	�L�Z����7����*���J�帻�
V�xx��?7j��J�2ȢW��Cc!�AvYB��D�&X�:�)u0���
(������$Dnݠ���ʗ@碦}�
�{�˭�x��t=��'U~�+,��*!�8+�7d/�M<��fB�I�C$d�@���ё{Z�ra��w"��Y���z/|��s�ő�s�*������`nP��f<)�cn�a!�=?�ˮ+�h�S5b�{i���<�:G�%�E
4�Thi�E�frt+u)v��6���u?�x����%p����������b�9�����>%�!���&9�(gQ����5Dg'k6��ݹ8hr�;�(� K���E�E�Ɵ��A=�يQfP�����(��>���#�)�H~]]r°0��u*���mA^�N�۸%`C4��O�7�'4}�!S�]"Ay�D���w,�}��"Q14\�	���zB٭q�3dp� ��m9�n}:H�9��� �,]ז��J���(S�>����9W�;�P���9*&�ִ���a��Qv��0<Z8R�C`g$\=���m����n��jb�r��A�=G*��|%p��ݙG8S� b�(a̟�>����CMѣ��4� #
�S+�$}.,�ݟ�}xH��N(���C��9gc	������U-�5Ű"�Ǒ&���anGr��壞�>��>i���:����=���!QW�[܆�����$���֔v�Qo�m���?�Ǒ�ѴwKn#��'�?�qhN,�|e�'�t'��6�u��,k,t��[���@�(aR�Ec��x�9���� <�tT��KL��P�I�[-���3��<J�6x�[����pY��)�Vw'�\��~y3�(�ۼ���������}��rd��R�t�녔���a�g� �vM�E���t�mg��.R��VG���H���%�I���C~��!k���;	�?��|O|���9�I;��v~�U3ֳc�E9�%})#<��F��;T	�=��Ѽ?ȋ��i9i~V��#`��%p���>�ff��M��v��v�e=�,���R�aG.��~�;/����Ξ�10�f�- ��ˎHr��v�j���|��~5��E��ƹg!0#�A�GMq��_nBT^%4�:@l+Vi1֜�,�}�O�6z�XXu�t&&�.�n:�;��"nq�����(t�:d��}F���$OӾ�r�"66��V*���'�i-^.�Nk����\RayRc�*%��]�Zdx"�R;H����MU,��1~�}w;�A�4����r��_�Zp]����"מ	�r;u%0]V��)'c)OF�CG-L��3�^��ǜ��ӘX����5�Ń��*�7l��/��z8�1p1ۘ+�'FHn�x'�{l���\�|j]�LRx�~�@U"���nP 1eD��*���1W'�����7�?���ǆ�aǰd;�����7��].�ǵf�*1"yY���y�RF���ך�?�_�ܲf�$�~�/�+���ٸ9�2Qm� /�Xɶ��sV�Ad%�����Gy��=�w��V>���0��}d�E�!ѝ�n�e�/@��[	�qpW^���S��Og�M]+����,6f�Qm�0����+3<Or:@�k����1�3�V����ZQ9�\�r�i��
rl�mV\��ж,�h#�*�+Z��ڙ9(n�~�����gЈ�oƫg�Ku�M�q��j��Z8� ���0�L�';����쨇&���'��?��HՠL-$G��:h�6e��Mn�z���E�2�>왂�vg��w��kJP
�)��R���y�&/Gz�eG�9�8}�`�Q�d���0�6��&-A7ہY}���umm�#�0>�Z��Hm����xW�5�S�;���_�r ���(��c�]L���Gj����0y�-]���D���FJ���s�ey>Q0��2��}M��bt�����V���闐8�w�;׼��99]@��7�}p�[s�������q�g�zl��4	!m#�ϯ;����͠���D�k����
U�Վ�y�
�O�2X���(�0�K�� "t�G�G��ju�K]��'V���MѼ�c�LJ��'�	6b��*��z���c�Ũ��G�%PM=���˕xĠ���n�����٘1��1��\��cԌ���ͩ(�7�3��S}h��F!`3�#��-���J����k4�Dp{��P������nt�{��v�\�
�q�/W�'�� :�H�ZFf$���V��@�3e�ח���Ȥ�)�R0J��CОd8%C�D��g�'Y5����|:	�v0e��c!!<�G�/����M\o(�v�T��<�S9�9�(��$\I�L���/_om��n�c��ʴ�b�^+Z��hBU��7�kO����x	-1+>����C[L�-��?��Җ�ڄ9���(�;t�(�p�5V"�>��Г��7�M����j�'�k���C��B�/t��84����{o<$���P��z����~E� �����sŖb�RZZg ��y��ʂ��E|/-�C��<�����-�7L�}C@�r��t�S�]}(P�UV�*)<�-�T�J��y��J��x�^�K:�eJ,�Q�������������&��(�i���*��cݤ��[5=0�I')�!/~>�'���n�AO�Y�Ja�m;�Y�S���G�z�25EQ���>F�*���.x�>��'�W�&�f%LA���y��4d���ÅO���hS��VH��ow��c��6�>C�UL��?�,�qϊ@�;'�CA��9�<Ց�@�c��Sp<��H�s��Ӗ�c���K@�W�B��Y�Q߆����ĒC��)��+��@ܘ�IhdA�-$LnUH.E��3'l�Q�)���Z^Ƨ(�!���I_��^��uu���<�W��'$<�G���Fb �*�53�)�g[_`����*�M�H��9F��N9���$_�-k&N����a����	�ۣ9�B9K��̻{bZNdĘ�c�O��4'{�2GU�kȶ�� .�.�d��d5�^
*)\��H.�܄3��zʠ���/;�ƌ:�z;��ĺU%��$O�Z�<��f��<
����(~~��1/�v��)�K���>���|;�	��,���Y5����`�v�*
���c���^���$O?c:�>y�D��XZ��Tf�$tO-�M,��lv�+<D����_��˯45�&>��9< 0�q=�;�a��A�4��+�؅s9ǫ������xg��9���΅ [M賍�)�y��>�K�$͎�Y�wZ���I��͂r�ڨ@ҟ�.�ٰ���Y����PTӅ�,���v}x�:!�nd�^��z����:����@�����L��:��a>x)wL0%% �Wʫ�	��\�yJh�FT+٢�l�1�
�I��2�
��=�C��Q�z|�j1�tS�P��T��N$����C�~�-�^3IJu��I���?�Z�4���E�h�&AmL{�	U�N��	R�AZ���Ǖ���G���ʶ�#��
:�
#2�`�}�Z��qF�E�`��&� 렷R�|= �������?��fh�X�ɮ���|����?�'d�uœ��#?l�|̲X��7�xE���Q������c@�w�0�8˭=���	r��~a/ӓ�>L.FBɴ���8����Q�&�Zp�z]��+�d��	#�ˏ2�Y�g��O؂0�����Lzߠ�d�S��N�/��d���������&q�Qbj�0�������
zR�X��:�\�ؚ��_����?!�0�V���^�A �L����"57��C���sDX4j��H��L��siߢv���P�����q��ʗ
�'
�ɋ�i�YP�#
���p���m[D�r������I�ldC�����=����9뜀�ː��#)��b[��~��R6�����6Ұ��Z�C�@^t�y�����ީ�%34)��:-�J*$Bv�����y��]+פ�ln��"��[�<���̻��59;�W�T@�	1�ū�Q�1#����=��H+�z����R�F�N�PgZe$o���aHڱ�~�'/�nxJ=I�6;�014��IX*8�
auIO�f�Tv����Yf�":�|��oA�f]��fb��U�_�8|/�Q���L�4x�s�V��Z=��U�0ҽ?���������z�^��b�.��z����6ij�t����- M�#"p]y�vDC}b�o9.	�JZ�( ��&-��K�߮_�,$8�k�L�j��-��:f�DK_�$jT� �e12s6_�8� eZ��c���g{+l��rƑ&J3���w��A�J�7'�I��!�b?�ň����c�	���)1/��8�DC�qo��,3�l4as;��۸�㺣ȋQ,e�?�qR��5f���_�.c4����r����-?	2 �D�����i`�()�L�Ϣ?^Fk��Cl)'� E�9��B���Bne���[+�?�W�4��$S�iO޸�5J�)���Q�v�H�m\��O�O��h��w(JKx��n��[��!7�,��E4����/��&i�+�-�l����Y���WQK6T���M�&{Z���u7�hw��FbCK���^��K���}(p����p#4�3����R��f�.��ƃ}.~��I�RBu|�}wC���Ჷd��µ85r��9p�ǗU��rri�������}����`�	S���F�Kg��_�!��XI��/��o
�U!��*6��
��h����kt��y*��J5�XT@��`���Sm#�s���i�[5���A�R�a��YM�&��Q��w�3-<9k�]����vĺA��a���ѝl�x�]��䓑��<Q�(2C�i��d�f�7N���xG�������`�/]Gߏ�Ɋ̩n���sOґ�k#I5e<��!�B0{��l�Y��N7�]��1��%��fw���*R� �玧M!�^�_|9Aj�)�����j��@ V�b�T�P�eҥ�7QY�l�+D,E�1"��`�IRƃ���Ɠ�I$Ǳ�E����:�eT�l���]����W%�fn�k7R֟ASД_�|��\ZШǑ�R(�
�|P__�y� �u��٩얃�	�����=�ߘ	ߛ�r��_�P$r�P�I	�T���LW�2�!O����3M��G��z `I#�D��"�Q�d_���m����!n�A#K�qG,��.��ߣۇ�:���<�wG�JѴ7�J�GiD�c��3�
E�����bBk�e�6Q%�&zB�Ncy�u�	ӑ}���R��[�}`%��m�bD/�!=�����X��,�9Xk�V�Hf��-�����q��5@v�gޱ_��c}lv"�ĦW��[�,�=�F��V ��6؁%)4/�Q�>���a6	��7��s2�++^�0�8X����xRPnv�2���gV���9�(����zQ_��XY�cGR��L�/UIw�A=D�o�ٮ�6�����2J��jjy���K��H�<�ܲn�|L��V��2�N�K-5��;�i�Dor{���L����a�uT�*�^�Ռ�6vӨᲥ����+<��kU7C-��=��|N�I���r:m��2�J�&&)�)J����L�+�/&ܻw����]�l���=M��e�?,�N;mfflp����:�o�Ƨ/@�	�1]L��M�=~3�%��=D?*�b )y�&���T[���A[�'K��.="?��R. G���R��������dIЀ�U�$�+�%�*���`u��(B����SJ�M�w�`%��v�j^�Pr�f�:Z|�}lYS�x�\�m9���m����.=�pU;��] 	�������Y���UkR�=�
|�W�{@�!-�DG����4�J-{����� Js���_N��D�"�^����3X���@�����a�$�f���U꒑�Q��V=�!i��F�2%�&��+���Z%�M;�o� A�#�E��2���r?��6]l�<�e6�w4�x_GT9�B�F.%C��x��G),�ks��� њ~'�d�z����wP��L��fbБ�xM��OP��Vl=w�X�����_���&��0ȹ�Q��֖�S������\��b��^�L��S����V��e����쮶���/-�}��0�P���ƙ�L}q�m(GvE�jN�Y�6s?
W�W!�������d�]]���Jz�z!����86h?K�ƅ����{����oP6j��d2��uaJ��.Rk3������2��]�o~�T3���*���D&�b��gm�����@�I����.���d��r�<��sU�&�+��G�~��"��9�e�#���N?'^��K�w���0Τ;}��+��s��'�aq�F@����VX��A����"jOj�fv�P{d�f�q�G�-PK�����^a�0��������j8�4�w��J�>9�]�?+,Ap�q;�Ӝ�a<�W��O��"���l�i��U
7DѺ�XS�W3&/h���I����@�?~��'i�/�A��$��ƞ����`���'.��˪�Uie_��ISS�]�]Z�������CT��������<;}y�>Б�c��%�pk�t��}a8��9,��Ţ�$M�G�ݸ��H<t�G�1�s9�M�"����1>^��l����n_ӲeF����ʂ)���G��^vGx����MF�.���%uHC�v����"\�W���$��������DU���<�ϧ
-�x����1�A~�Rf�����ʂ�J�y@ǆ p,v��h㖙rv������� -�7ǴK �R�M>2 |�q1�)<���,�r���)���F����CR`��t��� 4� 0��UiQ��l�ӆf��q9O�:���e��W��-��YFSm���ق$�q["
u�0���$����O��7�C�o�){%#��ŝ'��h"^?xú����׃�5�`���/���K͊iβ�����b)i#�]^�5����"����VX�1�0��Ϣ&ѕٷ��2>.��`us��8�@�Df�R��i��O8Ћ��A.�]�\�\��l��YH�n*Н�I�pA"�r
m�>����y��QY���O��*6:U���- ع)��{L�� �>?��z:�Wc��`���牔@���C��KL�P��v�����zl~�&Z��
�?���R]c��y��}�ٝ�����ʤ��a�/T8R_�Bq�1��d����Ȉ�6�Ҥ" 2�)�1�mC`��brc�+����33<+��?�A� d�g�K� �%��{C������*�-���F�x!9��u��!y[�sL����]��}���Yp�C��	�����+��~���ܛ��ފ+V����N����҇���YA}R�gi���<0>L����qt3
�����_���@*�*z���������9c�|n�����U4ψ$y?�T���M��"6y�S��:��
�b��K�� }�2J� �k��Z%����a|k�Lv�)�����(
�S��y+u1#`��78o滜eY���x���DW[�d���]�����)Ixѣsn�"4v�	�9e�Jpٖ���Mb��}�t��nL���	;Z��g����A�x���!ir.��3z	�݁��c٬�(�Q2o)�B��-GE�*�Dw��>�x
�~_��6����j)��cz���n�I��-��Պm�ٔ��x���,W�m6jWG���6���G훀�G�r0����
}B����,�>���
E'�����g{��{��B�/u����һy�7M~|j���\�cTk6p�ƾ�)�1	 K�p�@لd��5�Q���t��d���Y�v�^��u�S65c���>�D�+�����X[�ͣǑH���ĩCj�u��hT�Q��f���S��r��2��tգ�����i��Y�rB��{t�k�сyT9@RϨ���Ȗ������2�A���L;�M�7����`���!�^�rQLX�}��#3!�;!wS(W�~����3cNI'
3��	C��/8�d�����~���-(Z|_�5n���0�/�&�����'��u��}Jg(lM%�T��1��ը�8j��ţ)yb�-��+�y�1��4X[wϐ@�N��2'	�Y/����Nu�� z��:��6����r�Gc��~cH֣爠��}�E�w54D�]��P(���v�Y����Ux�*���98�Q�87��C\��ZPh��4��=��}�?L�؀���Gـ��vB��u���Fn=��+1�^��en��ӆ�����"V^z��!2�xJ��VXUIm4j�e]���N�=D����_�En:]�EV	��,%e��R���i@���S�(˚ ��U������gp�����������\[�EnIޭ��_4�ш�n#�ƨOI�֌(|��9����h�RN�eF��P.U}��qP�NC�.O���k��z�h7��ͮܕ[����U�����hC��S�܅ٻ:s;4���.(]:JQ���a�2_Zy����(�ct�V�"iդ��k���c��g"�@���ӯ+��%�u�ї.��D�3���X����KF劑�0��yE�g���@j��8^��!<鰫��Ȉ(N9�ӗԃ?��Sə�\�c��rNu�3�������J������ǝ����/�V/uF�8C�b��2Kc�E�^Me�£g�܂��;؛���d[x�����bD�A�.��
��א����Mv���ҍh�@]'1"������a�ʉ_د��m���,�g����P�����bi�m�-���#]�M
��2GlO��@Q�M�\�s��Z^/�y�H;9�� ?�H�&��Q�TI�Sz;E�zM���v��C�n��j774�i��Ύ�O:�@�@߹�]L֌w�S6T�k��G��~� ��g�k�A��$r��@�Є�u��g��Q������� *�:����/ss4oA��к�Eb�k,��̆�0�ޙ�[� �'�#�Bdޏ6��@�����%W뒭��#[�d�w�Z�X&�(�8!�$��>[�*�DYAx����lN��rб"5�_X��]r9E�*r�ͪ��K�c8�:k��7�1:����)�Sv��7b�{u��ńfˊ�(,Ї��߃O���7a��u�%�t㌇rB|�X�L�) �ů���%�ǯ�l����/*�S��Oւ/������_Jk�#9thl"=-�.7��A��E5�_8؀����6��zgyڗq��*O6|��M� �s�sQ�Yu�{��e����o�o��+�	�/Q"���}��.wM7�$�o�f�%|���w!��8�-�O�t��m��?_�|ķv1�_N���)FPxiA����1
:#�:�����}h�����ݢ����6_�f$����?)=;r+��ڒ�� �h�a����zLzCN�'M-�8nj�S�h�U��?Si띔#w�6�X�l�)+K�yݩ��"d��t���[8���Y������hJZW� ����ũ)D��[��6����L���7dNz��!��y���q��(`�q%�RU6H��<��2t�}����/�Ѐ|ux���<O��29+��L�Ҧ�#��q��k_�8�԰
��Ӟ�X���aiy=�s&�g�?�?K���ZΈp��B���<ݡ�
�XMS28�Q�c��=Ǩ
�4v�M���h=6���Q�
˶_�h{:u��{�-���O�B��``b�R�/�d���5�Ug*�m�Fb��z� �r�N��ƃ��\����n�I4���T���5Q�e����rDnaN
IZ /(q7�eg�Z ��ƕ�#k��~�"V ()&�����tS��x�"���,�JW�����8�`Fc�C�8�0Ȫ���}�7��78+cN���ws*�I����u��V)������<��!��e.�B�.p�f�Ĉ�~���� �b_%y�J���H�|������+�V�S��S4X\��ƲW����%��"��L�*-2}aJ��npΦ��ok!���(G�`L��-�J<�B��ά���L\.v�M���p�\^���6�X��5�>{z톪��d���w#RhM�q�OƦ��!��v�^���C�/Vp��荗��ggZ�\¹yJ8k���s�UG��g�i�Q�tgϼI!�pO��Y���6�UM���u#�-���s�F�1���yZ���W�T2@Q!2��K��t�K�O!e���=0��f_��˱�ji����ՂkQ���M���>��Uf��᰻!w5D^Q��|}����s��t�s��pMk���P�vȢ�6�+���͖\�1�� �#H�t��(R�Ǚt���w�g풛�N�bv�z�E�~K=lR�RO�^Q{�� 5���؝M�vc����,u���W�*Tt�R�h���^�l�
Ͽ�ϧ�P��2|2P�m:b��k�"�N�R~M�6��wé s\�
�;�Y��#��#i�U��E~��YP��:�ϛ�H� �u�|*�aIATbZd�=I×^�e���	S�)��wm�y�[4�6p�Ӊ��!i���K
A��{�hI�[�8�CQ�N���-��F��"Z���5������a�,;.��-xD���\B���'Pm���hF�P�*+�S�Lb��h��Yp��˒�0�=�n�8��_$H���������KX�׺g���Ē�Cd�m�e]S�r���~�
�}�{x�+�Xv����z~7J�j������/��%�Ĵ�#eɛ�:,��V�4������U��0�]S���c
��j#עa�*��k�!���oٳ�q�N���Z�B\����o�EES��x��b��`���bdk��E���B��p}�@��#�?�v�H�`rP��~̢��C�R%`�8�
d��:={G>\c�9S�#�-�OFjz�"�'�M<>�6��B�y��6�vc�V���w�X2l�]�+�p�d�a𧊗;�C���;�ÞT}s�}~�P���Gi��
KL���AE['�7Vo�|�J��v�?���{�1��2���ã�7�"���+;zJ����zu^�g��6��'��&V�
l��n��@v3��0���؎��5�<��M�I�ـ�a�p,�"��-����"L�M�h9��D`kb��$�û��#���P^e�7x��L�<DU�c�:�Wt��4�Υ@H8��c�0U�����{D3�r~���l������@κ4X:�J���	O, >�4��D۰w�� 4�${w.�5V&�F!G9��
.]B,�a��@��Pbm�Z(
qP-��;M_�!�?�;��^�.�V�o-Z,�ڐ���f����̡���
�J�za0��vy�,pseK.��ݽ�����6o��2�a���x��zb�ۨ���+iwx�
���O��O`S*������a���.X����ã��]:�_}P!�jM�m��碞��ho�!�Ͷ�>f��1@*SK��qƃ���>%��]x$��#�D���[i�����N�t!ǵ�\�� U�X��Z���a��D0���Zj������L�}�g�� T����Q�$v��.�L�k��b���}�Ǳ-�Z����V|T.l��i���$ih0dڔ�J�[��	��-���5&���%��SG-��=>8�x��Om|�=�^c���%�tY��K�������=���~�JI�`��b�]�*�q�Pf5����2�D�#X+2�g��Ʌ�W�2�`w�-q�H��Q�c=z�X%��;�!��@��[�A%��4O�2>4<���{��W�'�UpF��c��?��RA��u�j��w�<�@_C�dX�e�Z��gCG9|�>R��uM:�	"=/O.�	���;j�B8s�u�����T��%ߌ%K��I ��ɔ/o��%����w�z;���X��q��^R
JM`&�������7g���F!i 珟�Z-X�����\��Ά(�-��C����%��Kj
��|��Q�����㿶q} �1�F݌�w�2��B�l�B�}o1��Vr����Xz�<(1�S�˪�Nַ��E�Ly��� �ZOܛ��@T"�zo\}��(��2I֘=���/^�.c[�*�x�Zm���h����}��]��\�� +@���c�f��c�}e��Jj��6�Ćn�}|�3 =Pm8hթ��`����jX�ٲ0�'8p�w�'��e�fu��4�<]�8%�QRg�"�>+� ,���`ʤǭ��>�М_t�cu}	�6��s�z͇"O��M<�/����/��^x�����.���L��X�i����={*�X����P�-i;�釞?a��zB]�p��QGL�Y��t��o��hB��h��q=117����bJ��I����]�ƪ@�U~J�Ä=E5/nD���t�1�Xw�s�0�T�|_�*e����O:���Z�{}]V1�`�z��"���ߗwr\�|��l�ā�c�8�=r���r ������FM���A ���eJ�'��#��(���!��J����lvDJ/V�$A�19@��5���`��U����*��,�_&�C�Ԓ��`6�I���t|Z@�kD8^9�R���;3�f[���r�� �%<�l�z��}ʧB[!E�Z���:|̝b������w��d�FAJ�2���{���ptI�ë&�'�V��'�XTL�����f2vHY��lО��NV����$pV��3+�%K�?��K�>�Y�� $���CA^�O
�e@����9��Y6�K���7T��̆��ʯ�FUn��F���:�� ������	���v<�;y�[s��7��S����!j/��E�����!'�o|v�V���BJ��K�̽��h3M��=�p-ߘ ��-��d�#(w�>��Ga�ي��S�ц�ӭi.+��]ʳ�8��-�4G���*�v�l�-��'|{���q��t�N��l����d��^�TY~�dCr6�ܰ�A��xH}D�腄%��`�j�j��]��V��VU��sۗL��z�hVޥ�K;__#w�<��%�FA��|����2�4���m�\���By��pmP���`5Wi4���1w#Ȥ�'��S�|���}���0��9,zGf?������p�%!�B�tm�W�����_y����e�<��`i!ӄ�ADI��LB�W �'���˯]���ߌ�8���h)��������a���=J��V����zo\'�@{X*�[�E}أ�}���Q�r$�%qE����u݉��+E�iB�d��9eR�����?s�J�ڞ�J��~'�߷yfQyI�r��>|��0�A,9|b�{
t��oF�X5M��V\Q/�t{�(��RSyV�"��Un)�ߩ�Vz��F:=���C��X8��9�~�	�ㅸ;���nZ��֡���4��ʲ���YjB�2f2R�Gyr���,�d�ȴ�Ƨ�3��.�5����l�na=�4 �� 5��8��sz5_��"[���z��GO���>�Q���`?��(��6�8} E���+���|�����!����>���A#��rl�ա����l�ɱ�����ڳ�\ �]ǻ<�v(B��E4�NI�d��<���A\�	p0��90�IT?�� A�e�m]?��~<�k���)���!��p8����u�+��H��!���0�ǈB�r��Q��j�*������~�:�'E:H���+epx�Ox�|戊�C����B��;���>o5�T[�P�\L_�ML�]d��}�������KR����9h��P+�m=f-��t~^&��84����3,.�X���@�ھi#�5-}�b��[���`��~���<0X0r4)Lv�|�X�L�g]ΛK-����]bz�)��[���7y<�� �ioxF�PW����~Q�]k�?��37����ď� ��w�%Q0���{�P<�u��DE�_�U���)*O��D��!�B�}*�]<*�6�'3�%��蠔"^����^{���ry�n�2�e���Y06��?�M�k"w�|3JF���@pqΛ�tw��1_�N��}qI�i�}�we����;��n���5$t|��W�F*�t7�·#D��+�:��9"��>�0�Ob��v�]�ϲor����Ȧ���R4��MU�m����E��XZ�p`l�T�:���y����1�d�r�/��?K����A��v��A��(��V�*24r"kˋ�@4g�p#�I���{O�%�k�ss�{�}���P��-�T?�d�	�5m�n�,�-#��=��\�e4�g0p|?V�&�w�Qu��)x�e��Gv���bh�[��˖�K���3�?�fAҧᆎ�:�,:�	�
}��|8/�@���Ä4���B���f�F.�|�N�
]�X��D{n/�H�<lTJMzS�$�zK����_P(C��cQ6���;��W��c	�^�� ��qw�)�-o�Z�~�͟
e�w�k�����d���+/XIU�����Aדpx;x`�L����<�G�+
���s�m�2��"e*,N`l�P���I�P��o����	e{Ԓ�كڨOhڙ��u8��GPJ��+�H�B�}2ڧa;�h'�C��=7�-O0]��L��IL��匩9#��'���H��Ң�`+����v��RM�S�Ьk�h�j���-a^p�=��ۂr�^����$�h��E�pE-���f��3�C��T��)4���S+ۙ���@I6ʕ�UFָ�7��uc�s��I��qA�>���eB��vǡÐL��-k���O�+A���[A�L�R�~ T��4k�S�o8Õ
R]���pJ���`����[AK�X�H.�<VV2�
nS�Hq8�&��ա�I���ZQ�_%��2S�s�.6���s�����H*� }q���i2�.ͯ�Ӎ���a�����d�e����{�.1*N"q�?��ϡ[KVՄ2M�&��Ɏ�V��]�j���w�-+����`��i���~�qHe
]����w)X�^�y#�bѨ�$�c͏�m,[�,R���EL�G�K"���C�)�2�lC&�6r��iA�z�D�7��XA%�]t!\�Y�F�P���5EF���y�[�7���_6�w뼶�#�tK}�X�5eC�9�K�5���r��u�Kڙ���A�*E�)�Ȩ2��t�P�r\�FɷFx��9'ޛ���LŚ����$�+�7ˡ���}BW�]������a᱉U�����{|�-�/0������[z����ލ�.����l��"�%N {��F.�fao�r�.�c��@ͶlR*)d�Θ�%�t+�����d]��!��>�.*���&��ډy���	����x�=1�3�4���Pg�����R�%]4�w�.�콇45w�<ƠZU�HI�Ϗ��Sf�b蛣����V
��H�#@�W��s_kM0��|�O�l��7��j����xɥst�������ؐ,#��_��`A�3Y��?�S�����A!~p�L���g�8 �O�a��D�AV4(�8�N�f�ӃׯSg4�H��`�5���B.H0sii�EYс(��1�D������7O�Z���/Jb��T	��g�%�9$����'�UQ��(e0�d@&�@<���64�ߙ�� �&��JsMAC@;r�8�L,�[E]�Zz報�T9鶗��zJ����g�lU	�G���%���tu$a�gI/����iΆ�2�w�mɼ/�����Ay#�}K�KLK����\�2�]*�0�RŸ�D��|p��t��0�`��R~a*��{�:tH�J4L�sd
�>�j�;2�Ec���X���۳���׉7��w��r���{k�Q�4/����Wچ_�M)l��n�sIC����9�3h��ݏ��+��E�Y���09�oс��� F�w(B(>Q�0^6+J|�!ʢ����bc�c��$YM�������e���;�Gr�O4�$sQs1��1��WeE�����y�&���x7��*#Ǣ}k�;�'��e<��F����|�B�?��J"Z?H�����7>`7B�kyD�W����)�]Z��z�����j>�xu2�	��<"jV�<��Fb�}�8��C�����D�S��tR��hp���/Sw%�LE|=�r^�i�-eR/B�K/�F<�A��p��K��[�=X!	ߟ�'*�ːW&�a?��?�)K���Q�	������ f������g�:S�=^J37�j	6/���l�b��HzM!kwW��:����l'��ԝ$�T��L��J<�myQ#ح�L��K赙~�Ok���a�;*]xj[ʨ�ɡP7�I���}��CY�D{�T'|N��!� o�Bq�g�K࣓�09_@�w;@��m�&\th%�y��PAz��U��Y̻��x^�_K�{! Ӏ��Ԙ"�W*qQ�W��اNfD�|k��m;ѩ��Q��V���Q5tB��r�`o,͚ׄ�U�:C����}��0x�4�a��8�ڭ�0|"�� �;�0j�|$�4_�Ao�-*�.?&p�8R�v�j��P\�&ۀWQ��Ӛ���������P�o��oCD�#}W!WB_�~pL�-�t�	��*1y��t��L�b?�}	��<"e ��.�~�������\�i��4"�/�����ш�%a�9�~<��8�Gw;;��lِ�;�����~�Z�4�5C����{���N��	��<ĸX���23	�X���I�5L�:(��S��1_S.�e_���cr�~3����b�x���v�Vjx�,��)�9AR�*c����pf�
���bMGN 4��^ꗷo~�E��hZ�ӀZ��!�-1�K���2b�TEЗ2���3<rE��Zf��|��ei��N�!T���ݽ4Ez6���d����B��D��-�A;ɣȂsNV�d�d��Fw'	
�J�A���Ϫ��`�����+YJ���7�=k�m�Õ��cA<����\��jv lfs��>��i1!���ʬ}��i^�� 0,l6�&��TD4(���\���)z�Oa�ˈ	���B�ũ�ke���{�LD�(pn5�XF�g�;o9b��`�'�ϩ��$N����CV�Z?�@}�����<+y�M�Y9�\8QR�����f�EtG�2`�M۸����&>p��T��������C)��DD�t%��4�o��U������x\F��7S<����i��;f#Ʉ��ӗ��,f�3�_ˁ��4r��1<P�l%�Gt���ɢ�!J\k��� y?�ݏާ�h�
�n�$��NmmE\��+�����:�^�����k|u��)
K�Ն\��Ծٗz� g�Wt�y�׵�`q�4_�%�+�Rp�>��XCs!����vM_%�͜��bPs��܈�EHS�@�f.���';�;�1�y�+~�Q:�`!�渷��Q��0��C<G'��2�:�5�!X�X�W��Tkh�ʘq�Tq&��DL�w~D�N�~��*�t�q��i�q<�dD{�гF�V�E��.���w�lÂ��u�F=��5|�dL�Ä�֭�.<�k}0�j�k��u)a���`�����ف��!�s���I�+ܚ���u������-Z�6�5��|$������,0ᥪ�/&9-/TP|���%RqjKt�,T̇Ü|*���>z�]O
a;͛z��Xh��Rf�f��k�N��&,�4%���i|��:�&ٯ��ӱ#�Ad*��R�Ń�ԯv?�"�����a9>3�Y�����n�#�y�M�\��Ɲ��.�/`���Z�V�_�dM�z�&�-���Z��l�-{��2}��|`-�l��$9,��Y2g+�nC-�8���~gʶI�]��9���t�ײc<D�j�'��VtԺ%���Q��'���רz�2��XV�r~�b`9WaC.�+g	y���_�D���ҹ������A�ɺx�~ps�j2�d�$�b��vNG��&H���8t��|�d���qg��?=�z���u��Nf�[��ߥ�q����s�w�1��a��-��wo,G�~r�[�?u�-0}��$�+ȩ�=[�D��.���?��%����b^=^�/���L
�b���!���#io�f3�N�x؄�oO��Ȭ)���${-e���
�5�B�fY�����v>,PL�����1F�������C��R�����C�]u�����i;���V��޻�}�8ίY߀I�u�΢�/�t��oԹ0��͘��VτIS$d :l��~mf���X5���C� h���O7�X���H��~��d��8;���o� g�&�^�����W���x��|�Y9h �|̽�aQ6�~�c��0�<��Z<�ޯk��G;��� i,
l�,��C���̚��`�����B�a�n��i5���3����=SqVFMG���rww��A���9bޭ��I�r��>,��J��Q��-�P�L�t���9��>�[��$
�NA�Er"���wM���A<Rxf���P��Њf����Nku��-���2>��2tP����x���ѓULX�,R���v��ߤ��@pD�ڬl4\�wbqdQs*$6[�⊨Ww��K��pm��z1���w@����y�[��8,�+<�V�X�	t;'zHw�1J���Rm��"���4��8��a��<Kk�z#��h��U��?�����턛IW������%�.6�L�#��d�\5�PV�
�uB�@�`}<S>��@��#a����3���K��d�4bfIU��n���Lx���R���I����E%"�5�k�{���EN�5�d�_������"9���f��g�WiQ��>Y/3������5�ؼ0_i�l��J�L��$^m4�bG8����
��,�3����:��W
~Cn9��+wj�ל�����m&�H�M��0�g��:�{���:��3���H���w�z�$�YF��㽝X�g���cWǤ�Վ���2�	)_�-�h=<3J(���$�vgYǜ]��i�`N�n� b�1��趸�@������f�KB9��%JfUMT<�\�v��t����~Z�4p�+!�_������KL�O0L��cơ��ȺґՐz��M��)�a�"�5�YJ!}ƊtS�����v�>�>��M1� J *�Vl�ΗN��L��$0H�Y|Ѓ/��j�JB��O(�eGp�����g}q�!��+)u��=!,cq�D�v���`�����H ���޹�>>G��~�ƀ*9l|S���_ۯy��i��Kc�&xK������	f�a��,,L��oHm>1C�u(���N��8�?Xsܬ�n����t�:W{lx�`��f�$$�poh
�H��쏬'���dA`ؾ�!d�z���nA�<,@C։��ƴ�`��[}��ic���뜯��r���\�"1P�N�3���	�P~�+�~��ބ��X�3bY����������?�+u/����?���)�2f�wцg����4� e�xH֣��̈́�$JK�F�&&�k��vD�(A:�%u{�q�U���,�#g�|���#�Ԁ?Ǻ�u0rj|ζ=��\Ȓ��\+�m��jmQ�	ޑ7��`��۪���
q�N���Q��.����<����g�*��?�M,���~Y���HS̈́�׬�L�P<TZ)���c�e�R���CQVp큿���/}�>�2�Z������H;��DR7��0�fΐ��^�������,CC�4_�ؾ	�Y8
�]Y�D��??`�3�ov>��v�#B�"$"!�y�y�jæO��G�>;d��Ґ#�%�.���Q�>'���+w��UX��~H��ԑ
(��8�Y�v��7{��)�AY�f~;,��ӟ[^�i�P>~�g/a�u�n6v,�/)�:l��<7�J��y8�ƃ�g�g���nP�����ʄT��#ҍ5�!��3�Zc������d�� xl��,3���rQ����R |�d�/Y���e˝t�og�w sjR�n6��4�̎�X�������	P�/^�4"������A���7��c��&��̔Q�L�q`��i���������r�L�3�����1!��ɞ��Ґ@���F�xP���qj`7wܬ�C�{�	lC�����M�3N�JpM�p�}9G�pA�����|e�
�;�3.<�� K�
��� �Z���ȭ%�l�c3�����m����*�-�u���t�͟� [��mq���9Y!��.��7�=Ϻn�X����nvi��<c���Lct&q�#L�AE�������	^�\�5+e���x���D�U�~��-��8#o���n]ܟ�����{%�'2Z2�*��tP�̈́�ӒǸ{�#�>sr���f��
���euY�(����Q9\J��>R����d	m�X�ao�� �6�6�*�Ņ�E��_ק���^S*���Ѓ�<7���U��&Yti�2
����([u'%T4P� ��C���,�ʾ;��zƯb����o�i��>3v
uEz"�� l,o���Ȩe��M���ĉ���=%��7K�]�B��Y��"C��\��_;�D[����� �9��W�����fVS���&?�$I��B���&�6\@{;��������~�:ɛ�KHc������qKa7��~�P?�TЄ��о��l��>�"�c�N��QFM5�6�	F|>SՙAMI���o���5N��삕@��IUa3��	�p�=%�����h@��ǝ�P�,�Eրv���GWp��U8}W��n��D78HA�>Y�|�I��-�-8�ֻ�{i��$�x��_��άCi�/�!���	${���<fG������Ž�q}�6�IC����(Ʋ�Ku�e�G`џ�ZW�ٻ���u����+��$u^79��w��N�Xjz��]s*��Fh9 ���?�fN�eoR_6����c���B�X��Z��l ��S��[9����<��/2��=�����%�*��6�TTi���R'	�UA��.$vǖ�L>Wv5�%ҏlq.XK:�"S��~7��`���=�c���23����l�g47�
 ��٥8|�������l�s������F§���I�埨����G��5�X�����O��}c�r�"��V��*�bC�/���QrF�w��v:)�����V)�q�IOR��E�,�9�s �bK���vD�aO��c�t51��8������T"���md����s1����G�}>a��W�a5���
�t��W�^k��H�:Ny��EI_ŵy�Y���V��>��-�8߶�~�.�5r���_���?cg��p����u�.~���ے3y˼����u%8Wxh�@ԇ��)>O��͐Ҧ��k�FVo�
�@����$��
��.{Ʌ�H�ci$,��n��Q7�!��w�ǘ�R�_�!p&��׈7����ց���f��W�7��^�Q|]��k}�IHy�C�D�ȕ�!3\���9|V{�g�Z��)�뮊��E��$2��Q?계�5
����[��=�N��ύ/qP���[v}�H��8�����'�F�`�R@�;�i��f��1~3�y�Dq7rK�F��g��@?��CF��aE�i�/����b��iJG�ð��-3`\�{*s�}�h԰�JĔ�������b)*F3#�륬9/��ѩ����\����Ɔc&�E�?m%�v���dmxh�s���� �#�c��w����^�$>)��P��5�Q��EP�g�� S�q�� �miX3�7�0���4�v��oz�t��Gz��NL�.�6�k��`�%ѩL���j�۠�oG�v�����me$�W��N��Y4��c��ͧ�j��`r)+/�"#[�m���Q|?l���2���g|9TE��z�!_�ɱ�x�+�kiΒQ�C����8GG����g{Ÿ�~�?,�\��{��ǯ\YvjS��9��y]58M���m%��셸���.�?���K�S���q]�=Y;����E37����giC��eZ܌S��U���Q����򈁖�������	��!M�|�n03�@yh�����w-|"�U�����\���0M�^��)S�_�Cj�T���x;�c��ŵ96�t!a��Î}�o�m����o��2㹣KطV���\�6�5K��&��$G	��^tj�*�cUC��L|�;G��<[���ML\_`,�LŠ�y���8t/1�nq$�K�aE�AO��.s@���-�V�pyAH�����^1p���JM��D���s�9������]e�sɮ�A[��� t�=�|�����I��?yG�l�-&aXG. =Z{��D��}��S�V�S�.��K��Q�]�\Z��@�/�3 x5tx�g�/�����l��&�O>Հ3T�Ɉ��#�ҷ0|����e���(p �`�}r���_��Q$uev��VS�&<����Dѐ�Y��C�x���(T`�?���ѩm�)a{,��z%�O>X9�F�f���f��fs��ld-8ƕ>�gu3BO�}�{W���L�B��YV����_���h
��(��)f���Ť���\JL��F���L0t��͕�����@un3�t�p� T�B�(�N� N'�j?�h�>�4p��:�sr$��ny�V�g�!�'�ԋ��B�w<��k��ᕠ[�Fn�x�~�{�)�p��?V���8&$�Wb�b�n�Ht>�b�e��-Jxa�B�VjzQ�.�2�=� [�c2���Z��YJ��?�oFn�H2x�[W��,��;����p"�Hj�6��1����1� �~�+�hʪ��Y�" }�
��.x'n�Bp[.\��KQ(�-��0��ᐻo�)�TFL"�.��S	��_:�??"�+�VE?S �G��e�~�a������"I�Y�E�ጸJ� ����e�F�̩Ҩ��1v��`�/���CL,�?i��?Cm�h
���/�u�ޚ�P��m+&���@�P�Ct#��p�AG2�;{�orpv��`��"XZ��
�p	E�'����o�/�gA0�j����(�
�0��O��eX����������-"���Vq�5�÷t�Y77S��6:0s������7���w�����,�����J⪶̞z�0��Q~.�~��S�w�4��Oz%�p�y�;p�i�z�FcE���x4��DI_�5R���C��m��ްY��<�ad���t�A����+ľ�� �V���ǝ�V
d�Nw*�rq,��G}&�F#QV��"Q6�v/I1ǟӏ��o^����$�d$�?� z�W�B�tCdx�����A�@�YG�m5���=o�ˉ�@z,U��3ř8��i�X7�[�.F����(AѿHt}� �Z���Y���w h<6�X(���+^g��������2���Yk��]4tF[ lN�㌁��8�+c&ɭ�����Y��^Y�&��rpk�0�(Yp��� AuJ��/~���uwk2���Ac��C�<���-^*!O㒳)�_8����,�Bh7���>��<�`�g0[�[7j���9�	�8�v�������E��n��z�Cb�B�6!���ۙk�D�޲�>��|�i�7ݤB���I��K�H�誅h'�U	MV
(�����E�lm�R�;?�h���eq7�L� ����Q/P� ��Xy����m �s+������2�GA�㫹	 �j��s�Y2ල��y$��S5JCK��yѢ�W2�-�9Y֊M�4U� .$F�'�O��bp}��aN�p.�6�{�s�t�M �O�H�'t�5@�E��}���]��-�c�Y����F
&UP:s:��������i@ �.�J����Z�hk"����C%n`gQ[�L���.iQɪw�҆C���	�d�d4����z*�^Y�}s�N���G�A���o�9'p�*��6���"�h�#�o�,{7�ު�ݍ��
���]L5��*���Bb+�C^�-Ke�*�.~��-�)��s��ymb^9AfH��&	~��dG�I���n]>lu9ˉ)��ln�*�YχͤHem?MhA����	}9bg��yiu_��%���4&�J[���* �	ȷ���3;�!�40����J�x��cK��Q���]��l?�
�?vm�O��PsX�C��E��u����j�5�^rk�w�e�R���bǒ����]"dStu���|��t9.z���ׂd�� ��-�q�]�B	5ge��@/��n����ۜ���2,�2��9�2;`���l+F��?YQ�c����-�aI�#{�L!o��pI	�k���zy���Rp;/��cC�����G�C#��
S�/H�Ȋ��m4�������c�\1�ţ�͘~��K}&����޻��=td�֖��}����cN=���싞@�;p�l�wh��"��6  d���m���w� �C�����L�*X�=I�4��#v��2<�x�C���VF��k�d���D9=��bL�������}�L�����B1J�j��*��0_q��" Ee3CvD�J(��3�֧��֎)�D���w�`�kCV5�3��ʖ\_:�����6{��(���Mb�@�c�	0�M/0n�,��!*��k)�h��PS�@�(���ݼ� l�'�?TJUD�n24�h����zՑŠO�:�h�C!��P�F�O�	)����g�O80�v�Y�#A�c?��SDϢ�~��&�����	j����h�F�Ū����@Q��/e�����	$U��w������e�%���u�j*�?J �+�����,�|ް(�+$�#%�����fOCd���0�e���q�Ʀ�^�=���_ѿ��q�'ǰ]��Q�X:%� -�<�ȸ������"�r󹮮ʱ��V�k��"�w�ަpÎ��L���Y'X˳A��i�}i���WGh�ZvqU㉫="լBu_*L��q� 7Y\+�MV�9<�_7��W�� ����3����Ï9��P5�C�,��Ѕ�o$8�o���#������_�n3ؐ�(z�Bf)<C8ݹ z�HT=�i,�%��>��Haبe�=U�zs0JG/]D�H^LI���%f��Y�V�/"�=��Is
9+C�ə�Rk�X 	+RU�UY��n��A���{vi`G��l���+���d*��d�Ļ�;�_j���D�ߗ�JD��2W歌�
��hr�~(��G[����9#�7j\)#O��AS�ul�#�8��v�[.�cX��ڂ�0���b[�̅oV#��I�*�,	c�;d���n�Փ�����n�����-���`���0�R���GQC_Y�w��[�ˋ`�G:�#�|<e��Q��̞�щ����HtRl�T�tv�U���b�rб�O0[�ML"a���$��lK�,�XPƀc��r��q����9��<�V�����Cs/�:#��F�z�]�,"�t�H#�����L�5�I��r��ϯ���GC������X�����{�!���b�.�ׯO�\j�d�,��sO,�X1�ؼ Bv|uu�v�����J�%fx�J0��Z�*.Mq�=�7&v�:jM%���}�V(E�>DC�ߟ9|z�C���%y��g�����W�Ap+2�V蟘�:�L��g����t/\ڰn�.��	��o�cpa�G�x�&S�m<��D-xv�e"�cޮ5���T��hy@Dct���BRT���U0�:3펰^$��N�׊��- ��	�����{��DpgS7����/�]d�����:�X;�eWn�bU������-��'#l�ȦZ��G,Kt��r�����LqOjjR��#(�]�(��ds�Hb���w,0��j�v�&[��q���(]W ���Ǹ'5P�XI�gThr��}uk䆳�$~��y���
��2�}~0#,R�&�
,�b�&/ }xi
"'j�2F샢oȑ��k�Z�&��#�S�Cf��)���a@�/f�e>�%턅Q��1CTZjj��:�Vk{���iG��F_��Y�`-�g���>����TAw���#r.qsy��\�K�H���ԏ\�\����L�B��A��Y������Җ/ �6�?�`��g�K�J�`c�~�ԩB�Q۱�W�8��p�c����)XW��Ш�u?�,B�T(�ؙ�Aލ�n�� ���	��$đ=�Uh�᭎誂�@�w�i��b;>�Ⱥ���w�z�7�س:�wj����g�@�?n�ߎ!������5}U�7���{�|.�����ފ��;�1��6�53~L]�� ��>>��D#�C��j�z�.*ˠN����ٝ�&0#�~��o���;"S79
�����R�`�3M�͟d�s	Ǚ����HO��;ڋ��w���돖�l�N6�o�@T)�oҶ�,Z��d�wOV��K"-�ob��z�2��s?=�˛L�	��m���]j���<e�s����`Q�x�Iz���Ϣ��ʍr�A�Dh�+�jJ�v�+	���}:��<���Z�{;�$x�63)˂h��r�c�[��Y>�cf�jʹ}+p�6��қ�c4x������|U*���=�6U����h`<�L$J�ʫ�&x�\���!:g��$��/_�����6��ZǞͶ�u���R�
�N�]��/�1���t�؂��*=wDhtƍXw�����Yh�'�w���VHذcHr���{���e0�A�!�������l_?��XU�FNc�Px��B�}+ɛq����}̗i���FyA��q%I�L"���6��_!��7R�0^z9�#�Z�$�$��0SSQm���z�ƞ����e�҇K�!7�fr�'�Q�z'����S�po-�;��H��?9Q���`�B`�`��j`��lgK��~#Ljvw���]8m���8e>���PX������jW:%��;eܒ��{���V��DS/bޔ
��P�.�1���$��DH�l���e	�����R��sHR� 6�sgY��a*v�%�@�%nW\2�?F��᥋Ya]�N�S�|J��P�b�5a\�z>�[�@����t���ك��0j���?�T妜��y�ׅ ���TIU詚�H���;�[�+�����n�LE�S��Y��FQe�����U�x:�"��Ө��7
����J�A��P�*e}S:�f~8��[��&v�~����$�%�^) �0�͢ɡ���l�7�y�;��KNZkn�A|"!fuY
vh���Ri� �ooQNb�9 ���?[�"���@^1L����x� ��8J��nN��ˤ�H7u��=�/y�Hy%Jo���F�G����Mw?xy�H�k��0q�=*
-6��[~P�6���R��C�￲=h��5�oԻ���*@�%О�i١�oH�G"o��z2r��Y���|�*��L?b� ���B�1�8��d/�������aU%d? �G�f�1�z���O��ko�j�.�o O�e'�F��G^*��$�WL��(�! >b�S�o�۵=�0��7ߓ�K&����'%�g���eO"�-��u�Ȓ��ct`���8�L�x/�6w�����n.>r��~"%(L(��VW�3��
���~Ԡ�[nL�eܳ#L��դ~���{��9���*�f�Zyo�Z\�ʆ��H�{��m��z�Ƨe�ֿ���3���2�g�K�v�l�m���
H0�ɡ�M� �
�	�+DJ���5��-ʼ�w�OQ�Հ�q`[Xo("��a|<6�#KI��+���U3��Q�d6�N�>��/N�L#��e�G�eT#�{�H2_^��h^�7��]�M��?)��xI�|�g�˂�Gb|4�� {{9��B]�o" ��6L*7_3��fy�B��#��{�(5n�U��R�P�ɸ���1Q��I2�t1JN�r�c
�Ԧ���-_Qv�z ,�hmbh��.��)�4"���ѐ1�tj���>h�ld)�\Y�
1��DLi؂X���+$  ����	l���~E���	�p����' ��������{�ۧdp�fX���Q�����V�_eN��w�#�`�l2����yْ+֩���Y���jPqY�^֕ڰ~y���p�=J�)&�^���BV�p�?���(��T�m ��`�׻�M*8��*��n1>#�z��h�� �!�?�ߵ��D��s�{�e��ᎉ4��	 ��*��E$�k�)������Io�pd���Ѹt�фC�#�u�N��ӹy�J���i�兌�c�1�Ϟt�C[�0���ū��n���3<��x�i+jyU#$\� B��L�x�tO��u��v�f�^K}MO]k�(�U���<p��1�0H� .38�%�n����@���֙�cATPR�7p�"�� �;\B��]IPԬ��-����,�b�]�5´4`pg�
�b�Kt5�Z$�Dg��k�S.wZ�q����΃�=�}� ��,���E�$0�P$��F��J�u�F�ϭ�&�Z
�⢬{#j�CbX~`91:�`~-,�� C�7��[����#u�̭��$h�bf��l�9y�-�q���I�b\�+��赾��Ȃc���}'�uip%�U]ܖ�g�.d�#"���"�x��=�0�1qzq3�����%�Vg yo��Mr�6�n�Ÿn���We�{��d~s��N[F�N�ԝ{۔���s�%���˵ʋT |���"?L߽T5X��e��l�v���4i-e��=P���U}Tl�q��o�ؔ�w��'��lA��zS���!��=��L��3ӥd�MAx������NCS�X�I��vhy�Z����Am%�?�����7C$؅���p&%�{�jOccݸ �{
s9��2�Nvԫe�����ES����,m+�tX4xQP�]���\:�a]��J�9�7ɽ�Z��A��������O��Gl����'�sn��bٴ�n�\��}a�A��p�M%��U�He��I��+:Hs�^�^Q��MQ���_����ԅ����`��G�e�L���O	�mٳ�;]*�OK��3B.��1��l�d��U��b�b��W��o���D�穽±��E
h^U���P-~7�\����n&��L�U� ��f�s�3����Ʊ�[V&�B�hq^
�;il?��^�����)�� :���m����Q}�I��������=����i]��[�� �6Bvb�3�Jʵp�[�b�VC>�|����1M$D��=����#�}�)�v�ՒG�6���w���X�W[�<`��	���5��\��G�S�v��Hb����c��՟b7��	��ٶ��h_����Ko{��}qS1:2�[.�L���k�g��,��x	��i����'�6���ZPBMG���(��'x�~zf�X������:
�3H��u���`��<��=1�哌!}�}�Ri�MK���a��Y쭀ptZ������(������Y�e|�g��OUG����R�)���u�߁��WVOl� ��!���A+aX�qWO1���pJ�����:E�ph ������'��_Dp�"�������qR9���)�9i��=�~=Ռ�Ӣ`��e1[�By��qA5Ǜg�"��vdV��ZF����D#J�mr���ˉ��F��v+7�o#�%Hren��<Rq���Ÿ�8 �L�7��$sl�V>��zG����!4��=�U���O]�����֧49m�p;�M�u�����k�c38L69�����ik�V�:�ǅ�V���>sȉ�ce\^W/�l\^��I��[�Er���B����� =vt@c	O��f���`��["���H�����D�7˺Nvt`��fχ�J��?� 5�E�5�e���7ˬ20�G�=uv�r�5�B���J�C[�mk	��UeV"'��EE�����1q�7�s��:7��Nh�@p{����	��'tf��.=��	μ���c³n��Mf��s݅���o��&�����Yi��~�.��~��O�'�|\��Uza�?X�Xr���Q3��24\�X夘��f��r<�_ͩ��u8��Y�#镉�k�H��^�U�{2�db�n	���NA�8�����Q��^���鴂��J��p��p�,C�5Ri�b~�6nA��޵8r2ջl������b�L����uq�X�;����n��Y���7ȄC�]��k}\=_db�����E!gS�)�G���9�CR������l*?z���6�]L}W�����팑�^�h�ٓ�����􄛖�N��%�s2�ВI�Ө����`�mMxρ��:	#~��u=��?>YWq#�؎�����H�co��M�´s	e�A�d�n#��i?'�O=�0�V���+t#M�Z�Uկ�����2�� $�AI�#-�{̳	���*��Ӱ���Nz�%{��j�;*v��~_�^ X�BF�4GF(MG��%��	�@��Lb7<^*���Q����ǻ��z"P��#�!<&!���0֤�C_�"��	�`�](���?���,)�r�M	��e��ؗH3D�y��؝�svkx�V/0��u���<��������]CG����b6,n�T���e�û���t�?�� �gWoH�M�rt�8U�dȯ ْ�Ϫ�e���MK	�#���6#�V�f�-�Qv�e�R�6��\�}m}��8���'1T���m�{5��G�:��7w�/�d�����Lr�t���:Į�t�Mѯ)���EOp�Btt�Hb2�w�\�r�$Og���Y�_�~630	%!��,�pj��mw؍�l���՚jX��y�m��"�Ƹy:8:YJ'!�v^g�4r��d�VAs���`X���w�y���Z�a��'��ʌ����������m�g5?�wz���OX�2�q���͇U�(-���E9B��͛姭 �Q��U�x���#�G�����y��R�+c����}�Z;�D⨚�3�D�-qH
T�B7�Ա;���PtH�7��*�og���O�^=�y/�K6��C��X$�@�Jj��2�.u?����0wo0�w�m�e6P��N�4ȱwݷ�y�u�s`����q<�v���z�w�sL>s@�����
H�� ���;&0iˇ����7@�[B�)Ė�Px��k>a,^��	��ּ�ON.5���L��!}��w���N�p[3E}}*�u#�r�qBf5vĂH�_(�á�f�]���U�Dk �3	H#rt��=_$�G��ބ0^������Z��ZK�JN���F���y�3i7��"�ΘP�jD%�w�0��.&j�M������4�׳K}���7q��?A��5	w�r���缪1	�N\[�t|;�fv">��ܛx#�Dafi��8d� �}ɡ�)+x�~NU@-���Ձת��C1_�kj�-C�D�������`�Qg�����}s\�����p]����	�h�e��j�����D�C�ND��q��BX�o���r�I|7��ǕK<�$���l(#��)�&*�yu\p���h�6�2��S%�?X���9�a�No&}BU�����c.���pV�0�n��.�����Ь�Xb�{���:ҍ�R�x�3=A5�%��~�̾�$/�wXc%�����a~.Si��)�g&p���6�fL���`�sc.�^T���C��m�)�k�3���=)aP����hU��<, У���'�[��8J�q��0���
'c���s��|9PUl$��57'-|�P�N�f�4$W�0?�k!B<���Zp�eA'�fպ-�� ��\35D��J�Ƌۨl���tVW��#� !ڛk�"e�+»}	r�X�L����\�J$�!CC��}��i��Q�e�ʨ�ٓq'{%�ɴ�H)%$S"���$��EM"���m��������O�d�L2�|h*<�\y&̥��-:�,S����Z���X�,�OZ�y�N �$�t"y�\MTU���w^�m�����e~D ������)x�����%�'nVTCWӰ�U�(���\�l
�p�Aռ��6��_`�Ow����(�]�bscAeO_yon�ח����[�� �⫵|*;Z��m?��{FZ��˦�R`�u��ai��$�B�k?�*¼�wt��G��&��[W�/"Y.vұR/��R��������0�u�.4u6���,�ت�Yb�a[+�R�H�xY��#�,�rQ�M��}�2�g��a������F��=V�o�at�p��M@�6���gkR�hɲ&�aN
��~�w�QOI�[-�����}��,ÈP�����fr;�J�HR�����|Z��b�>��jTt�ǭ	��~�O�ub4�Y�(l��P��=�푠1��^��쐨D�00��j$�:�>�@G�J)����;.���go�^˩jHa�Ho��*\�Ʃ�c����;lX����g���'��6U�9*)�r�
<�f�5��&G[+�D/  ����0 �US�"GG���ʞVj����a��^ M�&$C����ʖ)��� +��%d�aO 7@�Y6��ju�Uh�	����L�c�.�	@�貙�G�-�P�g�	���r����@1+��|.n��������a���Mst	i�U�9o�O�u�[>��ZV�juf<٪P�M5<P}b�g~��7��;
��{�q�>�Y��d�~!T<��5=2@��L�����;�X�jʛp��|�B��H�O�. @l@+l��|�,��"~��Zw�����/a�:"��[m��$��M��] ��A�GS���Q^�̔��m�B7�Z��C���������ª�\�Y�gj<�K����%(������"�3*���%��t�ϗ� ��)(��,� �q2ܞ�ȡ�2�� ���x著#!�_���v�(tkj5s�RP�����uuRc�rx�D)!�Ro	`CvQpk��c�0mV.�����%t���.�o��	f&��2�B>�ތJ���(
��͐�9�,LN;�*�r�޵�=i.M���a\��l���W�@��7N�Vߢ�m�7��Hl_�A1<��K���פ���� �ȸ�}fCf�q�� ʩF��c@6���q�%�D}����c6@�%T�DT"�V�2%r�vz�����cD���f ~��@r����0�����N���rƢ�R8��J�,Z$���S�_yq��L��G��!E���w%u���;� &�Y��hć�H�y�(V�B5..�{�q`�)�#;��ڞ�a���_��C���8���<�E,���v��~NDYUˢ����G���#�J5��ʄ���{�,��G�j��BsKe)�K_���m��~T��m?�������&)�jn����D��k_'ewqao|�zʷ�ŉ2t��\�ٓWrU2��p�}��Lʵ�#4��������_�8e`�x��t�?��m��K:]uDD��q�]Kք����U�җX����)]*�l:ؙD��
�Џ�8����7�kTEnH�ؽ5����r��*����;o ���>��ē1��=�9��f� b� >��p4d�R��kg��T�<�랶(�4�G��h`iاcO����������`�#�@s�0^_>�4�z�;HOE�n�)�2�j������[��χNܛ���I��J�L]ĭH�_����(R(��C�ԟ���@Ip�_���:S0ͷ�RQ�+��7 CZ�J 4U�!�0�7[���o�/^[�R�䠖����@�-�ڮTب���$|���CDR��3a��i����f��@ ��=k����ԧ&�+a*����(�N\}�߉�u*��j��R�y�9�M,��K���1@�p��=�*u���m:)��j�?�Bt�g"����ɋ^2����f:���ʫK^E����Խ�K�8y�O?��d1��,��G�=ZNW�v�C��~�z�
c�^{/��D��c���!r�`��B�;���T
 4;Pmz�c>���ˎ�\vދd4���Ж	Q�vt��(�+g����Y��_n�tH\T}�U\���[�$�깹 }C��"�d_��GO��u^�sN���ZUȱ����'�;���Wnՠ��&A�Zqx��0�jgb�m����B�j�r�

�}����N��NӇG*��x�kU��K�K��s��:?5jx� t'r}�L&Z8S�"ݠ&ާp/��:���~���s�ڹ��A1w�G�HA��ޫ���W�d����������[$��D�z�J�H�緙���~�f`�Y"�����m�ݼ��G�,8�۴���58�Ǌa��7��^�r�J�0l���Y�!�XO����[�E�Vy/�~�'���_l���ո�C/uI$�ybQ݁_��T�)��25O4h�tx���Lo;��m�L�&��!��Wġ�G���=�|�o���5�Yhߤ���K�m6��V�D�ԕ+Y#�GN3�����H~e�!xN����=1�kZ�T��,�F�wS�f�3c6uH�v�	)uۈ��%ar�'X���b�7s;U��<n�[�r)16%N���:��E�g�_�[<�Q嵖��0�"��ED�\uD[jbi�\~[r��M� ����x�fP(_�1`S���M���h�zIp�.�#ح���~߉6�~�1b���V"�<�!��7\��[�!�l�n+�u��vi� ��f�����uu��������#�f~$k7u� ���(�������b��1 �k�ׄ8oW��<=�{���c�r��3�]i�Е}���(P����駤��=�~����
e��R�,̆z����P�t00��Vü��K�f��u�,M�r�F�Rwt�f_U�(]v��-��F��.Rw��21��n�}����p谀���N�2D0k&�� ����.���Ǿ��6b�׏�G9%lۡJ��(~X�}��]�(�H�y?�Ǖɹ"R�3�����{IW��mc�u�L������ma�m�Y��uʢ$��Q��Y'��|�����!2h�w�ܹzi�rK��mZ;�� ����@>�������VӪ-��J�]n�I�2��N�P��C�0$����� %mu��"�yʭ@�9��W?��e��{���(r5�>��9z���j	!rп��p�Ev+8�v�9�同�������C����V��9�������4�K�Y���Ш%Xč�t��䆣�����`��d^�<�\����\(�����|�A{27p�o�cj�Z������h�X�]��Z>� ���P8�M�c�����$�c���}����;�i�D<��*�='^���&O��r��ɠ$kx����d�_�����!����7���ÜB޿��-�JP�%pzB��>]�b�񿃒���L��$����N5�d�M��5��p�m�꯱�����E����Y�������6���s�1FIWLI�-9�Ew)�c	b�zux�VV�)�sT<��Ps�Ud���8�R����Q<Sr��s�wZ��S�j�T�Fΐ����d|�U~u]]$���$jU� �*�9�Ҡ�TK�lQ�'8�\x��Z�D<ؘ�:��l��J��DK�xQd��&Ć��}�@ �$j����5o��Qk��l���>�B��^�K�J+g�K��a��ӬHQ�w�����TR���kC�y7o�N���s����R4veޅC$* e�}^*2?̡��p�g	�q$����T�Ĩ�c�c�?�ѓ�c��n��xg�p��NaoS�Z��%�:7fp��MH���3�&�FO�8�ߎs,��mY'Y��a�k{-3�nN�%v���Am�}{���hU2c��t�Ԯ'uUt
�ëù��g����ӡ���G�,�<?�Y�#lKl9
-œ롲)8#Qͱ�a³!.RL=���������JJ�����G���S���[�g�nω�d������h�l_���8��4�X��%.���U@���	5YF>����#l�-ȷ
_��j�b�}d��9�<�v\!�(��IiHJ���}���dq�Cʎ������(�#��!Qf��o�tJ��'L��Ғ}Ob.��B���ƪ~Y5�f}��N��M�r�X��)�V����~���vNgo�9���,zXf�x� |�j�5���Բ����.� *���:$��D��rIčI���xa=p�z𷋺A;?�!�Ea��YT������SD��އ�x���<w�#<���|n�3Ӆ�ji�,#J�>^1N�-N���W��1RsܶO9�z���J�$����(z�+��(C�6ڊ��M�����4;&��`��|���b��^}q4ˏn67|P�j	�3L���:��!�bW_ƚ��s�0��G����H�|���y��f!�ֺ�+.�"��;�Ǩ+8C�+�1����:]:�8c��W�A�f�N�����t�*'�L����3����n�ю䣕����xƓ��'��c�M��R���D�������J�m�'����>5�0�u>d
1��bA��#U���<ﲼ]au; g�[ք��űL�d��hн˲���U�%���2B ��ȩϗz!5}�����;�~�x�W�3�+~ht2�o������+� ���ã�r��b�@��K�ǰ��sG*jUhx����\|S�����*z�g4		W뇴'�]�͍��3V�O�T�_$n��#̱+hI�]�XT������0KS^3TPM�fq]�&j$��]�t9���h�V�g@j��N�C�Ҷ�x?����z��[���Xo%��N�U����(tN!����rL,��?��V��<d,�og�y��=m�B
l�#�r�bs�ܞ��O��L:���H^Q&��;A�-��Q�#��a�E.���\j���#p�	� <-���fj�Y�V"gpH��;~v�ug��[YW��3D8��F��ѯ4j��2V�+���L��8��))�IC��r7����@\�LuT��M�%M`��0f���&�U�U�{�)����c@We70��S�¬��ؕ���U���3G�63��tny���	g�C�y�׽��ȋ���O�O)�Ϫ�"�8R����f-Gwا�o���������3��׏���yntM4��؉��b���)З�"�|"u���g��`k$<�޺�ƆI�]�~����}���m��%j&�ƛ����ñQ�\Dt[*���z�K���p��W��,/]+��"�(��p�T&I����4���9a*`kx)0����g3q�@:���j��e����@U���-3Iaǂ����p'M�Uەzރ�!���hc���V!1/��bK������׆��"ˈ*�B�4H�ꕕ�PF$�_z"��jF�v!m��@����f������*r��l,�
^�?J��N������d�IGY��� ��K��3�ڡ�1�I�5kI^�����81������F]�+�t�2�WO\L���HvgL��4g��m#��wnF����q���`��U9e�[R��X[��!w��RI��Ŷ��q��&x����LlS[Ŕ:��Z`�T���t�F#� �>��4��z;���X����"�,�ѭj�9.����)�qɩ�7"K����V����ث�5mιX��Yw�SF�tFU�b o��� �d�Ӵ�m�hB%iL�t�zܲJV�����ݙ�UvA~}�;.��bV��Ĕ(�>5+���p��0;[i�]��%_Be$�¨�X���M�@��ER5 �L#�6������y�k�T�l˄Dͣ�{ P>qH��~.r��V^EJ���X`�ڪT����B��A�Q��HO��M�@#�񞀫X3�!눠�~�g��·�q*^�tU�Ѵ��AɃ�&���F�:~��0�z���˓}No�[[�9�%�r5f� P���QI�*��ܩ$	_�1��.w�cX��V�������e�#���rQG��}�P:`�5�wa����;�����q%{<݇0L�#�E�oi�ͤ��v; ��;�UЎ�9{�'X�2����H���:hx��uG�DU�T�YȴĪq��+������.Ф;�Β�o��y& 0p�d��Իi|���sK���ƹ��
��#��Ud�C=���#��~��ur]p����?gI����V�GJ?�}"�=�E_J�����I|#�+ͨ�#q ��-_m�n�9�+tЩn/Sx@��5��l��l]Z!�BSj���M{�sX�մ��\ i\�P!���a/��^#�)�mpu��F�;Z�h�ǹ��NTΏPg+��gߦ��0���dc������a���3/�� �6�]8Wyy`]��'���S�7�`r��p2��D��=z>o;�
|k�ܥ������Ʒ
�)�s��#��C|3{��W�1��[����PP3T
I1�q��r<mМ������Ψ^6�S��� =衹Ț�� q���:��k����Kq.�N�ˇ? K'F��T��JS$�+�}�ڞQ$��y]��N�\w�xN~7{e��4[�FT+Hoy"�2Uf�F��J!AƇ)tn�@]�3���qDb�oѯ���*��6)��J@5ұVS3�a�uh�j�F����t��X����-�6cQG�K� d�
������4������æ,�2�?�88��i^	9�r�S1�a�oҭ&y9�"a�X��R�o�h���#�,Y����5�� R�����s��u�@�.���fD*-��)֫c�Ы�wcT,�ph^T��zՏ\�.�V�(@�\�H�np`L��D��ʗ�#t�f/ij>l)��l�-q����-����O"V�$���#C�.Qb yS�+y�C�k��0�aՔQ�l��2$he#Á���x��v��]ۨ�q�/�b��o�2`0(S\�������9�;B�^2��16v�^y�?�?��/�s p�gy�p�i�:�YJ�>2��X:	�n�\8��}����(8��L�r�m`�џ��nŚ���!��=����XO��?�9V�6?>P�z)���r�6�Ie�d �@P�N?���4�j0UN.���y�~I����#�a)N��r�sIs���UbqX���Z{B�,����o;7P�#��RSYU�W�Ĳ�A����Z�ɶ��[�5����Y����zsa'M���πFb�tz��(�/��޿�	Z� �������$�L�|��5sW�-~u�O�hF�~��~pb�]#(��Zirv�z�-bl˜�k����4����Pv|����+ᡬĦ�j���I4�ȝ֬wޯ_<Q�¯+�}:6Ѳ����zw<v�����wf��@����ÛC�p�ai<�l���AKc#��$�ԧ�{��y �P�Vb8���nż�C�P�h4���7�-m��!����.�}�	��ǡ��m��N�r7n0*�;8µ�r�y(�'&��\�����:���꾏G��1o��� P ��
��Z�/�
��
g�M߀3;�R�����X@�☎a�$�$UXS�>~���M�!�Cfg,&��vHϰ�乳$�%�C�n�>q��+]U�0gѨ�jf�z�t�<��ּ{�5��ּ�"?˹kR�N�ׄfdku�/ʏ�/o����̳K�`����.����cpq0���(]����֓+�g��lk�!� �;���ަ�o�Vg���ϱ�˄�F�6�Y"�o�3&*����Y��q�)�伦�ލ����}p���le�18�VD�٫ ��b���c�7�ea�R�i�F�9<�(�u���y3E\��Cbk9ݻrz�w��w� ��3�<���;���>-�e�ĝp�(��	2k�2Ώ��x8��>[���b�?��ӥ#d���8�����i(���:5�*rF.sFV�6��4�ݫ�c{>�T�7���Q��`2�w��q�Ud8��«ﯹ���:��7<��t�<5�e��O�w�u}��p믙� a�dc�2��v�!���[��x��o�n�{A�Y�}a����	�ݳ����=�|�.X>����������Z�n�xn�L�`\>���v�pZR�Nӕ�aY{W�b�T+;�����o������lU�/�.���}��6�N�9K��=}���+A�ȃ�[�(Wµ;®���/`>	Fz����;��@���"�Go��{T˙���ƙu"�섋��IL�mK��4_N�׷�H��?�L
�e�g�W�!��Z.-���`r@���H'��B��Fy��Ŵ��<�$D; �R'��>8$7���|�s����fة�
�����:�U0�X\9�������^��/R+muo�Q��yB�EyY��k�2��E��!�$	����p`oG�O��U4q���/�A2ɝ������& 7Z�%M���ᏠI�'������8��0��@-�;Zv��snී��J�;<L^<N@�]��#��9*�AM�ײ�0�U��+l�}F��M�-���Ng*�q
��1�.��� �8϶��s2���]b�t����Y����g���2�'�VH�i�Z�҉ջ�����);��6Oֈ���,Q9ԕ�ml�/b�t ��I_�P����b&���K[����eE�6i
9�ի{tD1�ra���>Y�Z��?n1-d@;�5;��;� �WS��JǨUc��<]��i�������i�	݅��IH>}���Y|K172���M�P��T**9*�, xj�,iy j��s�t(��6QZED	�]Э�Ff�O�uZ��o�u�!�f���eR z����G�K��s^H`vEލ:�P��ts7U�� ���~����[W���}�� �W)H��*7��fp'|~Br5Ӽu��Ώ0mw�T�4�.�D�^�]j	�O 1�W�Y[Z��E�`7�����s�K�����%4t��M�_1�h��)�Wְw�f4��ǯ4@���q�q��PU�
v���*f"�0h���r�Q�M-˭�����5���n�Ys�����jٰWOr>y6���p�����_����И/�Gy>�<�ϕOʲ��׷�>4������lyXP��M�B������0C�⹋g��x�,ͩ~��nKvЫh���QV��T����cG�D�� ��狑��J�k�ςTtZ�U�8<9�+�^�w76���M��z���hܞ��'�{�;��-�q	3����,ƫ k��|%�?-g� 9E�b�f��g�1�|�����2���L/v;�p��9������H���h9�(��fR~m�ux�6��Ç&�
e'2�)׹t�!y���&���؎�5����h����ǻt(�V�@�%�5��W�Ϥ_'{A�g��Y=Ĝ�q�l�}�r���E�[��p���K�"L"�?���V�_���:"�/�`���mN"뭆P�?�ظ�܀��,���� Ѹ�,/����֙��S����@�(?6��ִ�eч`d�S��8a=������X�AT���#���Uvt4�`�OB=<�6�U_�_�34���"|�Z�3�E��e��sCRc��mP��#��#�������w�nx����NV�.�: ��gO4iH����V�X������j��20h���u8��l����G�f"���u=4X�<����K�{b�뿣��b�.o��ҙ��J3ٍݞj9���<n��?/Ф_`}f�h�-EW��P��g)�Bsp�Ą㫭B=���t#a��*�3�g]��� ��<��˪R{�a�:�[����S�=o} �i۠��jӖҠ�*&r�sZ�[�����!�b'����(�g,~����Q�(�����W�{�-g����X8TlS�J�q��A�'�߮�c���RJ�Z�Gl�(C�����O�QPg�
���i/�A��x�lЎ�1$U|K��8'�Nƈ����r���C%�)WD]ۼ�����ª����P��P=��
 ��cW�b��i�f��^Y��b��Gd�����c=!���g[WQmMv	��[�����t;�G�l8��&�/���D���F���	�g��6N$l����ց.+B=xv�o��ZwT0I;�+bR�U���[ �e��,�%��	58'�s�Ӻ�@^פ5-y*T'��]e�@z1��������{0�;/<�)�ȃ1w�&��msH<���I?Z�λ����@�ȝ��c���������¬��`��5��`
Ƒ���Kc.;f�9$�7�yقz A�p{8���H��9׼ /Sie�g�[T.CȻ�b����:�{�	�Q��*�U���\}�������8�l�{k�����ztG�c(�9�'�2\�n���l�f����(�Cw������^~�>�z�I�H��(��eeIx�ө�r����䣄���#�y��;u��6��ik�;�r?ڧ��?�Q