-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RGkI6OGJg09ydt/BhEem6FEldffs1PH7xerww29qp1Zyjp1v6wcdMnXyxCHVnWoKi4MZDxe0hgGd
UCsEfmj1Szhwmu27++ik3lEh+h/9vEg+4hQubIChhIC9JgYeR7ES5HTplHxT7qy6uZ3GOMlO+Upg
Ua3MjzZeLI7TNIZ4DdgK8F8/aenWu8kzBdkpUW1NzbMJdRMSURQBMKF8QKowsCpvwFINaUTj3zSa
XIp9oyZWGJear1WKpyOLmQ7SyTojDDxaRMTKdWY0aeYqusGG6R43OqP84SdTUlwcwG/XeM1Rk/Kz
LWGpTBgFDHx3t2Yy/ZYzErgmYYE+tA+uqi2Urw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11952)
`protect data_block
hJvlCpOPqs9cAU9B9ooQsRFBd6cLI6LJZHvd39CPGiCLseGwLc88NrhpH67A3qgoxZ+zxUyVYERX
ADGAGsJx8h5+3TrVeHirOV34H95U3UWVyU5n/Yniw8T64XpuNrC8lX3kk4HTgBJr7WUFy2G0OuPT
H6u4GkIB8APrmnM4a+nOFA5wzk+liSAwsBCSJ0/gjJj5Qd1o1a2+Mz/p5UUFr0TheLmbLnTpp01z
FOchhfN4JSN1At8lHV2gzAhKmhJPes1bf/BZ0jHQZQLIwUz8uz0wlZkiKEId2RBtt5/owDwLsVAz
X64ZiVnqoS4ThP7j2T8P0Qf0Y1xu/Ma/4GXz6cMIgD302bYeiSWDzfvdD42iOTfnyJkCDdchWffP
5g5f7mrnp5t/p4ztXq6A+4pQv4Shog+30Pljf6dUCE6GoLVGRauPE27+MvCXppKXu8bxsnhvL1UZ
DssEFw+J3E0dJDqhqYJDfLzVdz0PZ2iyRsjM3+z1z6nqCNlDbnNABazOaEPj3Dmp31+/Xbdnah4K
Gc1Q5Ncz9X0un1AKeNvRnDpZqBDv9asrW0tgbDSgxO/1ycR/dHJv5E6EdhaXyIU8kZhFft/LTIsH
dftY6ytRMrPhHYWTyo1Ccl8imhqVkmNYOMIY0n7rVrNbt4G2gcS7X5Iu2/hT7FoQWD/u02Q9fkq8
yCQEIL22rre1Q9MKvkJuQB9xS9UzeI5OznuGUg6juHv5HZ1v66w+yYhyQJPNkYBCIr2uCeqFCItO
MchsX8Cj6o0qO6faI3kdQKpbK0HgPFzQFYTnqF1exRsvs8chqDhvYPP5W5nJZnvUrdq7EP7FyEbq
QqpbBdb0/IkL4vYWBfXhJ++b8CZdIK66R32NhTIQ9RJQ0kfrsVV5EiR+J8Dzcd3P6vkwUM0d5oVd
Zbfoea+oofmXpNv9UcZRA9/+MBoA+o8fHFcvoi1FNzBh1U3QiD7nGkklby/Pdg/oO2QasNQrokov
C4LX7iYhTVCXggN0LCydlkRGjvppd6r1WqmXZMXuZrw6fPEbh/BO2us/+wnJDHO0twDkOkTieWuQ
V2llJ5nkjkcvdydMyVQWEFyA+GPDsVddXnZi9ivKrGVZFZFhBtk5EgogqiSNXh3x6gmlWzxtd+zH
Cnj+YyOnW3vYIAF6uvXszggWUkKmvi6OOEljXyT9OmLNytJ/d4uQGHy5FtE1NjMBwtNkuyaSlLgS
j/wapNUmijs8eNnlDGAr+Ua0qZJ1SnSJKFyKnLSzSzttQ0XnckPKnRi4nVGIW999OtI00yiXsgaY
xcKDiQGCJuxRneLUhgLLj+WnnjjjwP3oZx7AujI2FT7B9SyDMec5DO9TPLzAypLR7IU7GO275pnT
e5Lq77NmNyFW7o3n2bYnRvQle5+FYPeG+Q7ranNvAeyk7jQtKr0xaXeZtznZxx/LhU6kGrA0NnUH
SpgkuOL7B+T3z3DqYeHBdi8ivHUpVGA5HdNGKz+qh7/sywIHXnGubV49gnGwXZFn58g8oE1PUvj2
jXm4OeBVBCHvt2hbMYtV32IucWt5ZMbS5zf6KEnPqOMuLeDNoXzeestaIKJpSRiH9f+qFF1W7L+r
bEYFzU5KPNH1DpS+2NBiR431fK9mhpQBr44mniepaFX1dP/nOD+t9BFrEFImAeAs1qKHPB0kFzUa
+Xwj2IjuCchbJ4cbIiQLQWZJQT0cqwhnqm0ZM/fG6Dib4CSFialOrWd5SgQiWQYvCiZDT+QTKBqc
1mCGdtWV+palIVBYZUcCEHuJrCTrjUyBJtxfblmNT0BI3C/GNIC8D+VDEHFDWbFaKxFkdJDgCFaV
EsEt1C55aMUBkKDAbheI6LqkYlViO3/hsPrSfoIYvMj/YdO588U2qV0fVg+yBbcnki+V7Wi5PLCa
qAVvygqfp5kKAz82fv1KM5gFfBkyxtgTuL9cQ0mm74UgwVgpRcWBlxJ0Ifr3nk5tM64sOBw+M9GM
hfVCgKUv+9Xn9v6Z3XfOIcKHCVgfmF7sBI0jiaVWsOhn4QXGpyJytbKgIe3ZOdl5vngiUgsVEQaB
MEbEa+U42GEZIecM7QAbvXOMsd5GaQRjT5t+yGkT1azJeXS7QxpErbDszlK49HlEsD1pIC1r3dc6
CXzkSqnQ8IzJAcy6qcgGjU3DoEvry9j1olv4/4On5+MJngRSdGkLwCaDoR7HassvEO4QBGXnl8sb
hfKIGQ1WXwjeZA/zDl7Go0PRh0SlA0514OziutgrY9PzF/TsRBZUT0ywjcrI7NP9sOnvkiFnqADj
QeYSeRo9KR8dMDmjLmd4b9ZbvNTcpQ+9xEuZ2UL6qXFeo4+hGSnGabH+H0Y63+pt/gRjM6d8uQvW
3B3E9WGT3f/R30nFJ/mfSgbE1XrwSukcs4f08UPIMcOWcqTNGepgPRANDvRUlmAksTbbSqP3w1Ij
2DaA8YgEascfrYe+45L/oc2zGoIhG7m6FyuL63h0GO6N1Qj0GFlqFE3rOhLXGpCvjkexlN54pQXt
MwswMiV3u/fQTuEowcEqkWpL3bcCz6ouCZrhjN3IjYh9seU0YlTZUV0pXZUv5hu14LcgY/ju5Qez
J9RCYrmkxIsqQ0mUyNKI+xNMua0Z3GeuftlOYtmsOiIJ7/OQTXQv30RIkWbYRnajh+WnB8uciXuA
z1NKW8bCr4dPGAwRJpm5nDeygvbc8UbGbDAzfEoevwbsD5yQD4Rqxj0JL5v6EduGj0IVhSFzHNTr
MzRQvPVnF++ZvkAVR03V+Q+3PojbuLR6f9+Aoy742pBBmVpdBchfjboU8O9xEKyZlVbaMyHOLZDH
QiEhjOUro06WUvLA0KGaxrfZI/Q6KJHrLaLix8QuNdrsQW/UlqbVoyCNrSznmG48bY11cDknTUr4
6Ihpjed77Sf+czCfy19KxybRa6onB7+nkzapIq4H1R7CXgHZcerYCnEBXzXHNPice6/IngPwt8iJ
Y92492bTEYik+CKTsOJeAsxzOnfwdsZpVubVVA/k+DUnAzS5tgOEJUhCEpGgbc71GxqjjNlIu+bN
PWoA07N7C7ahNXWpJNp9GNjzXuwSxop7cJJX0lPch8dK6OXob4KeA6hKKLRoPEEf6bUjyRXm812x
OCSNtRmTLxp/0ja415cC6Big5V/ad2Tv6PYrx097o2YYmK+6V1l25+UpiaSe+ZAHAsl3b0iLwQnW
sO9bhV1/pSn7SGkP8YAS3sChSdgONe1nEf9V3lXCRAFc+KxoSzqY1Kt+veZUHpt3aPE3nZICgjKv
WZBWSDRVIJJs4rra8ozk7AOwGe/ZGUviYaw9GD8UC/ig9syc2QoI72b5ZFshpIQw+p6t04VCCZPN
0+Th9KrCQra7wjYgYmKK44Xup42AYKqxOghYh4xbfvpPr0CxiEzLkX3At9rpwWTRNqaPVN+iNaWQ
l5zby2MBv9htpnNdVMM8MTxiopiAf7xbF2m+7Or2saNRosEm/8pEAKhnZgIbtcF4VhzCFlO3001r
E7JG1eHXGHrtlYMqaBShLqfUeOsZYevVBEDT03W2FN2cyegebnLDG/oLv81Kno0jdPJtuYRSV60c
DpktwdCFJ2Uc7ngzofe3naAKdG3g0qoMjJK6rCTehU86txU1z1BVOcfqrqfMTp5s7MfQ+bB9FDCp
y0oUcY380e/xF8X1vTsVKAInm9X93LvCoTigSLJ8+7ItFp86uWpuXuLO5xaoTUpqDppLlX6Ss2TK
C9Ku4+ha7jSlUlEe81TJeoh5IrnUGY0l1/LbRZISO9DkxnRHuLuBe0JFyvI5GcPPq/4WR8e8o5Kf
WJb5N6JyYfopMUrTi0TQlO+CfMW1+/g7PlChDQ59Ts1UCa3D89/MY2gPmwmklutIEKSBxC7poK+N
O9uDEVfLEMY0+zps7qeJfRzIggsvNQDwjnKNnZKt8CSadgDGonD0xvdgu/fwKhqd4XveXVrOwwg+
xZFoSkfbL/2R3UV9lfEKbZW6D8a4bKNUc8kQPyWUlOBSjZbFGbqZ8MJXATt5NjObW00OAyQXgdML
t9U+pD4/Bb/ZqeW/ksFyJkaj9YQKl+dUQNwyrmWpzPAmyUeuH7Vxff4Sk7l/yRsR2gEqvqBcneY4
lLwQr/VcsUuoF97kiKYgZ25BkWVvgsLitbvYU7M3W6KcxbOu2oUrmSzA6khFDIeqfIkxCYWftiRz
KhtmsMZOA2JJBTrKB92rXEGo3LBLzE0PK+IvKPvcIPM6Ax87DIftX1YOpmVb+Cjjvx1ykGn8kjoT
mB5vRmWZPezt5vJyjDV3NhKgofEA8elLqNFkGQPnUusBzakEFbkyfLvwc6LlVivikHd+jorVNYCa
GsiH2fCepLqEZBaKTHQdk+OJ4aLbiWwuuWsd1TjeV3tHxVGhds/sufKPtvSdymzdi1DUkFb09X0u
LUCklF8wTRVPwPh66FsODgSO/iniZQxR3eC09UDNrQSYCrM6Yen0OaadkDFMuiJkSBPZNDnZoF8Z
1lqJw/dDcfSQGbx56FbqRBmBOkPaUTdEz3gEAjlhGMAWqhSLM0CqzeCNKZKM/sF3+3T/v5Uh6drX
tE5g+pk/6D1zyG5+jXKlpbOzzBFeiCi3ydoMuUNlF3d5WlT5DV5ce0x8tdcFiwMb9Nsbt64r58cj
tUWZJnNJ/gNLz7VQksIeVjQf5iWEy2GA8s38ze/NpieB03q2m5jDPXxWY5o2RRWVd0NEu/pf0bwy
0JXaDjXuu+K6GRZyixW42eCS+AzVzrWbUS1ZqPrqvIgXQmzZj9fg6FinaNUSN0PAzawiOC3HZ5cf
hW4gjWgBn3qU/nUfUqoMmAgVNmf2L04okXtbo7IgRho73YbDSc0Jl2lhV3RRGG5g9CfRvh0efsj6
RsF2LwzCht7ZIqodrHYUM64YLdlVfUXlvJA/IuV9LY3/chffeQV3eIp+1uw6S9MLFS6rGD+7xprd
NhyIXj2dPC1ozgMsX40g2Hi1IDeM4sSKGl37ZyD/6u1AMII3FDq6RmutZmmevN8lk+Pk5VM7R32x
4Wwz54/CLBJ+YEDnzXhZXCS2EbNPflr5XnEbEw/YcWS21ZXRjMobLEyt98/5rG7VILS5pz44D2FE
ZV28LKN1vZGNjYdkeCIi9a/AQrEy02j2pwx5J5n3Fl7+Pphb47o0Smu0qSN1VjRvl87Sgblb7lqi
RQbQJmhnaLPBVUBiXMP2lBEDFtjeTLSvnzHElxfYwSLzIrvwoi8KpwodahGh8ap99tg6bxK6VO6V
PeXezIkOaRG9hv3c73/Vcm9oPl4IJsNHHf4kpP1yTqlOBP8F/usZjluOQGSQp4SoFXrWo9PyqOYf
hRouHT3TNmMOFlYC567GS1Es/1hdFBPaM0t7AkjW3bM2ZeOOBVIPbOvMR97Y0TUEV/5GWpyhqyHy
VywIYXHSebNcX2Im2obsT8ZUF7BhxBH1n9cHpU5jnRflz+g9DLsf1lnObQzI/2NAd9GFVFX5Obx4
5stauu581LJkmUMIZoCUAwF8gj1OWhdm6On/ypQAF3xcVbk+zklbSlwutk0s9pX5FdHFW9k0eDyb
dVBFyMLaNCopoz92jfIHekC9CMRvLBMLgV/l/TWWzoENqOPTZYPkWqRD6vO67p948Ox/BU9f6JbA
8CqidKB1YVN9G7uKPotDxOjlwBTCABCB4m8HLisqorLChy+NURy5uXyB2WDbUby5jcnVABrZdTCF
aTNn0PMxJX8ooPOG2qgxdUws51cxm3p0Xye54DOQWPSN1esB6NVfuvEL2cthq6TmmYJ6CMQH2puc
SUhPQsZPKEh+0hTB51DaHO1kgh+96bdB23k8KesHJXu/Dq9ZUv2Ttktnt1PDTSGQAIQyN7UKGUl2
LaAH3K3qzpmid9mHYweeqhllZpZ3IQal3JjvGDAbj3DkpcjTg+wNt3lQ86CYopiCla8qrcu24dhC
ZBodW4U8FlPtFTG8scpaw4B1AED5kbFJziQEYFPON6DwIdShdY+oyiSxonBLeZnwyiirqXwS21RG
UknHYDfW8qglxrEU8yfDWj2j/D+ydwpi6t0BzfCiZq344YRciZtnUo9m89bZeUh05zYnpDzDjI9X
IFIkr3Q+IZqF3i2J7VuaHUcfs5xycZrvFIICugvOevaTHVYzS0qEoGxw0naeTgu4oLe+j+RGDsjQ
AtOH2CuF57Fsqlla/ZMj32lKtcXtzQxRnyMyG/iSrO9IA9eMCa6nm08s6YxcxSXcszc1oI5KdWI3
0jtg+O4WkoYAgMBq25ZdZRX1ntBV84BjADDxwh9zubcK/ltszMZW4TkIiIytWpCXott/PYngLc6j
wL1ylmMzhLgI79y/gNdASAI1mvuJsIs7yi80sbFMqI3tib0fIVl+xA29+Y5ILdyE61tIloZBBC+0
8LxVFCd4JboA0cZnjR2ow5OqNgdV4WwEZy1qYA1Zd96MmDhAWgIZsAKXKsmMw6ZtK2fSG2YGSaCj
AqjnOSYtvD/zc3oeMUKfFz177y6U6o0Y1NLoWR4qO3mE24OEO6tWQAuqKtXzRt9bmcHfpOXRyDXI
g1ELH+Vg0aqQb3A0CPt42ZLLBW1/JptrSeo8lVeYt5Q3UnJLUrosP0aTagr8A1W1O3/sakuhXy7d
7F+nsiNLc+86HuEIny/F14a5tT0Qb2LQdnRxYFYqXoPzVwAV9HwvwdCT6Yzqq+tvJ1P8wCiB6X6S
43aRlW/oQlGS5nLm2E2uNmLCL4LXG3u9tDwbezim65dtkPQNMyqq5cxUR8kFFVUPEEmpLSRbsQ4F
iik8wwQoex1xB6vEnJLv/0kK5PshS3kD+Qv6mJ0YFtInAEbb+s1JShDR5vnmTmD8Q6+Prp4H+RjR
xxBWpy9fnn8DnactBGQDkfMMTmSBA2wf3PXhnJjUYp3dA93pFI9/HDxmwuvyRIGC28zgLGxLuxOC
uHL3aOGTLoWpdYNBjwAmAAOy7yDTMF9NiZT1j3AtQWRrDKEfcKU8nejY93Om7AosNcNK1H81IJfl
OIWGiLKoH/YbzsAVUYK12FpPHzExHWttbYAZXHNSJfNK0o84a33ZKQtxGVBEYz6oI72WKcuwe/xv
7eKkn1AP2nupZcKiIkWT6j6ZsX4IwxDKxLn6H7cd1mJHLrrt9vA8DX3fySl6sLWrHVX7W/TTVPbj
ZDH6KwLvdh1dD11vCwmPVKMuI76sWkPW825v8IIrj1zuZx/5c8Z/CxQiBImNy9jB3a/KTqpK0IeG
ce0qJWFX7ciSaRPtlHsY9jDd9Yy6m/UpUvfYKuyiZCl2cV3v9V41zuk9ZtMhuPBZ2c6YdOekBIqc
RBqpZqeJ8wBZfpD3kHpz71SBB012yyCadoAdV+qgF0n2uMm9Ec6LoOgEgrPMM0QTSn/JtLvxdq2H
tneSLU3xdrzNf+EqGnXd4actospLdTgBMCNUnOGpF6zsRxLTI3LCOFOtaeux54lwduOL5HpEoB+h
7LrMkBQwiknZAkBSWXUm1TT8T3mIi76F3y6aJPSs8MzICkJ0SlcNxQO2DAU00rTwb3/CX7mFBQtl
Oam3AcK7UvPqZa1O4RRalcFWHNAES/peggBby7t3O2xAjLuvYj33c2ot4OsjCgV2GCszkMypl7RD
I2e1ebJGN0aOhPIuTFIL5oGnTcf1DxuSIfQZizxwKkUa60VWl6r/cSUL+d5wLhnK0OM35QRV2hTT
+JYzls11iSPyOmZYtmG6Tk2anw3X0UQm9YmSP/Nu3OsQXHaEug5KvJQpeAC1K/l91cIqwkV+0BT+
PfQWiFV3Gtowxv9baFjHSOhM1gacstWjOD4HadIcK+50xuKpyoYk1edq55h11TGWud/kOt4boU3x
jcXR3YexaUQqNb48ia08TjGtqjW+72LIO2j0W6oHc9eo0T/LjrGALRXz3BQIeZTM8SHjWAIqgwmU
CJJBSa8kTRy5BnQZ1ud0guFFTjSLW/1qprMacZw0gkA1pzeIHrUT+5t5K8jdHCPjvteZ0FB/HByE
rf7OLL2LBkYsUhukfDy6k0fjKxVLMYBkDmG5K6dZl44Jd2KuOk0kHhQrhAnPis1k/TWXsSqmv+s4
K5MTi+pGnbIiGelo/HGarVeKoU3BW+GEGB7zRFukzW4I6XV073kAbMCbswEz0s46s38uyYEyUvDn
CjcJMCUiHyOCbXpw60fVPDyTtpQ/US1uvIE99QhgGv4kJGvUR+2E1yllLhzQ1px+uwR9CnbGe+hY
YdHd611ZpbFgNhiskefvDoYhLukP5bYdr1mCGxcsuJY6RciYUoZEcIGS1XU+vpzRsbX6oAFshnvU
9oj1bHia/cf/W5IufaXVbBotlVEkITtUr9Nf3D6YEHQOmyM6OZ0dNjOaKnXB29EjhS4rcTpB6IL4
ucN4O1xm06Rd6hWi0mo4KU3BqhryeO0GtfGi4Gd3Y9L7OM6stnott88BWPUJ0PcmG33CrkXOlV+r
I2KgM5z4SfrLQhWK5+eSjFnKokumnJVFzGngdXHqGQMlcFFSPujF6GZ4IU7we3ZY5h2tkRtu5N3B
ZZu95OqV/UaDXSv24uCOhyVIt0ETC3VgAgL41TOH9ynySTDlyIS8FRdvmOtpWQgzmSjkNcev//wT
5RijeNXDgktHXZcxurA+9v+Z6LBh1PB3xfrJCQlYlTJ3NhSe0f+Yvk7UVDqpGduXFI4UAyxRBk97
nxpqFwrETif9SzxWVC1xYZlpWzRgy0FWvpT5CoVU427W8Vuoa22stiVVIP+4zK9HHhV3gT/dTuOw
zkw5yNTywMBqU9ZkoJbMcgX0IWS0fbmd/nX/gRJCFGBDhqkaMF7RucOG4bHOgvQ8pBXWw/x3wj56
cKCQffNnfIHpojqOgeFgMhFlqLo3OHfbB8sQZau8nGiJCLaXdBYzKokLAvRtL6fq8QEgHzo4zkEm
Zk0Nil6c9Tj6If3aTC1Pc1ivJmAkdDME4FeP8TtM1drQAMniDcWQ7THMYZ1vNGrErEyMdiLkwABn
/pld2Kv7IOx9AZnWYFyNV4PseDZQrgN9ETsAgNYrxguEejhbA4jv1kM2JkhBbMhBdlNyjKaPTh2Q
IOhAT8GvekVoHhIw1U8gQukWsMZoKqL7djEA30Pj7oBTL8ANGedI2MlNG86h8aq+oSpr+phh9mlu
x69edeFy1xvyo3hrCHsuuH9PuT6dwusTiD5Xrfqdop2QyMz6Tq0linmq4pXGCEN2HNHtEE0ghkD5
ZMfejytAZvL2Z2ei7cmSf6dVFUf48w3EV9AsjrJD8Wf5NtcmuSCFbOqcgeQ8gbxBtoMD5sro7GVv
4oM6EpmPYexk4YGn5io2MoaABFXuJ+PI5bF4a2OZxTpgHO5qmm9zQa/EIX0tysmGEupZY4qfZ7NE
9QKMUZk4dNGIyChJJGAwkVTmeKKSSZJ/o25UuhbBIHGRaYUmEWl8iCIx04v2cdOWTvlbPY+lPCPM
P4h02emzr/u3hoNWpWeESIf/mtVtV1G1oxthFaPDvPZlhdAaUYQIDeBGt7oOlWT6fdLOsD3y5AOx
0rJmpR5l6yy/wrlXxO2tLoQfsPRi+6Ezj5ydA4lFTZJQbL+AQlrB6+l2Ivoa8QzgSpF46RF0+eU4
9FPR8ABcgRjOXXgNuYDmtWbcki0g5y0Jdt4yKpD3way07ak/6hiiQuT+q/IXD9fKTrl75CQNzuVS
+d4QQ7zaXtfJGGx9ngSJLMqYZ5wgNNDCyXKVtnyH7nYZSwbHSt4flTsniBEeUIdSmf5i30rA7NKa
qvgAG2rfRMQqVvP6Xld8yB5TXTzH4R8bSnXWoXRVBW/n3mnx3WTvhAw/wyqBKIeYgAr+PHF6Jggt
ywL23yZkxo6bcDoxhQt7HtgWxvtdImRuhjcG85LW6xvQH+nmcixwJ7S7Dfclh2NBQcRuBzOpEXCE
haaE7Z8ImLgINmUXZunwpFDjWBaVNi87XQR/ttwAP2EkooXIg6mJsmd2zNY25erl32GfT13cqvsO
rYsIegIFdJP6hl9u5k03SX1VjjhTZkIqMz9ThZaYK/rWlg5CMXyBgjnGAp5b32mVubqp9cuPNDw5
rA5mHq9Ag2qNbhS+fxGWleG7V6i4OYTq9pimbRUPatZBFoxAM0Isw78fPhfadLqclHSo/a2kMgu5
V7kgKym/ItBXfKggLY2FuiUwEzRjV7AY3EIBetmTVDxJu3BAoO5oulxlnwTRmFlUmPCTsHx9TpZV
dqmMuf8d2Gyp3uUhe+SlIm42RaZMGigmSkPQlvHeBb6/gfWvb45Ta8iwiwLy14oQsudtNmzkLdkZ
WoR9tfG+3KVbd5IqjH25SHcKIi7vd7JjPcF6uRHilP/ircB4tzAhBfsjduXFY9IwFVxaF6qO95Ks
M1AtY8fze6mt+gdwbyCCn4CpSrbkT/jvHNIrCcid4mFneaQ7Inx2dcxboiYozfQFwysSzrFYD7VJ
PCCQrOXXXdryFrT/vjiI2mSEegV44XM9AMiDjRsELxbM0kDdlht9xDLvHHCyGXg3xPEEKzWUHoBe
jXGbD/hWS9zi3NakPhSk8+IIjUCTNN60ZgtNHpEsf49Y45PvFz9+a/8JH4TCEBUujXfSQldsfvJO
I0sPRz5k9RcNMOS0OCBqRJ/PzkYkL5xWXD5NpG6y41X+S0FwM24Z/ZnBBoxmZu8l9nsVmm+tOSwO
eNQfvYEltNDn6+MFko/oQhftylodJya8kknTG+oVd6iP9+5aqhSCGRow1HgLOR9XhE/oIgbIWVtz
v5fwXe4ihaNUMLHpRcIUSYmPx1n4kzo0WDLTFJIsZlNZYbS8UWKXSnP0vksW/7xoU8XR++fnfr/R
XVdF/UL8Xge6PliGFkC5f3mrymWrma8amEZjlwbMVHktjO3uc4ldZTYHy6vDTMfdVRFEANdJD7JP
ikHFR4//LTqmmhBDqcaFtc/JWEfVC1LlIvcHxZkPoS3RlWCfVx6pEjmFArTPLpFC+jWWugVQjW06
Fl0njJSx5vtLAqIPAx7pxO0s7uOAuLOX1jo2aq6FThV4pHVMvVSQXoru+/sdgwOUIdbpI4FwbQSu
/9XGUdMShO88GDtQVXDs+FfitNzKYllYA6a95DGMlSjiJEj1mL5ZHO3chT2j/8vMmx24NtKfmK5z
8o/02rZBwbzbE2UrSeRcu7/ysAxXGBkRI6yrEJBZOz4oZbq2BsjFlXPgn16Hj9L8RHwOMFEoDc1G
8kaHhH2rmyrqrBh+tZtdiODGBTi2Gl6bIF12RbJaWPhPLzywQ65VZAYz87pUZVnVRwa0JnNIqD9e
mfXDSTKZnbsWlMH9ddND57MxXBSoghYRfiRpBA/WLd1MBVdV8uSpxdGvA2FfmGZmqDmGo5r+iuJo
C4zm0LRG4RyjTvgCAWp06t3dLyIGsGLhuA64Wa8rwAOfRk8MP+TzIaqoz8psHxlY/Gv4jx5kPTs2
FHgSFxAyPOIRRbBnpZouIkRSrDK9VznooCXGSW3chUpepemfBfwRb7KjxuyD+uKYYTDTrTGRwBKK
VHk7C5ov9PX63IUzj9hpoF+K4Lf1C1Xe/SZFepTSS8cWZGmPvutBLqo936fihA2OpF9Vxfw8B+a5
Y4STENmTDIM2LvK0ehg+TiGAAmb7YNAC3/tRNZdsgI/aQ52oPADlJKtzUKX5U18uluxNXzrom3p8
eGvTEvvrHGx9s31YB9ZJLUS0KjN/djCJ4a6B0K+Ap5WCE/qJilI6EjluEEEChmSk9fC/JdHbWjxo
NF6N1DzL+3JO5Dc7C9KIVMtC4BZWUsNIr4QPGnBmOrNhpA2kc68SdGT49N/FpQnkBqYqUdPLgx1Y
BY3qTHA652T4SiCLK/7Aq9ljTAu5Mv22/OCrBvzMWl139/GgjPbmVr2t/btV/BzNKtzzEcP2T61S
UvyShRN7S6M0xMAkC7WqC3Vrz1+0rtWRtPkc4egpuV8kn/1VY2kBCq1Ctm8IZqYE67dPcQBJqOis
ZRNT0QgQetHYWBbZsrL+go791HrRRrq0j47Di3uC+XtrUGQaANekVpVqqhDWjcn9B+2u4RsS/BPl
7SkoZwoTJB23ae6UesJEcVdDAp74KtIFxDiPReLmKdqjsBf/LmFBjuu7LHRTUTS5XpdjJuCmZqSB
YajLNBmIBnovN4+p8H38seNnbmNm7am2XJF1yL1/W4S1+tqNugeRWjxTralxyUmBBF53eU4DnLjF
6ZujQgR3lOtq+lDjcx312oJIfEW6MJSD8Hyz68jtUsmTpgbAKpryH1k+3EBFBjt69uQyJHSS5L7h
L5aYy0dxmneKLZdmHHiFHJP5HBiEQ7+xvIjSJ4Vc1KCjOvZeXa3q5CO1YfG/Uj0voaeDuyWwnF5A
+O199zs8BAkz6kLIFlF/Fj8cBShURiFn5zUbn9TunazOqenjWXs1c+5h/gajupNY/pxEybZ4ORYk
NdYtsWsjekUV5OndAz9B7G9NnYNh+5HIcsGKh7h0iKxm8HMWk3u5OObTj7ruYp67eMOt/1WUPrK+
OhDD9wSU4u+e7gX/NoADD1VgUXH/qYGE/zgmwFq5RYnnu5Ut/pV4cl8qzN/szq26J3w4cm+81rSS
9h5dxWxOPC6dYMmx4tTqfX3mtrNSLhfqFZcsY3Va9Y5AieaKYQVRNEOl/fiRiEr4Q1IyBwj8uo6x
kmGtuqgDDEmjePz/ub+MMcpXArZdEdlaJEgqTK25X98cWZL+s6CoW1+VYs3ZbX+bn8PAjU87QoLt
3deZfqQVi+0wOdbV76TBMJsv5N0aF3Ic2dCM8DlxKfQ2Dwg+uacRU7u6PAObotAFbKOA252VWTNx
L8PS9NIHopbIqkrU7HEezMJVR3pcZ5pLLui2NHiFp71l1/wAeU8fxZ6/fhj9jQYlZxDv017HaRdj
bbvwArRb5ybrzuc+QrrKwYhyW4YG390H3DXh+UcccuxHhBRlUGDPgh+pO2/dgYG9yWGd1aKDII92
wqfz0TtPJYC1b/ytsIad4rKYkHimK8y09IgE15DVlSpPiHQQQp2q+b4/SvYhLwEBclbkiBL+FxD0
9xJEm/lI1kMfz8tHBECI/BfZlECWLhYxHdqsVrnxAZ2+MZpBQGhQ8lIHnMAwIaFSa3Xsgf/4wf/l
kZTJplgPkq2GymWlWlr10dHTArJHTsSeX168wW78jc1G78WIsvM8x2xgje4z/Vpz0edhW/5qhuCK
4QEiglE0TsHk0xfus1xFQeIN7awEmSCIEVUTy7KdnQSYw9a9m0PodOs6dld/lrTJepDghMioxxBl
CD7FPMZcxMWV0nPqerPh/YYz6u7sh+5aHCOA2i6iTlHy/YX56zw2e6sH6obMAy/RLHROJb+fgZ+/
X6ECd/Cu1+H1dVW1NCYw/eiPu/rDwC5kqH0+4/36q3j1Wfl90E/HMiNotLmW2Wrk1NRoYLOCmp3U
S7sel+bZ3gZGWWwcQwCqgKTe2W7o0FSJSz4Dl6PrGAoCFqqKfLw86NAojWixXBo6lMJE8smVnRKG
BYFVlkSra3Q/dq9bGwkoOKBKKdqo83T5LyQ/ZmlCrBv//IYYKSSbh3gUmq/6yoY4zJPix31NV2f2
EaKtHsLBCm6zGHqtEZEf3oOoUQLkP36LgbZ0Al/d9qo/+UMNr3Xt1IM0wiV8CPXPk5LiEEBhnlP5
MIq2S30Rj9rEgKoW9Ye33Hk6Y3WggunFl0Kv8h7ACdSmx0ziwxI7e4NyJCd/0NFWtyUe/j2rgaLP
C1Xr6TtuT30MXpHXm3F4cpHVAx4rwnbvLoKApG6sub6uFDv1M/QvaeAIuJh4g+4V6m7UaPOSrolg
Q8OPv/vSrGQE6CceWYn7Wt6JFkZNG0HPzLTS47v0vALqQ9jH5XuNstClu5cvD0C2DRuGQslA8BAP
uBk18o6Q+kA2Trrsd5cvy0HABQUSxa5/k18uC8gWW8/UUck8X6OXGNicUp1iogzOiU3AMrhKxtjz
USdlGGs5wqlx3D/QSV7gZ1HiyXVt2/TGoRMIPBZTplUYdGIbibkmgqvTsyRpZad+Erwo33OeW1U3
V7etyJCjZDycKUe/n4f0f1MGHG+yNZDcgOhn2tNTaz1sRX2172Q1XckyPOJpRJlOjXMMhqr0jgOl
t6lS3rfXcjeeldgTltUj7wZRjYNo+dGY+ZLWA1koyZ3zhAYWWVA4vZtJILx7cvJg5mGZJyJawGKv
SQEEpdMAF4XCRN0AKJYbG5Yq1jH5kbEdCn33R1GvjJGzEIc5M58JiUaCFBR5ZCfCsU6OSaXuJmou
gWpYyN8lmZ/2YINEYtwLzrmk/OqwawLslwUh74n1hhjPLldRR31NOT7JDKtEUfN43i0457R9soMp
Jvtd8W2oZ9/iLhBv7Edg3uaO+D6WffRbgmtA6sPvXEJNu3VFePlJLgG0hV3lo3P8Z+c6DjnNUrX2
LP3Fg2nQhAN0NyQUf8wLSg7TPg08ODdnh6iZIMlLBV9gZQ9x4pgjkqSdp0zew7hB78u0h3fQ6zeu
sEosySz85sxae+wTV8ubWZWcSLrNuGPSslh53U3krMEHXrPMgKoRzX4jJgwZ6CaIvn+FLbiUcyDr
PFZutvJgmb+yfbqlD+cwlW2Fd39Qpx5vtg5dIp8Rgighu1KHyLmh/ddfhIU4Z7A9sU1YeXWpBqEU
oFSsACs9vuWbZ2pBjnNMp7I0Au7jSqJZPuEVKnz6ecmA9YMh2TAf5azFNHTG/Nc+HEC4s9PNDWYD
v6jt/ZkrcO8Tmz/7Wd96f7pzcr3ahqFl4F1XyW/U+3t/t8DjEHryOO8H0pEYARPNFcDXlvSkJkP1
qhUT0M2NGzza2JdzNdefKGRJKsPEvVy+G4epQlHsOBl86wGt7hDsX61PdcxsEMSS5lKCcOH+QBpF
rXNjP0UXGW0FKxe195kGMZjWw0NvIHB+OG6vL0vXO3HX/WxMz00ON2L4My+R81bZ9gtHNdQpbfRp
Q70+7yXeRM/zGBysP7kmM8MRvKPFvgXnDkh283wskHpfgZItlgSFgTi+pPilSPsachtHgO5pfarC
VX3Lg5+E8UEnH8ZgFLzPINjDHCOkm9a/a+kPw0c6WgYxNQetPIWxkrPrJMHP5tdzk2Sj6LdWWR5c
gS9Wj1rPzziHbYEFWB/SDFIDO4qAh1Fl7SjmRD4veTnwUSTcIHCMWrffBpjlS4sUznI/HNMTP26L
YVjVCaiYJs0zDRuRPOSrasJhznNTriVwhZbIXVAmtLW2dqYJEhfIsYXL7XAygFN67dcVY1aMkO6e
xtMytf8tEo8F4OKYIjLrmrmSdouE58ik4vIj2cxQYpWWkpQ/4ynOCvX4zTCJ82DQsZZV2f94rEyh
xvMpp4ml6MvWFFvFr/bjIpElyT1r+RkO+Uo3VoecEoQ2goLQ+H0RltBePvcjnXvDKkUlch33ZhbH
v9/HNzGZbEUBtwKP+UhwurabWHxUU8G3bqBGnaqxTMzmekl0K97vI2F2c18VlzujWkpWoJf1BU1R
dshIfY86g7zh+x7vA/WsnSn36OAwmyndWoGrxsxTdW9EmjXUctrtpsLFMsswI/q++ekqp+mEazTj
KPVRcu3L13Snrf1SsbWZ00s40U/0kQvnisS10cNo7G59lD5OPWeH63OrRv+hKvmuVxJ9PW1vih+o
/xDIaeYrVNzvpdM1w4QH9DnDQUuNsOOg77yHDNQS5v0RGWBnpQrYsl9Ubz/j8FRLLJjold4+w+RG
gns9SvR2nkJZ2Xx/CF7jfJVHmq3tDpfAAOtUolIIWFlHD/9W7s8bP7heoJrnYUEm3nGTGYgLGBVg
WJgEq1TpnzkxZ6o2JRCTb1Pg2IaelZMNPXxJTAyONeLEU7mbzBC7ieOlQru5uhV4RGQnYZIIZRuC
le1jQsFzcc3eS52RnPp822Lj9ZgVtIi3WyhGkgxhjlzLSEzTE4zQshKZqxZCSL3LdO+ywf3wnc+t
vhi3OKb8nCjEtP7HeGJAxFNXXZ+U/ij3MOpp/3f9+3KontKoy05j
`protect end_protected
