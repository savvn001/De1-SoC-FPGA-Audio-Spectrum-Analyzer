��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�����C�a_�h��f;�Pv�җNw"���� D����>i��CƳC+j��w�*%!U�Z��lyN���v_��Z�{T�w�¡�@����&��7re'+�b�h�J���2fV���3V�o�j�c~���V���9�!����;8R��!�6-dB�fC-�^�<gbOI�H�������G�'.���Eo}���H��v�r��:�g�27�n�����i���:ECT�h�S�|�/�#��k�������
�k�m�ɝ��JK9��Zt�/��n���O0�S��Ҋa������<��� C�-%]i�a��*���p1����?��nT���F�/��f�D���z5z�4�J�9;q�����vl�ڤ�5̀�A�t�o���^4������`��v0ST�D��;I�u�4<�/}�9���?���ϛ���d ����v��%��os���'�Cʌ��r�!��u�n� 
�(Nh�p%�WhbRj�Y�+s�[�:S����3K��1̢��T����7��;-�$'��AsQ�'w�6��4�(��`�{	5]v���ߺHd�2T8�,�]:��[ �y:.�C:���q�Kd���(����ťs�������(]�D��ר3)�+K�ӂ�F��|��i
������Q�)��o�g��%Q�I� �^K�{¸����WL�_z��I�)%s�� ��",U$��?�8��O	8�n'o�ے������͏,�L���A<M+�7�B��S��j(�7홨�P=��;��j�Q���&�3�E\��Kh4�Q$����9Ԝ
��ё�@��}x/El�%#�b�IG����b�<uɖ�� ;)l�H�_���>���'�������+�Y<2�@�܄M����ʉ���8��S��vb��O5uL^�/����ַ��+8Zr7c��Q�{��w��\��.8�y-,�4�K� Tw5����p��ѻ=w/<Ɂ�vY 2��`�7G��s��=-v��ݻ#:� mB�a ʑ�|�=A�D��o�ɒ���X�����u������2q����}Bý�@����[�*,^s���0δ�CwåQU��z0RT���7'�w~��㹵�q:���v��$��8?h����x�7����|3m�fX.�̗�,�`U�S�������T���T��or kb����㙤ڸ�0T��]-���Q��`�%�9�\�����4����w�6.��j�#?��2JQ|d,��2�_��'�ӤMR�w�Sx�Fq~�T�#<��1V��5�f�TZd�<���g肨�ѭlS-�<9
z��)g�y,浸G�<���Tڈ��*Q��LswY�/�i������d���c��0�� P���M���鋸��} �������n&-�K�F��6R!,��� C��8��\S���gr��ŧ=#��FM��G�����Ʉ��,FQ����"~���ܖ�*�ʄJP�ȗ-�_��=�QkI�Om�^j=�9��5�������d�Z^���}u�0���ߝ��Ȃ�����(�����X퀩�{�|W����[��� ��|��O`!(<rЫ}"r�G�D��u�2���c�Ĳ4�G�"��6[�}ꤧ�s����J��9�?�cd��K�Zt�S��:��*�5�!�I��xwT[iD�K0�\�&�H\&��*��B�xbqCݏ���Ş�_~�I{�4�~��:3�f(i8��K-�ň5��-�/��[�w�t�sywc#��N��џc�۴��y70��@��5A��A��g���J��a���	�2�՘1(�$9[���^�w#�8+.���([����S�aGa������~#��G�8o���TMT�W��nV�V�jhzCH��
�&Y6�h�#{���}�\?���\i����=�䤪*�\��q&����&�#�z�df��O|L��L�r�=��s3�9��#�;���I)�߰�:^��
`�'n�$å�u�?��8@��
�0 \���7��a�+�����[�o��Ю��ρ-���p�٧K: ���*f�9�5��(����D^q��rS�f3����ʖ>׌��rE$�� �q��v<��)�H�%�!)\�ƨF�dV����@���"�tۯ�ۖ���T��ț���E"*����Dޏ�U�����J$�E��+?^�L"�0�	1^�Q�hAd%��l �\���kW�"^�Ca�Y�^࿆�^���,-{�
����Gn��i�-�܍:�����}Ӵ�?d�(Ě�M;_m��b�H��c��J��g[�ȅ|Z�7@0|w�[�lbGQ���h7��ڱU�����z��:�X*�s&����.�U���̓/f�q����9'�h��Ǉ�m�j���+�p�h	���q@��>Γ�����hǳJMKl8y_���]7t�{J�fRR`�i�7�X(Uw�!�J��u����mu܅,��+�q�����G�߂g�����Gx:�s��,����'�� m�G��E,�/�B�DB������m7�&�p��JO�J~���b�)V݌�����]������N��l�3�1���J��B�pL��\�U�Q�+#�юo��~ÿ�I"�����rN_��?�С4iK�8�]��@C?��d~�b.��ٖ�kE��/�r����C�˅�p��U(��9͎��t����h�Hx0qCb�s�)Ӟ%�gl�=N\l'��8~`��.����{.�I��r�2jC#}���<���đ�y[�,�d�K���m�2�k��]�;:Y�0.I
��j��q�ϪD�!�� ��6,`oL�FZ�g��=��Ts�0'D扐D��q� �g2��;|3�Q0�Uq)7p�B	閉���ȷ�Z?fP{e���E���p3�M��c��˖'.�h���Y�W%���mN�bʭxmެ�R1�� ��#�D�'#7�&l�4��!�n�c{��ǫs��y��rFS��������\�4��"c�I��R��,��#(��b#aZH��5a�1rZQd�ͷ�D�B��c��d)�EC^9�(�l��7�#�sᐵ�~�"�����������c)�o�9~̀�C׻H�z��y-,����ѝ���7���!��gx�����>���*b*>��q]�����^�9�C����~-t���>�'�6/*��ˬearUD�G�H�r}W�=D��G��	6�%�%B�,{�uJÿQ���]vk�P��U
5��@k9	M�C{/���bE��0	��=
�-�hK9M�|�ӟ�����t� Y�4(�� Jʍ�ӗ10O���QĠ���Uk�V2`l�S�TKq�55F���xfi�v�r�6��dt���~b�ϙV:��^`	��:G$�����$�`�m��>�뭋�"�n��j���X�/"�ao�bs�L���]�$�٠?4=�PZ��I��<�셧��.��NJ�8��%c,=����7tD�	~O?#��JNx>��цf�@%�tɂ��W�}j���(՚�����7��z7�qq�xk�1%�`Gw=G��0{��ꋤ��gaLFp��1����ᆣ� �j�}ĭ�2F?�Z��e	����Y�{Z�β2قH8�\=�����6���<���X�J`�]ʒ�'=�n0u��US%��}a���l��N�B�Zi��n.�B�W���6^��7�ȘC�L`1�E�<z���U��g9��";������^��[�5|�zW)]7��!��4yD�I@��u�:fC"4�5h�Sg�uW�)uGX�B���F_�mh�����j{ �L�L|@>�'7��Kc:��W(e�r�� �O�XvLܨ��TYo�JƟ���"$х�Y����}�yI�t���v)�v���Nf/�[{�AR �n%;���p�$���-������O�	���^N:jKj �|%�ݿhJ�
�7.�6h%|LW�g�*���'�u��&tg�h�]2��m6U6%*�^T@��]�.�7I���h�"�zr�-��t�#R'2��%;��S�P?|mb�iUB5��SX�~�R�(���k�Z�(��;$\���M�A� +\����9+���>��`7�/y����~&���ɂ@ƾ���"'v��ͅ4@}1½���Ą�b���OK��Θr�Y1A$o�[L��q�PHm���4���0lT�����h��z�w��m#��!��ķdP寃[�e�L3�T�W�R0�.��NU��z��pwS�XC۔��T?����N�~�NJ/�kDsM���� ��W{��+��H��5ĸ��,Ax[�Tc9L�-�@*��50�qdΝ���:=���ca�%_��
���N�N��R!(�%���#q2WS���S��Sdӿ�ߩ��-�O>k=8/n�XyHc���Zf{�%G���)	{����7h�b����n�	Ɛ�3�#@�9WQ�;��;���}Ah�_cY�lFJ�-�:�|I&�[��z*��N�k��.��ߣb�z����Ђ*�Z���E��-���U�����7�t&��Y}�0ߨa2�9��Qpre	��%���`�L7YyH7>��������K~�,��cEr�'�~�|O-I�W��vy�	�$l�_H[^��$�T�	bt,HN��{�	J�6�H3Z���'�I���+��G���s*�:_׊��r������4ԔXXi��h�B��5�~��-F�`��Es�<��&���8�>y̘�#qع����ґr���p��m�T([�z�A������9 ��3[0c;��F�x����e �Bn�A���m1�2Ѧ]Z��rK?I��*F3|P�<}�΃�������宠ߺ���v�~m�4�Ǔ����q���ĳ�w�z�s�)��Aɥ�m�������&���#�;�����%	Pen��Y���Y�����ɓ���I?� ��kt F�a��T�-T�kM��7J���[�)��������g��0��Nz�½�R�~�\�S�\�p9<!��eH��L�7FxYk?w��}���[X^đ�bRO,�H}�K)0����(<̦n\�(!� f�Mt�$����1@˿��L�b7�d���^'�V�Nf��
�����2T$q�D�gJ��}a��ޖ���Gmav�`��	v�ڀ]
>kC	���H��=���ѝ`��ӗV�ݭB����6-��I��Ћ�]�'6i���K@o#��D�L���p�FϹ��ǚ���^�Ϊ��wq	�S5U���@(El�Fk�a��T�{�E ���2�i�ت �8��"�8�$���Ԋբg�	`�� ;]{�1�37�]�|>.�����ʮ�eEA��x� �XCV�l�}�>��</?�i�1hAW�6���Ǹ�=!��ߤ�5X6��{��#�v��(�w78�ʸW����K7�x��Y�����=q�D.��0Om�2�Y�<��s��ǝ�؄��Wgi�����ݍxg��F~�b�pRfv8�$������>;Qo�Ȇ/�`Z�$~ӐR}���:)OG�r��v�G&;6hɗe�y@lX�66�g�mJ�]���	�nr�N%�0�p������~�ȃ %a��N�%�sAa@�.<:<Q0ѱ�����ߍ:c\?�%�c^��U(��xm��ʑ�R6N�vd<[ѐv$�E���;FU�S9o�"ay��;�D�P��i��뼂����P&|�Ĳ�D�A����_������&NCT���FR�a���)�C�Os#�����85Ԟb�.-�.�G�Ur�@�nA���^������+������7�pq�b�$B�F�\��"_�ƙ��&ɰ�.:�'��4��ε�V��<M���.�3R��B���l�";��~�	@�r�c��5��������� ه�T�'ǉ�b���µtUyZ'��^�c:1��%w��qOEt\��8�IМ�,#�~�+�w��"�F�pɐ�[ͭxm��o⦠���4��DJ����x�'�7a���^�r�WF�{��o-���yRJ�R���Z�]��˗ԿO6%7��Ҧ�{����Q�<�@�찴�����[i�����z���-�E@�[?�u!`l�~X�b��d��v_���Q�S���n�,��0X�r&N�0*�H,��i1dg��wD����O�S!�_�:dS�ʀ�w��Q�P{��^�4
ˊ�.�O�1�����Ny�$�q�Y����)m�Q,�|��ޠ��/�S�� =��R>����U�w��3���r�s�����dbP��D���_�~1�JS��:8�w�5'eŞ��	�s���9��ޙK��+o��1�~{�|đ�(��Y��*1,ye�=ڴ�?���\kp-+�
  �<&����uC(��V��Ҥ⧅�*Hȹ���~�?1�\��Mޭױ�[�T3#�L-4��SP���?*䷸O��*��ۀM��%��6yY���
BEf׊!��k` U]�^[� Z[�f�?��3�nA�"��~�wZ��q?W}����DX����M�e�t�B�8y���Ru����Ju�^|�l�bt������&3��x7A��h��JgE0��,������$��p~�i��S�dS`to�$1>�al�Sy���IR�?�lde�Ow��d0�i_����K�a.�j��g��P1@#��2%K��F��g�O��'���{9:�ޖE���<[�u��E�E2��$=�d����~j��U�S�s����k�ё�k
?P��ˮ���$�"��ߖ�t��E0^swFG���(!ơ.k����%X��
���ZA��g�y�}k���@��Ñ�U�}(��*[�*X�҇q&��lE(�~	>f��3��3��#�eJdh�1�^9�| �Ң��DX�f��N��"U��#����^o�n�ٖ �(�6rcv�BaK�ɰ@��)�N���F�P�]��[���j��Ⱦ�v5�⡢���qo�:~c�e���;��n�3ּ�oyV�TM���~*�+u�D__z�Yw0�L
Q�8f2V�I���l�PZk���Z�m�
��ѳ_Ã׏.��Djw:��I�C�I��;���]�-���M�O5-!�贷1��S�Ba�����R��2ݻ>O��.�smNX�!��U.�_/-!J�7J��1	E�/D�u�*���/��~���/���;q�K�U��fN�+�V�S���K��4c�����s��+�VdH��y䋎�(��)	I�������<�:����ĕ�0ا��z�Bt��%�P5�԰bȋ�܄��)z�T�Zx�q-IZ�TBq5��7�^�قn���t��X��p'��iܐ������[1�5�~#^�w*�f]�����M�p������7�x�\���@�����4	j���p:;�20L�p��ݾ/莕.#���-����)-!��Z��1�A>Fm��5���*�LG�6Y�6b��xH7�����1b�O�������0V���W��yM	�D�R<�rݰE�s4{+?�`�M�)y��꣆L�.-T��GWj�� s���#dP�6�fg�W(rGhV��h�j.������=���b$!h}	��9S9r$�3�.1ck'�����Tڞ=�-�T�&e���0���_�8�q;.M�ƎU��T�J�!$@>���A���	�qSB�&��7U�B[R�@���:c~�ݟa���~+)����;'�B3D�	���������'~�U��Ӏ]����>�B�e�`�f��K��ǛײN�v��x4nN��þBj�ݵ�^�7��T��rj�U,~�F�;��C�qѮԋ�4n���evO�]�3����Y6u�e����@�mdO+�;dHi|UGK��8d��H�NW'X̤��,���< �aK���������E��8�CY�V��Hݚre�H����)Z�����}��pM����ט��%x�����A[z��'��%1[��.�4��U�9�t�n�u���
����Ա���t�h�������U����ɧi$��"���\R<q´��߉��]�ͥ��Rȝ�whv�jha�O�9l�)K�[�Q��"��=x�*_I;I�X�}���d}����g�	)�aXc����s�C�H�?�%�`>I�[�A�ck�F!N�p̟@�2�/�7��w�+T`X�E׵C�c�%�$in;�e�%���)���14����V?�:!�"�q�zC%J?����pY��:ap��_���ڛ��j�?5i&0 �mA����‼�B���N��곢��k.@�_�Ln{]�������v����/���p�78ސ�����qr��Ztel���Of\LL协Fy�n�Cf�
�BChχ�͑���y��F
�O�XP��n�r,��U�� ��q9�:��>pc$��s$�p2a�î�/}�^t�I
l~ ��;}��b/.�6�����_�A����԰��[)��n-�aS�i�WZY �-�3�SB�W�d%g�-7!����?%4���L?��zX�gf9�8���W� �J��"c;n�j���]5����V9�8&��4�q��#ɧ'�-þ[x�YͰ�Qn��w�E�l{O�I����B����.?7��� ���6q���e�tăjй����!����(T��^H2���p�� [8
ZW�vjꖀa f�R~u����U(�s�ҚJ��S��J�޻���!�"�QГdȌ��	(d����8�i�U�9K�՜ ki�BL��P-^�?��_�%�(�@��[;���Ĝ�R�������T7_3f�����Xۤ�V�^���v���Np�,��H�n��	,��F+�����sc�Ĵ��!�!bl��"D�x�N[��.�	�i�BN��������s҄L�[G���p<��,]���<��_`���A��e���߾7�`?֢��$l�+C�]��2�`sj�>:\��ݩ�d�31"B��z��������e������:�C��Y�U-=D�ߨI�;�z�Yi��W!nW|#|��TpRh2{������:�3�Fd�-�K�\��p�Il�O�!�3���v��Ն�s��.N������4�KL�LF@"��菺�������*���v�=��aQ�݄��b���Fm<"�5�@�""z����ɭԾ��d���L:��Q�$�tF0zQ�l׃%��C�4��l<U�Q�T*s��'��~��܉�[�<>��� �,��e��.������FQ�?�I«֦�}d#|��mj�n�J%��}�L�:��M_%��m����}���3�~�ņv�WĨ���|���*2�1�BJ_��- h�!F����8�k�ǖ���Ŝr�O֒)Z�ę�	ܡ	��z.�;�?�L��˽먂!!�a����w�o}7}T�QC��W�
<���]P7�e�#�^�����h�M���eM���� �Luaݩ�n�L`�-?�ۏPPx?���}�����nςc?4��P��'� ��;]��P{xy�T0����ט�T����6cÝ��9d��=�`�$�p�4���0��7 ����x݋�l����G[�!�8Z�zD&cȔ����0w��M�J#�_�I�ɡ�f�!�n�f#�V����W�T��_Lu�����.�"��C���ֹO-�/��ˎ[�uf� ��ѻ�, ��d��_�^:d�t���^�V��f��r�����%��,˵jq#�ē>�~V���	<��k�&�c>�)��D�����,��Mݿ{��h��W����\��q7�-_]�0�*]q�]��R�N
��M����Ԇ ������T��UOXV�BZ�'3>�\�xN6{���/��%�d7yu���}@���n#|��w��Ւ�0#aZ�	�qlF<+�?C�A����K�ěp��:
�PXY#�Tϧn�>���=Xr�l�$_M"�% E������@�
�0}(���1�ǅ��!X��;��UE5��eAf����C��͙��U?Uu����l��\�O��ZY��o��3���y�V�v�DVF�o�9�/�FS\�L'7׳����A�|��Tn�$���v���<��zCQq�d◓>���Ď��`��Z$eD�X� ��ԙ����8/��\)"�̚��'ԾSJ�TA�}���80�)��ݒ���"=x���!�̱R==�mS\�>�f���҈��V��ǆ�ǧ/��f����W��?z�@�Zu�0�cZuLO��%�e��
Ȝ�#YOF�O&�	��F�Gø�F�(o)9�&�M�	M���v��y�Q�C^ŗ'�P�$�DA�F�}�؇ӽ����U��Gڮ��X����t�3ΰ�	`��"Yj%UҌ6�8�O9KK�~߼y���	!�G��}L���i�^��Ό�r�di7��A�~b�������N�������[E�u
����Kܖ`L����7�hV����BMb0D�c��?����ge��5�:�6��?.�#C��,8�0p�-��d�[����?e�m�_M�O��7rӯ|p�EpqW�5��?��ݱ�����-#���^Z�S7�v���̅=yدӦFϻX�Xb��&�������WԻ;b���t�n���\���-�����f�^�e\�MABʖ��b^>X�"�Me]B΋����̧���"��ދ��,8���Cw,�J����#�5t�ڻ��hS�HY,ܪ6V=ޞl���^k��W���A��:�s�A�r�4����]b��U�'���h�/�3�����"j�l���Ό:�V�V +le%k�e2r�#I,A����9����~��W@}��.he������)�r�q�c3���Vi��d��5̬!W��ײ)P1�H����
�r�{�/C��C�F�'�9M�T��ʕ�BಧYv��O�Yާ�MR8FoK]�x��	���|�_]�yw��{1�uM$��Wg����
�xR}��rpý��7�)'�I���%1�+b`�G��<�̧�~���No�l}��W�լc�&���n��{1�$K�GjɊɰ���G�I�X�Ğ[<G�p�)��HW����cd��r$�=5���d���:o�sS�T�@�ۤ%Ş0u�����$52�x�e3��j���c�«��n�4��f���Z�lȥr�O�T�m��bz71�,�	MSO�"��$���z`Q�#����T��	(e�@5,i��Ϳ���+�D�R��+H��(�rۜ��߱�A.�����g��H|�ԃAWy��㵅z���:eW�S��7GSL�[P�Eݽ:W�.	�����5����~L�&:��|OM_iyY�H����~���k���%U]����4O�����=��ص�Y�ކcN�:��@W�t�;S����&���Ț_��%JF�]���@?f2�������JJ�&��̘C������ʥ���9V́���()�j�:`���Q���8렄��jA���ʔ�rJNi�ICg��ָ�� �YJ�CY3؛�Y��>ѯ�8Wp΂Z�j��CA�x]��q�@fgI�"u�%_�J����*�@h(6���#�jM�q����� ����8�?�2u�����<�?�CC��|Q�ϔ鮟j��|:�A�i�\Ƃ��_u�mgX�k�]#/��m0�[��N��SX�faymI��y������N���^"0tn�S_祰��Bs�Ei74����
;�|+#N�.�8j��(���*)�j��V6��ق�`HnY�)�y���e����̘/��*(ȫ��@g��!"��|��v]6Er��,�@��uȘ�ۈ�d��bad�;��x#�7�E��ݒ�p����-By����*>�g��1�
�B5�M����&E��l����ag�����ۻ�^�����JΥ�_+�h��:2$�+�o�S�㶝��6�:��@�tZ�}f�Ï������;�h��[D�5Ѯh��7�T�+�~�$$�N6af�ph�&U[dS���z�_1�K�u�Oq�s���{�{%%Zv����x�1>��\�R�h��k�$*k8�-�o�gğЙ�q�ro�	ʡv<�o�-^��n��_p�hu
��Mܡx'�o��C��������.j]	ą=�S�WZ����$��GTݚV �������}���a��6B퀮ęj�&���IRn�������(�tJ���'G�=��!]j�91Z 	%��Veݧ^%��Sŵ�b����m�ybZ�pcLEBJ�@̇�Q�9��Y��x�h��� ��V��+n�F�P�.TO�R�E��<�Y��k��I�A�����~�w���L���~�O��^�$�짜O1S�4O�U�-g,��Gg�q��n�eP�����Pi���F1b�3��ky>*.G� �U�t��à=9�����'O��Ƥ��u����R2B8�x�՜=8[���O��=<��iu��`syh�&���p&�/��@�?D4:\U��C>37��Y?o�5,?�i����Ű4��� ����,�\�hƫ�R�7Ĵ���d�9&���-�YmM\��r��\(��lWi_D����2K
�� ���,dI��u�1���MA�М�;����2
��7���4]o9�(a�S��%���%���
>�^}O�C���C����Թ���1|�7b���W�~a��)(G��]`� �F�YBi(�_��(���.M�/��u6�g��0-�{�?�B`Ȃ��\�R�Ѵ�v ��!��L���q��<��M���$���>5�"'�*}�mʐ�:�#ڡ��ϡX\	�oe�J�Td���g.��Z�}JK�3-�96����~�I��+,s������_%���m~�ҳ�-�\H���6��t�M8^Z`��	�ƒ�y(n��Mx�ŋ�g�}W�RD�Xi��RݕW�7^�^f��O^���9�)h]7�z �R�?>%��^A�S!7z����ǆy�	�V!^SΑ|��i��v�V�S��#�*�Ӫ�Aև��p� h��2���r Ne}Z�.dŌ��	@}ѠAz����d�v��%�Պw��!��ќ��U�r��5;r��X��J��eޏH�����Ib�?��hD)����14N ��G�蟾������<�bc�ƽ�-f�c\��a���.��FK�֖���~K�q�Gw)�B�%�D0b#��G�e�� I���_~z!�!	a��M�h0��j�`TnU7�)�N4�f�ʎ� ����
����}��3;~D�yԑ��b����W��<���-�I��y�$G7�t���s�C��NbE�R+jtv	���U�Gm>��8�x1�ga�nHST͞�����!��jXVN�Z�ق�K��1��o��,tS���'c�N��L��7ܧo$(��E#=��1S�/�:�H���;'���<5�&O�L�U��w�� Y��3���zK;EcT��j?����O}�mXGL-̪�c�TZ��o'xv��IV�zU:#��=
��ón��*��F5@�g3-��{�]�~+�2=�!�G��K����@$l�;���n�D��?� �@ �ە�e�l�+ѬR�.�N�I�S�Sk�$d�������s��]T���Q��`�F������k����*H��S]k�.ҎpP����z�5����X���*��6�2����yV^�+�Ux�E1�v������شʈ�t��k�l;�-���(�Xg��*nak�O�Y�)f���J+�����x���ݵ������+��!�����!Xˇ�f�+�?�w{�E�%�������ow��y3��39�F�}��[�ƻ���`E	�;]�*����k������l�)���P���ϠPSsq��E�j��mK��K��A�|��̺~�/( c�^ް�'ڤt����	�l���k�g��y ���۳�v_�	̤���!g|]�/I�8/�0T��}�1����	���Q�����4���%�s�q���2�H���*O�; ��G�v�Vq�f`<��\���-���8�?�& �ڗ��=��c�3�Y���`ף������<\]H�n8 ��s�(�p+H�^��-d>����#Q��?�R*���R��y�w�0��_���٫^��TL�҃c�+t��l�:V�J����z4�V�� d��sJ���hC`�	�Ż{���|.�']Q�Z;Q}ε��>�xM�oR���bos9�K�9"�#�Hg�4�������x-�yF����:��Z�J��;��t�[��ir�ד�ʁ���xG���Պ��*���K���k'��!�d�t
D^�!H���cG@��.�A�\db��9��jy�9�6�+�Kq���.D��=b��|b��\���#Hi�b��,7f���ږ�hA�F�F�8���O*d$�Z�d8��q��p��`��@uhe_T��,r<�� �g=[�-��_�u�!w�!6C�,��;��x�*����ַ��6�a&�3�|h��Z������U�x�g������g�#}���a���>ml0�Wt#[ȝ��^�{^J,�����fq�� æ�(���4SV0�����X2�c� MAz/.� s��Ѩ]����.
����^�AA�&‑�a��JW�y��9�(�
��a��tC�cB/�l��Ԩt�Ί>�Ӫr�:����-:l{��dPЇ��\ĒT�0�&��~v6���*e��@I���b4U��}B�K8gK'g�I"�S>Tj������9�j��]U�lV�NwЅ���Q[�};Eg
(|MHt�ڑ�!C�.L�`�����N'������ �fC$��a�g.͘�f���4���?���Gό�Gh������Д���)kS���m�JՌ7��K3�4S!�٘���g�R��(�s岁�gԊc0��r���`gK�"��}%��Ұg�V�{��Q��3���(��X��x��q��!��[�t�Q ����/������I&�:�%��!F�X��ߕ~�~�����uv;����I\���{Bn��<�Ws��~��T�f v��\h�.(��arƪ܅���d�N����r� �o��g�I�J����N�,W�J9p����k��c%_9n�-�ci����\��:7_��Ҏς�!�.��ķ9�*K}��MH�������iZӯO�'qr�$JS����
G�b��l�s��9�$)��jf\��6C7:�8�B�P۠��,@n�R܀-�5�B�NXyF�ǳ����*�.�S?U�����"\�ezp�%���u#����]� Ύ��h!�.%��I'/�-P2�e��o�T���kђ�sT����6���F#	K��L�Tî ��f���˶� ��eJ~y𩎀�̞f��i�w�/�(��i% ��x��W�NRnF��rΩz[�����'�џt�h�k���.$�e+�D[!���n�eqK(�Ϸ�����.O<M��Saꫦ�w"���n�6[5�G&�跘&�ќ���c5��0��ڌ�*s<�����,��x1���0���.�̲�|_�I=�yY�+��)o�iQ����(�$1I!:�7z�A���1��▅�)]�o�+��)����]��h�lq^�d�R�X����B�c&�uh=��W�K�3�21��>/!���5".ָ���Y���#p��i��~��X6�� �����wV(Kud5/��4�3j5B�$�}P	�'��J�y�jv�'x4�����<Ρ�mb�n�ғI&�"+#�"7��i�N� o�Y�u�,4�&v�Dw��B���Z(�7ՠ�.�QP&1}�8v��a��YT��a��R����8�;{�������zֳ\`�7�7W��(k6p>E���Hv��\����	�Dq�
�0U��׵f!Fc�f���#Gz�sx����]g����J�}�Uc �b32i��yV
��!J^_���P����*�v�n��n Tގ�3�^_Q/��+w�`&)�HG�Q/�h�<�D��Q�z��k4��{�E�@-%
4]3�x�d�@2rY�%w�Q�<O)��������)'�Vc
═M��z�)z���D����H;�nD�4p�iϴ؇3li�J��G�z�Z�4�e�C�߱��(�dv� ���!P%�F9b��pӛB9&��6Б����J���-�)(01w�bX����p�G��&���u3���eT���Z�۲�v��;n��㓟��Of,���K�ƿ��F��1H?�)�������#����I�}I��v4&��ȋS��Kݣ���f�N	��U)+��e4�)v�-�8T�������ɲX"5R�7�o`�v�ޫ$�l�q%�T#�!���>��f��9��.P����4�-X~����%f,q��Z�@A�~�ۑ&���G�~��+���,J �u���h������3���7$@���@q�Y�>��p��R�ޢ�Y�1��"�-ň��C?�[��Z܊FV����:��j�	E>C)�|��$	���t�|޺��͘	�ȅ#H��;Dsx�n��i~^J(a��vn��oI�xeB�l/]��Q=�X������g�¾��AEK݆;�4�&�k�́3����=�9�޴��'1�����؆zsOtv}�\�<�T���z5Vӿ2N�s�˳�.�Tq�����޿	��V������_�f&��ƴB�GXn�pa'���eS��P�A)YAأu��J��U۪VE����s�@�ܿ5��r�;G����1۩�a���=*w$j�(�O�����o�z�`o��	f։��v�M'�&n�"�5��g��Fu$ɱm���sbA����tsn�˄38�{�f���~-+U�D��7<�KK,1����:�����@q�;�PȞ[V��W�����VY��� C|����X���~�=����P�&�ȓ9��9�7y�5B��KKݛ.���j(k�r��s�������ɰCE�����z/)B�c��b}α�L�{F�^�Q�c�����#���ss�eY�A��>�i\�6i&�g	��NAo��t�X��)�J�	n-:[����h�����3
dz�D�3q�@r�Sq��8�'��f3狼��V��V��'�FD�s��3-8�u�q�g:����5�9��ր�n�j"y�o����y���=��vO�����,���V�'�6��ܺ�?�u��0ކ*T7���=j����מ|Y���\,E��>�\n�bm8��Q��$<z�1H�j�z�+�qA�X����\�ংlL�2_�����	B1DH�ܝ�X���>�҆6|-��>�71k��8oIs_�nl}<R���=Dc�^d��~��y����-�o��=�t���8�T~�vk��TpԞ�𬭸W�:�BX�z�NFN���MO-5ZGtZ�����O夷9�V5#&-]j��/9�����^�������m$���i��W��Xӂ�n8�L�'���\ݜ�ch�ֵ.�h(�E��퇦T���S����'�aJG���3�5��� f�i��p��)���lB̤;ս�i��d�\�x�'�֖6���S}s!���U�e����q�����Ǻ��NY�Y�՝�B&}㛭N�8�d�Ӷ;dM�y8v���󃹗!6V����&���x?$�S�8ՃG�x&]/R��M2�V��J��1!3�Wu�Ι�1H�2p���}�J���z����g���k���t��S���u8'S������Ժ&��k��"ǌ�EW���`�X���l��m��q䀖��\�E�gc���;��m�n�H9�Մ�%�@��{a�}l�4�ջl6!��®~<�^��+��\R����6|���fh	-��YΜM[_��*#���y8q��K|��hOx@��;�ޅ.���7Iol�u �0>��w�ئ����uw��\i����%!&w�
j�e�Hל��pF�/�U�D]��v�|@�h�R����J��������\R n�|�9J�:�����D�*e�X��eb����)Rh��N���I�7FOS��Є����)C(�ȃM�Ư���r�:��!�����,$g8#&+d���H����>�[�-Z,��<��HY�.NC�����������3n���}������;��U��v]�%{M�Q���!�=�P�ToT=�#���Q[Iiq���+�l���1�h�w����-��	��j0bV\q[���"�܁-�����-�Y��`
�I�g�N;c(]�ĸqK�@���|u#����sǸx��W�ߕs��V?Y�p���âզ�$$9���߁Xb�ѕ0��WL@�T�O��U=�y��.cl�Y�SXZaD���?����w �dM��2߾�ݵ6&oP���W\�D�VL;U�6�c��{�T0�U�R����Ϥ��B�o��b5�%���C�cJ��1���vf�k� ��X&�b����*=V�g�@�B!��R)49�}P��FRa$�͠ipF[ģr֔<��X:`���F�m��}��%��:�iY�����Ef��O�@��ZS�~rR{�xyvc�,)����-9	�>��m�����\�'2�x<�IV�4lD#��8U.y���l�ӡX�G���?� �jP��ߝ���ގw�T�;��쳁��d~\�����U�\]��zvSލ�1��/�Z��D]P�s?fO�2Qg�t��<�ApQ��G�El�����=\�����
��P�&d��qf�X/s���~`Ё�7�����<)BT�{�(�&Kz-�� ��-����J@� )���c������V&��H%��
�W���1�^���viA��"=�&�>�l�#@z9Ӵj�E��|b&��7$#���^�L���=3V5li�h���A��`�Pz��9��_�%��\S��J���R+�i��Ɖ�C�q1�P!�
��~#��>�=YZ��O{t�EX �#@���Hy��g\"'�en���Oe4k x�;�pB|���l;��"X�#�>�:1r��x���g {�뻪rF�~i+���hYt�=)4��릮t��q|G�*��t����^.��Dkϳ�V8u��ܤ	��c��
���0��c��
��ϐ���{cf�D�,�+��eYa���q���V���+/# �F��8C��1�L� �	�yB�>�8�j.P�lsp��A)� ��R��Ji����� U��,��Z(���KaP���Y|U]fG��C���+_��n��$��*�V��e\�dX�������3�d��~h���G:��#�N�t��1��P��pZe�B����-�آXc���~Oofady�C������g��L/��c�ÄP���2e�7��~3��?S���J�A�3�D�:��Lɪ�kD,\,A�+N9����䌓��uj���#Jr��(��֭ɶP�ט-�:a��l�	�(������=�Iڊ�q=L���1���ً�P̛ ������T\��F���Æk/��L�'��嫪�����b��%��{@�E~��!=~P���*#�]�)D���hm6,��K���u�t���F�������4�se��c?Q�w�?nP?l;��<���5��YnP�}<7&�8ͦ� ��cT[,�A��)~�*�)X�/n_}~��߫d�t_&��M;DX��sDɺ����1�z�i�6��(v�ʓë��w1W�<gԹU��UsM��*����5����.���}���!��~lFܝf�*��lf��K���ѓʄ
�G���Ѕ0N�!��t�X|15`�;�D�Ge7ЙI�#�����]�^iQ�zfɩ��!W0�ZR��Pyk��#�˟��4�Y^v���ߦ�l�?u)��t-_�N@�r���B��;����5�	��g�D���:��b�by�f����Mb[��Z� 6�K٥�@�k:0�5q���<���b��x��UJ�"Ț�EG?��D��>��]�gd��7�*L�O�T�ge��&��1�*(�W'SWɌn��cBP����o���*�vt����|p��.�颶�|@��#�����If¢�=��W\:y ���sKq\|����b��֦���6�X���m�R7�-�OW�^x>�o���G�]g����^Aܡ������%�����p��	�=�~�H6��)g`>�ί�]����Ʈm��o�kd�d��䪞�n���^e�����P��z��ɫb�o�h�Ñ>���0F܀�E��m,�UȠ��@�/�omē��G��k���B�|k��79�r�i �2H�Ha,^��q'�v\��L���]Y����~�e��i?x˃��Y����ķ,���G'�� �J
�;m�f��:�2�dcE`�j_Jr�����Xr�{�Y�y����3sh���� b&~�[�i��kӸP�%��Hd,���K��xǹwJ�@��#2�b�i���f��|��l���-��p�������YT�)�_)��O#�j-ޡ%{���*@�E7�֡�����=�d�P�׶��bb�����Z=k���M-�SI3
(��A���5j�[)�[��[��H�[����V��EeV\Y\c�:G���Q9�rd���g�J�r�:���L�{��Z���m$��t-g�W�%���rE�����}�HMVI����m�bлB.�����&�kPӎy�5G$Y~�ڬKU�d�g��s��#yK����+mJV�u� ��dX��"��:��}����.�e���
����Wq���H%�c��nadr&���t�h����;(
@@f���\���w��OF��@#y5�P�n���*�K:=�r--� ˬ}��rH�VU���(�?]�~�1Z�/�D����0�L�3�>�l]tT�W���[���W�ǅU'^,�Ԑe��RO�4�����]���k��e����R؟Ya\���������k��ЄxD�	�ue<8z�Ư����$��@Ń��^���8(� �=��\r
���!�f�-��#z�0���hJ����ɡ��f��4����'$��%��B|�:���D�B���oe�U�'��;�cW����Z�1���	�ěÕ��%�!��MI�e!O���*
�%��u����L��������k
�g��<�F*-�Uh��_��9ܦ��P>c�9��;�j(������ik;V{
6�s�$�/$��1Ovk�@�`�����ÏLZ�IYĩ�hV�T�vؠ�޴Ͽu��������ndc U���t�]�R&_���ؔn^ۍz���z\��,��0��p@����޽�k�[�f��Zs���	�b�'`�Q0��C��ļ�<�(�vt��ҹ �|��c?�n����� ���[�ڧ�[)�5�]+��r��,�����Y��a*�ZoxQ�̺yط&$��B�%~!bE �_96=��c65�]��X7e<�(&�>9����rM�6������=��~��b	tp2�C1(�y� K_�8Z���B΢���w$��\O��U�eCB�S�����s�ґ���#�T
;v�Ql���9n�EIJR�I@�^d���y���]�;Z���K2�-z��q�A.���`ٷ���jBo9���
#���S���q�r^1�D�n�34�S�7�n��4���Iȃ}��2��M4����>Ȑ��ַ��3��=��S��=������p�6U�]>��YGD[vS�-G��پXӐ�$/F�Prh�zҎ��m�|ѩR�Q2pk1o޴� J�4:��ݖ���uU9&�|��2~\�6�=)�������)��Gޞ͟��rGX�>�`��.�0���!�h�����l޷�ie�fA�aq��&F�3��F]���M7�t���[��m�����C���z�-��ҸC��&Wz���sh����ԍ�������o4�s�4�!�Mzl�4�m$PÄh�Y�G�k��ӺG���C,�G��g�CĀ���}��[�^���ץwu���=E����?�?�)�7����ć�]�|¦T��DE�S��`�����D�PD��ݗgb�vR�Mġm�&���kzl�2!��ǡ�d��������Q������Ux�#��3��Ւh�}��^�I#���V2�nI�З\� ҁ�מ�䲎��'(���1�K���Tz�g��!��ep͵ӋgmA�� �3H*�;
#%��ck��9\xX������X�o��y��I�8/G�2y�%�����M�w#����a+ټ�IE�� ��L�����S�ja�"�7��2���pDaG��_7�����4�����H��q�����{٪Ł4})�v��J��P �}O[z���qc�����.�8�:"�{���T�ǰGw��[�:�fB�a�u�wp���.s3��T��s�����ħsA����^�H詂 �0�&a��n/�*>���u��]d7�ކh7��C�u0�,m١��!/;8P�^��r��@H/N��.�j�ٯg����ї�@@���
`�4��<�h�ȷ�a���#��s(�}�~'������:.�"��p�]x���>�7�mDNV��m�{`�6/g�x���g��uM��+�w9�$�'�;�?�Fj�t�_�B`^����ڔF���%�)���$ـJ�/�O� 2utA�\Nl��<�j�:z06<�Ό.��yաw��������b�r�E1R��ڴ+���r��\7�v���S?Ш_�����b��8H`5,s
�~M�;����xZ�9ߣ��븠�C�O�,C��������Zw�6����{x��6�W�֦T�E����^�s�>�~=�?���?Cs�HI��Ǉoq:�g�+��߾����m��,�0f|c+!,����w#|L�km��!«(lQ��9Z���/r0�A�~�
�Y��Z�a�|l�N\4�1V�7+�.���m�(X,j��v����(�&) ��b��\On���l�C$�)����_���,����~��D�@�7�\�����Q(&��z<n�nG˶Zh�|��}���Cgyx{��wG� ��l�sP�1�C%�0'��������ǛI��c��٬�Ԍ7(��,K�5�yO��8��R|�:#d�a�9�H �����	������b`,��m�����3EljV5�����>�tpI�h��<v=����d��"�Z��}�I]�
�w����i�wj� &^��Jֽi�<69��ZWc�$���7o7yu̓w��M-���Q�$�s4��2.ω��G�iz7�A`��˝��=pd�)����/,~���ks���n����`f��Ug�P���zY��o�>|�|w޼��z�O�����7���,u��5;@��H�po��#�A�s����*��h7���0���ޖ�HkT[X8���y4F��}Ɵ�����k(�K�9	�ޯE�d�=�y�V����kX���W,��/q�/���/3� *X��1ͯ[s�^<�_ys=6jR/��RϽ�\����TL���\Ė��҂�qY�Q����c	 ���U�mb͆�<�R`i?
�˲��T�G�A�Ĝ(k<��1$����B�����5�]$� �frFw�K��aL�P��+��T�c�^��?½s���U��ߢB*�2џj�n���~��_�ݵ;b�#r��J���72?�')����k��W����c�=C��@)�èI O��g�{#s�GZM����'��>8�|���3�+������F�䵢A�pSb�����;1i��ߝ�E=�t��-Ou�t��>|*�ذ��gS1>���;�������B�ڢ�e���+=t@����y���P�1���L`u]۶�;�uLgir^v��u�ȑ�r�Y����O�:}���&�av���;2�s�j_��`	S�8
�!�bҨ���KU�9��x	F���2C	�߲r4�Q�M�V�C_�>���HZ͜G����L������aQxloJ��I7 i#Ճ�ݎ�vEb#Et�����L.��u�;Yt����)l�#u
�7�Q!��^9�֕&�u�rx�"|7o�sp%�V$�wN��S���l1deF���:!����Ą.�4A�_��z��g�1}g�֎-�-�ζ{U��Ni����N*�+��)Em3.2��U��M�����u:�ͺr���/�qkp	��8p�|��i�DGi�W����jT�M�c�h(� �خ|S����8�Tm`8͡�L?���=i\��9՘6M_�ܭ��%���%B������.��I>N������o�B��+�@4��=������:@׷ܓ!vc��u�pY����u�;�u?�Q�������ʵvN�~��d�Y$��2�l=&:�G�uF8K���{�"�ky��}蹓)G����b�K��6W��Bxt��M���������φ��m$��Ll$Hqu��5�*F��Ko	p��l�Sj��WW�d�v�P����N��ގ�e՛1U��~!���@"���L���7���*�Q��FKd���G���e��u�l?9�T�b�#c�2_����W�R@�z׷����;���:ʧ[)�Q�n�1�s�?��]<�@�0x�R�n�!I=�mZ�-�kPܯ~� ���Py�&��!��sw�)��k>=��!呟TH�kvZj� T^�[,�k�#��L
2�1v���g|T���[��l���WgZ�*`u�
`��(+��| �[�mJ΃)�y((�x�	�H<{2ԩsr�#NB�,���Ӫ��RM
���sm��aظ�?��"K����`���D�b��+�s���|V7�<J�Ի�!h��G#�]�Vf�?��ժx{�0������)�
#%�����K��U�e���Y������I^�ܸ�ޘYnC!���N��:SxQ�Fn7ċY΋C���,��(T�A�>M6T�ܿC��	�λ8d�g�`>W�S{������D�x 6�k�
�](-�}-%�"�=���6�8T2�{�<D�L�����Z�'��_��&[e$�B̙�zp��B݁���zַ��Df;�lw���)���"�x4� 
v�	zCC �cN�s�1;�G��O��4����5�g���J�w�,�	ځP0v���E�s�C��B��F�!G��Z���R������8v3_bl��ZL1k���%ņ��3o����<����L�X�Q2�m�ZR�'�$d����(���c��c-�%Sx�S��ƞ;L/ w�^0���ͧ8�~�PX>ɲ�D��/	��RzJ�ˇ/���^3������|���=����؝/xh�nb��(\!��9u�	�&12D	��ʌ;�Ɗ�)eP���z�z�s��Ҟ��4e���K����Ǥ��tjB���&K��f~�B�  _e�'�|�Y��vj��;P�"�]N���ƅS��7j�0I';�����+�|M��ҏ�pzn�����F-�c�K�:�]�������p܁�����sQ�� ���1���6���L�(�x�	N��eE[u�]��X������,X�7���l�>8ԉ�/.?t�gs,+���*7b�CѵP��f֎?6���JY���r7%�c��s�'$��"������J�݇����ȶ�/N�.�W���[�z��D��s]�w_���sU*a�i
��k����E��l$�������@0T}ZjA�<���?��\�Vôh���S��W{ô):��UV?eP��)ݾ=�a���3�О�~��l�Vۡ���VƑ��8!F:+�+Gz�p�?^ k芨�[`¸��qI6@&�W�vk1��ңJ ���!N��X��M<����I2Њ����|�X��&VL�9����*<�*�8�,�5��#'ЩM�+�oz|t�I*
���H��$����@g�U��g��5b}�pn����J%r��oƽVG���N�m�Q(�%h&��Q���3��Dz�ķtA��o��9s�x�L�[�P��Z�9��M��Mj�3T�Ԓ�F���;:�?���?�q�`��ҏ�j�T,���@�G>���-�s7|��Z�Ł���{��M)�"^"�wLE�@w�Z�FԶ�7��r~���'�6���hi<w��������I�A�D{��o%���b��O�-�C��DL�[�LK;�����LR07���*��َ�s�!gT�W��|L���+����v���z�ϒ�V��!�)��.�l�5ʻ/��+�Bϣ���!���9�)S�Q*��q�n�S�>��D���=��匜4�b��@��G��+όՍ��"��" ��a�l ^`�a��b
��H��)��h�2mt�Ԭ���෬3�� ��K�|K��[|X�ہk�FR�?;��e�D��l�P;�g0v�p+ni��RVF��C�[�F�>�wR7ĥ���:�Q[6~2����X��X�Dbh�tda�Wų�J�dT@ᆓ`��n���v�˽V�v��@a�іyXʁ�2��`����Ro�ym4�F��t/�w��Hf?��=��T������=U�m�2�|<��$����#�a�OY��jT�dG��LQ���A��$*����{� �oY�����D#�}�tL��z�T/a��Q.�-�e\��8kPv@����c��X�eV2~R���*�Q��
�e&���;�f�~�Ŏ��EkX�d��-�J�{~Dƥi������{j��v�N�o��w{4�+��C�_=�0%)�2E�'�=�*H���V��Sz�f�����;��+��ՠT�|��r�X+u=|�kb��Gd�S�B��3���s�.�t��Z}�?C��2wmpa.��2�NUz����kݬ0�Z��ʸ ;����w��=����<�c��<�'�MnY$��9��f��3��UnKʗ�P���݋͎}�"=P�HWt,u��DiE�"��z�	m��'�r]�@�>)o��;�>����6����@����8p���/�ИM���M�y���+��Ԕ���;�^�;��*d��'Qg���^���~A.%B2Ir:���qUz4O ��c�J"[�#Zd/į����f^�Nt7 s9e�RN�,�6{��[���� ��B���j��{l,m�;��)�O�ȣ��7�n.���B��/�}�)����c38n;�U�s��d9��6��I˽^�Y������X�W��{��	�s�3�b�(c��Έ�ylz]��rC����p-T��z��lؒ�qNa��}XݑRg�fBH�$���{ٻ-���tb�8��	Z+�������hs�J�\8V_���X�0O*P"s*��fљ��>�����N���\|�7:BV����r;X��EF�)���E*���_1�c�+oG��zN��-��j�a��Ӏ=��ß�&�¹�����+��(��x�Ȼ��["~�����{ʘQ���s��*k5���l�]
��ycx��K�M"99�ޡF�8�o�\�ݰGz�0��V=E^�f ͕�9�	am{:5,8�;e����l$�[`w����Y���Z4.���һO�0�K���Ђq/� t��=y&��!:��bݗ}�׋V A�J�4�B��>�`:M���A�# �4*.8.I�>s3��N����t���漓�$��R��S1Q"rpO�3J��,�!54��?��C[ZL��	�[v��x!���ܰ�������wC"���i���\f��b`�=���a�/�w�`7<!�J�<��Eڨd�)�,<���d8����	�˺��%Fy����/;��,��Y�ȥ��i*�f�f�N��	ke��~8�b[����o���K�v��4�;�NF��B����S�Mj9O wm��A?�]i��̼`���VD��j�#���4�NDH�a�Nsa���
f�����;�i�ﰦW��[�a�i
��p�HU�������$�J�$A<0�V��0M��N������N��<��B^�:f\���aWݍ�]��8�/z�]���vxO�ʹ����.�j�����I�,r0K*{��ZL�}Z3��`�^��v��n$�~yj���CCkHr����q��F�PH��'��H���j�'?�*q��A��(�X)�� �C�,2�UDS���{Cሼv��sZ���;�p�o�d !s
�S�z�OCTN��ynҒq_�{��Ը��1,c�_8eG�N�P�_��ƍ��x6W�&Mh�QX�?LZ�gR#͍v��}�� �\鼍&�9��p��Z�[�3��=���b�=*��Ю0�
@*'�'.X;B~��MUu�zw��nAܲ���}�1��a�v��EtKj s'��[��	�Et����'���՚ �)�|��N��5 '씘6�}��@�ΰ�n�x;	V�`��B>4<���z�4$�F��Mf��z���sr��x�h����a��BC�7����S�PO�>�])v��ʺ�5�coퟥM"�l\~D�J�a�b�!:���NK�s��/B�{�Z=��<U���W�hJ�[0z���I���.�~Ý�haAّ��J�#�C��?�>���Q�6����vm�ƸWv}�3ή�g(���R?`��vu�ǧK��E|��+I�e�)�(e��x�dAg��˿�&Eu�+������=g�^�����l�齪}���4R�A��� L$�!�����c�K��m0q��<f>��Y�L�#�
�˚���+��l���;S�c<�n	���|�w9F�/����8����)�c�(���Z3�7>������Gj ���S�l�.�.NS�ӵS��Pʿ�.*� ��m�r���)�l`���qs ,�}���5Ё�Z�ɳ��l(���<U-�R����W�G�nC6S�E̚�|�p�H�E���Z����ne9�#fA��~Ƃ��}Ieg�kl�K��3���2���>*�E�W�A��쥭o�O�~�o�����Ա����(-�w���g0�[wQ ��k�8��?��%Q�r5��7���WWLǻv��y��j �θA��q�u���[�d"#EϘ��Eܾ����(��o���7�p@C.fk�z�q��D"#�e�+*Q�M�Bu��+t#�B�g���a~A(��+(9-Uiڔ���\1�DLN.�9t��:�D��]խU�a��R#t���9�i����JW�(D�i"k��~�&�[r%�z%���8
�^܆O�k�m�}�8-��:)�����ć_��%D�Uiw����I��Zٱwq��OF\j~3��j���`׼id��V2}�>��t�����з�7#փl�&��MJ O��H,~�k8�,B���l����XGiw�L�eY�q&�x>n��D&��u��F"��r��m��j��Z֭�|��娘o��8�wZ^�G"���O-����p�g�z����W5	�gx��I���x��hT��E���T��]��!�;��r����FV(:���W�R����P��`W��×^��v�:��.�}�'fS�[��,�k�� k]k(�nϾR�$�������|�@g<��=��h���zf�)�Qj��_M(z�)Q�?B��>x(����S[�����좋�f��H��X��?@5[��� Odf?Ao���8��xCH��$~��^;I1���~B�Z��|�И7&��C,�c�r � �&!���@�%��2b�(�����=��s�����m�JLT� �cq�$#�Go��o�e�qV]N�Zb:s�C:9\&����S�8��0_�B�0�&�..��O/]5��Vp���7/��桺���m�
��e�IR_��T}�`�y�P� �
4����|B�������+�`R�1�{-n_���:�`���k�'4Z���s>��c�n�՝ȏ���nk���8
���� [7N$�h��q��֘���ܴ6� ]eLք@s1�*a��w@Q�2���/��vaS��eY�����b�-���I��9�1�Kw�E%c현��Lhv���5�	�'���;'H8�U��H8�4l`c[)��EZ�Z*��0hrJ�������X�XҜrC4���T�E�|��'M\z����Ak�c��se�]�YUI>��[J�>5���i�^��<8��b��P���-�F?=�
���4_���2�����6ްN�iU1�%��c��n`�
L5m���N�eE~�)��.M�a:U�c%�-��2	�����,����rN�}G0@x1����3���C�RKe�A���͟�QN���Dr�<;�T���²e�Ur�R�ڼ,轀��E��N�/��+���^&��ۗ���J<r_�a�6ج�.�D�)��`�X�$z#k�gU���@M�:��<�|HT	��o�ϼ8^�9���峠��D�(;/I)1��� �<��o9��?��ӰF��iТ�7����ҿ�L�d�Bͅ��nŋ%���sv$$�(�ظ�bh?_N�U{�&�>Sk�sf�ث]�)���h	bVW\2��۔>���,G�˖� sVכH��*^�x}~U9��V��x�l��%W�ZAƢF�Vv�<1Pc�z&q���R>d������@�\e�_G">ֆ&ʪ����S�1�y�-��<1MA�)�ץ��\+�T��Pr��������Xy����F���8z�a߮�z,��̟�Y�ˁ��Cڅ~��=F�����`
;������>"yA$3���c�4�Rrڽ��l���:%	\W��D����wV��� 1  j�sMLt����`ڔr"\��U1nB���E#�&F14`Y�)Xۂ���^��O�J0Yr�Gc�����
���/ءltc�b�XH���G�GV`R���9��F%n�>�N��=B��^���6���5�-��14SA���c��8�]u�hݚ�>qA�LI[RR�c�W<�6+9�[��9�p��-NM��Az���`���pЄ{,��6}�����;S;�-R e��]�n�*����1h�#.t�t5�ҨN�F�
}mX j��!i� ��>cz,�x6��Y�*'�����B�\R1'��x���yQ7s:��۬�=�1����Occ���0C���"#h4{� �T3C�C{�L/5ۈ��C��/�2T��ʀ��$U�W���k����ŝ�����d�?N�\{R�������1�|]g�֝�v�>�I`�/���Ц�qѰ[�w����yT��q'���M"��}R��N��t��s�ǐA�/Z2]�����K��c��5ӫ��rN�w���֕����y;w���&�Z�%я��8�M�z��<�Hs�tŞ��5���O��Ղ3�h�-8���G����o8��:v��~�Վ۰�)����	�����n���|�����sh|z��!���\��-�����z��T�B����l��)����C�{"��"�X�{�Cd���B@E����Mr!�0�u+��;0����Z�^m��$.I��A�x\� =4���~�k�IL�E��q� $^�N\H�,�(m�k���'�O��K��a����]��>��F�iVm��W�]Z���'t~���n��l�i�zپ ����i��;�]C���M�?�&�n��ٌ1ʖi�R~���T��9X�mӭO~�s�t�P~��{������X����4hZ���p��BQ�9�	57��Ɂ	�w)�\�.��0ڮ7���NzC�"�ӽ�#��M�CVи�O*3im~L4(k�k)�f`���y���!����|�K��Av]"�q�ge�̯*�
\Z�8�v<ߟ`��J�
V�|�]���er�u�:��]�߂��v����P�n·0Z�j5u�u;LuI�L�C�[Q�^��k�/�sl��L E��L{]�:�24��{���� �޷��C]o*��|J����])Tg��h*�^A�Zp�CtԶs
��_���%�a��R��VMrf>>!�FD������5�e$��,͔��X�v>�����
���o:�H��ӹ��麰V_8C�Y!�R��-NQ�=�<�nj�M�+�4�sqǪ�e�,��qU>�;u-����Mz�f�kh�$�&=�Nś�PNA������X�d`<�b�����]����d��S���u�����s���t@���Of&[b%�����ʑ���s�0�G7�\�*.5���NE�(8CDv�8���{�N1��E��I���[q-�8ɶF�b��=��U��tf�?>��j���LlI�2r73|��`)�(����f7ȡ�1yk�h�f�t�.m�M*�G����,��T��^�\�ޅu���=��������=qM�cd0�w���e�-��`"4[���Y��,�B�"�#mx��~5��R��A��.��B2�c���83Jz���n����]Q_�yv�&f�=Ai�%9aIl���4Up�]:wت���sL��)�����ɑc�&����jmO5J��ֈ�BD��ʕ|�z���+���e�7 ��5-t�����U�m�����������΃N�Q�%�	Rl�D��>�2�Y��ڱ��L_m���Q��s�zUdRl�TA�إ䠜;����_��d�����gR�\�$��%�Ӻd#�#��_S�ԛ�{�,^�6��BQn]��%�0���Rs���y��޺�����bwd�>���{�Rs���ڠjj�K�b���+b��G���l0�Xx���S�T���;%+}#vd	]�Lڐ���W�^3��~$B��S��7��`��=�|��Ȋ��@���Fm��^[��,]X�;�Fs�A�X�L�vABi�:�V��h�m�F�h�6�๮uKR�����v�bl?���+�h�3��'WZ0��>�Y��Q�QL%.6Ԃ��ŸL�!�gA�&Qsg �'������̫�Ԓ�ηga ��̬=���I_3��N�������y��;{�w���58�G�-�E����לi��ړ0�"ȓߦ!TԽ	%���H�~�5z�f�y.��&X�|�1g�E,����y\���=��;1�-|�5YQ��|����bk.P�.�|%��|%�}��n��\,�e�yy��ɨk���c��܆%����s^#z^�!�����F��8T�}���c��ҿX���^�Z��z�z���Ŭ~KY���qK=Xe�|���x�<��;��	�b16��
[���C\h����;�XÙ�(���Z�
������q�N���Yz���հ��ȁ��w��ot~y�O@B��-�bd^%{���E!�7sAZ����2�q?��/9i���2M#{�#1=O"Vk�5o]�_'��s��^������յUI�M���˨q�Xl�+���M�P]��B���QPPh�)���"G�k�Fƈ7�X]5i���y�Cˮbi��߃fi����N�SM'���ySٝz
v��R� �RL��i]�ÊB)&z\'h��w�f#T i��퇬u��=�b�`p��?q�JR%xsP2Dz�u���x)q:�V�Q"��Ni��J"�*�����s�M/^c)����OTc�𵤴D��'�cº݈M<�)��hШ*�IN���j���� �Ô0��Y�R��3J�2�v�+��VF7Yy�DT�a}2V0�sZ*���r���G�o1qi���6O��g���ee:��<�HL��r�5D���!����z>T#Ww�DLW'q�!�r��F�|����Jꕐ��}�\$3}ә�Q#�XLʩpu*2�����	�	ۢ�|W��>�ڦ>l�jf�������3V�%X3������wٖ��
5���6�M靪���/�H�E9|у����d�-� y�mA^'SX�Yߎʺ�ļZHǎ6ܔ�u�H��W�^_1��8���,������m���J����=f�EqƗ�dΊ�B���p�:��|����w��[L	�<?��r�8^�m� 8+vB!O��(�@�zS�4��� ��'�ܞݾjJDq%��A����l:�"]���3�k�3��cm���-7��0��/
�m�OEz\2Z�F�t��˒�Y96���(A���<8	�3uF����^:��#+��L�$��9XV��
ѬK	��e�4wT�gf����k�U�;_�����`����w��0\Lfn�s�Ɯ��YJ�d�̭�C�I�I�7���+-�8a�)ge���Y�>%�4���t�Ѓs�$��Q���ؐ����Ū)w��h99�E�ɿ��M����"�v����>�m���[b�)��p��>?F۩[�f��^p��Sk4�p�_���v�+:I��9�.k�֖K瓫���M�:a�H�_)k�ǳ�Dl����Y^��}��&��M@��JD2[*v��.䡁�m��q�L�����d��X��]M����E�G�i�� WXg_��`J����_bJs�7�Z��&�'_>Πj?5FOG��@c/�4�͒�f׷'ʏB<�:��da�o���&J+i�P�h�{O���H;@n� �'�O䢊r����g�@� �����������\!)� �E�|����b���ܔ)�\��ޯoI���[�OK�,��Ħ��,WVNU�E�i��4�3IWT��8M�o����c%&Z��)u�m(Į�ਃ9I%�;��(Vh���_���Z���F�ȹY�Y�s���jt<l	��eЏ+oP`�:."Z����mu�!CV٩��j�F��y�D{�V۪ԕ�؊a���ې`���"��$N�3�I�[|��q�r�
n'�<�(�'f�RG5�Lml���ݾ��U�eX�#5E�^�Ě�n�NA��A�����G[�|��XA�o�����lѩ�e��Ǩv����	�>��ޤ�{����2^z�8Ӑ�F�0�y�8T�Dc�Q���x���	�Bu��<�����X}���5/!)I���`	o�iej&iR8ɽA���ts]l��٤��"��8��P��j�[���*�Y��ɽa�����/�'�rE�����) �4^1ۧ�O4� �(4Ȱ�b�Rj��.1]=`�[R;��Rr^xјh8."��3v=Q��j����a(9h�D�?ʈ��T�)�.ժ��7Ƚ-*��G�T=�_�n@?EK Æ]'Q�gv�V��c �(�6G�!�^��|L���TC����=��:�-x���z�N�!k')s�8G��o�ۅY�T�^������>���q�>\9;�9)�~�4����!�������p!C�S\A��Q:�ν�#=�A|j6�md��������ީH�i�ҟ���L�VA���]�9W}�����6C�����KΟ:w-7�T�5�ڪ[�Rߴ��D���ֵ_l-��bƨC\$9&��$�����Z�i�׋BK>9��f ������IR���یg��UVdJ�S��5p��V�hE�4�~�Lu����(gT�ts[2�
���@���z�W�]��h����a9����K�]G�,@�ᱵei]����.����;���V���A5���3��x�TyXf/&�<��)�cm�)�z@�~G\s�d޳���
�~�Ut�/j�ߗ9�I�)K� ���Q �NA�R��J ����-EW�<;_�k}���i�7���*���ߑu��F��{�pM��Ǘ���8Aߟy��3���z*'���f�r�	l�" �1��A����U/�.�axE��y�f�����!Y�"c�� A���	;�\[�D�D["O���3q�T����ܾ��̰�P�8�S�\܁��K�<���MYJئ�+Q��&�[O��5f��kc�<q����V�S�3����9�7��*�qd��b��N�$�@��s@9�rJЯ�'l�X�fP�?l�{����>��rb�h�����lǄg��i	��Ek	I���-:
�� `������
�����������l�Q��"Դ[���X*���BF��#.�f�l�y�);8�yP��!Z��7l`��j/�7G� `4"��%�A�.�{���=��/z��݅��%�㝦��Ҹ��
�썹sCj�$\͵�HK���'�9�Qd��ӫ��&q+�!���E�R���4��=c�!Q�\W��E{C��m��|�!��f�N��Tt���H\K�Ou}�0��\�������7��A4n����	Aݖ��펏�s
��^no�]&C}�I�p#"�
��J[�C�y�m$���{Y�.A`M� �D�lU8x�a�_-)�*Q�p���F��}�����:5a�Q7�.�=�$���8�Ipk�c�qa�ר1�k�W��G�٥�柭�eڄ��
E�c�(8�z~o�0��:���H��6�C&R��b�ɺ%Lv��=��a���BX�w�"�Σ���!jc<:aȢ��W������9����2�3*��g��QȘ4~;tV��^��1f�[6��S�"��c�Y݂lŞ�m@�%�a�*Kɉ��&E�y�mg�������-b@c"e.���h��aoK2	���H�t�U�� �&q��.������a}upR�c<�ھ�3��A�e�)��!I�����6&��U�0��7J~�۴�j6��8�t�Dգ�[�H���b��HDK�y�L!nûQY�%�ˆ�@K�xm� 4� K������I\1�� ��f%Kj�q�k��W�@��΍�؅��K������bԍ�T�7��ҎR���6�Z']�gB��qP�}�`���v��8������"?U��}`������r�|��Um��pcS�撱S�H���N��.0R~�oH���ɚ׫�!(Ta*����u$$�)��pG+�诸� Tq^�/'�(�7+�H(%��탯�KY�FU:��7���I��'c!��l�ץ�#�u`�׀�P�s�w(�;�}%�E�~ە��P�1�
�J�	�� 1�6�D~ͦ(��'�2�Sl�t����������ƥ���~�6�a�Dt�U�C�x��	�� ��b�	���N�!rL��;��\@$S@ƶf'ͯ�,����#8�|'��2�e~_�$?��5�ó��U��z$N�-0>�aTM�̫m!N0��5>������H��w�0�8��t[�-89K(����r��B�%Y�4$E�cU֠���c�C>PG脇Z)�����9,�W!$�x!������ƕ_��G��I��H�s�H�K�,�XPk>ʟ)�s���/ �@�[��u0�bK3˩�r?I�-W.hs�qs�L>E��W��cw(�2*>��{͈<�A�]ņ�KY�]m��P�SY�9�������va�>1&43�^�,0�;45*I�L�>�(����=�9�7��[��Qr������hgI9�Ӂ=�Q���iq7^��T�8NLA*������|�Dا������Lф����|9��zq�5`y��n#�c�������us�8�6Cي9S������)=	��ca�l»C��@�G���!zd0���mE8G��Z�c\fn�yО�{��ۛM�6,�0�ny�/�?�B�[�����z2�䔺�ԉJ��E�bfŊ/����CV|9MreA���4���Q���J>[8M��B0a�I���}��S*=�E�j8랔����;��;�_'CŃ�U����u-��!�z�|J�7MT��xl�c�)��F�#4�^L��da�����=�Sl�.89�����=g] ;�a�.���1NfV~V����aU����G��y��t�$N>��<�.2��������
�!�t��%� M�6� M�|]�ML�wa-�\1���a��8��R�i��O-����;��=H�Е�w\]��Foe]|����_v;6�:�b�b ��\�n�I��:�x�'�������jޏr�ݔ��C{5�@i�?�m-n��s
%۲8��d��f���`�`��\&N�Ɠ�(s�߻��x'����5br�B�2����)G�����d����\��8Τ��fJ-�bZ<���y���lA��t������"X���Zc�԰��է�A��S��;Ͼ�՛��]T�3��p�<�s���0�A]W�'�F]��Boq���XdxTG�n~[�%��.y���"�͵�Z/��y�-�����@(3O-����:�� ⫛�W{dh)���(���_@���7�ޡ%?N]*���W�{�+������T�(3w_�i!��5uU���m��&D�11���T�,�����~jXF�
z#~�w� �6XT�W���FxM�l�dCd�*z�e��'Y�=X'����p갷S
�Z�k���36��Y�����I;�)kR�1n��SɾԍV �Q%��d�琳�1�9ٗ0i�����!fv�`�a�|;��R�6�����T�5���5L�h���Q�x�� ��2M^*��h�霅v۶.�d.�����i!�Ǡxfm�NW��_�{<��q�����8�a,�N��T��U?͙+e_>G��k�{� �B��0�N2����u��*?��κ�(5Ҹ1�\yE ]%��T�8�U���Fδ�K�^��"'�z�i�:������3s��)H[LԕHP@4�;�i��6.��G�GZ�+�4Q�˙���q���o2`Ĩ)3� a��B2����P�
��jO�e�ȩ�43��< �v�����b��2J�$d���ٝD�B,:͗(OS���}�*�N{)����p!��z�#;5�j�v�d)�\�b��5��Ԋ2�
}G�)K'qB]2�q#c4�C��(�G$�T���Ե�:�UA4���:ls���l�)S�؝�Xu��6�|�W2��^�~��WJB 4�љ����5��c����i�?�� 
e��������0=*b2%�(�䚈�;�������¡\2�~j�(�Q�ȗ�2k#��Ԋ�8�CM�Zhb�x�2�Y	Y8�r�gG�CL����k�a3=���q6���^�"}*�߁2/�j������>�O����HCj�<�>��D���5���	H��H%�tqP��ObCK<^���L�a��Ү|M�0��������pw���5P/ ��G��aD��v�1��}k�>d!g�#tƼxM�(-�op ��6�f�E�\0ѻV���Jf�?[���O _��]j�A�Y z�#x�����*�ł�(/UTA�2��KX�/����۱cî�m�ؖM���[0�-V!y:�����gu�_��j�[\ �@1�`����.$�T��8��`��5����.��&�+�Ն�œ�o��$�.<��h]*���Ȍ���^Uڲ� X^�֝#�j��@���晋>Dݲ:"a�
d��%\�C��(��$��r�W玈-��'3����S*bN�M�����Zl�F8� ��먟��}N�I�O�G,6���Le��u��M$�A�D�Ŋ_�eR�>��<�r@�zڙS�Z���C��Em�3;g��=I�� �gI2��?��u��p%�&[ z`\Ǭ�V�L��
�m]����5`N��+1IF�����1��9Ȥ�z|�j���bH�]���@��9Rk�U��(�?�����W�@�,^\ 5���駹!��Յz�xE��(��)�j׌�����ӢA�]�	W02��@��/H��\}X.#��.9u+,�Q�5z�z�\5�r�wG������$ �	Z�$Er�5+��'��8�\A�?,*� �����=ǥ���1n�G
�݀2���ԧ�l�;'�D)����Y��n�s���n���h�WyM�U �b��G�y�g���h�Tb�gh��W��oi�>��d���.ס�g��bF�(�R��-?����<I̜*�W#��Ԧ�,��;�W� �a�:�|L)8�N_�)���q���ZS�����O&�:4���}O�&�ք��r���b�Ci#�­��~J�I�%��L�l ����um�8o5*��F�^�r��� )4�]	�M��4����T�u&���k���m��Z��E�B;�����o1W�s��x�t�.~�cr�BT�>Ω���������_�c�����������p�a�u��M.��ȔF��<<�>l��K��k�F���G��Q�7>E��=8�h彰�7�З�-Ѻ�	�aI8�f�;$EJ`b���-�^�8_��v�wz�] 9�WO1��g=�A�<�8�Mm�T�I2ˎ�g:�h�3�̒����Z-`�������W��e����XZ3�-���s���o��C�ٖjY'���߈�!�!�mp�ܰ"���"�^W���z��$:��j��U�(��{��5&�|�7�!�4#�9�}U����ӹd��,o�k��6]�L��˧W��.�^�t��!�ՇhR�D�$�Y�bٔ�Au?Iu��b�S$g�/§�lG��
��̋��*@��(�wO�f�ec`=�¿����ljOx8��y����J��k(�^��}���&Z0��k��b��� ��/C�rWu��_����,�J����v������J�(�+mO()����X������&�S����D%Y����dSaQꋛ�o/��pO*v9��NR��Uϟ�$��A�E����ߚ�J��K)�T� z�����r��X��U�&ū�]��
�ye���L8q��٬%��b���M�ea�f��@(�c�|(�yt������w_ʅ����]����T	��Љ4�0}¹�@U[� ڣ����$��9"�JK&��@L���IȕQ�l��I
��FV&o�v�]��8��N�`���%��m(Iq�%��7k7XX~�P�����q���])z�2��Tld�����Y1G�3,$5����ӂE����B��>E줅��QI�LP�rs\C-Wa����G
����1�ŭa�xy�0%�c�$�Om�%3�u o��_I��7��Ď�c����?,�z!�$��^X��S���Ϙm+eXy!׋JK���U�����Nc�O=�����Ծ�\�#��*)�E�M.,nlL�I��������
�'�T}qEʛT)4<s�D�m�ɵk"o@P{aE, q�a!�'uU��y>���fC3h�_�B]����Q��g��H�&�=F�}o�����o�@����&�ش�rj8pוY��
�O|C[��Z1�F���SW?~#���F�g���:��?����
�k}���Ү���Z�J�tX�����$_�;�e5DB&��~�ꏒl��o�Q���&7��!M��CK�(��V��$�%�v��C��q[�[4��G*�J9�?��DQg���5y/��>�gj��y�)�:���HN0���|N0Ίrmέ�rX�d��1�o-�0�U��G�ۦ�i�Bf9*(1��	�z�����u�r
$�C֪��R�j}s�ۃ#p$�
Q��6�Et�[�A�{� �l]!�?�X'<.��`C�u��[)�D��9E=�B��������E�n˽���WaBm��䩤zA���I |O�:�A$��o�̋�E��,��YN�)Kt�&��Qnd5�_�R��,�|l�/40wS�0xf��_tJod]���[x�ѯ;1��Qkؼ��MG�I�&�ti�G�1��h�8��k����#�� PF�\�p͖�(�����]�D�-�m��ƺceA�̿�z9I,)2��!r��A���=����8�y�h;�璞I�XЁ�� �x��*�r�#}�����ȿ�$��
E�@��iۉ���z��4��Q���=866�R�b�.��I��9�Сآ{S���5Ŋ�-c9��{�*��&>�@���P��엪/� �L?[�T�0�u<���]_��� �I���Wi�仟ګ�!Y�c�96��g?����J/���F�ɖ��dI�B��;� �3~&c��9�O�5�7���W�%>燠�Q�B[�5	K_��lU�!�'jt�>����:�T�z��\�jT[*B̞�,# �7���{H:'���dscA���~K����%��&�XxП���}ȼ^e�
5�e�E�)-�
�U^�I�U\�F�<�s�Ѡ�8w��vL%J���c����F��oCT��F0�f�%䟚erB]G��v=�J����M�>:�8�n�zU���Tc2�'�N<r�.�dA�tB���1!�$���ֿ�<��]-}m��
�&��e ЂJ��$��9w��:���z��ec_ T�h�Ό�z ���8��5� ���tDvp�j֑�ˎ���Dqp7b����� �O����H���t�O�a�^F�s;���
"��%C�@6�-��ˈ6�K������g����FP7�	�xp�I��x�0���0�����!� �kV !��7� -�<����D�9�X-���|׽�m���0�;�F_��}2�?x⣷�5�~۟��7����a���el��aBX��i{��%N��f�8�H_�yL��G�?�	�n����-��n�J�̎��:.�nS��L����|G��/=.��6G��wʻ7l�Y)D���g��~cF>���VTU��q���8�H�k�GN���\p�f&�+�:�����d���pm��y�)�v��"ݲ,��Y)9�It���a��z�(�f�&���,!�"���#��,}��5i}JO������t&X�n�(z��e
l"���,��P-ܽ����x�r~�$���k���v�y>CL�3�M[$3��q�rN��ָ�O�H������En??K�2,�|^�T�zE,��!:�0�.M0���.8#��7�TO��a!�ӧ[�ci.�%|�5Q����Y�d?�no�%b�>t�Za���l�X4Qx�NԬ����ۚs���&0�	�"@5�o�@͙�\��J隚������N�WD%lm	!�>�P���Y�04� v��ky9��fK�`/���җ��`���	&~��r텓rk7�P�
!��>�"T��EMa֮�f�>�$4R	�_��4 !JU�6�-?C/u��־tɁ�����jE-a�JD�b�Ez�����m%���J��?���:2_�g
���"�Lp^_��l<����c������Q���b4r	�������Ƶ�h�p�kz0}ŏ���q�{����hŏ-� �Q�OX�ZZ�׎gJ�H��
f��`wH���3���gW0�n�Y%���ū�����i1�5��-.�b�!���h��v0,��ƿ��{O����;>$�����,��2f�{=�'O�;�qq$�#g(�C6�[��bJ����������\Fr����2<�	b���F��;5�t� �l�f{���C�A���'���5}Ww���1v��{j�}�	g�8��r�F�����T�S=g@v��n�_D���=����]9���PWA�Bff�i4�兄���ot{on�C�&�Nap�z���%�	vu"��t�?~�$��"�TYF~������E��d��(>-���{�[�0�`��'��5O��=�	���h��Ҭ��j��f֤/�]X9�n�k+!ˍ��ɌD����8�u�-���N#J�KZ@��z���R����fd/*�}�h_uiQ��*���IL�m�S��:��m�m1?�[��',nbeZ��3�R�c�*8�e��BE,T}�j:�{	�}�˵�S�/4n-ҽ�J65q�}>���%�Z��R�\�.��Z��n���[k����[�J2(����%"\�AA�U�?���xW�Z	�HT�-$�����%	+�����a�r�4W-��rx��.3?���𾺞�T�5M�BOwC��w#�Ǒ{L�ö�����:A�����C��/ŀ	>G^��bT��J��n��BP�N
s�oR�E����:E�k�UO3�I���_�9Le����'G$Hhl�Z���3g�w�)Y�y/9��d�?q,�+C-^Ӯa,V�2&�A���7��~�\�	QƁLI�ʅ�����~C�$���g��&�8��=V�2A��h�<F^"�3i.EH��i�B�5j��HB2ŒA�S�����P�Ot�($O�B`�㜍�TM�:TUDJ|��1������ii0�uR��D]���p�G4���;�/kOaU�b�L��q��c�+7�o�GH�Y�Qw�P�7�>�� g�a(O��f��k�7�#�����a�������J�fZ:��8p�i�A��~��O��	�B+�e���FBK����SH@?^'3�uX, G��5�
ا��vPman" ōh��t������-kG)�f�G_�S�����	�e�� �ݛ]�ؑ
���K�^�f������V.1o#�f��e����O�[-�ç��Lҍ�����B�v�0
K<B��U���2���4`&	���?y጗U�[4�{-��n�������H̸�`�*�ħ<r��4��q�h!����O����TS)�J0_���=�އ�}��G�a�0Q�JPC�k�ь˽��
�K~�������xa�ߖ��B��Dd��b�#�n�쮓$���zw_��!��:�h�<�W;X���,�"%	Ƈ|�uv63Нl&'h���i�����I�� �� JV�2bV�.�qEg�5���n��9ӦCUT�#,�XY�4/�H#c���C}�?��QR�4�iĸ��S�6���ݽ�B.?���(�^6��6g����ҝ��;�ChR���RM�N�4/}@�m:���?�����޾�����_w�-eޘ^�ɹ�`�,�����JR0TJ2 �UͰ�z��K�ۖ����GZm%CR�nB���,i�$We�f��#�J?�0��}��ʞ�ly��)�XY=�}��M{';�մdO�Oɀfk��sp�c��ñ�K1��,WW���4<��p ���Y�P��ug(i|���������uF[m�Pu���6P+��6@�Z/�����8�[�c����~B_�D�[aȩ�d��@��J��`��ϖE���<�������ql4���*�r�h/?`։�h�/�m�ɝ��+$�4�K�z�����K�R�*�f���E���]���}E&�����?R���f�1�&�1�K� ��u-ܴ��>���%��{���.�64�������R�,�M�ǆ��TϪ5C���R}����%��ƹh�IW��'&oh[t�z���1���|ޗn`ǂ6Uj�a���i�]�#D0u'�N�N���lG,97�IܾD��`�=z�����R��Q���9�=$~�$:m����W��Z��C%܂ߓl�9B���de�pҝ���E�Sq��_@+�T�ͱ.vӜ����3Ek���܈ ��)������� .z��#<�lLg�h�I]��h�~�xb:j��:=��,�3v�NW	�� v�K��_�ϵ�,���_)�p`&� 7>4O0�k��ZG�h��,��:l"��wA��Ul�)4����Y�x�����渾B��7����9
����Dַ���]��҈�7X�5^��ٚ�"W;�C#�ȋ��[	�M��������m��5'�G櫟2�9(Ml��BBkv�2ٮd�E�:-SB���0���~y/����P�� �٢�WHݡ,F�n���sp�;4��I4֠�V��Zל9�v��^�����6b�z!;����0�3�q�Ux>%�>�
| ������0G�=��OD5�6���Q>����y<5M�&P�q'�b�J�e����#\���ʶ�B���a��B8��@7����4t�9�
P!���TlO>��JY�)\U���Q���,���3��緸�("�rx�zIғ�T$���M�ur�Ҭ���Kr�\\N�	���w�KU`�L3���Ӎ�[�Fv�H�E�!����W�E���U��;�z؂(*��Y�%B�%���p.��A,~ĺ^	W��+kXpߵ��<���	��L{�K(�goy8�� ��¨V�f��1f��_��N#����5he��Q��0_�����@^	�hKcs�#�-��'�ӂ�:Q�G��׋�����SM#�5}�%����Ə5���~�_�П
S4�Y6�>Z)�)q&�@l�D���ӑ�p�@]k'�������`�6�3��ݱ��V���@�ͤ�u�'�j��x���>SgW��\�}�y�&�oFrn����"���pt7�Ђо� t��)ܪB���jE�wn�d�R�e7�R��j��Pq��e�'����[w���� �e��_}�CSFn��������~�_�r��M��{�dg�����4�s1��o�"Zl��/�S�	y��B:<ﳀ�kZ/OD�~s#9%[�_M��E�{7�m�K̃����=!�,f�E�<r ?��D�?�9&��\����el
9yRe�p�օ�s��冥T�t���qՄB(A	���5�U��Sې���r���k�?�i���ؠu�F�eh�Ă����w�=F���QUY���)͍频y-tK-�=Ĭ��tx��K��uiW(S��Cm&!��'^���*ΔZ�
� ;�WxA�.��w!�P��1B��b�{�sx�R���2;�)���Q���yUc
�t��]��4�,��B�`0�3D����WW��\	%�i�x���W��5Z���\��(C%�ë2��2�W\$�0ܿĔ˶K�t��n������B{ =�a����[�P`yB�݇5��ͷ5D��@zW���Y;b�2��^��J���C����lh [6,V�x���Rr�up��$s$�r5u1�lުс����1�����eB�C�R�ԋ�@����<�b7��v���~b(_�+p.&���?bϐe��ȝ�8��V���ti��(�X{KFun�D����|�+k�X.)uE�e�vy�}7�(�h���<D.�P>|�EQ��g%���M8�c\��ʾ�C�Hc����jV/��!޽6c��S4��$w�RߜQ�F�tb�,�v�~�_T ���l:t7��Ά��	iL�Ud�YǕ&m�v=ߑwHq�R��[A���=K�����6?܏An�t�"��-��C�5G=m(5~��`����h�[�P@��=dg`��c&�&٧	.$U|1�xLXu_l����Zх��P��V�G�42���BJ���Rˍ/E�������0H;
��9��6�B��x}�����X���V{nc��pB�x��o#&Ż���n��� ����R46�>F]�l�>��I"��{�7}��� �F;�ޚwk$(l���߾�޽���uL{���I1���\j{��;Ȅd�QO-��Χdܨyv�@�Z<�t8б����Gb��F����oB��������5�ǈo�L��m@uD�o+�D��G�q�hâpK����$l%Ll��2�e,8逪������޸,�M;������I��M:���1��+]�'�߃����Bb�cnw���F�v��Bsp;'�����秧��,�MTF{�!p��0a���'���t���W�bJ���3�*e�H�[W��Ĳ�]餬HÚ�#B{�V��+����H��������y�9���n�-R�s�H�jQ��gg�H��g������|H%�������_�Y0�p���oX`�����󄒜|;��z�/S�o��-��~�?Q��E�fvRR���Z'	V��vq}VG([��~��Ms������l��j(ƈ���Z>���*�~��x-�c���u5�x�7�����Q-	7����5��=v�*�|�^�\�)��e��k�|)sh��"�b�x�F��L�g<O�2��J\��`E���K)���;�8�Q�o ��b����E��^p�Cת� e�T�y�������z�{K��t�{[JrPyU�԰S3T)��BQ�Y!.#Q�+?��<��} 6l���
g�# ڡ�<Ob���a�Nr��=��
IfJ�Ϟl�3o��;<���p����y+��������fB4�*�7��`�*x���)R�8�3M RU�dx�B�E��&|��s��Cq�P���,��A7�#Ϋ$G"��]�k�(H�����.$�QN��u�H4gH��z�r�
�mpWWV-��<�Q�4-�HZ����6�b����&�E��gI.iᮑ��ߝ�$��KipGD0a���q���e��g��\,Y��{w1���թ���C	��|VRx�3�ߚ�ry���9#��en���lԸ����m����l�fGK��H /�{�# @7�炌�a'c)HY{5��]T�ƃ�S���.	9�.��4}w�ό�!g6̀ʹ�o޴��-,Y
v4���2�shA��,	s�3����d�؂řD�^�-Q�%�[�V/�0�Q%8RCFc_�X��֋k�o�����S f�t�f�!��7���H�#�8�������%1!���ęe�n[�R<D�.�X#/4Q�ě\y�c�v�HԂI�N|	����,S�f���
S�z��q�Es��\��5SB���!�f�tU�|tֆ�`�,��,-�3�bp����
��. ޏ1��b��n\��=�hF�h�{#T>^�@)��&���g��&�c���`1�f:,�p
���e����E4[�A�%2U�.��Wq��>�'���;����9��x��Y�|M�E�O-u.���JL���'Kmμ��96�1���M ��x̍ ����\
B�pit�gߎ��?�ww�sK�N�9鵴R)~�Q�����/��G�C��4L�hTG�!>a��F�f�0�:�Yy %��/4�&O��0����BEƥE�	ԤA�TYr���5���u����|��0\m�ԕ���c�D�q�s�T� ��n�sZ[�!��<����-T���t�ːV�_�g�����q�ELo�T��q:�}6K02. �>��hɳ��6@�{@,��	5,�#��h�z��Y��� �G,�^��6��슆�lau}��xԽ�&T��
*j�96�4���'T nI�,�{��5b:����)�2&���ot����-�h~Qa9�m8g�s9,�T`��Ϥo�s�c�C��Hj�:�o��4L�a������,�9�5�Vq��]!'�Q/'e����a�p�$F��	,x�\(�	
��߳�R:�I֣��m�fMq	!%�	��Hh�Oz	�X��� �}�}��O����_�Q��l*W���<�U�R�N��w7OhMg�	KN8�r��켃@7�iJqq���{��{�T�Vxr�P���9�����]8�Zl��<���I�i�tlk���������j�e�e�~���� g���ji���wy͔�`��)�.bZm�4f�p~?�����V�Ͼ|���E��?�Q���p$��u�.���
�a=fmX��&�b=A�y�zaJb�H� �RF��wR�q�"�B]�|VE��cV��&E<�&�7��L*�k�jI���,��XE~��^�4��������cQ/ R��)�U''�1�6:��wb�\;N���v�/�K�0G�tn��\���b(̬�bmزq�oT�`5XCjD�?�5�������U��~4D�4�] \��ǉ��Gl�g"we���]�q����P�	?�u��^���*�M�͙���~�� ՃG��a�ay�n�����%��c�5Wّ�GD�Ђ�$��n�c�k���S,}c��y~V�\k�gԕ-H3����#����M�r&,�:t��DO�'N�4=�?Qr��sj���U4�?K�$5��.������cKV���?^r�m��l���.�m�*3�FR	��
�l
3��;�գ�#�a����i��Z�������ZP3����ř��f
 ��]-ug*x-H9	��N�&�(d��+z�=Ȳ:�J1&�ۚ��6o5j�nٕ�
�t�&�Jp ;ьτm�G��7���~�"�r,GRoxϽ�Mx�?�E�%N��~"�l�ސ &A���F�a,aK�}���տԸ���g�(�N�;�z�T�J��j�2e��'1Q�D�[C���rՃŸ�
�
FY�64*�q'Bl^�ji|�k�i%�����!��f��XP�����Ɠz^��rr(J3��||u�t �c=�g��E�ePlz���+�WB�Q���ߔ�6X�/�psA���*J� �	-�znA���;xO�mY�Ue{�꫒^�P�1�Ɗ�(nͭ-	�`B(��
����7���Iݧ�����{2N�Xm�'"�զm�Bk�*#N:]��+v��AF���ޓFQ_v�
�*x��S� ������yZ�k�xuZw�r�7a6�1���sl �6�/��S��!�K����x�!{�YU�9ݫ�`E��l��5oa��F��~yL`}�����9+T����tr�N�r���r)9�;G�����s��#��}b�^�6�C��C��_t�-��q�B=�"Z.,&����}!r69�mY������O�G�BuNB�g]{���ܟa%��������Z?D�q�U��U'����L0V�����"e�bv�o��=�>�l�-��R
~"�i���;uah�p��Nh"�Nن�����|#��\���F�|5�K�u�#�E�3��*9n=p�iK�/~�̟0륧4�2���'��g����U����G�Dh5��6�n�_|�D8�TO��XJ'�j �N�&1Q*���N8���%'�޶ѷ��b�+!R�b�]�o=�RZ����	��2�ANK)�v\̞v��C$IiT'��w-hR�y�I�ө����T�|�ڔ�����~&i1����=n�K�?�cVJڒ�ʧM$��6^3ƫ�@1[���?N��a�˯$sL��,�Io�q�������QJ2�B�դv�-A�z���7�ݯ�t߬mJ��%B��]+���7���=�62���x��^����aB6c��9��ߍ�������(.\
�t�`��B�gp��NDJ�)QXw7n�gT��5�dy�q�Zp�ߜZ��N�y �Z�õv4c兌467��3cPm�6�Z�gݔ�����Mv� ԡ!�
�oy�._�ln�ū�{ަ{���9�^wܬ�7��޿H�k] v�$�l�V�=N��T�΄f2l:٘A���|�����lK|�ލ���Ȓ�~b.�����ۜ}��f'o���`Ȫ��[���$Ӡ���SmU��Η�'�2�'�QG��a`�[��+[`�?�j0��O�(��~ܐV6m8RG�v�eR5W��9�VK�S�:ŷޡئk�� '�-`�Y��!��xm)�žj�=��Pw�A�:i����H��ۊ�<����4ް�6��b��HJ��d��jvf���7R�
qg�E	#�>�����u>� ��	/.�_:�dקu�ߵ�Y8LUob�$�t��w��}�@�81�Y<"ʳ������4�;���Nf�$mM�LP��?��Ն�'}n*�Y@l�xY>Q[?"2.j��;�"p�D�����п�e���
j8����$��1��xNr��N��=���e�!�oa=��)�9��;�p��xwĢ�[e�t!�<�v�g�������%�Δ�_z�io���X�51����  ³�}:t�D��i�{�˰Dwki���E[)�>bz�SS�+^��x��U�RY~�����0q�P]���6�!�J����
�#-�}5:���a�W��?8�k1�)�/�8̟��SnL���*���<�>�1����^�1��Z��=�5��/�%?�����!?ԨӪ?qb?U��~�Z������� �����m�_�lݠ/:�X ������E���B�~���D<�Ɛ%K��Y�a*MDdk	|5)ߢ�����jk��N��s$�~����;�@��즀���L�*{��cCU�0�_Cn��	�S�++ �E�LcZ�!�A��փ�S���l �]ժ7�+f1��e�\i�F����vހKl��T
gľu��W�W�;q�-i�:��'|�^E3��E�$�JįY��E��|o�9����Z/Pm:�؃�@���'"��(n	�_��0��_D����早�%�-�BTqt � :T-6Ǳ�f�M˨���l���ޯ��|Ժ���R�(���� ���[p�E�����a�ʘ�U,iQ����m�3������mBp�u�e#�+��dE�Bx�7˪]�#���>h�l��U�^�M%�n4<��?O���q��Ȉ�����j�i9f8�ً�����E�M�oAqWŭ�P�p^���P�߮�T'��p�
,7�b7�!��1��o�M�1_� ��:�����>�K�dR	q�rӣ��N�Iقt�-���\��*�3�:�#*d<�2<��LS�13}؊�b'ڶ8ā_�-�tOBaF�v�j>��b�b�:��t���(��EY&O{/���ɽo�}_-�J�#�w[U�xy� E�{c��X�.qn�<��i@,Pҳ7%{�	(C��f�8ħN�h%�3��s����c��h)*B��S�&�j!u���l(j7{��+�O]%Pd�x>p*ux���H�j_�̋��M2�}�`�$x=��f΢�� ���x�+�$�������W�z2�%��Q�8�����{�p�2�ZЕ�gDF9(���/>���#�Uc���0�dj#ڕ��^;������:az|�ܡ ���I��k(��¼��Q�"�:��]s����)���ܧd����u��!b�
qבqJv�Z�1Ӵ����J?P�MYH�����v�R� J�h�k�ϓrް0��c�k���(�6�����gʨ��x�N�W�ʓ>L�����2�%s�֕�j��.����֋`�P�/7s������_���r��̳ݰ���;Q�/���4�T���0	2�9x5��)^��K�)��#��F�i2��[]��W҆ti؞����E�X"�Lp���s�M�����w2	(��X�>��R'�D���u:���l�������j���
 �&������S>5����|uA��뇋��ǎ�B['bUZcA���;u��_�װ�%w�e� �����_����#�H�Ys-r��G�;?b�_鏔���P�Y�{���	CS^sF�*t@�nU��&V��O6�K�0t��l"ߤ�L)7��QB�_'� ��	� �y�idD������6�&�{9��ڱ�E/N$�#"hR��*{����PꂠO��mHu����J�"/$˜�I&hB�|��P�K�sq��KLݔ�7!Γ�9�E�����<�a���;N����r��юa��3~c���t�<��6�)|��<�«i��ڴ���&��mR�~s�Bb����<.j�Z�<@���2�G�3頩xMc<�#�sFÙUa�􆛛_u��9zW��pI��"ض���3//">���a_���P�_H8��c����WJ��%չ@�]��$���s�|8��#��k���#%�)�t��Ԭ��xzT��6�L��ys�<"����{9z��h����*�_�mM�o���Q2ۑvJ��8
[�&u%v;aғ�۟,$�= <V��m(A��V�n���K��D��r�D+%z�%0#��(���i���eb�P�=����Ce��N��3d����q��1�ݩ3�$��>{�T		wg�Ȥ�$�Y�(��K�O]������w����g���h'۞F�~�����2m�N������/���a��/��Z(�Y(󺐒��U�r�]+?s�@0j�VU��4�yzk��\ǋ�� 2
�����*���:�������S#q򿒢a��������`|-�t�F���R�P%�+�,&Z}�#4�B�_wD���� .�	�����d�(��S����`����U�� X;U������KX�I���c��*�^52�#G�!��Ⱦ��"^S(��H�}�5�Kk��T��=[� !�(����ѳ��U�D�U�{g�l�u�=��`�OP�PnJKX4�2IuΝ>��䬩���˱ř�M�x�����)��F��*�e�r|�Ĉ��+-âq���3�ա!���p��y�����7N�<�҉rDCw]���غt��0\���k.{{<���ݔ���6p�����ne��e8��h,�
�B*�� 37��`�M�m�S�`y��I�7�|@��6>ܽ���-�X�a.I �%��8����C	�U8��_��,1y u?7�Pz����B��wniXp�6�A(a�� ��b�1�?�6�֞��J
"�xx>|"v[�j��˼C	 
�ER��"�"���y����m��Q'@�]+�ؗ����		�zT*��&�h��G�9���i#��0�|Tw�T�!�Nb�ߙz��k����PO�a�4��q|y>�+��?����©�o\-��4�H=KrI���ˮ�V���x��s����"_����^+Ʊu�$=58���8�+�», �晰b��~F^ƃ=֐�@����r�j�,�R�7q��0��%��
�d�r����#Y�%�����_/s�\τ���]�k��]-�����x�HQ�7�P����\��(����.f��� �������zI v���r��B���6�]:}��ڐ`�p���/$�JO��b���j_��,Va�)�% ��V��c1O�@�
B�/�0�N�d!�µ��$�an�m�R���
�֣�׵�d��n�V�`k�����#�	�l�l���f0��=�Q����0M�#�Bm��-�JA~����]2ˈzb�)קv�U���Z��}zj��H�S�)��ٯ
m�E|��%����A	*-C��S��P�Np=m*c��[�If��(5�})�|~��'L��x��U�q'��-00���x��_�t>�HT��Fo.���򑉘�<���j�X��>�vR}�BI��a����JKp"&�V��P;U�����å���n�H=)��J�KE�ZW'��Y�%3%f���p��u�qEĵ���� C6G��У��`����AϜ���'*�V�yh�	�	k�9D䖢	]���F7������4N"�*�ײB Y����D�k�;�� ��/�e���>�C#_{��z���c�[��H��&`o-ӚK�¹�:��о`dZ���*F�4���S���T����O���1(�%��x�tL5 �4I`�i��Ul���7��=�X��៙d?`=e����6�]�B���(Bǀm,m~�F0��}��
���*r����N>3f����d�H��̋�m�K�_c�����֧��ӡQ��8���pR?�����}O��{Y����{�H&��R-�� 1@_)���2�K�eҘ�%�ے)�����"��s�\��sK[��P2�ėC��Ә��[ܵ��ͽ÷^���
��Y㏽ ��B����J����~!�(&q�l���������?fD�<ҿ@�(�U^
dp�i�K}
Ç=p��,Q�R��Zi�>���l�{��{~�EԾu�/M�iR6�7�#KD��7Ѫi˲�.�)�2�d$H�c�C��B2ڃ�������@{��̳�j,���?�����==ʂ;��v�a���?cI���V��).}��8�tJ�Ԇi�=v��F�	Y�#��GE|���
�L ���5	�ޏo�j�{�����ی3lX�6����"C�� ��0�l#��	)�xO&N�;�_*��w")��qF+-����l5��7ņO<҉M!k�v��?�n�L����ⶊ���:����>a�@��.�lmS�f�g��X�.�:Mt����i�G�
r ��ku:� �ڑ��Cv�ϐ�ڞ#jc�b���C���K�S�od��&�یq�'��e�H�o�(:	y�s;�7�z���Y"�d�ns�?J��E�1���N��1qJ���/X���H��d/
cʙ|�'�W⪭�� 4�T��/+�|�Y����t#����g]��C0�
 (��d}jR��w�\�]��.RA}t;�ǋ�L�~���H�a���R-Т�'K��#���ȂMe郧|��&�����Փ	Gn� ��ߊ(<T.X+#��ZpH�ί	չ��{�Z���#k�n]�G�C?�啓�^�)9aҙ�aA��p��k�D� ����_Ũ �,�_"WҌe��[Dd�þ�^�a��="��]��T�x�|bᓶ���z{�{x�ʞ������2X:�J��_�ɳ �Z
('���@��~���nC?Dקּ���s�����g7���[Q��a��W{���5aw�i"�FM�z*S��{����u�4*eB�2�a��k�HM�c��Q���
��'�҂�h~i�3ZJ�S���S�^��\��,��.�_#u��2���*��R!�Q� f���J�Џ݆�j�`ƨ_f�Ք��X�9W5��L����Iq�3v?!���)GWc���o_�9�e��W�fHQWc�郉[M�DM��O�ЪW��� %Ը�ÑV�W裠��©�O�:�h5���R��^�g�O�ʹk*M������-N�'�i�!(�ᮜT��4u#�v����f4�H%� ��U�91t����v̛ku��q'����� G�0U-�#Ԣ��ً�^4}�&�������2K#�Vi])k������!.���]�%�����?��B��m����
��I��	'k��6�	��k�,�* b`��v�*+�z��9�*I�]����֝�v��ߊr�'.^���=���R���U��|Q(�G(���S�)�py��1����|jW��bI��F��cZ3�yu3%U���PW��+랿�a�q��z��L��;21�����~>@�n�_���hQS�0=�$+l5�t�q��eb%4��ZXݗ��c����[�e��`�=�O���{�$��o+wD�|a#��S�����|}�^�Rƾݠ�Vl�R�؀O�ܤ?"7�$X>T�}O�M�u��헂�3AU_����A��6�fj&��Ig��
2iK��Mo?���x^$���ÿ�秿���-{`N$r�,�S��K�����61?�� %BGR�mū���a���{D;�.�r�G#�/O�/i��껥k�5PO��5R����R����pB`�*t+ �S4$Xf ���A<n�5�z���O^єv�rZ H.q���M*����5�0�DT}��(F
��z���]�Co�j�M���R��"3�j"G�J�/����+��M���]�<��]JT.ҏa�}��C�z�z����5
F�c>D/G���e��E�sKV����x�� �~���z��G4Ø&�`���Y��U@lnS/+��OY8*���Hw�N _%#�t'uv���Y+W�u���E�yR�|�HiypQ��,,�,�{�����ŉ��)�ٛNx�����!�G+Q���]����]�땗�D��b���B�x 9bɢ�7s�H�3YȭΏ���]������ߡ`�A"�x��PtA2�#qc�8�"��!.��yԲS���`�������2�l�#����6�b޷�M��G�w)tA����u�g��d��Շ�{"��#e�H���v��{+/�o��"�����I�G�T_�Z�"U��)����c"A3	xW��&�|�C1�C6 �$?�/���)Ȗ��
���a?u)��QxG4y;VT���:]�k!�OєB�Pygc]g�x�V�;#�0�ʛl�I2�.��u����0�N�ά�4�t�hx] �0��{PW.��S?γ( ���(�۫t����ʜ)�����_L&��c���̣3�v~͖�Dp�X�Ms*������������q��=QT��o?C��x�~��b�\|����~��R�zX��VǬ����#+BQ��Px�gw;7���1�FT�j�����x��w��Z�db�#:\���� R�d���Oxx&��Tc��t�&[sn"�lG�-�j&h!�,Gy�cf���}�
��c-�3"L��`�Mb1�YI����eK��m�"��9�����1=!��"��s"������U��Ū;��-Ͻ�����T���?2�}M��+gf�}M��䋌�"�DBΰLޱ�I���k�'g���������	'?/�2�;�ֲ�&�����Z�������ߠ=�j~���$��
�z����T��j����w9�K/(��A�R�[l<?�޼�}̒
��wk�%����v�Ha�r�C?9�%���M��Swh���c��	�y�NeE5���j��h�� �T����l���f
++)�C��+˺���֧Y�O9R�����Bq���.z���+�j��^�OU�00�}o��5-�a�W�xz���G�q:�e	�A0���v�zܝ�c{:&�ٝ��ٺ�@tC��u���{�,R��~�\ �]mV��K��� |n�.�.e�/��D�K+9��n�V�F�W���`�)�1����l����2l1BR�c:���*�R���D.Ꮕx�����`�gk[V��	h��e�S?q�d�Pf
5�}7xUk,�̖r-�`��k�7�=[������ ŊOዌ�]i���7c���jJ��)$��]�Ơ�N-��zA�ssS��7���=�5���rI�XO�p�x��i����4[��R��R��e�;UET�ͯ�kh{9�L:��6�
��D�Co�&�f�NW-�u���}e��5*�RK (O����l��;�T�S�%�J�âz��'��$�V2|fC)$&��ѿ�ARN�뫪 �F��E\$��R�ٞ₱�?�K��1��@@{��n~O�8��!��@�H���ɽJ}���R�YidёZ�ه��
p�/+P1��˃%��P�.��b���r�R�5���4M�"p�R��C֚��
r>#O̚#���1�S%Ԟ[|`�Ϟ���Ҵg���`a�з��M�f;�D������a�#�o4?��C�ch��%8֮�3}i�>U�yc���?N�_���M�В�2�ӊ}��<���p��q�"�s޾�w�?'w�ѕ�2�G4���3ob�F�TvF���W�{����|�!6T�on����m6�^]��Fp�z�?E�.��=R�ޔSib�������|�{+��|"��Cj��yD�v��r����=�������D�?�td�r��3;���=H[�vظ��hr��aF�*�T�h��Bm���ܖ3�C��ޓA�e��ޗ۸� ����X�-?U�E�cE-(�(/RG�
I��h�L�u:y'׆ֱ�v�Ӯ�4A���Ǟ�r��ƞ�z���(�0�z��Vrg��d�;��1���2Rw��S�әI�S�(�e�����K��.(j+M�`W�Lƙn�*�8�,�v�e\���s�űT��h8S*�L��g���G�݌"l�ԫ�6�~y�wz1�2}�P�`Ϛ���R���NO����R���Tx#I������"��~rc�P�D���qy��=| fPǔ�DYh��&B�f�]� ���33��e���X����d!�Y"��e���]w1\���I���9Q��	�9�"���VoT"t[ƹ��Q5�Xg��8Vx�;�F��	ޙ�HY��Bv$����1��VI+����z�U����D�_��N�QT���Q�L��c^x����]�wǇ�Szcb6r�9����ep+ߍϵf����w}���1��L��5I�dn��I��'�
�b�$�{�����y�ЭZ#RáA��)Z/��Y���?��f�´����h�P)�f����H��@�S -M�Z�&R<�ھe!l��2�l�p9$5c4K��.ק�O�o�2w�t���h�U��ꛭY_��}/įu+O& ��A���0Ѧ�9|���i�U�!N�Z��(ŉ(��{W�y�r��������2��͘��@��$�Hڌ:�@5k�D�A���a1]	���wwV{�0�ۻ�����h0�࿩�C8Wv�h��GK!}ޟ�=����e6����C��?���Ğ!i��n��[�)ֆ�!�%�8�[��7=���	 ��[�����}��A�\;���O�j�z�-;$ N�����|�'�)���U�����w= /���zbŶ�F��Y�mD���YZP�øߏE�}S���T�u��jǅ�Z#�i���X��@0�8���F�ļU�T�S1�{�zv�m����A���Dզ9���Dj��W{$�c~~��W	[�g�6��9_Psϑ�1?��r����kV̼Z -䧗mb�T��OTꪟ�;�W�KNe_(/Z�~@1jR��:�=pg�KJ��-���^�b�|}�&q �Y8&�	�B��+�L�8��C%����H4�j"�]v� ڡp�V���v��0K�&;[uAK��N���Rno�HN
l�}H�k9ڹI���<��T�D�S�1�,��+e|�UTz&�R�c����/ǥI&'�TΪZ�]�����4�h�'WUi[�h=\�r�[ ���h�����Y3+з����^~%Ոҩ�s>�Q����׾�*��>]i�蔃��5]�b����.��~\���R~�i���t��k�_��F<Q���6G���:�Y���t	L�ԅ�+fv_�o�P��t�+`)�.x�Ӯ}�rb@���0���Bi���6�0蠨�0�l�z��`�P{^��m��Z�E�p���D�io|��w�	6vX5�5'�2	r�O�ā�6���[���t�X�hrEP�\��'���Q��ݦ��m��Vg�D�bӡ�>�#����]�:փ�L���a�}H_�hQ�t�|��c�Q��2�;�N�B<����%7���Q�#�g���WNȩ�	Sw���z�v�#�{�oˎ\��1;'���T��g}��`4�{0��A˩c*Y�wAr3ٍ�̸}2����	;��e^�~�I}'������U⑔q�D5�8���PQIKk�ԋ��԰����<��M7pFu_yҐ�2�E��T_3�����!�{��~5����΋ �W��E��x��]I0�r��,���/�w4Ʌ�A���DP�d�n�8g`dBLq-���h�Ut���س���saMc"��m���7�T���Dq9��7d��;K��dpC�tk|pe�GW��WM�MQ���	��аahp��Y�� P]䴋U�e��EߥX�?V�4��	�I�Ƽ<���
���g���O0�{eN2�4��m>O��R,��(>߷S�i�+���h��\&)���S�e�ż�"�_� �`�䨕�*��&��C���H"��@��@I*�Sf&
^AY�+�Խ{�h�w`��Z�����!�D�Ҧ�?�5i�~d�D��G��M��_Zm5�����W+��מ��D(5�BQ���v���X�٨2�?0ob�^H-���kW}���Y�8�5FK����H+4� ��ԭ�\
k���k�#��Ý/,T3�~f������N:��@38m*�`��@t���L�_ o���1á��'���1����&`�=/rl�-hZ:�T�+�V�+-��0DP�s|#i�6�]Z��Wp_U�q%��`t�=M�K�.~!�8 �Bw��k��Y����.�`�}v���L��V��C�S쌱OxlAv����[�/Q���%?I��Yݛj���a|��L��K)Z�	n���*�7ި�PYd�$�Ď���R3�5��bjio�)ي@Ǖ[���a�$�P�՛����p��8�/�]� Y5���GG+�����N��>���6}н���3a��W�;�)3��Y�9h��Ų~�)dȪE����߄��M��T�� _j(���bZ@Y�s����Ö���4p�IX�*/�U��?zPN%h��'(va�$�s:+�+������g��Y���9{��k�u1�\�������3}?��Q�k"F�{�h�k�: ��Ȏ�*:���7K��v��4���֯����.��0��jrYx��C���̾��Ϥ	맭h ��R���j3��Bv�=��$L"ۑ�= ��'���<�����
�� 8i��<�"�,�)R�Z �d\�q��U�,���
J	�e�?�!�{����+��2����y��8H�k(�]*��4��c�_�LU	g蚣(V�̓x�20�I�e9����h����� �KŚ�q�^z��2�%�f�����i�-s���+�$�đ�Y��M�/�f���VS�\vc�B�Z���z+�
�s����;q��M�(�=��l�*ny���rY������X�O:��vN>��@s���,��ھ6�X#3H�y�i�/M!Q��}�{)p�,���e/�cةm�uzxa��	��`B�N�H�ah������-L����=�MC����z�QZ��r����WHG�䴊�S��.�F�<���OחH����\*��R�8i���d~:�`9��R5;�R�\e�:�
�I�0���2�OA�g������=2������Uhv�����, A}��#�?P�G�����^���/�_�[t�|�_50������!R+&�Q��"�f`�¹�'���2?����(/�1Ò0k���wN��7�(z��ڙ�t�Tn�k.�I���A�9�e����)�"'Y}u[1d~5Sc?wB�f�~�$��F�g}������\���RE�"���C��]B����_��10�\�����w	y>Q��,�����4�Hq����tF�
2Iv�����^�#.���1r·M����9-�	{�J8���[B���2-O�k�9��U��G���E��Vς�G�@�S���4�5�n4LI
�?���܊mu^t�Ľ1��k���0���ʻ0-�9���)]u
�;�}t�<w�L��n�i�8nЛZ�����&k��5'ѫBÂm���-�:t�0MQT��F1�/#6|����x�9��%&<fܹ]���;�Ul���~I�HJg$S�N�E�w�07��O�������Bw����\Tm}*b�-�洯���n��˨�A�Գ�.H➴+}:������Qx��$ؕ!���8p�������uYl��AW�>�b�땙���L�F�0(���w9f��-����)���	g��ۘ.NA �݃���W�RZ�����M4XkO���-�d�ғ�[��_"2S������*���/��Mnf�\.+��� �V9O��mǒ�� &��-���ӟj�����ynx�Nϝy։�ߠ�fc� >J��Ad>.��d�+��A 4��Wqͬ}J�g�;kd��IB�@�x�3ܐq����X^迹�sA����B|��91��u�JC��ҶL��ZuT�|8��4"Y��y�@\�
���zU���)���E�g���S�՞*^��n��m;ʾ�����m�}n��.+�`��d�)4�� �1�����C0��V�����%0�$4ݹ�o	q�v�u`��w�0��&�H%~����Pc1��	�@ �nZ���P���T0�]ܤܑI�I�]�:����[Gl���cG�m�!����q
�oQ렱|������ڻ^33=S�u"?j�VMf�`�D:�<n�g���k�����\�߶�X�Y���#Ѕ��;	�a�r��" ;�PN?$����$�ӡ����ŠD����7dj1�BXo���TܱZd_��K�_�qW^�?Ķ�-���m�f��_��v]7���;5�����D���ᨥ�;��sXZ�b�aW�釶�p�ź4������-E����	�8��f��n�I�4H�Sq{�,\�9]���l�8�m�7LףG.�Ȗ��%Ќc�)Ƥm�]1�ʛ�=��c2��U\R��ڗw�n����꥓!|oG&b-k,���1��}Z�B7�e�9����l�JQ�,t��Q[�.������DmF�,��	f�lOf�1,�<�Կ�)MQ��eK5���o�R#UW]��f�ZU�£�\R��i���dI���R������Ɓ�c�Q�3Q*c�9�,,W��Cg-4�}W��,�|VR��J�=ɪ��g"����X��ic��������X�صn�]�c	��*���1�����cU����[�������	�������c�c<�7R^8`� )"M��Vq�N(�Kjc�bȍ���0��-PN0���V�G�=F[RC`���S?=\��|��%�F�Fd���YWrL�+���*��|�s�ou��L�>�U64�9��t�Q����3��$WI-��Բu��ܛ�(�}��e����pvӦ_вA�6�į1Y�x<B=Cr��?�d��ƛ���H��b�x�$��m���m{Ȓ��`?�~��_T[5�#?'A�e��E�-�f�TY������\'=H�y�u�;����r�W�4��L��ͺ��V�ջ$nOھ����9�>OOF�J��/�X�@����급(������O�P���_�k,"b�^$�tS(ߡ���)?r���F�[�Ў�6�X��7'�F���d���cT*]�u�i�u��m���:��6"��T����4����ָ����'\kS2	�Y��y[�O/�agw��bٍ' �B�v�8'��V���sG6R�mC:��
FC>s����%�AGՕ�9���Kq�=c[|>�/��҄KWCǶ��[#te�˿F�j�h;(��Fa�|��-i���Ro*��*�C�w{��e��OS���MO�� b�h/�7�x��I71/����H�����D7US�0ѐK���R��`�U����Bw6;\f��7h�ת���	R7�����|t��X4Xu���%:x�g�D� t�����T� W]<{��F�3�j�$�W�����!8�X
�H�	�A$򇊆7�ed!J�A��QO�m&�nY	;gN����Ș�:�D����ol���Z�ف`+�;����m���{[JR,���[��R���b�t8o�+�o�ĝY�]��� �r��f�Y�%��]��.�/C��Q�3�c��j�����¬���(
�P᧌�����.�6u:8�ř1v����� �v���}cI��(���A "�(��]5�E�l�B�.�ք:�8���ܩ���i˵d��*��o!�'�r0�����g�9�a�u
a�_/�Ԓ�� &`�K��\m�a�-���Og��p�z
�G��H���๰$ ���u	=��4��K�)A�PG��Y@��$/�C�nk�.�ɋ%�ǳ"u��U�ݞ-9�GV��豛c�)�����"Թ?7�6ꢒ�;�M�l#�CO-�������+�.�M
��Ճ�;G���T��pd�!��kI;K��(��ߍk})ʡʙ�j�-�p���p_/g4��1�w 
��!�~^�=7LEI�f7������.�<�/�Gs;��,���)���G���$L���"*/�M�)\ܲ���9d3��2pNdjH<���/J��ҵ��f�I;w�:"��#��j�3Yє����_�ț�
���+y_�>�M�ꂥj�0� �"	�veD,���H�E���Ά`wyZ�x"{4�]�Y�~%@V�_��0�
nZz���IM���[ܣ��0qsdr�҆�r��M�HY��,oWO�
��P@�*�P��iW�H��tN"MLGG4ڹB�4��-���4�%au2���l�(:Tw�#��=�Ǝ�Kv�`_�l�LJj\�������O9ލ""���x��C�E��K�&uC�y�nEV�G^�� پt(9JC���z�'��uǝ{K;_A/�u�_��|!2�Y�EJ�{T���~l�T��"
_��Y�fJ�6���\�	
y<��<ʅ�t��B��} C�`��H�Ě<	�R�X"�,��F�%�vF$��Lw�\�8Q�c!�|�o��3
��J��ܥ����teCmg��L�n��j	��}���+\j�wp������O/ն�mB!����ԏ�j�9BN�l��z.	:xW�PY���,��w~?&aKI��/'[v^!?1D֛�z,�D8�x��ǝ��b���[X���|�$&4�b�:�p���'S͝@��]8���5fb�$�V��Āuo���s�p��a�C���Q�������H��v��DޠC݌OA/�q�L�'�$�M�؛h�t>U�\��,�|{�O�	��Z[��4�v�%|{~����¨l�=�f��a.K���`l�3�T>�{�f����
fk�®N����-ȍ �#x�jL��*;��t8�pl ��y�������J��4x==��ewq%�q�r��K4���穤���˸��$$
��#d���,� � ��Z�8�U�i�m�iM-��@�1�9;���T�ݙ�b���j�H?.Ɵ�%4`��2�0p�! 2|.au;+��`����h62�H�3�(b�=�\^�#ɖ?>�s4��C��^��4>�!��s2@�H��@d��G��!sP�+����TR^�	g"A�S:}#!60P�i�TSB���@�b�y���k� ��,e9oA<L�`xIhأo����d��I�W�F'A�4�5��TO����݅ٝh�9F4�����-"�h�l�b���gF	� 1㹺i|���jGV ����џ�	�Y����G YY&s��72��)�&��fIP93>�5}l�E/�.������Q����3��i���zw��ԏ\��,���{�,����R�V;���y�t�x�>_Z��NKہ�^��#o�-��'m��O�}�̶��ॳd���Tg���3����!�Ze���jeY�0
���b� ����5T��Y�����b�f�&+v�=xp��R�T]tSM*!���T	J�-v�x咔	�)
��h+b�x�%=����f����!(��]�ܣ��U{M�|���ӄ�c�
��}4��1n��E�V	�4,`L��/,����RNe�O>�;R�E�>�2��E�*� 5�ӔAM�&g��ػ�������2z\�*ԝ���k�Z��xch�z� #<�<7sp���(����0�])!=օ����QWN!5-�f���ꀙ��r���4K�ikm��'e�y?΍Wt�4��Y��}��`���ɉ(��ޙI����#"�����yϰ�>�2���K:n<�D'�*�M�f�t������� f���G��R�D��P2M�����P'm�3JY$ox�5.�ѝq\M���z�68�����y,W��(>�k���F1zT��Y��V�qL���6`�W�p����J������J�iK��z`�7�d���;�%F��1M��=�`?JC�U����A�WA��-�z0#��<G��/<��t��U�� H�lxF�o.�z��:6Xg\�� ��aF	obQ9N�"��y]I�w)��N����rY�(�AQ��R:������ \�)d]S��Rj�&,���T����=c�H�S�F���Bse��I>���o�爱,�
��&B&Y�g��%̒��L`���������c�*�������mvڿ�:����B�ޚ{+Ki�%Ҟ���F�?���/��H����V�i8�B�\�c��Cʝ�"�J�t��N���hV��Q��,�.���Ľ���a
:z�3�g6�Zn���e�C�l����� v�����}	1=��2D���k��;x]��Û�Xۯʖ|�Z�!T�r8��5K�WD��Ӄ�ΐ�{S�29�q�1��̢���'f�0��{�,x�ߡ���T�f3��O���e	>�#��̓��7��ߔ-�c;��4�ܟr�P�E�e#�7�11,as���a���"�	~��Qbv+�����-8I�	�!LR�BC�2�e�#�D��@u	�z	Կ:����=Ĳ,�U1�Wo�e?ٹ��'�Y�u��`6�eH�ZJ�{������EL����K�Otᯠ<�@V�*l�@�Vdv"����0�Q�_o˦ɱB.N/�f��J��]R�ޓﻥ�0z(cM��;�|���3���|:m�3@��)�`������ҵx�η�{�N��F� �NWέ%�R˩j�f�k_B�E�G���� �.��:4U�`�Y�\��ͯ`�� ɪ><j��e}�v���Ď��~1�Qo�:�ጏ�mW�n���L�?`̂����H�5��� ����7�h�l� ���3uB08͂�yj���2Ȃ�J=��Hn�@�T��+�|��X�%3�����L �Aћ��d�����R�T�L'�]�a#�ZW��ܭ�=��݀Խ�x}�z���}HFc�������[��� fA�(�������uY�����a[�7}n'��L�Ç�L�E��[=����J��œ������f�~b�g��<\�\��d�a[9������S��c�eb�a���t���/T��	�%����������Wcs�< /%nʆ��G摨^?��@
>H�V6B!W�;�ۛS�U�q�3s]�����X�i���sl�/����n����\�R�6��?�D�K�lm���-�gk�v���h�˼��"RH�7ا�Ts�v`$�?�jq+
9
�����s�T���M��U���P��P	0�Ԯ��*�.�sη՝̒��K/[B �"k�l�pi߰JtI $0v�`C�5��uģnz4��<o�VE���k�¶'t��9X�oZlt�OvZ�pu	l#���m�{����F:\SB�/,�c$���EJ߄fH�|ݾH���|	��*aw�sՖ�x�%�oC#9,
k*t�"�b�3Ƨ�=��1՘)Mo��ap�oC��Β7F�x�B��פ���;es��A�DI���>��n�	����57�/��>
��>!o���d�ۜ�!1ˉ٠��p�E���}c,�~'�@�����ߊ���镬c�}��K
��-h@�`�6!e��#\0�6B�+qg:�)�[e>A�R��[�R �(�;hI+���Y�	�7����#/G���4~)�����4%��k��-q�7 .��0V��;�Y^
�eOn��X�@�n��_#����"�N�Fʪ��n��Í�k9L���i2��{L��nK�������ruN�-Y�R.���U���9hpa6NDs:�v`�wĪ�D�V��p�����b�I�k��:��i���ֈ���7�t��P̘sS6R��=-w�m>s���_�9y�>y�����0��~�t_�&�J2_"g��*�~c䠲�5�E�܉ c`or~:_��#OuǴ\ /�kXo��e����%$лpwG�!�"6�6��	�sv/��>�?�*9�dK��}�>��oKI�b$�l����8,n;��[���UP�e�#*	�]̙�c[@���U�/BvO��qmX���S�ze���R�� �eM��A{��G��Ӝ~�QL���6�:Z�&�H�b�Gy_��Q����<]9��*���;�b��3�|/����U��t�gX��� 
Unܙ�10�r�|9\�1C��E�GD:X�<�����Y���ͫ�|u�q���o��$�`�I�����b��n�!�\�1��!!_N^$Qh�w�v�y�ى ���Q̦��BJ�<��S�[S	��	R�C��D2Ǫỵ.3�:�S��C�`0��t��̌�*n�7�A� ʷқ���sE�1�(����C����0S��Q��+ƺ�+OPI>|0C���s�Zs�-Ԓ��j�ި��#�8?-�q&��D��k�x���=d�b���.[����୐���D�8�9�޿�ھ	��c���C�=�ㅂvCj��U�ɸ��\���;�t��)��B_�ђ�B��=Y���U�'O���3K� ���[l���E-�Ő��lc\E�՞�3fm3ň�7�����k�0:��K�_͞ݑ�����dTNz#X�1�0L��;����ӍXB�`�ǜ�Q��3Lq� ��)�_��C��^$��Y���ɡ�m����]5�V��!��;�I����l�.�t^ql�epzB|��Q��G��1� +P�ʡ�T݁gx��R�#t�D;o���Fϣ��(�Y���$��mxmJX�*/�:[�f�׸����o�;���$�mO����(�������V�d�ȅ{i
��t�ƚ���&G�i���9�^~[Mv��DI��G@[������#<;}[���2FA4���;�0�u���p���=Z���w���z��q3g\�HW���ɤH��L<��j�Q'qr����M6���`���[
t����h�#��@�5rG8G#�K�G�e�1��~+bztK��)���tl���	l���@t�}��Z|hi�|���(Y����ə���n_���R��2dw���5/&���+��^�P��&������:,����˭yʉO�N�Ӆn���a%���/M5�xEH]��?$�Rr�����
��?=̡��}�<f$p|<vMd0X���]@�̱h=g���z���=��Z]������s��x�S�;c�{��뇝�M:H�%�)��m9��G�Nb����(D�i�����ć��yj��7�V_�ckh��������%�٥*31>.LEϸ�q�{�nyv�m�3$��6݇��I�i멮��pF.�{��p��>˲4�m��I�ތ�i��?9�:�1�%�6!fF���G�\Vo,5����%Q-#+�9T��>4_�=���?���M��7���br��w@�E�2��߽f����/#�3�Md%�6?��0.��`�������*I�&�"y��
ZUJ��$�=Jʗ�0w+%EP���I�g�6X{�S�oq�R��p*���2�W��ˏ�	�4���i�h{i���8�8]�HͰL�c��Zr1���&�/�ut ωIK��k��Q�,�djW@7o/a��"��ƵV=!��&/U��F���ֆMj����5S�&	���]:\x���֒����h��:Us��K��1.�?�N�V%1r	`���^��hp܍DKܖ˚���'�Z�6*�沸����:q�)�>����l���
:��D���`�rW��]�+<:cDǱ*eMh(�>K����&?>�y�}���7_J�5=9��	�i��u�,��_��~���Xm� Y�h��K.,ղ���w���lM������C��ϱ���I�ʺ90&K� �
��艪����{�¦%T�85�-�׃n~:������H��_Bv��6��%g�e���)UOL<�"����g���HW��GɁ�ॿf�7/?�!yG*N�8S4e�=�<��V[&��3Y���9�h-R�)�]P�[+L"�e0��G�Ɔ4盐�E�(S�=��ܥwA���$Fj��$A$�@�3i���CF�	���S���̯Eӿ�i}��'��WT]'�NQ����1���e������s$�.vo<V��D) e 6�
��9��Pn+�G�؇s-��?��q��[��k�'���|w����v5�Mm�e�u����h.T�΢�N+�ўܵ����)y-���&�-����[�Tg����(��?�aB��{J;.�;8ܳ�N�F2Gg��ް��E�´����W��&ݖR/|vA�o�0.�O+���S|�)O\�m���}�B���[Fݭ#�"��I"�./��Ũb��NI\��w����px�%���0Xh�آ��͵�zRC���F�σ T�L�tk���>{O���SW�-�u1Wt��y⣍ER��0���9�CWMV�%��bǰBf���8��8���[5���������h[�^n�Fw໘�$x�)@ҵՐ�Ʃ�%w���m%ٽm���e�i�L~��C��LB	Hn��|*Zp�q����2jS��G���@A����8�c{|���wys��yNet&��>*)w|'�[�BA�l���\̿����2�[���� �'9�.G��PY�k�S���	ȴ�eZ��4I ��V��@���W�X�8Q�ߍ�@�Ѭ�,�'tP��ҾQ��t���
��P�?F&��@���j�c�{<f��<�b�P�~>�ܚu.�<�!�v	/Fف�C�?�~�y��t��y��d��o���|�&.{�ag/�G�q�p��Nɪ3%g����>FuZ�I���8� ;M��A&����tW�V/�wk��
)�n�l�1����jR�y_��Sg��>��l��-��U�l$T���p�0ֆ�WrL���h h�C2�g��R�U����8w�;�ַ����rAo$��q����k��� ��׮+R�4��R���$I8�*��k�)�f��z�m��׽z{`�4�CY'���o_����
�/'�23�!֟*���z��n����+���l����3��U!G���_�����0����(�Z��A'�"�wbI�=BPH�>�^��3�!��"��g6��\�P-�����j�s��\F���F� r�`��>x⛪oI�>^B�
��Y)�m��:޷���`:Z��4��jf��g�?��\�:u<J����ң�.p0y�>�����u��F�2��Fw�o��L0}���z�q��l< fvו/�("�Dp3��u�����+�P6sKso��_G��J�N��:#���z��*������1U�._n��$I=?�Vs�#
�������RݥV�e*S��B"��V��,1�j� �p�YV��r/�J\����ޙ�FB�����O0��e�L����;_k]_��5:�f�X��C2�#=���oS����	ȳ��F�a����.w�x_ H���l��;r��]D���~����F�>�z<&���a{���Q/���ՠt)ǝ**�8��b+/����K��:+�Shڭ����Bv��At�	{��SC���f��ms�g��Z��^xDs��%䱋q�}��ήM�M��D�����]<��>��_�� ���>��|�r 	!�&{�0�p�j_qR���S#L˰!����/̎�V��-���a�.���,��	uc%<섖�9k ��v���j�_�e0Q8�����"����!7ȳ��0�fdEs�U�Ҝpg�յ�iE$d�YᢋV�Q��Ϡ���J���.�O��咯u��N�Sk�ﻳ�А��&C�>��n�V�u��J����vx��u��ka��8���	���O���[�I��0�v�/<� �~Ձ$e�p�岈�����C�[�w�Փ� �R��ηɲN� �Z������'PG��[�e=��%&�'
GmV�:��3�!���M���z
��M��{�b�=��9�dx�xޱj��S��#5���K;ܽ/��,Ku/�1�i�]�9�{H'������9�|C��Ϝ�ma=u��"�q����YVk�g')uǍ;ȧ���j���f��/=v�40�����a�7��/�s�b	ϓ���nŝ%4V�����t�*��Ʃl�}�BE�'�%)�̴~����Z�}��dL��-�?7�'��\`��a�Va�?���d�d�N��'+�F����z�:�/k�j{dv	��Lz34hΗ�SC�F��*Cʕ�{~�g�d�z�X�.@x`��~�{�Oh+��!J���ڼ��i�J�Q\���x_��Q�CK}���)a��=�j�ֶ!`)��ê�O*(s���r�_�/��S� �[]���"r>���-Hs��:v���	C��÷J��b����=�|�vk��w�����`ci�L�m�&+=5Wy����S���:qLҶa�jN�\?�M��r��?'����gל'*y�~���S�����,ϓ�����(Nƍju��	�oϤ���Ƃ�Wf��!�,&^{�&_���Z���W��i�'�G4�o˃&$=�?kX�J��F���WO���qϳ8,���������DW~�
9.�2��ҙ�Wg��M�*Q�?K�D7*�<��w��T} �s5�S��6�赛��i�����?@5֜t��cp+J<T��+������-�7�^�?�/���.�R$M���|{+<��SU��F���¡!0�. n{�L����������6��׻�$��WE�ʋ2� �4�iy����E$�C����bӦsI��e4<���B%��vKT�dMH��"��`#r
T� jWGL��^���gt�b >��P`}���S��9,����\���l�E�!$z �Z�Q� � �~�Z�@C�Գ)���-�MS͔�s�޳v�e�"�d�	ɋY��O"�*u�-w�Ղ��;�n�k�����.̼����O�(
;�,̳M��a���}�����GT� �Ye'��_���3�5XM�ds�:��K����I}|�8<0{�D�z�R,"f�n��āW��ܐ�P��x1��]}����LΙ�j��q���yĬ��G�h<s�r�b��e�WcJ1PE�'��%�ө�aʗ�B�|b<��:��r�XѸ5��{�8�b�N<�=�,w�`)��Va<�O������q���n�@\��0�»9)(�	M`��wL� M���P�ABI�|Vc��'��V�[�����ˀ;�~I!m&i���Bs~ܒ�%5�2��R�"��1B<ض��F'++%sT��5�"m�4�]Y�|��"y��xъ��g
�Z��_� 	?���"V�Q�%pWX�5��5��c	� k*������2��Q ������wh+*<����2�W�#
�6@���	-�>�����s�R��%S��|�C�{=��!E���W�y^��O�*@���Ƃ�`Y����Q)���s���K�ķUѕ�_BV�m&��K��\�W��uq�#��j�z��|��g�M��X����׊��aK��!g�ߘ:�uO�֗��)��� �Ay9� �l	��m%��K��&����:cA휗="��0��%֝��Gy��Hx��zf/Qu��oo1����3{X�����&���S+.x�6jBqX@$8�����t�E�Z��b65��?'i��G�|�&S����f��K& 4Od41�N��*ʌ cN�떻�}r�~@a�3������f�޸Y꡶��x혬L�9�2��ـ���׸�#H������)�a�G�Ԓ��@�/�����W��C?p��3E#��n����&�(3�b���9�	��ۚh�����h�Pi'8�k
�5�l~9� ��ь���GG��m�'S�>h�N�VW���;���}eg�/���i<Z��3-/���W���Օ��}_�ڃ�2 ]��f�ԉHNϏ�)�gc`p�i���I❳Y�<.�<P���ߦ��;g�G;a����EB��г���m.�Q
,���].D-��t|+�|��K�*�ؠ����c���T�|?;U o�?6�G���B���־��O������L��no5�\�&�*����,˰���.�kh��+�ӫ
;���Iq2���n�l`��)'����V��?�����"�I\��7؜���*0��\Eu>2$k�Rų���ѠׂTmY�}`.W�k�)�����}�~��m�OL�mM�u ۡNб����3��v���9�I��F�-!��b.�;m�1���t|1�l� �@�i��-6b?;�Rfam�W�o.����Wi�����;���3%�c�����]5/���wO MW�������;�[k�A�!��u�G��@6��M���=�uM;���T�N��i|�O�S�
��a��D`eS�ז��B3���7�ԏf�q��H�He�K���xeS����mzs
\.�3��4oJ9������ϯ���p!�ڰtH4����U]����JD���׳ڡ{�b���-��f.[��k��ۛ*��dOb_�s�5�k�ӂ����H�\Y�1E�B=<�*;ʴ\Y��5�2Pqr��Tⱴ���d9�L
VY��(�ƾ1�5�,�%�pTz$U�m���u3A,ۢ����乒�ax�B�B�������:���Qϸ�c�w1[�钼e���R�潈{��̛3�%)̂���6�T�<R����ٞ��E��uN��=���w��KT�B��j����(N�|���*�>
��L�[H,��|�9�]��xzͽ�q�Ͷ��'�z:�q{���k��	�Y]�v�!'`$
����K˪�i&��~S�﫣�]8q�û���I4=��4z�t��V��^x�˾Z^�Z�'[&	[�8V�[7�.���(�QNX�:�u��x���9>a�fE,�N�rܘ�)�Y�0�Z ��%^m"y�9� �	 �lp;��(Y�������9g(��_!�����9���yQ��i�5��_cvq+G�[I^�f ��ɘ�՜@��'}4L����U�C(9�(]��Z�]����H�@+��'0Z;n�8H����&�����2�H�6
�
��aY)��]�2����E�չ��o=�g�&U�E*Ŀ�z��'XD�d=�gj��E��i?�n��p�N'�y��+5����A9�������!1*�3 �h.���V����vλ�Kʟ�*4)i6Ŗ�_����a5
ln�&��aC�|~��W�RӾs�p��Z�|)��d��������(��\��=��5�^5p�h��4������Fb��5+k$�3���}nn���q�tKM�X���`Av���-e������Nr�[��6Y�p�M �����H���}5���O�N8PD��"���Q:���?����S��-���@<���>��=Q0�<��-d�"��'#�Y���������?�B]���^&2�9U˒o�g���7��xD%|�$�Q�U3_`��	']5<A���y"qNGg6�"a#���y=T$�_=�׽����bܳ!���B���aIں���~�}?Rf?��^�O���l>�7�A͓pb�	�Uw�==���{Mdq��]�r��ǺN��p�8u����sӏt+��9ւu���;���<�
_�j��\ �Zb��	,���r�_}6o��e�*�*
�V�H��E7���H�'�s��ݶv����ݞ�!��"�x��/�s)ڤZg�?6��]uj�w(
<6�F��H��BC���M�y������-���N�@��0*#%��xi������;2*�FL���q/ׇ����a�����7���M�����~��	�J�Cԯ~t&S�W�U���Y+����DM�A��S[W��?�<JI�>�V�]2�He�5S�@B�?y��o��T������;&۴�S�?�ܗA~�����w��/D�K�
�w=F�Цc2Ȥ���e������������