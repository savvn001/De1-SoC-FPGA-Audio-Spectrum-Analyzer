��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl8Z�e���'�����U��PIb�?d����1b7���d���`�����
�@K��̊nA�T�jܕM�B�M��*���3v���$.�{S���^/�����~B4���w[�I|Tk1EC��� �k�j<�	�� <	�ȝ�cp��HP�X[%#0M��`��Ń���RC�s:�)�����x\A�Q1i���9��ym�
_AW6��\I��"Bq������|mH����IJuM~��G�AM��c�}y(��#w�O�S��Ij6A�)4a��Sr�A�)R ����I���6I �����!# ]��wE7���K�?
$�92��9�ů��Eo�ס��S
h�8��S��u��5-����:`�`�&o� O� ���n`�W�?;��"�&�OK~���3�����L�'r,5ؚLx�%X�6�~��.�)�����<p�/�1�-V���b�o�?nwZ��r\I���kZ�V3Ӫ���}���[���򣺦]�S ��8*���nß����� n�DxT�.���|	m���]eO��2w�֒�ԝ�a�P��1F���_~n�i�8�?�^ �>V�$�^�WCoM����jא�P@I�����v��<�R��e0�D���^	��|���\�fu��1��<�W��L�M��k͖ �k\���_�O���WX���â��9Q�գ%lՇ���Pc���9� ]c3�@��\7�ъ�i���H�h���#K�hG�����9s��J�mQ�mĚ>��(�<"��9`,^=�9%�P�Q����R�H�åf���yݻR-����o�	Y���{E��J���w@ ?�">ُ�vDC)�|�"�m4e:ڏ��os��:�#߶#jR|���R�����%�O�ܦ�����v�ݵ��c�������In��EN �9d!"*�Nt U�9������ηJ�r��.���E�韤�	R���AOu:��1N��t��Gfhey�[\,C�����E�#jt}ZYAVх&��$~�F+եe��pKA�����Ҹ�?���ݱ'�`�q�^������M�*f��Ÿ�{8��&��R���)R��m��M�+7h;�J��u Cݟ���
X�DQ��2��.��Ё�-޶�G����q>�?�����)ū&�w��1{�o�� ?d9��+�Z�y�ME���0�v��0f�B��]ʡ�7	�˦�&:V�=��@#!��ݜșoY��[�`�?1P�J�]3��:�~	�(ը�]Mk����P�۞4*�x���T#�gvȉ>e�\J?������H�-a�'7;$�'h���3>N�d*_�'��W?�"�n����K�^���Oe2K{�/�EF��Ƴ��H8� �뵒��0c� �<0oCq�-�c;�d�ӑ�I�X���� ?��l,sFw���+�'7�3`���Fi��Y��+��-VJ��m����/�n%9]߫N���T��s�ܭGo�ԅ���o�^�tye��L,��٪_u�_s�:=8��dH��j�?�7���-���K��8���=�"NV������8>���W��|!ڸ�Uu�M�hO� �_渝��!U�	�9�!W!����_�����"�..�T���n�3ux٭E�>�* ����g�(ǉ��İ��3��A�¦{20�n�xIm�n� I�.�/+-��O��h�AB���q��N.M��=�ti�8����yiw��=bj�9��T�s�m����� �*�>k'�����@�q%�~�ZY�4-�y��3�x�~�`�I�{�9�� (��c`�z��/�����o�^l���,|�"(x��TW�EM�ތ���k�������+�ao�`~ǔ��>�Cی�:��!I�x��˛���� |����p2�h��RH��Qؖ7֯�Zȁm���Ӹ���� $R]��'QmS���Cߒ�v׍&RO&���L 	q������쳌4���OJ�X@~�I�6��O�J�@���f ������A�ĩk�H����te��LZ���\Tj4gmݦ��'|�&l�T�N1�@�]f&a�0��Q=��i�+aY��t��1X�
�� ��z��E鴤��#���-1��yZ{@�@�$����Ba�I��τ+���&��"d���ͷ��_, eE�{�r������������ ��u�PG8 ����#(xǪ�=b��ńǺ�\r\%��K���6���\� 	�{RDϑ�Z��R�:�"9�B��ⅲJ2��[��(�mU�����ΗR&_Z�\��?�Jߴ��2R.����:�����1WL��9�2��g?��X��:��h�D��{UaX�ZƤ�˅4p|��A3�_�JO�I�h,��&��F��{C�V������,K�����8ɢs�ꟻ΀�~�w��SE�5���TN`��z!&귳�ԃ�f���t��N3����y��� ���]��Y��?�1�"P�gm�*5�.����.�"K��Q�@|{�)_���ɦ����*8�]@P����>���*!���ԁ'c֑����I���7���;�y[0�S4nV�Vr"`B�-�Gm7�o��H����M�s�q�ع?{��(޺��{�0��̘;J���b���̾�����"
fm�A��ႅ�lg�<�n;��E�T�yR�f����������қ�f�琔��E��c��h�]�!c>ƿ���7��G�c9%6W7���F`����򠔵/G�&��?v�L�%>�ob�R<F#XJg"e��6��O�p��#Mg�(��·�[�)D�I���ez���+#�?��V�2-�V0!F�����Y�J�V~�0�j�I��lM5��& !�p��>����3�O�-��4?@4y�$��Ɂ�{�t����9OG�� �ǰ�RU�P�'�՗�j�|�A��<~�I�"5A������}f�w��v��iR0Z���Eq�M+���.'���g$D~|/��%G����	0fw{'6 3�YR��>�35D��D�g�%u���8d��3��?����2��B2_�h�.��8)����p�j㜑�1�)���}J3�}��2��m�*%���u_���� >C��>��7���Iʰ�*{ʸ&���f��Ѷ��(mG��]U`��^b�����w.5�Qh�i�\�RLk�l#�n ����������oMl�p���R��r`%�;(|��t=����Q�� �_|��zՑ�r���'iD �#�4��%�"��O���E���`�����^��J��x�&�A�=;�B^=4�z���:t,E��|!&���Q�k������;Z#��ڀ�ᛣ��4���$�D↤�NB!
���[��89dV���l����0�l���Lcf�ތHU����~Ϸϔ��tJ����0*h�ܨ⬭,��m餴YN����WQF�����(������F��0���hoe���L��|]���9ș�e�I�,�S�QgԊ�ϕ�vB}�F��� �i�l�E�v��jw�e{K�Ch��ߛ��D&'f���!v�60��Lb����u���0������_��e�iz�������c���c:u+Ͽ�ڋ��4�Yl%Wе�	_mL�&V>�a]e^Îb��~x]:~���*Ps4��:��m�{j�֎W�t����'UG�bŭ��J�<ma4�l��;V��]�{� �;��]��B)�de.-��?��v^�Sb���纚Sc��q��.���b�+��Z;h��2�6��Ν�\e���[^u�E|�kc�C���؄��9��4� ����d���gj	1��������3|�3��q��׺A��1TpY��6�4r����r�F�E5�N�]C�쒞��z��[t�]}���pPF�(�y<>\���>�|@��y���6��l�o4��w���?żp��	�#R�G��5���Y��+�:� ���M>�w��J}cL�@R�7��p����&|��>}j{�?�Wɗ���=�åMI�-6sC�K#���T%:��pn{"�����P�O��aE����i���F��F���6bR  -<��f���ٿ���v��?��lz�`�~]^���׈�H��y3By�̺����������I�BI~|��a���GW��t�2*c�]��i6*/�?���Ug�K~���'
ۮ�_ڔ6�]���"��g�޴	���(�ԛ����.�!B��.����.~V���ݱ1`~	n|WF"���:Z����J�̻�i�8z�V-=_�k�5YF�6�%y�\g���m)��ʧ�2e`	�v����C&?}�>@�S��ה(�/�W�ƆK��>��^��/+e�!ڸJ� 닍�Ӈ%��n@8HzO�s�����^t�/��X�k�^��B]�9#�xD1s�	zo#I���ȃ$�p�����������T�$t	CC�}���lk�����s��і���C����o�a&a.���w7wE��$�!�_!�\x3JXU�xn�߯&m�%%ȷ�E-K��
"��q�L.�hiE�w]����0���VMr��4p�ڃfR�&�����([��'M�N~Ln6�^j���^�ܿ�rL�k��X�/�1_k�%�!���<n���/�.�&��i�L[�e^̪fZ3��5�'+9 Re:$�B.�H���|l�~��xI��8�c�fl)�c���ў��fxũy��=ݎ�Lf��@� )�q�� JΕ�y�����al�a���N�%�h.LM��P����-0��;mQ�}��0Y�D�q6�|?�r�E��o>�@�Рg���Pv�CR�������$?��i��B��R�=�x+2e_��ڄ�JQ���@�M�4Nҍ��ثm��\�8Qj}s����/��ϸ�F�ŸVf�H�JL��{�9|�!�U�WР޼�e����e��&t�aA����ֺ�.3�Ncf ��g7�pgdg `D,�A
+3�ƙ�~����u�Z\"���V
�Y1����r$p*/J��H����5�b���N�w�*���7�p\��
����;���^X���;���,6SB�]/�䱖��&[x�U�l���`�ĜP/Eu�������pn���R{�-�W,�:ۖ�5�ӧ==�K�(�����w�4:'�p���Z�vJ���*d[(�`��62����J��G��$_w[[�`���2x#<��w�P8将��Oh����Z3��q#d�`_�ў������z:�}Fk��~�� ����4����������u����?]1��e����g���	�I�>e��$��(�.\t E�5K�������r�	J�~�ٵ9�VU�v���n���'��������hov�n)��J�����n�Q�X�Q��3QD;��K���Z���@�G�����R���_��)&9:���Y^���"�P��c����ڜA���	ܯ��n�>� b���Ԍ|��s ��ZZ��>�a�m�v��*�2�&�@aEG��vʸ�ab��*}ͲoL<��q,��H���1�)/4���p!�J�>N�T��\�SBQoxA�E���;��bQ�n4�J^�/;c��y�BS�<�},�s�?W�)��&���ϑ�<e��Ć���D���kO0�$j�c����Zʐ��K7�t&�h��#h0�<�R��,�/���`�ў�tχ\��-Qx��cb"�⺴Dm,��Œ�4BH�����ry��61i�mq��L������bFP8���̖��5����bQ��.�?a������\��P��[)sx�a�Eh��J���t5j�qU	��ɓ��ȟ�� *�-�څ��	?���ΎS8�[=� k6��M��'h�sM�+�YQu��-�6j�h�3o��.�\迪D�_��?|iqf�f �[_g����AUw��4����_w��B%�Ճ� ������¡��m��z�t�Q������e�&ˬ7OpL�ɯ�V�iQ{d��͉@�o掣�Ăq��]p��r���	���