��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	(IU�iֽ!�h�S�1�/O�N��C�߹;�䮙p��c�FE_m����1ӎX�T�L޲	y� 0��/@��S��e��0.����c��J3m��^���V�F3�3X)�%���6>����S��E��u_���CƇKUH�W��2A%�P<���3F�e���	�?����5����$�e�K���<����Y�G��k��(�2'#�B�G	h����Qyq�K����.�BÆ�.1��~�{A�F����d�\��$ɳGl#�f��?
WTM#$���k/I���K���($��q�7�h���ͽq��A�A�y�wM�6~YQx����n�j�%C��̔ŵ�-f3m֞�o�I��dxΰ�f"r���w�b�p�I)md��ق=�`�D�74�
��|�$lo�������^7+w�;�P�)�4ތ��Z�1Cm4v�'���r����&vͅڋΧ����.��R�«j�m�o�0�Ļ����
�q� l��
-�R�6p���jk��|j���]�?-�d�\�d.P��sܯ�^pi~���ه��ޣ�T7Ђj�z��N!����G��0�pL{���p��T��_���G�������g�X���s���(+���rV�Q����ٻ�1\�z)UIkR�������F����ΐ)�ao�
�	>����}z܄W\7�HL}�W4@�q;��m�u✄9Nϙ�"n,Z *��D{}��[8Sej�ˋ6|�;T��-R��"���7�^��٧��"���OkP<�N��Ǉ��T��'"��Ia ��YW���ܷ7�̔'u����	�B$�n$�Y�r�ڬ���d��^�"��{r p"�a�\�Nuٖo�5�/;��z�Bo�䂆!4����(�[w�kI��d@W
�[�b�EFI<���)~�	��	'#�}V�+�g�Y?5?���;F5��"@x�'Tek�� 8��w��v�!,V}�j�x��OWO�n�c����IԬ��3�-���%��U�GO���H��?�a���v����!EZE8A��s�T(`SF�ڵߚ�C�+��cbɥ�Ch���Ӟ@��H#^�H�gp|ȁUj�Q>���`D����j'8�:�N�[F����L���*�����hz��j�S`�N�箮�yq�t1)v��Q�&^=��� ��.�qP��_�ZО9n��w��q��z��
y��"Jq�N���S�H��Z�%��:E��i�a�5��,�v���0~�瑪x�Y�$�����%ȶ�w���O��0)�I��}��Hn8�L���BF�ʁ'8��g_g5.d�+?h��2\���1�2j+ D?:4��F7�]�z�쐥(���xSD��˖a��	�Q��6Z�w��*�F��O~{D�& +���6\t�7y۬�y`�$���کr��.m�1��%}[�yn���@�|��ÈE����7�@�����0�s��pm&��̨�G�*��#ӏ����pm�h�q�+;�68{���k���Yֵho�~�ɉ�5�Wfhb.Ӷ,l@V��j��ib���J�����*� .��Kv��8��>z�$O��Iy�XC[zr�)N_�N�	l���BWrp����+3t�շ��u�l�(ͭav19%���� n^Qo/�XR$��X��G����
���%���җm� #|9��s�ڼ���E �~��9-���^	rV'�=�!�I��>�.���U�ؤ�A�G��6�
�oQ�h{���[R��_�X[��G���&��(bȐW���I�
y �=��V��$7f�À����Ot�<��i�u�����,�	�+�h��,[���Ю�-a�r�Z�z�d���+�=r�ѝ�4�8-�i���|�[���g}-;��{k��4�� ��7�dQZ� zT��������1X��==u��Z���6^�rF��B�`�a��#���P�v����aa�̌|�Q�g_N|�s�Dk �
r��'�cT+]霗�����|�WP�i���`법éA�hz��- �U0ͬ^�9�c�e�H ����UV#�h�/0��ŰA	L��q�9�F(�cSM�����~�'Nv�Xt� �i�4&�$�A����y��X�K��)����C�Y8:>�p �a��<���\���\FWP0����n��%����>RN�lF6���o@���L ��������g�:��+E�ؼc�D�p�FJ�f��*pp�HӒ�������!��̃Ӂ/~�i������=��Bjb:�L�E���c�I����Ay��iu�׮B�h�8~�7J-���:�R��=�#��;�/H�z٠X�r���T$S������u-x�6$4  n�=��I�����@�Vg\��k����f���U�$��
��,�zg"�f��3UO_ǉJ�}oh�'#��}rƲ�/+�S��9�NE�f�UU�%?��t8�����\u�"�?Ǳ�ｌ��ۗ4��2��83;Ǖ�/�~@�O>8+9�ʙҠL>Z��#���U�o֊%pwn\�	�/����AQ��sm�P���'ּ��ވ�o%�#�9��5Y�6r��M�Ò� �s()�^g���t���3G��c��>�O�+O*A�Mw�~�^�
���W̓�8��)6��l��>��eoo���{Sl���J��^�c��0��?�E�
C��1,R<Xϕ�.�A�ƺ o��F�}g��X����(}�1�:�u�ʱ���q�C�	$L�9�A$1�Q�D�͐�@��%��&J��uk � ���o��x\ZN�*%(R���
�tZ�XA���f�5ȬS�2�џ�-���?S�?�P��]�?���a��̭�[�xŢ�mJ�2��OPv�:�ztϪM��G�uP�4�M\�}8N>�7P�;��$1�ୌ߄����N����=�/�ك��>l8E�0q�\��,$1��.��;��~�a΢����72�C���1b��4����I�I$�J�ZT��1���[�m�<��Og�L�{ ���@��{�e1meJ��xgos��yH�+d<7������t��"�˺�j���?��J���Z�!����j�]b�����Rȿ ��c���q?�]	vȳ��"�Ly9^�z,.4�j��<a��Q`�]�76�k��ֲf��ޗ+����4��\^UX�A�� Q�@5��sR����Q+c��F��COjh8��y�[���;��j$���Q�0&��SPrg-,�:	v��s��#�󫂳�� ��ϐ{A9�Dqpq^ؘ^�V��F}�@g�*Z#E;)X��ȨH��L{�p�=���;���i�hl����*�~�������z��G��Cf��]��\���4�KC�$��,��� ��H���AQ��g#(�����X����ꤤxU�\2aJ���1��'�*M�V\��ۄ�u�����#����\��"1+-1X y�+�X������ ������������ Ly�}k\Vq�{�Q_.	�L��ț��@ސw�i���i�C
�wƁ�F����:"�_9O��lb�Uҗ��a޹��|Q��)v/^ess��c?��=�ۆ1���^}Z���s`�5"P��5ڜ�c�v������<�	G|�th'��}M��[����NB�K@)|a��B���{h�؆>I�Uy�~>��6��_��V��� 1�˗�v�yjP+�h����QsM��¬��N��[+3F�
��E���j�S}zr���2��CF��Ag���k���cnoe�=�|t9e��khJ����o����;f��^ ��QG�mH�V��r��P^�@^244�̀�{����F�,U��So������&(*�y�E��鞞�Aa|F`�neQ�����LzK�U`��G�gs�w`]ʮ�"� ��i���-ф湉@.�I���1�&S�)��!�hn�%]�T3�@T�%l��^��*����\h�]�G.���"(8��i�!Ro�pF0�r�c=��	�c��2Ϻ?�����>�4�R"����tq�"�㉢��4��iW�*4g�;Җ�"K�"DEϥg�:Qn��'��-K#ˊ�0�Hr��,�����R߂ab\��X�_Q���=\eRn����%S�7?@0��WDw�{�mb��f &V��Oa�����ZJ�BX$-(�w�;�[T��*L��z9c�:�z<�	9ť/5N���N��W
�~��v-���1܍��%7���,T��)/�s�[���6+�ʻz���q��G��-Щ������Er]Vub*�|�
	��"���	��T
#�}�(��Z�l2�RY���Q~B�$^�s�N-\_eO4��C�|�B�	
��*����{TCT���i�$�I��	���
q����W��jo�<w�	��h�n����h�r~�ޛ����=���x�}�nȡ�|�PIS\z��۠;�p�+_�i��J[E����lB`bBF�Zۭ/�Dh[��Z����P������W�(��Z��4�l�J$�e՘r���]�JO"c�ӂ������m�+�W[���{��VYŭ��	J*��)�7G �ԯ�UL��w֫!�D����Uh]�g�E�#1)
�����z6��e�'��!ݼ���~���qJ; J�iw�����U
�(� %��*��;�x�SO�HP[8o�q��vP�p��GF4oeQٹ纈ġ�#E�~�$c�>:�>%�� l�9�$���~^N�k��{���(��gs#µ>��,\5'h�@�B�˹������vǩ~_�9�=$Ps��jc�w>ĭ��x�a�X�EP����&F��I֏�Ps�b��":o?�h��nT�?>%�}�ہ=�Q8�µ��pB&HZ��´�tO���^Aѐ���;DP� �w�y|��	^�C��n��1�ǨN!�Cn�gsȱbS�1�R�U6/��H.���dV�8�Q�*ĿPj�=�\���EA��DHt|�!e &���Ē�-]A�s�c�ڍ��M�)AB_��g��Ft[�(�娠q��]���=��kc����3��R����LY4�aA��R{�s���sHs�z_���
��q'�^����|r;�n���y����4W����r�#�9WZ�&��dz�f���F�jC�gi��4���s��v"��Q�?�K'C;�R�,��BQ�#"�g����{d�9�Z�HX�3���6at��6ʯ�@���W��Ca۠-��nia���}�z�W!�t��{|飸�܏����wo8�Y~�Hyg���+S�0�Ҿ���mvb�_�����YM�;���yM5�O7D8��$Ӧ���A�m�p�v"Čqz�*�f'I�Fy-���ZX�
[oR�B9��I��IQ�;É�nH����[�3�\"�$g
(�4����pƜ'	�($��� ,H��;|@.a!�2If�g5�ya]^�$�1;W0���9������iK�P:����p��n�f��\�
��e��8�鏳�F�a���ʛ��H���Km-����Hu��4��a��8��"/:�kN��- ��H�ϩ�؄)�߈��k3d�i��n��N���s;K�+<T��E��)���m�,Yg��+��*�#j�Z�H�����:��U���\��L��fû	�pE�5��0�U�e�
�c��z=A�3Mm�����[�?M��g�'V��j%�-0z�S�|P)���YY �n[�I�q�×-w�D(�0w�z��p.2.&�MW��N>�� ���1w�M��� o�G *i�2\Zy.�~?��PF�_7�ɱֳ�YdN��:6�s|"���}����l��f����v�,߲�Z���'_�r�m����W-��5~��1[��n��_]�glJ��>�f�ߜ�@���P��8�-�/@��?��	k� _�� D��n��;����m��<g6�a�.+0����wH�0���	���zz+�2����jh�W'�-��EW�k�����UV���A֙[��b)�����L�[E|Ue��i�vq{#-#;�cI\���[|�����_���I}�qV�W�?o]R�;�I]�S�UJ��V?�Z'�]�k�t��y+�����=�?}OE��vp��JN%�ӵ��:�eٚ���V�.K@�r�q�h��r�a(�d�L	�d�������޶��-�ƟW	���z��p��4�o���4ޙ�*R]w�@x�&�	�wPD�E�X>@����>e�r��Ȫ��,DC��b���1��;t�|�{ܳ�]j8�O�6���ѓ��lx���)%!�;@BD?����F�=t��������ܟ<�/�S'�Y[|[l&�)�7�Yd�C�D�*0iL�j�W�id�e��#n1��f����ꐻ�P84l��[�U�pC�2|�rߛ�x�XR�i0I��l�*Z���R9^��ez\�0�ɵM�!�f���⼎�7��]��d� �>�BT�d�)���;��A����L��ښw�l��>|dm�9f�%c��qc{y,9\��0���=|�6&Z�?���̀�� ���C��8��G�#9=wS(<�����uj5�� �	��2��'tt�l�G��s��3P.ֽ1��]k����A�����E!y�ͧ�8(�_'�W�����o|.���t�i_:�N�����o�G���D?��rIxB߆�;h�!�N{�?�f��m�)�W����N;�6K��R���R����2jE'�Z>��� �Jk�<�܀+�0Vu���߸T$�;�^#��)��.�^��1$Oޟ��S��l.f?
�9[��[�_C���!k����ps��|��+�0E��A� &NC�[{Ņ��-\�/��Lt�����K�����m:н��͒S�2o�����U�޿L�	�t\�W�D�����G�]v��>Ļ{�b���yR��=� !o�)m�9h/�n��	�-�Y���D}b4��mp�(�vgw,פ9�͍2>R���fq��r*Q�< /��շ��R�,��e�3�����U9A�c��.,��G�p2�%���!�_�XD�ԪJhf9�m�U>e|�C!ݲ�2e� fda5��>0~��L՗ 6����K�,Q]W/�8����PC m���k\q��3���)v��<�U5O%΄��k�^d@�Qg�l*�F������$���Nj��,����*#���KN�H<�����1B�_�Z�(������e4��ݱz�q���K����YUHW�N�|�JDT�XO3�SD�oZYl'a�������灣k!����:ʶ�}3ǻ<�+���ݮ? ˢ�lu�'�5��c���i�	��G�?�3/�w�}@[��N/"g�E�9�[Dj;�����Z�,�s�{|Hv�`0?���e�K�B��קL��o���,<X���5鴄�[d��{��E:8B5"^�>�w'�03Bɢ�X�A����WAN��%g��|�#���g;�������6�6.�<�6A��.?�ɬs&����j�o �q�"zdC@qrx�S��d�t3+�"8��#���K
m/?� `��'��Alm������*��G�N�yu$�"hΗ.�<BGӭ�Ӑ��4����{fp>%���w{R��Rl0H��$e�n��O��{��'5���1'��&3��?f�~�[vA�(���;�/���۟Ty0w� �Z����3���t�Θ:"#�r-����멁N-T\�D�EV�m'��j�-����������(����D��r�%������هPu[hw����1����|}τѡC~���C�n����g�nDӄ�B?-E��<dVw� ��y�oĴJ{��g����A8���S1��9bw�m�%���$��R��k�2�@�k����	+��i;�UL�ۻD�K:�	�҉�4��g��4��.�n�E�M��&�`���%:�`r��SJ;���T!��3��F��D �ps���]�%3 �J�פ�/iDf�y��A}�R�c���.Q��_7vm��\�g��á���M8�3�g8M��|�V

���	�7��s|З*�C�ʤ?_iȶ�W�N����i�/�F<�( "%��|���.*nC'� ��΋�3ff�YLn:I�1?u��ɘ�f׸��Ĭr
�Ym�x(Nl쁮 �QF����)-F�ޑ�8��O6��/c67;�{~N��0�i�FG��{nN���b;�S�2�pc�R+��D�gܵc�C���x�N��oy���JfJf��!z�g�L�{oS��0j5|}i����ȁQi�2P�.���.�)l�����s�Q�A'��3��=��PsQ�QH<{a�e2�p4K`K�Y�:At��ֳ֙;��V8t�^�
��|̝L�B�ڛ����yݪ��:ˁ�����B�Z���Pv�
�'{���<|����Ac�P/�F���޽����8��|P�:���s׮��&��Z��n�K_Qs܋��h����Oƕ,�k�]P٘q3y�Z�	��f���ЋٹaEz��2+@��2��6:��J�1�{�|�1P���Q����-[B�*�ȥ����O�)�X)�Sn���1F��q���]��	a�Y^È���N�%lD�o:]�l`��>�x�PAF5��fxy�v�R%@o/�G��X��ʌ�2��p�]T�Br/�"-4���I��ʪR������%h�<�kdG,Y����=�F�@y����Z �i�%�&�ʠ�h*���Kn��Rb�7�`l��&ּ�?˺��|�.��[�w{'�!1����W{D)��"�VW���h�֡c
�U8��۵��2![��9Vzu�O�ry'��]�Ѵ��H�a	���c�I��׭���F�*Z=��L�S�7,�B��N��i M���Ώ0$^V��P��4�F-�V"��X�uo���|pt��I0`I\��v|9Y>����M���P�@�xϬ�%��B��wE��]�h��Z!?sP���=�XU�]��4��S��R4������x%*�Ͷ"��/���ڨ�%
%�mnʣ��y�
�Rݏ&��o"�W���J�gO��m���8'�%(��� (��k��y|E�Ǯ+��M|��
a�܋l������)ַ*�r��mq�r��s7Ԩ��h�x�F�L�c%�FKI\�ፋF��d�Ǖ�4�|��`f�l��6I��N�>�z�:�4�Nlu3�8+��kY^C�ބ7�6����0���*��X���a�5�d�������>3���,�px|eި��8��#�犑`�*Q�{�A������Q=��C	���Q�ſ�f���P��u�PDf5cz��9���L��OD�J~���/��,ր&3�s_�Vi�I[a�B�r��P�tGQ�`�'��>J��J~�ly�5}T}F��ɠ�7Ky�6ڿA�s����ṗm�]�-X����J�#�u0��8��M�97��Ŏe���$<���c�x�3������	�l팪�I�/�\���%�u�!5��7��	�YD�4w����ߎ'�5�b�ZRb�9e�n�&7���n�l��bE�{3<��S: R�K�nC��;1�Bg#�O�C�W�-c�W#����
�W�}�����h�avb�F�|�R+y:���|U��N��{:˃o�����D��1	��=��7v]��g����ȡb}���2����SE���4x�x�/$y���`��DS&!���o��x��!�ݏ
-���F�5v>��g����k�]Z��>�����pD%Q���tpX�<N���ʪ?uҼ�u�#�j׸Z���|YӨI�(F�{@u�b�hr :�1�:�y�����ҧ�XU_�"�������ң�Y�U	K,�}��J,1F��z�Է��s�Xm�XaV��!�g`���`m��]��2��MP�����̓#y�ߌ+U�����mNp�g&5\��arDDc�"�֩t�śҋ��	�m�o�sBX��CK�'wN�����Ŏ\����b��c���[C���M�c��������k�[J�aۑ/ꡅWd
h���(I��G�!u�r�C;�����
Nۥ�Z�b��Ӓ�*�S���V���qr�wn������a�.�շ�ݔL�әd����ǁ:]f�G�圑Qx%�R|)m��e�
6�3���G��7>Èj�h��6꧌ÓJ� �������}��Qx��BM���<��,��d�L58#��J��l��{���eF+S�ҙNeQ�	�}�=ѱX�A6����GD�*Ȋ/�%x0��|6bA.�g��v
o���eF�rB�Q�8Ӻ��b�,!׋�.b�y=Bz�d?;�{)�鷴�1�k����op�v2�OU���=�x>n� �����A������w;M��q��쏖l�}��z�}�&c|�_ہ�S�k'N�3�SUc过����w�&]'oGL���dIA,K�� ��1�҃Ǭ-t�쓉L���D����!5@�R�p��M4)V�i���/\j���;�|�4,D�	�?�����c~�׈��E����Q��/_�.�8���Ǹ>���]L700h{��-=���%�s�k���!N�$���;� e/3��C��ג�)@`���ĊS���Sq�@܍�#�=p�;
���-�p�q����Z��?����	"���aD���� Y��2L�L���A6ʤS;U_����}�Uy͹�x�u?]����Y�@�gh_��L�֠#6�@{U�9�C�i:3��b��MFA���ɑ@�*��LO�0K:GL��*�ء�?�r����z_�#�bv<���J�9G�X�I�{.�ew1��j��|#��$Z�&M ����7�<wd1ō����N��m��b�Ӑ��HG�={������2&�͚����ytƊ�\'F]UGӺ8�7	��\�/���Zw��H�?�,�ғ|���`Ǫv���'S������<��U����44�Ke�VQ�&��l�5mp�\��T��e_���pY@u=<�W{���ƴۦEXdއ�7G��(����1�;�j\ �� �ù,��7����G-��Z��#��*ы%�$�Jh���@*�oنi���$���s���8'7�>���j�����Y�7�=��A�Lg��S��|e�Ux�l�7_��T�p��b�ϔ�j�����k eRCf-��PP�})d~5	=OI�5��w�si����xTф!28��^��ّhJ��з
/*�6Tˁ㚷%��ޣ�`$�Φ|����8���/\�x/_~�^ ao�B@!�@U�*H�ˍ�s��Y�p�bT(`Pe�2����� V������u����,�X䠥��>0|����� I	�c��t�)��쩝lp��vϓ��-�š�鵨6���F��3�ds���
l�hxv��|4n���������=�k��:��2�?k��^�UTy�3�W��q�=J��?7a��5��ZL^3\(��N�e[����r�IccpM:�[)�Y�����n�o��A����P ���<�4ѳGR9�is��_�lJc�P��8�ڍ����:�%�[�Ύ ���+� dY��؞��O�5g♫�ޜ�rƇ�8 �!�����"���������WӠ6U��ly���)����a���vk��C:�������ں��X��.^���^��J�[õG$(Fd�^T��Q�� ?�"w����n�l��u������:��p�ER��7��8��̲��V���_�E}%����t%����H˶H�2�j�5�Mc;�j,Dӥ+��$���<����E�(�2Q���'��rڮi�Y(¸2�3H�k�x��9l�ǡGغ�����k���{��A(�LZ�!������?]��S�g�.��x��y��PA��vH)�ý��u�J��`	��uA��<��=�oTe�82�ID�>X$�����~��د�3dR�����ܲ�5�|۝%�B�p͐qA��nq���нP�Y�-U2����,�1���{�?{nǒ� �ՙ���>&���ֺ�Ӏ�ޗ?�C���T�Jw,�F�D���E�!
�~��B%t���x���a��u�n�q����q�H�y���x6���鱗���N��I��cL���]�ݶ�1���z��ܫ҅���N�6���S�enKlgG�6z� AZ�8��d���b?j���g(�������vž�OľaL�j���nGL�	J�p�D1;I!�Y�\ ffW�P�+��2���C�+I�]�\uBZ`U�X�G��,� >��xEN�Zl (0�%��c%��JB��	҂F����@g���7ƞ�Sq*~]q0�#Y��G�$�a�yƂz#�2��+)}zQ�7�����������Y���.P\h�F]��t��V}�r��sh[I(���j˃Y�~�N�gNѴGԎ�Hs�aл��{�r��w[�WUL�s�R{�����9�Cz���B�q�� �ʼ���	�a�~En����hW��l��1P5B[��|-G�E� AT>�Pv]�q-�[���VDª�m��X� U�O҃����x�w��o>�%��[7�O�e��<9��M$�ۓ��pm!�W�pj�4������K_Cq�X���w;��$�Rdx@J��F-�2]�+~"���=��ؑF�;�'��^'*.��ёgI��ɖ~��j]'��~BFw���= � �f�Ʋs�V�����=�x�kh���p�=�Gcn;h]��kb���$v�W��E�e�_fr��Wc�|e�7���#�,�Ki~0��AH���܆���q�W!�e�t`6����9����N�EWz��W[�?��<s����Ѵ%v�48dGv1�=D�!趄���ޡ0 z�5�˟��pL+*{���̔������T�U~W:�MP�悯ۋY���4QP�.���Ǩ �� �{�6w�'�yK��I��*,�K��<�h �N1F^IS�h�<�w�Ml�"��*��gW J]�i�{թ�5e�Ǣ ԝ�k�iqS�|>c�A�����(�Hܜ���-�G�3�㙽�{������&v��Bq��_k�d�=�N���,]�c�ۗ����;f��f�P
�R ��M�Š���y;Kط<�����>���@�
	͢���n^D1G���A�E�.��]��y��$0|B�`�1ߔ/;]�u�#���_|DR��|�X&��L����T�>��j�%񆌼}��U����C��v��ck��:�'3joEw+.�͵]�/Y�4��v��j`r�F6G�{=���%�XɌ��B$��n3�����P����G.W�{�D����rb ��
��o��a3ҭ{!Pa���>�$���s��E%Bh�ñ먩�c��u8��'�v�g��s�����c��X@>� ��&�DRK.�ШA����N����ē����X�i���g7=��1��uɯ�z�}x�1�F��R�ѯH)©?��`/]Ex�Y��و��4�PP��9��L��[51��Cn�mĚ��K��0irKy�C[U�KZ3�qs��G�!s������i�,��������#B����¼Ư�T�2S�ސx�\�"�vK����mL5R��ƽ	uኰ��z�1C��)ﭰf�p��[�|�/�ƲE�Ψw �՟����9#��`w�G��?Ә��)G7��H�98vd����� -}}��������.�?��E���� 5��C��	s���.�������wy�&!�-a�Zl�2]���۱!sp-E`P��2_����.�]c�z�?]*p{0�HЏ�#*���a"���Yb��4�7Qv|u�����C���y�U���+��2�CcT��sx�+��t�F�D�x�J��iӇ�d���e??7#�5��ՠ|��=��kG$`�ʴ%�U��sHV�;�8�g�m5HM!
F�!�<�eY��%Ԕ1i�c3�t�,��0�uH���\��O��iEp��1 ����$�R�֖T��ӧ��eC�`=L��p�ƒ�L�i�*��0��1ԿXy����>�����E2�����ĕe@&e�W5��@e:ST �u�Ȣ�#��� �n��7���kn�|d�(iB�poۻ�DR9�u�ڨ	�N��8�y	�p�3˓RR���A"c�7��U1yu|�n�����,M�pW���U���{�t��{�Z�����:5���߇�9�X����G3
��O���"��d�hڭ�aR5̌�6����I�9ɈCV�r0|r�.x��]�����E�*��Q]}�
�s�\�J=�w�k�m��E�h����;��|�����]a��zv���1vD"��l<eXw�&����M�6s�<j�"�X����m���FL�6�)g
p��M���J
@�^W�r�w3�sc�zyT�H\L�Ҝ�,�(���%�pR��F�U��"��HO�<���KX,f����=R4n`JA��,�b�6�eB��u�)f�aq��Yw���``��-^���5�+b�D��n�� 
d�1s��6%�	��r�����l�f�n7�WbN}�44_\����c*��k������i���6N�	��0�"٬&�T5^�k+�Yp9`��}l^�H3���Cro��곿��'u�?�i�j@F��[�i�^��{��X�U�$��p�o'0����07����� �2�.��僛Ë��:�`}�%��E�ܯTպNa�7��蔆�|5L�Seyf��#˩�}���"�����K͔�x;l�&8w���7P�l��$Mo�y�9oǣ��bt�?`R�8o ��r�c����y�׾d�`d��3��vV�䃙W�u��y�]c�e�4�P�͙\D��;6,1�I�a��6/*%���m&�����zQ"�r(�g�ULʥ����8��ǭY����V��`TIB�BA�lJΦ��]�)$��=�t�di����@���Tè!΀J�IB! 3�/��/`*�;Ta�F�oy�s1^�&���y�	�/	9�}�X�>S����1?^��~_լ<Q�Ѣ+x�Xþ9��/
_�ۡ��+�6s\�.t��tVa%�|5�� 	O���Ć�4o:j���^&��>�/�ĳ_I4�Y�&�	�u[ؾ���5?���?q�Fa��]ԛ]��F$���/��%X��[� ٲ�/�H�k�~蝼����5�2�[P�WG%\M�W��I��h���ࣘS��}T��������������f
� �c8,���U{�ucT7x�*�iU��IV�[/��hY+���S,�A9��}5��j���#X�-Ì�T�O�RA �����S�Z~;%��od����j֫B��e���#�X���!^f._ܽ�Xp�Ѿ>H���߾���\t�����̭p�;Z(�^07X3���J�$�n�
�\
.��cY�{�sf+��+�UZ��@H���I�郾׸ ����0����:�>oP�lzB�$b�����=,��tg��� �H�oG&#w5}��4�̠�ٮj�`*SGi�tolRM�
W�HN�D@��D��9�W_�>7�(aWO��Ri5�aޑ�.Bۦ�sAs���I�ƥ������Qs�VcJ>e��]ft��%�Ύ�C���5O�<�ԕ���h�)���r��~(?��IX������1�y��Jx�c�m>3'ܴi�2������_�g��Ղ2��,�:&���2 �%}���i�j��=V�ڭ��� �8�>��d�~}{��?[Y@���Wť��J�����x\���	OUP�Z�g����<;c���[�sȍh��g��MhXq߉q2��O���%�.\�F�!��G��z�ܣ�� �go`6B~�W�R�H����G���W�ˡ8�?��������V��J��v�cR`+�&e(u-�n%������SE�fz�z��w�t'�~�A�>��ܸ�cH��@!���!�/46��5��Z��^l��)����(OK}����X�3'�X8? s��N�gk{V���'qPS$d��xH!tN��0%�'K���E+m>%��~��O��tu�;~�J�M��hR�8��	v�a�7xWԎ�\�u>P�2vq~4�I��l�h3eK~Q�yU��m�Xs;y�"z.:����S�L�d�ud=��8��vy���h�����6��&��}�q�ة�EL��Mt���z��r������΅Ziߩ�B?���}\���JbP������C�ølz���7t�2��]�[aI�o�l}���s���Ѓ�k�Na�)�3�#?P��Sg�Y�g�����R��h^�nb������CƆ�vG�;�����4T���X�Y�ˀN R��90��C�X��ͧ�a�m�֐��_r��ͤ�k���?��E������`�F�+_�k��3�G��1�~�M����		E����

G�$��O�Xz�e��Я�s9��w��Ћ�4f3����TJ������b��v�+��*P�3�p|���Z�d�y!O������O���LG���4 �=j��&.��79�;:]U���*�5�
���I�y>=0Z����D3�7��j��X�U/����[(�(G6�pp���w��&�!A�f;�J�� ��J���Ql!F�A�[U���:�+
��'LXe���"�ؔ̏�Bq���=�2�M꥘�y+$���\�{I_�k^8��p�*�xp�}�X� ��vhB�R�'����;JN��*_�7�n�URk*t~�xo$�����m,������CՇs���x�Qf����1��@�Y@Ŵ���J0� ��2"�#ʫBQ��]�r!�1����I�E����P*hs�u�2�����S}�� �{|�؉Ϫ�af�/�����Ҧ�K�*���kQ���뛦�L�ǆ�A7B�����a����!r��gE�	�,3��|'4��ߥw�� ���誉'��8��$h�iGr���( �uK�L����I+')k�wWtbvN�qN� �T�B��M�3�P;8���t߲�~�x���tbT8��O �,D�*���=��W������*/��ȔC���W/�
I���zW'+tc�(�d!�����N{�?[E�Ūda?�h�	À���Ž6]����	��@�fgZ˽�7{�s�����)R��T�T��򴸂a�L�tP�:o>�Z\<�������^ݍ��QW1�|��sj��C5��C(G��HX�
�Sgn�ҟ!,�Bɷ���>��'��TE���@�|H�Q���ضXvNu�]xa��8�2S¤��+�.D1�.���렽�L�hA�>���v�	
���K�eOƋ�0����Y�(i>�Wo�����t�q���謷9�ev��S~�t]G&�\{�v���j
i�u��__�HBȃ�J��p���y!��w�r����@6x�9!)7�"�(E����8�>O������ò�6� rg_��Q%
����"����#��z�_
��r�>b��%xe����1��ψ���7v�|?�?�>]�/��G�^u[��H�,ky�����p����3��Խ�l	פ�]g�l��<W�6���L��|(���)�i7X��`�I\�`�V� ��0#��B�!
�p��ض�oxx9{��������3���֦��}����L�%�XY<�k^m ����
&)U#��p��my��9ϱ
�F�^R'6����َQ�Fz[c�qo�xg��]e��-k��@�r(��j�7��lH]7�����.��of0v�Zn��wl������_y;�ڡ���A|Я��v����&=����<��'��e�؝��̠� ���\{����i�U�	�н���:u��r�u��cò�m1���O��rr�u$靛wZ&6 V��x�����l��2�N36WE�@�2
K�>0qJ��}���1��x�f�wI8,c��AoAұ����Y��b��,��s�s��$ ��C�D���(+�
�n�|�Y��"�^�	8.b���������'5���ոcHE�Y�i{� "n^�g��ΘQe��DUI�Z�Y��������!����7����/O���'��'O/56��\swR&6;���FݢG������(BGL���t*Z \���
��b�ٶ=�&�%�E�G�m�u�C<�y�� cb\�d�k��#���d	��%$c%H����kjVSK���h��[:c��a����9k�r��%K����	j�{��$� @Ӯ��ǚ�Ә}����2�~KP���r���%��Ёr�cg����1�צIضf��~Y��Sɂ��o��̙ʃ"�G����ީ�*Q�b���1���Q�� ��$���>�L�v�S����Un�	�bF�}@{�3�[լ��UA.c�A��dQ�¤w r0]��sD��)���lG����M���R�S84cČm�R�B�e{;��1��Z�-G��@*��KH�{c����>W7J�w�,N��*�}'�B�W$OB�؈���ؖE�,�����BO&�p�yl�Ob<=Z+��Rs͸���gvL��^�TZLXƦ]�"΀�k�'�.8��^c��_��'6xE��l%Q�v[���ON�1�WY>i|��٭�q>��pl� ����}����agw� HpaL�Jd��I���XX��T����?S�敪zfR9
o%r��T�p.�!�̾V-?F�Č��0@qjs�|�z�^��������y2�3��Ō��f\�o����q�}P���r�N`�K�3����Gs�f��:O��7�߽Cq�x�ix��f�S�{������D{{|v�7���Hl�L����K!S����/��SF9�5�M�!��T{5��J�_����Ly�'�䙜\��uԱ��ՀI@�u��!P�*\�kl��xi�xh�C��y��R �L��j=�P,N6�o[`�pdY�����V�=��J���<�eo��U:�0T
���P���'�\S'�/z�ʖ��N�6`�Mf����W�m��T|mA���4Å΃�&�q�<���ٱ��)��=<3E�e�տd�2e����)'��Nk��]���[���&k��*�b�;1�IK�*��A�)��Bs�e�ӱ���������=<�f�`�����,t
���,éɽ|�':�kZ��eD���v����Gݱ�}tS@�:O�m��G��H �-��`e�E2�՟�
�-e��ϑ�Պ�!�$�q0�@u�{m8�hf�q{J�,��+��"d+��uF��Q�/�J)`�����4ER&=k[��B�0)�\�U�T��ش��AZ��Z�aL/�� ���X�ާ|^X��x� �e���d("�cmuJ�d�-�����8�ҷ�Q�w����_/��Qj�=!sUNJl��.����"q$���}�k�)Jt/(���ـbI��X���as�r?�~�T��%G�/�2����N
�{ii��:@���c���A��v�5�b��+CK�[�ԣr@�H7��$�>�W�+�S҇�G&x����ߖ�k_�bzW��ߞ
�%�'�Z�Ã��0F���pB�]��Fէ�a8/�1\���$��42���m�v\��`(�	fV�h�Ԏ�רj �՚�,Du	�7v�2DrB���
�b����L�k3i0޺2*]zx �@ڊ��Ž�t�:�ಁ�i��@�G�k1ŧ���KT�@�狯�>Y���uZNnkH����T#���D���8m	�-Gh!���zdf����Q`�-��+����H;��/ ��b1�9����gH.����y�|�1�zI�O�ʖ�l��t��?�{���-1�}�j����O��b��4?�w �|fY:w3��HT�� r�]Hm��؟}F.R=v���P�k��?����w��Ǒ'�w������5���4D}Tx�]��?ݸ_c��T�v�]�K�e�n6��*p&����a��	�7<rت%����"�r�#gJ0`����*T�Y	��̚ҝ�;1%�޹Yw��:���&*�c�z��GSW�
)c��J`�8�z�*D��Of��^��:�s����� ��kW�q����p����%D��.	LU���V1���?r�e[K�k�g`�sS���+&{�R��r��~;6�r�6@�-���X
��o��pÿ�2O�r,�@yG����
��,�`�OI���t��_�T�=�p�PŚ���m�i������%n�,c�R��P_w�����	*[*V�z~��@T�7g'�!x�r�L���EI�9�;W2�����h�p�@LVi��끱X��9��@��n��[�GK_�I��t'v����|�8>������LӖ��,L���1b���B��jU�zjO=��8�\�*j�K�5�g�)��|!���3IJ�δ�Z��{��,̖��m���\��n	��i�<��k[��%
��PW�y�a�6 �	|�)R"�\w^cS=z�	Q���K�M�(�r�33K�:F~5�!�i�m�E�,�o���?�#�z ���O�p��o��A���B�&퀃�x��K��w�ͺ�Ju�_�s��H�~c9yN�m|Nl;x�;�Iv3���2<�#P_�v�)�>R�B��r��c�#?�ڬ��CcY���Zo�Я�E���!E\�`�:��,�r?4�$�Ǚ;��5ƹ�i���Ɋ�!�����jK��z^׉�U���ز��ܦ�`d��9l��P�X*�R�MB���:!�d�ܰ���H�>EX������<�����i��M������w�a�Q2�;�k�\�J��r[���åYi�SA��G�T���e<��
�M��J�u*p�<��-���/�#%/. �e����%�3��r��H���4i.���U��=3E�5e�g����v:�w@�4E?	b��1+ۋn�������ﺶxGo/i@���R6D*a�!�@ya��W�!G�̑�_4{f��sy˫æy�5ޓF�FOh�%2�5���o���S)S$^U�`;�N	�r�)@��N{tK���%r:�ww+8A#E�S�����P��1�<v�U:��
,mB�eT�m���%;F�s�)���MJَ��\�
�����6�M%"Ġ�T�\׌��BK��y�Ȑ�O���֏WW��H�}x{>��}R:����ul:����:P��x`�Sߊ��m�t=�o��y�LG��F��h�_�n@�3@�R��ܹ��p�ԘK^��#Ȩ$��8�p��bf����FYc #�/��l��<&_��Ut�orO1MO�5���O�򙮷e���P`,!F�0g��q=�&�-�E�a(�.$mx�7>�rp���8pWC��]ɎK�Da]×q������*�iJ����I�%�Z�p��pXwQ�-�̄=�)�������������	�K����Ka���@ӲM�H��!��^^Ns2Q���֙.�����# �ˡ�����@��c�L��F�:1�;�Q:X�AQ4d,�g�^)�����;�:�O��P�.I���p���_=#�f���3ydd�'0'��;�B6��T����F}��1�7��R8��X(mB�)��f�T�~���r��/b��`�&�s��}��D��k�"��^X)3�S���Jen�qK�u$΋D�����	�Kz`��ضu�[kǸ$�0�>D�w��=�{�U�7:Q:P�#٧8K��^|:=J]�.U��>�,Dd(�ةIG{^��C�3P�Dn��Ұ�TL��~�Th�� N2C��d�|��&Ly�z"��S�W��X����"M�m�Ҟ��4��u��<�7c�`�c�mj�u��	��>M�F����+�m����ǋ�븟k�nRB?�[�+U�h�7�u��k3D+�M���$t�AϿ�u��p�@�0&��	�\��m�6lkm�9xv�H�	^����s� �C��b�:��{4/4�#r��,��>�I��/Ɖv�v�V�g���J��np���l��?�s�Ӣ�w6h��7��(O�7���F�a%O�EB�E+~�*Z�E���'��IR�Q٦����4�b#m���4���[4���R���Y킧Y�[�Rzi���_�:�.�7��BbЏR~�%��}#�ד��n��ߩzѺ�� �LR	�?� ���F�N$���� B�S��4�K���(Hup�t����}���~�'� �^�F��V�Va�n�?�c���{���Y̍8�<��յ�l��Z��ę��ւC4 ���d��`Xv���Y<��1d� JO�����'�8�f`�b�]��u�b>_lqc�Δ���{��YT��31WRo�^� 1�#��ڶ�f�}�JC��=��r�[Wв�y�nl�ˎ�{5=6ȵ3���N�ɗ_{�Zt{�r�\�����Xi�����ȿ�)�U�dS#��hKœ ��:�_����k��t�l��2�o����2�́�"��V���1]�8�x���jc�OM�h3�Y��w�8-�9bP@l�p�T/$���~>�4]ջ'�מ ��2���ɽ�}��`��ڸ��}�0g��x�-5	�fC�<�tn���q~�R��5�����1� ��P�iO��zǽ?�tpxyC)���*L�D� �'��\�M٠��g��A�}4���
�yc
	`��v��eK|.�G:;I#"�YPdz��D�µZWF��b�T�9��5o���S{���	�"z�򕥙ʑ�6W������L�G�DF Cm�ה��*��K�hF��C������YS���Wbf��-?��`n�/p���Uka�L�,����?�]��I�ݣ=z��|������ C����<�u����\���Ϥ��m<��C��^���ř�	� _��m܀r�)�� nm.}�	_a�Q�Noe�(Z��@�b�w��vg�5�8�,�g�M�~B��-�.�b�sedT���"H�F7�����~w�K3����퀐ܾ �F&}t��q��4fd0�s���L˹ǊnRW�4G6�wc;���	@�ʢ-:MȤk���MWLdU�6��� Xri��	.�%NOַ��SE6'����v��cӣ�RԼ��UX�޿��m�u�/��w�
���Ϲ/�	�y`Ϫ.����"t���ļ"��i��ac�&���E���g@�M�&��_<�������^�`ӊ�}q࣯�o30CZ��BV���\��cJ�	�!h�qK�5�(�
z���&�tI�)a��B���s�E����w�_|�i!� FN��
�4D�&�q����W-�kR�#S:N辘HM����0�5�5�ۥ#Ɂn}�2`�ߺ<<�z˫Y��ҧi�ܕuy���
�e�j��D#zH�.Mb>��ӭ��bP�M%�_�6�-�cR��>ԛ�d���c�
�w�+�zlZc��1"ve0�`nQ�Pд<��\~&Q��<�T��6�=p�3�Z�U]�����u��F�O#�u���.b|������ױ�^ѩT{u�S!m�N����?�s>��S��g>�Y�/ͩ�8�e�i1:���l-�?�ޮj4��#P�=j�%�50\-���p%�$[�v%-�X��N��E�eJ*?����7��*M���TE���s�:1Z�M�O�XpZ|��l3�Ë�V����:QО�'T|�v�
n��GA�^m��K�И���^�s���z�+��X�g��4�lr
��( �T�*��#���O��,(���]`�6
_��NNR�Ro����(U5�%Lv�j�3��C*=;ۄPap(����~�����rܸ�r�`	�<��I����A�	Զ4뒭� �~L��F�|6Hb�L~���R��	�x�a�����5��IƝi���/Ls��
!���]�|"ROIJ?P�v���τ��1@�:Z�$��3�y#�/l#�6�.�>S�����#'������,�]UtqJ�,_?�7��=���?-D�qRj�uO��Q��/vU������[�\�#�MC�<����I�tU���/,0�	�6��E�b�`nNzaq���fH	�d�臿����s����ё�X���0:���$$-)���ߌW6�.���N�A��c	���*aU�O9Ý7����nGbLb�RX�ĳd<$?U�]�9���u[�~�
s��U�5`�Hcت#�R������%�Hd�c��$>�~י�y��F�>��[��ݻv�{�p_�Ƈ���ɡ+-����G�� ��]^'��B��W�<K���=@�=�!��^��D[A�,��$4��+�V��KFQߣN�тba�17�����O�����S5���+�f�%�����\I9���������7�� !���?�68��Խ���T�M"�Ex�����܍�ɬH��&�����ʒ�4F2�4��1s�Ec�0�J�ֺzL8�}5	��,��7ũ}--8?�$���G�G�~���!񜹼b;�n,��3���'o�!� /�{�� ��7�X9��S5�M�m9Mbۛ	ҳ��L������Z��/��X�L��fR^<�3��+��!�ʯ��^e���NE�>�9�72n�����4��=
�|�-F�A~�M��r��S!X�oTx����j
��/b�C£a��(kYc�$Q]������xD2/
bƪ��v���گ�P/O4��f��x.���YH}��ʀ�ʛ��xKf��$}&���5j���ڧ�+*)��P�dU��.�x�1���Qi� �%�>�B0����+Op��$2�@���&%A5��G�q<�طXV�*��1�q�	t��=%��_1�QB�uJ 5(��b09]�S��2geY?�?=���&X�&���kzT��檴��#;�����d���t"ņh�*>�����G�i.��DF��=P�Qs�#��nw"	A�����°)*+iQ��.@���z�⎣�-r�F��,Llm6��� ��g��^xL�M�j��@�u��xQ@�y�v2���Ԙ��Ɛ�J X����ۓ�;����"���gPe��3�t q�;F;�]@�2�����(3jo���r��Xq\��\��aǰW�@� @�P��O�>�傎���`�
�%���X�+�	����B�x��G���۞�{Ӛ�==��֕m��%�I~-���9������4~��7J�e���k7~;� �ݾb/ShF@��'L�wM��1��&,�V=|}=S�IA�@[N$2*�ɚe�x�Wɰc����0�.�~D�;O�� ��`*�d�o�'�-�jn�/{/.���|��j�4J���>Y��^��	6>a_?�ze�kx�W��V�r����}�w���9�K�R�lYoC}�ef��ί�%y�����HOn1!W�f�tA|�d��^�Ι��eAL�?E� ��7q�!Nկ��*>�c������,�κ�x{�XYs��H�ԙL�h�m������ͅ�R��jh�/�D�� M@��5R�fԤ����h�]�"m�,<�me�f���	w��ɫ�j��rF(q1ߋ����s�u��k-�zbeoV�`���)���*͝��z2¾��~�/�n�ߌx��ڂ6tW4��>�v9�r֊�P=}�i9���_�����U��n�_ �Yu`�i��Ή5z��{U<���F��-1�80xT��֧��\�@�t�μ�!7a�y�&�p�ً�4�D�F�Z��*���g*�z�}/����(�A�1�=F��6��}�V�w�M��}܌�"t<1�(b'p�:e(%�;.�qݾ�!8+~?#ctm
�%>F���|V�
c��^�0�'������������v�"���r��)�Ye>��(�*�G����aw�ao�(�=�T�Ǵ0���v�_&���lv��.�q�'��o��Ag%��� �|N�,�����+<?C5��aȖxD�@K������M�y����F��pػ}"��$���g�·t`�_�~���׆AЃ=f��d"�犼�j�Y��ϫ��D.�8��i^d��r�Vpn,v-���bޟ�6ܣ��5�SE1Vj��9���V��ߘe�}�5z�&����>�����?�9UZ����r��A�|��1+� ��Ͷ�UP�E~�mo'N	��,j������E����T�4���a�W�N9�;�=�����Ӆ"�p�@)%tb�ln15�r^ᘇ�]c_ 
��������.ߤ�Wt��9tc�E��.>)�P:��A2��>2"q��;���%vl	cr]�8w2��pز`K�����݇�#���J�圻���UVr�׍�_@���p���x��L�Q
�7�@J�������"�
�N�E6km}}�ϲ1�Mb1���8W"0o�g`/�/�/fkR^�^��mpK�ϫ4���i�Z��*�1γ2�@��NN�u%.v��q�&�F\�79�B֡�����0�����aY_/L��'gůh�>�U�Է�é*���~��`��F�у�<Z�AiPlA�z"�!��CUZ]w�@���r��{r >���6����Q ����wJ��n���!6�X]��ǒ�9�
��f���̏hO�W�g���[�m�ARDj����LU��yo`�i��t!��AƦ���t5����nsϣC��.��>��ɜ�u�)�N��d ��L�C���sR�巶�3�2 +�Lm���������L���3@i�G��48�v�w���AGoʊٺ��9�� ��{�ɍ���^���a)7�����K�8Ϥ�_����2�
.�3,J�A��Ŕ_���n��Ώ��N��$������{�B,�n��b
88�p^v9S�Ԍ�W��2t��҅���$���MѤ2�0C�R̖k��	ܱ�`��rM�m`�,V��e.�w���K�G#x�)��+U�p`��#�9�O�3�5�N���J^��Y]��rhu'�~��:cM��-T�I(��x�S>�J�����LӜ���_+w��k�!)Mn ���ݖD�x��ˬ��Q*g�����H��B���ֈ�3�׷c�2��N�pnq���x%R)��(�A=���]R��j
n���]1eP�X�(�᳷4�@9��W����O8�+�Τ�����G��C%���]A)+[�@"*�Q�R�v癰{9��o�����{a��b�z���(^��YRR�4��_9m�5b-Ct���AU�[Z���� �t/��%K��v�:߅(k�1;�D#�j�4ozu����iI�͍��r$�A����q��/� �!X���}YES��Y�3uAPOZ-LeV�i}0YR���n�dP�,�����{<�O��m{���D.ND
JBU�AFv�s���mC�N"��C+���ݒ�u����Aŭ{���;���GwQK�K�� i*�����oOq�i��qj�����=c��>�r��6Ȁ����WIv�^�8QK�~jB�sOԒ�˙#{3�M[Y'nf��>23��$/��a�('η��������V�Q��ަ0��ؙ�Lfe2��Vkp�؛�l?(�Z��v�Ĝ���C8(wo��׿Gh��i���."��>� ����]�j3���EC���yux�p#h�hi�h�X҅_py*����6J��ǡ��*�t@I��;8�q����3�5M�2n�� ��xB|=��J�@:�r�RS/�������Vq�[��O��- n��7�%n�p�U�Ȏl@+��I�#��F�|�V����O4�ƨ��~�dt�R�T_}ԤQ��@u��q�mW��I��	=>H'�,��.�F�z_xs��!��0EK�9��4�dH�":�DR��FL��:����6r��ė|w�Y���wb����дe���-��xy�p�a�ʉ���YJ�̜�^�@��^�uou< ��B`)7^��S��e�X�(T!ѻ�;�B��7�R�i�*�v���G'@E�-|���n/O��F��^�SJ>�G�@���	K����-ʺʓL�#��p6���͍n}s��j�Ї��\��#� �@���}�sx��!d��~cNq����G��&v�@\�?��m�W�[�#�E���e�;3;ш���֩�D�5=���!�($k;3Bo��vи-�tIb��˷Z��K�ݣB'�X���K#����\%>3ujq��i�<+�.�^NLZ��n������l�?���r�
к�b�a�����C-��}���i�h�J��+>�;%LHr�	���.!�3]�	�qTu��D0!��K�d� h|��j�6OBu��7Ęv��ttoi(��3n+��h��p�`q+�/כ
A/�.��:��-v���"��p#��B��/��!w���x�؁bx1z}?�b���Zn��d���c�J�h�k'2����wOsZ�>���/�]�=H}0��#������~ɛ�������1�5��u%Aٝ��Z��@��%�
9�~�"��.G;�J��
℻r����r~���>����e�8\v<�F��#���)�0�ޯ8��@���rR�NE�l�i�Ό��#㪽~��NbCk����F{���l�bFKdq��Q�O�:Nw�z��.~�	�@KV5��v~?`)C�ƵdU����tv4�=���%�N?xhE����J��;���S	jd0K���1���Z�㳚.�7����~e��j[eT�0�찓���$t$�:�f�$��厢#�����a��vƖ����ߝ��5�wq��U�jO�n\�@�1��]q7��r�%-���L@���d�к�pβrb�N�ܷ8�Ta5��@��M�C1�h��V��ca�A��h1��Oq`�I�̧2��& ���0x���2��/_��&��^*��4�b��k����"z5�u	zx�Ȗ�#и���6: �����B�*�>���wr��C�Uq��L����i��T����rfXn���a��~�p�3��L�&�E<�5�� ��R�)]�|eU0���3
��KmF}�9��Ov@��u��d��b8o����V	@o3ljl�®�y.Iq�|���5I�K��!B��v�:����`m�p��~��2�:ƉO�s��]�X�]�P`���w�]����S;6q��\�T$�oh_�.��d_�� $�S�&��"R:�7�����	�,�&���zB�M9�����S��M�Nƛ�;;���v�`e��C�6���u�Χ^��K�8���&}��*���$ܾPq}P{�&o�7'>�����XKN�$�"Qn�
�aV��@�4�h/f;��VN���mM?RB^�l��l#�
B��t* 0Z�ȋ*z����N
��c!Ad�=�Φ7r;*�z��i���D��� lP<4�e�����������uuZ[4����k� H���	4d֌�;�ˌ�X씂%j���x�a�MS7���a��K�����ᡚ-@���������t�TK̍��i�9�$�W��v�����@�g�(B5���Ig��d \�N,��_&��U�&�uJ��� U&�=ّޫ�g�&�X+j�c�o�u����PD�ci���;��wE�[�$Bt��D	u�G���f�;/�>4�޷�����f�vO��|��l�o�z��m��Gp�Jm�������F�`�(Edң%'�(�`��� 4�!�U�� Q��m����^�&U��O��B��L�ԲQЙ�3�hZ���.�f�C����/��+P\�����C�s�k�-vŁٿ� ��[B�x-��'5��1J��Ң/fL��'D�(v�)��s\�ڬ��<(�Q\M5r^B�*�%�e�c�ţ��&U�;���ka��g��� E!)!qř�N4K���w3`䧏�� ?�
�kD)����-o�[��W����1�����bC��L�rU*���(\�~��Do�i��M���F�&�����mW��CS��w��ל�n�B��*�MĖ��}��KR�2��R#DywS6�@�����	!+�,�dL�U���WDg-㩚}qܚ��jb琒 �ؓ�J���{R��|�*��(±ʯ3�j7��Pj�yY�d�e�0\�~�֌�ۍHn��q���Nu����=�����}Ƌ�r�²"*�}�<�_ڒ�qP�qr�%J`.u(��<�6�Uv}���QZ�A |�Q��c!
Zx|4m	'NĴ�0��:B.NI+�\�8=��ɽ�A	ـL�Z�M��̥�K)� VfvM�9Rb�Nh.[�v[k����ﰧ����e��`7�QTMl$�#�:�l00�/�j@����P'Iv���f�H/�n�b��"�d\�Ϊ��f�B�$L�h����֊-�cg!�kAY��X���d�l/��
�hB���10���>v@�:X���1����RR�V���d	F��"�G�u�3�e��k��C'#�V�@�,�*��������$F\k���B��K+�DZ��8�ˏ��$R1܎�?-9�t�^��m�C}W���S���xIy.D0\��Q��Nt�Ln���x�h�����\h��c�υ�XBݨ�"V��I~�x����J�������̃����#ly�,2,���c��� ��;��q']�.�i<�A�.]�nh���,����6Ǹ�p��mT��i��]��9����o٨%M��}t�� ���Z�!hV ��_jz8�R��aϷlP@�X�%�_&G��XH7(�Ӷ�,\9(��qrO`
d}�]����55c?Q)4��+u(�o�;-�|!pG,�g^�j��l�\�%������
J���%�q� �l�E�	|����k a���N'�<����^�nβ�`	���[OO�pų �߮}O}��z�� a5�A�%F6e3�=��\��"��.Md5.�Z��q�Iϩ��9���t�%�;����愡Z��+w�a.D���Ue��eA-���thMm�W^��+*���+V#��������T�T^zNN���؎�R'z�+b�xj䖲��4>���.�9"�GX��!�Zo�X&�ey�������о��3��i1hF�޼��m�e	ml�CI�O�X sͽ(K.u�K����}�4?t�����b�=lG�BGs�?,����ߢ/2û���e����IL�ȉ,�+���+�����<FB�,c��8cV2��ͭ����=���*�(v��h[o\��20chsw�  2��B�r8�X�ν���PUvԣ]-���C*x��bfy��͆}S�TS-�⊦���du��{k�$�z�V�v)vhe���bj���c�-:%�*�o-� �x.	v�}�Tؖ�p*�0�\���
�϶}��Y���Y���V�1�����?>;M�pE@��%-���U*�2G�~��s��C�:�3��A�-��j����n%�~���p}�)�$޶�f���\C�@h��5��^�G�����L�+r�Wy.!�h�0�V:��G�A��V5)���r%U25> ��
�����P���ae�j�I�����.����
}�\����!L%��;;�k�G�2<-�K��Zƻ�]f{�������fq�����r�5���/d gNڃ�{k�pBk��"��@����ղ:��<%,9G(u�� ������xk������:����~,�k�W� 1'�ª����������h"Q>�X�`�s�`2���}�	����O���pC�=�J����dmN�Q��&��~�A��uљ#����mo�J�����8�4lH��.���6
�z�aNJ�������&4����g݁K�+�w��hR��S��u�'�Xo�PN&��Ӝr���R��Hd�,_�N�K3%l/Ɲ�^ae;���Mo�Ԋ�穖��,LƘ�~�I�l�a�U!�G*�sjI9�����w��iVNj)�a��GG�����C���=4�В>E4��
䘧����m��ț��82E��f��f�,X@�0���tJ��@��V_�I�KT�r=��3����>V��t�T����I	ۛ��*���V�u#��pKҡa���X��fd5$�Z8v���^Ati����-C��c��.�m�o���vq[Xc|��t`'G�I�R��w����)_4��5�{q�bN���i³���Gf#{ׂq�tGO��*�M�*'ݵ��-����Mr��e�,�h��-�h[��Y;�fr��\�Y=տ�,y�d�A	�)�HoC�ٷ��&bD*q��1	�3��aRQ)�jl=�A��� M8��*�u_�%�*&�͒���y�Bp���$1ez��r}��SE���]���R(v�k���c��Z�#$�'G�Q85]�ہ���"f�73n���=�t�����#�/j�a��r=1-�T�_�ɔC�1R� �;��Ks���7f�1��?i��:��n����͒�����k��jk K����y���7򗩔�o�$���}Iq��%=�ɋw��3nrw��7���Ǻ4�=�n8z����ۥ��ݣFF����T��s�U�P�"=N=��>�ń���2S�
7B����ܱ��^��=X�ӨS�]g�uoQ�O�3���yB5�|�jRS�@�Vټ�����%_�����<)0:��_�f���wW���-'����xt��I�����%94����11�� ��0\9�����2R�1��P�!l\�/�F���5{��Z���Bg���.e���H��/yWNs�5O�"J#�AT�ɓ�|��DR�,Î��������7q#��2C��4\v�L��ce:)�7��7�X�Q�y~�°Les����2�<r�~[��K�n����eR���B)%)uu�pCۺq[I��,|!�y�I�&�b���!����W@sz_�W�PT���KF��}�Ħ&�O���lR�Mhl������{n8�d��E�M��]��Ma�K�J�-Q�����|�3M7	�#L,�y�#5Pds�%��E���+ ��m#��V�bIʾ�{��U _P[��l~r��o�0�6�Q.GkV15�XѨ�C�Yf���/Я���E�=�c�����ז&�<�tX�Kc�}1c�F���F��0�-��#}p'2�c@/we��=h�-Z	5��*�6W
��E�|�Ȣ��?ȋ��+�5����[h�R ����p�R��=U��PO�?���d_�c���6�LO�_��/ݕ��'��T"(���Ŝ�|� ���oq��#|�)��l��lf�`',lxhD�1���_����cK�8��;�d�u-���t�]J&�MuO�q�b�z�*|�o� м��拎'}���y�;��ߑ�6i~�k,g�;,��2W��Ң�KjO�!!.W���A�MFɼ�Ҏ�=|�{`��{��,1���n�t	���J��D���x�����?i��d0�P&p���G��UC�&� �'�&27�W��,�+(�M���F�y�I�jsjLMP��c��j	���i�.Jh�F67��R�KS�4>to�U�t�ml��9@Ճ/Gf%+]\� iS$�tQ�fl�[<{h`����q�g�����)4�h��!]�E�QZ�q@�/���B�
���"��E��>{**���K'���á��A��˞�6r*b^��@� ^0�RPm簈�Dg���Bk	P��&���/�|�G��f�"��ʽ�o��5�k//X�WO�Νsڄ<g�P��y���G�`U/iJڿ��S�������,Dm�� w�߸��Ě$!6��:V�}
��ģ3�-I�NJ�����G�2��ǭ�7�fi�!ic�ߪW<�k6[p�>��r�-�o��ް ���xA��1.D����2-�j��@d}��!�Kï[�j9�����=�*r�a�\f�����TcM��3�Q���](%sE�ᠺ���~R6S�e�[f7�W�4m+�����һ�;��9:jk�oN��Io%��0�W3��u��L٠����U�����
q��MSX������1b�:蕒�����w"�� ��HJSV�&�&���mI�4V~~k����6��P=��oEI�0���P�?;�*/�+ˢc�hTb�OR��YF[��+�AJ$]����7�����N5�i�K�� ��*�Y
tzX����_ăU#g���d	�f�8	K$���[r�H�lKjͫ�GJ�&�1���k A���R3S�}e|,���r���ͼ�4�������مLw�#�fP?1�.�e
�O��[�(���hm.Nw���~��(�Co��^2�F��!�4XD.y�r�:�Vٵ|^"7D�E�����4��h�HI@�c�ܰ��IL�O3����9ŧ�S�C�e<"����Oa��P���2�6�Ɓa�$c�lo�D^�,3��v���c����\6i�H��
�4��a*@{"�=��g�h]K���H�t�^�<i��.��M�3`$��i6��?�ʎ,qz~F8��xx����e|���3�ִ��B*��Y*t]���D{a�NR3������;ˋ��1�
���)&�"l����E�l�Y�i��%�ۂ��*%���+����̔iM���e�w���f8�_([wf��U�������$� 52f�:����%����c8�=�Dz@X^�(���ϢD��M�~�vx��*�h:����\��a
�&�3�UbL])�8�{]��3�-ca����΋�.��k�S��P�92�-7�	�j��7�^?+z�vܵh�(���W���&��.�bf��)d����~�� ��ݨ�Z&�tMe^v�T�wo�������'*��.]1�9�^ 9
�G�Oµ�c}��靏������L���@ 07B
\���H��4��U�*,Ko���o��PE�O�ج���m-)و��w:���8:�Gn����ǹw��=�cxJ��3,E���>{a{"�������X�Γ��)��F���'������[�qsF!&M0��\l�w�g=���Tc'Y,5�h����!#ǒPݣ�X���ҋ#r�alTx�t�ѵ}pz)��/�B��!M@s2U������8e��i �oi�t��n��OG� ���^��<� ۶�?Gz`7����v���
�D�Yߏ�裦;�a|i��w���-�n-�zаYޔ��d�ܤ�#�ޖ9�,-��IOe�����݂g�����JNG*�f����ˈS����_�ؘ2�"��ipk3�Bԕ�1�5F��R-כ𙱕A&& g�MNs��i�WbGS��!gFW�xEO&��eӴ�t
C�i����8��-��C���G��X��Gn�۠+r(�U�fö����#���WjU�	�8�oQ[�W-�Ee�8O1��>�r?����<�q�3�(�@�aF�4ˏ����^IkL��"(�����^��t�y��cg@�Q�5�i�2+}T���'��7��7�M'r?ۋe����1�7k.�u@�x��啳NI4��6g��Dt��Ll�4�����E�?��7���`.��pB��]�g�ٵq�ſ&���_3e;�bV�zrvY�t���_�ل�d�M�n��g�gA.�iP������]��b_�H�7�i�a����qM�Ip4kA����뜛Ș��p?I���RS�;���<R�7�$�-,�dW���N+Wk�C�'�S��� ү.�>6ihD��x�zyf��������������6�d,��� T���7��|^�}ݿM�^n0���)���r�&���+8;m�i]wU_RP�)���Lraxi�0�Ob��zԨ7�<��h���:;,�(j�ߘ�_r6Q�!�/	�$��5e������ȱ�M�b��0�/��Y���'�3��z|)Z�/��/���s�����L���6]�Y�LCD#",�z.r�2�b�|��_Ei�
������@�&</�>�p�G��Lص���eme�����1!+E}H�\�HgR&�`�h�Z ��o\����7h����|L�L����6"�H��nQn���p>�D����B���#8��KW�%6����/��h��6�oh�(8���MR���G7H��m0{̿MVA7CH�_L�����c:"��B�G*��@�3�dyvoV��m��	�����`1B&+�:Y'����4�/2 X|���!|z�
xX�@����ɖE�m�zϩ������1+9x����i��Ew�݃˼I<D+~~�+>7�FRL�5@�$�󁐃�,ѠΩ��L�IkCNm� ��
ũ�6n3S�.z��YGdNg�	x�O�-�j��U�m�y�� g֚�����0�@7H|��àY�6Z�@:�U��f�a�8��~1=��%��g+ܳ=���R(���Βp�����/��k�6=�*��&�w�9Z�=w��2e�j/,U ��!��y�xE;�K���|���4�����;��<%�R3�ԈK�����^�[P�BeA$��T@V�V"�ڣ�4c�+D�
3�
3譳̈e��}*Պ53����r�QX�STq��Q����0A27���L_���"|����e�������g�]�wƾ7eu�Y�s������(Qk��n��[�=|ER� �$@��]�ˋI�=��'j&ְ���4"�j�,��)�G�gfE���9�T��Bp�@���>�|K�s�Z�'���y�I�rN(���@C�&��:�q&0��R{�5��������ㄲ#C���1����	�hE�o�1<X7�KO�lԻ�]P1�s�Bd�=h��{�)W@8 ���8��V���,\ݢ�� >��t���Z\�O��u��E�K���]�n��NI��2���R�쪂�c#Qh��$֠鐲�ΩZ�u�����{�ᛦ�>c���u�_s�j�'�Ɏg|L1Z��,�K��Lr)�TΞ���"���g�ĸ�Z�i��߿�c�بU8��^�UYR��A;�s��L��)y�� ��t��	�b�_� U���C�.�R�\L�9�M�s���1�%�O�c�w�t,u���辶uV�<S�;�'�x^#���W�bGb?�
���od�_R!
[�R�"���쑶���wB�!h엨D��>7k�g	M��~~t����w=�I's��z�릘o�)��#��=�߹CrvU���gz�J&�um�iz�����C����ך1Uh�u~�OFq>(~�o'xkY4�=A��|hw���y�/H��hy~�@�h�dw-�2h,J�m~�t?�$�Z ��������Ln�c�%���<�$�S��_�S)���B���M^����9k��F�d���@y/�5�Q��8�#�p�ih��(yUk���[��W-���&_�����(*�b�c��hhL��
�j~�[��'�W.+�0R�E�4�������j �'azz/�՜��v�t���R�Ǟ��I�;G�w߷��1�� _�A3
�,�#� 5Zj�U�OL�h���N3��` y����[��W��gsBQ����}�+zռ��v���(�복�ʡ���q]�P�u1*��Ϛժu�e���j7�����器���.9�+=H��~Its��K(|�(E�2�j�J�w����Dy%$�/���l(���R���L�������w��Ƣ��nh<p�+��<#
C��gH�=��Ū�`������,wG	����BAh���0w�^�1W)�W�B�;��,<�id�bF��a��y,���x,����/�Rs�E�ehJC�Pk��S��T���nc���窴�X�E󞩛����a�~�.����>�7�q�v7������	)��˱DیHȃ>}��wrr�������1��� 濤>�U�����Z8�A����|���\k�k��%0@qJ����.��UZ��ɕ��*B6a�|PL;}�ȱS��+�� ���/���R��G��E����=���`\ۖ���:/�H��ZpA��7�*&M�.��o���u�Gw����M�6�������@��d<�)�p����s$(.��H[�Q"�A�myEe���S�=�T����:�D��e9�a��V䧝��{Nz�������GHil�*/��H�!&��I:�ʐ��i��?�� Dhto�-��yR��!Ҧy@F��3{�͚����Y���'B )�T�3LP\��d�����?�����2$)��ooy� �tw�t�Ŏ�zU7���M�3�P0�UE��V�A�����b���F��[�C>��7ـ?��M�WA�����'&���;74?���9�- ���ޕ���;=6�aO�P��l���w�S��x�b�:
[&ո�,'�.*f}֥�`X8o����j�'� �ü#��&M<�4��2=�-u��4� �U$,w�X͉DD;>;pR���̶���^O$'4eUӹ�zSM�ӵ� �:)}��;�YG�{9�V��'����۔�ƻf-��������&�E�auHE<Pk?ǔE��ɬf�u���l�"iT�1w(�]rB����fw_��N��ݒx�u�r�Y�奨Yr��?�5�Ʋ���*��%�A�0�����'�)v�r�.h�K���%`;�s�i�ς�F�]������[!�l�,rV	;k2����-�@a(j���`Y�13�[�
����v*Fa������\ng�{�E��V��Ĭn��t��5��L����9��~�[Mv�&�[U�ɍ�����/��	��<>�	X�5Hg��W&�v��Y��>�v�aSg�{��f0��#��	�=�X�c���0}��x0_ O�jUg�a}v�Pi�ҿ��C2L���E�2;��P���Ej�������O�εe��Aa9\K��_��6��q���q�S
>�_s����x�heֻ)���Mq!���T���r��w^�{�ZBUTm[��(o���i�|*Qo�bμ�@�v�k�52{�AKn���X�p �qK�0Y���\����n"=�yd�I���R������h�9�t�C��)p$�$��ɒ��/cY_~:F���V��C�e���fW"w�7S1�X'����3��%4���#d�5Sk�[�d�9(��t�;�Y�@S���D%��,$��Y_o�u��g ��v@��~�d��\�c�%5�3]�4D=���p�ұ�,���1Q�n)3�J�!ՋP�I�3�&#���x��HC����j�:��,�R�
�Ÿ@x�nwi��<;�)�w*F���轀 �'*)�tf�ߑ�N�T#�t �����|��n;?Y�����UiN��CZn�;���]���߇bܠ�--���N竭���X���Bk��Ǫa����q��«����r6,�~�1��R��|m~$��rA��R�삌W�i������jQ�X,q��Ԉ?x&g��.#����O�ˁu\��������ȗ)?!UK�@g�$�ݰ������,Dp�0���w�"�G��$O:��d@�q��hx�UPƥ�3��<�9�.�����%��L�Y��� ��)A����/n%OĞ@68�Ѩ�����\�7���t1�z3"�|���m�p5��I;��Еа��/��9���K@$��a���l5d�����=˷�t���2g���(II�7]��d-	��|Ha
�~-�:���Dzq�0�ُ������<ĺ޺�R�&A�J�ќ������q7W��E��.�s$HA
���2���+еvd�x,��M��J�h� ʁ�l�!\�/��+�%�<��D��cM�n�v��������u��г)2`b�O����爆F/��v�nZ`f�2:gU�Wm}O�����j:����]�싺�K��2�JaiW�h�8UY|:���<㞕+\E<{�Rb�!0]*���mŅ.5Ŵ��ƐTK���?�{�5M'S¥�U��;^	��t��$xM*7��s��zc'��>v�a�>�KY �V�I������l��4�S��,���ayH\����#��i�%(_��z�,x	"�[S�rRo�AO���[�f +��ߑ��M	�إ+Z�;`���Υ[��J����&Ɏ�����c����n�a =�'�\dm(-uQ�cp0�-��]��'���ț�����o)�c%D)�"}��3��
B̚UL�ьŠ�[�p���!��Z��ߘ�GLSr��2��a����	H�&��g5�gjBS]���l�um����L����f���q�O���0bR�m��� l���F����m�(_����7iܑ���>()�ݦ�ؒ����v��L��-�P�ͯ�T��_��mc�X�j��t��������sA��S*>�f�@�[�إX֣e]�g��?*�hZ/TᧇE�F�S)1�+�:" �9�5����j�	m��S`�K��B�'���Ӈ�tU�rM����+(w��x2��ZP�b[�� ךE^_�J��N7�6R�$S�����E.d��$��u�g�N�S��󱢜��kؾ!�Fgiꜛt(n�ۨ�6�\'�Nq�-�e�[�n�[��BvxW��4��wM�7h����w�����G��,�0��;"@���X;�x?sƧ���+E=��)��]!����$�Q��0�����k9ѠK�i_��[������8bp0Y�G��tԧ"u��G�!�VU�����A��V��2w��U���`��7�oY��D(�ZR$SO�rq��
�h����2���O�
W�aN���4;o2~�X��I�AVOCY��Xz�S�"v��/��JB(s�f0[T��l�~�9����(LB��_Ej���Q���P�"##�W��{���O�����̤���J����eL�rc)/�� 3UHh��FkZNtl�#mĘ�.����(?��/��Ŏ�?�����!p��r#o�Aꚥ��V��U��E�Tx�,��Aӂf�0
{ZB2L�ω�	�5Uw<z+գC��a����25*��J�+�A������h�s�[�]����0���IU"1���6��E����υ�NX�����|���(?2_y+��:��� ����(�ީ�����%6��}rte$�"�Ҿ7�N�x��;LwN�0D���u�O��qL�{f<���e�O|j^}�����yx��pG�:8�6���GY���A���\_���"�G^���i,m�o��r�X���<0�Q1k�����
\�W�Ҳ�Pn�*u$
|�G<���>0��ǯ��jx�I&^�����rJ g�L��Zƥ�9�z��7(
���!�+4�0��T:ƔW[��M݊v�7%{�u���td˦�3�%k���U��	䄰׍y��v�qh�+T�YJ� B�9���,<l���j�G���@�y� �	Ȓ��-,ɡ_�a@�\����B�a�
#���Ƌ��b�������g��SB헑���[�"p�K���r�E��n�'�ÞC1���&>�G{�l~��(H}�.̻�g*����ֳJK�(�����(u��Z5���P�q���~�����q�����YSդ�s�,D�a�h�ů�}K��ht�� Չ��).�&���Q<)W�Ф�SJ�k��v6v����Os�]��������֪g:f(��&G"'�D�d�Av�����!�?`B���<?�5ǋ����
���.� EtT�BɪS�.�!���P�(L��H�kX?ðNg�OR��{$�͛�+�>�/"B˰V��k��U�Y|q�t&�5*<-b1MVr{5��ee�=���$N�h�4�]�3�X�Q��"w�Jbq��<�6��5<�#F+�l!:X����\�E��c���{{�Lrxv�����!T-��i�E�'�'��D~ k��r�%c=S@��g���Ip�F�9�P�h�d/����aߚ����x��M kSp�ß��|��4���<\�����})�E���a+����t[���!��#��6�(9���3z�@ײ��EF����)d%#�7h�]{�A�����c �/e_��-H� ���X]�Y���l�m��|[�3��'�v�ۥ���Y�� )v�F���S�Z�;Y6�¡t��݃�H�._��yc�.�A?���^&#��ҏ��s��j�F��3r"'f��ZcVq�L�/�+Z��{������b&��~u�O���d���Ž���\�;�M��Er����Ҳ���G$~QŪ4�}�]�S4�	��83��WQ�N�[����V��{3�``B�a���L�O��R�Y��zC������`B���g��%�V:-:b͒���rM9�e]��g�9��"���R\���tC�����"�33�P��fY�|�<�C�9�C��
�1�VP!I���~�ߐ~�H+�X��fM��9T(�F4�g$g���uڬ��T2�5�6���r�{��o\s��0�tV����b�)r����Ga�Ex�}�ü�S�'�WE�����I��*�/}��l�l[����G4	� 2�J1�PͲ����E½e���\��L?�O~u���9������=��h
}�E�J!�s�Ȁ����T<y!L6�Up��l:^�ɠ3�$ĝ��]K��,��hX�[�}��fcXa���9��m��a�3q�f�t�������;�;ƐylA�vb���>�N�CuI�B���|G)i�,�;�f+��p�� ���6�4��k�Ş�{�S�v:6���N�d���Z4i!*e$�G6�n�'ӣ��O|+�O����?����D\�J'�a%|�5��WchA	�!.�N*�G��8�,Iϻ|oEՂ/ۀp3�|�����ud���G�ߍ!>��H֦S��]���N����$Ve��|��⾇[�{��|�4��"���֨�Â �)��"Him��^̗��'�Θͼ=����	W��̺�i��_�r�[2P3.�Q/4$&d>�����}�8��S,�Thxl~��UO�/)S�����7Q[�����פb���#ߖ�����3*ヱ���y��B[��k#t�r�*~T˓�� �����έ��ۙ-@U���ع�+�!F��]z��$��je����n��_��T����-�A�V4ӊ��VeZ3��ka��wy���|J�5��U]�sV0���CH��K��#��a�qT�Cm�)��}�C�����T�� ��C��e��6MI�^rr� ��&�����_G�����f���,�E${�������zC�P̏4J��G6��-־<�ƓG�/��틍{��E���n�P���u��ta"Z�<�G���%�7!�y�2�
qd�����t��+��6��7����E��Qb�cn��y[zb~�r�JSv?���bNb�2��g�m�����F��h&T[��u3���>}�=�%�k&��t�ʸO���.�$����$kn#ѓ�ޣ�D�k~����$y'=i����������`�b�&�U{��2`,�,�@vE�O+:zN��fȩ�g�-�.��i�M�O�;�
=�5F 1����-R}�
$Y�!t;��QE�&�%R�-S��ԫ	̎~׺�3J�F���30�?��	��˅���:ʃy8��{M;��J�������{�������҄E�c;���GS��G[D#j��pQ��pnD��|*�6<�_X��Z�T�p���銝=;EɤJ,�_��!#�05�{M���`b�C��������1,��^�ƟY$R���U���Al�9�/�H9�Vpi4�X<�z���-��9�0MX��qV�͛Nؙ���� 2˧�]�o}�
֓mYB��XKE��5��~2�m�M�Te��f`��T��$��ؾ���y;R��V'y#�iw�uR�_߇���i�wU%R�G�}n�`��q��Yp�*_ٛ���@��Œ|�4�^�i˳1?O���r�~ǒ� 5�����j��.�V�ZÝ@�Bܻ�l����צ����J��F��Un��a�!ҭt� g��mU@[l|g�J2f*,�C��u9D��R ���������;id�$c�Q�	�FC~�0ʞ�J~�Q�P}]b�5rGH��<.��.��s�	S�&���� ̨����QS�<��䔎����C�w�_G���îױ�hh�w{��~�̩���(�Rq�z�]<���Ȉ@ų�X�?��I��k��<�����Ui����[+���XC�A� �iݫل6[@b/�[і�3m���v�	�h�'Z�T�T�)���:�)�ʢ	���f2P|.�l�ع���H;�����%r�����q�}pJ�
�����Z|(T�S��E/ �e��tb�>ܠ���������+�1�:�	:|���z��$o�Ϝ6�V�+�bæ���ȼ�l&SG`L?��-����˝I�z�I��Z�: ��v��o�uV�̉^���o�C2�r�N@�V��tK�J��uϙ���Cz,�>.��禊��v�`Ns:�?��Ji����U��4q��S��.����t�Ur��7�7RfG�雷M�$+~|��5�_*��Gw����X�x��,\n{WD���$�v�W�zeeg��$&�ۦt�M�����-Ј���ٚ��io�����M'~��P�ܓ�e{�hI3�%Y���D�e��g�@��x)��	��4 7z�|Tm��.(�|Dx�QP�,���y�[�oL�$����X�O�~L�vsK
/Uqd$���<$�	�L�@�j�6L��X)= �o�iT8����l16��_��R�+����va
ȓ�&��rwyб�����q�����K��j����F^��V����D��l�&��,�u-d���]�ۂ'�J܎�"N�@ �F��Q�:cX�����壙-�4dh2i)2wp��J>��J�������B�l��ہ�U���0�sk��̗� ��rogIs�?�!"�n�"w�߂��d�x��D��_��#���8��L�P#����4.
xG,�D��X�P�k
�L+Ɏ�����$7�N���Lv�ڟ�ۊ7}x�����R̥��^�tB��U�@��\�E����������E{E����W~ɇ~;�-���R���o㪿y�<� qCQ���x`֕D8zT�^�EE��j���>�Z�o7p��T&��)��)	;�\��X�ũs]p�e.�isҏ��ɧ �Iw�=��ϋ��Z�d��k�>��\7~��k�[�	���W��@�-���A�Bv��MRj�Χ��u�4���ъ��(N['tH=�l��"yLJ=]1�����kP��?�@����iG�����H�ۨ���u{<s؇P&����?v�9?�%�w��+�,̮4��x��&�<�ӎ��_4����W͈�HZ��(�v�)b] �����~�%]��]�q@_V+�p!��.��Y.�=��w�<u+�S>��q����*Ә�K��(�ah���磶0���ᙪ�v���Q(%�t6bA-�KS�F�t7S�[qE��D���?M}�ߵ�C�ŕ%����Xo�_�6�C��z5
_�D7�'U����Zo�u[(���z8�s��1���Jc�VK�{ n����E-�hz
Ƒְ��Lx�C��>�H�pL��K��\��z4c�c%^Wv}�⟳������}|9���Ł��8�(	�4��L%��8Q� 鸲�6�����!���l:eV�ߊ4�38MgKTj���ލ�hg��+�+8���8�M*o�Z��� �ك.̲ K��|	��J�Z�0�5��F6�N"א.`��~_|��.Y�n?n��F�#	z������OIR������ȃ�o4����ގ�kL9�����:kДxtL�;��S��  #��[{R�O T���i���ZB���&��K>����P�^�x�d����l"����6�1��E�'��-�ʄ%�C ~�6��w�v�lV~��V�a@���
'I���	Z��.��Ԏ�����w]9Ahp�s2ѱad�~{~;�M-CD���i�v�@�4�����P�����7g��?��`�vD�����}\�B>�;�i��٤e�u��aX�+��G�!��� ����0�_�!�[�b#1�����t��u�@�E��O�񒚥�.l�hZ���U+�5n	�`�=�`r(�Z�#�gfԐ!��e}_c-�Q���Y+f k����7�}N��.���d��D�Z�;◹��7n�� U�� ����=��e?�Bl�^�ːI��j�k�FԸi���2��xCl�G���~��F������̐u T]��˯Ld�5���:d��F�f>�~i���:�5=G̡:�^a䔂O�S��@�s6m^�4��YK�����M�*����NB~w�ʵ�3�]�΅�6��/|j]���I?s�2����wM�5�YȎU6�/�8GT���2�_����Q�V��(?�+i�s�i�ÇI�Vz���6���Q�I���#�C/��f�|�)^4C]$�֐+�i�WxH5���C�@�Y��4��x���v��j�	�^�AK�*M$��f�v�Ê��SQ���6�Y�r�qA�9-]c-y#���	�p��&2Zf�ƛ�1�����m��d3+t�����B�*/��,f�rr��$r��q�@e�E_���.\<�_�V�>dUU�����s~z��x�:��r��oR�|�����KR�[���Y�R��}o��S���s��z��|�^�(�Қ��3 �'ҋf��H5��L@*!I��W<o�NV�0ߌ��o��ι���4��6[�%�cIQ]����p��X�6��X���1�ߦ<����6��0��G�9F���w��2o��r^t�p�XU��v��Ic\�Kt����L�`�XERְ D����X9؛4!X1x��l�/&zґ]�ո�ܵ�W{D+� x��*�����vCUP@2l~
���86�%c��\��Ζ�t��{M�:��}:1�Ӕ��$$���<�YFf�Q����s$���ՍDK%��,��&Ԇ�G����d�Ǘ�)�6�
��o��;�6q�l���z ���9�ʺJJ�^�k���j]�t� M=��Ճ�5���r� _�2��^DŎ��f]���3ؔOݧ��=:����'($�u5��Q"x8�a���%���'�G4H����V�e*�D`�v�E̔K��c�U����%BMOEJ��%�Өޤ"�����$+�Z�R�e ����J5\S��G3�p�đ�z&��(���ň�Xd��h�n�E[��j�R&p@$�OB	>>�]nF&r6��Ks7~Z����3����٩�V��d�$�щ ^������Z�v�u�2��,�M��&O�C$���IZ���wބ�ր>1���݀��?,��Ax��&>��H�K�Z��-�f�m�dxf�� g�d/L�aF��x���gyv-�J3��$�'��u)�x�>ĩ�#����Bʢ���d���f�����d�y���=����B��]�m�����f�Ԗ�u�����S��)|67y�m����	ha@瑘�k0�(�e�2�L�i��<���zW�u�g��B��H�c*b]W�,Q��5=�m�{�_)s�x,&s��Z��Y-�irgG	ؤ����Y�"G�_�ʂ�p����R��h	)��,Z�E5S\3<���U��.����%���m��H��SJb�+��Y�瑿��K��t�<+<�S	���^'[j����̑��	����́�M+�j��L�J`%+�qN���ߖSx�G"������iI+<����'i��r���F�� �������,�l�ri5�*�o����b��R���C�ڪr|�Fk2����)�Z��lRB/Ψ�ޔ�Ƈ��?Ï���b,��JS�~��BQ0�b�J���)��71�#у��ipR\���-��r̓���T2Hε$�S�K��Ϗ�(0�6��}�U�b[����ca����$9٭1��Y��^@O	T/,H���J�@	� Q^�>,�ӆ����6�
=[�4w��#3,7d�Y��[mQ���8�K������"��"j5ءK�ߒ48m��P�w�b(���-�X`�����(?ee��2k�TQ�4'�է��N��v��"�wQ�w@㚼M���Gg�{�n6���A8D���^Ɯ�΅���[�"�<�Ⱥh�|
H� nd��������5�!�#���p8�|�(EAQD#�`��*�5¤�����!H}�&���agh�m�������s��|��ar/����Y�aSE����^� ek����_W
�Yg	6G��L��H�"\׍�d}FvX��/y2#�giˢ�ٷ�&+(��_AT�q��r�����Z`#S,����0��m�FJs�t}=膈����C�o5����^K�}����	g���Cx��!U��XIV@���R��Q�,����,�M �[v�"��O�S��E�WT ��w�>G�/hŅ5���$��8Yj���޲-�;DPob՟ZY
1&��v-_ Y��g�7��.�t=Ѝ��a��ç�(9�6���Y�~ {�D�tw5f�@0�|a־����F�gX߼��L��T+<\*S���|��-	K���,6׫����2��]nJS��d��y����X�'����{�^\̨�o��^:�U7�!��{�����{n#Q�S8�Tz�
�����!sVCð���`�����}��T9U�y�s��7ͼ=y�9k���f�~>C��BEK~č��F��f��@��+nz��)�����Di!l��>���x,3M��w��Z��`�*���;�@�R�@���"��".Ǚ��|F�dH����)	�@��N��f\�m{����J��.ߊ�5���%��[��������ţ��1O�R������{�P�-b��xߜ޴���`AIU��io�ޮ���q��"�-Ԑa+kG��T�������L�Y��t0�d�4P�r���"[���y���\R�I[���t�	߽�M���*�Rcz�i �U�BH�H?��ϭ�b�G�D�p��\�+�`����d}7��@hF�S�����Yo�0��k&h��4�Pf=�5+}s"ķ^��%$�yib�W�M�ЂC���a���a�MW&����+*q(�,7�S�w�/���6K��S�j)b9�l,�MZ��,Ƿ��/��Ԏ�_T���kjy�C4� �b��y:&?���d�\�<�����FbG֨���A�<23���k�.�/I'F�'���Ҍ;�-���!&�gP����)�#��ɡ��x�M{t�ä<�L
��a��FJ�W��ɜ��Q�%�O<;KS��˼c�W�[�,(j��/BȤ��������0��YD(w���*��´�A??pB^�2L���P��Q��^���c�I��$�w�e�j{���U)��~��P��k�h�ƵƵ�Z��|ʑL��s�G���������F��Mɱ��0�Fu6ӌ�C"�h����������J�����D��z��	Q]�ȸ_$\�vF9����Z��9���P���p~@?�yx�_k�q�Z�[���F��[�k�.&��m]�%g�� ��[�tw�gv��t��O�hs�=�u��:�d)	��w�r;�����*9?��o������B��p���]�ϒ��ؐ+��+��ɪ��\@z 6�����@wP�	��;~Z���S�&z�f�e�;�}/�E���s��s��yƋ~�&/��/�.�<�-)�V=��Y;����r�Y� ��[� ��:R����푭�;X��Ѕf�[�{�Q$��z�q����9xH�Pi=H2?F�}#V��t�o18i�}��=�F;HC�,V6�gs��V�������ɢ ;S�ٟ�ƏAs=+��f:޿x�!>��^�m֞Ϣt���$����|u�9��?�vM��ר�s�M�@�o�J����.���q{?�l�n�I�e��mme��ڐ�H��RF��qz��_x��l����!�1�0HlȲ"�͓i��G"k�4�w]��8���7q�4�P:!���O�עr����7�~�,b�ڋ��-�t��J��v�^������[%I�^����bݠ� ����|k���~��|�ꐦ�&������N����S	����2�u���4J�&�KEj�S�"e�`lfK���k<�H�H�+ #�-����C���gq�D��;+��K��Eݎ�Vҁ�ֈ+��4F׺C�b-��]�Yfw�n��oy;�Z�,5��ϙ�9��՜����&�9�c�:c�O���sA�x�"�%pzIa�<�	�p�� %�;���P;�0�~P�P ��9*��ñ���J�L���KǷ�@0�뀅�Z������M��irs�c5X�ж���b����Zcs2�4Zhv��D'����Ɛ��kmD�� Ƒ�F���{[_��)�wI4�p*�$�9?j���)������Q��O�&�x۪qr&��(;�w�M�����Mh�T��t^��{�+k�gM�Ry�L�k��+,$wJ�~� ؙL
���B4�cE�G�@j�0l�R���(+��� �O���q�)o�ӽt�H c����~�v�ĝ������c�ٸq���:����fi�ک�_�w�����������~W���95Z�Tм�ڇ�Z���k�&˟H^`�@���"�F��~���<J�H�&0�5d�h3�t*�t̜�9��]3ȿ�d�d�"�$����S-�:�u���.u�.HloLP�֔�ɧ�<�ɭ�+p�q��� �a��;v�U�$�V�㻛ƥ��z�H{;{�oO�C�+���le;�����[����U�Qc咘�^���A ���h��ߙ)����?���0�$S�W6��2���/��ʍ��(�F�<�	��؞Y��W�r5���w�Rr�,�3��	j���߂e�ai��tTa����ᾖs��X�3����Y�+2��	!r��yэKU�wM�'�7��pu�˿�
��yW�e2��f�ʅ���IV�I��oG���W��2���[���3}���~z�}^���$A�u�S��R6>f`Z����q\@4i���`�>^+�1MeÓ<�h��.��z�J�_��vL/���g�p�ii��>4y��d��-H�����L������m	O��p$�4 ��g�޲;�j�aw�ї�y qKL���z�G��˲$a2��!�������fxvs�G��v�Ϫ�$c?B�E���]�5�w��t-�H̜�q��\	��w0����4.��^���W�3�P�VI�d���⾆��3p�C��mZ���Y����jQƠڣW�E�!�Pȅ���kM�����ߚ8�{��<�m��Kv�� ��F#&;򆳭�2bf#u�� �ۚD��0��%����~�P�lO�o��j�"wz��Qw7TD7�g�'����p�q�P�>��	(\����Ji�Z|/��C��i),�ؖ��>��e����&:�b/]����<k[]�M����<��J�V���9�-06P�a��?b�nSm��	D�-*~�cܡQ<☘���@;�x���Mg&���zGJW��΁���8;׻�M���i��D�%�meA�7Ն�D�F^�:>o�rزv��U49Y��&O���[D5���a�y���Aj$�Ȃ�SD�bd�F�.�5&I����A��3}{�7KbP,2���s�z!�Ӫ�Mo��s�D7��c�`���P��-��[�Py
R!�Δl�JC|�u�6"���e`�4�&&���
�^5[�J����6ł���?b(�z�����-��w�zE9nr�p�����)x��w��F{`[�
��=F�Nj�!����-O][*�XK�XYMto�i[av�_L��~��6��iDd��De�/G6lL�Af&�>v�O� ��.Z��hkZ�y���	6S ��f�'ҟ�U$���ZE�CRe�d´M�U��Y�E�)��)��˥�Y�{�_���`�0�:@��}���Ri^A��خDZԤq�Ep�?��"��і�ǧ�h_�����f�ל8	���tz�C�W��E�ͫ��w��ꞛ&�
��^7w��{�
e���(5�§���p: 7	��E���p�Lƿ>t�s/JD�C��ۣl�[�s"HnJ�u�iJ4�吐r/yR��K�PE�(� �96��M��Y� ap��w�&�[��~O�z��Ls �kZU�$��	۵}m�/~`�s�t��I`U�f���@�Q�C��5��}����D�pv���:=�K?a�b�Y���9���O� �:�o�T��-?zV��J���e�*[�}�-���hx)��o���"�_m����
�?�2��n�`�C`Z�h�a��<؆`�Cs��'m�{�~�J��7c�e�,�:Z����|���	ۢ�S��{R�6Xv��\�Ԓ:�2�ͮ	�q����4�eb�U����J�~�Fڣ���;<�����S
Re����HK��+�`Z}"d�%|���6ԥ�,��g�܈+z0�P��?�
�C�����,��ߡ�'��� vUs4�
��^=�9*� քVךj�D�؀��H�ŝ��-�!6ga��S,ɟ:�]���Q&O�A+�rcg�>����t���V)���k��?���Yѩ��CFy�e;���z�}1�L�֋��~�[q~����3�YS��iA����I�lK�{4y5?,94o�"π���V{VDLG��#�C`�n9�/>���f�%����S?��j��p�_��%�7rdv���#�Њ���P��A�g1�����£|�ip�o�^M�����M��}�㸌�ɪ���s��������(j��"�>,H�M�輦!�W~��i��v~�?�~��2��A6>����L�[ᖛ�s�k8�)<(z?K��J�5��m���қ>�[��Y�6,�S��d���{��y@��`Ï�9�������Zwe���{�$���@��Nz�l���iϾ�\נQ�P�:ws�ǚ�dR~i��oa�:B*G؅TN�?����|F9�ֺ���d��A�&R|����@YT��Tc�Ǻ闄F�Bo_���j��3|u|�g��M���I��լ�4\��4m���(˶V��t�Ve��s���� 0���e��G��>�-(�Ż5��1m�n�!���NG�Y�,��/�W��_�.�k�7J�����0rArN�E��q;h7�L�ި_Jcy�>z�}(��@����<���{4\C���4�̈́7k[�QEYiXH�UF�v��$����O<�B OϿ���k�#��C�c�8z����+\��0ݮ�V:�����S��Ѥg�F�o��|SC�,��GQ��d�����o�~� jHY&�tz��R���������:��^��N_�},P����"ɾ$��ʀ�f刍k#��YS=7����i�J.���������-s��%���$̕d��VT���̣b�}��
����B{�����Y�1�܁�0&8�T0'R[��	�l��5�}�C���Tڢ�H:���`D�k���p% 
`����=�.&�= +,��U����$K%b��#��4p���3PO�V �i t��g0�U7h "%�0��m�J4@�KZ��ͳ7�8�2�xs���oಎ�knz���lXjm���I��1�W���!ɋC�h��4�`��v����sc�-�pMiWs$i7 5��f;G'���b�L�0e)ѥ�- �D^��=	�>���Eh3��Y�hO��z9� %$9"ytm.�o?N�L�/����k���gm�������X;�+�D����0u�y��<O�D��8{_�x� ֳKn���V&�,��@y&";Pw����u��d��,�ަ��*gb�]#cei-��f��#j�v�d�@�t�-��)Ĵp�}�׭-� $p�Fz���z#g[ƪ�\��Pn�3[��Hc�P,.x3��sB.:AV������eROs >8��ƙ������YN@����6��X��v
O߶��l���9%X]�kq�<�i�G���J`�S^��:��0���4�i�ٽlBk?�J'@����%P�������w�u�W�7=��"���*\�b7�S��^�eD��w������h�7�J�~c������`Q��h����f5/�@�˚!�≍f���˚��>��� ��W�Q!��W}��΄ >j��U��;��*�Ͱ�$�ja+�� Y3T�1��2��ձt�rR}V�j6�h��1,qYI�H����ҕ��,Lg.���T��rv=��9h�Fm�,�ƞ~%��� ����f$p�v�����!6�`���4w�l�]����<���`;�U ���q]i��:Q��Cf�w��~B:J/���j��&�4#�� ����������ti<���$P��	��0m�x�)�NVck���q����.Զ�M*��K�GxN��lJ���hL���ޒ��tӨ��`��)�1�� ��T8���5�[/y�\v�H���z3�"k�MO$L�/5G�y72��J�+�R��3�e!n,8��w|{{Z>��X��u���5(�P$�~�X�}|�����[��T`��&iᦕ��_�it
=Z�ˀ�C�S~����TmT[$����km,!�yК���r��^��X	�#��|�Zo8ȟ�-���L�	[�� �FZ"�N�Q�j�uO�������u�]�'�p��8��P#�L��&�O|����M慘sW}�����Ԟ�:逥(�d�*K !2��u�r=�w���l\�{�z�V�z�_W�K$��(�-�S�&wy�ƚ�85X\�a����)Qa���c�v���Ɂ��{"2���ߵ����Z����j�&*�r����͂�Id�#�A�zw����.6���8����̟�o����g8d��Sj�7,�!���-Z�N&��8��&x�b��U)G3��&�u5��?�\��}�^s��[w7O8���l�č��Qה�3s&!�z@\5�pc�C��W=~\�������(�!HXA8�7�Q�(�MfdH��d��'�������Ds_�u�_d���gb�R�^@D��g��h��y�u|�|PV�t=�הߝ�5��*P۷���"�d�]�R2X��O��*-J��J��M"�*�1F/8l�%b��[@�
�U|)��tP)�S��un���!-�H�V�K���ۚ���%,"H�%�~�?�t��
�f�u� �#��iԊ�&�a<����1b�/�a�I�s���+x�꒺6Lg	h���j�j���aX;����)��W�.��5|�l΢l�gPk	�����6{@��1R��am���Q,���?ѩO�Eo���5�JX��̱FNphZ��Z�wڭz/�$�۫k��?��MH��wT�VDgx<��jՔVܤAx"N���~��ĥ��q::2��G<�o�����4��ܓ6Q�-#�(krY� Bl^~:�p�)�92�Aa���#� Ytqy��na�[ �<�`,r��Uy����}���狩G�M"�6YTK��*Ye���4�A{��&�
$q���fU*�0C.T�tcpxǑO��F�a��V,�0�����}�ݺZ��&��2�D��$7f����⃧�CL����s=���(���lD0���*���|?2�[3Р�j�C
�:�~:���	TS���a=�f�ga�%�⣣0A�����n���b�����S𽬊J������v^�|�=�9��_����~�S�6?_�Dq��)߃���S�_ݸo!̒p��O=Yp�(��-�#��<8�U,ǣl��;���<l��_9D�-�����V1��T�
���.�&����oB2��-�T��AH�&:������ �ދ+�,#��t���g��z��MN<�)��9�7��$���6��l�b�ڶ�̩�V�v���)��^ōA0��&Lw��19�&BS1��rK��RG!�6�i�C���Fmt���u�.�l\�O?t�;ܠ*��v�f!*���aυ?���8���,׼ܿ������m���7Ɨ���e�o�JT5#�o�wŒ����\���l�"����?�7^��x2���DmHZ�n���~7�E�;i������X�[��ۊ&:TwZT���ΧrՎ�7����&@�{D��B�A�4�_Q����u��jX
w4�@b�.�f�Q�[���LS���X���l@Ǣk&�QM{�8��7��}Z���h��t�L���1}?w"�걔��:�q��;Rj` O%��S�X�csR(�8\��Q��%�2*T�A28��Z�R4p]�ކ?~��h~�7����3P�@&�"�[�S�u�8�s1�jh��bFخ���Sol��p�u��?Zt��-���-�� Lߡ��-��(;W����ε,���]��iݓfߐ$�QPY!��Eb��XF��~�ku.0�Cz�ָ�]W���l�
� �I��j��~D�kr
r	���J|�ТF�bVgc#t��`�I��.6�9	�G	/����$�5t�=X{:)���h���j1��G�
�Q�)��+jt1}l� �Ӑ�jo1��F ߹_M�trP�M�2z�����3��:0�?F'��O�[��1;jSjp�SJ]�IZF�m-2c�on��_�y�׾!&���m�!x�e�a�c�����_Zi5�s�\���]W�\@4�J��v�3��W������'4g��V[���k��cG���tLn�6�M�U<]zE�}������~��2@=� oi�i���4	�ʂ$-O���0��t¿�U'_��S�Z(g���h˭�-�a�Z�d�i$��:��7��)�(6I�"?|��F
C�g�d#�m��6tf��E'Rp�%|Җ��d��Qy����	͝�� B�a�/a�:^� �" J�- n��1��$c����C򌭹��w��=ZO1WerR/&�R���F��,ۋ<�L1bU�]�DǿJ��Yf5Z㹼��K ������|���[{X/�;57�����㪫���u�B��y*J����-"���^�/B�҆C���v�B�e�K�ו
 '��KH���L^�-�r��CH9%S� �� ���w�O@5��v��e'�8��K(�-ëp��Z��E~�����v�����E��{k��,�Pv��g0x��i���i`�j�'߻շ%���}�67ۊ�'j����D��ӹD���&�k˛�V��u�)���Mw3&4$Uƍ���e�ip�n�fV�+D��53�M�	���̐�)4)���i"���?�~�M$b$�r
Q0G�y
tVƮ�Vv,�a���A�Z���`�o��Wg4�!�!ekF\�C�)�x����Vx��b��<A ����e\hO�{z���A���� g�y�;�'\��E�L�*t$J���X&h��sZu�'�Q�ם?ǋ�*�;,�� ��$�BŅCXm�'L�MmELKq��cp=<E~F���T*�R�<V"��s����"��뤇�Xb/��8���~�2v�f� I�Va���3�o��/��G{Ҩ��d�!Z�D��T��`j�Pva�5�TN�>]���_�/a0��V�
�	�.����QM�՗]m2�@�� ��Yf��F�e���ݒ�����7,�����,�S�쐀m�y.�s��_���/}B��L�Ť�Z �"�pT.?,
CD g����Dw�i�[�v��F��jm�X��/H"��8�TJ6�:YH$g[(.������6~�Wg��&Jn1���t]�
��#F[H�Ό�|���LI�Pi~��Q��M~@X��B���3���4�+�W�e���8(�V�"��lc��DM!k�!6ϼ��ท��dCt�o+&G�f��?:�Z����8T���%]��R;O���^6z�++�;���d^#��������!LyZ��,n����U n�$�׮ȱ,?��:Rѓ��F�9���"��Q���q���L{jp�XK�T��8��娹9��C���
�I
I^Z�aZ������:�8F�S:����(��O�Q�����e��?�je9|u$o3�1�8r�%}�.R�ᆵLau��"*C�|��ԧ�<��f�E96A���u��[4��6չ��懮GO���<�N�ި�o�ۧ��{5�O��Na�SN���elf�m�Ma碃�)���C�r¥�M���ȳ���+��OF:����;` �ܳ�i�7�3�d����wQ}ԛK=�����_�/FG���'P� �����ò���� .��wƟ��פH'�����0U�������9X|0��9����쬈��w�v�=W��#gѰA�R�ٍ�=�M�
<rf؉2�4�|�΢�L�!=���g3j��H�7���U��I�^-W�8�Ė^ʈq�I��o6)�,N���P�:�#����W؛x��%��0C�́(�A.��%��M	/ut�1r�Ō�^q+I�y0x3v��&��MTqҪ�}�kQ ��P��h �����`�N���|(1b�,ˏB�	�i��}} mS	���T�Go�����g=�C ��*�C��z��({Z\~-t ��We����n�N0
O�
��e&��(8�r3JO�RmY��9�T�A�pjQ�L�-�����Zntq`m��?E� /I�]���n�0*ݲ���}N}�f<��݈^I�+VygBMҷ�n�s8y�i�������ڙYI��L���Ɛ�.���F���uTJ# ��v;7J��;gY�5	��>�3N0��&�����f:��H.��bn��O�5���.Bn�Eo$��a*��0�v�c�B��Eb�9����1/�Ig�d�<i��D�����'�����!����o��	�ZU����B�Bm�\1��fw��俔���+*%�1ڈ��D �LX�#~�N��O ���nS�_�}�ހ�LY^[�K(u8��3\�)��͢f���{�hq!�>��+�hy�%��oѠ���	���/]Tpl�b�;l�dV���'<��b�,� M�,�V�c�x���|��@m���bȶP���S�u��T�>�1�`����ѻ1�j�@�_N.� ����p��d�gY�4�`���hku�������?A���/���V�N�_Vtk9z�?g�' 4ݣ��.���j�!Q����Ŕ��N�,.::�tp��+7�ޭ���N%��8�Ǘh���+�! d6�t鑙:��@�K�>����t���q�St�����՚�Y�E��Nƪ�����⓶%t��̌H��/L��\;�:�%i�o���f2���N���v&��n�<su�%�T����;�੏�D�9�γ+r�M8"��
FS���k8>��JI�gc�A��UZ^h��łQi"�"|�8FRq�t;3�o�WN�T7��f@Gl�����/._��A��uAf��������SM���qc��8�-W;p��	�zw|���9_,��I��3:�-p��D����lz�}�n |17����v�x��+~����pU�B|����� ������1�ua�#��o�YA��}ө�^��^���!���#󿵚YE�O��H�O���X�����aB�$�&��+U1TN��]���Ҫq�DR&�KoY�@j�3��wR/ωC�oN��##���S�c������9A��5ic�9'܃"��M�?}��fNJ`�x�-�wH][-��vX3,�7��U�1~c~�o�v'V��qg%C��+�m�HhBU�=���@l?�<�ٝ�f6f�	ZЛ��\�s�G�ܗŗ�X��D	��sJ_��9R�ض���lp�����g1QE­nm���8�y�̞:b�W�#��;0Вd�;4��A��)�5�!b�5�Bơ">�r����0B�{�	��Y%O�) ;X�TAd�s�n�AM����TR��`�#CiP�w��[�3�������M���xFw���C)�?{���B[�n�=�)��lӚ�O��EӃ���<��;۾�Ћ9@�6��B��W�+�T�#�1L�m]F(�m9�h��8�k��C�%��x�� h���py#d}_O�s��oA�3�#]n�f�8)��Y��<�'QG��7��j�R!tSI'�,WX`^{E���2�d����/)6|�kq{���Mq��ޢvB��q%�Bu+`*��w����[X���ow-˚W��"�H%*Wt�F��8q8Q��E�.ez"*2}�f��OT��X&6=�bX.�!�(rp(z��=g�MM�iv>���a�1�M���Hv;�!�_���fKa�%4��Ni�ARq���DK���"����n����_��5��~?��\�G[��@��&$Еk6ef�k�ClW������+��iq�aG�q"�UG\y��; N*���lN�M+�
2<���NaY��ނ{s�F��#�X�ң���<t���y���sL�ލ4tw��+��8��A�c��9��X���U؏�L��%*�Z�wo�ʸ^�y(Id��n ��8I-�������t��X_��μ�T��~zP+�&�WKO�I�D����/qC���n�Ц���n����<#s��bp�RM���5+�z��.�L4%�4�q�:��c�����5'�zr��X�V*��s�ف��NRf5N���aľI�	59Ր��<z��:��Ҷ����`֫����]��|� %}�q�Q�+c��(�/���M7���T��d4:����|�!�#M ���\�[4k�+X�P�����W����>9�^��]��!�Ns\�+�8�#0VTȕ�����߃ѵ*C67.^�2&��[���S`x�D{}� �ͬ���ӻ([M�VVt�=���!�a�J�d�����T��nҗ 9�#Y\6���L	V;�=*찢�>�Q��p�P��5꼧�\�L��np9�1'��mr.k���ʙ/�>�4)1ٮ5Ҙ�f�iA���F��RCW�^Ў���HT��-M�O��/�Ԫ�_����\�"�� ΃��<�4� ��� �9_�Q�\`�+�x�z���S� �	�*{�C˪�a����"�E��>��n�)��Y�ؚq(�j�&�����%�%,�����2�����[�C=��-�	���@|��Kv��!l��J��O~:��F�Ny��3����H�d l6K84)��%��fG���4�@Xsv*p�:�l�B��Ή7�����X�؄��X����=2�
e��Ȩ�(������MQ��U��WH�����7�V!N_x�~?�j�L(�Ýı����B�k^F�UEF�T���i�5m>�^Ǵ�*Z�?~H����Jo�Q�Ÿ�e&�H�L5~ʞsy>{8���ӌ����	��:Eq\7��5���25f���F�� �e;l�qۤ
B�g�"���G!�R=�0��_�!�pB�3G,����*�,�(m��Z�R��Jr�7��L]�v�g�����GG��E����6�K-_��H�@
� ߠA	�b�^�w�)��v�-���s􏀼�CK��B�����Zz,a2�����������DN�����L�̺��͘ϡs��g�xazz�0�� �W���p!�����2xQ
�R
KJ��%N��r)�P���>�r�9���zDѧ��sZ����!n��$sd�[E��kI(�!��G�x]�9#jYP%h��W�7�>�i&�f�x �����s�j .�D[p�~�p�Z��6P�k�~��,5���=Vs��[���cέa7�&ҡO���*�^R�l?���S�a�ڍ�f�p�9��e*z�y,�Tn٥�N��� ˼ެj36�hשy�4����%�
,=��;�,>X�~H͋�E����_Z1s����������&��7�[���d���3���.(<s �J��W�SM�c��
_�t��P�Wk��+�E�	x�Q�p�p��.f���<�PoUЀ��|�D�X0���Oz<c�� ��0kgEI�������ޡ%wN�,N��΂���2z&6Fm*�R�:��*�CÌ7*��WB[���������>)q�t|K�����Xxa��6 �"E9���#+G�����D�\�E��=�,��ݦc@���:6��,Q��m;j\j:MG�{�����\�����8�o�#�O����׋WPU�/9P%ek��;c�A^d��}��tfV6[�O��_w��s%�� ����n%���~�n
�H��?�&ا����
�3�be���t�R���e9@���β|�'�����Ν��k�1U=�5MDK!�5���@�,·������'��Y��S�Yc]/�nA@�b�w�D�V՛]lz��]��,�Z������	1~i�c4w�h��ר15u�.�Ѓ ���d8��G#h�T��o �v=������w�kg�!�H��7��=Fsaǥ�e��b��IP�.T"���a�`5e.��OP�Hf@�p�$uv��SZ���t�x�O����D����w��&+��<�:C�~��D���P*��d�*l���>mw��y{uR�/�r��N�/�Gr����yh����9M[<7X��_����C�l�&�Y����c�@�i�I��յC�w�I����B{����?~�#dV������VZ�NN��w���4œ�nWy(>��E\t荘����i�3���;�?�\�3��ɧ�r�ұ��*��2�m�@� ������S��n���r�~�L�1t�w��6����P��с���D��Ϭ5����z�k�k�80�<��&&Z p29��-��Nj|��������Yʺ�X��DU)�v�y6i�dG��b�s6Lf*O��D��l��/�^~\�]<�e��]�wh���'���޽l����x%�{C_�~�_q\?�V���_^!̄*y%5~N������6��߆������z]��_�jɋKbT�"�|�����4����-��-���w�E�V�f�x�Y<3UM�,V}M\�6F@�R�O�j2�q:�]��JQ���f�mw��KB��A8A�P�����H��8nz��cx�a���$n�DF*�b����x�l={|����7f��\>�&���b("8��>���^����A�F!���������bⶭ��m$Ry��S�d��';�~$��/��A!�uz�L�V!���N���ꅽ���e:�P�o0̵���Yx�3�x��"�20D;����|��N6<� '/��E�E��Jq�\s��C�a �VEU֝��\r(��`Èy��k��à���+0\��Ԅ��qӈ�#'.|�j���DO��h��t�Ӡ��iyf���Q��F��nJ��1�i�g٥�f��]*�'0��"���٬uۨpO��b��Q3nu8͹/���{���� �2w��,�0`���:���}�k@��L�`�`�F�h��l��tz�l2�f�LO956��9\�1�8�P7-�O�]·ݯ?=/��5LT��Jבr�qp�����mP�-��v��V�"���Q�w��6@��g7t:��$܀�q�o����6�J�Ek�����h�|�6�E3pi����'�w��)�0	��ڎ�VM[��4���R4Q�cC̀P(�=����z��
�&N%�k���t��ǂJ�]6�(�K`�A̿�U�_�G]u�ޔ-[�2�x(OT��i43>tgS��J�Nk�\�:��*�� ��<���.GSE.B0<؉�ä�o���9������j���������Ĥ	�pC�q��B�b��b��}�C�Z8�6y$Q!�Ҹ�_˵�ȫ���9�>�I�(�i��:�ɥ�Y��0�����6(i�Nw��/`�IaxV��x��}J'ڐ��7��`}|`
f�s��}i2� ��/H!�Η��W���K§9�3���}�#�E��-�I!�W��q|����~ҥA̒��G�lI���1O��
�0�}���G�-���vX^�F�_J�(N$<m`.�b:�z=�rʘ��MNY&�ώR�o{X"6pe�}�|?I#\z��௃����:�*Z3}-hi��`?�����<ZI���K`W���c��6��f��߄��WDTX��_KHr���l)��E9v9�xM�s��'��Hu��@QŠ��dG���?l �	Q3�Q=C��8��DU��	^ك�B��(���&�ũ�A5imQ	]��[��0��f���2��'y���*�K�_|�)y��m6} ����R%k,Ylg_Ϻ���rB����T9o��[$��>�Q\�}�'�9��K����[��i�oWl�3���c����u�}��X�=����M6vlߍ���5e��7:\��Z}�d�ǋ�L3�*��� H��і�'���%s~�����M��|��rٙ?�r�Ñ��-��o�Izs��Nɮh����v�u����V9ˀ�C'^�Q��p���:�f������6���!=/�yqn,����>���Zͽ�Y�v=sK�Ʋ�$��2�՟6�#���/�V|�̌gs�bbF�����<�:�����B�/��Z�B�G8�S�8m`��L�No��CW2��I�&�ov��6�FR���͐Ȍ��F�c�οP[W ��X�,a�zz#i���8+�N�`B�.|J�.q�T����f��X㞓���@��	� �QI0�/���/���V����:a���OT>^�'�0f���`zfA+��jX�W��J|���-���i7Q��S��2��w'6*2 $�?\ow{�dǐ;U[Ǥ��A�f�����#����̣d��w��C���6������(ڬW�BE��"�^ݳi����W�2^*y��(x�����*�|-�^�=&�������	f���y�C�����K�	��c��-�X�ԸUㄓ`��|{�r�/kx�峠�<�X��A�˯���z��Q��=����=�}R�oY�ؕ�V�;-��D=+��I��`$8H���F�T�Y奇S�S�L|��	ܜ#��/a��V�j_����WG{-��,��PFR�[|m��@~ɿi"�-Y�PӸg��]Q��Mt-y��f�l�D7�u=�}c9�3�O�/K���)�&�7i���0��$�h��j��9[�$����P���_mn+����=��o�W0�L�im�^Y���ql��K)�,�8 :��P>s�"P`���b�3���� ��`��� ���h	�4��VT}�z�'(�7���J�wT�y����$��_�I�F�$N�y�9��������;�#MD�~�uH��H���f~EƢxI&��)����i%��i��zL�Z2F'�����e$�ߺu�%Έ�����ͨ�yp���oA��e/f�M[݄%�ɷˊ��Ճ2��2����f��B��05��� ��a?sE���~��B/P;���Y�T�z���a���95�% nvoOM�\s8��_�QK�ة��.���uŦb|!`ֶA�m��ݞ08F{��V��q�}W����Y�Z���!+�8��W�`k\*1h
�3�C��3��zgw�.X����I�.���W�I�p6ղ׳Ǯi��҉Q���R������u�d���kׄ�\��Ls0]=���-N")��WM9�v�ywٯ�{�Ũ.��tis���Y�|f�O��CT��9<��9�9f��F��,*|w-yr����c��-30�N���Cr�{��7_rڗJ��֧���~65.<��*Y�����Ƞ��NYő׫��[ɖ�xN���cPD)��F�e�3�M���1���D��=
�f�#m�:+3�]�F�)@|�6�g���R�A" ��)C	M�����m�jNT%��\X�jB�zC���v�+�4U}#�n��I�g��H��h>�a�nr�k�%�<G}.��mvr?����i`�L�{ܹ��NĞ�]������NC �Z�l57􂘶�ƪ��q_�"}�$��B6w�}�Gs�~�Ǵ�e�V:�dFL���U���i�����-�[ AB��n�,_���ߍ�����A"�f[�WC\c�d��*�����Me���8��c!�֭��g؇.�=?��Rq-tiXԒO�\:KF���U���=`�ԣDdH�#rK��5o���",�M�I7��� 0�2(�	4B:�	�4��}��6D��Ӟ]ٗ;lWH����ʫ��u0{�;�W�)��J�3�6o}�`Mun ?Gr�L�\�_ٙS r�{k��E�L�5��5�s�p�?����$��Q���n�x�F\
-���K��c���:h54A������;��2P���!?�"�(���]:M>z�ƲP���nN,5j�N����tVF���C�(ߣ�g�1�h?�;~;ѷV/�Ɇ+����聍 ���[� �(K}�L�����&W�	lyRfP�+<�g��|{<�ii��z�tsrb67	�4(8�0"ճ�{4��=%�:�u�g�!����*��Y����g�mњF�4��)_m�!�"|9��˼o���c{���{J��|�j�j�&�W�b��^���ɔ-Ճ��	�� ��J��
��R[��ˆ	�J���`>��z�;T��sפ7������dJ��%����U����j${$��sD�����D;,
Ŧ�[�{Y�m��f���!q4�v~ ��D����w�s=��}����fk"v8w�
ۄ�y8��ș�����p�x�!�aȿ_p\��,��|��;��a��kd�iD�V��T�w�F�둰��� �9 X��i�Ts�2S���/�D���m_hF��)�o ��1Ky�u}X��u��H��χ˻��80�G��ZP�8�[�h�C�$�ȷ瓼q7Ať�������*!�Ű �V`�rXc��'Ο�R�S����N��
�xq*�O��ПD��E��C��J/���G j�r7F�)�"l���0��jo�I���cH/�O��G�d�\�y���=V9�^݃okA�d�*�9��؁��[� ���?���Ќ�X1�ԟ�
�+�{�-���ob� W�A�7���J����l��v�GǬΝѪ���|U��v���PA�Z5�
jl-$�G�0T�ꄻ����Ol� �6��>��~i���r�U:Hd���>�+������#�A=$f�k�6v��W����A�kv_�(�φ��0�Ӗ�}P�y�:��I=wk�{2�><�ı���"45]Ϊ�	bA�i���|�̬��I+�4;Lh1�P��4M!����Ѻ�>�a��Tp+���x���S
������vd|�#;n���¾J+Z%�;�7'ʐ�^�b�L��3%,�F.l/N����Kiy�tz���.����ݬ���H`n{U��qwΐ�EQ(��I�{�Zb�E�	I$C턖�|DQ���2��0M��}&9�Uu�;�4���� R�إ̹�P���~�dT�
�`���/;��p_˼�?��L�\G;��p�hM���a*������K7wR:�B���ex	c��i�\ֶ^g��
ƶX����X�yk�Y�4�\��L�!q���u���gV�=.iϺ�`[a�:J�&�1;P���\6�����@&��������,�����lZY�E4�8��˻��'�)p����[L�e�L��.X�x��m�ܲ�R������3�d>�6.������Ӱx)�!��z��@ߧ�ݻ�p�w9+�'�s,l��S��5�&��ks��� �M�_��+v���V��}�' ���j�쇳�_��J�y��M��M4��<�s/�<��`K����H��y�b�||�L���?Z1�!�^4�
�= ��p\ŝ��?���x!��3)�:��|"
��p�k��r���[��;m�}� �����:�����Nw�j9}�T�jR�%pW��:�S#��PaX(�	�:R���6��8	�mD?�m���ʾ�;v�20SQ&���~3˄�y. �Հ�߁�2�\������I�qe�گ(ж��p����6�fT��������!�LL%t�z����]�>^�t����86�/]74À��.W�&������+��㧋��sF�*�!��؄���+��9��׻a}����!�%�Ǫ)�]�8J����89�b|� 0���4_�d���� $�X4��������YTYi>�L�����]�I����-/BG�9;����}���Gfw6�f��05�%�,PAt+��;���A�^�VCB�f�����G^�L�*�n6� ��4h���>�=n�Ε��:����b����s��(M�v�cO����~�27:I�|��ʜr=o1\�,�u�t��Ϗn���C ���K�q��S��v�R�Z.�o�=��X�
P��K��P���"�L+>�6�ט،3\ձ%�o-��ڏTs�
z��	4+���]���B�! }���)���K6u���q�jck�$ :g��V�oHf����h�f���l�齙�N����JRTjVtQށ��G��P����"_�ť�-�$5��o2�R�S�����n�8���gM�j[�c ��M��Zܺ�,J�O�&��X�O5r�vL%?R�~�I
�`v�I�{-���CD��<���~��:r"���1���0KU���S��5��׀C���v׶�?֟8�>.P�PFU^6Q��c#���餐G/�0b5ugS����ȹ���_�h��S6�$W,����N��� ���%��>��&E�Va��^-���G,��_�s��\�qz�Xă���ꭐٞ��w��yn��k��d�c%�9T�	�[�~��:sZ}.Ǔؚv����̫꽬�o�F�Fi���S{ZNj�L���y�����wq��>z[./�O}����阳�����A'���Н�5�� )�n�Z�����Q���!�_k�Vܒ�ysU/��&�c�a�dRp�N$*[]����L�8�A�Z6������R��5��[BB����'��j���9w{���I�5FL��e���|
E��u�E���h���Ԑ�W�ɦ[�ť�g�}�`@�geɁ葩�)���~\�C%��uy�`2u��-�n�~ ���%J^7��K5V�޲��{W�h)��|���*Q(6o�׽�Br�D�J��+��Z?r��3^�f����Py/|fG	<l�޺�)<A[����hG4�� F��&�D�'qHe����[)�e�	-�VWR��c���x%Mj�u��,1Υ���� D���||Dl.\Y�x��7(����\4�O-������8���e��?^^�r!�q�b������/���I�	P6��0Z�3Gp���g(�/,B���\�iϏW2#�?
\0��>8G���"q
��q�/��o*���&rT��g���L��j���d��+EA�1ί�?;|[q�o߆B�U��fP�&o��[F���
\�K/fP��qA���b�~�<�^�v��0?s�Zꞇ܅��AD��?�"j3$�X��s�r�	D|Zj��Q��7Z��x�Zm,��*-��1�6�*�ŭ�auFTo��x��q�E����������O��])�#�w����zj�*���O�)
��w"��5�ČdM��h�,wŮr�,�S��ʬ'���Y'`��5��r;���N�:ARG%�ac@�19Bc"7������
��A"Wx�0��l:�JߤW8�v<�I��ִ����a?YhiN��W��}��SEQ (-hi� g�U��8��)w��`u쮁���������2��6"Ǥ9Ie�ɲ�΀��6�H��v��߇x~��������[����g(�p��vg����p�R�����9M�	$=e�x�MZ�9��Qr'ZwG�Dd1g��Tn�����[gf�oU�����ϳ�n�`\��Z/|09ʂ��T��u�LL<�z�I���8z�O�,<p�;[�C�z��L'HƓC�@R�3�w%�f
�ܘ�ڜ�MЄ�n2�M��-Mv�{v<m%�[�A�Zi�a�Y3LGzL�0z0v�}�Z|�[��fg�/ȝ^ 7+�E�0�l����ڕ�1��G�A�!$����[�?�6�{J�{�kҜ�z�6� R�Z��/�@���6S��E�R��]�aR��7-8Nfv6B�I��d�D#����������95�3�OǨ�b���#^Jr����L�:Դ��G�C���%3�1�F�;V�6��;�o^�v'T��н7c}�c�����+q��,Jc�iZ�����|����[�\x�y�De-��7���I����k�uވG �fez���G���7��ĮSAٜM���`���U�s���ƧY��)'��	*�oq�+B9����ҊQY���M	N_�d���n��k�c-[��L���4�
�{tx�������k �*3���y���`���C�?u�v���ں�0C��>[+�>&K�g�x�f��ar�%fH a�J㳉Q0q�1-yٷ<k�y�84���Q�^� ����{4.�خdW�;��˩+��"gJh�g�	�"/��E�V��5z��$}J_�^c�Hnz��mX��S�l�G.��[[�A�[j��f6�W!6�G���t��w��n��H�u��ah c�+(�w����� [ګ��\@h�K�]i�ޏ�:HC>�?A��&���Z)��جP�1K�q1w7�{���Ƈ��O-z��ue�U��	��*|ª�ٿww!�D�x�*ȃ�?���8��i�Ȫ�����C�m�z�i������G���g�x mN�'w����K4�Y{�,�>���XٳG�+�̶f����o�?Q��ދI=� l=��kY�Coc`��$ };�mK�ë�{�ik�F��H�P���B$���]����H�#�G��Ȱ�ƛ�0����z�:|�V�'�e��H;׳lӳȍ����}Asܶ�Ђ ��'l�1]~���9tOu�q\�����U��3z�|�yIxm��$e;uCXJ�6)~�#��@��ĮQ��{���µ8CY�v�|*}�o�8�����0����F�Ye:bJ��k���v�њ�][y'%%n���m��Ҩbp��.T�pa�Æ1�Ժ�ʩ 2@���^z~?� ���34����Zr_��*�����T�.z
��c���@N]��2�8n�s�ia�tx��)5-�[yR��2C�]���������;bx4�kG\C�a.^���6 Zv�=�,��o�h4_��78D��l�j�</���aV�"��`�L�D+e\��#�G�(� �q&����
rݳN�����{f>E)oH%�Z�Q�� �ߧcoX��L�J�M��j���˥F� JE��:"Q�w�)�V7Ot��?K�DkXEP�>�ؔƑ������%�(�j�!���P��!y�c�cB��!oKp��_�����β�g�	w�6�5��Is�
��#��\z��X�|�l���ӿ	B��,�6��>�	��:�N���������	��G�չ�Vv~���E;J�R���,�%���.���k�ܙ���	j��XF�<��ucV��p'�E]��$���1�h��yS�=���cQ�w	h1�;E��Eq�����������uvO�(�u+H���gCj�x�պ�'�6{�[�>���3� ��K)��D?��g����h"���DY�R@�����h��Nv�I��Г�u���K��K���G� 
�S���+Q����:>3�$(��h��P]��ړŀzV�r#\�	|�z�,��OBu���e`��ѐ�L�eڱ]�k3�إe$��5��;��&2�98F�]���[���*Z6Dg��:�.��s��p���7��n����� �Q`%�>P�[��{�{<^J՝�|*�;�?����P',x���0 �C`�oE~�F�Te� H�+�^�!5��1��|
�S�
��&��*��s.Z7�d^��➤������^{ ^��u�Nȹ(� �G�V��F�ENw��:*��k������"��}A�=F9C��a�᧲���JZ�O&��6p�����B�7=��Gjy͚�_����!��ѿ���Ҏ�!6��{MJ�U��Ѓ��E�M�{ja V�W��)~kБXFu���ؓ=D���L��
�=��XHtsZ�	���:�j�]��]�4�����+Q�n~`���[��]b�j�׹�;~�Z���uvo�sWl�x�A��Z��ȕ�	��_f=8��	q)��9���@P��:��ƞ��.dq��Y�����z!�˵h@DL�����O�s�ü,tz��y��>Be�3{iGH�o��@�~��j���<�v^�"�¹:�wO6R)��t�f��I��Y���E���.��|P�F�(�9��U����1I� m����"Z��V�=�	�8�Um�qL�@��{����s�4rG�M'Y��K�D�bC2+�:5c?�Qe�[k���_��o���9�Ui������T�8(��oJ��q�����V?�(�0V]G�P��bMm׀&���������|N��mXڎ�o����g�%�V6oc�?ԇ��Ol����h�o͐P,�sW�@H�ŃTde0����%�`� 4����7�kw7*�tn�+�:�>7�H��iG����eY�[����
Z�wډfwsI��Vy��{W*����U�1�;�k�k�uWv�P�,��:"��V�i>w�C�p��'8b��'k�zM0�P	�Vd�%R0T�zZ�uݪ�T���Lʋ)NM�G����)�X��E�Z���N�]�N�M���՞�k��B$��-�D� #�XG�y�d�z��ER��1Jb�����|v'��}�#����<Kt�~�G����3q0����$�I��O��M] u��u����=n]7n����S��Ƒ��|�l>*X"����~F�?��ܨ��ǃjX�+���^�Q�&4�Z2K6)	>R����.�l�����e�f'C*��?��{���'�&��P�ᄁW�1P�q �yQ2VF�KqeM� ])௃�u�CeO��j�%lMU�s!��-����K��?m�^���	rī[z?�[C���y�Ip�=V��/F��yC7x.h���hWtN!������/B�[�W+���g�h��O4����E�/��L�Z��u[3��S�X��5�Q�U4�Ob�Y����EoE2�$��ܣ�#������EUE�������p�����rDq��x>��wo<gyIկ���O5 &%Fd�ā=�Z0��y
dr�z�@�(�,4s�q7�U�]�j���W�@>��k�p�l5;D��ǧ�`;��8)��R���T��ÆAx��w�d�/���8��x&<ᯌ�8_��gU�?"�
�PT�CVg�r�s�={g�ii���7�MA�P�z�
�g�>Ė)�;B����h��D4�O��ͪ?;M��1.ժz9��D�������K���k[�T���&�ِ��?E(S��J���{H�=Y�	�W�$�p�zá�IH��(�yJ�E��I������/a�����X(�hɾ���p��E�Bj��n�L�!{�I�6��?���咋�1j��ud��iC�4#����V���ܭ:��=�=���_�$����9	���)������xEJ)�[�VjP��o����D�w����Ҟ��9SD&�Y��t�
N� n� �$��n�� H,
m.;��}w�{��F ��I%��y�M����N/��n,pTȐe�!\n� �!�ס?'�	l�Y帜Y������j}�4�a�MG?��&�<s�L���2� �\{�z�^���i�A�6!:-��y%6k��Y�"�jf���;�O���W�f�]����vJ�L�2@t�܉u6\��bh�v��L�u��=v�}涚�9�#�n�$�Y��D���o+�]�R?�b��e�KƕX*�]扤D6~�,e��s������: �y���L3�}���0�����!MD�F����Z����*|���lb�=���=�m��S�2������b���=B.��T�l�3�"�q�vM��'n���x�Ȳ-������xO�'cc8H6R���
����h!��#
f�c����R��ӳ�k�CJC��)�>h�
���K����*�����\9����:�]㍏�53m��r���� �;-[����DB �$���9���Su1��!��"[����(
���+�Ҫ�0�c��)�ՠ�-Ue#IT��NGպ}�Q)�i�X��0�m�[�%7^�6�\�j+J��}Cʝ���X�0R��� �R��7^6���j�����CE���e����P�����U���ēDJ!���X�H�]�mF�������x�(v��:��Yu��o�mZR��:b2\tJk�a7� �b�"������R�uv�]Ú=����Ѥ|��X[Zz���xѿ>�^�U�$�m�l�6/"`$���wf���N��T���F�a##z<�k��$bqQ�{V�F��y�����~|�wF�������=
k <�
	_��1A�f�s�ؤ;B^�'��ܗN�t�%���"�1k3��,��nY�Xğ����ҋo���3.t�0=��W�4	G`�q%#X����m��O�H�����9/�ƲҦz���.�BL�d6o�D�Q��q�j�����d;�?��O)�[Pc����2�*&�Ƅ�67�P�]�ѭ��}m߯�/� ��x�����9��O����ȫ�xC�[E��+"�t���!��%�7.� ��^o��`��	\�o�<�1����	E?�i�[��7I��P��Z1����zl�ɣ��!� P9f��|��Y�d�K��i���G�����O���A�ar�J��w:��4�s����\O.wt~԰:�xF�?pWH���� �)#���퍢����V��,�q�}F�����`׽b����W��I�Codﳣ�%����#y�N)�ECä�u�x\V��}�_dfH�N�/�p@X1N��8o�Wğ����-M��c��Lp�Ԫ0<W${Z�q�cB7Zd ���=�z�<"4-� -^���s�$5ޛ�Uu��$�l���:yn��K�Dp9�|���v����]���Ey��@��J�8���q��$W��b�Q�z)�结�g�)]��ؤT+���[�W�����Pl'��WX���0� Ò,x���-�R%0'�1���&���U�`���y�c�N+�>��r�^�Q-yE��A���l��ku�I������@g�&����Tp�rd�_�����v�c-�g��3��r���z�-?�49vP0s�q.ORH����P��;H�z�%�����,G\�"��1*������%���n����ҳ��egΦ�#J�(u˻ר����w��{���%s;���\�p�9Hۑ���W3׺�����q�b�$wP�/�-t�`�/�Q^������G@�&m! *�{}�h�x��o�@��N�i�<�Ô*��*�x^��Ĳ�1p����?O��j`�#Y��e����S��o��gK(o<K�O��4	���i%��O����I�H#2�d.���E�
jP�h���H��`���&V�g�UT ��1*�j��M�K�p��ؽ0�D�x���\I��F�
 㪞o��Ƃ|�mB�^�q_gK�����o�=��*3SV����K���w}|� wF��]
��5�3f�s2\z9f������n��e��!��+��ߥ�^�-7��4:=�mC)��m�W�6�7wS �ww�CT���)�F	O�u��Tf�pp3U�'����il�������9o��9BѤ��R}�`j�%@l�H!�E�z�CHD���9$�w��	0�ef��j���f��4;<Cn��X����>G��r9xV���]���V�Z����gv�`�c���eA�b��-�}�CT���аx�_^F�=%j����1���g�B�b� ��j�v��Hׁ����(���t�ZpK"[�lB�Uh�K(*S���ja�˞�i4�y��P%����������J@�G���c���2��c��}^��R�QP�����?��D�\l,s�ǿ��h�<����p7�ž$7�hh����֮�e��i����^�k\d�`�vڝ�9�/D̹�|�l1ś��+���f�1���j�$JK�;XL34>�{&RD�{��P��Vl"�	j]�������U���%�zCiSUd"u�ȱvoS8��i�t�r�ϛo})�`�^���sד�F�%�e�x��*�4�o`�(��&(&F&���c�ʹ�y�ťA��4�>�bE�o�X��+2�F�a��*��lp�����Y��5�w����r�L�ShhYm�v��gM�w��p�M�ﱣ�H�)��C M���Dƃ��`B�Pu ��EK�`������X��,?\-����� v׳#�H��� 'ܨO���c���d�%�s_���64���-xZ		�ǆ���.ɳ�5guD�P_�.?��ݵ4��$@!9�K1��Π�ZfG6ű5�G�o ����M�wi����W��]=w����� 	�x҉�&�P�Qwu��LLk�D~��3�	�����!��V�7�pf��e !;WPы�0nŢ)]�B�j@G@'܂�*-��Ւc�w�Y������
���
�$`?��I������5_*`Q�b�(�b˺�|(�6K�=n26�U��S�ʡ�7�	z��)�cZ�u1^��N�%��~������N⊰���/C�0����W�$+z�@&Ls��z?}:��Ao�%����Yܒ�c���L�$�1�bwrT0�žY;gQ7�B�¾�����
#;�1VU�>P�v����?��#z!���5v����1 Wi�����sk��K�$<:=r �쩕��;=�W��[��g0��S���cT6�~�H�t����(`QУ����� �C*���%�x�c{�'�|'<��ϓ|i��R?�bN�/�_We@����cРU���"��_��[���.�	nm�"�*���H��?�����r
D�	t&gtEᄐ]d�N���E���o�(�>�59$��}����V�w�������'C1����lߵ�Æy�~��s9�e
��E�-����IJ�+�4sj6z�}ŏ�>�����2� ��)3[-���\
9��T\�:j@����X�foOm?	�ʲ�YF���@]��t3��'?�&΍�;�!.%	)2����F'���K �pK��NZ�R��@��p=7�)���C�3���z�Rӈda��������C�A��9��eV.'M��?��X)���obSp��?��"����>�4M\{�2��4���\��b�w�*����� d��y���̘"�r�C6b�:� ��X3�;n�C��&��f?��Ρ�ԥ���9�����z�+�f��PT�.x�/��!n�@ܷ��1�A?<��N �>"G�����.%4������WX���a���i���^d�+@E��/� �㎈<���t�sS#M֤i(���8�+�zI�
tC�b�g�Lಗ}��m��L�E�����G��I���WC�A���Y~� R�ݒE��ծbc�1�	�L�T���c�Ĵ�Pk[m���ʷrT�H �гO�bx�i+Dm�q�P0�n9za".�4+Kwٻ<ak�y��%E�`�q�Y��T��[+t�QRz#}�L�����o�x���N��G��̦�M�f�!�FhN{��ݎ7nQT��?�G��+wM�c��j����v�T��������+����E*ؤ�E���/<Xn�$��+j�n3�{֑:�Jx1_e���I���e�Ŏfڬ��)����i�F��I��U�p��`p�~��;������'�"4n҅��g���r�p�Z�������`Bǝ����g��3� ��"��>^o��n��:���YD'�o���M�y��tSHCo6��:��·�He���6�kiߌkM��/�8��ߤ�Y���p8��%T��k�5��u�gKm����@�Y2�Y��)-:~~�4�q�#��������j��gF���؜��������F��*����	J¬7}�jU2�Eh�!��j��v$�?k;��ߑH/n�Z��7	k��K�N��H�S�$�<��`����84!��to`o+�Q��tA�8Z/�FX�}(�0+�*#<�붖D>��(�|)Ý�P|��@(��AHf|��۟'QC͐��T/�|v^�KW�"8#4 p�"�b� �J��</,��K����������e��ª�=]���G��#\%pX���V����h���yp��W���pmDm%�ͦ=1���1�l߈��Ao%�|2�q[�K�ǃ��# ��;=�D�P/3b7!Y�)�"�@�w|�;�k1���j�����+�������ܜ�Ϙޟ�E��>+N����E�X�8�h���Wf��B��l�6<����+,������a�T˺$��X�?�-y�i��k�ȴ�8��i��y��T~$?������5w7FU���;�G��/BEDO�	�ªg�ܑ�Ν��%�I�G����5d$�4���j�x�&QT�
�i�Nas!�,�������a�՚��W�?���0t�0f��4�ڰ�s��o����8D���%�G}@�F]���l��n���k�["����?�mb���:� uHSے^�D�j�m�cQ��uj֦���sX���Y��=`a�a����5��>�?�4(�jEN�oNV�F�U��׫R���FRf*=���g�AzV�(
�4S��_Z��B���=�	ЋӐ3�R�J�W+�ٽ��}$��p*Ic};�ء��#�y���};�eAQW&���Q9=�c�S\��8�x����\!+�EJ��gC�e� y>&d���^2�Ks�D	�;�<o�Wu�
wW�I�C_���	;y
�?���E���W�b���"m3��*��f���	k_�U��F��%|<��_*�X��bT��(}����'���{��O��ۑb��o�R�#0У3�l3O"���.��;ӕ���M���|�Zt���z�������k�>7�ze�J�z���&V+�r��Xۏ�Z6�Ძ1m�,�W��C"cV&��B��ᔊn�厧:t7��'\��5���B�E���+*u">�d�y6Z\ S��?�4��_��R4��f}e��;V�ĢW�y���5s�_�N��&� ��],��@�ۢ�`!��}�X��PA����Z�(�)4J��I�:��=0�����/,
��pʙ�R+v�ⴱ�ſ�����"���>%�Yf��Sy ��˲��a�|cJoh-�H�-bz�.��� z0���}�v��ޭ����oj7�r#�*,�a,��x{�5I�88Lfu�k@��q�#�j����9$:C�E�p.n$��d��[��؎A�������RK��9��)|;5BC�Ecʿ���T5���^�����0��<>�c���b����zr���yZ���Dx���i���7��N�ݤ�QU$������P�8�9=��1<r��U��"�-�6O�6�0����4s�)K�pQ>�w���d�3nע���J�/,3:�,�����1&(�� ���s[��'?
R9F�Ym~i&��;g�K{;5�/�pT룽K��' �sS�P�V�b���w���#ݣB211>�d$O�Y���H@��\�;T��K#^��1��ig#�HsR�~�<H���rPeT����R�Yz4�(�KD��R��3�ڮ��CE��&�!�:���9���R\tց�+�{�P�A��Ax�!��P�}�?0��tQ��#�	����j.��@���4{��$��L��!��~�:EL��`�!���r�B���RB����LU��@�l��D�t~�'}��=���;�g�!E����C'BT���%���"�⻥u��t�H#�S�,ZNy�`c�F#���>�47�Pu#�*���\�z�����x�*2T!!1H٪�V/(�#��=-jw�f�.z���/�2�U�&Β�q����8,pNF�!�����?᩻�s�G�f;d��р�+i�r�e������tි��R�fک�;G~R�>�9���"��J�}Ҳ�r��d�$נd�O�	�2�!�C+x&3��ͮ����8����K����-�G���Ă�"�v 'P���w�cF#���k(�dwB�v*�)�xk�ny���Y�����Ĳ�q"���,*c��p���i�w��E���r.R�@��@Bf��:w���gq��G2�'}�����6�.��������f�h(�bd���H�7"L�����m�t{+Vf���6��m��$a~:}�R9�
-�k��I�ˢ���E%�7��ͨ|zէ}�p�u��G��O2�8ꉻc�e-���om|�E��<�l����-Znm������J���4��:�v����f��2ޠ('gtc'��Ñd�|˪�b��3�3������:��9���5Z�Dɟǆ\�b��!��H�����w?M�C!���鿷�ϴ��8�{��Cs���l��X������V�����r�_����I��b[��~�>�4G�A�p��a��h���ȂKN� ��K��%k�m�ִ�gl!b+��<&��ߏ�da��ia�у�ш"1�o�R	3�ĔO>^;���^��Rg;��z��n����dA&�M��E3	�
1d�m���?���M���ݧAeL�4��6p���E�NM�y9
�a�W3���s2vζ^ܿ�Z.DX���7�p0i�?�s<P�5�LW���9N�k-+s�dIz�3��� *���QQ�v�/��tx ��I�.?�a`��zk9��h�/��VLu|w�A��cϛ:��Ad��xE�4��8�KC�����H3���,7�ƚN�4��Q�~�Ǯ&E�� CH��4ʌi���yɲ.}y��	O=S�P&s�G��!�b��ξ[S.m��?��L��>��|ko;՘ulb��Pa����6�uZ4W�a�o
G�����@(¤���G����=J���>~��G:�p�^���#�"}ZV�z�Ð�<v���[i�k.F5|>/�wo	��}[q�`ZT�������\��������z`�6�T�E
��:���(:�<w_�u�C�1��(�'��򂸔�J��%�6�8���.6��a�O�r}cB:�8��)+���ڇ��
܁��M>,���e���]�5������=|6T7fA&8�)W��vUO��[s��N_�����u�.�>9)h0 *I~\��g�͘��?%Ҿ�R�hɕ�n7�+������P��bع|q�,-��*)K��,G��ib��sh�6~	�m+��YZ���iP���J���������V꘾���B9��c��:��퀣Ϊ�T�R�}5�����H�'&���,�~r�T��)ȍ�3�/�j?��l���}w	mq��^�+{B�
�5��5����Hm=�ʦ�M���iY�
f��v��9�*��J�R���3L��%����:�r�?֬70:���h�8M�+σJi2z �?Rо��J�ݡ���$\=g��w,{����M=��|��t2�4�U��2
^L���lu�F�[���g4�?��ۭ���d^>�l��L�����!��N�_�6�F�������7O��P�����I�.�,���ـ���(�-A'�b�S�E�A�ޕ�Q�b�O9~&E��*��G�-��!�&�?>XH�cE>�Y�>�K����9z�0�T���c9�|������׌�.l�i%ǠI���|70��+ϱ*�Dv[����Ѫ�F��5��R��w�'&]8���|��"�zF��d�D �����}�����ѹ頕-������ �&b��w��!�C_� �"��B�W���}kF��� ª����>QC99���F$�5>�1o�L"����+]g�C,9�E�6n�a�����G���$k�r�>˵2Ft��c�7�[��j=ǟ��bӬC��J�������IM]E�o�����6��(�c���0��&(�|~��P�����ʜB����$��O�|N�Z����\A4�
���Y�?��61��ި�e\�T��O8����F���{���~9��`��o�Ou/���r�#�ENi*�pʟ0��)��D��p���_�Rvs�b�\�QW%���G���D�ס�J5��K:tC�|EX̏��X�l��@�HE��x�B�ՙ����(�Od��2u�K�������K���q�К�E����}L]>�n��anYՄ��*�OI���0~"d�`�
v���:З�����0N�q�Jt�T�9
P0GtK8�Ů�P:mV�7��_��|?����͡�K��i�<�[����gP�z*�`*�[O���6�k��4�sc���6����,�K]�w��Q��Ǚ�;@�y
���t��}� ��R����B��T�C��B���Ջ��a�{��y%ht�
8�����v��y�4�V�e��_�hq�+��Ey��[��F`��#C
L2���Z�ֵē*\�N6@��hQO��x��g�e���wW���k���篛�}����j:�<+g�'>��]�b�5�Sf���_���͞��YSY����{��U(�r�j�d�a�s,�o��k��Ć��y#F$��7�ҥEB�:�K��U������Hca�RH�c���02[��x�ߠ�h���C�t�\p�g��_ӛ.0��!M���+V_�=���������,�'���-�+y;I�n`�Saa��C�j(��:����7!��%|	�&�P��Wv�������mf����ByOw�� ^����EDnV;�R�m�tl����Xꌁ�� ���,�v?M���.F����lN�	'���F���]`��X+`P�wڴk�z��_����! ��/�Y��~�(8�s�߱qP��� ����C6�4h+I���,8�M�i�t��UXN8Zڴ7����$-�=Ӫ�<F����E�ݠ3~�'J�)6T�݋���悸T$��x�r�fȓ�<i;���Z��z;���^B/~X�y���Um����DVz	����y�	�-}�$�qi.i��޶!��!�39b3Ƹ�Tv��#8k�L^�5�Ԫ���zf���✗U.t�ɼ>��(b�B#K�H�_��+�\�+;�,�9�����|���_184k��}������rZ!,��?��`��z���,���<#���&A� �{7K��R.~e	i :Oi�O�k7���iE�/H� 2���6�:��K�Zz�O.���+ �5��sa�4�@�0�˽����'�B0@�'��GxzR�0C�2
�:�.ծU���`�Ы>9�>+/������T�"����]�	t�J��UL�+sd��������L�>Nw�f/D�=�&�:�Ji|W����7�L�Y��6�5{�-v�GI���	8�V�#���[�'�q�G �z���Oq?�\����x;яT�Bx������q�6��>���b����=O��m?����~z<��C '1nV\�{���Y+�8hu�%��ݑ/7�`S��e��~N�wc��{׫���z�ω)�TsjL�辬�d�ڜ<���5����;r�B�s�X�\AlB�mq���!a�K"�K�O OM�:�V�~��4��P�[Ke�maJ��Mq�#�.���|���
D����_Zu�|4/1��_��2����B
A��ֲOr�o�I��6B�ޠe]{��"��T�7�wRk�A3k�Ԛ��<�jfe�Y��^l���C8����\%#���o����Ĕ:���jή�c���~���?�˜Է+.�ݪ� �	*����}�O<���o���������n�9;wz��>!B�����a~G�?>���� wg����T��b���~�tH������^!0qd�v��l$s�sA����	�
b�Y�(�o�E��4Q�k��h�PW:�V�	9���<�C��d�'��wɁ���X9���-��>��pmY�qtÿ�x" ��uRa!W�r�U+ͯ�(�Ac�!fi���t��?aw5�����y�7\��Zu��� ����y3I�h>]4��)#�����I��K�\���26/���x��g�֓�91#�#b�\�8�3x���w�c*�g:��r5ZcRt'ezaw�ǧz�ǯ����_��(���)v	��3f4��U2��.7ρ���6#j� ̽�#�V�a~�0�{�7vUf���Ԩ�G���	>�-�.��g(��83�L��af�w�J���#�;R�Wd�n���)Pj$��@A�.�U'�W3����)���"yQs���4YR�����SP"��ؘx�  v�@>�2���LQi`�R���M�d[�OT�~VR��B�̴�;F�փ��e�����ee�7�Bb��jȄR=����@P�`$ə���kWT�,90���W�	�Rh�C�Z:���i ׋oe��фY��KwN�m�y2Ϝ��P�KFO��_�1�-ѱ/��g��ʿz��B�ۂh�ʖC�Gr��=�����ڌ�9����qݟ��4��7TN�� j�
���[�P�&0��e���#���]�b���WM�j���.��k��J1���;�z�3��+u���'Ҹ;u`rs�� ��@�*�V\����DR@��l��E�.gZ0Za��e��B>h�6-��&���x�{�w?6V;ᱹ{c�&��2�R>���Ѽ�S��������\ᣖ7�]V;ټ9� T�i�L�\o
�jQ����d�	�V�(ӪX�M�a�篩]}�K��)�.	�����ܵ�k��}�l�	�ݫR�C��;������|5��J�樅O��<�
B��%���4����,������A& ���m�~���RA��Y��t�~����2����f��cce�d�y��g,U��7]F����##�h��^���`�c�9{XLQ��Ǭ�>�"U��ó�e���:%��o�W���m�T%|��Gώ@�����J�ZA���{s��o+������1��6���"�p#B��^�!H����J��q[�D45z�Fs�ҥף�0����ܷ��,h����M�v-[w�?�6�����5��q�I>�:�7x6�JiO;�\��+���:�*E.�=U��t�����i��[y�*4 &e�M-x GD,��Z��y���wQ��>5u�ZP=QHUE�q	j k�]/�]�Xo��2eZmlm'¼��r[/+(�4�SS��{t!�	���䞍'x �[L���]8���{C���mN�S��>�#KUz`���1I�����}DT��;{���^h�redu �m��v���<*�]����TS�J��b]�.��Օ(J�T1��z��u�
�u���Tގ؃�����B�Q�C��N"���u{��1�v՘�[���<��j�5��fp�X �JN��o�r�t�:��#$љ}j,GR�@,A�sX��m*`d��|��'��U�)�a�.��q/����.���h+�xh�4#GR��`��.���=�W�cA	S�"��Ќ�e?F��tI���O0����4&��xq�<�#�)H�M�����L�����4l�Q�|{ܨ�g�М�Mn�E4�<ʙ>�-��k�}@��J��R1�\��|��0��;G�dX'R�Q�?{�-X�UN!��q͟2n�Aw��:P���Js��+���a��t�3��1�Y�B�ζX:8vWMdkI�o��c�ݟ8��cڍn���s"<������������;�-šuf�l�I��!�7&�.����D��� ��A��d��o�؛��\������bk�MN�ēZ����/�1�ş�k��bW��'�a��Dj����,j���3�7G�TC߼'��L�2��}^��c��d<�b�(���|׮s��w1�Ƅ�˸� �����1�H�g��+8u�<��5���p�K�2s���g�9{Ԏ����f2�ɧ���Z�V�R{���.<�w�7�i����"�$W��R�ɛҩ`2��H������[����cɝ�-�X�}����5i��ľ�}r��HD9�
�q�+�z�;g�(×�{�J��2~K�Ra�s���Q���Ќ�Ԕԍ���%�d!�{j�c�s�GM���mW:w�Cq�-/vx\�G�ŋ�	��V�� P�}:��z����b�J/:�}���z�?}������r�\��uk`��)�k�R�r��t.l��XoKK���ϻ���B�T�VZ����=H�,PC�q9&jq7����0+*.��������^�,յW5�a=c���h�{Lvy;�l��(��M�;�>��Y=FO�yn�k�9T�Jw�y-�OD��F�m��dJBygu�����%Rkgk�*���Q�� ���H�y#��NtV���+@O�r�\��p3eA!̉��r"�[L��|��t�;`m��9�����H��p���i�(wp�� ~a77�����nE!7ͧI����S��ͭ��vd�����yb�nk�~��x�؆b*���+�(��p��^�.|>{�����>f��*�X�fFP��TRH��U3FhB��G5b�&�Sl9Y(^ǫ@ E	�NҰ;cx�^+���C�R)E��5[��M��`�su�	$�A�`�W3����[:�Pb�(+��)�@^&����yy���\D��x�H���������@d��9 ���g=�2	���Z���L��Ґ ̜&�o�
�bl^�W�V/Go" ��޳�P��VW��}vf��:N�<��r ���n]��@m���?����u��n�l,2�^g���%]��͒���/rܭ؞�u�۬�?��&~:!hi��!�֕t����%b����X��s߶���KxW�d�rVy�[#��t��P����h6�K�{ې5�d��ᜡ[�lNNd �=��K2������-iӔݖb��v�DC�Y@Na;���in����ZU'K@=�)e\�De{�Ō��}�u�ꓶ,�xt)�n�l�~C�:���g}7��Y+O36��H����oLʧ��X�s$�|&hEd픖�^�g=d�bV�X[+����5mu.�ʃ(����-�SMC.0�5[͓�g9�g�O�u�$�!�gjO��c��Z�ą3�93z�HH?:�{PE��y7~��"�{���V(|�B����g�(�P�tc{k�v��c3�7�̙g'>�}.��EK{F �'B��; �M�F��{�x}�Zy�V1qN�X�g#��Cl�lw��>��(^F���s�>�<@o}lo�k�LA��v���%��>~�4D��2	S�kǋ�;��}�P��Tj��zV��9>} �ѭ����O��!��MA��a3��8Ey> f�(������[ݬ��^ �5A�C���Y
�Ǣf|4x\�V�5��1fG� �n��&�J�2�H&22�"�>�RS3Z@����b^�����_m��
���UlIA`�-N6B,^m��0f
�[��iqrL;�	�8�3g{����+�b	��P1��:���ٺ���ضn��y�w���:�z��A��_8�Li�����$p�V�� B��v��R:�xt7>�akʺ̡��@QZ����+y,�l���k��Wޅ�y�RՅ����LպBsGY�.Vx�z�$����%qZ�+&���¸�,�-�&#9�[�%�`���6(A(0_"���;ŕ�R-��S�D������\��Ga<S6q�:�\�(ɦ���>�9fTs�	RUz���]>&wT�|=���*��{|[/�qF�K1q�E�Y/�(���w�3W&5��c��#�H��DR�@�M��� �&��s�z(���(Ϝ�el��=��n�K��g�
�䛭���Ur:8�&'�%B�E<��AJ�ML�@�_��3d}����4�3�ۖ�Ux>a�<�h��K�B�-E�������]�4��g�cy���8P�ȹj(Ԙ�
��aK�zj�Ǫ^�*�w�.gF�du���-VyKm�lY0�[s�8����5���]u�E���ր!�$o�a"8�����0�h7���T�gJ;��D�)��ނ�Y� ��$�g~���Z��3&	����rP'2�<t��Gqu�t�ME:&���O�\���**���%E�������O�F��򾂾���ek�(1ISl"���'h1��=fiG�;us����C�q��1���t���f>_�����kB�h����?�!��(��t�.zV�؁���01�!d_`�J��w��[�K�Z�^D^�U�`QǨMq�[��P+�|�	��`�L�=9����Q�����۫�l���o��E,{`��U�K�?��M��\*��\0*"Nl��l듀g�Z��|b �'~���p�#�����8�:e�TJ���A�=��A#�������|�*���x�r����R-�?D������&͍����;|��)�q�챀/�]����_�����.��8%�\U��G��|���Hjhwh�[�=�e�T�Aci$9�╻;�P�Μ�ӏ�T���y^�!E�{F���{�����^�16�U�D�-'neܩ��m�p�xm�	��:�^]څ?��2xO�O�`�;;��t�s�]H7�m��D�o�K�C�g���?�a'�{3|m�:e]�qݢ)prk]�(�j���[M�3Z7�w)w�#l� �D>���g�;�N��3���<��P�^k�w
l+_��v�[C�%�l��"X�h��`w6U*�.�A�`�x�~��p�_�l���P%O��Z��gXHo�{�M1q$6�
��M�@8�A���ފFuj�Ψ�����Y��R?�Z�f��;Ց�LebV8�%B��T7���&c�ʤ��T��`Ǡ�cv�2}c���;��ڦl��ʙ[' E��;%��(�����,�8��1
�P8�@�~��u]��y��Pz풿�J#�5�^[� ?�?O{�J��#�D]���()~����_%�Y�������omt�q�z`:���y�?�,<0��v/R-�}�qG�v���sk�E��u#�ߦ)s��ӌҫG�����љ�Y��{���ac�P�-�Fy>E�'�~�]aћ��g���D�}�93�ߟ�M�`���2'K� ?*�P@Y��7��%�.��X��w<�"WR�^��
*|�����_�|����O4:&�u�xXQ6T����f���m�j��v��?�߰/�/���E��!V�ٜ�]q]�Lut8���Z��
�*(%{r��]�xo������^X�
�F�SUP ,$*�n[@��k���[�����qf��-�߸��H�@�����*RY�Ȯ����R�$o�沞Nt��}D
�@f�t���_�:ȼ 0R�_4�6{���~�RN��	�M$_���j��i����D]v�����x�~n�ќ��3cc0��q%�V/��Ұ�A%�M�Y�\v>�^��L��SN6��\�N�f�������6T2�����0���H`��϶�g�@'���B�A�`X�&,o�����3"�(E�y�p��2-x�mK~hF��O�h	6V*��u���`2 �?,[�LKa2�,�;�n��튻s���[$��lI�-�j�y����,�$����]A��(4f�m��'�ܿ�bf�]�w0����a�ut2���b6
n(ܥ��`��1�[����?3�T�ߒ�	)�M0d|�-�!��@>a.]0V������;�+�������/T#������K�t揬�$)����!�~�6�7#)V�p��L���E�՞�	��p�As�R<������甖��Z����P.��G쮈��(�V����5$��D����:�Iw�p�>��)��q��:*��ȧ5�^�S�U�j��Q�BB�5�ٻ�Ƕ$R	��e�\�����1$�����N�AWw��~pI���^o��}��)��ˀ��dˉc�\�t	?{�����R�PW�|u��Ǒ��_��K\E��!�>�6M��_�b6AJ9⍩W~��L�������_�v����Fa�TUz��;�Ϣ�F�&�>s��sf�Ԫ�[��g���Q�}
��91�~��{v��Si��n�v��;ڐ�����'�EY���^�{���,~5��D'�n/piLm{и7�wQ����X�]�ͷ$��WlC>���T!tE��D���1�w�,�s�,�҃��'�U�����6�+}Ӄx�xxq�t����eבo��]mn!_8���e�7[i���(7�؂�u�Y �
ż��ф��K��n��L�����}�/��7ra�_c�V���(�{d5�ݥzdd�0�&�'H����\c����WY�ƦImM�*k��O�Ѳ��e`�/ޫu�+(z=>K�����va� �ũ��@r~�3 0L��$Z��XM����Dl6u�4t�����#�id1{0�tձ�ZW��ϩo���'��m�H�D �=t./��-���#�Eo��ݿ�?�!��<�H�\�KT�'��Z�7��2�5����CU��:���JD�����'�s�0���2���b�t�u�ǐ�3m�38=���X��9XB��5#f	N]�ex�nˍǙ�[����T�y��4����w����@-( �r{�P�ꕃ!�rΥc�l���B���CȢA��~w�phT�B�y���u�q�7p
l)!t�M�*�S'c�JK1�E���*��]�;.���GT���P�١5Ȇ���&�Y���"�,!��ˏZ����D�AeU-�Z�������<�J�㱸:;�O�+ͱ��NE-��ϸ �*,2�<��m]

��緷
(hJ���������3�%�-?�6�ص�`Z�3{o�mh�c��~}�i�4�������NF�{agѮ�-|H�6���j�o�Xf �;�'��,K�|K�f�����n���~�[]|-����iM��y)��*z�z˨���(Ё���6f�F�B�|�Q��8Ϻ=��X�'�ɣ�Ձ]��B!���i�W߼?A�'#m��K&��?ڨ�J�IXق�Zx�@	ن��P�?�<�]4�M�e�=Y`S�5��:�q�)������E04Tk�j��7;��_<Lq^E�fRF������W��i��X9�S����>��eX�t�j��T�����v��a��L�U�(�ۊ�i	�T��1��*�����k��4�W��oܿ�݌��-n��?T*u=�l?�1C�J��oLJ�!�@J�ߕL:%	���@���_A�󵴎r�Q�e�pɸ�8����;1=�!>@`�60gnm1ĉ4q������ ݹ����� H	�t����kD�+$��L���$�QQDԮ7 lCA١`����Wa��+Uwe4"�_q����B�Q���8��i]E}����t���%$[	c�5!�b����eP'�;a����=0�G,���Z�dL&&݁(���Н)*�	�kI�ĺ��a���J�r��-9+n̥
�O�o��������tA�7����H8oޥ�tʪ�ڒ��<��d-�Wg�\L����,�๲�� mg�e����;��|;��r�!�_�0jo��5$bK��aO٤�kl^L����3�\]~�|����"|]�S�t��H�#:$�gE5>Oc���[���q��ɇ�Z���Vt�D;���3o:��=�+_[.�Ҥ|#M��JFI��Ա�~,e'0V-�Bz�j�+<�+ۗ�����*��6�^}�LҦ��F�\������6�p�!*�U����n�M����,(��(�>f��J-f�+�$��(�u]�@�Oa1B�9,�2�,T�";�V��d!m���'&�Ii�#�&[Vl9�Y����2Q3�*0�!i$z�7	u<[1�U�G�	��˴�����Q� �\�ٗ�<3b��Frɋ��	@[��!3܉\A�mHxiIO�?��8��캦շ���Ȅa(�|��&O�˄8J�V=��*m�,�G2�xC< 9`����� uVh>��J��rbu���-+�M�E�����e��(22p�&�X��7
E���ߐ'qz�.�����:q�S������IkU^���DQ�\<R>�RcF8%_p��6��&�d�p���?�܋al������7h�_9�+
=�)<=iT	����P�_�]�k�����=���?@'���Fz,�c��'�,or9>I>�`nW�N��ߌ�W�N9���-���{�4wd�:߰��ڋ��Uv��N�ӔU���RN�@�f�6^��*B$5�#	�)�I(�f��~e�ɛ��@��<�H��L�����Œ��\,SѦ��,�b1���}h��h��^�D�M�StB~�0P,�C����9�͌7��|X2Iy�cX��$��ClSN$�g_�_�Ɵ>���߅�e|�^yv�v��{l�����7\�8��
��Aⷶ|]��V�'��S^��uS�K%���kJY��� R���C3mGW��N����<�n�s���K���ji��6�;(
�LT�w&�����tԮ��b&y��f�=�F-9�un_��G����\%�GE�FZ ˟4k/U��r'}6���M��vR���j��ZzJIm���m�b�;����	����7�R�_I.`�����6Ž�ShZ�r��3���T���4��o=���Q�d�`���(���=H���v6*i��e(��ss'[2YH�Nx��xU�+��Չ�9#H�y��������?�?���E�Q_Th�*׌���.���q��M�Ӝ/W�������r���ҥwa��ʏ��̽���w&让Ǖ��JG��5I*Ҽ.�N���ߍ���R{74�ֹ��̘�'�eP	���pV`���fI���u{�8qun�&L,�䬱����7_sF�+�HA�����2kȿ�"N
$�g���EE_V�@�K�'8E�cg�#�S�'�O��1m�_]�8L�d�	.�L��M`��i�!��Lf��0��&"y�^~+�t\�)ڨ2ܦ9)���P��� �s��dvr���D�}����#	I��{H��M6ƁJHr��ͪ�{���h:��OԕY�������<C�W�^ݚ
{.n�+������ep�t��.������_nC<R�E�oMޥ5����'�D1Y3�I^&/Vd�y%��v�,�(��sp�U~��n��-��C��w�W�[AԽ������z�XZp�3:Y���ʉ�T���)���b�|���d���O��8��J
��hn�����w�GRʅ _���7�[u�_o�j�����%�	-����R԰O˿�a9�̮ �%^��f��ˡ8~w4�~����z�q�O�a��z��ދK�Q�/aRY�
�t�����v,$�cMw��1��մ�C�i�{_�9 �
�p���/޽@?���F���%�Vڳ�N�6 ���.u�(�ni�<�N��n�C	������ex�)��Սo$�JD��8�AG�j�;�`@�=%ە�XJɖ0h��huhn)���?���C���?Sd��CZ����H�W��]]?	r]� �^�����4	�Mr�\jV�J�i��>v�U{ٻ�I�zcO�D	��ӄ�$���.�oj�J�{����<<�s�����MAw1I]&-���zan��?��G������#2T<�y��G�B)b����tb��fz�0!������eE��<n���>�XB_ Va��Si*��o3vH]��
����I�0�
�a��.(u�G^u�<A'��뵩�gs����t��"\�8t�=͖�� w4�0�.d�Y��*5F���k?IС�%M��V} ��=?�C��(�so\�&��@�+lPߥ�?X/2��w��"�/��U?��k�1m;�L�(��U�U����!C��
�sqp��.�d�̂Qm⊛F����	��nXt�=? #W9�� i���C�p?_x< Ő-��a�.x�t/��4�;2t�1���*��JS[�\/��iH�!P	Q+�o�$��q��ɼ��+h}����ޜvZǑv��g��+X��A���2��,&�#����8��x�֝�<�~A�_���B��v+u\E��&IDLg�T������w���A��S��0n�{zZڍ�b��/V,����	���L���Fp�ZZw3=*���<	��T�>��lyb���ѝ?���`�ܽ:�B�>�f����5��8;2�UΛ��%\��)��F����m�M���φ�M��_	u���QI��P��[1�,��V�2��w����AK4/�k�%�z��_��a��o�Y�<���:0"o0�0N��r����m�r�ѹ�1���LT�`�� 4���/���v&��|�
x�jɳ"���v�*�ݷ��- H:ńHԹT:"�Jd��_��Z����s]����4z�ׅe����N|Ȯ ��R���γ��AB@���}c�M��x^0�_�g����U8�����^����̯��(s��u�t(�h���V���dag��b��z߫����s����Ǔ�7����⩸h}��X�^q�?[*���јŚ��ǿ��lr�k��hkq>��9X�d<�~������9#�t��x�/�L�}��EF�� �-�̒��ŉ��'�Ņ��Q����DX*��׋a��p���dCzO�2�-?��q�mP��ƾ��N^�t2S:���mn���醆ؐE&�Wi�2xr�(�_M	�D����\�2+�T�r�D2O!����l䆫��W�s�4�SU�^�YY��E�qg�$�F�$��Ќ�.��15<qءp0�ZMx��`s{g%g_�q�MϽ"'A�>�?�����ˆ;���SQ������H����,&���,WIk>)�`E5n�C���9���!U������,�yDA(/�(&��=�n~�{�ʧ�>�'Z�%V=����!��MB�y�Ex�Rפ0
�iU�T���� ϖ��_�q�W�TX<Co�ΕT�l�C�td<=�����y��TxY&\��X�?=�>�0���
�
:�{f
S��d�xVL�|��.[t5S�Imn�+"���1O�%v+_-�E!�?"��+�CJ�Vg�,�d�ѾC������d���^wK1)3,4�V�G��<�Q��]�Z�O�"X�=]C��걘��U�����HJ�>Nߘ�"�ۮ|lu	�� ���cɆ����L<�j�g�Qi�b8��Q��'�^�l�yQ�򩛟>9�)�� cW�VɅ�7O!��2�tŋX�F!<D14��N�1�k�5��+n:5��Pk��׿�4���7�9�D���H2��� ��
"E��	7=�	�x�pᶩ)hk����ȕZ���B}���[a0�ͽ��*�pir�X��֓�sEM����n�nҙUI�q�ɉ�v^~x�Sǡ���>��.�^����z|�Q��f.�R�';��ܧ/�E������,Jy��T��\s}յ�u���ԩ�@+�a�bg����,d��Ӑ���i�:���E�$nAV�J�q<��<�F�r�	rq�k!��?��;�(<FY��[v���$7Q��GG��H�#�haI�s�5z�F:}��K���~��u�ݬn�� �m�[f��Y �̶�L~`0H˨6�+�����"��/�.`�0M�H�-B���f|�v�6YT�h"��2��ڽV`K��u?A�Z� �F 4�
K��i��o&K�8��%r3��\x�h,~-ܭL���T��O`c�/1���2ZI�����=��N6��;����&s(o �<����7� ��}����)QC+����!����l[֛DAБ+�c�1�G _@&��j7lpB� dC\k��3y(�����/���]�0�a}���.����ל�zB��w��-��{Ǉݶ-t�}�g�~��t'���Ʃ��Ŝ�R)5����9�ᇹ<$~�<ɍ�\�g���@��5�n=�X���U�@z3!���i����[p[#�%?<m�~�O�e�70��s�z��rpe}�h�>'}���N��(�Y�M�*̌ 3ͮ�Q�*ƽ���8�^�U�37��
�T&�:&��}Z������p���t���Z�Β_��fā
�w�V,�8��D�k�D������-lp3[;q����jF��lhl��A�=nHR�rٍY�¡y�r�6��Z�Z�M�f'1�g����c�t6�K5x�3,�=/�&Mo/d��C�(>?%Mr�a����y���.����|yb�jk������!=���,LO�7H�ŉ��v-��.��Np��)��H�V�� �&Q��:O��굀���o�\�'���QrZx��_�k��D3J�v*:s��;������J�3C�#�~��T�9�3�i��i��q�0*����Pr��xOF���;[*��pA�H�z��~%o�䀁͡3 ������`m�����&򪲆mvz6��(�߄Œ-f���c������bS�ɨ��̉�qf���q	u�Ru�ǟ3=��am�MyޘÙD�#�tJ3QE{c��r�Ʉ��L��:�[�ȟLs��'-�	_4O�=l�Z�PG�u���{	D�������ж��<)T�F�Q��/t,Gi.�^ijuj��3`r��z�7�W&�҆ڻ���S�$ţ������W-{�Ѳ��T�!���'�,��A��@��H�i��\���5���
�u]Ką��.�o�r��Sw��v�J��ؼC��$��W��o�����:�[,�ȫ����?.��Ts׸3p�̿�K�r̅�9$����k�
�x�z�נz�����\]�m��y3��v�� �M�	��"��:��w�/�Ќae�ߙ�Bw�,�J=lб�gXZ��)nS�o���s0��=o�9�G��Ƃ��w�n6�����J��jdz��]�&ܡlߦL��L�+�\�����^kc� B�;9iq,��p��t0n`LxT��O�2]��²��;~&��-~D��%�� Ƶ#0��$tTϖ(�ϙv�/mk����W���	N�D�S[A����4o����}�ı(���"��d���չ�y�]�G���=����H�7�ޙՂ1�@�\��lq�;�;�6ȗ
QK5@@�}���	�{؄�P��t��/P%�/A-�wߝ�"%��_��z�^t�F���p4#{�$|��������}�D@�Yz�R�=_M��r��t��QGЄ���|�s5W���g�c����o�D����r��O4�J(ߒe�E^��p �>��F>����b�[���3e�0YdE>��|4��ZȑG��9e�qM���Q����eEb�i�p"�&�{$_O������Wg�{�H�sR�6}4i���T^/��6�c�aȽt ���<�킁?Aa�
�\�;nj�ّ*>�����e.��fK���iP��?A�Z�� Eڕ�CO�/�M�ӣWo��9 �������������O���!#��~=�o�H��d�D���z48�k;�i����tB%Ĳ>���0�#�Ce��Ņ��a�Ls��sG/�[o&�xG楢؎6pl��(B��Qb���Y+�:�w&����e��E}}�erO�<L4I���e���'|Y�Ǿ��BtJ�t0�^�lf���A
xa��Cx�aL��i/f^j�0bMne��"�j�_%����u\"<9&�B9����X���e�T�BLٟ����4A����sU`i(��!4��m
O���_�<�g;���cO˺�	W*��uL�K�C˨��	����S�n�<n�[�+� �?7��[�Y�� �VO`6��A嶎�Q]�S_�P�8W�ԟ�"��~��2��7ٻ�7����]\'"��ɦ�sA(�̭4΍���^U���������,u<��z��' ���X����:��tS�9+����򃌶CD�����
5��G&.��4�mV�yf ����3����	�[��ns�QB�;܍��=�a`�C�S�Ф�`7N�������C�Y^�'�W�j�X�}/��qEo�(���
�J`�6�)�
��pԨ�����Z�yǅ��P9� C����7d��Y�+�U���U���3zЪɫ
e��ߴi���[(�����ko�0p�Jʷ�h�����?�j<Ө���0��)��%��{��ih|4���x�&��NQLD�z��WHq����P��U�˪����8;���9�AM�M�֨?������h4L؅���H��h�	K�ks�b��8h/�4���\����Jecտ�3]�^��!�sq!p��}���W]��>����J�[��Y~mɎ�^zTEW�-,/0k��j&���[N��OiO �Պ���d��jNC4ȡ���sd�s���+��sԴU~�-���h;`[��Q��	P�9����&*����,���Ʉɷ1v}�Sʶ˒��^5��B~[�wl{f�fH����C�AѺ����s��e}�p�!q��RE�,<�HP'�7�VYF-�@�=-[U[����!v��^����Cq6����3g�V4��@,P����hW\�m�ͮ�o��q��f'NSK}<\/���"H�,@�mbӻ������{u�R'�7����A(���'����n9w��]+ŖL�۾��c����n5iTe�8�:jHu���V���J\*ͶT��b�4��`.|��X_oמ��-��t@ ���d��]�if���ۢ�ޜ4� -M�6T�r��U�8	�R���|�![��[�@�S��+�Z������kIy+A�-!�;�S�m9���,��g��⦛v��N�Oy�&���~���=��p4�vs���Q�N�ZINP�F�+_�Nr|���V??Ǟ��{��(O����D�s��^���� ��kae��3�[80<�%��^m�9����gL�j��W!�O4r�+O�L1�6� nt(��=ۄ����X�Lg��T%x�Q�\d}5��|��n�I�^��Ϳ߾|�W�}�ӈ�-Vt^��)b��I�4�
��O��B�3�=X�b�|0<��0�@�-[��2���?�ay���}�B��i���z{���+۱�l��oQ��P5�`��I���L3?�5f���q(Y.��7�t)I�-R��~��_���2L��e��
��'>�~V�Wަ ���4�𓷔y��!_�z_��%l�<d��El~��^J/�,*�rb��-���yy|�����f�yM�W�>{�+0����c�����3��_3|A:���؋���/�\�@�~7f[�P����my�=���d�e�'Ӑs2%�c4�5�=A�3��cə6c�!n��".Cf��`��yA�ֳ���B1
h�A���/�.�& |�1gNRe��4z�_A��o�#y�{�R�� <o�Bvj�xjBa�[���iM-�
	>���$s��5�hϰi��պO�;�A�6�ٍ8כlui�a5��[NE���d�oV�P��7�![/�^��a"��A�"[#e�,\*d����.����Sq��㰥�a��J�H�%^.�P(V�|��u>Lg��j�Zװ����
�e,I�|3Y��h�d��1�g�px����\���=�����ػ���Wi���ˀs�2��T)�.3���=�ery�7�2\b?iD?��,�6)5��������L�|���آ[�	t��er�j���J��U	�8�X>��Ԫ��B}��_��ْKT��u�zh��S�H"�Lˎ��{%��#��5'qe��-�LP�K���_���9�2�gJx)[8@5��B���O�
�r�ْ���~�r�0O�M�f�)�;���"Kլ��x?��("�<uLm�����on�L�Q�͋�ٺ��x�������J�7ʆj֐#�]W�}���Y��M7�f\ܖ����%����^f?��\�tz6��Hj�V�o�RL���@c���i�[=��фF��d9o�}2�ե%��O:�q��jr/7�3�"�Ǽ�0�7Q{��7�k����`�����,l؏�?�$H��$�����UR�3&�&�*V
y�c�0�o����B�wa.5{w�}�#3�w6M�����Q�N�qS�� �!��r&y¤��ͮߋk�#4C�)�#��mac��H��̻��OÜE�!٥kG�G.����-pq�=����}�'���|0G���M��:>��t��ތ�/T�M��h
���Y! � ���� ��|~�PA�7���]���6��=��˔|�G��������PL�t���Y�jm�z&w������^��K�$}f�=����0+흗��!�J�N�h��qH$��J&�'�1��̣Z�>�x���o��A#�$Җ�"N�|���ozIQ<t����D��L�Rќ���v:�9�oZ]��u�l��'�r�f\�Ùa�Lwܽ�6�х�z�|�;�H�x�l�a��pF����1�~�~��B"�!%{�Gs����p!,���=�Ktxr.F�k���%L2�Q)ۇ�ˈ=D�I�ڣ0@N���ܘzN'�a��!;��M?�ax��������/l�)���j���^w�~�P3���w$@�I��p!	��
v.��z\OP��#���u{��e��I���fJs?�<�O]50��J�^���D:v�W��P�|`�8iX��s��܋����V��Cz�z�X�	|�!qzR��f���"T8i*#���3��-ă�7N�������p7M@���(EYX�@�r�f�Br.��d������Ծ�1�����7C�!TM	hꗈ�����v��n%N�j�����X;6�R��pm�3$�hcUi��E�o5�7����Jj���r�[�6�z-0似h�_X٭�<ɸ�3�����'@A@3y������@�M�剷�#M������zUOe4�D��*f�8߼kF�3�;n�&9���S9Iɂ��\����v!�9�U�d� Z��hcq�.-�]�_؋[���gER.�%v����o�Pqg\HdlR؝��fPo�)XU#�on����_�c�`���×<���Nt�4ż�u�� X�Y��:۱����$j���0u�^ٹ�3�M����1T��7��u��ّ���WL�Nbi�e���>
��;l������y�%��_���F��/^�6Gh�2گK�������G{��8z�3&���s����R�j�����:b��>��,Xn=�!#�;]�(�����t:p��+>^i׷ �[6��e��1�a)p<<��v�&�_� �\�ߓ���3�r�
���я[F@�r,�k��	���"���3�;�vFwu��Ѵ�L�*p�[0���nïe/zs:b�6��������ȝj:������I�� �.D���3ž<��80�t�x��'��\u��#��e.�MQ�}��4Uԛ�*���h��,�uWYc:Jd�쪋�㍥����藖��I�(e�B�%��E����:*��W�+�^�4�V��L�
>~�@����ƶ(l^1�⦨Y�>',{�~�?�er_��0� Ip)��h��야���Օ+OV�{�Յ#�Pg
`�Su��3�ΤPM�.0�#� /x�tp�噼��ؼT4|��f��})	��K�Ƶ���4�[M~��#+�K�1�Q,�t���r�qhrT@��7�+0�]^x��mfP�ɲj�����_�d����L�޺� 9+��L�lU�ʹ��O�`Z��{�	�L�F��Sd��'0o^|ǎZaf[HG 3 ��B���S���������I~�F��r�\A���{��q̠!��"����g0��l2�h�]����t�$N�,U��"º�q�j�X�a�S��\ȸH�ĳ�hXɘ٨�^��-žC��ᣔ,�M(�������s�{��NDD�@h	ǚ��۟��|k�s&�,=���l���a$]�qRޑ(ɼ�|�4l�!�`i���Qs��!t]i&�E���shA�����`�8#�^�p���� HÑ%�8h��^ �>3 dnLD���&8��i�u#h�e¶IJ�W&��-��6y}:�o��y�]�mQvj]�$k=�Y+L�p:�%A]GPn���0����J�F���b�T�<�r1��z9q�?V!�T׎�?�(�eC��������9�*�;�m��h�m-�5� �it2�������R=������̩-7��6�)�N>�,��������CJ���/o]�b)�W���wD
 >�37_X��i?+V֑���!.E6=A�U��`L@r%g?etpu�\�ODͷ���t�O�c�yul�v��ܗ�5BU�Mg��<�Pж����Q{:�t� C��.��CY���J�q�l��F</Fdٝk� kR�]�łe\�����U��I��-��� ��eLO"��x�T��9z�L��N�t�{� ���Ǘ�Zs9E�d ����̧}#���Q��cB�H5��2_ }ĕ�4�@�.��6v����O���&��Zk�5��x_����шv�
U��E"��s��[�~Ӣ�7���`��>n�+ ��x��vn%���:��a
m��x��s��B���)EB��ҋ��͛X�}�S'�)��jr[���$�W�V썴��b�*0��ށ���˷��^R�/"����1��#�T,9)I�kxQ��bPB +���ܦuh���Gi��<���|��JJ`*i��Ke �\���*��e��L��s�Q�ѮZ���/�Q�g����7W��3k�(;��~9�L��C�e+�w�.J�fv�7ι���P��}v$��������&z�t;��0foZ��w�2�e���0��z-[76Gp��Lr�5	ra� ���9�/�� �"{����Յ����޶3��&5;%��x):^'���j [}V��KC��y-��~g,xڲ�����	Ţ��
<wC�ի���w�*jU�@ϴO?D�*�G�;�E�N�{`/�U�r�P�}�鰨�cn�f ��b$�+�N����ܸ�W�o|�W������}�/���A栔�<��[B���1�]���w7�89��
L�zָڂ�.�D��ZXn+=!4=�)�wo.2ӇWT[AT�T�V��א�/���R;m�'/b�k�XixD��aAK���.VF��`�������l���~s�4�k��*�d�c�JȌ�3�aX��E�ږ����?���������׫�.x� �ܧ��
��Љ�5�E�x*n{:� ��2F�)!Վ��5hƿT�%XiBRz�4���
��Ҭs���f�hx2�W�HTbv����dG0D�VH�`q�FUĢ#�<��4&
�������l����kF��~~� 7��E�� �!���g�̘�5<��*���0�1�IH��O�p}g	���pq �$F�R���Ps;n��3�>�"�ԳZȅZ�Sh�X~c���p��ލ��)��DW"����W��|7��b!GF�������%����U��"��39C��8��K=�"��CN��S��#"Q
x�C�0�ޙ���*fRs�Z��R%���r�����<%OS��lvɣ���'���K�xհ ��PE��P��2}|{���̝g����������R}?$�K<L�� 0������p�E��Z�)by?�j�)����[�ɧ$ �3�`�5�j��+��M�];TA��_FI�[7P1��8��c�y,oN�c$�Ӧ'��j�mj�'�tJ�-��C'c�5���+�q���O�)��r,�|I�|�F6��?ׂ�zz�J��L�
\H_�,�$׭��\e<c/��uپ{_X�>�,�zGݢ��Hg�j�ʠU�4&�IV�� �D�~� al�x78[�廴z�@ت+Mۃ��0��v0�G��#�Lt�N3p�1~d�C���h!sI?�&)��ȑ��Js��c�����&�C���k[����D/	6l(@6���0z��w�����U��ڿ���BŽ�?����m�u��[�jP��%,?x�g�܌��93�T'��)�[�9���bv�#j9�����A�`�lߴDd���<9��.$=�L������m���8�%��i�A��\0��G�;�,
?q�����~�mA�Ķ�.�J�R^ex{��I�:�;��p/�+x4g����&;�C��u�oW4t����T�|���g7��i&�.T��)�>&c�4��\����\�u-Kfǂ����k)��}N>���.`t�޳�A��d��;I5(���&�W?�q�S��j�����/ޞ��S@�VYa�4�kY��U����Š�(������z%k���1�
�*	f7Y��	D�!�Ơ�KR}����Ac
_
����<���c����1�T$8>"{���F���:�K�X�$�o�_7�0��a�m�:'���Q'zv��`����A�S#X�����d\VO#�~�Ti[~E/b7^i��X4�29j�#���x刅bI��@0B�B���8�g`�������OJ�ϸ��v�Fi�8{U;*+ge��4��X�G�7�Ă;Ё�yh�$����%"~FCFxb/>�V'6�o��W��u-�*�����x��U�ǥӔ�҉zUU3BZ�jD�(�r�-���a�atf��^T����ìl�K[<c�d�%�+բ�q*1�͛��{�G"�v3E�9\Q(��F����h�х3p>��31A��]�X2�sr�h'c�1�>����I�e�q�����L]����O���S�ZU�	eA��0��r�C�	�=,H�il3��W���rpJ�����5�9O�;3��}ދ�E}����2���?K��$C�:҆�rB��؟�w2Ll}X�� �Zb�8tύ��Xb���WŤ�*Q�aS���鎍Y���� ?؋�6 �?X�����,�㬬���3r�h���G�A��qeQ�����������(�B��Z�I��N�w9|�g���6�	����$f�����<#o�v����o'"��[��3�c ��M�k$?&9���[�ڸ?O�����Ѫ����~=K��x�A���;쟷���*�2]��r$��Ҷdp��|�S��B3�	�АI�3�A<{s���n�o:�.y!gU!\��[��������MN��3���?��h@�L���8oO$��"n4��o_P�����yI3��� ��OZX[Z�G��ڨ�4�𠜝�{�?�)��G#�L�W�w��YVa�\�$����NVb�n�kjK���+�6�u)��A�|]���tU��Q�g��@��U#θ^�D�H���e�@����"[^��g ���.a����?y�-8����w�఺M����,.��������V�N.t1���lN|�v�1�����#⌏�n�@Vȓ�r�|[	��T�;9�`���\�bc��~��?j�9I�_� ������c����Q���*�y�J�~C"b��.�F�xW�;�O�x���=�_foe��
��.խ�v�5��n�`Ib���Q�9�lK��WC�Dlo���1��n���`��^P��2��L?K�}u��?��qN���'��5piV�����!�4T#~?�\ږ���Y���d�C����G�X̢%Ի�bv���z���DA�5��'kE�H���5�.�3�=��^�����
�d��8�O�\ۚ��Ϳ@z�ۻ�Yl+L�M�n�����"�6\��M`�H����^�3Q�ֈ��^M&�*'�*p�����	�������@��S�'w�=PI����D�A1D���qL��uWqC���Ɣ^#�[�?�����}m�3K�G�.J��%���S�I7-ŵ� �����u��.��� �|����pm�IE��Ir�-�o�	��U�����p�T�Ga7��@Y�d$�:VDL����wE��m�3(ѐ��&%�� �7����ĞW�v�HX` ��$ �6�$ .�)���|�Su �f$��5s5� �54�� �>U#"��dv��r@'������+�����,���9��PbB�G�G�G��Vw�{�������_%��wq�'u�1�"<�-]�9�	��/,@��Sk�v�S��D�y��'zlkpJ��6u��$���u�b�
3��hC=H����-�0���z�\�\��J��{��=q��Z��XNod�gQ��k
<!���د}[\�'Y�Y�j��wtTޘy>ġ�������/fR�0�`1�S/���n{DQz�h��Θ	nk��c�,X-��:�)���8����gEo��bR_����M�\9�H4�$-��c�(��e5� \vBզT���&T�!Gd���z5p#�ŕ1}]ק>e� }Fk�MN07k���Y�o��ڒ�XʝcT�"�jX��s��&�T��� �R��c�v��J��?��w��?׈��I��e��LMS"꓌p~�D��Ă��qL} n��O�u�U��PCl�������p�ɦ���4���F̜T���Tݫ��t�����4��n�'x�ƂW�)B��h�p��8q��0J@��D\' �!0�`�KV�At���*�߬fo5_nUXk�j]��?�ְ4��qC�]L�9Qo�{��/=����b�b�z_�}��W�^�g�L]�y3a��^�8�Xo�9ޏ��jמ3B�Ҿ�^K��q�}XŎ�خ�j��Y���p+���(7��쑦��l�B��,���������J��>��'�c`�fT/�;�\SV-�Yw���F�6#�^肞?k=�����0^�J�%������jdA�D�2	�yf��bX	�
�d�$Ժ%�cbH�OxҶ!�VA?#�66��>Ax��.(,Ȕ�-{W�Y�4R::��/��5�W�()�~~��F�p ���(x�D���*f�s*��k 7;���Wzª�2_�-���#�?�C:��{L0�n ���͙U�G�D�:�N�T���<P6I�
ƅ�K�� ɻG�2�szSHǗ�Z�����2^8���v�����ޅBͳNE��E��R\�}�r'�(ZPS����h�ɩD|���^&V�u��Q;���ݤj}L��̨�p�^(���+����V�0�w�r;��)Q��)���9�Z��"N�K��q�S����1}��xT��~��O��^�*��#/$��C�R8l��#�)+R�i�0��û��t����9Tn���[.�o���"��1��@���X�e���5ܫ���Վ{��ܹ�,��V(��~t<�r-`��͉7����&z�N�\���k�`�v�>kZA�.���ߟ�C��`T����\��D/dB�l���=��?b��Ҧ$��z�:�t`!j
�<t�_x�>6����2�O �}�%E��0�W0l�����j��O�>\& ���ѵ��k��;��%Ͻ��U�[�ێ����@�����\K�.��U���N�wR�;կB�.4!��F.��-�錫��
8�/<�)�ߴC�k�.�i�)X��a>���V�g>B� ��lT�B����PԮ��ʇ�,�����X����s/c��6��
�a�t�lJ�fW�"�+>��l Z�՛pK��Z��GTk�h)����ӊL��(n
�z��Z�����N�3��W�JP8_�ς*��j���!:�F�d���[P�z�s�L���x؛��oї�Y$�uX��]�$�K�{��AXTI�7�/ʧ諏tDb)�(�W�)���`�y�"rO3�z�;���s][Bs�],�\E�2��JM��=?��,Q)�8���u�]��I[�tS�G�!\��/ݸ��Ӹ*�NU�MV#�v�j��e�`L�
�z�7̬�X���=B�U� ��3yn�Je>7I�g���[Fw��};��=Ze	#ӯh}�E]5�;�O����,&׀�ݯC�?�	���}oy�U�7O�N!��pP�
��aq;�+3%0�gcjb8o M�kt�#u�p�=)���6m��r��������S��vP�x[&��x�*�Y3��xC��6}?��=@"[e^����n��aKl͚�H�I@���9����=S�Y���*��.ZK,�D��rBj�7�!�j�V'4OH�ID��9љ�l'�	
�:�͐Jk���H٩��^���,��ߚ��U3�΅�e�F�a5�������t�&C����@����n�	 O�eC�G�U
7���.?#��}��+D�X