��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���� n;�7�Ov��@a"��3S�(����=�[�\l�|�$W��5'f�vWtX���>#ߏ�|ǔ��k�q|m��1}Ps��S�{ܢ^XMK!�_�����ľ�У��J\{9К�h��]/-��]�37{W'�1yΤ���נּ=�m.'c�Z��a6�+'�WX����qg�Ȑ8��Paȏ�8;��Uk��x/ȶd��gNc�M�]bE����p�B���rďe�Q
M��r=@�����C�3�U��i���֙3�n�A�Y�]`9���2�E%P�~��_����U'�7P�&���A�D�u����Z��b�%#K�Yă&���.3TA)��;�����UӞ��c��f>�5��\�	�0~���uN.�+
}ۿ����NX�f�q�(׷�k}�Ϯ�o2�Yډ������)�MO:�w�&Ph~+|ě�Z̺�\鬕~A�x�D�:�+)�h�[u9��+�g4<��jW�(�9���+`�;*�����݃~�+Q�����O�2HO�儁53[�e��B�$�=��UC�{� ��fu�3�Y�Ԛ��1fB�k`�8����u,�~��^��_�Yt��' �E[��������6��=�2�~���U<�D5~4f��SY��7��f�h��²ʋ�:���L@�ȗ��c�4�*�����Bv�a��%���'%�(3��ZO[<��!<��Y&����8��I���cSkȼ�!YBۦU�i�U��qu�����uҬ�eKy��k	e-�*�	h#�WZ�1��S����}����
b��3^�a��{.��{D�ӯg�HgG�g,@t\w�`g+g��W���s����m�����a�Ks��De	�|����;�,i���	"sD:����İc�����-��6J��J@�;X�'/�\X��iQ��:��PN����=��2�M]�Aw�yp���>��OS=4DZ�d�T_|9^�_��=��.kCV�?��!A�~��(�4�e�u#��|٣������Q�P���3o}�9��.K���Kh@aZiS(p�G~�z�`�#4�q�ak"*o��LЕ���w`0�{�)S�����[�%'b���衝(���R5����r�U�_�8\!=�烠��(%3	��٥J���P�˘7�lq����}R?�M���V<�G���#"���~ٌ��֙���G���Q�|������icqh���pd��}��d�Ao	lRg�4`�E����8�uxn�Y^�\�0	zNp{[[�%h9U<����2�����<|���6`�����I@q��˯��3��"#O�Wz��y�5Vb~� ���f /X�մ�l|�Rr������Q��x�Z�C�[�E�)���	��\h�(X�D��Lq����nǣs�Ŵ�Mh��%�Y_.�i�+֥�P*�|T��L���(7eE�=�T_�.��U8H��`D�8��]=�7�W3S��RW��#]u;f��.�uN�R��k�`P�n$�K|3.F	\Z\���ʰ�&�WNGQ�I�))n�aY����s͠%ظ2d�z���<��:�Q�����s�ͩ�������9�E:I�B�|
�+�R W��V0��NU
-\S��죴#n���ך�������;��EC!	��ߩj/Fbʂ"z��Ǧ�N��E�̴Y��(f�~�+hvJ�����"	�E��>�G�IL�nT]p�6��sMLւZ(n% �O���u��jД���o'�gy 	@4x�Zo�շ'Ix��d
V�v�a�ݔ[�{�E}��f���+�Vw���d��C�����U�c���I�S�f%Nd����ap aV�ѓ5�%twa߸�n�7�@s79�x.u4w������ݣ���(V��QW�ޜAp?����E��"�.e	v��p��Dב���ƕ�
��ec�X�����6A2ˉ���.�d�+Nv��+�o��[W��*y)�]�-�l�,�es�UF�k'"!1�� j���"�y%SB������ا�
�'rˡc��G�����x�tQ���S<�Ïr���;��r���N_h�B~��Ӑ����/��f�G��NX���ٖZ��7����IC�t��d�.�b�؆�#��گL}Cs�9β�$X��}���9�~udUcpy�,r��tĕ�P�9���˒TB=�����=7�8�3���[�q���l�'�AŴRPǂ��{��+�N	���.xq֭�̅w�6/�Dj�'��@If�5�l���w���U��i�!D�a��3�#�n6'�f���n�J;b�̲%�=��q%������*?>�%ހ����&fB����M�@8���T�E��|��d�Ӊ� ~�Yك�l��د�=�bӶ�(� P�d���M��CgF��uS��Dy���䞔6���\��l#�6X�i�ǿU�.dsQ���*�6|��EC��s�t}܋�����)/���m3���Q�b�����X߲��m'
J8�W����� ��Q�#q�Ú��<�/�9�1=�ʒN��,�����!�|��!4˥�*3����OG�ۍf�U�~oZ��;�:�����?�͎�9'v�ѵ�S^�6�dL���V�W��2W��4������K;��X�Mv>a��7#�ޮ���1����L��L-AcU����ű-�޳�F�Z6�t�E����~v+!!o�Go���D+6v��F�����	:�g�Ӽ�O�������(bU�_��.�����2�^�����D�gs��\2n�ꖄ�w�S�9�����T�L�����T��-7]������A~]]1ҏ�Q|�4���r�g`����!,xg�4�k�?��{
�!L�{P�̓6�[�����e4<ocˁ�`^Ђ��=V��L�=T�6Z)�����.�q��I\]��ى`0��H��M�Juh9PLn'7:����}=JcC��`�,�yMxS�����5e����h�Y�F�(��S�{��b	�z� �`��8���ߜdQ�eS�@�f����= ��?��W����,�����on��.{�"���Ȕ7�*�)���symB0K����[��m,T`�1�.�H���գ��ew}�r0��weZ�j�<�.H��ޭ �`j~�ٓO����$ЉcH�U�WB4'�m��!3N��ѡu�g�zF��W�BBd��QA���?l��!���9�`��<�����{<��Su�G�e�L��=���]���C'#��2H� ��?Q+��_	BB_ܢwG5�Ԣ��I
��{��������[%oU�4	��2���/�3�V1�)�3䑻�-^�ۚ�D�d(A��cj�ւ=!v�y#N{�L>���<��OJ����9�5����Q˹B��M�)�Q�R����G��b�y�2�WܒZ������n��`˴���8~�V�6s����x�X&�ύ<ڌ��G��hױ��u� �ᖾ"�L��sz�����7�ŏ�ݘ��ui�g�����<Pz���
Gm��Z��qt����������[nŭ
�V7�g��ӏ6�����9k����������nC�1N��2�=�Ӓ>��q�/��Ie�Q_�����7�,~1҃Q�x�R#��d�
���@�U�o%����#����BrƑ뻎F�"�N)0	�$M�o/�J��4���cM0M�!e
UM1U�ˡԹ;�9h1>=�j�5��i�x�� 0�(GR�T�)�������F(�]\���s3�Ia����ϻ�()c!��IHp�P����>)U����A��H٫�F�P0q|�G������1'i[�g��7�]$6{	�͐fa�Mxr֌�s�������@�F��U*
|ypM�̪��AH��{��X`.�Z<|Bлu��e �d��e�.�!��?&J++���Ld��g�{�_���q#`\�{���C�Z���TL��x�%�ۙ���E?%�/�l�M?��M��	�M�L;���bm�����&���:ot�cMj�'˨������y�q�����D�ӎ��hD��e.��kS�JY��������|�+�k0)&��|��m֓��A�c��v-F����W��m[�&�7B�!�GG��@i��<���L-~0�10/\��v_&[��*b