-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
biieDqlLXOD767RiOOrjmw1B/twea3Y18D6rC2HEGZhh4nuy4uuSwun5zt+LvnxwtFxTBtbV+qiT
fQTLmAGCPoCfJSy1RNufZmxs0bZKFJqeWreZSTYJv/6NUa7AFA5QWgdg45MG/Jm4VvIemSs8T7de
g8+AN0xjujXjX2Y4DuoMqIXzSR2vcI8TwK65zqf9hH6NeuF77Rsp/yXUytJbHNO5ZkeRuv4cme5z
rk3cZmEm8HXG/MvEz1FtkJVIMIvEUhGFOdccfQOHU3SFlt8U8Rdk4RTLqbwqbtJerBqtm8CBBYrw
U2w3rXg5XAjIg1ySXcMOyjYd5/3c1VX7emtA0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
oos/+yjYJiLUuQ2UKNUepF94jRIqDTkT7ItnxhQGVcEdjhYt22QDDbjUeNmOFuQp3zjPBKp2kAJk
fzBKMgdqApgnMgkt5CKO7yI55U6uwxHUlj5lNRr1M/DTDcAkey0fOe0YvcX7fgALBM4cdLYgb3XT
GlfD9tkAMGRUv5j+tZ4UoQL9WE913RwGs/sSYkphqxaRXjd2I8LilEVeCyzyGXSVlBCRpqnq5/7Q
L646oSZJ/SPWeFDbPFJ3XWlNj5KBMm5RNzVVn/2ib2/VQD/KxzxroSX5lK9te2HFQzJXfRSwYGib
Z6DkZTDQZCno7/afqifwNFMi0H4JwVDYILYceHdwxXqU1whNihbavvQyI6eYb/2noDdJBzV1KNzW
AOC+MuPGO+sBl5s8am3bVbpCEqUHzDLOgeslocvZfcYmvHbOWvOOTZY40gDxVhjoTTKvQ0ftZ/I3
j2KD8IT+Rfh1lRjO5m54++Df319Rdesce+yhUhxyUHhRihSzh8o3CjIDlVVY15obAjd9UBFJjuUW
rdsqfucjZbOgGCK1PmrxgO/qSvAE5H2Oxf8bcqT+Dppe9lwajQWN369xW855ex7COA8Vd77HX7k2
0r4gO6yFgkvA6UgxwkAumVaCCCOF1Ea4nz7IE+PHfbOg0BlWKdbzHhG4FA7SwnTRKmbM47x4Epy6
WsiRz78AEOx4gA9RDinXQ3uOSvHZmrh+6V3Ho7xX4+/sdUHQ/1lhgS+3ZM3zpaf9/ZUt9AYFQRN5
MGOKHDNLNXDoevfbCOklQNYyqOWkDjHTnKIZdKv6dlvE8k+CCCI5JkPoreYx7Jcf18PeOr7QYPy+
YJ+X53cryCftaXOYub1zkK789PRjA+WwF8SYqJGX8sNMKy7FK5vXhChdkJk8K7mwjSZ7v+7OgbX+
eVB1puY14hHua6tsRp50APGXUOTP0aVnnl8bRZn0YM5iqR60RxO+hZ1QEIujrY7x8+UROFqf707L
l8wqd2dYdf2U+xY1stzGTRebBZNXuo1kQgwgfYD3MZy5J5cJOZo9nxMdXTyoI1FYtks4Ayw+sBvO
lRixRRpnF7qc+NtOO7GTYPVgZ6tkHje1JKKjftWfrH5V15N8LWa1QC4Ki0heEta1QApXHSYsW9E1
Kv3KcXV4gir463AfxfGHbzq62OlZO0pZwFfzbmHZO+V+jRV96OcoRAGzr1l3v0BlPuD1VpUDcEaR
1uCJqrEVLK/ZU0VVzKOeLwRFASov6uUPG5ufIwAKQzyct/I+GqUQRBtpNpTqq0y4fJdMryB4L27I
t2A03GcnFtA7txsCaIIMVTJ1eDa4T96GpHww+Hh1MHW8GMEfUq0LJ/UhVMCnmCFKmTKkS1kSZ47r
2pzSlPsS7QE4c1w/Q/PDfpgwfhfF/uEV6GRaeoc/j8id2D7VRznf4Qv92o9hCxP4vUGjV5YUorBl
yQQrDyX1i2Bs8+H7RCz8L2GnqrcvuRg5Xh7nLOrQs9Iffb6grRP87Hrfo8jZCtv/nAZO3ghKTZcF
FYTn1gWHzG5qOju51w4Y8TfPBgycOUYc6s1sQkLjkNo0NRfZidslnBb3lDY6qLdo7rvf5YoTdqDP
+77Mt32ivJunyet9kT7KEvmKDaT7/gu7FTlqhaG00Ik3Z0hUNHuulKCjAuBJf8FQRvrmHyhs8Gs5
PVgdDIOIrCnSs5b8zRH3kqydBFCBTSDMovDC7poyoL0B9IDd63zMHP+4f+zEzEYA2ECLrrPGAqD3
auStAGOumLS3Ejxbr1rAzDoWljCG0CzoQhMdS5Hie2JwqHcfAYo5xKjf3ii59t1T7bbhp7fErv8b
FHCSNjgV67YXoFU8KHwt5emN5tZ54PsqN0XoRPO4dTvVOAL/NVAxsFeCl2Z9DpwIFITXTcnqhewf
zj5ewlgXseW/5tmsqy3/eeZJGJ83i60+bIvit87zk7+rAu+x7Nfq5SOXEKofdjRn5OcrVME6p3R8
iIoGV6/vMuVJFYyjSdBbsSrmtn7vOoDeHz4KTGOM3RdPaZr07TI0xjnik+AofiiGb5qPcdfEjU3o
Jg1KGIzAlg//EeEICKNC2xrWJU7RQpfodokHw4yjZODsmgrQf+Da5QKu5U6yrf7rtS9D6SFj6SCe
99eX49if50lXPNwELcj3bNcHZf3RW0IcINGDjlO5XYSYHSCUIH3HjTWB9s36vHCGwvtt/V3aPIMm
bNpRKNk3i+kMDmP5rkmeUuEvAOxv+oP4jN1HcvCoi9hse5m80AnXeEsSvtwg33ypOX5A4IcDYuHO
X27c3sJ3RrdJjrMZTX2bO4o9p1On35qzTS4p+hQOwA/2M+53bKASWOOUJpXccekoTvmAtipomWjr
TIAzjPFcjLadVFcl3UgYF5nTCT+78o8FOxg5AOBdNnENPS13UhyA9mOVmFlX1lZ/H7MIXjrD4flH
kXQ+2NNgy+crouNwVLsxwdi8n4Mvgawc6hnNGHz4mwBH6IVhqa3RwHDGuP7R4sS2J/Wn9fZvcfGI
MC2Kt5WxT94YuxWKa6ak77JE8zCdjRpqTAPibIulQ0bo6Avg7l0dz3n1bH2QpJ9Wsjy26k5LZ2Fu
LU3kcAoGhaTXRG1KUXqoEgHcbFpGmP4zmBSCN8QQ7NeC03DfxLptHj9SzxBGI3CDOexZy4A1/308
tc50sVUS/dd3qAsGvVzcgtvVoE+GvX2mU/4f1aUy9bvIzqN97PzS60LcIpSaAQgI7PhfNVqbvPfY
DEgdI9nxHcyosWcWVHxSFaOg7AVUnMIj5gPKRa+EitjogNFKP59yrNnZGe77wJz0liDedplp4Z+T
vPKcKyLpT6hD09xcNSzeoiB/t8XhvCemGAiO/CCQktf5v/r39xgEsNzJ4NHR0SsHOo73M6BMqvpi
qjxCv9iGCeGwYSrAXC0OkRFSONYD/gTU8nreWdtUsS+p8r7K2QRrCFC9Y8y/KxJ/xM/3Gi/TNVkf
bvLTM7XqcmAtSuLG99p84XVh0OcY97ACdWNuNGwKhnBTPVSSYEc+OHT4Mvp0HlaXkbw0poaLkiqm
rwqSpPIvPPREJa31vcQHO4Yp4Ckc74dc05Saj0Q94mdBwd8dXUFPNxLpgPa9wRPXhgvpkUuUee8y
XNU0vi4vN9o6V4eKVZj6VByP3RgCFaRNdeKv5Hn+PIVllSW33tJd5dlWJK9Mb99/hqFsd98Hilnc
4YMS7B6Xj5RppsTeZg3t0xoxH2FiAcICWMHB29SISv7dME5lbU99b2gEwPJ1vYCYSoOv8+PCshVM
wSQxxeExL4yZIQhVbmq2KnYo89PjboiUEpVsPQfKqG5Z7JOlh3Bj1sTVDHzKIZkHIxuPHFck1USS
uXKnvMXWgKU7QNkpb8n1xiNxIiTT2xE84Y4W6ZKznqZKp5jYOCW1RHGZpY7804f92r5WWDVNisjU
slV7eM5PaD5tvMilJMnXRc4c8X9/o5+Qbq6/tFxM9NQi4fwjMyFfIGcqMfuKhbpsFKwSLn2ETfKw
SuR3KCgP3mEoAclnZOSi9n43UHeh2clr2DOYgulj+ovIUkpy6ibcs6HfkwNErN9rx86X3QEBF379
KckwnsOFB8kxqlNk2t+cfjswBcydIhAsr9hlIthbZfPWK8sNLaxW/HBJhKKZa1cc2aB+akOgfU/J
ntQ83Y3yd6jxW+BClVJGq14d6Y0urgao3dH4UtCD/uVl8nmLH7rScFOEnfm70PAKopO+ORa+AUqc
REaaUeJQ1oJd1ISS9JxkScvlLxogwHmbR2y890Ipw1WWQA89C3jANXatBO/GwDoJhsYMX51AtXy9
+otSXq9GIdMpB1lUOh2t3FjltZ4hTXdCeeCKcprMiBaVSo7wZRmxSriCZUs/42gvRl3rSr+kLQmO
pM2OC9iR/nj8cV64KcSCP5LocRZ0uOBEd0OTbrvTT06+QjaCdEjQ4m3z2yIlJoZi83HTg9nwOK95
QRg+//pC/0ifKd+h9jn9VjcCLIdo4nyrj4BJIAg6/88fiz26bhUifmNlc04MGivWW+ZspZKDgMqE
mN+5OFXWnbf1GismHDactWnSDtxC6rLoP0ycVktVU2w950fcyI0v70Y46SnZ4Y7X82M8bIA3ORcc
5eyi8PRa4ry/n5Qi1O5Wh2buVlPPcDw1nOyZ0i8p5vXfz+PYiyKIRAV2UiWuFtcED4uiEXY0QE41
A7H6Y3YRkzjESTVKsHQ08DhlRhahmkt9ETUFu7CG9FYEB9XI1U+2e4NUwyPITUFyBt5CVXidYczC
88TLdX/p59+l9d2IShKd2sud4X7KwbLGyWGh/LTWXbu6E/6pUkYN1nDl9ZuR1v7W/xMFR2sE6hlr
aC4kBA2PE0LpkCT6poYGuGQ1afIljVGSoFHo6HcpfCnPyYzlsnu/Fttz5Xf1MHlstvJH4VS2KJRq
Ibw/hCJNcUVVu+BM02Vt4byv3eT1etPP/6YBbEUAosdcQzBmEd9xszhwt7tG4kIrBfcgdsTGo4Jh
k0YGkrHKFuvGhokVQsxWroEtaqhFw+nq0VlgQRm6Yn4JaqZFd6l8et/W5SK5V3AT7qygxLXJ4vuh
P1NYO335zd9DECbkRsRt1Wjupa8wc0Nv9t9SXgr10HvuNhZ8gYJy7EkjsOXmK5EW4LXfIA67+y21
DaLjTwJA7GfEj0g9KiutdpQGZYs9wkaa43jCRJPkD+GNwfUnRt7v+WiUmBbvt7rK5+WYHZ96zie3
+6+GuOVE4JtqYmz7imApwXaWCZSpz2sjKUe6znCCDsfOcvTZDl1H+pXYQ3CQWO7duaxWoPXrjN2r
IOL5u7fxqdc9cniGJHOr0klm0h5IY/bbVUAYSctREiGafSWoQWqg1SW2ExDt0XOA7TS67xxmk3SL
1aeAV0Y/C2QuQy8+hn/U6S2+TbGTJZQjTzPn5Zhq5eVG3YobdAc+s50MI7rkWpJfnIdPmYngQxf5
FpyAKtbLVjbUjHNvtmUozWCHjLzOUjeBNPOiTyYY+85U2u2GhaEf7PGwMy7JwdqZTtU4unWZWe8R
VuziRs/K5/M5Aqa1MC2SlfWoNJj9JkDqtCM+610W0yBnYqn4q21kfp2Ucg6qIzkgN13n8LOj+mGu
2c+54g73wLQc21XgyMohC+0zXkQ69DaxfCBOyPzB09OLRrgI1iMtdUwnoEUYlJKEyV9SpRzDIWqg
uwtN6+FemNs9/k3li0TUqPz0GJUtPd2EPWd9NgOrtOLLswawtR8e4VABE6X3fNtuiLkg1yK8AjR1
ahGyHK0sZcRLzSVpSoKuJtz7GQSANgTSeXKlNOlmflnplYLvBTYg3NjhdaVW9XHiuEfCMKJlm+uI
Ab2AP3f/MiLOxHXJYIhKlx3woNCtuXMjO5qCCXUKGjpmL+QWCba5fRazXsSkYd70XA6zUhhnjKof
xInbt1SPzlkhGmFdEq8uq7yVo3U1qy3BIXZCEfrbaplJSf6wQSTddCpxAQwPjyaTTg6TZ8UScAMF
6Z1Z1qF74TeILeAWGQ0qvlxPixzshrXWrLlpx7+6UVf90b/lbonT+d4g0V7uuaxHAK7cbtzWhnTG
2MXrHBUzU/U8JLE908D1cWRL91L5LsSobdDtrlMk1JpWCecSBL2xvoqPxIUIQjdwtgMqPZaAJ5Hk
Ktsxu38WNw6TMc+xjPX7dBG5gDZ0wtKyDnPT5LpjmMhBenRhpGBubnGTTVSPQDYzPJLLbbeLjWKg
Y02i3e+SYTBYBFVqVwLI0hnlKT2RZ3i/TZqrByKXrbi6HAuvZUnPk3YB9xAQBhITpLQabCxyGm8a
k7lxPJVLDX2l3YvQ/7e6uwD9c6DL4dDbHt+s346aHijCrBOkCbJshWSDKscO87hyrOrlW0bW5lUw
VXYELu2QhFHTSyWrxq1f7Sy3sgRsVhoh+JEhFzQHzoJIfDiw2EhwiiyZs+ZivEBk7n/f95NXfVcr
J3H1LDPbxV9t5RuVlIVo2lI2pVXMWwOihWdBDjqzUFDgG8uwJBZTUdr6lBzsM5GYOa4uD2Ad2ISX
1LtExntATRHQlP/xuOdlscZbRMTGQU8Pw+x3sX8dxnj62JPnj1cY9a0RmDDrGBIh5NxYwuS2d6H2
pJ1cp9BzcGiSSnXI5tFIKwhKEMm9sihH6qVa96alEpFJbibaJPgZ1xACQb2+Co4LXzoHI12PMVP/
6NaUQ7FvZKMfWRbRs625g874VKsNonB6+NYC5t0/Ttb+wPkG+Mo5WKGLKUIfVmXtXMRHEUw/50K0
mdJ1AOaOyYQGzckGp/+5+trVyyUk4HiEZRJOSEB7owinYVywbezETXj4wo24iPejIf101keaWjU8
uOJO0T6jIVL52B9o0TgVexaypnDF/HmUqx6l3jPhyqZo1RtWwfQqdyABddPrRfK/lMuNDwLWq8NW
pZous0vrwHxGbXLKsM9G0GNTSUcCVsoNu0143TdqsobcGWCYspemY5nKiLvzlgZC3bET9BkmBhHH
XDXuzCnZqcNzGs61PgaGbgNjwrTJoJUOHS1lAW1hCVN2rb4xRlX/wnl46uPshqugvpH2rYTDnwXS
5TLWqAsQ1yhw794DliCSJChT8VZaZRkG1AfaDVrkTwNVQYJKsFbfmJVq0PmEBJmLIImxD6Mvy7xq
AAgOaaIJ0eUu2rNv4wr6bh1lAAm66xE16/PbPeeVqm3d3gOZtPN2a25PXpwKWklOh6Nceq4bTGMd
elBvTndS25QRB9rYax5nVAZXV0xzH7QWjhfVbX/cVLEh5NW5LvUZEmORnRgyuDKIdmtMg1J42w5m
G/PMQaVfomBdK1f42AttSCV8pCpVH1rWOV0/VOsGMFK3PJPghusXC6Ln2AKPSyP263WVV/snbwWp
IHTFxFofep8WOyZDtoEtJV/3gaQhz/3xtORjutPyFzUEeerJltOXHgwmbbyU4f/9X+aRrqQiu44b
uOGaNMD7DnZ/KutifYcfJQXs3Dm7RzshFtYnU+XahweVh7C0Eez/vmxFz9cX9GDTd6s2i8fCZkAe
oHdVh9G+sRRIGv+dBfUmnHYirnWbcrXDyyyJz4WAuvj/j1L/uu95efnLEmeBaPqT1CjaNjXDo9+F
vHajxfCRQOyj3v05p/M2rgtg61TLYScqfH+ECwCKU9nqoK6V+BNr1e7n6HOhCUFCcHNCTOIV7d/w
zuhRSLctdXaeTUzurmVeGBtA1SSdAD0tudyjp2H4AGvuyiFepTKq+X/jg8kqicIr+WMQs/wZUNsx
zZccucO4U+9nzHOQjLvHjtW+19j5mmtC8YkB/o7Y3Erm0LE21bzyafuFe+8xbMsP7dfsZL2xJwR1
BHWHvC9vH1m5urMEdWuv7/C792tbUTdzoEL1E8XAzx4njxFb00za1rmaBYoNYhZR8KBUWav2XFjd
WcAD1XTd1tkphlllt+lGIjgCJhaquvBR0ukx2Kgvd77Blx+KG1wWV62pTp3+3HQ+lf7qsLIwGWtX
f3PKZkA8MTOY3BGML0RAnhAyrlRAtqipNlxLwSpj/JhqyoivNiOrmD9l8vTkWYkMYWfDj8PszwWg
Dlhn0TZF3aV1aYDKBMmGEkU0eddWdT5PyThy9YqR7fWi66dhBHgvSsoqK+zDLux2nKC7fJThfnuJ
fQjVCEGrgm0TSeJ3wxwWD7fqdNH4pdyvrSvpiLdbWimgZsh+hW+dWD1swEvJ2ZJu8B1kB3iY06Xv
810LsThdm9oEnZVYbkJGwJlCq25oW5mYqVuJonMPN7/A+vovShzPBgtR/vB0ITHm99p9GKZUwNJk
R7DE/X5P5Alh+EDPeH/AVb3ZrneQlv+U7jk4cUypTs1z/wXOHUMbIm0KXkGPgaj3A5j2bG6sAmoH
vEraPfZkg2Rv3pRyFQZPx7PIuNqE+XHCR9J18prR7fpL5g/YkEixagSpP6VwzkZCOy21r9cQFBIs
AIxcGtxIrhCxveBuvKSAnWLfLvgZFA+2ZQMGLOR0b54uC8JvN+eOOc3HWoWdMYeIezga6IgviGcl
JiHiB3e9XYodui1bsGvwFIDBD5lz+C8MGCbwSeebSQZc0ncwkr52tJjHgQl6IYnq+RUELorbmOWh
VU8ughKjUc/y0Am/t3uvXaLZo85syaaZ0x6lMetWDftDlIkqZvo+8o2OL9iKIV6XsREG+fwUTxcB
9isvUrFxxOaB5Qau9ZlfAXVy+SM//N8Z7pDCjX2fwEKnPmFfdZxPYiNJL6rAZwRPrt/zyILYrq01
zC7I+LbfgXCMOIxDAEem2Opb8ViZrzQBOLZT3T/FN1r/oFOxjgi9DflY2a2OOTXPWlrsra6uxUfG
lL66k+nK3UGrXqW6MMDcfgMrPRPRaxAaocttfo8/6MTqQrDenH5MVj2X7U0KaeDf0LlXZJo9k/sG
rHnCFD6IizqQsbajUQVuPW+DkiTH9xArj2NxIVX1hwgJ5jAmm0mrz+TgiLpPyIbFuArhbL1FNj+p
RmtgRa4yFhQQ9rM16q/nWO8Zh9pFiSBM55rFuvn/betG6f92Hx1hyQA/jfB5IauR7oIDjv2j/ox0
ycUHvP9xqwMUsuqH/j+pDBrHSO/so8t+w3x/XIgYo2XCRIux/AdY8fEtv+f5nwHnHetIpKo2FKkQ
sbLb+8UFHtbSmMIXyHE6hdgBEP+kWG6wU53kMM70ZBSG4vrrsBk3VKGIT5FqXsMnyfJkBn8tibqL
y17dCj5WEbhNk505j6HBhlqn8ng2cb3Qbh42OgyHhsHxQe7yCHVeKozJ2yFVlxxD74g8G9fnOdW+
zIs0d3C8aRicgX3sFjfjcvwIQmrYepoulqo6DmZRNWNDUpFR/gZG12D/6Pj1/WRiyTfJ6pS/i4v+
wkrs/12aOdI/nNVKVVyqTg0wyPe26Iy+dV3fa+TLtG47LB5DlRvfdsaioVe1XUQ4ifKDUd/pmhL0
rFF/wyCKOMbbTCAiQoZa1DO0YJQR7tN1UYGv/tiZ1VrY00bcKihhh1cutGM1qQwyDQ04+sc49mGa
fv8y3YmXJ/g+J2i2sEXcmtg/nBfWs1ULg1zMy6XFzsAO/IuS0/AYWMZL1mG+3jEk9wXOiYDzwz/P
ciBYVXTYemLGYYF1BFjwGjmnJaUaishrOJ9irv1d1Bd8Jx8lNlj6B/LoxW/R0/rI7akPpvWU5Als
uqBEeiWm5rVB+YgpeIBsnz82sWlb4VQJINNRQFK/pJ99B8+qQoFo/lkpk+zYMk3vDwAK5B32tCr7
URXEEsdDLiD7MEeqRaLGPaZ5/EPb0XnOfw/NI3qZwEuU5WbLqEm4tdpeu2DVJghqnbJnimCnw8As
G/h8d5jFIWeJnT5GGWJYtX0Lz/JQ1gtd3K6Z+LVcMk2QHLXhmyCMavO0EtjUaK/FdoQWnKMjrToK
drJzwbW/SUaLvf1CYr9fxKAa+6062MD9xlLvHMyvd/HGnZsnhMgZl7vkv67MGzPmizqCiaPi63VB
Bhg7aR2Bnklonp38WTGwlxIgNHi+01a3VwqrWyRn55p6++JqoXH50Lo5L2K+k+1imrumwM+g8+G1
tupgKRV1sPOj3vyNYe82divS5S9m1kmcRclB9wcy5HOVfd7wzjv58dRUrRXoycP9IBwTPh7aUJcK
4E3T+m0/C8tODDFrYCXcOLZmgFfk3HifBsXEkkj8LZQgp1cTo80B0Bc6vegfaLtE5C1+kVsqBfae
jxfF0be9yZy8Sr4+OdQ9yMYUboRerbxp67unrW0uNId7sZmUgk3sDPtJ/vIjJkUtWSnJZJ8ALiB3
JzPimE5enQG8X1pQwOeYsUIlM72wgz5p9SA1R86O1lVUYO8YEt3JACyca3+MAjPfqXYlEpgnX07O
cM6UlWrPq1Xw4FN8lfoEQ9qJ6fIAdOq6Vt8TOd0P+I1aULkDuTdczU9Ik9gInnCD6yL9wjCOei6M
hqO2kqPmRxjFEDXaDyx+AWUWugQLSauyEA829ZzRiuocs+QYwhaAW0OolWtfb36d87+jSmVISuqd
GOMJm6A7LLz73ZDuwqdBiyEThZ/en1KkQFxIwJFhOI9gIgdjoQYhmhYhLvJK23tHTtbOmabYVyjq
y9SnBpcD3c6iLjdxo2NwLXqXAcdVUia1CVZ8VHDOC+tAviLDoc6qRB6G3OvR4gU8NcdYFku+HKd1
OwqvgbM+SXPQec2CxtLfZkl3Qw3lab1tab1qWOazfuvwcKJT+sV4bd3HzNIw7fh1hvDl0g7+5v1T
G/SK+kgFeaWzd9pjmPoxd6HCR+WFBmBhNlg=
`protect end_protected
