��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	l�-d�S%�B�O�-��H��W.:U�\��e��@�#ysJ;PF��8�b�HTd/�C=7NZ�a���r��B�l	��`�DW�4��
J�8�ak;󕣈����yk�t�2-��aP43"�[�A�\X��
����_���^��֦����K���&�v�dZA?e��8�{��:��gA����N\*�:83+�
O�������J�����*�.w�q��F#Q}on� �@��c�^ļX������Ċ;�aX)�#H,o�(7S�;�L�.t$%(勅m�:�qf]KD�Gn���\?Cχ3�#U}�e@��CU�����]/jY�����m�Q�͂}�&�LP5�HT��I�Ţ}
A��u�g۽݀��s#��G�p8�}{���H���U��?Ԁ)���C;������nO���b��>��Zʨ�{�d��^�M�\�	���>1p��cHAl�ÄV�1�!y@�+��z�`ݦ��R6�#��xd��#�\M��.^��z�$���ß6n�� ��|��`Ct��'f/�u�ش�H#���9f�e��͍��F���<e�W��.��z$�T�Ɇ|F���߹����ڭ5vs�$)4l��%z�BF��\�!PW�! ��+~����"�IMhS���i����B��4��ಃ �=-�#�AuN*��a�������Zk����+���:4��o�s׾8�	�Ln�B�
�v�nC�U���ZU�ѧ��v�����c.gLx�&w6a�ph������B��[���נD����L���-79�/�x�� �HU��v-buË�ڲ�Ƚy��"V�������WXzj;��TYC�������(��MF�:4�eF &�
��NV�Pi���������I�>�q�6��03�bF (і+Cr�$>����7G� ���t �6O�%�mu*���p�ژ���m�'˺Z;E�?r�65ҷ	(��o�j��h�HA}K�D�PB2X������Zs���&. M���j���DM4T�OF3r�����<�[��8a3���5�m3��
����<t�� �#`د���a؝�#=��%�����0��h6�ϱ��}AT���ވH��R�NM�r8�ks�f���0kOA��_�i	��I!9�bwQ#������!hJ�����ʑ���ˮ�kx *�q�����9�;�!��4�r�K�WN���暲
(�*�ڱ��M�Co���u�����06��p�"�nS,����L��.�;�3�+~�  Q3�0�+��c5��A"������ӥU�bػ+��K�"П�(ѩ��J��fG�$|:�����`K���Y}����piB*�Ǻ�6�U�
E�3�vb�Q�R�#^�s��·'�Cv�	��:w�u�m�b����c��_c���~T��o��/)t(?�c�F�^���2_����������~p򃍅N:m���/�+#/�2�xh]D*�(���}p����
-`8�]��m�T��܈MA�/�����dC�����h�8�I�g�a�q<���`3�~������fݸ�lj���>�*H���� '���ؼ����fJp�۵LNE �Á���D�>��ej 2�x`׹jbW+�ӱ�mg
[�9f�m.ʒ�|���|*ڻ'=���^ʁî�?8<+r�n����z��5�`{\�]�oI��=A-���lmmݗ1��7[��vG�h���_�]p\kxM��S#�X'�Y���,l��U����y�q]���;?$�[e)�Hp����O�������qr?33�E7oӥ����t�ȋS,z��������ZÊ��GB�W����V�L�d掏��L�8,~��.�'�)Q �W=���Aw����RI*Q<��ᾝj�U7�׷֊�2N�<�rg��fc����f�%E%����ǥ�	��S��	�)S�����*�����$���â��H�`4_��t��_�`���dͧ<�#}����>���J���/5��Y�*F�72�p��7#�,I�8*JZ�=\d��M].����3DC] ���&C�>����F��l��k�ט���J��aUY��1�{����P='��C�Q��l��(�4V~.�RqLUᨀ���!K�-��ҙ��zy3��b�0�>�ҥ9� ��#�p��/cL���>�պ�D�Ȇ���#��+����Q�J�%�H���YhZ�D��gD�{��Ӫ}w�k[J�\�=�����5��435X)60~��ʒ��t3)��gE|nk��~�N��`Q�`է�ز��D�;L�]���is3�r���	��1�ʡ�nk��׭�y�l��t��s'��L�2#����!�t+b/���&����\^��&�r�s\��G�ۭ��Z[>���\�je�ѹ��Z �%{V������D������U~o �t;�S���������-o段W$��ҩ�N�d�S��R���sJCLqV!���Bf��>Z�锌�;椼��:���M������6$`'�V���
#��G[�@ᐟN��c�b�Ji��]��%�iH��~�~3ǊN���+��M�6��Z�6�/%I�69P�}؀3Ua�x��|�N�;�U{�c�Y����Vge� >�����B<D��v���>��B	��B�n�8��1\��!�h���E{H�'�z](�)_L8��&.����L T%g���F�@�.���y�A�2�U���1�!}�;Gώ���})�9.�Z��L�^D�E���) ����q�8���2��Mw�L����
RC\@�����'5�mt�Hjw#��8/)��ͅ���h�PL#.G POקXj�u�l-2��J�(Ϡ��飼��"Z����v�+�)pn��z�d(��:a�ou5�$�c�����Q�e酞C5�� �KAq�T/�w>�������^�e��3ú� Zi��2��wu͢����G�
��D��O�N�O��X�%#�G!1j�ޘ	7�����2�W���:х�|"H�����Q�K2��=�+Ip�$m�6z7���:�V?��R���OL��V�;�5Z��61lJ��Qb\>S�"����"6�5�����k?n�'6>'�
��8E4յa�N\Q�Ԅ`M���*}=:����~#�U}�;�s��@�:8FM�o��&�^;�>���uj��z�
�]��T;�omZ�m侊7}r3�*����AR���流Z~ų�Rr#N8��r h�/[,�ء �Y"�Ř��m���}�5/�$0��X�P�#�f&2v�Vm���4�	hu
���47������Ⱥ>/є}���1C�d��m��89�T�Fci�4ne�������k�B��'��T��z�`��H�R�� k�2s8ƥm�*	�6|�ZLqM��:�d�$|��,tj�Ƹ98���u�X�Ya�n`�4Jc���G����Ajn�r��HzK�U��å���1֞:]{�.n��$��θη�vĨ
!��bD�&�`Vg!�k��� �^u<5թݥ��:�\a����l#F�62-�Rc�^H�N� .t�E�w�l��"�E>dٶ['���r�X�$�q��3^�A<�4o�u���Ca�y�f K���bmn�������c`����Ɍ�M�u���(t�ϸ"�\��튧��`�<ZJpX�g��~"�\���u��֑�;�p��qE	&����.���
ҸnCŉ`@�H�H)�)/%�����'�Fk��pˮ=hZʐm��Y�4���!��q�R���Y�¬!n�7�e�#vn=>*z7�rI���	�o�.��G{*P�m7cf7��`�����w�l�2���x����.9T�����O�Wx��iZrQ������C1�R&������o��MV�%�l�55�3y[�xo��C�.���
���d��%�Fvl�+
��d!�ۼ5�2����Ѿ=�ۿ��,�92�j��D���0��T��e�,o�3�x	�4۲=iϷ�1R���f����e{�n���q<���8��s�8H)�<������-���KJ2���L<���_�-�.�8��؏���O�c��W$9�b��~e��������Zg^dE���~3Sp`j�1�@��� ��D�}��O7��V��qqvH��2?e:-�W�r�Ձؠ�1�+U;
So>"$��,h)E����`��ql30ʵop��2tz��"DY|�e5zԻ�-r���t�MtU���چ�&>���-~\��I\���t�����d��my{��9b�;3�?�E�h�7���yV�����0�U�Y��n�i���g>M6����kJ�~��ߒJy�8����;�'|�'�5az]{��"]U��x�O��dY����8�jl��[�+r�1b,�VYY�?���%��D���)�9
�v��9Y�z:��+�`(^��&�!��3�2�{��]�ِ���\�.\b�n1���U��5(6�ʄ��x��u<?��k��E�c,�_V��Z7��>N�M��B��*���"@��<�$�Ua\��St���G���ch�&��M�J�@��*�cr���6�{X���P���ڛ�aǐ��T�PRe��G�������G�cr1?8U��c���:*�A9�*ݪ;�JY/5s�y��w[��fݽܶPL��a���%@���v�W2��.�[���W��3a�>�'F6��:vf?d*�h�@��ŠO�\�q��(�#x8��霛�X�<�/5���jE=�5�����<B�����,����l<�5��zک�Ⱈ�X1���ɲ��-b>�/(�@Y���" +��b��:C7_����km$;+�r�Hbf�|��r����?�!\|����%�M���[o�������4���TaJhyH/4��3댁c@�~�q�G���tH),a*�?��I��}�(�A�KN�����Hn�\s�BM�B��ԦyG1�8���<	S� ms��>�����D=��|rf����)?�&��	��nR����S�3�+�Bο^@װX�:�������ؠ��&&�����%��ф���fc�QG6j4c���!?����m����dn�F
���An���O+�C��HԵ��aq9��ԕ��jG����Qiӭ�b�����Э��!/ť�~2��^�z\�5���X}Q~z�k�!���+�w�"?~����5I�7�Sdd�M?�'��x��	�!� ѮN�u��IԦ�i\���si�}И}�������s$}E]�z�Z� ?>��]
��jA5�	f0����B�^�5v��'�@��C`m�фOtf�V�ڦdqw}���U1��dWm��
��{�]���`-�K����f�O�̧�g�2��V��LO��o���7��S�=zhy�D�2�*���}��h�;���t󁛩��J�Äo|��:v��)�J�vho�Z�8,�8��⡟i`)9V-�WBW��~�T�^��G�K�(20�Cv��>�΀���71�]ƌN��/�L"j�b�j$�O暤��2H'd�m���eZ�/�]`���ʚg=��m��ɹS�I_y��{Ȥ�p�Sm�5M���~D�ϰ�泶5���੦PAD[�#'�o���tf��� Y_3&�nD�ܢn��|4��Q
�O~�9Mtk�2%�!l	52We��\�����TÐ&�k�s��`ԃ0mLRuU&���>΅R��y�O�OI��?!a�b�1�baL�����a�Zx2	�c�AҜ�ą��%u���NnO���*�X�J�����[��E���S�I�y�zu2P�=�ۭv��+��S��$]d��d�~�O� �]A��u�4���a�V�3�^��g�M�'
x�"#gj7p�y]e��Zm�R� 	WK���]��3\]��1F(Y�M�x:B�d����G�^l���O�}T���8���X֒��dî>�k7h���K�D6���u���Ӭ��K�9�Bc[�Nz�`�˭ڤ]D�!�w�c]�dX^K��S����n;i�L���&	�5c1b��?7a
���15��N;D��2�D�����(����?�ݨ��T���;]I.�&[o�G��xG�מ�@�ؙ�f� {��bc��O�;@��/71��C��-Lv[nV�$?�C��叢-�9�&F������}���K�!�!=%�#���A�@f8���XF=&"����qM�U�+�M/�k7�y��P�E�"!gO-�|���[����Q���hh��/)�>iS���UR=�Fk����ƛ�/Vמ9<X�$ԣ3?��k�!�{��w�|Ш
H{i^��g�-� ������)�t��[b���'9�u�G�d}�ʌ��aj8���b͝YX�!*r��P�������!��"��eW�J��@ϳOB]�������A:��߭бA�)� �_U{F����˛�@����K�Ҕpy����)ς+*�
B��G��Qܛ���z�ߞ�s��!���~����9��<OI!wq�.��S�>�t�ٙ���,��}~�7��bS�]��d������~H�ogەy�� '��_]-R�5�y��r#G��4��Dw�R ����Z�
w���͵�>�w�_�ՈUD+n�7�׵�	m�?��6&=uO	j��W�z8:�(C.E;��/�7��݁|����>�#�+\�/b��d�Կ���j[�{�rd)1�5nSku�ժ�������pNP�bܟWz� ��vG�$��4i�/�$4 w�KŹ���E��3��9~w�&�5IJג���+	��e�So���}�}�q5R�Ü��P�����ǄH�]&��`��2�M��031H��Q3nE�.U�@bb^i7}��$����X��u��`r,S�M"S����ʾe�#32�Yv�I��Y�S�F� )���+ֆ矍�<c*\03�6�!�"����=b�>˅.����M��$����x}Ry�q�i��=ƘˇT��e:\���B���d$����D]�8�j�#Y�<^�S0��URƷS��YNΑ�2������өx�s��E��Z~'z:R�@��U����^����+����z�UH]VkU�5����W�K�2����L�����V� �H��W���\J�7=6uq�6~����{���3�s��:V{x��F��\�.�(2���m}���auQ4X<i��2g�����ݽ��^\����@u}ܶ���3!r!��x��+�PDj�s�4s(�}�L�*����g� �+u$D�Y2�ӛ �ژ� U7 ҥ��ͤ����OV��3&�Kz�`��q]�H�fG�+(X�D+B����TV׆iΆL�;���Ifl?=��0�J����
�i��������6�:�����q�g�F;E�a&�
��[���ˊ1dܪK9�S�48l��̳�i����=^���!�lf>��=H�Ź>\��Q8�	?��d��� �ϙ�u7�z
(T]<���l��]��~Y6�a�z�z�>I6hznΩM�u�����+��]]��чp��tl;��挷�0D=L�Z�0��A�1�?:.i{e�"ķ��)�݅�rpki0���s�
\nx�2t}$�g�^�/k�я�SS?ö�I�_Μt����J��W�s�N�B��~��f�L�0��"�,r/`����m�A�c�-��+F1�GN7��:i\G���������y��jd }���Ui<}��E&nš�X��.�F�-q��Y9�k�҃�`F�+�� B�M�XX����׭���U��T-Յ�����)�b�R���p�x�Da�*Y������vRʬ�Z��!�#��p<z'�I4��p�l�G�s�W�.�tF-[����5��k:��[�U7�%0*�%��nOE��憅��7E=�H/KB(�h���	3M�j��%��ʞ�O������oW:�����9>9];fs�{��B��az�z��hS�|}�����",C4���Y.BEX	g6�AYE���mG�����cOdr���	��V_��\QZk e+�=8c��['��P%��TA����x+���%}b��:�R��frU�t�s�����b���2��x�v�^����`v`���c��遇`k���7y���V��c��e�6��|N�$�|�W����eYu�Vk��4ûf�ʧ���tj��2�W �}�F�7g��w�a�<KR?{Q3�6�����h�{e t�V2�o�9��%v^� `��Q���ro��/eecb�q��	l ?z~�.8W�&k���(
��,���S�p��n���� �}m�i%}��)������`i�� �wg�r��ɝ��^C�B�W��ϯ��9!)��+�Q�V>Mɯ�Yh&op���qjO8�s���}���M��G��O�;�P�S���	d�Sw������Y�7�2�C(�%����q���Gx�c��>j���h�f�yk���Ҍ�B��E��r�J%�kx+��y��!������[X���\�uw�PD#��
�D�pC���8U��=X�>]6�A@���l�dy�f�:�z'/�����N�*�񤿹���m�1p��~�ޘ����l�Z'��xQ��m�i�0dM���el���m�tYF��$�R�46�G4q$�h����E?������EQXս�����J4E-��0� k����.��˅��ipq=��Z_�Nf�8���-��$v#��&r��jL�o�B]�;�ŀSA�h"��B![:Q�ե~57C��C@�7��G���=DL�ffO� �$���0'�x0e���pWɜrƥ��C��F$����Wdqܬ%Ur��ߧ@�%H��H�C�d�Wܵ�hNҷg;a���\T�����F%m�@3�#v���)�F�����(Ȝ�ؑ݌g��.bF4�8ց80*h���a,z�`�,�Ӽf����, �?�pb=�Ú%�j�5u����Z�|a��.��F��"��q3�� ����&�-�݌���Y���*�0p=����lsR0[[��xK2N���G��.ŷa�~O+���N�
=������r��Am�= ^�*�}�����q��ׁ���RT�/� ����4�I�4��M��8��߸%`ќ��i#@�AC�p� �Ȝf�h����mp%��/w?~�8����w�'So��kC��R��	|���u�L�=(:� ��ԥq�j�z�&��ȲqA"�(js�Ǚկ��NvI��b4d�)�ё�K�Y�=珻n\�e��7�z��!�H��&�?8�>��
+�vs�VV G�7�'�t�ܤG4�����S���y1.�T=sa^��f�����i�׳nDPsS���wNG A۩DQH�^�V�d�˺��_6�N�nV�$ȟ���@���"o�/5����-I	4�×|ڽ�ؿ��������1T�sͭ1��?���A�9)����Py��ކ-���B�ﮈ�;쵪*x�0s����h���9��@��,�u�	����"c�����h��?��w8���}#�9S�I��~�H�yB^�j�-�O�L���հs����J�-��0k&˵HY00Bw|#J�$*o!I�^/�>�+��d �/qp!'%��R,�e�J�^J��c�ͭp�2m�#}�jHd�U� <�T�G�G��� �[��6�2�=� 	��(b���*J ����|.��D�w(����;���O;&��-�SRܟ_�X��U�&l�c�S5:Ӥ������;c`ݗ���E�2�m4ԡ�~U ��/�	��1E���?����?���XX6��}R�T�{�j�*nj��\�-��)NT	s\1]�SQ��d}8c�\�&��X�HK�N�c�%k� �WL���)�z F�6��8�(�x}�-�O�o�=~d�|2��=��B���1�$�U >E�:�Fѻq�?�+��E����\�BJiz����v[��g��'!f���A?��;(��6fC���jF�664���Qp��|"�]�dW�����&����/� q>���hE�?��m�8,�\J£;�2�v}<��n$&�Z;u��?��|FMlO2ӹ��6@��f�;��lj��"�G��
�Y������ �V�ň$��y��7�G���ȅ[f���hE��(!L�D��E��T^��Ҭ��9��V"��<ֽ�
�D]b@��c'��,Ј��P�lFy�Cg�~��ࢶ��Ƞ�}�Q�h�H�#I#yvRƱ��㻗B��.�Cy$��욇��X*�zX��g�� �����1_�[\Ĥ�ӱ〥Fx��#ܛ���M~���0��q�+sP0�O�f�]t�!
�	�����,����4Z��74}�-K�c�=VL�؄- ��aՉ���O5��/W1`�8[v�(z�oɫ��F�8����m��'qD,fA��O�׵��eh|��(�hҠ�������U�؜N��M~-���r��XlV�D�%	���L�R}tyO%秴ڦN�<��`������RH��#���xN4[�;G%=J���A���ޟ��!�M�O��(Ȃ��+�5���Ŕ��J��a?SЀ��ʤ!{M}]�+}_��[��g�r\!��0���o�d��OB�����14�°�b�Ql.�qN�Z9���o��Đ��6V��}|��(����cwm��s�M��@=N��4�O�)�+��dg�5��������TJ��=3ɱK/�k1�ck&a�Qp�n|@��Q��#���S^����Y��}��s���
9Wz�[U���M�_��2�e��`T̀�A��K�%9�w���eAdGA���4���R_��"��.���J�
롪4=���<��G_�H��\��[��tB���? �5�KS��<k��l�\KC0 �h�,�;>�Sh4Mֻ`�Q<�Ԗ�}/�W*2��5JG���l<��Џ���a8�`(!�˽(�Z攣�y:�O��K���D�a��F,n�����T�H c
����s�*��=��-����a�wtS��r���6�>;	���a&�2�������ͪP�lM����r$��. �#l���HC�h�\6.[m�A�Ғ��~"
c��D�$�#Z147���}7�{i­ԶY?0�<7.������D~'C���]|��y�^C�	!��I�2-˺ςݤå��yރ2�� ���r�S0k�"[���iH"�/��B<)�E��hvR?g��k5
,ؐ��t5d�h���D~@699(���n�/���nzU
%���8�7��� �J��=�	�T�l� �>�%<�^z�?�N8�*�аgv�Gd9��B�'EQAS���6�n�D@�Cqm�Jt���{h�D�Yq�Y	�����V�sHhp4��	p���>�����N\%ݞ��ģ��#�
�R���,7���ށ��ݳO�b��W�)۩����*��yʝTt�\��g��,��������5���Caˈ���am<���Oy���Y�10{T��w��}K-�%�u
d�1��cK��P��T䀍h�B�}��);���BMc:�	Ɋ�x:�S6>T*_ĿIm,���������u�k�6j��6�%|�C�R&`��
A��2=���>D���ĸ�1���ϟԅD�NfP�exڌg�N�!����K�4��t6�=m��S�Lؙ|ʝ$LH���y�^�_��������%�z���ȧEn۾).K�~���{�8��ŋY��b�t߶3�u2��,��}��6�����R�0�z��Sc�h�?���b2gq`�u'�t�Vu��ke9�ֵD��Ew���d1��@[��mԼ�r��QٰSq���*��ʹ�se����J��=Ï��dF��d�Wj��V�2Ӓ��[[��h4~=�:]��(��i��'����	3=pe���U\.3��S�C���Q�#�:�����PU�;��O�=�ì$>~�	#ux\T� q��Ex�qU����f�W�g�e���.�GaI�1R�m4��Mؽ.%.�j�	��R��x��7+����˧V�Ć�p@����t6��gO���?.�Q� �����b��;gwX
�����A`+�����'��NX��WwB�_k��@J#�.3����Ҧ����J�s�Yk�G������0S@6n�)�w�X	:�%_��n�0��kB�I�;e�'��ע7A�6��ݫΰ�=�]#[ }(�6wO�t�����V�K�g䵹���U`f��"���ǚp�?;s!��^��^Q�<�-����P�+w@(���>��/e�=٦�_�.@V���-Mr|H��)�W�Q�hN�?�ù�����P�����u�bf�+:o�<ܷ}'�����f�\C)?v�S Ծ�����^����N��m��N I��Уt�1c&��z�l�U��A��x���q���Y�Ǭ�>r�bˍ󵓘���*�H�i�u''z���L�,G0Uŝt���S��2����}:�!�s�eFv<e�6M:
�CK�+�����2Z4l���g�:$G�s��7ꑚ��?���")c���؃���gE�b�B�]������v�(&wʤ�V���3�����d�0����˴��68U�4����1·.���9'��_��h�v����c#t B��߇iCse�/��=x�(Pm4�p �ql}I�	��iS0������h�"˲�f�5��]�>S��I�4�\+]��<�n]�����~�p���
�;E�c��8�[��,<�(�3:�|
$)���h?(Q�n�Hăb�	����VF�n^�$��l��+�!%��G����<��{����O"@�/���*�ǹH5EU����Θ�����r��*Nw�>0�G��WR�x�!�Ӯ`(��`�w>F����~	�{����Ą�C]]�ı�Ię��8��֮�[�@˳^�Yʨů��d�cԙ]�+��g���g���6JI���'�.�Y�@ct������ƆOV�ց���x��;:D�y�4Ī`B�t�|<v�8��:=�!��b�%�CEXKʿ��-�q|F���1ps� \��FL:��v�խ�-�,��H��%ٚ��Qn}i�i��5a�J3�홤�X}��>��_G#�L��Z�g��a'���t`0��e6�.� )I����Q��Q
�<�/[���r�S�8���T�kM��K>��攗F�|:E�lۦQ� �*寈�|u��W���|��sH�-K���}P�C
:�'�n���rB�»������"8���?_�7���ТO&�w�Jb�[��H	�yX�r�q_Y��IA*'��?B@�2�����0N�����E�_�\��!.l��)@i�2'�	h ��̒$,	yS����;�+5n����Oyr� ��)�dY-�����*t��i?��̖
_�1�9X��a�J$Lp�[�Ar��d%��X�_�`xL&{��r�Q�<
i9 �j��+��ڶp$�v����}!��bJ�6��w�>/��sܠ3������S�$�]��&����Xʛ	}p`�4Îvu"�x<96���!(D��Q�3e�S"Ş װ�9�c/ܚ��j*D�=g��e���G�W��bz@��ݰP��=b����un1�<�[ X�jy܃���Qm'$܊sz�Q.�'�(�̘�=G��Nr_�%������ *'�1C,��`H�?�����<�d���Rs36q'5�J�ɾ�eیU�ş���):5|��3$������
����|")�ԕʪK7�kiȱ�-��&P����-L�l�8 ��'�W}l��F�'y��pe�u4�, y*�J�(�EQ�)��W���q�LҔ�W&����i(�����B�"4�XDy����v�k�i���"S���-� Ǘ�3d	r^͵��ȡ8�[M?��Fen
js��#Q���V�Y{��^6x�������L\�5F��gkV��#x�*����-�Nn�T�l�taUR6�q���W��P�j%w�|���z㈦�����8-�
@Gϣ�	��R�6�m߈�x
�6%>���}�s��l�T�M���@���*~y(f����y���
Iv_&�};p�W?�6H���:�s�ט��p�2"Tń�,����${�!�q�q�^�H^��%H5t"�x��pP�����rM��n����GAyOm�窣E�EX5��_j$�T���W�2�� h��a��\</�m���	�h���W�(#3(:���<%�����Oc]@]�,
�]-�N��n�LVS�Tf2|�x8�&ƫP���aαQ�<��β@��-�[ƿ=�I+�!�r2��4����� ��_�k62��4K����Ð1~*˧r"⊳�b���SQ�$�;���'�0ڣ4W�@��![7�����a��@\��$4o�&�pA�	O���������C�8����ˡrgG���k�4�.T�@<�̏�����j�ٷ�$H3
��}��3���3o[���b������-l����pS3\�;9��t���wQΩ��r Fz�|{~�%�XO���}�/K�/($�LZ-wI�6��L���ME��M���J?�fdd\����o���)띉��
n�#�Gj�D+ض2:��#��1 z��)�_�k�������?�]�+��L�Q?�̓Sڹ�I4�$���"J�y�@H[a�AT�:�!>��ʪ�6R�-������e����y(D&t7G�`�Xt��<x��ۑ1Z=�v�������?�'�������W��ZN����}� (�)y��V��'q*������:��	�@��;�ݺS�4�Pկ�]�ARN��Z�(� c��LJ^�	5��l��y��Z22�z��׺ͻ�/�Ņ�t@'����� ^i�fI$'_0+�]����4V��p�� E�;��ѯ�}�U����<	(�����;�7b���on�όg��P�CC�-i���9�w�`����rzQP� ~�3��U~�;�x��Aa4�S�H������"��ѥ��Bۯ�[��XS)y˦���2N�a���	��F��uv�8E׿�����*.2��T�3�5搢Gqq��-@F*��X�jQ�eN��P�����-~p�8��_�'�ߍSԬ�8�ց7����M�GI��M`WU�l�^�0���]�/vr�j��~Û]p)l��� ���]GO߬" ��שz1J보�i���w` ��DXc�_-֕0݉@�\�;��so���ό��	�ۡ3u֑2�(9�h�^̉���e�` �0���4��)6���Ί�5����I>����uq�I���F�dWU��E�ƜX'Z{@�5= 7�
ތ3k*a����Sy��+ށH����'�e;����,���g8����
��(,�`Vo�AGK�}!�
b88����͎i�x
�pZ�a8�K�U3��*E4�<l�b������N����lz��q�7l؎�����%��i���[��A㶽�nv��Ԣ]̯X�MzI��H��K>�P��9�"���v��0bg���Z�8����p����ڴ�i�ד8�x���!��x�"��P�&�-�)�$��G���2�������)�==죯�Nt��r8]�Rļ*�8�.�*��;\���C*���h��!jj�m�V��ܒ���s�81�L��Z( ��i*`��ࣄ��J���Y6�ʞ��PU;��@��⳥S6�}m�er�:��`r�%�V�0��|ae�jT��%�\]���8�F7�}�(I���MpQ��F�T�]�����Q��E'���ٶ8Hz#��ۥB�m<�z:ש�}��;���3�p$����I&��q��\�c��*t�`�#t4�ߕ���t�K�?zw	�X��X��x
�C�]�e�&������R ���2�¦���]�1WРq�zr��+e���[ǩG_�^T7f�7[Tp�w��h�1:�.؃�|�CS�|���7�]�v &؛n/͑m��b⸺�'@�d�s���p��e�n�@i0���z�6<: �7� ^����
�O�j^��@�D��X�)py�S
���0�����A<���[X!7}H��A)DUR&V����u�I�gI�8Np(/��z����Lf.�S)�_�F�/�m B[f"�\(;Zaz��5�e��7�}���q���(`��"�x��KWaP�U�I��7�����6�'����<���;�>�����5�*���\��Oz�oq�_C`!1۴
�[ֈ��V) �cs^���5InX�\�Xo5���ZY�JH6�	Zi���7TU��@����e�-��"o��
�<dM3��9�"��H,���`x��P1�p�=��9~n�rD?�IfѴ��2����-��Wz���UZ\���z!�,T��mH[����p�Ú�!��)P�#h ��C�Iִ��������ԡGq��sQ�)Η��iûu��:��=���ӉX��K�v�KX[���-h���	E�����k����r�꽤dL���ϯ�R<@đ�Z��ǋ+�d�D�{>W`ߜ�U��8��ɚ d&f|^�?3�zy�])�%�q�;.�rz�gI�d5G�Y��@�e��l���c����Rʘ�/pY��,�0+D�@gZ8�z1%�#E��^�/����s<��JPȹ��Y.K{�o�A�I�5Z�K�5�� ��_��oV�O�)���Ԓ���½P��W�]�O�"/߶n�dl��?J��Ujdw�:���hO�!h�b�ttSH�a����JY&q�5	x&�\�Է��4{L6�����8g�mԎ;3$�+hw����dCYϳ��zqc
�.��22!��ǓD|���B�Vr�B�{��8MKL ciEu󮯲hoJ����R�VQ�n���Pk��I���N� p��v%��P.�ʶ������R��n͜��˝_�wʤ����'��J۪zM�^~�!�(M鵔��h���Cv��fC���C(��-��n������\[A��cI:��{���������[��O��dI�|�tb��
�&;�z����Ϥf�-�-�F�ϟ���?�'��<zwһ�!_��'!�Z0����A�3X$�#�؛r�����$�ϴ�/��<���u���I�(1������1�ϐ\@��{vq�'P�ę�Z�´��ת���$T[c�A%�iȳ������d�7��uˏ� �Q�X�x��ͫ����V*.�I�����R9�/6p���unV��,ei �y��g:��}���j4���/z��~$��5,j�cP�����zn�r�bW3(���򛴶��q�)���rjl�W�����,Ӟth��2T���<7LCu�I���=�{`g�1�?T�1W��W����bQ|1���%�=�kQ�}3NZX��.�)������J}�����	�,/�J�)1J#�tT'V����C·�C�s�h�$�	MvnG��`��:���)ة���TG'e�u
�i��m������G�
�*�� ���T�Hf��t�[w�vĐ�h�XO�l�#u�z̜�ii߹�D�jf�m�5��;�^*^��9P�|�u�`�t(,>*i�K(a]�,�4�a��Sב8��b�v|t�tk�������^l��6cŐ��s˦�D��]Wfù�0%��7��[jiI��1��<�2Nw�����Jş/������pĢ� -f!K۶Jӕ^0��v��j���@�X�pR�c��5��;I�`V������UD����� 8 �=�<D��B��<�~�L��&��29�� ����s4��\K�5.�3r���s�Aᩗ��l{�:NO�j��[��811J�8�Ƕ|w��?P:|u�&2��yP���#����`��X:�\�$���s+�I�fl���2�?�%ba�����2@�)=Dy��k�~�g�o�d�44��v�"�5jK��RX��~0�@����p��z�Y��ڋ}�1B�������zO�싂@�e��$U-��"��f\
*�b7���Q6׊Z�0��/�2����!�a4&�BtW鼂4�*[c�>�քz:��
x��_@%9Ɍ�;��3W��fB�  ��5�=SF8pPD�������ڂeڶFTFL�m�FPFYQ C�q+�ά�_=�dڊN!���G��#2��;7mz��%���ˠꮅt��w�X-G����Į�kV��u���#��=��b�BϚa����&�6�F��Ɍ%�顗Q�,p}D�t��:ƜXy������o(�����4���������,�m3����ґ^�Aw���"N���uG�, ��8�Z��O��uM-��p�;p��Vhc���"T(��+���)�])����^���qْ����l�A�j�@��m	�a���a�kN�p+��2_Q.�~��j��f���^D�MϾfvU��V>,��g���!e*�$�0&�� vtĿ[DUeω��QN�E�X>v��㾵��	%j�B�?t�'�����&O������T5��ٜK��������C�\�JK>�B�ҟ<ߕ��Ị���)�n�n2Ӹ`$��PQ���r�t����]Ɲ�W�v�Es��h�2w(��P���#QH��b,��j�}k0����NB�n�8$Q�>nݡd�K���ST��%ǫ��}D+=��"�c{�>�,P�f��N�0)��7���aGZם$�Ӏ��x`L�z�U �\�a�-5u��[�a���#f��Z�����G�Ɠۧ�q� W�¶@F��Xi�Z�×>�1�-4�K{i�%1:w~�}%O�d�Pk�4摓��� �����qIM�,�!�����?���tx�;��Ee͂z ;F��j�)@��k�Mu�)t��%վ�Fѩ�Jo�LnB4����/�Q���"��`�
�u��~�ރ�{}�m	��,k��eR�r�+�B����>&��<^�
d��ұ��2f,�d��3�KbH�D_�d8k�&5��v�D���U^�C]��a�S��-��X��ْ��*I�҉�T�a�\�ܭȦ'�T�Va<�������g��G?�r�ɬh`C |h�q����x���[݊ �̺�X����V��ʖ�B������JmA�z���$t���t���N�g(Thl�Ǉ�*�uv��rwh�&*?�$�$x��	G�z���/,ۙ;��i"�J���<(��@����R{$���L�4�����ɛ����0�����w֍m��n��j����#�}�Ԣz�0W��hT��$,T_D�����B�-��B�+�Z3Y�ԗ�v]505ѝ궷����$�^E�̾�� Y�U��;��Ǟ�6��)�<"T'�L`���Gi�EW8������x� �����"�w�.�"L�)Ù��	�&禬f�b<��SG(}N�����|�����>���
s	�6NQPW�|x��)$��\*�R��)�HVP7�o��ä�
i�{p�ބ���OVx�]]�9B'���R�F��wZ�XQ�<D�Z뤧����k������𜝅C��c.иcuHKV*F�|BeA�k����˪�Q�]�k8AOƞW��ۈ�1O�A�$J(�+��tq�m�w.���ȡ�D��k�tL����hB�*&9w���㹭�J=7X_R<W�V��ӭ8�"�d6_�����Ȉ��:IǦ5�LM(]����2�������Ϋ�C�H���T��]d
�[!�>��{H��5�3���w�~ĝAd@��-����n#��"T��fO��66���r��ϢG�~fq���UK�i�jɭ���jm�ٚg�m�mdN��3f��&]�r�Q��k~������.k ����n���]L>�`��biʹMn� x���>����_Mq�|0� ��a�޷��f�z%�U���>*�-c��\�ưG 9�Y}�� (�0�Hw���/q$OɎ_Z`�sY�)9��
�����")D_A&��^ǖco&%���M��e2��5\�����Y�r�*NbG������?8T<��8b�>�GQ8�Y)��� a� <�Si3I�S���7��-�w,:�l�Ś9�Ri{���hW0�Z�,K���4ޓ[�I�f"�{��6q�?����t��0m��5��� �! �f'� ��ty �Yd�!{��a��K�c�;~I�_�H�R8ZB�����)�Nd>Wa�ϔ�ģ���K���c{�T��Ȏ>��������F��Cf�&�/�ܰѴTr�4UF�����+�=u]�O��2�K�7'\�B"� %� ���1��q�!����\{wg���>�$k_Jh�d�Y���i��zr vQ�~��G,�� VK��ƼM�����hyH�j�e�H�L�P�����i]��G�-��.�����d��y.�2䓜P���9��q�Ļ�p{O�U&&o��2JiW,&]�ت�}��ؙPK+����먘��D�s�cT���>�~�*1����a�&�o�	�ǧ�ٳCP����x�Q��\�߃H]I]X���'�VB�*���}�� �Db�>�]\&a��6����Ӆ�ܔ�;>�%oB�/���W�y�y�x����~/8��O�y��h��a��3 �x��.`߿yE�3:6�[�[��/.��5��p�O�|V��]k=\	H(L|>+�ͤ*�E�瞞_F]�7�j�I-#ڸL�E�x~�y�J9�Ipĉ?h_^�LH.��Y�y���������7�Z5&��� Í���D�`�|�o�~ȴ���mt�<��u�{�Z�p�	�7������+��'��Í4�cF�-�Z,ܑE���L�^�Ďm&��
=ڪU+&�B�{��:\������n�C����F�������X�7ǆ[	�_ �w�`M�+ξ*�gޞa.o<��GЧ
��"��(�?V���r ��wW"����X�"b0l���ĺ:��>����mE((��Y�b�=��'�ȹ�BO'L���d�`�7!i,
���_�$Oxΐ�pQC|b�����M��j�Z���R4�1��mN��0�(�y,�ʁl�6&�@tNh�D�� l�~��g1s����D0����E�"�eʼ�l�ҝ!uie�T���yA��"�o��uJź�mi�̾;KN��DA�nZ,Lh����4���U ��L9�Q{�%�ugo_�x��Gk>w?���U�@\
�@�Sl�4��u���ܡ��H԰> �n�:7��2)�BA�b�T�O9բ[�w��ϳU7ZxܶN\n�w�~�IϨ:�4��阻?r��M(��D}��V��������(�����6+z������ي����ʒ,���0�3��N�HbK�H�kWh�}@�D�esQS�$p�6���*\C�/��n��{!PI:�:|��nI�D�!#<���*�}�S��?{�R7�������U���,,]�N�s�0�o��}�B�%�19,CE�)�~�g�\Ŵj�P����J{���l�/���̂E��v��:'_@��I>����D^���s���T� �7Nк�Z`bi�f"�k �V쵕�g�=�Z������~���-rFL�=��޳p��_�`PJ8&��$� ��3|c���R�����2�����Ͳ6�J4ϖ�%��)|]��"��3c�ѿ#��߳U��t���g���=�Q��)��ʒ?�����	}�!;�o���u]�IԺe��W��ϩ�B5��2��K��a��v@){�W�ѧg����u�hɩ����J� ?
��ܖB��e?/��zD�Kj!���E�j��b�"�e�D��W���+>���Ŷ���A���� g�>�+%Q뫂)$�����0��c�yW�6���EPc�y�+���϶���$�wD�2z1��va�u��yj�V(��;�o�H9�Kz�d���z�ޙ�L弞=�ֲŇ`�ڣ>�S�,{b=���Q^d;�-F�|��ɸW,�;R?�̯{��� ln�8e���~�^��&R���zk��z�/���(�:	р[ޢ0�
O+�����4���B�g�;��vɚ�W+ˊ�/7�m��kIވ���3ޟ� ���`m*��a����Q͕^���ݝ�s>�O�h�V؟�[���;!�U�����iT8� y��zKOS�(?ޥ�Ū��*1Y�VP��({	��i�doI�M=\*l9D�GcɼQ��2G|�Rq{�z�֒�ֿ��9��H9�qFZ�X�����r��O
--���W�&���;�x�
��Y}qJ20���x���Q3��m��*� A��
˸Kll.���3�r�3X�>���dF�s�g�)H��!A�����o�l �`\��}�R ������O-���	�}D+2VN�=l���eYoI^�`�=.��L\�;�%J��8����!HL��l=� L%����/����V�ȴ�$���t�s�4� /����Ш���o���#	�o�2Z��%W�<Y�A�R��C	z�r�m<�5�2W;�{]������ �Ƣf^�Ԁ\����|�q���ƃ2W$:��d�3��G�cS��i?�n6�2�;,_���-{2��&�.���<U����; �rN�'�?Pe��)/�W��$��h��I�BU�]����N�z�O5��*��ËXq�J�j�X�t�xt]��6dv��rM+�;�BĨ�
�|d�G�L p2f��j����e���Ͷ6,H�� 'iN�%�� �qhhx��ȶ@9���Yܧ��i���I�����B �$r,Gч��G�p�9�%��'<Qё�H�ی^+���3�g��ri�h%������Æɥ>˘�#�O�I���(���5"����m"
��,,�Tg�ԋ��JƳb����6N/�����T��Λ��y5�k:R�TԥQ�D� ͉B:;6�:�zh���7ӓj��6]���g䗒.ş���i��K񝎝y筈:���|��9]ņ���䭨1�!�J��*d���cr��h�d�G��Y��M�8��qU�!5��<�_��S������f��n�C���Ҋ�ooi��gd[���Xe���l&½v�g���P�+���i)�5+�Z��H~�bx]E��v_Z�4�4�H!cИrt7Q`r8 /�g�\T<�WV�~5H�Q�����^���)���'vb�'H��;��^������� �=t�2�����+v��ކB
^�����q+}UP����]�C�������(�����6��ȱ>#:��X�I�������(����4N������n	d�ٶF���9H��-YeL���ˤ�M��O�/�Sn��6vqU���x*�@��2I͛�ڒ|�8��F��C�αH��)��R�'�-b>R��BHj�	/#�!�Td|�����qAk=��&�ߒ	V���� grA�`�L�U�����7����T�U��?��v�	I��?�w\�'��{>�֭��Wg����Ф�w�v��i�����|���7�����rN ؼ��pP��)4��� ��2F�s�%xA	BG{/�I���f"�-��{-qEf�d�/2ʃ9���7WΟ����,��M0/T���yi
%�X���s���'����T��v#V��<7y*ϥ� 8�:(�����(�}�R��K��qr9�N�k�ب��9mܼ4�k���L/�>��������!\�p��W�1m1��r��כza���PRO����a��e�����A�N�i�#1cȓ6��ƀ/ы��2!�RG�u}pw��G�g�j��@�O�� _�d�����7\��6�d�6\�j��!aD6��jrL"M&�A����g���T�!�S.�Ҡblr%|r�-�7�q��|E;�����>6�;p�{볩�ڝ�8�m�}i���qy3�Xߔ���oO(gquYHL88��p��4͌����g�SW����>E�-G|�`l�#ͽ�s��V�^��[��A?�+��\�$D_�U3�,����0h΂8�%�_�t,*�`'�^�3V�xW��F;}-^�hz�2i�jM�,�����cЁj(t�.dW�6�A�f	��&����wK~LT~!��c B$��)�M�e�"�mL��7��ɴہ:h�ߡ?1��4� �};"%Eonpg�")t+�'�A'��1�h޹0�8�Q�a��2->:����E��pk�޽�Ol4�p�t���C�����:)�/���<�u���;��%v�A)�98P(��"
����ă#�M��o��y��Зf�5�ȑ��]~��La����V�@���H|�"Z8g���j*<�o�dz����톒�r�k^ M:��Q��ޡ2C�bּ���cz�ds�̚(�n ��E�©���_�z�}(�0iP�)Sw@�@՟<�s�l)g�)`�v�~
w�PR@Ӯ��X�.[C$h;� K�D�U3e�E�FltE�!��ܘ�L��A�Y��-�aHE��+$�7���F� q��S�����_�<�u ��1��X�g$g|�y QR��|Y�� b�!�=,�������̱�s�j��7�#L튋�\`.:��K��a3�.�#����4;��߭�"����s�j#c�%y�8 ��`��E������va9�#��!׻z�苷@��F��HD������&!Q���aЇ	2��}�sż2YEoF�x4^Ƌ��w�)2���+i}�mRR{b8zl���0ƢD�P�%�����%F]�ɐWS�=Qꊮq�4���q""����?.��A��&�^tr�[N�WJ�D,h=]d&���SI0���A���\e���O6TBo�%ȰO�)޲{Ųʠ�
)$����xM������$�5�����D _�72z��OCy�0��q�}پM�N�[�Meh���i�ya)BQL.m��m�'G�����s�N��V(�:�N.�1H�&]��Z}��C���<�z0!�(�����b[��}�7ñ�|"&+��(�o�I�<�L*��v�C�!�	tIc�r��﬊c�X��5k�����
��ۈ郪-|,_,m����*���|��v8MyW���Ky 2�(}ƹ���,;胍�@
mD��W��� ����J%TZ�k��7�^s�T�2��/��Y��隈|�4ӕ�,��o!��d;	&���˕�����۬����L}r����z6Eb2�qUZ�+ßrD����0o�/f�l����6��5��\\|h���Efr��
��<��{�#����>K}9G�<�)�9��h�@��V+�wE�thi!ʑj"Ad��CD]`�S@�R�1�E��3��L~�!Θ=�kct��ah�-4�v=���Z��mw��@���ފΑ�{�`�7��T��|%0��xJ"
��������{���u�
:릎TOB�ɞ��%���Źx����_�=��XMZz����m�Vu!>��R�����b���H�*���.I2 ?c~�,�6x.u���N��p�_��X��}��f�d�
�>�o߼�1o���u�AZl�����}����%�ʍ�/�����r�����MXܞ�����b.��,� ���Z���=�/�F��5�J�-��C�%�4Y*�:���D_3��v���0/]?�X���g����PY@�"$���}܈pGl�b����z�f�	�j�3B{�?	f<>t��8v�}B�c��̣T��a���`�M��l��8����zQ�%����tp�
��OX	����)����y���Y��������r4w�R���S����6�(���H,Ԧ�:_?IM���x���2��A���dq<��h�|�eF]�UG�M�#�{�,�֭��&�����h
���!�j��9�8/�������u5J���4g�t��B"�����r_�����N9� [�C2�ռ)l�~����,|���r��c��)��ƀ�EN�5�K�ˠ�b�������H������qw��qM`ˇ5���)�M���k~�V��1�e�1� *QH��s�G��v��F���H�)�x]:v�/F��Qk]�%�^xeM& Bʢ$�B0�iR	b^�m�JO���-Qa�<$6"zڦ#$�&��{ϕe��w���#�v��� ��`�K����欇��yeso�:�`!�p�WϽ�C�n>1j���ɨ��U��n�n�!̆,�n�.0<�d4-�_5W9�+>IS���c�@"�L�:��toύ���'B��:5��bhĤ �nn��i���OT�"�8 m�¬��x~�(������-�vrF�]�� � u[�B����D������NE0���}G��Ņ���s��d*��Q�$��!1�qؗ�q��W���?RvPN�.}bӍ!2aC�򊟲���*w_>���s����vJ�E��Z�M��B�:��?�SL�`y��������V��%�=ֽ�Ă������������w5�<���I0<�V/�����1�f�0n�$�ud;]�]�]�,ɐY#mw���&�1�����J��wl�m��C�[%#��Kxy] �֬������=I���;�D���!�c�Yi!AΩ\I���g��vb@C"��qo�D��b��n�^/����@t(�ul��a������|�g��N�/�3�a�|1Qr��(oS�����oT^օ�`�V�P[x�Co�C�{�j!�}��$�����;��p��Z�r�q@r�����d���:׻zx�cd1��=uh�O?5����
C�G�)bp�cqT������Ph��d�zs�� ��4�<�J���yV-b�_�|�Γ_����ۣ�j`q�&�	��B�}��]��a��PV�*%Eܚ��/ p���7���@f�+;^u{3�)�S��0�܊�?(��9*�������D͙��Lv
*�6�N/��.���� �]3g��^X<]D-1��(���Q����,�l���5Y>!��t�̝�*����8�>{Zo��x߭��a���_ޟ43�9V_PM��=���t'|ԇ�d[i��0�2��h��zm�S���j��6�U7�v����E1O���5�A.�lc���QM4���������^T�XYb�p	�t��Xv�?��DAcn.Jb�S]괮]O�e�.�f�Z��oW���k�,�AT]l�	�2Q966��G�ۅ>�I{���֖eiYq��$X�4~u�h�qA`@�hV⢝�o.L>�*�d�f�E\4v{���QR:�-2�H�̽|�� �`P	�E�2O����L]!���Ce�]H�D��M��Y��l��%4ȩFn�C���8�Lss���Z�Sºǅ���n�I�s�J�W%z�����uK#�C�֩���ݾ�kp���Lw#�m6X��oB��<���ϯ*������:�a ����H���=p��`��0?8�l8۝2N$��1�-�ȩ�.͖�
�p����7�Fh��-_�1 �}��2�+2���	K���e�ѼX�Ď��QB�������4<�#���x=U��rĿ-�0@]Δ�����h�&Ն-ڦ!��C����X����;��\�Nd-W�tb���=Tv��B�^��Z|������;�d�}.��I�5��Ibp�U}!#Rӌ�*5�*�]A����R��'"Z�;S6�?�o��m ���YR��F7���F�H�I$7�s3���ouO��9V�侟�g����=<I^�gZ`��xn��Cя:K��M�nܙ���#;}1��F��N���\���5�e��aM�}�"���i�x�VOξ���=��Wh��;��i�y�m�ҁA6�ד�~�2�mL�w ����[s�"!��q�m�0|��iA��BӅً%U剄kVKP{�;��N㦍�R4�����!��~����q�xI������i*Xߨ����ʃ�08� k�>��."{��*D�p~2�PB�V%dZ�w�Ƕ�����F��'����r�m������S4�|���D��Q^���(�Xe,֕�p1O����	;�V(�1h���ã��><1?ަ��Ų��w�9�Y�h�w!찌�A�4�3,��Є�A�*����v���u���� ?�����%��T˗�_���UzIk����a�>��	���}�~O��`�p_Ζs��9���2�X��y��?N=ՙ/"�� ��Z齟iq��u�A8����-�C�{�v4�h&�qi�R���r�?o������'π�_�f�,�̤jݔ: '%�g�̶�u;Tq��+mi��xk�9����+73ϟ�;�nq��MZ��\\6�X��~7ّ��_�����I+�Gj�e���B�\�� ��J�-��q��ڼ���(x�+���'���/�S���hR6(���7�M�mD���e�65�������3���[�������_���km�>Ɩ��
v����ڶ��>s{a�]"�W�>6�_��J��?O!Ƽ��>��ح-tٟ���'�fP�����2^�}x��34�~#��6B��{�(*ׅ^`�����8=�Z)?�2Y�
ᅐY����YF�	
7�����t��si9w�td����Z|;sm�ܤ�mV��+X"'�����*T�Lzw`��C�
� q	�}���s��Љ���{>�PT�Y~n۱x�G�P)�p�f��(,z��������(��:�{f�4A�$�6T=ɦC�!�|=la�$���j����ݾ_Y��R��Q�"�O�>5꾡(�2�82�h�o�y�{B��KT0����H��TuS jo�C�0K/,���L���k���9�6�׎$�r�Ɉ�fO,[�a�������M_���f�� �R�!h�j4�ciP�t �@��8J�T�	��vk��q��}EY����r�,��R���l�O�f���NP.�4��nFė<� Gvl���ժ�E�x��BI�e�}�E4�yZ�f�s��<�Ч�)�+���U��X�1�2� ��G/�o` ^� ����f��Č�j9�n�ֺ�vQ����?�p��:�"��\@QnF4N�$G�?��f�pս"96?��}B���ix�X�i�ж9�d������z)��o/�$H~�e��W�1�9����0~�ճ�Wޣfu,�y�-#^�J���vA��kwB���&�*6�s�����)�s�$^&�"�e�{�Pݯ^��6T�D�덝�BHv#�WZ)���^�_%��WB�.��봾��:����f�`�ִ�܁g��e
u�Ml��L��C1��
��r�ݶ �'��P�yzfs!����H5db^��XYXr+m�u�yˢ(Y���:�l1��]��ݷ(:[o�wO4�H.��;r�H��{M��XA�� ������zr	/��(�j��r�xI��
:h�O[Ǝ���fv�C��G`[��@r�ԍ�_i�}���A���������Z�~��熿@���Ț�Hm��宵��<�=�R�����#�L�.�4$"gWF���!bfx���{[�i�~�
`������0J]������)�-hO�i_�c(��æ,x��5D�v��.�/�H�ֈ���1ɍ%�g4+8��l��/P^�/	�0��8���a����<UM��<��9ԁ2oɶ�-,�t(�lKPm�(���3��x�l(���~e�%V�Di�;^Q��10����[�	�f:�������
��z�}G9���)R)P�}JWys:�G�%O?3<8��N��]Q�=�g�L!1	jG�T��=ά�1�vd*��#I,5%�.�T��eG���`�e���;,����Q�G�f4K$;�~YJ��N���D��˨ɣ=���,q&7!����&�}W|$&��(8�_R��0}�k��C���:1��rtp<���I�{�MQ�K&(��a�ݸd+�\)��`����'s��4��|*#�V�	I6�ɍ��Ob��,���E߄JW����`4��N���&x��s kؖ��l����z�&�@9�
s�A�Ba��8��q��0�Y>��c�M�9�t�����AefWz=�O�øv@d�}x�>$S���#��m[Н����:��aCh��ԁ��%�7�|:z�$����n�Q,*��k*5Y+ �WY�[��90	��^k�S�h}�-ӣ�o#��\�ɭ���Q��Y��"l(���触4�7��؜��"�u$:��^�ZF���YT z�_}�A�!q�Fl4 Q�ҟF��%��o�B �#M*QJ8䇿�_K���J%2E?�e��NJ$����k��G�:;CLnIr�6��BZdH�ax��k��sɫ�
#�2"�v���J�۟�ߏ�NUvn�3�&;� -���H���y=�d�@���k����45����M�&�� p#4���x.�'W6�ي���X�����C� ��}�I:/�ƽ_�#3�4 ��Å6�מf�60��NϦ�Ϫg�'�S�%�KQ�7JR�n�Y�I�ġ�+�:9���!�|nv���t"�p;f�=<J�q���u��c��1�z�/r����*U���a���_�V�7�����7$����R��,+kH�,O:{�h��wST<'R�:���%�<�l���/�%E�$����m�Ց{(���?�;s[}��}�e��Pus��td�]8��p��=�'�}jhF��ۡ����!r:�~X�B��־(���(�/���&Y�a,�*zmb����Z*�.�Y '�2Q8�V#}F�-�P��]s|oB��5g��^ǌOWk�_j�<�Nr4�������^��1�k�M�����Tߦ��!+�_m	g�??��k�Q����� �JE%�����>�Vu�����!$�j'��5}J3tƒҧ���6�:X�?KT�J���	W�Z>wl�-�l�gq��I����e A�������F��[����s?D^H[p�΢ҡ�͹^,��+��F<1�l��_{P�w�1��r��5udܹ��a�a��)��W���81ȏZ���Ԟw�_0
�8�eDf�O�x~ �+���屍��zy�Z�+�T?$���D�ȕJ�H��* �B�3�Hj����'����r�Q��e����/( z'�J�qòQ�Z��/��)*�R��E�����U�jP�
�������uA]V��C����a����I�eXf���PU���DHK�+y�v� k�"g���T�����B�t�>�$ٴ��.�hO"�4)�f��7��\V7���7����QR @��bj6��t�*�Y�%h������^���i��c��U��TW�"(Yx�k�8ÜV-�{�ϩ��Y6r�?��Qe�ea�A��ǖ|!�7t��!>x��[��h�=���:K�L�ż2YF >��$�yk��%���A� @F�WlH�b���f�=����EAm�l�L2y��d�X��
��x0�����qN���Jv��f�so��iⶰ�(ͻd0?�QsK\��)�I�E���/ؚ�g�{�Y�k��߈r9����2�Re_4z�\�S)f��g���1���s�1'�H���D��!���^������O?x�y �FX��P�wvb�	?��60��o���e��	������3�p}�ƪ4}�51E*�gR~]�N~�I5�w��uۘp�9���Mq3��!��`���a��R��n�PE�l�m�8i2S�+����|��P�˙U�$���V�K˵h\�&��ܜ���d�.�E������jF�`��d&�x��o�Q�p��W�̤�iG�n�կh'�R��C:d.pbѝt��]�f#�V��i���xͳh�kd��.ԯ�z˩���̅���_�
��f%�:��.��j��qX/.n�|p��QZ烷���T�d��!����Ke�#Ϸb`�i�.
~K�%��u*8���y�[�#���w��L��N�W�V��E��S���9֨h�h��g�x��Vv�!��,����*=diw��7��"�"����P�p���]�%����7Y6�N��ꢶ���|8���&�N�ӧ������ώ@(D�
���5!b��yPz�w�N��֦_������$��X�؆S�0rt�)z���xK;�����(����z�&��ʑ���R�A=7+͑��%���dg.�����P��4 Wni婒w��j!�����U��c-�_���v�ǟ��ir葇�J�� 큈b8UwN}e��q���35�z�Dʺ�����a���#�������K�$�-���Ϯ1�A}*,߰B'��b�/M&y�~�B�Bpi����T)?�i^o��=��܇��K?J+��|	�ڇT~�X�m,3E��P��{ש3�ꐮ�: �0W��O�ܧ"�"-M�c������ϧN3G��
��-"�`�+�����\��;3�Rq��@��_'���'��?
�5"�a�T��D��,����7/\9�D�X�-ff�&��8����	���({�O������f��5"�G:`�ܓ�#(�Bi!����Eߘ���D�4�\`�aif0�*|�"�z���V?�׊�~������pAǿ,�d^���xI)��S)�w.
�zjd`��n7Y�FEϣ��hg /��sK��)�5m^�7�b{�+H!l��^~�v<������'�|�乙]��纺�Q�:'9��L��~f�e5%a�P\
�tq�BV���d��e��S�@_��ú� Q}�$�)�2�)pRg�yE���	�����k%�h�o%&��%�Q�p}Fԕi��%da5e�ҟ��Z�|�Zh���`��bw;���Q�Zu�0?KU�w��H�z3���/�L�?��'0n��IK�x

�}[��b����4��@:P�������*l���eMf*Ý�)D7z,�
�2m���	FcG"Ꟈ�ws�zU�.#��tLA�ώU�d�GT-; ��ֺ1��)	z�u4+��^��-pI����t�(x�Y&��#�]��������-�Lm�-�I�g,���\A���z6����ޖ#���f�K��;�|AO"QX�X��$s� `j���[8Ѓ�̫��`��!ϗXzo����7�34Ze�4�������"�,_=��7�&����C�6e�ۼ.���;P��#%��,J�c4��N=��J'r��t�u`����ek�YMy�]��$�7F
��7�G�k1S���:��U����T���Ϲ$A���G��3|	��xʸW��i�����ɔ}bH1KY6�^/�exVN&�u��sϷ'ݟ�����4F�F$�U��%<���ܾo����aq�xƭbWe��(��K�?)B�+�3���D9���F��v�^r��/��oXz�J�<�����Y����R�[�#M���"�.
0�Ԉ�ټ��xp�.J�~o~�(EI^yU�Zq_�}�e'� Kl�>UX��О�0�\�$�c�!NZ��p�.0�!T#.��o��ǡ��b?���<�y�>Q�}�v�����րj��C��$�����W�n[�<�I͓�
�Djx�A��d�/�-��Y��kE=��������밮����S>�a�{ql'���$W�6$5���x�<��>>2& �\��	R���r���|S��|{`��&��"���%zٵ`7>�:"���K�����8�F�dޕG����j@*�fpϫ�ˉ~�^��w0���~3����;;�y�g0��F�Dg��=N��I�B:i�!MeQo�YG�F-���b0W��e"�uk��`��(CǹP��e5!d^`K }�
����)�������&�
���י�oA֬�9�TP���gf�"��0L�iьR-6QRڬ�	|��gVƾ^L�o!:Z�uU#H��(�^���lJnC(��j�.��0�U/KP�μ��X�Fk�������$��v���ؾh{4`�h���=$�Ŧ��G| �ݳ!�Y�R�K�vru�����Kz�3�X<@����A	���v$efT�η����t��?��<c�����0jz�yI�G���?�����z�c�֥v�Er��]�Z�ʗ��q�$����%ͣ����>ZLi�;ɼ���\�u}�UU.�"�Z<u(�k{����Ş̂��OH��M�ם��]ň��H�0ϡ�Q.��o�ިnS�m�C~q�W�Cq�AҜ�6z��n��nL%6P̾�	J�)!�~/)�������.���%bH���0�B}�ʚ���v�XJ#i�����/q8n/��?<��ѻ����AK�E`)y0s.ar�
I�2{���N�ؾ�8V���g��wTUi�S5[qrOz�&��2Sˆ���%b;�� ��T�0$���a�u�Tթ<�A[j���<b����ѝ�f�?7�9��W�h7Q�s-.ep�����~Y��a9�x�k_0��&&�i��zհ������̋�R�N��*]?/Æ.��qj�����$ �]P�e�	G�j�O������?zb3��{�f��W9+�m��ij&B�9���yԜ�؝�DQv� �	��<Ry��k����Π��1ߒ���hܪQ������d�K9;����E)����:��%`x��Ě��ʰ��-����s+�ە�$=�Q�M�z7�+[[W\L�C�TY��t�|o�w�v��O�עk%'����-ަ) �L���M������σ���s�_�5;�3�����(�rey���>���{u'����3}j+�b-�k��ZF�3�$E������PN���&�#m��1��s�7�9\RA��wQ�|2MQ3�.F����H��u��K6U���};8�\�$s�Ot�k懻�E���W�����'��Iz���|��H�R"��n�n��͌�^7��đ�d�OMz�t�&���f��z��*QP���V��L_�'�c�˯���>�|m��
�1f�+p/���AI�6����ՋS����h�����Ks��+l\���^����{�8���49"��I'+Q<3eY>KLu�/�ʗ?��%�˓8�M��3�;lI���H�P2��)�z�$�!=�ޯ�~�z�"�U�5���Z��ȏ��cQ��t.��$��0uR�uV�Q�-b�3���[X?��?}Uc�-��|��w�<�k�YG�_��3=���i��+C�g�+K��rX�A��H�It�T+�1��i���Si,!ƨ�|��׈3S-F,5XC��2�ϼ�ݘ��c��C;`.]���;H������p�Ő���LJ�
>ְ��X�PN�w�˵;�"6����(��l��C �#8	�p�3���e�3��F�jg8yJ����4��z��-�wf�x7�M�4r2M������l�N���v�����&iϔ����n}DG�&Dp�7�,�B�������?\�������g�^�b�d��{.���葠����y�~�q��W��\PY).�=����sgd����ڍ�i�W(ʼ�3-E��3�(�����q�ܴ�P��g-	Ł*+p��)����6@n��(��Ԯ�`B����a΄ް�).W.[�GS�I�����>�w$��`�������tL*[ׁ�V��F̶A�Yyt��	����>Y��"�`s��P)Z����E<"����CK���!���0Z�'�I��Yʅ�q*˭� :�J+��G�-���s�l$����bSG��q��#�\M�t�|��{���<�z�z�����W��F���!Ⱦ�R��KZbJ�4 UQ`^9��n�����dw�F�mK���6,�B1���(_&�����WO���Y��9�=ԫ,l��.��@�/wY�8�^?�G�׳�6OZ��q�(a�XVX��ĸl��K��ۉ�eX�����h������tj�J�������v3��-H1����PtBԚw��l&B��A��"P _eך���|'��b%',�~�����)���/�?���/L�B����=l�9n3)�c?���&fMD
`�`����DL� ����n͇2OغR8L��U���"����N���e=��M�9�tմ�2-�B�Ҿ�>ȩ4���J8�/��qH�̳�E�G�Ran�x�&� �Q�Յ��s}��l�?�j��
�vS����+���t}�#�"n������6�s 暜l���`Ş���]_��x��G���u��tG ��1
~�$t���m�60��r�V24E�#��t<�|0q��`�*�Yם(u��ٝ��N�3�����o�>B2U��F`���~�AzL��~��,3��v���$��v���ar���K����.ed���vy��P����1q޴��aAB���O�r	���g�2��9G,�3�S���ВcbP�N:͒]�7�G���U��_���S���ۂ:�t��m7��-�z�CF�`d��.n�v�x��� �Q��#��R<�1U8>.����m
�d��Ю2Qת���Ԗ�;�%f�Z~Y���_|\ ��2�͎��SHn�9��뼰'ƨ�Gn��coaJ��Ɍ��օ���>�k�s�^�)j�����(���8#�@B۴a���W�� �~AU�+-�؃���:O0�{��q�����i����xBs}C��dk�s��K\ej��{��.�����h���Chv�d�xL��^kgjM[_��U���ٴ��HT�ҞC�^�C�lI;�\�}ۺ����7al+�� C��5Fe/x�{D���3%�h#�#YuL>ro�P�l��$��G�qR}�����
�`j-$�|ֺBϺ�۪�	�?��ޥ��l��|������m�{�?��%�#k?W8�zŘ������n�ts���y����_:��_��&�x����'�`��ޥ�˒�Q��β�"���:ҀSB,6���F�R9Ĳ�F�\�j�6
������0�^�K ��Ƭ��a!����mg��}�˝9����n�؎p�օ���+��@ ��#Q����P�ɚ�#h.�U�ju�%�����\C6�,E�9mg���ޫ��
��S����� >�V��G'�sj��'6��\�I�|�aF���H���$E�
U_�S�b�T��ac�����bE��H�3��_�U�f�M����1�o��Ͳi)Hj����y�f��]��'ָ�(�]���ۨ��QrA��,�ٖ�s����$a� ��W�)��c��?�����D,5Ok^\[J���tk-?�M1�S�cy�"�9�ǢЋ3ˤ6�I]5��@w�a�k"4@�����Q$���r���y&�	<�Rsc�#-��������nS���з��@��d]��E��,&*_oT�<p��B���q���l>n�������(��?�[w`G&���>��m�j�.�&�\Qe�Q`��v3 �	�D���`�~�Fƞ�%U�-�/X�� �a8� �mJ��'c+r�%���y�!M�В��\��a���/?%y��o~}g�dz��������o��У��x���O�*�^�n�ݨ��=Y��H�
��/�`��Aˎ����ݏ΂o_�c�ۓ���QYI�D6��:��U���*�����b�\=y��"�X��{u��qd��~<(���lVdX�ٷ�&%@4%�5�>C�Y�DeՄuJiYe��\}
?���Tv >���)�J��)�!��h���ʇ7�s�}eW��6����u��=�^fE+� �B����4���ǳǬ�7! #����D,�!�}��W92�Y&��>�����?{:��v�2�i �E=��w�[.@��җ�.L�6}��;6M$��t��o[���:9z��Ǔ2��VG�t��E*W:�	ج��\�d�� v��S�m�F��@��!��N.ף�F>�!�opP�����NVD�b�U��v���������\�{�p�:����`��0t}>ͤw݄�s$W�h�����ӣհ�u�)1<%��sna��Y��� ���#� 2I���Cj���)�J2$�^�2_���W���S��Wlի򳉍f���ZP6s�teQC��-}��Ξy�c�5Y��O�֪G�@���i�VT��X� ��;|��Z��~땓�r{_<� �yJ�T�!�wn1�qz0�Kb�~�S&�X�O�f�ҁ3	w�Qv��'�E�,�34{�~7�V��rq	��^o/<�5�?���Y!�I=���=�e�����rܜX��>f5F�B�(����,���u5j;��Bk��{���(yt2�Ǎ>�v���W���<+��H�LGٛ+�η�n;5$���FYe?u�����)�?S�I�_o��qQ �U�`Ћ[a�#f+�+\D�9��ӈV��d�sSc$����Eg�0�/(���^c&� 6!*����.����&��LGE����\k���$�Iv��x�dKI�Zu��0rA�5�8�T�w��{51��մ�I�G�����y�q��R䬣ŎH�!�g��� ;�W��� �LӍ�yO.�2�Ư�� >a�b=��&X������d�����)�,�:6�/@sZ|Anރh<����{���ū�������ou�o����ț���I���]boH_�bY��/9}Bcs�+����;L%��	>D�G�L�M�΃fT@!f���6F\��^��?f���r�Y�Zh���������v�ͻQ�#�C':N�:���O�k��W���7���hI��L8�JU"=04���u<> qs��Zn㾘���w'�_�|�h�V��ʈ/a4Xƨ#��'W�'�N�.����+��8�m�D>cKaG�R
T�`2�W�~mDln��4��v�稆�Mf/�ҵ�2Dp���v�7� P�H>{�U}3�X���]"R�"��JN��������#�����:����H���y���.iW�,�*3�>�D��x"��� T��QgN��3Z؍�u�?,��m-�0�?�S# �s���:�3�'p���k�0À�_��lw��q�������oT14���ڵ�H3?��Ѝ�m�1d�
�uX�K[�����}�,�;�y�R[>���������;u.�F�|�SH��V{ �գ���Xм��Gj2 �>�/v�z�k5�'�BYz�, 8%��ն����p.�%�/�����y���-q�yL�����m?1��As�mb1�~ ����waO#����F�*�Hm �u*�,��iET��ACW&���L	�T�q�r =�5׆��G^g�� n�Yx�#��50c�Og��ţű�=���L�	��l�'[,�1ˋ�M�}J�$��E2�y��]��P%٩�$�^����ߥ�i$���|w�V�������A�	��ԯB��">_�?����F�������NZM�a�˻`��]oP�_7}����%@����`L��O��|)�}�{�q+��c �oS��e
SJ�����=���i�#�}b"�u��=�/�\Pf�\��!I��İK���Cې�e�L�ڽe������~��seP �,Cȕ:�EIck�%�Vt�L�U��2��@�>e�c���XyAc~�(o���8������bh��Qb��#M8��vZ�,��7s���GV��=�4T.ǀ�D��f�@���H�����ԟJ� 8��$MO����ԟ#Ҧ�|����4�b;��ʤ��2��;ت�Yq�����M�m��N"�)�>����$�^��z���3�|�&:?���`�PzG_Zx���
\�]���%B��Nn!�IK�5a�2�VFK���[�����&�=p6��w|6A�;�y���,NVɣ;o��#>P]�ĸ���f�����ny1D�J���dgJY�=&Jd6�`���El1�n�Qѻ���B )�
U��!�ˌ�ap��H��uL!��ΑL�l��E�9,p�~=��_��j�5�':#Ha�ζ�K��B��d�	*�pb�[`��q�E���-�G�y��H��wI��X�I����J}�eՠ�Xj���}9�Z?*�#y8�s�pC\�5r/ Ӫv��_�8�`f �o��^n���W��h���Y�G����U����� �l�0���ۜ�)�&�í1���ș���b��V��]�qU�  w&��:fǃv�e�� �'��j��v��ɝ�Ҏ/�Z��9��+6/�!W"KH�m�ZI`��C*v�yۍ���\��?a����X�,�<͕��p�j>��z0;=��09���bI�2?�Oܘ�$��`{�
c��c�Dg"��ܪs��t����E�
39h,���q	��7D�؄	�`�"�?��H�"i����r�ЏB��3�����2`!�H�f�M�5�!���DΈ��LT�W	�����!
���^����0i��%-�{I~S���p��"�a�$�0	��G��vS�R.�����,�du�0tM���DD<]VTe��T>���ռ����9~))�+�S�H��6a	�]�����uSb� Zd$nR��D-�p>��mTY92<���8FB�e�U*�vV����z��Qי���$V(�T�
��ݒ��e�f;CzٿS`ω����K�}�;],�u�+��>Uu�xY�N8�pê��*� �C�yR�d��p��*v����+B��E~ϣ�$�U�?�})V ��9l����t�{�TZ㔂�	!��D��F��}�3b�j`=����D�5��<��� ��)�5���H(ￒ�Ge�ަ�)�I:��݀�IYIy�E�ŵٴ����p���(�+��ՌP׺ԫ#��/�N$W.��m�Ci��X���$���#�G��'nV�X��f��WH1T������F��'��b	9�Ew\�����e�g�>f�����d
���y��	q.BH\l�
N%P^��4T�k����+�|+� �c2�B��2P�������H�G��X�,ؽ`��9C�HR��7!b� �]2oT�`Ĭ1q�a~�y�`��9��!��7�lt�$Ҹ3*cS�3bJ����� <�R���}���}TG͈ٲ0J��D�����K�bÜ������	�?7E!o %l����Svpv�-�"�n��|��V�-���>e�T�)����(���LB�	?�M�L�e����:/~a������2_�������I��g}�Ţَ�>IL����y��������	t&S��:�aj�R��/RO'z$~$������Z�KM���n6��~@$p��x�����\�y˗ǅRsi�r��K��h���*P?�J�+++�j`�V��� �z��z%a�&]��6m�	|'�/�)s8�.3Y�zxg�}�@+ >�v�n�[�4Sd�70K�>��C@��X��3��7Tɬˏy3c��ʺ���lԎ��/\Y�US�mQ�ֱH����ѨȀ�Yq+�H?��"�
��L��옛/H�#�|�&�+�n�G(���F�bw]�8�3*�d�1�\�-Va���q
g�J����ApB8��z��`����m���=|��M���^/'j�/�}郸o�8=�c�N�|�a���Z�#I��p~�˪��S[/�Ҍ���w_�}�3,D��B�@U�C�����&�W�s����;P9']��R�\
���*/'h~F��/�{���8_���0�F�f�8�s5GEe�dyp��}#�P=
��&���ٗ8z��_�^3CĤ24��X��SO�1�V6�zT�7>�R��x������"[�]��Yo>�~�:��� Q�]�`Q{ƝZV��O��Yj��3�r��4��M�Z�Ӳ+�I���$e����������g���^�<��oA�ζ�$2Tp�*0)�Dfe(�.��yR�7prC�B^�k^����7�å-�UIA��J�
��Z����O.������`+� �3������[aݪ�)�5����D�x���=��;|�Z�A+}]q���֣a $��F�|�,�.x��e�A�c��*P���M��l~YE3tWl�*�ȐsQu��R!���&����H[�HA_�D3v,e���2�9@[X����@y�z��YK�>�����bF�C�[�����)8���F������2�\�v
� ��r9�"nQ�Ղ^��$�ɵɴn�E��66Ө�?k�@�B�zb�k�}Y3��2�ϭ���ѧ�z3�[��,���"F�Y�X�I�uM%���
�h�"_j`z؝c�N�����f3p��TW�آOaz��-�c��e!�P+�m�֮�FB��2`��>7����:mg��ݍ�d$S�����4������󧀪�OtY�g����O,X��u�E�5z��jq�3̠�����C$8�`<���@ʓF�X�r�9<��vX��e���E�>�j��8=z�IVb���p��4�YZ�rOC��ݭ���#��Ƕ6�59q��:��X��i���J=�&�ft�h�+���cR�g}��PLׅ&2��[Őz#�S���{%&}f4�DL�I�;�	��X#���������]=xp3I,����Ҟ�U�c��z�1$����Z��{QR�=U�!�x�2'�� 1����ٍ$�hA��1����K��Z������5L`�*pq��griu��_>ܼ���U���3�Zz�@署'��]�E��$r,�c I�*���[f��֥xq%�/��w{�
�}:����,嗩TEE�i�i�tI��y��o����EoJ���m�j��������\< ���Y��3$ C��,��D��d+F񄘠������A�2�!�{�Dv5��0u#�٘�u�����>�oDk!�����mơ�\w�t��
Y��F�/��Ĳ�	�K1΅@��lР:JG�{����E�,�!隑 �>�l�\���7�%�t�}ch�V�|2�ade�}�uC�a��q**�H�����j�Cw��F����W)'�f/�Q"ЩW�U�� �^���5��g�����X��jN<���U
����)+����7���9��"�F��M���7����ɮ�ޗ+m%�_�mC��͌	���.�7�ߐ�_���beB��丶.���B<�������D�o"��o���&M�ޡ����6fҺ_��������C�O{��8�#�E���^pON�q'���6��-�C����x<XEݫ>l�(��A2o�c6 ��"��*݃�K�7�y��zc3琯`��QW��Ȇ-�\2&=e����4��w�3�~G�*�8��!����5R��gyS�M!�4h0n��^޹�TF�N.D �Otb�>6c��`��C�ܮ���p
Gd1$Q�09r�����f�C�}'�,���2��%����;=3�g��u7$1#S��Z����?���)����U䓐�W+��-��K����nn'L��+�Uu�/0��ꔾ���Z�|j�����ۆ�);�7�v9��!�ϜF7[*��%́[B�K��)k��͎^0��dA>�&��)ht� �y�Z̧�����g�`jve$�0�G~�a�q�=�m6ڛ����g�׵߫Ӄ5��Lp��,	���R�B�\�4���d��䆥g�La�45Q�Yg�a�7}2�`;?�䪪�8��1�-���O�;U�W�~���ɩ�(�8���y+�BeqI�ӍX������Q� �&���?�c������b�2����rt�fv5%�6�A�R==�)��l�:����f3��H��J�v��%#��ݩWT�?�n���J	]x�~?klVG�c�d:��5��)�ۛK�e�0pӁ��J��X��x� �&Cd:�a�J@Z�t�MG=~����� /E`t?�;�xd;V��,m����f?�9�!c,3��S�Q��I����� @($�d& }��G4�k/����c����Y��mgY(2�:��|�J�c�E������H��N�����,^��
6�C�N��3�_��3�m���?�B��?"4Ȁ	܉:!�N�}<��^�j�9�.������i�&�Z�r�˪'���T����^�ye�% @V�k���|��Wۘ�
�p����~�~�CQ�Y�c�
�9}�������|��]>9��R�S�=\����N�"L�sD�����3/"��\n���0����<�l����5����3K
�!���[�SJ�zO���6z�lc�Lݵ($HDM�$ζ�"Zs�Ɋ4�+}���$���h�.P�P)w��2N�b��FQ����ra�@��r��
1&�Uĕ�f���MN�?#�"2τU��Kfh|�P��QN`���A�f����p)/��׿.�a��P�I���q6��
t�����07ȅ�c~=�L�[�{3^6B���	�O���L��@����lp��8ѫ�����A}��?�Ń}��m��$���^ {�'y1O���Q'���\P!$j<���!�7 {?m-�����0���Cy�lk�2�}���L,�H7�!�kP`��C����y�ɷ|��ێ��Æ@K)��}"�l��]3@��9�
l�*�<w��AR�mw�܄��3�I�
�h=ݢڨiC��O�P@̚t
`�C��j���W��vܷ���h������I,��� C~���P��Tș�;T����>q~���:lл�pe`� ���۬:e��8_Ikʷ4[�[`Hp�Wu�I����aM��``^S�ex��Ca�v͵�s�J�٣���f����A�p�����!:]��׮#�)�	�O��Ӷ���%�z,"�i0�N3��<�x����讇{�S���R	�O��(?�;׎5��e����9�W�+@��!��F�Y�*n�)�*� ��| � T���f�~��Az,���%	�di3��:��������x�RK�*�y��pA"�e���cv����7�D+Lt<Ri<��`-
��P`��c��!�~H�;�lkW�fκ��P��17������4�'��,(��y��Ępa�q��k��i����J�>�<�S�H���nPq�o��Oܲ�ɘ�֬�7�\�)��p�/	QerE�?��=Y�ߜ��F��hB�(�U;�X��F�?=9,���vc�\�]��KU��q툞eX��x�@�'q�j�c��Tu,�wq*�*="�@U�Qh�X���S�ۼ?���g��n�HM9B|'�)�s0d�8�c��"�l��F�}>��O o�=0��7z-�&^͇!Y��
�c�:R&�C��!�$k�j�;/L�L>F�), �c�&�����/�;	��C�!�u���l؟hv[�ƞ`����E��`��`z9��贏��3����"[��]�I~�=]�AΝ@��][��"C7���M�Y��%�yv����Jg_����� G�i��ـ�\W<a���'����$Z	y�.�o㙟	�6� _��>�Y4�G�6v��C�7p��%rI�<��,��9�Z�av�	�9�1�b����������s,
�}>�^�>��:�ӂ��"��.����i��0��+{#%�?o1+�o%��XZ��$C}���*b�	ph��_�Tqλ�ؐ�P�6G�0��:���֏�j|� ;2A�*�#V���9����$ti���&6�,ORAӔm]��9cVTK�N�k>�����z�,��qn��J��D�wg�K��SO1�z"
��}��0�p8�W����,��N�εS�8��F��EnvJ��L\cn�����Dw�P�F�00�\����d��E[�#Ŵ��\���b	W%����$�F}0�Ay���Mr|nAV�o����Gcw�6�3��!tx$]���*�(mFv�C"���H�G���g��fپT����s�Ig�����3�����ݱ���t_���/����nH12l#.k9����6`��s��}ŉ{K����;���ȋ�M�pZ?XJ���+����H���n���~���W���.����TC�I>b,U!c�4�OrȔ��g)z��yZa�*����lȌ;�mm&I��
�Y\�U��A\:c���|�b�ԓ��K(�*��6o�  ����6�k��˷=x���P��H��vR����҅�P�7�f���@��X#H[Q�H�EڟxKؤ���ԷD
+������<�͚(�e"B�@Q�6U��c
K�q@+�`0����ٺ2E�/a5n��� ����M��O�9?���?�}]�U���,�-�	�~�.
>�O4��XC��R	���P(�>�8����v�%_?Es2��5��u��������G���t�1a���Q�`l�`��π��bI,1�ߍ�d�7f���ف�c4m1�3����4���G�V��_����ZA}��Cg�<�hF ��8;�d���b��n�ȩ�U�}��e�lҡ2<�=Ȯ�c̐ �x����$���җw�@6�=c�QC�v��A*��څ�D5,�3��O>���'N<d(�#��H�&�Į��5��,bh�t��M8�G��'���j"��̪�){���T،�?|�c��Ħ�Q0>t<rx~(m��"���˝ʤw�頹��Z���tng���g�B�o�����7y�M�L��za��8��,��:����j$nF���d� Q���b��՝Ns4`˟��H�E��u���0[�sԨ.��k�`����|�2ד�U��Ō��y��Z@>���|f,�_;e�R@�����M����(���S�ȓS�s�/z���\˨���Ĥ�L����u9x����l���Q�ws�m�J����eg���y X�[jno��"�����ƭ-�yk(�f�*�,��dM���7WNoA�I�jK��A9���/�a���2���t8�8���#��<�H>�E�|�*�;N'Kok֡���nA�^��j�àvX^��B��!5���8Dμ$^=P�,�,��s �*���m��g��v�Y6 'F)��5ል��%B��u��E�	��6JS?.Nq�~�L5��f� UQ�:���4Ć�[��$×�"^Ɂ[�Fm��h(���R>?jw��|�0�I��ٟT�b:8�Y�9��M�X������U��r�P������++S��2Qc*�?o:a���r�<x�1�x�2�Xz�=�g-Gt���w��\���>�LkU���h�3��n��P&j`��9r4���;$����R����5���rz��!��-�A��'��t�WU���XE�wN�����oB�b���L�����4g����ݵf�}�P�G_��v����v�}�s�OW�����#T�8N���O���VX�	�K  �v�ґ���쑨@��-�n�� `�Z��a���^�F��}���o_1L����+F,�`�=^�cx�̕�0y���+`�,���/���U�1����ګ^\|��B)�h��<�h����yl���!����=�ޯy���BYV��K_�^�{�jm�iɼT�W����+�/�Q��"����9�4� �(�wҞ 7!�	���QHz�Qu�7�m�R|�g_�@$�WbǎjG��F��9	&�ߦ�Oq��z�
�)��c�����]+�"ԝ���*@X˷��eT|����;r�ʀ>�6���/NV��t��28O�!�_½za�񒡚�/�¼)���=�e
�\�T�J �I��y?$�Ƒ��]ŵ��ٯEY��~������LT|�K���C��Q���wc��?�˞�N�H	�ݩ%���-�O%a`B�^����F�ۣm$ߣ��Ck�E��T��X��E>'��YD�z-�$���`�I���\Q�F�[�7c������|�<�3X���yG�s�q�/̓����ԝ��~uP�go8��oz)��$��#�X�+��R1"[�v��傃)|��e@��fꩵ�2#���1��Ȼ���T�N���dBI�m �M�(|s���D�r�:�M�,W-(���8u�er@T8\��t,j��6��@4,
���p"QFl�+R�/fb���W0.ąo�DѾ�-}�1���o�TS���\���0?�XF����m�T�A�=�P��1�^?���|��_��i]�!��O] >���PNrN oi um]����"�2�6��T����S�]�]�H��>��4��xP�cD9@6@�(���qUĹ�%�2���\A�W�����.ӲR���g�qT�G�L��:�)čP�t��7��
���kRE���� ў˭���5�����Þ����G@��V�PRs������p|G&��)�TM�5��mO��>QC7��`�B�4�G��}��E�����B��1wV$�Y\z����_�=�e1��	�5�ЀuX!�,7�h���6��]�s�u�j�qKj.�"��5g�ڃƟ��T��E�c�1G��c�0�P-+��f��`��cl���e�nlO�<,<�Oу��c��^2�>���a��ҥ<���=Ñ�K!�7͔֒@�͆����5-�u^���/+��(]b�7v�N_R <�w6�T�i19k���$ё��ϙ��<S~�� �1����m�!8<N��zy�Ez�= ����FM��X��ޢ�5��rZO�Z�Z'�9gX�9)�B~�f�03���[m�z���8�H9��?"f8�Tr��f��S$����rͮ=��2@���������R�2\���Hy�2��
%���dJ;���=��z��Cc�E�^��1���䞍���A͒��&uŗg_V�o��	�h��"�![S�%%��;�tJ��k���^[�s~��؀�F��́-nU���p�z�����ׄ3�s�b\tN��|�O���m�\5b�H�p�=��1��DIo�<�Q�FĪ��'�A���<�����q�ϴ�SnP#	פh�����O��hZ+q;�[���}t����G�P�fXS�l ��u<�{��#ѻ &3��_fM�M*$>v̉tI�Q�%v\�^z4yu6fS�?.b�ICSֳv]��}՝�+lY�ӳ#���W��%[�KP����"��K�%}�BVX0q��teΎ�����X!���p����G��
JP��.77
#�g�u���䨶�e"�����0͉�4iCա@������\�gf����][�i4R�G�c��^��`��J�S�\.���6��ԟ���z�H��+0�����c��B��9(�ML�8/��k���D?(��WƝ[��=`��x�d�pb��T*{�?h^pu�*q�����<&�z ������EW
KR�� EQ8g@��|��T6�`0Ť�IB΢�?����Vb�����rl�C���
�&�	] _9)6��`KBf<�H�@ْx�&��Sboo��ޤ���"�Ŗ)����%��-'r��W�@�*uM��Q븿���kD� n�e¬��!�$��/0�Ļ��zF@���_~��Ji'�����h�2��x*����#�@�<̿!w]`���>�yU��`n+ 7�/S�[�Bi�.ӱ}�$N�V�R��f�����ǟb�;���
���>n�eY�N<C�!pa�8���M�}��43ـ�j�CU��ѾG�P�@���#?P�E�v5�	6��&�����-?~�[W�@�y����Ͷ}������*�'G0�.��w/}E�����ڢ��/�Y޶DѶ�騢��X�ڲ)���Z��\g�<�|'� �4]�����}
��r炓]�V-,hJR9����S�TR�"�v���t���c^0�*�E�ְ7Zp���U�d�\��=���t�,�$�L<Q� �H�݉��~�B�%f�I*��:�N��K�ٻ�M��=*���dΑZ��.
�hsf/PD��VE���a.�����������vK)GA���w��Y��&L�����ۯ� ��uq,2,�s�A��fy�{��1��G6q�Y����ESz�9�Cm3u�n�Q�_P�W�^,w�����Ac���m�F'�0�~�,׋҈T�Pb6��M;�>�l���
^6��+�92"B��cv��>��eN��3��K�&�N�U�"9W��`�޺����V�Z���;�ڎjyL$�s�^��!�Ctŧ�:���C�-��ռ�:S.���2c��k��ů�����2��&L��vR�]�5i/�5"��4���K&�X@�������<&�]M���eѿ����M4K^��B0
�Q��jm&���_%��������X��kqѽ����M��	Z��H��8$7� �b��1�JA\^����Sc���W� ���qfz�ѐ�پ�!�I���-A��VQC�rBIz��50���iZr�g�Cr�~`t�ۥdG{��ܗ������vDx+y����>����m"�ܿ�ȋ�HF@���Y��{�3�E�'�NS����R���*'H-��}����TY#��N֐A�{����6t��,�����$�B,�HI�~����a�ʏF�҇�,}�I��u�6�g]���̗�����Ur=����z��i�٤}"�t���ZzF��7@��=r1�
���E���ծBD��>�a�iv���)&���sj��'�'u��~�c7���n]��I�
k��_XEM�恊����a^�i�[Ӧ�~ε�.J^�@뛇no-8x�E0h�[
t���.򛔋A+��Vv>�'�aJdmu����-aP�t1�GU��I����\dU�d���ȥn�rg�����S\k��M��O�]`�1fF�㏽Jbʌ���}.��/�yj?pp�����t�Ѣ�����|.9�����og�`�� �.�"��y:�����[��HC��k=�-k�A����Z��'s�sS��k���*5�[(
���r�ە��#�9����]ؓ0Њ��Nx]ɅsD&>r��tU�-΁Z��¾��BV�H���4�6�_q�;�| ҊX��P
��(udq���F�٢z�a^����'S��YF:W�獳�
kʐ�
R�[Q%�=1��2�] �����'�"�"��<��}��0%���h�')�H�V�i���?�o|�n��-���#�
S�I	i�`�aJ�C�},��Y�xt��6%���t+ֳ�x�D1�����'ȁ�G��N@9Kg[0=���h���yZ��*�)mM�|&��1o�d����_9L.�g��_%�;+K�-�9���p_4g������P��: ��'n}X�������O�y,s��ݺt:we�Oc(�L.k+���6��2�1]�;A9��RLbjܝ�M:Fe)���7�^�h<�mcQ��li�4�M�âm�n/6���1����$���FƢ���]�Ӭ�7��8	�P�D���<�jm�!����{'0e<��fA?!0���Y0S��oq���|��l%t"�l?@��U�BL����(?r��3J�[p�H�Dz0x����h���X���A)o0ƞ=L�S��c	�Fa��d�^X���Ѡ�yR�~��W�xe	s1����0������z��C�}�px�>�/ޮsW�WV�`��l��1v,
�"��Ucw�mW�<��q6X^��8XCD��R�[�\F����[���/�B�a�8	E� w���3�b#��7:��sY�e|�J�,(H�`�	�ϩ�����<�)�����dR�&	��"����62w�!
�J^Ԭ?U&�fz;l�?P�'P���O*�������4ҍ#���|D����	U�_��]�#I&P��}���*QF�3τ�?��b�e|�{!)s�Fr�E�\�����qؘ1@�[��3q�$�I���
�l���&���� _#o!����.���d�L�Z�lV5��@�Ү\�wS�R����@7r���N�/8�`��wE�5�+Ӝ��(�o��H�o�K�r$�a�ﷵ������R�hZg�r�v���p	��{uD��٬(w�0�>{�@��B�}�J���T���Un���c�Z�� �(du�o�Ky�p3&��2d��[���%�(��V�Y�
i?,婡��x���g*93��G�S[�#RC��Rw�����_�QP4;4�r��?�3tY���i��e�yy~�����H�?�ƌ[=�"��������ߴ���)��k�o/���d�C��BF_�nHn�)�վ-y�X��Q �b 9%#���<5���N�J�|o����H�
���7��/!ɫ
�5Vޜ����_� ��y�E��)��Z���CaT��o�0�+�����*���,�fK���&)}��� ��G�{�JW�ǖ�-|�O����sS�G���p32��4�)Z	ma15����w.KW�z9p��~��̩*���Q����;���A���ǹŭ�1 ��P�z��~��(6�l,]O��C1e6�ܪDn�<"�FN�iML�K�P��6���������Q��I�N:��B�	y�gR�q�#>9X�����q�,�g��w�7��1Y��JDv	��q�
&nCl�����*M1�7���ߪg�蓞�� 90�)T�F?lHU�i�AQn���A(+���i��s����9;	"3��r��o��� 0�bp�fg[��Ye�̟��<Gpq�%����3EzFYq�gj
�!:�OG���t�n���g\�j:�Z-G�]d�x���0!�}�߄Y�M�~�uc��ϊ��Ǒ��x���|b�ȅ�4����;�b��L�"�)l�z���}x�e]��r��6 �#o�%�
��!��0��01z�_�]DrƸj�F�HNTwa�M����Ȧ�FS�ΆM�@v��:'գW��%�,�ۊ�����Y�O�Qr"ATo�A�&]��"���2;Xv����t:��5���� �n�w7�x��H���<�%,��#���Z�`Q9+���oK�n+%�z���S]��~o��o�6��۠o�r2��S������-LGo�V߁���٧�l����f:o=���;�s]�<�����%M|=��Z��: IK�c����� l�y,� �e(�4�f�GJ�7k;.-���=��[-�35M ��睜v�Ř�}��F�=b�l�#u�����x@7�@�1B��\[^�~Tj���.:��C/��ۚHc_|i3�M�~��Ku*ȴ �͎R}:��t6���P�7�٫"����"b��vG���U7/��'��/�->`͐ �f1<����!��D�L��Z@=/{ǎ��uS���Mf #�b�z���谧R>nU9��R'���sT:��R��[ZF�E��`��� ��r��'�ȡPb��%,�o��/^V���:&��r�#��a3)�"ƲO[$�B>���*B��hO����{,� �Iӱ��.)U��X���X��k)UH��jg >1�{��C�r~��G~�����1�T$s�4x~&ʀ�rzj�����}�ڢ����1���d��U���gmh;ʖ�� Ce=)<x�,ǹ�����C��Y���'e��+}�����ә-T%�����Z4د)~�S����![���q:��|��~&X��.؁V���kwY�1̜3���:x|�9;O�W�"�����s�CN��o��ޫR�^��?���K�?���Em��s#@{'��V��ŢFw�z�q�0������w�ߙ��j�;x o�Գ�X��7�&��Q��vl���[��ߎ�K7��a��t�����E@>y�MIn0�	F���o�(�����}�AoET �NQ��y���u8'gꥏL���b��%�TY�@d��� �L�́��us�v+\](|��]/�ע��̆9۬����${k���x�є�Ok�~�]���-���,�b�%Fv8���e���(���ZV8����VJ��A�*맶v��ݦ����$r^����Fוb�"%�GԎI�o��*
�:��˲w��t��ܡW_V_��V�u\i�#��k!(�Kjkv^����%�v� ����^�:ۄ�2ܪ��РV�)�FbKL�%h�5���`���2܋QT���xXL58r�,.��n��C����r͛ho�gE��*�S��#�b��2/��ؗ���8h,L՚FX��QD�K�ϑv�h��.�����@�z�,�WNҌ��k�͖w�
��ytD⥼wi�HO���:�9w:�9�������b�NΒ2���3((�r���ț���=���H[�8P��p�8��x�.e��j���G;0-�O�GV?  \7�P���7a~iׅ��
go�Rh�E� צ$�+�0&���ЌX��WMn� ��'�1"^ʪ�.�{�ϴ4]�
�.%�,]lo ܅�� 	�W̔������Zn>�>�E,������8�%�R�E<��"	���&�ƅ�\��$j-�g�BGh�d�TcC��8e}�����Pz_�2#�����$_r$�?�m�Y~�ῥ�N��Z����.W�ܞV�#�]@�A刢�	�j�ie�>D#fnJ���r$"�̊]/���J|��������c���}Ќ� �M)�H�	�{��F����"Iք��a>��;����sYR-R�G��b�>I����zP�s�[���w� �.X%C��-���'Li��ikY���<n̲��Q~�s9�0.�ޑ;���
������WMr6t���>�`%8�je�KD�]6�I��׿�ymᏑ�c�3����{]�dY��rk����kώU[��d�%�}��Њɾ�ޤ�(x!�����vv��4�!�R�d��,��5�Vơ��$ʛ����̈'i�z/�$��6<�TL��/�f��7��s�
ʱ7������ʾ��AA��TDPq;��j�;ڧ4|�7�B+��EU�e,h$�����B�t�iƙd"dd � ��*� f���)+Ne]/�r~:��f����8IBa��Y��"4�^V.�@f��)$SƲOm;Q��"exB��!�p�&�2g�e�����[��į�.p��Ei<�!�,�'0������8��ЀTc9}gi<��p�f�N� 'p��ȁ5�G�:��,VJh���ܝ�Fz ��-�Z���R�5�D�3M0�7V���f��?�03$ϘW�&K���q���6�Mh�Џ����ts7�I�~[��<:�i��)�]��w��k��,2��.����D�\ҍ?�nL�@��aY[>��?�X�E.�+���v�b��B�s��go������<��ԗ*�s��{7��������}�-ұ���8;��EU]�%��x~7�RBc\K�����ގ�D>:k�h�vȘ��mZz�Ep	�J%f<�6�D�S�J�d��
W�r��g���q��Aأ��8Hp[2,�#�`�5H�«B
SLT~E��P;�5� a#���ѡD^�cn,]�� P��I�5����S���6i���|r���[|�[t6MOi�LȚ;\�{7$j0P�~��#��~ik�7�j~�'t����ni��u�F����m`���Gk���a�g7�iF�:�N3���B�25�Ґ�0Rt��8'����bS	�YJ���̶��z�D8�:�[�o@{�J)��F�׈#�$�|W��ה���.�'���^�i�Qg��j�^a��u�^�����Ӓ�¯o��������,�`�LE�7�?}=���W��>�{B�/�2��O�4�F�y����7����r(m�?�Q/�].��'k�B ��i@W��Af�
W�� 8�ߵW�i�W�X��j-G�;"`G�q$�t�V*[�f��� �F�#�k ôϧTӻ���U���n?��W�E���~�
����^�Co�ǉ��9�%�jʍ�]�PJ)���RXʶ�{G��[�f��E�־P7������_c�R�]��������n`��nv�lѻ�XX�i��O$(e��2v/�b�g�Q�>b�Z[��K@^����w�+�,zu�u��[� ���W�.�Z��2���E Zq���Ϲ��K��P5i�i�%fT]����E�]�&��?��<����O�Ş��3�(�}sGus�cު�v;ޑ���I�r"��r�L�ň+���
C���,�RG��H�t-u<��q=IJn|�r�8F���E��U�qmzĴ�q-Ҙ(�u�+�x���<{�����"Kf�qθx��y��Հ���(hVfe�K�0F�~&$Z����Y#��tǛ�r�PK�w$AMZS�k�h�v$x�b�ΧT��R�Ԉ�i
��osP����g&Xԥ�Gh^�s��$1��D��Ax֫E��݉\{͕�r�����iV3�0�P?�hpt?��u�S�G�D��U�m��Uc�i3
��r}t~��Hո�)�LR����:���D���+3�C	��/���<�X&�^۷,�a���l�
��ؼFL��E�����Tߕ�1��X��h�T߬��o|@P�gF5�?�ꦤ+o�������CL��;a"Æ���g�H�W/_Xc��h�#[�/�N	�jK4dk�p@J:ާOD9`���9�I�T�)<e٪��S��������[AB�lZ�:���Uy���H�~QL��҂bW�§�6j#L�-9�~ہR���6��
=���E^`�i�ۍo��my��Ȣ}�-o��<T�g	�#�x�Tf&ئ�d(�W�};��p�1{�Lz�}ܨ1Y#~ڤ�[��*�E�[��/Z���c���6�J5?
� ��D�59$�1�m^�XX�FގB��$�Xa�9�-��(<n�?}�l,��_ ��1;�4����>�O��>jP�9��|+�����8�e�P�"����3b�X�/���k�T-W�b/�����'�h\x����YA� �:(�+UBj��@�	�2���"�͑�H�.�Sz�����,��d�UtV?��$��򫗵�\q�u��4U�v.h,GY\�hs��g@Bl
e�(E�$f0��T�[7 's�e�y&����幂 �^)�Q��p+�C% @��l䐝nھ��
��s6�ϙJ�U�LV�����/��$���ښ�O��K�|�B'k�ߴ�C����-gs3��cO�i�����&��n��!5w��&|���n�������_�A)����a�2��0]>���3g��{TP�ܸ^�3��e@�8x��b�iHo���D����żr���VS��ѳ1��MΑ{LT`�	��w��V�/��B��^Ң�=�Xe�Y����Q��s�R��'�%�YR�V3G�딝���sj'�����	k�e�>Z}� �挩���!�8����H�憎�O�A��Qq�:�R
����R����}�ԩ��X��M?�5~m�
�2�kN�DG��!�!U�B.�B眲�/r֍&X���T=ۍԼuA��d�{&��V o�⬷]���5�Jm1��j�¼Mff첷� ָGM�v�ؙ`����x2�j�\��n,�Oj����2z�Z/�xx��:�蹏�z�:Nw�*S+�ԄduS�C_�K4u�P&�.�~P�z���?���ml��FO��:��;��m3��pq��T|F���!$qrU�f�&���pO_tw޻�,F2[����W�bXP"��Ҕ�j~���D�8�,닃M2��k��;��A�Dj��8�sP+�~tV/@ѫ�v.�������t�/u;�7���VtOu���jq�yB���w�Z�7�1�Y���*��-��H��h�yeO n "�T��+�q��WJ���O�܀I����fiF�J�I��W�k�q�o#��UD������~mK$F�h����,S�(z���/@}��<�2F�O��T��9U�a�W���OH#�*7��w�'�$f�&�ct�Ǯx��gӼM\�o.�'�?[;$���@�c�D����M��[�<��v��Z1<CP�fB�/���?C2}�QD2�i�>����6=��%Tb��eafջ=���������"{�s��LRM�"ҹ�k�;�8��~�/�����}��3Z:3[����B=�ss3���)a���)�5��w0#q�&Ba�s ��hz�O��(]b�쿣� �I-�k*Q�-ז��w��㨼|�b��N,e�� :�al�D���O&_Ν�C�2{�w�&�P���s�K���E��3��g�{>vz'��R,���[3���d��Lݲ��-� C�V�*�)� �a��?SŎ5��Z�������B��ݢA\8,Q8Q��۠�����2:g-�[Gf>�w�-c����3a�:��򝜏���R�*�H�7i����H����q�xW�+Zz����J��1e�-��l�4�[pC���N9�@ @�7�i%"���D�q��9d D������%2K+��n�m��h�v�`^`�E"���R�0�,|��3�o�|���^�e?��������v���3T+����)��E2����$5��kF�ˎ��Lf����(}��� ~]���d)��^'nO�	�MY����dYT�-,P'_�����1v�t�Qa�KQ�J���<Q���2<i�v?��
��C]�;�7͕��ޒ#)���a`M��7��)9x��f�N��yT���v�\�aR:�0�͟G���c�r�>r�Z�. &'���K�(ೣ��*֒�`a�D�F<��Cn�aB>����<��pF,�z�6���'�O�\�!�8|��樧F���'E�k�B`4��U��'j�<=l��0��V�"\d�)�ybk��pib5�Qr�rh�\��-��Vp?A�$yI���:�9�8C˲��X�b��{��dDLJ
KB�G\)e�-��-��g����)w�F7�K��M�YX�S�F]��I�@�O�<�N����۝���Q��ϙ�6�~� �뼘.�g���i	�캫��66�"�muR{XWC	���7�%SJFhR�!����b[.~K�S���3Oc�C�|���P�k����X��ϯ�N}���kt�Gkh��	�$5�3�:T`�}��8�,i�ט��X����������!�g5���7_�,��;]�u�5n#���0���U��b�,�����J(��z���iS�+�)��t|FC�.[���R�����o'���Cj彧�2
���C(L��-���m��h��[�G��k�U0z��3��h1H�S5bȻf�%�����P�٬�T����#�W7o�_��tAΟ�^�P[E���+%����%dMG�:����/�a���4 ���z�!q��x�鏭s�P��S �a�9V^8NQ�#t���F���3�o�B-?�O*�]�
+�N+FM��i̯���&�Um�i�*��.ʇx�_S"���8>��ǟ���H�r}�R�X�r2�Qੜ��"�)F �&-�e�a?�7]�e���n�f*���8��m�ݘW>����b��7�Ϳy�y�+�M��!�Xd��4��4}���z"���sS+g��I�@�ߒ��~�_e;�]A���_ ���Ƚ�RB�/�^��@��K��_!��dJy��qP�z���T��"zD�wS<�A '=�6ZM�K���"\ �xv����.+<u���:q�����2�*�7�d��g�� |����6�x�G葈���˅�ox�Z2e��� |9������CF��,��Ev0:\�1!�v%-S@�l�q.�[H�D־�+�&#A�9����11��2���.����Ϡ,��7��V��n���I��2�����$:B����T��$�(�nL�\d}� �br�y��ˣ�[y��a�,�������P$��UP#�F�(����j9߄�E6A��[�b�V+���|8J�7�z��G$)/XL)�� }3�H_4�q���_''��/y^�q���F.������3���]��(��~�#������������J��s�M�7�_� �2�T����2^d���cƘ:�:�*��i��Q�ʬJ-_M�O���*�/��^j�X,CIw�QWi7lf&9�Ζ����0.�X�=l}�ER�O���d�{`�LZ���Ɇ�wy� �w$�uKx̑�c���=���&��v���X��"��W����@)o2580 
}���9ڔ_%�^��ʽ²������>�V�:���`s��qVW}���P���z����&�$b�fyEr��}D��)5�����nd����|\���)/n� �eHic�5 ����xQ�`��b�a�^��0=�)�`�����g���jQ�ݩ�}B�˼Q��B���?�0Z1l[�B��s��܍dҘ�?��RԜ�w\�ljq�ʸ4����Yn�<�TEf���g��� �+��Wܣ�o��ݞ����(	��1=����h�g$�ks�rC3��Ad����T�>�&g$�W���2�Hp�Hk�.@vk�4|�z��.�Er6�e)&2	��j¯��c"�kT��0�����I��(G�S�c*M�O��D�ն6z;�$s��@��c/�& &�w���kt/����}�p���U�����-�&Zb��Ӹ�_~QN�X�� �~_Q>ޏ$B+L��#�l�Pk��[�]ꭣ`�,�ӫN��
�t�(�9�"������ib�������;���)��Y���[��r3&ހ������d�i�q7��t1�Ks+���4����cn#e��ʚ�Ԇy�����`xc�p���Actӹ6����wL)E��D.(v�I-����T��K����wZ�K������>��c�~f���1����a�q!8Lm��&$!�4���tjy$�T̵*ڍ�����P�ua����y�U��_4��xbÀ^��؜��=ʶ�O���@<�n�B�-��n%��O��m���\}\��R����2;�6���y�$�s�A��A��C����Ϧ��G��?d��=�h��_$�#��J�e,`��b�(e���3p.��$umy�@n��\���܇d��ɭ�������N p�ב}�>rX'���U�ʝ�JH�d�򉱰EZtA�.���%a����K�t�9
���A��<dS�N������V���(�{���U�'�����~�yѥzyl�ه������Z�LE�F�|Os�by�A���c��@r�2�m���H����Xۍ*I��r��EY��p�m�'P7��I�� E�l3�sĻϒʹ��t��X�La��ӄ��T���N;9�V\J�	�
�s����{ՠ6��0��2ذ%$��k�k�L:!����>�#oz�!�~����%��-�x�8\Py�06̅�!�\k��a�jg6Fl�(+Zy6H�n�x���e�^�Pp�R�΋�!冷ݖߑ��ŏ�QM��K]]b�9b겭
%�Zze~Ŗj$٘F�Y٣�)��<�#DOK��`��EN��I�[��$�Y,�;֊F�o/ѵ괌�p#9�W 窌П��.췐٪�a�5œ�G~����ad�t7�AY7�e��Y^����Qq �5�*�n��_��B\5�T�h��x��(��X��$�Z�fd�:�Q�ݰC�����S!�*N�	h�π�˔�?��scm+�!��H��d���hky ����k��m9�u>r���4���σg���as���W��I�7�^�d/+����j���#g"��.����[�Taʷ�p���k~q��M��Ѹ�@�4\K�j����/#u��r�,�〵��8�A��n[U֋e~A>k@�y,K]�Ɇ�K��؟����T9tB!�y�Pp?8D�K,����[���U!|���&'�}��-$t���"w�;�2�M�)��X�7���?ʝ�3����#}P��Y�,��`��7?���Zhz�Ģ=�k��b	ܑ[u[�r��L�_|�� ��/J�r���$�s�������\�A�9����{��L���L��--��l+	}�JX}�l-rE%�׃
f��|�;��r�u�~Z���P���jv՛	\�{�}�����̥^繛�9�e�K�8�ǌ�#�{t�{��cW��a����Z��E����hV��p�=߀�i���Y1+�d@Y][�W��p�l�4\ʫIOb��VY�UU��V�#�Օ� =1���u�$,��:�w�<̇�@��B˨�� ���4f��g�+��1����dNM������R����ٽ��t}��u��}�ӱ�a�⑇���X��f-� L�&������eіk�2΀�7��,Z�Ku��l��S�]䱊M����IF�7��Xg��� 嚄?���I�:��ӭ��=�THc���݂���<̑q��th�$���~�� a���ע0��@hi���nj��,P�lҚܼ�Z2�)��V(�1�b���Z�����Z]͙Yw��:)��w��W��~���^�� ��܆�g��
4y֥$Cs�"yܐߛ)�-�s��؉�
��T�&���<�XZ$��/]S����v]P�|L[MaL_��ࠔS�d,�+�}�g�˔tQ����t�:S���P���!ӝ�a;� oK���O�_ɞ�-3J���m���v�5�[�;6�+�G&M�-�!�/x���L���9^�ҭh}i�YZ4OQ�n:Q��&l���7ƫ����ӹ�93J��(�")?9��o��,�Z������������z�kN����A̚K�%b"����4H����H�O88eXtv�vCy�����]�n��;���t�Zf���y�ם��7��Nm����{�t)�ֺ������s�	c,�;,�(v�)�]٥��PFͼM�Zg#�W0��ҟ��\�(��b��e�n�*��fݗ+�����%Ƕ��><lE	�u�+��z$z�(��`oX�x�U=bK�e��~�a!���; )v֕�区��S�}�E��J��~�43���*�:<�3u�%�N{���W�j�ޏ��#�+2°�;76x�qw����)Q�(+D�"��h�b�,F��q�W�^e�g�q0jj�Tp�
�I�$��[Q�F53��N�|��B��y�WTi+3	�U��!�∹�rh�{�v��(�X�{(Q{���^���K��f��m�������s�j׃��� �Q�TOE�Q��?KS���`X�Z(r���x�m�w�Jې/����EZ�L��K�'==�ԑFj$�邻�e,R�\y�hT!������㼼P��)�c�N��ͭ��ĺ���@�>2S��M�� o���Cl�$�t����̚���R�����my��O�_N3�;��_����>R-"ޅXm�_ϧ-!�\|;���5^nu�#rFc2��y��Y�������R��q���G�����'�0�G8�`�S��=������:gk���i���i�
�N�8�܆��'���fi�N% -ݖs9�L�OB��`&�D��(6�BB����j(��v98n#�g#���.e#�S۟�[O���#�mN͒S��t�'�O�
+����G�ZWZ��R�!�'&:�"�QE$��NF<3�[��!'��i*�9<�=0lL)م6�
M�TPc��z_����]���@��5�7 �Z����+�S��g�Ù>��}�����x��plۘ�E�ݨ,�F�_H�v3�KV͵p
img��x�F�S*W�n3Ƕ�?t"%U��v�8Z� ���X7�MQ|��i>1q��ѐ9B��{>�RΓ�Z�`�z�]��&a��:���}[�a���`�ឯuߘ�7�`�}���c;�
����dKw++��+h�?��f�ϾW�Od�]sƷ6*���
5��~VYo*�����s�?����n;1u>s��Z��3����#�0�1ӂ�Bi����̢I������s�ǁZ�X 	��PI'��[�-Y�HP���M��I�`_K;E��%K��d���IJu�?�����,���%�ľ1�_�y�I���Q6v{O�,x�����$)�^�&U֮򢙴����V<P���x0>(=���HX(�1�/GJ�[��}	^���n���j�u���v
B����'�]���B�r�͹�t��TBh1W�!iGK���Z��ݶ�W����oBb<��^cG:��Yʹ�2>h���l�0��
�a�)rU�M@z��g2RXųT���tar��~��+w$��-!>�d����
��2)�Y�9���J6� v��N<��M|�ۨ^Y�R���A�u�������P�f�����4���|�f���,��i�C��xf����xZ\�$��/رˬ��x,��qN*,ކ#�*v@[�>r�W-fk["���*ӷ�/δϲ�E񜗊iH��7��ɟ��ٴ��x!�
 �z2i!�;��4�ںF�D��JX��f������zK��7��1�l�WXP��0��� d���AU�w��k��w1+��e>�;��u����Q{�\��f�j���0�);��4�$뭌��<��b|�X�Y�{
^g����^
SPf��9�D��7��5�FCk[s}��h��BRd�����c`^�9#��[�Fn"�5H�O�M�
v�¬sԋ���ﬨ��y
rD��P�u������Jx��2����RF?���/z�ύ��]�F���I(��K9����(��p吡���S�3Kϑ����LӲCf�b�BM��v{��4��E])�%ы�?}e,���u"���$gEB�B^2|\%��������}�U>c,f{��!r{4FT||=��t����HH�+#��wc{���F��TFچ9̈́���	���R���_��ld�����g���}�kv��q�zoh�1��4��R2k�d�W⎆�l�ݏЉ��-�Qu�պ\�\Ep�t����7�[*�F��&3���e�U�����qZ �pN[;�$��thN�_� �V�;�
�ݷ�����å#�U�;���TaPk���.����LSОR��]�y.��>M�|�LSU9��h�6c��K}��E!�i,J�z����C��۶r�{��{�ϲ�"�K��Ш]�Y�q�Y혣5��0}��9ߏ˓��[|�ѾU+�TZ7���ᩕ��a
����[oF,�H�̭����n�u@|CdX::p��
�)ʵł,�4U����E[��#����g�')�^d��ӻ1W���&��޺�9��♊~�gKo[��
"&�G%�e�%�"e-��B�r��M���Cs�b��YP{�N���v�Jއ����-:��~�6Q�&*���3�7!+�U$���gY��@C�_`f8�I��|�r�8b�m�}�65��zv�ZBJPX�s�`/*���	Y�.i5+��O�k�q̀�v@2D�����o��Gw�B��<c�~ۻ�	,�=�<�hQ��B�5�ۨ�̘X��&�
9����5t��;Ѡ���0����YMh�H��$��⓿�(��Hq�����A���w7���6�x��\	"-0�S{s�D���G�9�1[�7��K�Qi��j74!�~�������V�����Ǝ��Ef롯c��r�S8�� &FB/$��x�lnT���Ƕ��'�A@���N��06�❦�Z�HWX�xM0��k�����������,���Z���y�C�8-���OA٣�
�_��⸁�WU~�rZǰ��n�V*UE�����$�!R�D��I���U����w���	7�3�^?��EdN���;��{�w�ޛ_�«��S��<G!���
�2��R����q%9Cf���{��W��ϕ�o��%�Q�B��aX�I�5���r'��#���
�X)F�&�ڙG�����W��%�R�N�ɜ�J��'�t�a6#$I�M�p[Gyo�ϰIyL6i"�bsf4�ww�>��-�Ϡ;�y�hW��P�����HH�&���c��
m���0�+%,��ޙ���
�1�5kT52lw����# ��~���d�f�b��-c���]gS~��}˳�(=l=+t²�-f�T�)Ӯ@V��sD�\���S�P��o5�����D�S��[���ٗ�jRA�]lȯ��Ox����u���"�Z�q���P�s�E5'�����q�4���z��PM�<*�iJv�t�S�
��]��0�����xQq)�#���&[�㕻��/=lL]���c��}�3������R��Y�`�mk��Ӡr�s���H#<�5a���<���zR�����+G���؞A�,RJ0|��¤����bђ�D�������n��MrP�ݛ`����o��Ȼ��P:<�}) A��2BPې��
,��D�Z�j��3�
�@KB��Ov�b]��z���1t%_2���p(P�䫃`����}�Z�*�Ux�pUY������h�`���WC!���� '��������W�+�й8��P}� &��[;�2�R.#кA�4�#�OQ��\eF�=��y�������┙8}Jd;�O����y���T����a����Hv�L��Hj���kBm%����4b�;�� �;���ލ�k�^�����b�0�j��@jt��Q�#�go�17\�Al翗X�H�@��F��%5���j>��*���^K�Kz�d�-";�1-;x�#� �Ȕ���D�p�Hk'�l��}\�F��ZI������<gE���.�]�Ng�vw��x7�#�B��ЩM.NSMX3B��~]�u���U�~o��ԇ�K���!d$��o�n߬s��6h�iEz�#>2��2nݜ�o� ������Ǫ�i��2�I&'�3@�Y�,�|6�"+!1�c9�v4!.ݏ�K��5u�1u.hA;�$�yF�n��"�b��Y��������%�F�!=6���Sz���9
��h���1����!�ԕ����
���dM�T�������"�-�9���C��~d�H^kUP��F�L$�$F�ii�^ڳcf��"���ҫ82��K�����7v@*��PU����ɇ~�HP�_%�D��V�͈���%#Ɂ A�=�"w�)p���э�b���6�Ijq�`��#UMQ,���B�}Q�������*UT���%�<n�Jk69��!�H�vh�d�=������|d�[��`������{9��64Gʗr�s�4������d�^raӅP ԍ�8�[�m�"���p��zC�4)�~���
:a���Pd�$�sៅ"�b��x��	�>q*�`p��>��B��|�S���wcS/���kU"F[)E��]h�*�*Y�	Mu�J��^�Ўa�8�d����0w^�w�ye}���m�����X,]P�a�4��l\ƪ-��L:U�[��($�2�_W�s=1b��,�M��"X5�R��*E��k1㸎}���)�1�ELF�ߟ��y4; ~=n����q��_�	ç-((&�߲[?�k'd���/�bS�EʳH_ܶ7X��oc�n8��@ݬc��&�i�3�v�����&�X�Ma+�a��	 ;�[ϗ42.GF��ƛ�6�\���k�S!����-�'=�*-L �V
��6lo2K���h9 �g'��x�HD�?��!Lh�)l.�tn^�]��q�p(�P3�gx���s�m�*�����1EFY��*�d+F��*����L�BL��?�@`+%	�p�lĸ�N���/�]�6@ؼ�V��埅�Q�X�<ZU���`�4(L�k��-b�޴�Y��o\ *�jE��s�nZD�o'�_X��v+���\?���H�����������%S������ǽ!�9� �K�m/��|bj[%)���y]H��0~�{����s�k3��*Z� ��FC�jF���q[B��'ƺm�ў#�]�37�L/'KK�R6\�_��.>���G��&)�J.i��y$�����Ё�dW/Pycl$ނG�3�Wo�hF;����ao�ge>:r�&L�����jһ`"�ř Fm�����У��k��ޔ��hB���u��ʙLL4�-�����S�Zf#��4pW^��56�ts3��8o��N�k���a��@�%O^^�L�
��K3����P�U��V��7���1�p�6�R�&�Nې��sU��Rd���mu��Y�7��L���'�6O.�S��]��5���׵P���70�zX�3s&#iCF;��d¹��U�C��$_��>��t���ʠ]�`<UA�Q$��Q��1�1�mTb�
���j版�Z-�L��8Jw{ڞb��2�)�bs�c�G��M�$z�#)�7��!W?�7�7�v7�S]QRG�!�X�!TP���}t�Âg�\>)M�k/��5�� ���=0��7��5��њ���vl?�\��v�+3�z������Ǐ��K-@`��[��V̙5T���n,}FÚ��G�фt_T&�V(�p0Aˌ�)�$Y��;@G^z�D���%aCm�E�G(�<��s�0rD���l����KPr��`y�uA���˲i�3�![��ty2�x���z��c��_|�O�2�*�=���C=~�ǵM�eVN�,����]b�"�Q>��Ar�s&����U߶��;K���e!���Z"���eo���.x��hyP̵0�)��/(��w�j�ȵ�Su2.�P��.6H���$2�{!�����aM7��rk�$�UTvZ��e���Z+��3H���^�|7��})�|U��t����y�%ˏ�������v�>R�E�e4%ӛ0O������z� V����ןh���C����)��G�e�zx��BRf�	������	7~��&��3�Oأ���z��5���E�D?�W%D�/m�$�F�SC��Q@��Lf���C8�!Nk�����ލp�,n��#h��j�z
��O�K ���IU�'S��H7I�")�}dL�ǯ�j��Sj]�uܠ�񝮄&�W�����q8˦�s�L�J��������	�yK"I�F�쳟�o!��7��k�����PRMgڂ�dpB�$���S�m�%| �^Ϯ�pC&4O��Zƕ,^�m��s�V=�MK2�P�{�%wiF��Q��3��y�QJ��偆����m�`m��X.�GV����Q�\�V��>���/�8d8�Ѷ�4W勲����04��`��bӾ��10�Py�+��0O~j"�����jE����J�o� ��)Ƃ/C�+�h�0:f8*�͇zQ���)`�b�����e����ڡ�h�(�P�� ��ѕ+7��j�d�S�a��AB@�.[]����a�;L*ʁ���Q�*N�h�_��j�B�.��<>aq.�'�\�����M=e#pM#�z�W8��a:V�8t���2$����hX����؆kiԧP�pZ��"����i��t-\�m(^����.��Q$R���¥�=�kW�ʳ�� �����$�9�Z�[�(j�Vn��T*w}���4NnL�&x�1�#��.^�@G�) ���T��������/YI�Gl	�޻�ܩ�18m�Q��PH�-H�%�d�����L�7I���F<�D�Z_ �ee�(���DYA��wRK��ЇP*��*��-�y���!�FR�Weͦ�yQ��L�����
�"����F�����<t�C-�
Mh: ����S�_�)����Sg�̲XD|E�����hJ��@tSRp���_�d��F�*���Yrʖ~���ʅ�2�	��*I0�Ο�kļ�JX���8,�Ů�~�(���ˋp �/r�� ���#��	
�'e3�c�3�yI�A$7-�j�U�8B��̬Bc�N��o.#F�ۣA���@i�Ked��@�pPK���l�JtHpK ��M�d�����w|��]1 �l�H�E���[oT�K2���;K<�f�[�*�]�e�3B�6�W3�uu�3�5Z|v��eU�9����r�â������X�v��;Y�Z>� � js�N���R��v���Ƌ�����<V�b�tA�$�8�c�����i79���<#nD��(��u��od5$]�N4`�UU$Zd��
U��^�Vy���?���u�o����94y�O<����q���&]���|8G��%�N��-*O��)���-k�r'���5����7�v�R��'COR���A��;���,s�A��:��s����*���:��S�qg��P�Y$R�1�@\��o�O8���!
b�d
�!��,�)�0��; " !p�hG��JI�$�<=7�}{<�c��SM�'h�FVS�%���d;B�g�N�K�k��=�-�&Z,`.&)�d0������z�͍��L�>Unr����������
�=j����<�Ɯ�1��R�H�N���L$9a�	v�Ҍ*/��`����W
�|0��L�����==���Ë��i�!��L@��7��c�<N��w�*5$y�
G��&ޠ�N3���ЧdtZ"��0�v;�(������7��}�5��pK�R�j����6~���\���@��[�];��������xTj���ev)g�߯L	'����d�@��ke}*P���>ğ��#\�g�_�;ȧ�ȯ����v a�s��m��D��~G"�`��vn�l�����%vm#�m�&��'�{����}Ψ.�,�M��Qʶ��G_��O7ޘ�0��P8����^�u�.�z� ?=�����ޱ��^�vsL*���o��cs����-�F�d'�9����vLx��z� �/xBa�N�I�d���y���.y�"����`����G�A[���Q���p�;� �σ�DXf��[:�HK�%K�����@b~<ʝ��D.�cif�06e���{�b8
Z�^�г��n� v����Fdc��!́>��#){
��C��D�3T8/I��-[�1������#}y:ڥn�A;�]��E66���ъ�FJ7�'�߽{��jz�E��&�qW2_n����&S�h�_��c�?*�(�� �+|9��eSv�l2���8�-�XPH ���6V6�x��FO"9ki%���l8����uXѺ��xv���Yx3FU�;�"��U{�,�ȷ��������O$?T#�ŎZ�uC�w(3�,ks�B#߃{&�8O����Q  i̾Ԏ���ĥ��[m���s�0U��5�l�gꃥ��U �UKl�(O��uN~a�w9�X�ޤ,Xv��	��AzN�c�{Mݹ�tx6��"�9�C��X��L�E�'@1WO����Gr
!37)����(��(<�8=�L\�߆����\x.ſ{��>�`OBqB�����.wbLų�2Jr�T�����I��ɾ��3<a��_־���������-'ٱ~Z�G��-�*w]7ۈ�R ͺH:\\ >�}ǉ�õف0-T(m�TIJ�{�����@���"8XH)��٨�h��:���I�d��YZG���\c XU��Gk3�cpV��S�
��r��m�4�w	�|`(��oA�cr(S�(�{� �Z��|t��M��k�e��L��o�#��7M0������C��k^o���y����-ӧOD?��MyWX�`V��P�տh�u��k� ��:���z]���#�jx䎍ܞ��A���ņ�F.���ݡ1x)�<j�}���񼛵 YZ�j�?cJ�dL�ؔ�dk�x�"%*��c�~��"b�QM���T�̡�s,	�B��a%e~�v�L�ZH������sV��E���W"6��?nAk������x�k� ���p|��is���� "Q���ď�f�]�-�CM>Uvj�� ���e;bW�M3���;zG�d��2HY�嶦g�6��z`�'����r}��k�'�]�>v~�:]�	9����P% �?ϒ�*���̘���ڀG.�X#�;�~v����w����e�Pߟ����j���XX��U���4���g�n��w���I��a�[��i16:CƏQ��2��dt�q�)\�����^))��^ӳS5� zJ�xqY�T��S�F0ӗ��MM��7eΊ�M �/��	&��l��3���@%'D�,̇U͓��cѭ�����s��"-��LW�L&J�m�Vr����41����]�W�
EY�禳B��Ն�q޲����	¬�������bu
���d*��yv�46��$��$GY\���E����kv�����00����5�Y�,��������<��|k8���Ƚ���L3#dO^��Nս��ĥ�vo����M��H����¯��P$`T��~������xn�C����u�����H�v�3¼}%$tir1l�q-�X�EB�4�S>cR��^��"Ϭ��皢�;�6���qnDÞ��]R�jJ�r�����s���%rD�2�\�{���[�ϔ���ito�V�Q��,3�J�� 0�!I�[(_�z�=<R�8�'�#��\/��n�nަ���/Ƀ��3_N�,�1�^"o�e�_���W-NIiT���l�y�k6�4��X.$�����}Ъ��Ѽ�ʼV��h���F2X�Ȗ�~�5<[W+���hkw�����.8��<Ŏ���L���qU��ӗ1\A�CNR��Yp(��J�k��Am�~`>�Q(�n��苲|�	�{Y6Iȃ�W�e�<��b��gfP!����єfo�:_Cx ط{�cV��:������t�5W���i�Z=��I��s^�Kl�l=[랒���kS�Z�VX�y�e�����:RqҾ����Lj<�*Iz�|:��P`6c�t�T�H��jS=�C�IE�bŬ[]g�a�����X��S ���<�����H��zߚ�.��VF����k�A�Cud��WxA�<>�Id��Q����޷ϋ�&ڷ��;�2D�!���-JV��+��	L�Ds4C�
��Ky*:v����"���C�,���>��<w���V��t�ق&A[���K����qa"t���\�D,�%����)@F���B�+� �PV�bۼ�n�T}��y`y$t��z���������@�W#���&Y.����.`.S�$`o��!�cIY�)4��}���1��_g�{�dP�.8ohF�u�,"/��%�:8:CL·�Z��
mT���:�ˏ�r�=����p�Ԝj�e�po}�����(�����KP.��S���N�ًr�_�Y������ޏ��*�|��R�yx��.�cd�dv�������F�����0�^��o���F�������[2"N���Ĕ	�t���s���z�PP��ʛŷK������8��ban5�FaҶ��c�ճ�GM>���ug�ޙ�0�96��THa@��oK�\�~���ߛ�r8<����x���P��a��Bwf��;��%g�"5�_���;Z)���:l�0q ��f���n��_�4R�B�l�K��U	#�j�96x-�,E�.�k���������'E�I�}I`���Wv�!�5�=�F���01�2L�25���孕��Y��G������j說3��]И�B{����跹�3y3�]g�/(Z�@���G���)e\�'A�_�0_M�y���3`�X��KGtt~�������X�����|%�^��>����L���-DV,����3m(������f0K^P)D�Z��)��:��Ð7���`�Z��n��?/0�h�d��G��9LD�\�i�S�6a%����n�aǎWl��8�oʼ��#��� W�����\3��jɨ"w M��N�6�bT��n�\����+]?�ՠ����c�:�$Y����*9��g�m[˶p��F6۝�rL�Dzc�X}k�J��I��d�A�p��ZQ#�l�`��Lkv�>S
�
�V�I�[�V��xF�����4k��Sʹ�[�e['+-�5նa�b,erS9.�d���Ө�Ϥ[�6C�m�W��ф�D�j��Q��8�S���W��$��@��Cin�2�����f+��FA .���ԅ����w�6	,GU�w��/���I�g�]k�
$��DPѴD ���4I���e�#f�e<�YȿDMU���9$��C�{�4h��а�;����+��S���I���p5'
������A	F�a�/j�c��p<�D��z��Η��`�f^��dE^�b-/����rN��tY]��V��C��*h8x�jb^tj=�5$�j|U�s�o?��A�yN�ŧ�y��%�����x׹��!.~ѩ9|�/�.	�eނ�`J����I��1�L��[#J�=梦�� ��}r����u��B9�c�Bz&���mVb^kGCD�)����H�ri�;|��Fۘ�I�Br�%�|�eΊ����[��:YYF2�ma�w���pXnFr;�G����� y���C��q,��xZd�qa?����Y�4X�������}�Ҵ���݂c�*����ڟݥ�sm��6�U�Gi�Mw�,�QrZ$�J��9з�;���6�m�ߗ������>NZ�n׈���4�j25�YQ�ؤ	mr�y]1��S����7AP	D=?��c�v������d���v���M�U>��߿�}Ew E�WEX��\�K	P�[��p�F���F)��tn�\�S�%>)U�_���߃bDc�MX�$��iGU:|���\�i���N�E���6�.��KAG�})�G��!�:��ME��H U���м�j�$���	%
�VZaG�����-r����~�}pr}�	>m�t6��4Cc~�X�-d���y%�&��gFnC��\�	��XBTu��}�'# ������O��W�->��<�+�,@�v���<PU*;,9�a��q��j���NV�e�hN2Vv�̵�:�E���1�V-j,��wj,q=fbá��O�������=�'�*�ͭ�����G>���NF&T�y����X�ɱM�$�z��.�n�B%�]_��3����e
᥅��$<�)�$?��Q
�}X�\�G�4�L��B,���QsH)H4b:��/���c��>�\l���s�{I�������EjN$..0ٿ�r�&��E�!WӚ��RF�JCʀ�hH%+Z��0p��7�=�S,��$�n�߅ ���w������%��^iZnK  �TIgYT��*��Ķ��E	~�X��6!x?b) �e%����"����ͧ�U����2ް�}�㱵�]�&��@�&S��WqX|n~���κ���K�������N�����nXWA3���;�)QV�ܿp�������W���T����m�1��O�Z;�j�5e�N���֓��0ډ��7k��\K,ب۾#��a��c���h��
�t��^D����J��mn�ɏ�-�s}�iH�ݓ���HȻE"���R+��Ti���>Rn�*���-{��Csvͪ�}DiU�:h�xT���k�Բ��|�
�L���e&���
�~w2�U�z�i,�nv\t�/�H6fd�T�̱E}abUjwiOR�=�o#1�����Q�7bН%&N�<��ߜ�����Rw��� |k�2��1�F$g��`����}�զ./��=�?�(�E�rc-s�`�uE,1��p�f[�cmt��9���<�X(-��i��ib�[6��P������@q]�}��&��$��0����;�����PŨ'b�&��v��v:KSy�ii��̻cH0�m�}'�(*��{m�
Z�0��@��L:Y�Ni�y��p���0�A �i�(MG=��Y��?���1I�Z2Dխ��x'v-�|��)�J���ɒ�)�e�$�)�,�0m�D����G�����J�;�]�Ի�����$�X��5�(��_����c`���=��#��8LS�Ϧ�w)���+������Rҧ��DSh0�y�g�h��l�MC�H=���1cV���G�*��c�xF��V3�s&��iw��ڿ؈�g���HJ����Fx}	d�?���1���=:i�$��,l���VW�����|}��<��:�~�<1E�eb�Jpʞc`J]��GA�1����7�cI1�Jծo�E��6@�d�ػS�J�e��(�iysJ\>���mT��s��!xr:8�#�q1�Њ���u�bhgg (zԔ�<�|�\Ά�CBk�rjH�
��v�@/X����׃{�'�곭��A�,�������_Ծ� O�v
~"Jar��9x�Y5�s�_��Ͷ3.�}B�G~7��+�`��Ɗ8ҐOt�����g�d��A�t�yL��6m��7Z_���؊�N���r��ќHx'f�oiLЖD��A7�5(�4���篜���I��6��i�;�����?�����;�1.V��f�bq���'?;�ޱ�b���ΠIGy����$�5䠌/+��a�cg$_3���i"�)�ks?*^_W� Sߤ���{Ҕș�B^6����BEa�c'����9ND�
�*�N���L����:�e�� ����5 �!�pΏ��9˴��]��ՍYR�)��y��"a��*a<.@�B��ςs��Z}"ƖU\���(��?�l$��"�\GNi���W�DEb��>���b�N2����0)���}��W2+Y�� 4?@��)Z����_a�<Vcg-����=��g�*��E1��9���޽Tr�/+��f��u��5�Z]��t�[�-��U��,��ىϠ`��V�R	��7���L��r$@�nȳ���-!�в=Tz&s����0�'�P��BR��NY�c�t"^�˟�2EW�yR���EҘ��#I�-]�Gs�z����cz@;c�3�����ni�)NQ� ��n��3��s��I�Ic�g�V:M���2�$�� �M�C�+���{���������_X¾b8��A�@���T��m�{1���)�0p�A����ن��]F�r��H!L~/��z�����9q��9h7���t��
Kd|���Q.���x����cHzt�۫��[i$��,C�x%�G��TY�'krU�{?�5��x�9�J�Z-y��Wyz�s��x�Q+�9A!����g���޹��r��MK����F!�{�����s�~r 9Q\�H���N�'�?�E ���nv�M�{R��k�j�2�����bG��K̭��<�e���|vV;>W��'�� pD�1�2T�dAR�M<���'�ߦ.����{��u�c�F��\`��5b<�&�-='7z��k9\���x����QV�qx���'���a���#DR}��|���Bs��{��I�x�D{ �b�3�j��{�ͮ��c����	�����ɼ��4���^��$cK��Gj�A�=D���V��\�����O�v�au�y��T����K���c�N-�<2�
G^�\��O5�W6b\��}���MO����<�y��S�]��%q��s�J�t
6�w CT^���md�ie�k����2b�b7�p�#�!���\�,��!�X�	�I�O�ว/�� ��j��Q,��uD6��=� ��n��a� ����=��I���Lݾ����dp�!� 4@�3-d��Ep�� ��ќ9��֟�Y�Dj�� ���UP�.uM�j-���'85ܗ��$����P�hX7k�3q��{)�'��.��������q~�����QQ��E��~0�Z ��=I�q�j�0;$T|ڈp����dӝ�ӥA�A�$�����!D��{6�"���9B6�_ZQ��'���1�&i�O�����xc���k�y�L��\���7 8]��_V���wեS�!�l�M	ኟ_�P�/�ڰ]1;��0,�@J�����
ᶇ��<EΌ�Xhh3}ь�⢘�Y)Uaa�E�/��G!E���UM�b2"���^�K�h6�"o+�C�=1��Ez���皺8N���⸤;��2�6%
���1�����4	t]��r�FLsR���7�!4� _�a<��u�I��('A~��z�?w�<r��w� x��s�����{,o�l���H���<�Vj�����pw!����'C����f�>f���$9�븱�}ƨZK?���;��9�=p�vj�l����<�F������~�X�I�]�_6�Eph�����E��;*oP�<�4|:F"N������n�1Y@v��$"C3ä~�u�ں$�y�g���R����yLiI��}�a����3.�ez��)�io\8g��H�Y[�g��xt��ʵrg����K����eD�/�ϐ����rov�/H\q��^d�4dߥ�C�8���wl��R�Z�R�= �7ZW�9QY_�{�W��1��9��6A��9p�V����l�b��F[-F�$--��S'R�F?�	��\��P��Ư�Z�ѕ`
��߬YuXI�ɪ-A.��?~����1���xd.Z�Е�Fm��>�7�H:�)��K��n�[�d�I��R&ª��]��,9"B嘬&%�0Ab*ʵ.��H��3�4ܱ�:F���3k`OF��$82x����c i��r0]x�mE��+\O���)W��tp�O�AP����V"��w���B�	�-������ �p�J��P��aa�訒��^�5��F	PTz�d��&kX��N�c,�Z�c��o��g`B�D^� o���3��4���A@!~0�U-�5�΃��,�2! ���2L������\�_��z��$7���1��Wl�۝��ݛ�ku�K���trK�\��oewǸ1fw- �$#W���&��	b�\�on��7;~6�EKwYN�/� TRq���\B�9-��q�1�3�2������=p�0�̜�{����s�B�����}�Yy�*��Lӹ����4�	�q2�jb%���'&�l~q��1�\�S-�*�k�+O�
������K��Ty�3^�����#��>aۙ/-92������s`6V�}<z������?�q��n�m��da����Nxc�k�I�b���@G���	���kh�o��]�94$����^���?��<tT��s���&}d�}<m�$_��B�ۏ��U`ab"�i�6=8�.v};®�v�CFLb{~���6'�>�T`]22JO.t)7�����Mf?J)�����ջ�U�y�뇯��RT���>^�I��	�*�B�X=%���������1(*I`�<���r�2�_F�c��%��ȵ�RO�� A-��uE�~����{�������*�M��$ŷ}�Q�p�M�!�/��;r�K=�Q�3u�RR��,�>j?½����˄��ˮz�kEP/�6� �#(~���'���{-,�'.�h1���4�vۘ��햝�J�06����(�O���dn_������jg�Qy#��U�:�|�X��ѤW��n�m�Z��ʏ����)[*Γ���lG�;>�q�*�?R�E�a��/̞z%��<*��fUF1W��D[�˹���w�׾���F��A�q��|�j%�S����=���Mo.�7w@&I7�7�︹	�!�1ֽ^�r{�[]�n�a�l�2O5���+������������`-ǃ}��:O���oH��2H���G%�V��þF��,�@f������Y"5x樳7t��>Y�ܱ����ҧ+����p�bZ)t(�x�ݜt�gD9&�ʶ����`lj�-����g҃���n�p|�#U$(P�Ah�+S?����aE��=t��wT��z�&� ����K�i7}q�����7� ��9UxVq�NF�Jl������eU�q��(j��kEzV]��,E� O�􃹑�gW��~y%(~C-��K�gFL�Wҿ��	b'�M@�̀�)y�
��t����c�̸?a�ɵ�}���̋���o/�6q�q��Kխ�#�8Xg4�
zX��CLI ���F=����[��*!w # ��m�J�O�3F󠒢AəÏtY����lf�ƅ�d"֊a��ö3&OY�%��s����w^QYV�;lf��N��U�t�.CCo��̽1���?V)�2�Z
ݛ�������h�:U^Z�P����ׂ�Ȝ�	fKp�^�o׬�]
Bj����V+++�$���UP�\j�Q�ұ�F^!c�}/�����?�Z��p���r�tw ƈU3|���2���>s�:�Q(�6����^���`{��0� �4��ܵ&p�v�SdsNj�x�n90���� x�{r$�`R#��<��A=7!l��AJ1��,���u�,�VT�]���wAS񬹇gb��_�B�%�3�D�i�
�q��~��(��� �O m\�pi?���[�rh�qa8eGZm���#�+�pr�L�Վ��& Q��i����3J��%�p����*|��-�]�Qo�ˀF��s��P�p�0��gmrQ46�l\�(�.c����[9"�Ѽ��y�j�����Ոaw�F�+W|
T$�f��ca��6E�$��ʒɖU �>}8���c�p��5���!���+u��]�F=f�
Ą|�Q�9�6�<�-�q�9N��e�yo�S��n:������gҵ���y�zYj�y���{���s}����d3U��~�pܬ%��\"��r)�2RF���k�J���e�&_�/�m�3�$��W��<<��������^L���ZB��<8�w���[TRQ�%��r�f�����M��0��8GxР�nLv�^�Ȑ@F8��Z����8⣪�[ TO�A9R��[�������F�5������,ƛ8J���1>: ���jC*�q�ij��ϰ��3���|�p��<,Ќ�����#���H�P�r�DHƬ17����E�Km?;���3듵��(�!�$����G^ ٢Yy
~�����؃l��M�I�������1��������޾o�����2��f�����Ih\ �K���`���f�ɞcXM,�Y~o۞l��A7���w��^DKFi���[�)ݸ ¯A�?�$I��N]�(9� E�ǻj�|�!1s|gI�ER����;�H�Kn��4����R�ӿg��h�+q�`(�7������G���֩�t�X��o�H�H";��{��8��^Ir�yU�X��y �h�0�?[d��&?LĀ+Uh3$�yԋ=a{M�Ó~v���
�?��t��%i����e �Q���O����tf0_J��)Q�|�y-��J�DT�g
	Ĭ���Jk�i<��0�'��ͫ���M6�Ǆ
�W�_��B��Fkz��~����ꗔ���	�Q���"�s�n�K|�O��;0��!����nx�#܌ɒ�jZȾN����WP�|�R�4780�������� \<9��\m[�|��_8�&AVY�h��e"K4[#��H��Z�U�~�a��x�P7��E`�,�o�
kB��@�.����rt�� �Db�f��M- |m1Q	����ׁb������v#ܪ�U��v$�TK�
v~�A\VK��l������Q#MQϐ5@�1Կ��L��`'m���3S?�Kݗ����Q�}��(m�1���ƞ�2*��$�Z�e1�R�+�3�B٢���DiK��5��0	/J?R�w�kN��u����n�#i��{��Љ�t(�R�NDR]�!���@�4��u�kL�n
��/H����R]Y�֤Q_��_��U��>��r=�o���&��W�UAY��ҕ�)?e-q�E��r�ɟ7N�������/"��>n��{�����%�=�'W�8$_'mgȽ��-���jM��YQ�j�P�d��3Q�08�p/)n���i`��a��XM,v�|?3�N("%�5jU�\9�����4]�#��V�5Ci'���~[jF��QP&|	D-�0���x@ȗX���y)+9�J1���27_�D���Q�(&���(�����lf8���p��
��)�-t*��i�� fy]�z"n��Pp�Ez��6D���x�/N�
\iȕ>_���5�#�y������������/ �J�"F����.0��B��Of���NZ�Ԫ6t��?p��DP�x�TÙ5AM�2�۹����9	A�5���O���`�,�Ad0'X�G_C���gv��{;��'��G��eŋ6*�øN.�>��r%��uw��N��󜎳Ғ��)-��t��2��H�����	C�� ��s���h<���PC�$<lw����Ye�Gg�\�I��nq�@��j��U��!�u�4���I���d�b�g\G�ш�j�ۋ%7�1U���xI����Y�_���7��3��L񮔝�]����`��@���@7�E�����C�
Ϧn�!���1~�՝�}�4�]cIWVu�C�(��_�
~�>t���3���q	����J�V ,j?(��D�L�f�h���B��2~0����0�`_ݟ�~���-���K��4�ư����+�4�����½7mpU�������6�Y[^7�v���"K�Ệ�ɽ3����\i|/����	��~6/qG"j����z��*�
���g�<�6�d��5$�쓱�b3��G@Tx򇳭��1�)i�ǘ~Hɪ>���\��56� #�WA�W�t%��m������G�(�G�g�T�>��d��_+���U�Ϭ�͡!�4pA��Y�^��\��{튽l;�a~��Xv�o��AuN@�q��^���L��/ �p�t%g��F������1%h;Dd�L5t�7��[P�q�l�`ӛ4��w�G.p�JbE�k���p�)���dR��wL�n����N�(ɠ@]���,��!��1��y�Rh��*��z�r��7x�K����L�����?����q�4C���R�}��a'a�6��)�g[��I������X��.X<Q|P@���0���π?.o�x9^�t�́��˶�	�Vb�a�tu�I{�1�n�|Zx����[��A����=��� ]�r�����vY|�H�`f:�
�N80��hy������K� qs�P9���l�՛�W�
�U�3v��^]���<�*���L9N`ͱÃ�ˁ�<�Y�j�lP��Q�7�0��Ie��w�,�G�2MF�7�''G,�W����w����ghE��D�q �m�-�8/�D&y��(�	ۿe��y��<D0�Ǵ��E��Q�4E2�J�5~Ĥ�
-���凔���l���9���g%�'�:~nI�С`=�*&]�� t���JI��-�'�d>�Cc�B��q�Z~�n��}�Ɵ�әl=9֗m��"�]��72��z?����;�R���f٧C?DsY��DQN��:������7�ϗ�R�Ś�pN��K[G#�+
1�e���l�>�-yA��}:���;ס�s緄���_���7}��v�:mq�Δ�P�����E�H�ӏ����?J���,���j@�|���Z�5���`�pҍ_?�6xa�­d��ؾ��D�o[< �n,-Z��=K��>lmR�_7`��E3��8�!o��Bɛ3��;3K��Q,زH��
�T��O?Uܰ�
�3>�Ӄ���lt�G_�����u�zkS/���Ր��x,6g�0�v*�%E��x�y�����<����@A4�ٶ�'�K������|Ѣz��## �v3l��`&OoԅA5Pv�,��E� 碴
�vz~�F�LJ���olVOMߖ&3�y�S���E�M���q����:�Q�Ľ���>o��-�3�0����~%�� B�+��T�,eH�J%BR�I2qՐ�w1�(��{c$� %�}�PT��=z��~��
�4��^J���H��7Ւx����G"�֛E�/�Â\��"t:�Y����������G���4��	csNW��j@����7 f�`Mɼˣ�p���� �Ơ���q��%t�RC�����Ⱦ����K���>.66� !-5E�m�{��Q��oK�`	~����	�H���J�1��(k��R�Mu�,\Oy�3���r{ �B��������vXY}~�ע ���ܤ����\��1w��`�S�i���L�K�k<c��՜69�sB�Ls�"�|a�h��pLcʌ�R��,N-��S�j��w���L�}�c�Į�i�N(�x�g�|����1v�u��0w�F����2�8��i��F!��;҃3?�}{�_$Ιtk�Q������6�q�]�&��b�����&V*�9B���� � ψĕ0�G�S0>#@���� �3\�k�����O�S�?Mr��_�'����Ob���;�k��km|�g�gޣ�ѪJ崉�-�J�3^�U�&�>�a.1�. ��u��=8v�ـ�i=º��c��Əj޸�+�y7.7D!��圇%dra���U����$+��|�V����r�\�"?uVK(VĤ���i.������qz���� `��;_�	�����e�G�
�fB`P���],A�>0%�ވ�u��_H�f,f��_h�C^�4��߭Q���.� o��'qhD�m���Iй~�-�im���YWwb�mP~Ub3*�Da�gO��
��UC�?k?4%���R=�h�d�ɖM_�����#Z��х��}�[� ��]F�jR�H@۪#Z�%;����5����v��8�4s��Ls$�N�y�|I5N�����i�6�5��b�Y��ݓL�g;���LYl >���.����|��jZ�g$nH�V!�A����R���h����K,^예���bc�
P�V7�Ը"池�`���W���6T=K����6�m
�0�� qHA3��H`���
�/n��p~ys�X¤Xׂ��Έ�}�Ld_[��"�B��eR�/�<�X
O��b��Ml3K�EX�Ӳ�_��~�{��=k��5jhl��Me(��^��Bn��(�� u��������D�s�� &O�㊨v:Nӥ>ݩ|�$
#��2�Qi��d��)F�;QGR�)xŠ���Q�Ӫ�G?��"�s�fm�fFuu���� Pno����\���w��`�k�[�����>��`�$M�{��OI{����<��f_'�YDF���_���>zc6�B|�=��3��]�#��㝧?�?#��rc����J?����!�kkq�W[��]���F�T=��)����t�cuXP%���JC8�$0]��:"�n�N���*{_���=m���^"ۋ�l�Q�V�=�gX�PL˛����"g���Y?�8���r��/eά�UH�i)�~��bϦt㭕�������&�X��M<�}Ѿ<%"�s��L@��g9�g%!��\C��ȕ���0s�ʞiJ��`�X���>J0�������7��B:�ic�w�\��?~5L�R7>�N��{���,�T�<%
r2Sܬ�G���򱺅p,⃔ s@��w)�(&f�����ϟ�7;�,�	�H����5�N�{3�!�3˙�|�^�~��gi�DrDߥ؞/߶�_޹�.��8���TeŤ?��@� �s��nP��cQ�:�R7���-��WI)�%C8<�"X��na������̭�kǁ��<<��A����������-?sRY�=�� �V-|b|+�,�i$�0�n|�OH��w9�J��?x Ĝ�䶬�/�I^O+|E�ht
$aql�=�\/�7�t�n�R�ʛ���&�4�Y�����yp��[k�¤�D�g����J@iΣv�Ӣ>(���6PiH��zo:������^��*�M�pi���-���`�����6bGԓnt&XY�qm�&ք����`���>�./e�)�=~��yQ��\�]��,s�7����F��ũ��g���tͿ~��J�*�zc;��9�����>�ٲ�뾾��md�qf��u�Y�$�%۫�Q�G?�"��Q�M�%���T�?��wMw|߇���q�@��4\��p�uI.7מ؞�5|���U�U�0o}����������@%�.�Mo�!��΂q,#�
�v$��58�j|rԧ�ң6ϜŒ���<�;@��k��rȑCϞh�����K��P��_�h��d���\�,$k�m�3@�zǓ���붖�ED,̠��i�����h�	��j��:�D?�P*c��L">��j9-�X�5��&�>��U߂^���E�?�׌	^�g�@����m�S�T�ß��YO�S���4��n$cT#UUH�?"R/	�C@ĥQ�FBӛ-0aF�P� &�N��ރ�a����iS�,R6���By�M�C�!M�w?9t�'.�-=�/�ǅ$ѧ/��D��:����>T&��
�f�(�Wq�h�Z/C]�#��v�5���[܁�5L1������i��A�ul:��,�6�7�A?����x/iޮ���)�(s���Z���2o�RC9��G��&���΅�(�\xq�x�yxD)��� 7���v��kyc~�|u��D�.�wB�H�T�dg�"�w\�n�o�'�\v�\_p�*������	^��9j5n��k���������'Xt�+�� �oQ��9�5�Q��Z�Ձ9��yO�����.����Gn7����<��7���XXdn6�#GueϏ��(�H��/��2����\
ÿt��I����jlH�Z�Z[I �#"D0���@�*�8i>Ͷ��U���^*�{s�Y 0 �#Y���yp�2)�'_���*�O%5�����2�X[���Ӫ�
G�lZ�?�8�ŘD0��?S��l��q����� x�l\΍��B=����T��+��z��Y��Lt�ĭ(s����s!x=c��D���)w��fu��YT��a�c��p�,������A���4�%����3���渰
y��Y/'TM%�(��Fo����>3�N� ��)u]]�37�rl��������l��
NClS�/�r�m�#�c,|�a� �ݖ�h��!Q3L�7>���n#�e�I�2:F �4�f��]��q'��<e����R�����6?�]�x��5�Tۡ�;5�p�e�-q�'��2z��S�����=�e��\Kr���yTl8��������3�3g<K�z�yX�FggVY[�}j�e�O�����1�Ǧ�Z��3��U�a��2���@x�D/z(�`�2BcW̞�;��x����m��Wpz���|��j/^Z0ƭ༴Ld3�2i]�iS�����EJָ��N�p�,�)ܖG����r��'��2�Ó�*�3�H�_�)����D9B�������X���v�/6e"sS9^��r�z��X��R|q�W�o��*(�a�s�c���6ȅ�b+];��O+k�d�b`��70��>��M�f�0FMYE�H"����r���e�.�� ��-��j�35@
�I�@���E
��+�|!�$$i����i��3P��z��P�V</%���	OX3-���_o����Bz�Ɉk:n����'h���
�:;�`�]�?���=����?��jSJ$��rY�q�6[�Xy�����+�V���}���>����/��lľ�꣙H_���s#|]��⫕��x�[B���l1�z�=����H^(�h����Q�v�i�=�N�%�Y`�+P=�5���N�U�H�r ���"�$����̪�'�����gA�#ѩ��%�eqt�'�#�m�Oø �f(�_,�LD��^��]��-'�^͢|�Qo��I��#
e~��-4��&���ʙ��I�f��Tad{��ΆO�S}C�\�Q��;���+ؚ/Ɠ`��AN��Md���v��Ց=�9i�:D�ߋ�	�W�gYφd��a�U��f�>���eI�< v���*��Iޅ�S���q�C��j�cj�G'�S+¡^r��C�I'�p7r�)'�%x�>�N���;�Bx���eX��aQ��'2T�pk��#�枴~$�Ҡ5S�[֥�-PV���t1 �n���J�!Ն���b[����%�e����I;(gjR_�麗��7�C���Y�w]�i�s�s���
H��4'.����b�G�i�"N��I�;�u��~���4[E!���G����!�/�0ך��Lɦ5�#Jg`r���'��~tk�o�h��FF�Z�W<��N�&|3 �V%Zb�<�bw��nz؈0Pzi���jF�t'�5�0+�5��t��X�ݏ-#�};�W��l\B�����'\ 6�N�8�"�}��`�>��z�����ץ���r�'�����9t�oF���L3?o���<����s�d5��2��(&��*vA�F�>�Rh�1�VZ���$J�p	�@����`)��&��y�,�&�]AŎ��J�qTiMd�6�R����d��TÙ[���9�jY�9O!k Ɛ1CeTb��.9v߽��DV���oY8"��SG��đ�����*���D�0M��f�&�lӻ.�����_4G3�7���wk�y��(��?m��9�VREO?��2��LA�#���cp�c�"M�2�S��\W��X�� 8l71�Х~NGlm��nh�.@,	
�n.D�m��#=#�k�����z�����O6P+Cv��i��M��L�Z�c��+(�&��U^A��D=�ϒ�$�>���
7�:�\����{�_1��QBEu������pt��W���^���, �+	�ޮH3z֐���{�ˎ� x�ݷ3�y�,9wE��S�Q�mo��415]��;��Ӧ�]R��^��x�U���O�m�"!4�K�_������ T���HU
I��F��6O7=�	g����6-�N�"<I^�)��_6���u�CnP%��c _m�*m�
{L��n�S����n"#K�/���6���V� ��0�ᘎ�`�v�N�F�,�M���}�)�@j4b�
�E�y��H;�h��,E���3�U�ǔ���A�����c���\μ�+����7�jG�RL�ݲs��*E���L�_�l{���*�k@rC�]y�S-jX���]K�A�jl�ƈ�&)F��	I�˼�ڕo��F�q���h��~����r�G��W�;~�	��0��l���ZY���Ǡ��iԗ0[O��+����S���'��(�ܨ�Ƴ+�E�Q��`�l�)�&��1��?�$�i�NX���s���1 kR0>L��	^�,��!�5}w�/�����U0����R��������`>�Wz�4~^�A�d����]MzQ����p���yu�R�&:�tX��f�F1Z��Բ�`5�:���B�3��װ62�����h� �ǘO� Z@r�3�W�w	�Wi�BP������y
�A�4�'�to`�Q�s�
O���2�0U5�E3����c�]W� ���\�ي��� �j݈BT�vAa9THܐR�@�w�ՀJ(������n��I2�f=S���������S3�w�����a�S�,�.�	gC����x�i1�^�JB6p�56(Q�V?�۩���2C��a��Q'�|nc��k�\GX�XV.U�
��rʽ☀��S�����O���́�ߋ�iR�1@��N6Ѣ"vy�*�w`N���^
Ԧ���?��G�U�"Yx��_�_ݔUTa�����D��O���V�:�+����/�mi�ǿC��UH3�k��+O��*r�=k��+��Á�� ^2�<T��V�|��$5���җ&�fVP��ۂ��O����X��JުE��_٨zr8>��6rŨ��K���c������7��?*6�<�f-T.����tC4���ϡ���%sP�7���4�p�y��#ֶi�?B�Vl3��{��F��bq��2����-p�;��g�O`{!�0,_�VK����-9�p�;�*�ЩӘ�X�$Nݪ.������(Zc]���u�D1���~�P��`���MK� Nsa�8�=Ф�yc�tS��Ｕ(�<�vc���Z��|�(��P|0�װ^����!��W����s�yzv�˅M5�������j+Έ۹�ęG8��'|�?_p �!jz��\�, �t���gZ��$Y�^K֩{Ȃ/|X��)睸~���
�.(�Z[�|S�W����ё6���ň��l��ݛ.�Of���ٶ���	z� #��5M��U�q2�t�2�4X	�k��CꝌ�R
�{ğؒ;�R#ߞ��|p�0�������<�pC���3��eͭ�hB�3}�����K��;����WC�ga&H�%�|B?��0%6*�Y�kH1j�,h|g�A橊aj�9�"PQ9� ��KعpD�B�V�'��U�#�$#�dQ��� �.���l���*fm%|8Ln��rY�Ef�'�;��5���*S&�92��+�;($�ϧth�ROV +c)��M�B7���bѿ�d���c*�3i>&D�Ј�&��~ːI�������Ǉ�俒��bP�q<�9�^ъ�9@�GV,�v�_N���w>/��-�R�YS;�ޖ��)ny(�տ�iRՉoz���X��!o �ˆlQU��{�lĴN��T6��a�5o�5Q�ˑ�.�3T��m*`=����ZK<�H���G���TJ~�B[���#�gs��[�_�?��w>���e��'(�
r�d��e�6#b�f���֗��b�;!��M�~�k(�{����p	

��x�+v��qُm̩��(&>H�u���ߗˌ�`"�$Ȫ��w�>��TQ�Nt�@]�ch�="s�W��co�ۧu��M��V0=�h%�cQ�ߙ������+�>A{�J��I�vu�=U���u� �/��0}�e݈'��l��4%������&�Z��G����Q��v�֩��!��B�Ye�O����A3��5ᆊ�H��V6���ӯ�Y/����������������-m7a>��a�c�V�g���+�������Y~T�.����$kT�	����f�����$2�0��-4���eM��O�I{��_l�^�q��
���P��.��w�Qť�ͨ*b�P�~��V�5�)�8[���S��x^,s^8,�b'������Q��Q�ߘ�����x���&��I	�g��BM)l��o��e�^�R���2jg��*+�=ٌR��,�&Tb�D~�������/�Q\�����'`�^��*w��o: ��L��A���A?�dA�Q��>%\i��+?
����A1�E�h�iQ�xy���|���΍�ٕ� ��]x崞���l8�̞F��7Or4�HY�
̖* �E$�#�*!V��6h�}�{9��s=��\iLqU�w�hhb��,�9�^Fť����ý�X�@w��DQ�zr/�_9E=�ao<��� ���*�EQIF�~���_v��O@p8�1�]���fw�jC���.�+�I��j���>�M=zκ���[\V<30\��l������+Q��_�=	k`��a�.=_>��,�sa�&
���W������y�K �RA*:xZbeS�~L������D�cM47Z.&�0�e��ӹ�m�i&�G�{�:p���������l�"�XH��5IVvь+�����K��r���W%E�տ��p�pAȽѺ�}�D������� �0��}�Z��2���M�o�,�qC�ZZ9:���
�¥����gȕ���I��i��0L�
���� �-����o�����U�~�)�0F>x-1ui)S$ӛ998���sࢢ��;1��l~�T�ͰCݵ��Sm�UD�K���_���t���h0�ż@�܁>yp��Y���t��V��P��=�����R ^�`y
�2��m���Ƙ�TI�N���d�eA>�ː}�7��Z�K�I����	�����-�O�п�+��.E��Z#!u 2,N_EԢ���PU�X��W�҇�U6�Ey��I:���#���'	�UGnI�aMmӡ��3B�L��G�j��}��Wr�_�{JC�c�qZv
nݞ	]�4y�Ig�3����fu�l�  T(�M=<#�(�c��������Jm�=���<$G��5� �<_ҫ�ի��]����C �������'��ur�s
�t����#�&�yN��l�����'Ҋ����d��MKA��8��KLb.�Lq����j�M:H��MN{�=�-?�u8X��o��mK��P/HN��C�\m�N7�o�C���,�R2<�;%����Dr\Kh͠ӓ����+�kCȊ|�UѧKfM��:Vt#� !l$t��769�=�3ϻ��(��H��K �����D� G�+IL;�B$�t�I)��]�������[�W��˳C�6��D�?q�:)M�[T8TS9�^��?$D��~/������t�DU�������V-�1D��T�/�Q��g%Y��[���S.^;͙��, U1݇���H�8(O�
�G���[(�X�g�A�3����9��F�gJ�Y �\l�y���{0�"�_E�>@5Ҷ^����ú�<�ܗ�ѥ�����M����=h ���:&3e\Q�� c��jV?`�+����ږ���M�R��-�V��|�� ;����Oh��?��Ul�ⴔt�CD1)�!U>�.�Ө�Y�Ԅ�L�0�'S���Z*=yK�W������tF��}iG�~V�OO -Va�KU���z﫵�@���R������~��VΣ �	:�92�*�gXԒ����U{���?o�*��	��3&O&�c�l��A���yd�b&��:�䎿�V+��7�c5��H۷{u��4X��[�:O���p��͖R�Lf����q*[�QH����Zޕ6��U�4�桬S>�#�r��uY��Qs�H��D*�|��M��3�L�t���D��ӎp��hgŬ���_k����Нõ��M�.����6���I :�a���@-0^$N�T������¸�F|�桓`tHJ�_���#��Щ��7�Gs�l����U�tֲ&���7���//.���Y�]*^r�e�g@�}�ef�l�ؖ��w�2)���M��Z���0�=t�h����b2}Ա\<r�o�̧S�{�v��k@46]r ӎ����(�l� ����D��mY�j�9J�<^ǀ?�3�唘/����ZS$���a������~�u�t)W`ex{�Itnj���MF\&Ԥϝ&��i��f����m�����8�%1����h;=���N��R]�{�x�z��)��w=ߞ="�#!�ݠB��i�������d]V-5�Sn��!g]����xG��=տڣ)e�
z �E��ر���z#�:�O%/�U���hO7���:~n�l���]��e)>n|^�<Nv߹>	�+�i�B�W�9��aN|��B6ԉ��'���*k�7�{�f*�QX"��.Ǹ�$G�2I�D����l%_��f瓹3;���<��r���Wr�	��ب�^
���B�3��	8���]0i�6�7��:��黖�?�ۯU#��u�1aB}HP��Ӳ��46��ˡ��O�r�����T=͞�4�dwGgh�5ۗ~�0b`Õl�jJ�p������AG+&(�
P�ȉ�i�ɂ����BPU��ZZ��g���H�~�_X�����1�LS��������ѡ��P3�B�E��tW_(%�R����O���*B�Y�׏�ϗ��N+|}P��Բ{�e~K���%5c��ew`��� ��
N���{�мE��09>�VP��!ޢ>�Yx�ϙ��+\1z�1��_��m2�Sy�C�2�?���y3>����ja�{j��4�#�}�T*G�,^V+#Z��(�����s#�(`�����߼Z7S�4�"�Fb��3!&������[+��["�O�X$��&���ja1��1g���G14Σ,�Ix���a�0�Y�rVas����o�\�a��}�_�j9����}e6�=�5���2Ҏ.�D,��GO�����i������#f�Q�ܞDg�!c��͜�"Bu�G`5���cZ�v	�/�F96Uж�.^Q'��F��SW��QS��߲���wGԟ�S�3�4��~����IMe�yx�����܃<Fl��:�|���h�D6@�N�d*���
t	%�8�q[d��ط0H
�6ҺH��L�x6��F�[V��2�exA���N�;�[��%�Rl�X6� 1f�a�⹜���)LՄ:��.~���߿݃C�� j^�x�ZP���9`a���X4���&Ym�� �.Ď9�Ί�fRz����o\��~C��;��/Y����	*� Ϗ�󡹥�I'`t���ٟe�� ��	�����4M�I�C�"3!q�BV�U���P�0�5g���`���4L4��	��~��3���"�F/��&���*��H�Bz,��'x(��9���c�ӳ�\Q1<%���Ӷ�`��kk4�0���v�^~�F<�~-|n��4�)U3���n�;��;yd��������nzQ��)#ʷ��N��:&�FX��[�Y�`:]�[��� ՗�+m`��@_�3��5o���:��9Y9�>�J��7�UZ��
�G!p��lB�V����ے'+��#E��j�s\�f^�ů�/�� Ua���l�fKɑ�Q>� ����X�R��t���w�x�N�s�S��x����՘����7ܢ���y�j�U[,;'�����Z�����ض�dO���e��k�6���	���ɞ�$��XޑG�)*�A��ىO&I27Qʥ��9����͍���qE�����Q,t��1I$�w=�^=}�tD�z�x�X�l����è
�ߤ�7�z� x�h��k�U��BOBQ3����PW����y#� `�7pbv}n�>wbJ���)��vpາ�
��C��s,u�&7ҏ�
��px��3�ϔ����{q_����R�qmE���<Z���4�M2��z�rQ�ү�����"Kk�7i�#���k� ��⦨��`��cZ��M��[W$�y�`�%���e�j��!�y,��	yJ����Xa��_e
'ta���(rV�uMJ�{���\WD<bށ����<@gQ�<����ZU�۬:Ũ��ARH���&� �l�1�^�u*���+)���z�O�V��U㩒ǈM�����~���s�=e�sP�P��H�?~��( 5�+Ue������3�}���Ǵ�9�����3�������YNd���<�;�������^q�M:����&�����>�[�<�;%���dd,�����us�.�؈�`�e����f�@�8���z����novR}�P*�|j��_Q�~�{Z|�M0;�~�G����>k�Ũd�^���Y�1�&�g����M�A�b�zV�&��$k�_*��5�?sG�����R���d���g{�IAW�7�k��N/
&:�x-FՖTv�R�;f`i����\�I�K;`ڎt�����	-�6���sPD�����N��qJ�� ��?�v�~!�p��H�k�8��O�u�;��f�xm��SG����ӕ���S h�|ђ�\]W6�(9p��5��{ht��F.�C�25
��h컉�� K�~���%���D�r�B��ω���vh�y�;s���z�e��z���k�
p���k�'�U
#zЁ�@��R�0��Z|�^{{��,~Z�V�!&�$��J��A-#����I�^�i�0ź�f/z��*>�A�۴Vo�/�K�| M�t�M�m ��1%&�Y��S�B][��V�����zD�ƝA{Bb~w