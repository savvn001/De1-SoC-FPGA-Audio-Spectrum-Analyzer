-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aITfLCJRpM0FtLJ4w+QsIfWGma+54QYBTueHuuGL8ybS71hoSCYWu7VVxzFFbUJL8/P2EuRDYLfr
hOTGQPn/dFuXBv39W6dGYe0rfReUxBwQkDKrmDmdHvyZWrQ8G8IVKZTd/y03r02G/blixGTfHiE0
i2OPGM8x6OVe0nIgUbSHSWLsVDFMrrvuiSTT6tl7pdHR4p6I1d0QfebrzDVUTo26bWiXtkqKwpMz
IGBJGsxs9szp/eA/Mh2rw3BOfNJSSvENk07E+3XVVpwxha843UmEXhyGtJMSmb4LzDLldRKfg/WD
HB4KBBxUedr9//toE+dmomelI7VHKkaUBsDHbQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
XiFTDEVeXk3QWCGdp11Z7Ie+dx4vxcXpKw3QSd+G+uc9qXKzPYGmMTyVPup0litS0FnRRAMgCGsw
BIO1qgsgKAlW4Uy53JDtxb4UXPRyBIogQEwwRZGXpfgB0sOqqZZKnlrCxFS7byBQSmmNA2GyeYMH
Rj1ERRG9dPf474I7uiX+/J0uSDDIFV90Z/rdxxms84MQ7EIjlmWAoSpq532dJlJjHwORmlYv4Pxm
R5ethEzrTH14yr8DQs2Qn/pCF1inQ9iVcbzTzpZr8LzFs6cLPi0IniAG23rwDt3QUMGTyYoKqOIb
xu367VBmwNiP2NmAk/3jIKCMaS+f735falVApQ9QbMVZkKJVQNx6UvA+acdwjyUbCJDVVwLhs77f
5i6bt6xKrMkyfD82IDNnP6hGwnxU0aBiOro3KWmx0syaS//Jtcw4FUSrMGhyY2Mxdd1Mcj6uzAK2
EoYSlViZ1oxVWX+4nSJxUxVa2FYB4VzMJALwfHI4fbPJz/klg5mTETda5wCC0K8GnJCvbc5fY7/u
gxr6bz/A5qk7bQy/7iKm+1acRHxUkxx6JlXvwtB1rE2pSbyDkjjcOo/nd3j5g1AZFIwx9POYfe+f
c3Lvg9wV7K2P2sZxH3o6rlsnOlXCjGVUFyS9DcKKGrhv6kzAYHIC5CRDUVupb+SUzuYKMf8xFbhr
NqEjJ2j8s1K2Y8Q0Q4XmKBH9k77wqaDzwmNjgkQ0FimT++TIa1jjJ+fQy8D/Id53wdA039qXAdBW
wZbmIipnXGWNha9zmqvyh1t9cSvoRccF41MjvuZNtMd4IjH1CWJLGdeRo25wSxsklpgiLcFQvZ8g
WzLnTEh6Zq8W8rhvWutCRdWABHGSiqjb0oAB3z6rjxUjTE1sBDRMvCqWjTkmp9vETqQERPD8Vh1s
L9Oa3FUMN8n3afRNYedaAOTCMcEC5aUoiVqBuyDcU4r+Gv79/yRbrVlUqTyiBa20kHMWpoLHvQyU
gbTNOpDeRo+o7DQDF4CdNjEuBPcXjpIi+MwbW7Iq2wQAuAArseRxeSSO+QoY8Gkf1oR7mKZ+AXR8
XMHQvHDvWpjVpeLoU3B79dJDNU/3C1q/amUjSXtVsoBxaJPl7hj5ygxXVMmAM52oAsxGwd3veNrE
JVXJpBIDVPKLtXZZc0Moek4NqNa0SHiDn9kdmq1swtABw6dT7rcz5J72TuCHnw5k14aIQv7CeT8O
21wmlOfZ/37SiOTxTzJLyAutqxPE2lig93qfNvmEpxVckgT6uIfd99hCg8YI7oGqaP+k49uz0jpl
MPh8eoUUEVFl+G/VU+xODN2iyGfT33eGO9j6LDtiiMklN/5bthTOlb9PVh9tb1lT7Nb7Wl8Lb9fx
KtS3Sp7ygYVeHfRPUvxE1cdEEESBu+JszH4Dwkgf9VYWYVn+XRTVa3kPx42r+G5+Iq6YEoB3uy1o
rnDtVnTJ3cQIcvEu8IzCb1OnogFHzZxlYAofc6Lk1X//Le5g+nghMELQCewxewkWZudQ90w+AS7h
vah3UypT96043ssiYeDbr7YOEzIjfhk3+uV3UKO7rYPiAlUyx8swlJ44yd+W/evok+pco8sKXBSf
aw9plK+Og1GGBlJOCZtP/ehRePR1DoGRagDWRHAnXfRNQe8w63uos098JJ2/nBbXOxx3ecQLGFsv
72F8Day+nIhfLBzHOwwNe/DBh2gcXo2hB8NOEZpN2gUTls7jgnkdqihbmimYmrXGhvmE9sD3JPHQ
75v7lZ92HzBKTireXOHrtv+TohmK+rqsYLue5KFTB8f32BQulXCsaOM2oUFEbh+8My8ZLoSM+hOQ
LZPkOCSSI/wOdvWawIUmpdIzR3vZzcB84j8ho39yJaQS66eKDn95DqHqKs//RmeMHmcYGY+VBHMD
a47bRS+rG2Wyl6mz2su1BNxibSK2xgt8VHqQK63uZUtSVLLwk+VjHq6uJ0EY3SIiMAhBgsC6Bwj5
B3ilAZhQQ3xtyUVRkGkKkbacUJJeeu8Fag+QjLu0lS+5AB4i6d78841voWIlC5lUQ1fDUrhUkq4q
/jYLKj9YCsa//ma2rbGJqytvFVQ6Jdq5EOSrV2ceELb8/cqTj35R4iHS6GlFrlKXeG+kLMZG7FuE
wQqctgDpvnzMM7EEd0P7ZJotR1qx3TxpHTXEHxun6gkF8K8Fi8bRhvYQEC4g/BO5Wa5Qzxh6CQnF
SkqkZIInKt6LXcZ/YNHxPXVeOkiSduRVJWkn4Ltc2o8Sapco8SU57MaS8bN4cdhNzRt4a+Hj8nmt
L9ODu/3qKPkJ351z5JvuH9893KtdB3oyXV3ilLzoeb8v/gCpSdSiz7gui0GfkghHNthlJlALawsg
luKbRf+SulWavpI+kR41eVlanfkAdC7A/NBzaTvq1bCsXqki7xWhLjnGlPNK4FjDXdNn7BnJrdIE
n3RUp2qdQlhmo7NTZ7oZ8l5Vuqv7xFWdMsTa6VZHi+5VfqzhetL0Q+42EoeeJxgrHCwHGJHvRwCL
TdP5a+1lnlTIWYlJHY7Xt5WtMm3FG1Kxj7QcqwW6cZuLhPGdyYvIZFWEVvpGJBFuiy1aw9D5iebv
ObJc6F3GPJKoMv8Cpn5kdPi5KBCHgpnQchIEwxJeB4fqL1lXKzwKzQ10QXC5QQELYhff52sN8kqM
Aj6i4+FY9RGe7LIxBfIYHxDSrmQw7ErIpn2JUlO46E2Xw+uwp/WOIyAgwjMIeXUZhhpBU1AasyBP
uKpMPOngBVeEY2fuJY8kffDJdH98g2BcA9mCo4CMDvTUlY5Iu0WPFzqzQSX6//91+e1F13aiU+3b
D+BGL203n4cTngfqOAnR7hzwn2TJDspBz3Gb3P/7Q3+kqv283oMtRl2P/VyKBTidD9pgOfycmYD9
Zh/VxSm6SodeSNFtxYJTRGnuEUW5aD4UhzxXbdU0P5XhvzPnVfZbrf4ins0XYY7D3lx2e771/MHO
5f8HgKAU1UdGPgGFwTzDCqKh4PanVfgd0UT9Edr+9EYb8b8YLoSAiecbVJqHngZdUyaxugBPMH+B
oIY+Ax+9ESkdU9gw9l5RJKFAdAk/bVs+QW73s8PWB9nO1Fy1xxN71bl3Cpz6dh0iwpfMYF/4QNV5
/JLWL5eZ8nD/dLpvF/E95+SE12KIQFDMmcyYxZSOr4BZmkxccIck6VDpW3Ntytcc8Nk3OVYFQqkv
Tk+s08Ab/QWYXXXxdEYr705zqE2NBxSBzkAUWPtVFJbLOGyDiKL4RZN0Co9IskG4alB92k9RBzWj
shPOzexPEAsOQiO9PxLm8M/vspDsoARqrz2DollAhl6eD5Ce/PARHruUAJQg0NSA8A2+9ntSo2tN
Zt3LHFJ4bLzTsS/GK8TYO8VH5jZzU40NU1a+aXPJrzHBJ9gFPo+4YU4FOcvfWgoB7yRoYE88Q76k
Q/SIQelcJ/SRYWXufnftMZb/bt4JznR0SnmWk9+d+U2WrbhvwUkdewr/MK+ZCkZQs8wJPklDZ3vB
FKnxqNZhPbC/oJBdQZLOQQR1HcBM1HP2J9zafAxuidn/DGNiaBh0lZOlurnNZ7NS5Z2uMfGjHwGJ
KOhBMxn5aiMTsY+hYfSwQIfKCOlY8Ka3vwcwYQbOcF2+ps7nWMOqUjmX6GBsgqPGCCzewkCMGBDa
Mma/TbK9g7oVdFPT6Nabg7aR9QPuvn+mPBono1i+D53Wy8KXzMFTp1E7BPIgwDgU1PeP3o98XqEe
tX4kJ0HLN4mTCQh5SRHNxp1lA9bGjJzxILDDu8xvYxg/2vjBB8c02OndciCSyR9NIKJ46j8YMaAI
edVMiDNShdrb9AA62DsGAETnrpdLQmYjCufQzZ4ANP9eDmtljSJMkLaq0WJLXYlmJgwBb0Cta86Q
tdATlwwHn9W0zBG1JKyF6Ds9coubyEsq0nz5odtNkAyoAuGgd6YlpA7YRqrOPNKh0FAkk6f3yPor
+Sw9jbxDFPLv8m/9RDQr7cfdzc+r0Y/jkqLL+e7FibNNK9Rj53XfrFNNypTgDBqvGpRob/1q+ks8
HnksfFTgmv531DDKgBnHCyz84P6uLJkZOnoza9aiPKr4+BJZbcQ3flfwcHbSGj7F65KKgeDX3sW8
sQ0MpQv7i3aRVQD9HgFo99rKtE8MTnP8V1IHd9EEd0f9VwHL/aruqayYpS7CCAE702hbv3q+6quZ
N/hht+tn+TeKv6FfoS1y5hEQbmY4AtFAqxO1+mgeN0m82Pa4IsZbnN7LfGtozNXKnOPdguPAy8Dt
FVoPxKjeS4GI0cF7nUdUnRZt2uh2JSvJdsUCxtsnz5hGGCKj+b+0HMdz9I1RjrhQmvqN7/74dXnf
Aie9jVaE4NN2xyJc2mg3DyRLfUxwjxO/li7ti6ebAzigS8qRScWkpgAU6G/jqiGDK5t2Adse4YWq
QA3GgPIxzQYTiLbmZxcw+wCQeF7Ycw2D8e+sym12pYu2QFlhs4u/q6lKxUpjNsHNkAV1DbJEeETm
Keda3VjHoILUTCoP/NX4nlwVIKbFs5MtPjGwNb+AqyVRRokM1nzkaXf0EekvdZSX47mMx/k1X1iR
m+m4aDVphFL2Dw2dzYyN58XPGqFsxudatEmbLKiBIwWGktqjBF2cDOT/Ghiu27ZtRpAnbaoYVWgY
zy6oMTqrf6aHMheD8haZFZxBtSTZyt92N8euEQix58iL4F9kF8A6q80mqkp8n+NU0618mtWO3FpB
7Nh61oXAk9rkFMNaixpBcCRJZIzu3gG5BdCJwjebYwV2PeSoVTCe2KXbEQzh7RS/QALjOvimFWEQ
U+oUvAyIUuH7591Q2H4x//GkMH2yhhd39vlC5e40Nkb1W/fF9SPHY9lo6KorXDc//Tw/maLtjFlI
PH5j1KgnSEzNWOolINWAd3LQCwq40El4ZX93C6Q75n1oSjVrfzqSnWIrI/iE3pKm1+sjW3FegqI0
z0V9OdXlNYhICCebdnXLMgYASQ83QHHaoXigEdjIdEBXuRAAoSPOT0PS00RFxWaAls99pLkHTxyq
D3fh+5QlchqWq7090Tl+ZbHOy4QQZ5iX9XhJ0ZUijJ7DZwFQYWR95t9Ry7kC/0yOe4Z4nv2pVGRC
W6x7VjVzcfracg0NzRz/oCRswPmxGWdqum5TxfmCiqC+bkcGAcG7nC4+VCiW0KfqUPWHN1bBWnPp
2A9BiWiqmcUJpxePcbu+ilOBzpzTQ406u74WfnBD/76UGsbwLPiOxoMRWmwEJAjfoprx1c7rfAmJ
BymwwWTKjZNdxkyLCuswE2opRwGONs+YTB3GTQp10Xp3JtmukZvjtS91OSJJqnaLE7rrrucRWevP
8RijWRRNtGcjF5xR3qNMHY8b6B5k7VQfc+4ORheg7QJfG3y9BZONPNGxc/V6SY3kLzBgTqt2Vezz
u8cKBEJ0apYA6laEQokDa0wdPScf9AsftbxTR1hErX0mYwOxqKdzt728fNLDxwPSzXqs2cw7TYKI
2nonEI66Lj32vijoc6tMwUXFGynu9hxRgKrJG03sJyDCOq3XSoYAumnJ2ykza8hkTXRp4d7ICrr/
A0M8ZQMEwE+B8WEly4dEPwqQKMaBLe2O9heKLkgiz3wZMlMIJF5BIJ4rk7H3jfOLymTz2hUH6I60
aXq6mAoRB9MSzL1Btod4AciqvmVONw9xrvs3O/k4d9AyUtHZ4kkpnSVJVOLgRIwSHFvyNWwcW+1P
cR6PsFovOSjQfCqdIZ8aUc6b7GtvcJCICzqMaC0/1qErE6q5nXHUGR0ELuGN9YV3xkRyq0B29ewr
K/EAEanDgwCJkFA03zLxPWzg357QGPr+Q/DzYuAzwEzfDqyWhD86wM6CprCHBbMf7To+9t6Ff/iR
Gb5m42ArNuX8+cROeAhPg31mqh0h2M3nw5hlpmAGseKgXblZ4i+UaW5L3p8fYUJj+FAXr4akqaOA
2g6vs6DDQwNo8BYqplZeC07R+TWierPOyp+TLy6+c/r9pCuB32lWWwNsW9MoroalFx7MieIbHwzC
9C0kieQ+2wvXjmhYHZ4QSThnv/N4qfKCOrxHQ0e4wFUyspsqc+mLRqNYpFO3P2nlH/r3hDyc96WL
aajbhvYB0Hg22oB+PXpis/IWtWfp+b9nJJJ62xYvCgxe2RPI4bJRETEaWfARtJXssiFsTk+GserC
yc+dtgohhmrtEPbOPesoacBFwiKsWiF9xJ/ZZpvHBYiNrPSN3xcu1KfQT4vfZ5obT5xyXLUvF9Mm
fbPWId1VMNbsg1xvMMQJDjOB3LrsLETlAFGWIIspNsizoItsAOhZ3izxVbvQaUY802sDhqKabdEp
lycFl0KINeEtfvOcsDp7RbIEDzD+KVnjoPGlj2QAuw2c8heTEBdHKBOtYGzKsjXpRrCTa0WxNdDC
dZX3QCh0fCn3EXGiy6czydCz/66iwo/RuCJAXDEC9rkVCEA6pp8AvOq/VpMmO4sn2w5JCWjVodtv
H9rX0fYTehIw2k9288xuG5SLYOJaTKDY7kidIKF+m6YIUf1aNIM0qKOB4wIFvUCf3/wyCghpW+x3
a3b29W3idKvMoiws5wijw1MfwGdZZPdwtMJIRzCEXiwKX61AJhpyRjEhd/LHM8mITWDy9ftfoR7x
fyADQX+NeSDhkNqrw7QcEtHIC7XJG1PsGPs7KPqod334iLBMvV+PVJp2PfJBxuzfwTFAwRP42ORW
XLvGdCjZnORQcqzdnjQqybstqJ1u3bgM1bCe2ZLtGlHj6z+XHwWGh/RGGHOTaz9KCaM7+FgsWbGk
mc0jkjDrhb3loZeBEN6mRcK/TwpRF3yg4RDsQ8MTzIgbGMqa0xYONpif2c3XmEC8QH+QfA53RowR
jxBiC4bxAEznp/Yt0uQZmws8uiTVn7PYLIJPwFoSI/cYufeNgtsRghAVFSHhlYpjhEloxTdAhxWL
BaRal+0lmBcHu1vT2dgJMuZZMgwGvy8OgiK9aV4/3N7vDYbTgCLEqhyEWNI+PRHYyF+YWB/AGv+x
dkUvqJlgjzxLuFZCSH7g1o71wM38hZ/9u4o2Zxbd+gui64Yp0UDx3G1o5W/XLqOegAkUxzHPkjNm
t/f/n3VK41Hx92vdy9BE9nlpjfU8sUAh18H/cRDONYdIreB/BsFg9fP4oIgmj5pHEb+mbr9Ogwn/
+1T1VSxY/4zeWjeWYkgKNcGrOsfJwhy8ZLuJ6FwDw14yWInDjw/fAR7boD8kOt+v4vt6fQ8dmMA4
2zbov2cNTGRh+lEG4UTI5gRtxf3I/bzJ6cBN7PEzQZOtOpPrmRKKoy5lfV2r1bR6GkkbZyrlxtoQ
yC1r/l831btB4siMV2er8r5sgAL6uxOjFT35hQLMWYtIqVjv81hyIaG5U+KhU1MP9Lg/dfCOb/iz
kuYZVaGESMH9pgRN7YoX/CMBJXmWFZZX15WCEO9APyYKOVsw29XZA1bjCqB6miIxZMIHV9VXarA6
tt0Mc8nOrf5Z2pGIRscmk56tIQwEWbr+34ar9EyogZi134bubRgKi9SM6FC/AZ0bLT7RdxWQLnBw
vUe0yn+VxoAThUoL5EV17DlIhSu6qCyoAkjjaTjKDyF7M9caroVBd8RfoZphGbRJ7ijT058UKyaI
nPViaVVsGY0nivdGduIsWQZ1OIRV2lFSQF+IYdTPfL0NoUatiTfafz2Jvu0eb0GJRTChbegzQa+8
vIDgvXD7k1ZDyIRU9vl43cR1peaI/5GMOT7xZBTu7X7kI5zgYjJIUidnUJOjJccIhx0Q45Xdmnxy
U4hrlCiss+YSZhszD/wbP/cmAm9JMn7sTnTA+nKAcFaGsnt9He2j6OyuKTJ+hrKBQ6jSFvTGfGyQ
Xgn2z1FU6CaLbN3B3DKOPRNupln4BhtuNVNnmdc54zNOX39eptoAI+W69NGmb3XfLUiBGeKBx8OZ
4EKVIodwwuL82e0L4JlG4xu9/JuZ8eQ0csBt8/u8voiOcIaVzIZEMRH51I5omMmI6Td0VP02hZpd
etO+D2ZrI+1RsAaTK7/dm6UYsdQHpdxNuuovb2dlqeBOKgKi2Ipx0xreaM535WC2kfVyHRTsrW8z
YeHpmwPDl2sVf7fq2so5kZuxmnGfaIpEb8UkJhEucLzPdxcQcIjjr4T6mqahwhH+aVwEYAxIHcsI
gKF/eYN14xuyzgfRcjzTGBSqX9zB3m+BgWaHK2oVBj7CRGJYXvhfbo3Mqd0cxgeXXIfER1n5G44m
zfq0XAWQZoW0+PE3gg3Wams3Q4di1c1jNjcvr2N/xGIGz61H8keE5862Ky05pUYU9eCb3SpwHug/
2Ab7lRMM4fR+3oi6fUOg55TRaGRWkBfPaiG4f69kbskP6259WO/bn9CkgBhQ8FCcFSbiFRGZKZQC
n2eGtjmZquy2Ya1UxvJLGskgfW5vge+tWdKzjf1oSZRZXjEObZ4iGsBFslN13zrBBsKF2J5cf+ji
N9c+V93xR8I1NKx9Uhz0qPMqGCkeAbO8PMBCsC0M5thquN8S+DAx7gAM0sJy4n7Fu4hkgKZLnRc0
XfwYJIIsZRm41ZtQvtopLoYaHcw3x9+NH/dGHuWBgnIPXzXp/drvsaWOyKJZQBcL1KvJ4cNxID6f
kBy1PtRsh88FQWDVDZgspcxtJS92wLYvdBC+DHf0l3TucHPA12PZgVEeDYREWNJ3OLRavJnfskhy
w8oaPZ/hr3JI/PEhAQHPymX+AGVP6HllizgjSJpPqKBPMSrpFcH9spIolbPJnLRKrb6ttxuHEWVX
ZDXnxtOZ364+YrlliHa39D7i0eJZz1qVSrw6J/F/ivJSKmy6TIgSxu4w94+HI2Oulhhozrogl9pi
5cg6GFYlM69MfNCfA1IKYpx1EyVqJfVLpjAW2gLvwtQXTsvIfAQKNXizKLdH9WEDUnjTPRcHM8sR
AOj2RVVfq+r/SFCSCxrqxT/PhUUZunLJCPygsHo823c9xLy73qZ6bwaA/+XgNPZtq4iUGiITy0d8
JjsGUQPj2HnYb+PpP9icU3uRTcx1/GrgvKTWMhiI3l4CMOaY+MqtGXad8pAyuT8/A6OElK4p8Xgc
bCq2GLYRiu4E4LSEn4oYRCsqavW6IFCTry00QSyxs/xzEgRmgRHd9gKpgRm2DWRosDbYPY0JkYrE
VPDOREJ2FV5paS6VSdI4NoLsWwvAFaGDYzhl0yGv0dIKBR0wFWvKC6mp2AZFYoy+qlkMLsmMUI+i
w6FvvPaiA08Z6NvSU5bEMAKvDGINHODxwnh+BavWSjX6OLyugkBIQ9HXvjVNTJgEsTZsJ2Y0QG0g
uA8I006EEkDFAFJ/4oFW1BqTW7LxweRLt0Ej8IHteoyZE1YZa5q5XRiJnsAb23rukVQ0sLy257h3
+ChCO++z123t0zvul0TKzlt/9FmVHQrxHlVjLhkuyiRvFDtd6qP7JVx6nhm38sKdcSvxT45+1nlM
p139RiYWERuv/gZ8IIJh4EgZA8c4m21pw2LZ53t/ENU6D7C4HIx3pvvloA8S0bSvNtM2lu5bNtL9
j5osccuxSGmCxLk+kZjp4dDsEoRFNXGq1OKOjCUajnxyAe4bfJ3xbIGOsewwu7T7ivfWb5T2MSX3
e9b5+ya6gV9jtQWiZPpHbTvpSzPH3EP9JXFUdDbiNT4QCHiyfvD6+GcmNX+Fjgl7ep4jxFLftAG0
x/4HzXyJT2CF68h4OxB2dSKh5qHL48tWY3M4kXvO0w93mJrTywLoLVFy0tQ60IlbSWkNgnkB6vpR
02Ko337uPKDhIsj/mYvkLRwyVZGi2GI6DXUn/USMcC4JVMx8HR+QQsajPCkFXsq5lLv8xLR8uIik
+JpXbJrwMBHdsUX2672RJSf+rVkEjCyC3O9MOI7PLLpMd9+eC30A1e6bToypkphseydUUJvNCgnl
2vbTQ+89gTWLKlHsl300v5djBHtno6Qmn7f78fv90zHPXSZ0YA1q2nR8zMDtp9Dz4+IGHhsbYDWq
FA0QIssmhYcMRfUsy+SSSjRLxYCEB9DGLQomUpdNLCN5V2qyumhvl2Vo9jab+XYotT8PRDn+xo1S
5GO87JXz0Ri/8YNHyjpKpkqe/0yW70WCCILAPwHLlxNB1W6pUYE/zNDJS7ptXIDypL1XRMp35mdK
Im9RYcVy9eVGkA5v2BBGqDbvtXWhgdd7dUujADZSL4WB+vZHhVI4oD/qacelAiULJfRYxFCyPTW4
KStkQIEBUKjGbUbbC98DbXoU0xSh+ouYMg62VwhT+TKzgcQ2JRLJkAFweIRdZcHCdc3B8XXheclz
w9QKeIVTqcWfww3PZ6KN9y/nhMhkpNCZIqyPiQjcLUIQhqZeHbpu70b6CD7oEjZGOHJI5cnS9ena
VYCLfMfQvuOGvTLUUOkYTEJY38elDtTEy+2AeJUUyJDYKH6CW6EqaqWTByQr+xKEKmvkt+szdTM+
UASgCwN61T7/7Xrb7bh4x/gNe0eAyEUG/SXELf+5dj4tgrDqi8gMld9+w55+Wpp5xQYRXQV4Ozbb
sboD67JOgU2cNchq3TymtN2r8giW6Q6nmYml0kFsk60fbINhhqt/BR+LUWfWKvoqMaSMt9eLuBkT
f2SEKxHTH/9IyXNmelpZ6dVFP9lkeOIFz4yE1WW02hGIpy/1mdg8HGR62pcKqjXCvmVrlJCU0JIC
RU6tLqoZrY6fZFF2ndLQ+tNZiypxWKpbdqT1f4gnNUFAatXWNUelrX/roFsO+bdBE2JV57NSVzQR
1JxV7Se6mr97/eurXJA6loTRj2zoMLE2jEnGJoKLAujqzdu2RN87Sy0LdKHfajmvkM5tGLLj2pGd
Wv9gYecll+JwcjA4Cuzd4tjbUvNMYGucsaN3HE/vJK27oCEioPo9kB0qchIglZE8/k71iUQtfcQh
Z4SZsOn65Rypc8VS1woS8Ue8O+sjvroWtbla3HaA6HT5G3F3qv7PoY/BzLGGoEywoNkiD+tcET2E
xWQV9SkFV0vsRmghQj0/blcdQFEtWkZrCFQPE88m2WX9Deimv8ynam29N1vfW8ej0N3Rm5xLIYla
KLPiWaSJpNjXbTRAYiAEbGAiecfuVteJRRBn/UyVI0laDMlK99AWZP/sr4XR7cud9n8s+M5CdKty
itStBfBvfBJlEIR55RJt7MmQZIwLN8cwi++MW8jPAkGYcky9oPAeLxWZMGlB6ldeYQgmo6QTZq1e
3fWcu2N63GwkBU/TIx8Vk5VqwEcqGsheP3g1iKwXGX38LH+xLmmI54unnIeeF1tvzDQ2Uei2tBQZ
hsEnbkReUZtSwuo0QEzXlDuUW4sfHPfeO0YxDnoGMK7o1pr4xoJLWKlfILoApds2nTzv0XfrzGrV
dqqoW0swcI7osxa5pyW+u+xnMa0yLVDEGFJOG4UCDepPoUy62OwMGm9uNHLzdLAQfH2qSQVEZSeQ
7Va+uIqKOvgQ7mZiIFOjAev9JeYrM425wnGIhrz3U7EzCsueyrh/I86zSbLBGGV5Lp+ZqTgDoHaY
PU/GPh4XgCWKbJn94ZMJyFvLY5oAU/TfYOI64fnDeaxnW24Ql6RXEGgIhClzgmMNpoiZCUX2Q+JM
OYDK9t7J3HW9MT4Vk38pBGZx9DCurk/eyWCwb3MwYPcfFObuej1YHEU4uwf7Q8Mmx26+8mOWEXww
pMweGj7pLoRJ0HxpM4xg2u6FC+ZE/AjGR21QfqChNb1vsHs9JKAAYxqhap8MThP4AXR9mHkrtgwI
yK37CPmg5imVlWBDjdfcW/rNllo5OWZggjes2gXDf53tJui60yw2sYm4mU2BCgcWRtHWbEVLi/VR
Y8JuC3R5L/xAsB0c4S4RGKOnT7Txz1tIf8w6m6ZOLG5fqSa2Dwpy4tuxu0eTtsCuinmKJB5cQ8SG
5WlP99BDPTZQUO967BCyttuQbD6EKpLzpbHkwLy1wmKrU1Yv7CQsXP/lsJ0FQG9J9I6IHdzU9lXQ
r5wP9TF6B826KrtJboT70ggqBr42AazNdE2rC9HYDEjpY9VJwOMfqZSkOVfsDl2FcjOUae0xWsOO
qGV4oMZf9vItzfqb0uE+EOFGK1L3iZ3kU5I0FP6PiFbrFND+2R5G6sZ08GEEWrkzVflyF9M/+9sD
XY8qTCKXZ1dR4muAaBYkAJI1GWTQe9Y5midHcZT0RJhocHdJa3o5OBl68CopEMkUxOwg+t6ixxAx
ReQV+zCPJSrOgjui/gc47ZHLmAgTcaKrdwaNyhr1fD8eQy11mMNZE0v4PtXXD2plqNKPc9SvXxmN
6mk4xfDlmgjRVv2As3CP7J85viFl2XtbZhqcQ3z7vOV4qOOR1jps1eCgtknpKuiMZ3nfnExK25jN
Flzp3rl3eSoZI2YS2AEL+VDrJh9mLAyjY3y7s6cnlVe9PFNLNHQjR89tfkioYQPQuutZ1eCDVRSt
0yOw1dQWG4pU40wdN0y2I1EbktZyIMFrsXFKq0dvrL1FwJHrLGaX3SSkN936C3J6NXj8XVO3JutR
scPypDCbONRPS6Ne0pE3adZyK2noeH+P77qqQ8ttcfe2PtaHxBSiLTB9KmA8W7ZT+PgY3iuEWw63
eRNiniHJHVomlufW179eWTLL8o+iHAaLDiUIsQABIe8uk03Jagr/kVdGnJRXHSfdcV2DjQARsG7E
4KowVYDmaaSh9EwJ1x5qZKf14bWD528r6zLHAgtVDfa2eBVKOCeT/0ATiK6Q+PdtNo8yOoeZ/uWV
VIMaDYRJX7pZkYIzk8/xsa/uRjC4nlNbNrh5S0CmTYIARfeYsvzOblI6bypZ/63ZC+/mWz5ye5QS
F7SvZlFjowaCuU0pfQzYaQpu+zcCbAHJgn+iFItS1fmSPll02VowN8I/9kW6CHIoX28hkxDEgwG2
r7EFGDNVpPeC3KxFJnaYv02eNwuTPcRpdlraU9IC2YxW4MZ2ngY0oqQ19SFqq9m6LFjEhMO3ujLD
U/CMwfdmpHuYvuVGQA2uMFjf6ZXD5XscxMLG9xu16gJHo0F0wKaioQ6AscMXsE6b2A+E61XCwbcf
egtzvFT8x6Naz2iqkVojc9WlD0CsAbPL36z51nyQnTleUUKRCrnBMU+vm/BncjiX6VGpKK4iOAJO
uMamu1dhWtJbXhH66hmMPkNVfHJGwPo001hh9uXko9LM6n5Wq/B580+zIGSnh29KZMA5cGRB7Ylx
31Fswlpw3YfHl0Uo4/ddEz+LwoJruyXzAFYoy+GvHUPw+6fCdND3Ba9RyRcGT02/pkg3Pf4hqYmx
Zb06JjkSKSHJbRWh5aqrMAkLZRShrrrJiTfQWSwRXRfVfIWtfyZkVaKf9n6LHTUJpfLJdaxOadzI
60v2NO+h0f/8Lrz0JeNmt7g8VKeDO/uL3hPKTyJKjR/NCJ2DEXYntNH5s070rV+w7p8t768+2XLM
xP7HZ/mgkq48IW7hNdrpMXAYPiOmbLJUVfNc/DjyaytJMvcavbb/EmXdRXB4KuaCSAqrsomHfSrN
+oMQ4nWslNF4cUJaftcJsnhdzsnm7NrvBDjYNbCla8aQ7jMRxl3DoEcsMjdop3fKSi9LofnEYpi0
aeUPYvnxw+blXuzbc35ZSX7agb1PRnQ8GRfUEP+84QAqyM6O+B+/EkB9HslqcnDaRIFfs2iXCs7B
SbbYXyd75WU+5xLD4DsDxH37mkApESz+06vT9p4PIwNBzHmRr+OXe30l/ckQp+Frfr1Oue/xTen4
C3dYJnZUzNZg4C32/exBPvycXRZRdTiJwfP0oPWScRCCdkU94MLnn74OImA5YkTsuTUmcw3gapqa
aehlqhmfHnT4Q45M9zjfkFIqkPf4wBlI+K94ob9ZAWztgCwc+U+/BOIU1Q/ewC4xZWvDMJNunqid
SdDZxuS/uK8H/gZBlQHuNNVUjGh/2Q0OlJRsc2YK2ylUGB5FOrDIhvOYl/5c9e9eSKCAR+j/s+rN
49yv2bZnVc5CPfa8RI7Rm3dsz0ctxAxZxSmVrpcac6jVBYhyEIXFtgi1SxCco/bAuz9vEpYKb2ap
PPxd2hX3Nfg3Ze/rRi7kewGOwm9xynH9OItcvUitrmMSMds7PD0anFOpHspIm/X7I/u6P/j7Kly4
BLDsv3HB8zLJTzRDvoRVuz9e6iDZHJlIlNPPktMpP/srQnI2J8/1pchK6Pup3YE3wzoVWTaHMoeY
Ll9/M1I5343pQEqAurvYv7NGJNzmeMdm1p0pf/IYtO9SE7c6s8pomsY7pHgOHyKvGOnIVA96svRY
krAkPmAIWpOaQu9RWEdyyJc9TO9pnBzY/9bCeuWRBGlplEOYG2dspU3IFFkuw8S9vIGNf+Wz0j19
qRJpZ2xog2yWiPyVQzQ/r0EjV2Y5Kh07uOwewS2vEq1E0WDz/Bq8kHSSHVdYl0Elnp/iWdYIz8Ju
dx/RhxrLNBEp+umopzZFcKcpdbRMMipgtdxuYGUAl9nPprYijfq5BkBedPeUSbUjm6pMXqgZ3EFM
uRXlxZl2B56fLDw8DyfQuWftVVq7khO/s7sIkUGqS9sfy46ImN3UmhOFLawnokRJ/sOHKmpabkYP
lNIszTKlGYeUtrbabC6M28MDyZ02XFCcWHldP4ODPImpQovezluYZcJsQUfgZzGntzJ934bnZmWc
4NnFqKHLScOaUwFIw1y7nW7Ogg+j9tdClDZqYBEAxoIFfmhzTYc4JcYpIzNHVB2YqzCmOuc8Ig+t
pQyHXw4cv2RJofvn4nVSTPgboNLp/ygdLXZYbk9EcuD2HwVfhqj9Uh6MQ4xVDPWp2g7ZNgbD1/Hs
ktdOd/qSagliFmHRJjKBvXHYzT73qrPVivcvmUHyJ7vEhjrz5wyWm9PfNsRlxv09uWtfyWi9qWZe
9Fw/uF5iO8RzF0mtyNCh1rFNEDKuCkKMHfv2wBj0fjsynn53viwCP2tBfsvFh+b1nAV0qDb/FkeB
JV/uj+RzMmH9vSNbMVOJHRQIFfSKFe5gDX/9pgAiHgFZyeerksT6gOu1J8rEtJbRM9gZD+v5rXyb
Bv+zymhSzYyqiDie7VjHgR2XTqPWNmeIbp2HEiV2tM+A2TRtiDZukEGtLrWpnx2HK0BFPWqDtyBC
KfIyeSaK9CZLhcQS76gITeJky+F8PYzx3NaiOg6q+k1HFWDAdGZOMX9oh4TAgoXKMVzB0mEwxZTw
TUb2c2K/8DidwVUg5KkjROENJq2Qyk0+Z0LeK0VXSVgYruIaUY7Gef/1FIK7XJitX01j2KEhRjzB
WqKbabE8P1tACTg9EPuLbf+25lHP0WHYXuUy9ICW++zXbx42mJ7MhIqFb0cZymid8wFnCiCL5DBN
gSGUdWi90AW2OG8WTVaiDzHFcYgTP4w0HjduQtKsW5oC/1LB6Dj3Fvk1rr+RllvgZWJPBciy0OhW
wp4oak4Xz/T+rm0Df6uzBUrLYJg9HOIabDdxG75d28QdJDNkNOYI1HITRfxYgoEJsVJTyFo8KjrM
388J8T7JOTC7mdjHFRSLJ3job9HtdTTh1r1fVcutgseKKxEYaiW60XLgMnerFUee399xAfcltLpP
zo+42+/UOnMBO/gZKOeS3tkIt7PhRvKuofVFfeE9bwdCPwFJpzOG1K1LuFY05ppNV+jqQXcYFVOi
A0vZ12sAdIy2egYC7m4z4528NqOBpTHkn4GSQbQ8n58fra0tUEUaNhUKZK1tUYvxdLT5U7gLJOfg
yhsqtf6aVG5ZsbD06Swm8VXEmTtj0sJexKQtX3nix7ORAEL7NRfTtiB2RDi9UjVTrU3JXyF4X08y
ttHZ2aksV6TpKxDwhH7QAL9XmjoyymtsIo91sdsf8JLOg5Rpse2IvJtSrFry+5jrp0MPT1TLL3d3
gA5XQsqRubwgz3BmCnmQudQbd5w04ic7+XBkaT3GhOyDxqyV8xwTnpCUBwiEfUeOY9jmo9WPSlBS
aPo4esBFiwfnKiovaE4t+ysTfUoW0XzO6WvivDl1LRFx9y9eNJWwyASV2YgISY4MwoDWdZgd+St8
LVEbGSisnTJsF55CvpBQjnnMv7B9vrReIIDRt4dGoS0bmhBJ71ste3MwtqY5GrmdZArMlRJfEEGs
oG5GQD0yGRy3GYfBIkXG6+z7bOCN757cMu9DuJozc2YLK7GgFjtANX29cLK4oJPzM5lYHLAS718D
e0XnPT0hTEO+43UB5zff4i4LsCmmVk4r8VPhLq379dqldOmuNHxHz9f3fcrCUNTyZ1+nOuHat/gk
ZwzbgD5rNaSnUzAMeosUSXKMpnHPkqiERpKpJfLjuyt+XqXE3AoDk4QKjcZEybKYucEzf+o+SiP+
RFG5MgHNHMvZY0XQckX2kfJokez4utaJvZliZuHgFO4RIoUdtv2Pti13t7ksuf+xykfeyDbmEbjq
pauJcEX3HwqhvNDkmmmYoeVh9quXtu5jrvKIvK7ECi+g0Y7D2Ot/i4mKlvoPdvw2R/hDmbNzTjbV
42RFD7SRHw+Ko3wZG60+jXTYifHgns5VlJiPJoKn3imCmtWLi0MsbBvkwuRkOa7+Aeo8hqXlTQMY
l9FzSdxgjHYkxA1gYZoqOyy+xQ0DuK7pkf9e7dqwLpTnCSr47P8Jdd1zPPlevYlwUmPkhZosj9nY
wzOESYQ2EnlsUaCntlznYPwId6reCVAQa6/KeXUVYgPuzvrk9WsQjADCKxa20WSC8I2RtfHauudR
pxyL+AFqw0LpdHkV9/a9gMIssSX3GOgYvly4uHbTrHuh1qIPd9VWS86ra4zu3VKM0Cwxskrl7MH/
sj3j4PMyvzdnvloP2g6sZAcyVYp+jk7/VQzsn6uzLgU18dLoIb7PrgmsjOIAxI1MHS6uU4f1K9yu
B+okHKATKHPw1DT2FoO9BVJ/bmwHibcVqQP0kn20hvBHxTeRvyf64WdSBXm73luq6rZQy+46oeBx
TUnB4A9cHsEMiyFcC9EorAwE0qbebpp4MoPb3bD7pO/Zz/ecWMeT2Lg+rF0FP5WB9VZ1/pujQGev
WoWV+FYzhy6Aatdc57WvwLxnJ+a8IjXETeFnWJ/7JDqzgcK9ZaTGav/0fa8rgHuP8O4X0whzeIFm
Z0hJ5It7LtDWWZbhpyp9ujIIsWEZSNrTYTeUeW2rhhZFOS3v0apmWWmREB2Sn3vspWrrBs9nqVBT
mkYS7/aSBFH9bc47bxMZdI7H88jMXaKBq/phQ8rJSg1Qp+QvV2M+kbXDLt/o9q9Auce8hBxxZ+yx
HBwUHk9hePEz8wjpxKGlQYNefz+mGoYDx9jp1XmqFfb2UBqTJtKXE9V6zzdzRBAGP8LhH6hf4CLR
OWmZP+nCplW6ocq9iU64VilmjRF/jEyAL1pYa8/EvcrMo40mFnaAaUxgPxM7wMSvWnMFl1TCF9/J
fmGqiG7zP5w8RKqWlipOBCS4PAtLSvTjeEwRa3tFWgIZiA6MWPWQ+Dcff2r0xW4hHmJ4ucjHlKGb
GZMJVTWyhI+ONluI1uFYi448u9WT2l4QDpbv36SLcXV7DMZZW0JacU9EI2DDeZCZM5fBkNkp8kBy
/zz5qtFUpHh5aB57rCu2f7QY6/Y7rIXzVF53EUVGi4qCd4iNc6l1Zrdj8wAOS65TDpl2ktl+g6oZ
q92YqSmY0L+yzaVP1IpxZIDbTwDCPAbsV8gj8fDebH8AInBl7gR5dz2lwiDkLjEDVaLuPkL0c5o8
IaKlozo0tH44qw6q4qziMWQHOeVOCLAlHvnd3rh2UWTUGOxUnZFn2LHXyKZ1cU5VAXx0h3ybsa05
/uJCpX6LfcO+MYt8sgg22hB9KmIgbjnw5BZviDl0RBgHHC8b8qc0oh2Fwa0aRHILMZYEh9Bb55LC
/lccQJpbTRp44dQma5Of2HiY2zQNyfaDzcwkavTcAYXMdIMG6VTQVfvjoQl05OakBs/1MG6n3YWG
tZX/9zW1GnbbY8Ggdf0Pr/wrqVevdfsAMI3Po/KLXRlAybUWbk0MGv/Y4HidCSRIXg5lKwhW6xJ1
GRKxgBZzZP2uWQ4LHA2EL4bnNcYClFMN4K11XjZcTs42ZFxgs3Zlx3bdXefGNRRuaMgXZ2YdXb+T
7lj4FYgGB9Xj0buF5ajAch4ZP2zFby0Kwaug1RMa5fZvr+DZxaliol3+WO8XIeagpzbXHE66jaiy
JF9k96nPAqsRWJm4IQ3I0ooobBRvFYsD5n2BOJl4Mc0FEVVh8pUl7bBzBGDfliSv9Jl+c1Jcz4/E
kU0vhWq/RiKxblfsoTBcurnSCtb7wdkY7ddIFHCyNV7WEQYPI3MvlBN4dXLrAaQFQDdmO6gGLpBP
+5HnJqquBfh37hJgrspCf/x4tQ4nTt32cowkproJv1ECo94otKU+eLCCPVVv+AEDG5mh0ED0Vcja
Tdwuv6vrGjaziEhMKhqBGpo8nXlStfchI3eGABPs6DCim1G8+3heTal5OtN8X23ES7ipxgiZsfdZ
T9BZw8J8EYtiIWZ4k/SI5OXw/ZXh4yi/jAGM5+eRB8/7lxRvfBY2sFxrCPYQxXDfKkgLFSWfa72E
J4eeqwgqUV641DIbY0sgH93CXalMRziV9wiSodlC9LXajBQLD/JAhnCT2Vf+fjH4uPRbbiUYdNqy
JLbc/+vYYzM6YAJfPOrkkZnol+3ebETHBw3+npkYjre1Bl1zzJLCToM/MP26Zp+1UMZOQhF/xJzw
goo/9br5+tLNckuQwzfnORo278uP3Ziz7HSAbaG/73f1dAVSupMq7WPgCRCtfgYdftodAkyEe6Ms
Ok02D+/EVeioiS6+JPNGnWuIWsTYylFelL4wFrKAaoP20MQCQc0sfnzq6rqkugePCZCdaW6jfMta
Q5Qz6ucbaEQfgA8kzfgP2DNYgQHUU6o6JaVoRgvm35qIYXuSstKcYvdzgK/iY+n0kcOV9326cKgx
3Ao7a8gPSHSNsryv7jkoAjQ8chhXZgTeNiEdxxZNN3Dfxs4t9dMPg/cZkOscTlg8VI89AaTSCdTa
lIfGK5amWUwEC06exMz07P3RrQU67KdYDzI88XN/20oTZZ4ChQjWJxXrC7BYYxA44V6AjCtDYQMJ
0jwFEOG1qFggXh/MetsyDxYoRqCeyWzETXFrhnbzU/vqin13Bgr7LgoZMkLg5g5QhT2edW4HCOfa
b14hokoH6TANufNHn81XlrIY565SLJAKAsyoWeagi7mB6XfP+x/E764FJHYY4CCDUBXtoBdslNYd
+pkqt0FKwMrREO+cgsepf0G/A5f6CWW6+//6wuyStdt+YphPctbPdnQNcHrBJJIWmuwx1GZ+AHf/
V7Qa9ScH5+d5YABCKwhCG5JV+JrRYEQKYi7+Ck39VFEZAk0Aq8e1Bx+POfOrZv+KxvkCXzyXqx02
zMpc8H2/GyVd+Dz6qtCmep6SmoYXRU0G+iD8vWNFFRo33sWEZY5xC1MMLTRZTtQCqnRpllsXAuFX
MTp2AD51nKfkwiuWSWfe9UrXLPwQXdUvQSOzyFaxeOuY90kcGwRonzP/Y2teqVY8cqAw6X5SyNlX
EKnXWx5DRBoYh3H0ahGB02VhZZA/sLfYZq62uKF4yosXvlT2DtbfTgBNM9RTm/yd++qeVfhjSzfL
UPbbu9VZbdfA06QmBRuGgM4rZtCDgudGl67zwFPo2RxInUbvxMDB9Kn1p2Qq08cxJj5rk8sQFmze
FVM3Y6mPgMM2vZ9KQgC9EjLz6FpdAFEA1d5PDC1fH6nt83MHqi9pDwmzBIX4bRJYAGfN9IJPuERf
RdJ1PRwIJUv8GWjoPaQevCqsx9eB85+UR+TVdeOCF/taAHUTcjpH+JZL8+Lm7yFUOOhMZaa6jG2i
UNlH53T44cUNjCZzYQc7SFAOvqFVsbkeSr+NoJh6J+y9qrSPzale7A7vZldhhgDZ0xVROb4tLXVI
GPl05VRkU28bSTF/VjMzakpBZospjc5BXtia1m/g2ORFu6lggkb7BsgNUFQpmiwWAG+foYbElNEA
HtS3AidFk0/4vpfXpFapRverdXdZL6biy5M6IwpKDkaCWgPDc97Lx2/4fhw0RA9l3oHgTO8HXtRG
XmxOtgNnM4WREWE8Bn6vBEhouB+/dUiYGCYOg5DolP8ze8/OIAClpE7i5KROrIzi6T0MRCduOM8v
mYezcdnDfHMzf7/K9gBRezZX61wiD49RkF9gxbqvk7S1oboF1yzR4N3on4IsyATZJy4bY+18DnUE
uUVcUiloeD3lWr/2nmsT4DbQXMJokVUkMdZaJt4YX5v/OApOKqBEf8OXz5Cym+LxPNeWew5hLBLg
2QJgrHOpddR+8KgevG/XGBDlCZ9vtDMQlx3j4H4Bx0vyzb6ldfH0LJaLhws/WgqjuMDB5fsM6CBs
A9qit8nfTJx3Bo4ygiMgP/qqraPxipDEkchZcJCRLzXjvBccYrbY8J2BIvKGoFBQTfDDK2aAbtXt
Ai+gs5I8tJqWfo0PgDuDsKM+9qLKCt9AHLtH57AgzotXj2HtKDUUWUKYjQcnkLptYQGrt5KOd0Id
j2fv4mu9AOQ6WSXQM9+ma5Jx3YRe94q2TwtSyxJJhsPB+O4jARMP5V2r8/RNHZp1XPY46KCTVdk2
Zurs9rhnhDThw/oUF6nv82duKirAZA9HA3FZsBtxbE6pKcmo5SPWqsWpoPcxWZVNMjJmlu/G4FYG
Lj7U3E+rjfpsOXkOHPqqddoS5queQSS6QiWxFTqBp6A5FVJQqvXu+o8ACf9yGPcRoLmQs5u4hS8u
dUO0SmzT/fVyTErkrLI6Pnp6Tdj88Wzxx72xraLjteUrKp6VdNIUhQzjx8flNdp2Y6okYvNBBn+S
Njsr1GtwR/THmHMUHPIf5PgHUCrKLODXCsVGQQBl82blRNuPMZUzSxTdGEbAPftMpKyw1eYYF3lg
lDgXq3DmpT1pKgP4arG6WwGUV8GUJ4sodX/YGcQ9Ca5LEjRd7bLh74HWTBxgrfITrWRJ8eQdPvEH
Z7PMEgMOh5bjwO8z3B4OhZyF23Ufk1taU467dxJY5zfjJNvAhrDygDvuu8z9pfYa8xHjjdSmqbke
v3smj6v1RHJNmEMu6Et5aPuBBfzv//4g95yNeDgnfL9So9SvRwZgg2VUbKGUUo6EIoAqe9eke4Jj
G4dEPDVGC+mFQtOiAfOuoGVrpCwVVrqnGtuORikajXXkj8uyrIW1mY4+HiFfhBECx+aFOmob2Y3M
ZwT43dgmdb9T2rx3IqLaWIrtkGGfaEbUj4HrS5gFUCJlRaSDKYvxt7XLAe9s8Qnr+h324bZmVZZg
GGBYEtpfEBAaaviQcj73ksMGf/pUOZVHBCLV4jqpZvLr6CjQmE5pdvrnqlnw5RJgOWp31V+cSz93
iDbvBrLl07IEvN3qF+R/73Wp2Cj5U5lVO8cfVxGtFpMoBExPrC4ZWPDIksndv2YbgZEtKUIn3zUv
WAwV/V0wWtyYuAdt/61vdrINO9U1mrgYAiveJvX+H9HKzDDhDtd9P1g46NGNzTMiAtyx2F6CGbtI
agD9DQKlGC07d4tVXguqup4q45T4P4ahNBn3tIDNr0XWiGtXfks9uQOBwEw+BHMq7nyWb+/dwe9E
lVoriw6uHNYrj8peJLBY6TXbQRTGbrOu5ienxkfGn6W6G+xP2NaCTI22B8KMrVITm7LMNCCSoWg6
3RdWZoc/IdDzidTZhMN18Y4gQZeCT5o7QpiHjtO9ot4ZPuPVnQarRNQcuvUZgyWfNAvN40vKYJqc
8Bc7vfkBB89vjdaDPKHu7v6aZHofecGpbJKnn+oh0n4s0Lf1TGRMB+KnvhQg8HrzYCCjhpdKHakD
VK9ILaHo4tD31XfAveBF1ovCk8rml+PUKMLNYfEf4bPmUYM6WNfOk/7N3kLzxJsEmO+gXwQSvHE9
6nn02acZ+0vT2R3NuIZQZVecO8L6/YS4+YkcnXqjdRt9R5eNZNAK3DLZtzcnHOe9TNLPeBMN0pYJ
6xs1UMm9/Ssx2sATHSA+tr0e+uTfAM8h6Lr0pGKdg3/F28uJ3d6lGnbk/K+5Y6g5WDEw8icBRhKc
QfJe1g6jlgWKcixVFtCbgZXyT7BsONuEbXLhI7+0SN/6dZATwxvycj1mOs7umpLB3veDaZSbTgFW
XBlHQk6TCCp/2Xevlij3QfQOjvOS35O1wnf9xcJNvRiGMKGUdvj78JVlp3X6tiYZal5RPM2OGBvx
N+paagqtlnLxsM21wMuARwMIIzaJ8M34he+dnOEykBSVn+f+NOr+/0V18fAj05KuM+DG2H/0GJkC
u32CD2rPeMZvoFnp6RBJZ040DsOKzW9sZSlk0H2rdCOHQmEzUAuWlm++1Gyy35sbSs9SeVxOp6j3
8F8WAwGAkn/8BWIPsEPaiXBdSZTND9frk0EjBYRgQBRvLT1QigqLvq3XGgZ+UqNnnlB76PA6z4/s
nCBZjnDyEFTFCffljNbLU6mbxo0C6XoZroFyhRnLSzmppkdT7nu4KG6tBzuD6tv7qk8CVoJ8zg9F
lo0qGxpGvThqjZIJzK7z9eGk3H6RAcBH5MZ0AuHunLNW+eRpmQ6dWN6UAKuM4TcP+Vg7HAkGJoe7
ZvqWnFvNFu5GWvVNfojxWZa60iSGkzJMMvmJxeFGZagkd0HUGZjncepSfALjjvOKT7YHMnM+opRS
U2xqplE4Tk1BLsHTSNIZgmdd4iwxiZxh7RcBELJyxG5nT1kqybbOWwibUcZBzvRZvVqmR4zXCNp/
Ok9r6IkWz3QtqderJ8RNsIuHup1oU07o/DK+xhQSbtcgOG4qqjyQr6/oTjc0DIapbs2RepZmwO+g
MC+tl70UTkWY2CW7xzMlnrPz5ZqmLmuzxsU2Ji4pbr1LG+N4Mg8ubDPM95H7pgmtsiQhYVXjzt7p
MTqoYkFrtJ9a5bcULl1cZp4y0lwbPcXaht/1DBYaF9/cFTlhYIuLVOkUwMXubSYUOnvgqYFr2soN
mdu663nhDlAmI8C8IVQ7yEyECmWoNIYE20zFxIieRN457eqEoB+UxnCoWpIjsRmQo1l97S1nszAB
rnXqvgq4yujZPaLMpsKje/PmRJzSHLn0Q/wTv/3C32F37U4+X6Lwu/nyfaQS/9sm2PNuVmxlNngo
KHyAsjd3emZERs4D4JkU6ED+brbk4tz6QleW8zZGB+v0YyvaFwpdTD/XXLPr+Zer9qRTWSz0szsk
zDClL7f1Y+CZvs1WSpkdF6viAUyVvc05dw9MtYZiXodU1f3UW8qnqhGK9k1RKlcwAEqsSzRRIoaQ
fJ0DVHZnGeavX7qpmCfmeZ0DCSpjPJRyt6wnLZ5IB+fXFdrAV4EoRuaYHUmfUwDD/3+S7+xzMZtt
wuPpyXYGOnRSlez1y7FHo9AfwM5S1TvjJllSkiJZ6wu0EsJ8wZTsDy5vCOPKdhPLhLvQe37ToSk+
gbTtLE62/95qFVy/+88xxm8i450gEj1VFLOWc6uBmeB778dHUejXGylWWChmIa3Er0gny3RWRVxf
h4HROduj9JRnior4Vb+0gjeXpkJwT/QYA7S/NVv5daLI0XesDt0KJaiQTH2t8DLhJXmADo9jEMkw
GeEJhP+HtcOfsqLKsr4PTbQY9wuRngjbZMY4DdTCgtdsVH8KnZuvLT2eK82A47+Vw6WNkgXKWd4n
6J7VzltPijGfZuomn+FlSV18WgH0KOGIrHvcu9eI3OddnCDNUGjbRXhRUvCsYGf6F6F+LizHWHgA
1orA8rgePIwdw6jxI0X3ElijK1JAOySFY3SPW/6KMF9G7In7hL0i0hyi5XCqGrbBtK8rKmbbUlA/
Kijd2tDQFIcRlIKgTIaG9FiId+2JavqoR17h5s3FEhMsuAzQ0GX0i6EYPIwtyvDZuPNQsaji9+uI
HCS6wvZuucYQwK9fyIoIAHv9Dnw6GtPfa8PAIAEVGvAT6xt0M8YKmqO3Yw8FUytwRnDpS1OPuJiy
fsU7SZi+gBVJb7Gr4UJ/p9I/lbk7+xuVL+SMX84trLBcng+7KwnUVVz9O2ApreTPZtUbO8kqedq8
E9tAZkhMOu3Oe5m0jX+MZczsZpzj1U6hz+rYzPPDsIKvigv74OkXFXpVBbBmiUMmCLo10MemJsPi
J9o891H+XUIR07VFCB5BY3yTiYmh85LWEk9FSgFQ144PoYRZ52h2UeXBZUDDV6UgV//6AQEaA+Ad
nBw7O0mgBbBj7W5QGfp2XmmBQJ7X2NW/BmXWyWjL1meI3QOdYttoSe2WuwyDBoTbsibegRnIJxju
C4NXHpM+RuZTtYpHYMyrbPBV2Ce0m+023+yHZSQmjLifcFjs591BE26uP7NIRvLFEmWcZ/e2qTn+
sbg+0Kt7iVugYkzOOq294/jwCslNMbf6O5bZipxM1rnqWmQdQvyYIxfYuH8WMR/WIEgOc39NttOa
Kaxtd3gnHwsTz0aUqLTwjoWPd6iWpXlkk0X9IKBjgawCIWovFRxzC/6RZ38QQyjM4ky4daY/nLRY
5Etm4BhT7atySqsMnqRbco5zSIqbqryEPQt1z5QUCgs2QccRidSrItOoka86xWRiTrxxtdM359e9
V5h5UEIdD4gd0MtILwUgBstoxm/pawwxwvYWYbWzJV60cH2mXDuwCfZNMT+q1sv0YcgM9yCfg2cG
QoAQCuM8ffBs84RVoSzU66FDCH3f1ZdeufPgL+i4K0zmtpieuw8ZuMZKhGIhP5c/N4eTO642LgFq
7kRWYtw70XrLyEOXR7mSKzJ+b56XWKrnK4iYP5YMjqID0vMDjg1xZ29H5gxVM93D1mqGYr6vuTNJ
7RGCsQ/1XEAJGr9XAG8sIjlogvjYG2MRcYcUK6Q5zD11fXYNAOfTy0YvCD+7WKgj1LR+FcqQKNst
HczXrQrHKxMotVAt/1GeTqJTEV9mRJgzpLtWKhkDqgJiK0TePu41xTWjvcEYldySOww9wFRbR9Gh
7BdsqVPPTF4Pv1x+1KZ0Ujt877LRGejrt0GwGJ+GkVmd+MW2FXTlyH+bUdlA6u7HRUy77eYr806T
V6j0QhgcoTdeaOm5GolFMHZA1d9GicNw4moHpm+z2RZEfAzU41p7HD8qr08IGZB992S/afeZyW3U
MpJxP0QnLBF2egb3b6zALfl7TwnSn0kuB/NyeQHLwkq+x6NLB2mgNFZnGVmdQuKjviWi4+8yY4Cu
N2Op7DSaAdh2q32iDiYLcTBwpBqCFqjWMV8YSP9p/Z1QxU9Kgy00aj6cvEey5SwFH7NIgKen3EHw
L0umPc9GsF7FLinLGqV5seeGEWmJPXvPt0C2bCKI1X4+vEMp78HbwIq5xw9f4ZvUwOwkrFLErGBJ
AIyr2k8sMj+045q6G/l7+6FWcs5399ud0MIyygVbsAoPNx/p+/CjODaojF1SiWu9s7YK44Yk8qGa
lzf2BFswlkwXamOQR3BrUdruuO3awVXPjKZseIx63A+9goz7xioZFzKAGZ/B2m7sdK0isjgszoXR
EkbL9EAK0VBVxi1YLLht1JVg3JTcJP856pKC/RwPFVImGsk1aBfbQpR6xbl6MMxfiO+zHTeykhyY
OZT4fLHdOUydrboG8biSpviALG2qREim+XoufIkMuB9lqC/1I7g+aUWmsY/DbTi85PndMqF5Vr2W
NtISsenIztRpP69T901kArQk5nrb6kA8vuqNc/ULwU/bHSkDR/kVa8E9PXoxOLWEfmci2Ah3KTiI
fSvcF5bZIvkBtraQZT1/ba+Lx+qMtNBnQJWGOM0NLexNaKKUVCXdBQCAqDuFfuefISU93AmUqybW
iXAMx5CFr+6tZVcCPME62K4eMerU4Ix6w4FkODTys6eOAZbz6RIZNXVosDzPByIBI3RUPRlKEjlI
RGWpbTZ7QHVZq8DG2zYjx+cEybIPfgCAn8C3EqJDBzST9WRyu0/I7WypbLG+5uIRajTxr/82BjDx
LOW9JsRiD4HV8JEtjTHn4mWhXKoqDkVfraCUttii3DpTH6YOoReXFsDpmIX2d9wTh8B2fwP4EVww
tX/Ki2DJJYQwTxI++z6B6iQUWHoWZZj16LU65aKSUIMpxRZBnMxF7LIinTyhUel4oT3UAR+wl0nP
iw4frtjaxJZOLADkl4fntgTP71l6NyESQ8rQ7Azc1cRdnNT7Q4VUH3ke8exqPhwR663FIXrSH+X/
iKXV25Po/dRpaJHv9XBIXdZ+UDAGxBSQHuf0xnPdCDW7zI4OONQxF60mtfxUipt2FI6PI5HPLXJe
GzadJ0X5F7rh+7YEQTjObAp5pmrbHxcvD0fuT0Jowbe0yCxotnJ5HE3OVP19FUY4Tmdifpno4aIQ
yMi/ONrIi8aEvzsSbr5dNhwq48k+U0ZZqXYaW4ngowQ5ZZSlex3fuW5+jUsHiExlVeWdFut2ZGJF
Ce4G3rDSvo72d8ns40a4MevZzuAJfc58jRuVm9zNRY9iz7MXvDdnB+NZbgZcrYya+4x6pcGI6Jyd
d9JlKTtsJii0hOzdTAerlrF5E1Uo5xnXZaDavi7QcPjYARLcsLUZzrJcZAGExVcd4XRCfDS5ReL+
Xlj2ylUUSEzfj/rgr4wA6fuQWizJXLUHqvrQhvO6aOZNjKHBYkpetGX0+E2ZkbawXSUacX1W0+/6
tKb9QX6mwGQMaBBGfQeQHxFoxIoHdTb+QJMakWZNq9QjvCUx6zuvzsX+zNjPJkK0mQdUMb4SXxal
+0tjW3aKPl3JkKW0KguR7r9Bfu8qYxa5ghLqAUyiT4TpIXgxkuMON/t/jSWo8IMEueuYmvZw7Lvq
lSb88TWDK7JoKrFljmCl7kHivK3AI/42TU0apuLYcBnSD1ngx01eUuc5sVAGRbCah/LZGVgURyNa
FNOOfxpqRGWY1A2hvAUu0G/Yc04kWvnaWcNggH45lEWHaH3u7STNnP729Tr3jme5GdWZ4cIw8I8J
8HokZd9VNGnIxliptZ8fUf5mIGAlprruN2EB12QxsxpqoF49glw7WR5hpuTLgSDxvcQuPMTFyeL4
xYb/YvhWdI524O/hdkDt4UUvs0HntOfpFyHpUasjsv6l/0Uv4qy2/d4PEp3EC2G169IaE6LG46D+
+5Jm0l+sdagYkCLM7ZCzBDy4WD0awjHlRYbaa0NTc2kwy7tT3/Zmnk26wkc1k5wHe6F2lwPV6JRm
tMyaEbqRIU1pzF8a5aWGGgOiYmEAjutFrDEjJ2MLiaqDTq1fpGNeFOTaajYGFz6+/TCHswkGmbo/
YOa65EZtS4bJgAtCS1BpN06HbE+xyD0G3lFm63KpjqvAiGjSFVmynMGYrWRaxjtjuYUtVVi2Ceqa
TfLKCc2vcHw/KxmMpnUVBIVWmr1jBvt7nWOIsl9So+VSKd8X44pqKKn5QwvqurtvPpPPBXTGTT59
Pyy5cyKkab0l6lecb55zSv67Ngungt3SWlRiZ43XplFOcqExY+qtQ/XuI2Nu3HHt8Np/+tumyUws
R6RTMDalMsLevHfrGO43oqqLiFSoUw2c
`protect end_protected
