��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	Zà9,J�Dn��� ��|��{U�g���zf`��-��)t�F{�Ǐ]@�R�:�r-`�/�$����^��<r"S?Gi&u��a�
�h����.q�u��(Ǫ�Լl�ol�v�;�	����8Y%��OVC�'8\�Ԗ˟]Ͻ꺨��`�F�頩 ?�%
�}yM��j������k��������WӅ�]!D���1�b�79!��k_��l��8���HȐ��$��2m�9�aWꈶ\G!?�`2�.n��ގ~�0(1���"�uȜa�zCz���N�n��)z��CJTtN������X���R��ӁȾ�Qڅ��$*����a��$����s���X�p�{�W�5]�s	����N�?��l�"Z�\\�CmH4�P���K�G��W|��K|N��K�%80k���U*P���w�CH6}&]S!8%Y��!Y����]eI�	U����8$��6�\;�me>���E�3pq}����}�����}s��=���t��9�q��T��(���� ����xD=p~~�m�&�`�%7T�j|�j��`h���byg3��M_��*y���L��%[8� �&&:2I3A�P>�F{b2����C� �&
��W��D�Z��Ժ=�`�6�2N-%��7�iH<=(06�}�6,�-�P�&�z�$<�a=}✢c��E���OI�s�]v����K�*�,SW˱�בLv���i��.N�NHK�(#�C�%�����*J�WlJ�*!S� 5q���	C�������Md��=-�I0#'�v�4�ۦ]�t�,��*&uj�Y�'7��aJ[ޖ����(8|�2��&*�� �@���F���r�O�S��x�K�|k�	F��L�@ZM��t�X\�}X�& �D��i�}C��GDL�"��SP�%���݌�v8��-�3.��=(�N��������$&a0�T�!���]�QG�,���c ���,߰�R��So�[S�J�.�Puf�`���|��N����ΰj��HJ9�f�#���?B���-a���x�)�8�42C��7����3�QLs��{��A±.�i�͡�RR�e��RIN�DG/��7���e�큒�R�A�.�xi�U��'���4�����N���^���|3�r3
W���e�OL��u>?[L#����@���KY�,;�iڊh[��۷؆ua���e>\�G�P��~B��gF5PDj	�G,��n��cK�L��>3�j-w���B���L-?�>��+�)�1��mf�%��@_���%�1��*��;�|χ��-� �רb�p� R��<�Ӏ��0�j1�\� ���ꙙ�IZ��HQP&��&���4<kgn�8�s>O�i��7�k���yT���+kԟޚ�2���4��v<l�h��AT�;	��2I�)��ŗt
<+o��Ȁ�)*bD���5�.��L�#?Z�#`g 5��Àx�?཯<)f��a���6�̖}�����w��j������"H�"1��IfAS�#����]lr�
��G+A����,�}�3\ �
'�UY�����(0�3皾��`X{�Ǻ����I����-��4�	���f�mv�lu�G
TG�U4���B����ٹ���x�j���?�������ÿF���+s�z"-%�^�K�DQ!xM�I��a���;����N����eW�l��b%������1{��`�����fN��%,�И���]�+`�������� �ϐ%�����B[h +2`;I�ٓ���^��H�|e�)П�,�EH���M\R�)�ͥ�}P��7�b�u<v�@���5��]M+V~�h�y���DU�ώ^.�Q�Q�����b��q�I!�V��5dR�1����֜���+K ���2�ۖ��;�މ�kp)�rƙZ�5��v�!��ֶp�hN��h��]U�2Y��Gp��V럖�=��A5�8��-m7����G�NE9�b>)���Ϊq���b�'�尚��
V3�Z^�HZ`�)�#�^��נC� �)Z�>��Tek�#Lm���1ҭ��G-P��T-�͕�F�����a�����o�jl|����N�T۫q�'[�q�,�µ��q��,)�W�BX�N� �ǀɞtu���Џ�9�A����?���5�}+w���>����n���M�%M�8��8aH�+G�i8��m���p��|D-����X�>�ϑ��+a�xJ����i�6�Yw�,1�g׶�i��]8@Z1ַ\\4㏷'�!�8ت�9����c��B�sG݄��X.�j�̉��L�\�g��.4�/���U'jǡ�Х�HÖ��PۣCg�D�sl�&����)N����
���F��ӝ�����Z�2Ӫ�Asr�,�X�ӑ)T	u��"����f��Z}��DZ��{��)�؃�tH���#�$3������7�{����9*{2Pc}4U��/Ȟ�6�DSP��l���u�˩��X��k_u��!	�����M�yXf�����@�S�o$Q�yZ3�΋*{���ә����	�K�l���W��x�2���ݾҴ�r��O�������o-�m����b��I�_@y�/|��oE�>]WY�¶���ZuC��5`KmD�)"`]F�w"�Q�����Xmђ�)�N0J	c�a��+�t�@��X�]J�/��ד/���`G�j�TK+�{Hǌg�Y����.L�C�OÉ���W���,*g2P2(�,��PGԆ4��1;���0gGȍ��+
+Ŝ���Ξ�Af�̪�D0��*꯾e�qܩ�?��,�@���/�9I��+�ZmkS1��j��A7���Lf�j�
q_ҡ~Ah6����$���p���5f���!x����w���i��-���߼�Zǘ��ʚ���y���f�Ζ
���^E n\>��T.j�/4ch�q����Q���B��_$
��H>\��̉}�'j"s���x�Y�ZJg@����/���X#x�Z:�0j��rP�ĥp#�߭�J1��7�;��ޜ#�;7 �&zu/���+#5�gb&8Ҏ���e�p�iJ��$>�8�����q[ݽzӋ�l(��R\��L� 
�Y����ó?��z�.Om����M]��F22����Ps�Ж���&v�S� ���Bm��G�|Вd�p�?���[LtJ��7�����{�=���u/���.Xz�!)��|<�c�8uпG���ӝ��1���$n1K���s���q���Z�%$�o�$�" ���U��&O���m�x⽤��p��n�ÂMȒ&&;� �F.��d�Y�^�M�-�vp�4��<�F+ik����B��c*o��=ト���;�e5���Ձ��Ëͱ��\/�q
+�]'-��I�h_ٲ��R�NԱ�2R��B~��r�{�_%92#�p�Ob�v���z�:�{׸չ�����W`'�y/�tm�����}�rã�Q}��Id]Gy�Ig�F/�1=����?�i�\�A&� ��0�V%}���A����[e��ȋ`�����y�l�T��*LI���
EKM�-���/%�T(�51�(h���|���@�L�y�Z�e����<
��H)�%$�aNؓ����J���`c�r�5��H��ʞ���\�_�ȣclr��R��y�r�
���%��dZ�@�e�UUg1&��+�	B�<Q:�˲Ɨr�N�c:������w�A&��:�U
�Q�]�H,�r?"ݿ�F���X�FJ�%Y��%@��� z+�X8�8Q4{�?���� �7�P�~lүl?E�a\��;�y+�uL�x�ؐNC��D_R�8d�}�yoUM/b< j,�_%W�kN�vW	��-��S��7i�
��	�{�/L���m�����ܶ���QF"۫��Y-�@���g�vX;�mY<#z]VQo����5P���צ�~�U��h��e��Z0�A�����B�ɻ"��nPL��&�l�!>1��}�l��w{�+��B��@\a�$ɒY���~�)Y/;��@U6��㩘�VC)�@ED}������0l�A��ca)�Y�y��&�����a2��U�»�Y��j!h:\�۽�'��x`O�.2t�c�iiC3�/�9�E"�?��Z�n���f'B=%(�:{�^I�B@W��ʳ�:��6�q��M=m��`,�a��̥v�͢&��T}w]�n����P�)�����@9�)1x�
���_[������ � �-0 ��<�^)Ʌ�
WS|�=��&������t��p��K��7�F���FRi�w��T\��}1�<*�GU ���g��e�8#�|OC��Ğ��s�������f��7hu���>��LP(ܒ�l��!�EB��,H�;����6��"�3B�	0PI+4��2'��9W��X4c�Н�y@!Y�mP��������KP�jZE=5�-��B%���Ե��3Ra�YCF&eW�tC���n_b��3�~r�\=���;�|�X �Be�q��������\+��C�ד���u��:�+n� ��#Ϛ���*nPjđ�Y1�\<��?�IA9/��3�q�+���#0� &�F#��Z����$aۯ.T�,���8�)��r�G��Z���m;q���|�]� �7T��M?9�A��[Й�K5`F=޸��g�8�!)��/f�
Z�:9���Hڃ�N)������9_¾��4�ѥ>�g�ϭo�0�W�`�L��	g:��rd��h�扒u��-yq;��nzl�A��&�$O�Ӣ�L��K�^��FQtW(NN��m0�	�-��Ǘ,��n^�J0��σ�� 8^���f���V��N���%��;��b�f����zpY�:U$gS��E�'P���^�I�ds)p�(�K���o��_��rYm����FV�����������aKc�p���2�u�I@�ܷ�MwD�?��/l�tڡ�͵:A��r6�Ut%ߴ����A2f�F��+����T�1�Qf�C�>�y	�!�&�}�-x2�#�����&�.��q!��vD�����R��ǆ�#�w�>S�r�z> �6�(��>#ۥ^��w�HR��Ν��;ʚ��x�"�Z��	����	�qQ�#�zB$ �S�$;�k�I�0�>�k���i�l£;=�&+L�W�~�>��j�Ő5"X"3F&��}��`X%/����6�*� ~�_X�����V#Ʉ1tUU��5q$k���C�� x��dӭ�,���/�d�ˉ.ӬZOV<��I�?���I��!����lL�;�p<ؾ�"m�A����s�`e,X�x��Lo�&��jPuN�k]ӕ?��8c�^��ǃ�{8F�����Ϗ���/})@LD,l�ܧk��l@~�1����;����Ĥa?���<��PF(Ք��3�{��ƿ�T�f7HI�N�fr;��D�G{�9��ޠ!2(�{8k;.D���1=�& u��fx/I?���Fz��*h�[�W�sb����8���@q�p�+�4J��	�>?PE���wF^
z���d��>9&YT)1��;w]�{����)�݆��G'�m"ni�W�(6u��=޷�'�#6,�SFp��۾�?d����	>�i��m6G�kD�wLR��>w6>-Z�bi�n�3`�W~���q{ݏ�?��*���Ʈow[��?���b���ή��rE������~�U�-\¡��8���J��e�6w3~5aݝ��	.PH׭�S_cr���D5�Tʩ�[��)�w�u�5�e��gʬ�P�'�X���(����5�z(�U0�r2���u������{x-#�;
��`FF"=�7s0�gt�W���vL�r����~Q�]�;k���f'>�wK@�xp�4�Z
��{���r�@�ѵѫJ��:n�Y#��"�n:U3��2{t�RC��̓0�ꉤ�G�v���qd^~�Z�Cğw�L���iv�0���+6az�'Q�i��k�4E>jY%��}JH�e�_��6
LRCk\�:l[/s�رjOQX�KD��x7ɢ:ݺFH<����`�_edd���z��h�w��屓
�~4M8t�^Y��C��9�K��U����Ai��в;ٺ߽s(�Q��K�'C�Lʾ�=s��H��%!Eg�E�͎����J� �Z�`Q/O ��%�x����3�D|�=�:L7����l�*���L�%v�to�ذZ�)����"t����a�f�� �b\����m��y����g�Ҽp쩊��'T�D���n!l�!w�
�.�W!���Y]����{";�kR}�55?�,��;�6�=�
z�Gt�+Nİ��^;$yZ�cp��4����z�<n�����nX����纲��o�ڡ���"��xݚk�"�R#�7y�>M�b��5*�8R���P��5F|�Ԟ��-��W�7�^��Kd����5���Ԣ�j!�&j�Jb�~�;�<[��g��'6g�]#e^s��e����)�����@RqJd�?xi�P^�X��ED��Y�L���������#\���f#I�(w��Zl�C�����g	��,[^"O�� t�b�}�R��e��ү�)�m�I���)h���jaյ�b�3 �����'��3�������s���1�����%�)X�X3Ү�V+ǰ5�a�Q��˿;v4�B�aXQ��v4�;���'IrC?M/�֏+Tv�&��@Fs��7;��[�*O+O�5>g�9�>$bP��1�0j��}�Ě�-�kn�!���ѽ�ǰ_��#6[���Ì�FPbб:"`��U0�	�^ݡ�@��.�D�x����EK�����~�g<n����x�kL�$m������Ma���Y��N��"�<�cS�	n/����˲�Td(��IJ���Ir�l��X���a���G/j�9%�����x[����=�����_�`�V�����O)�Yn���8E��5��w������ -��Z�����shWG�@�3Zt$!A�VT��ͅt��|��?0���#�c�0���{�a�<]ks�C
��
��h��
�����%�WOc�O	�g��v<:�(�b��ZYD��:>:�Q��)'�,����>j? ź����jE���S�y͟�qG��3Z�J��p�l&���m
T=�񹫸���2�t�R᪩���K�?C^[��VK�a��Z����E[)���>����]�-MB��|���_�^���B@���g�f�T'եE�ÿ����������A.V(j
S�� �UI�� ����MYy�j��6�����0�� ې5�2�.~O4ֽm#A�u������
{j��`i,(JU3�Ə��{�lS�|�+�&\v���'�)�hu���ϾO_gq`o��3ޮu1h÷�;�y,�Ҡa�]��y�3��X)��׌���}6��
x�{�%��(�è�V�zp�Ϟ!���I�`~C�0��L��L�wxߙꭆ�F���!� $�<%�X�1��D�4���eum�N�1/ )�DrZ�Ƀv��P�}��,v�S;Q|�XK�^�@�H�cY��/�G�7o?U�B�oX���N��G�L#�n,r�Xz���ߏ4����w$q�T/��:1�e+�6[���}q����������?4��t�������k��B����A��<�O�W�,,n��tͦBrCAX��-�]�7 H�tV��`��0�̷��Wl$��9B��|?>L|-�,f�$cl�ٝ�G��@��H23?R���<}�L>�5w�_RkT�ab5����W��A}*7G�ĳ��K]{�As���{j�l&תN��ſ͎�� @U�s-�fz�G]rtL([����c	������"*q�Q�#�*b��b�A9��8;�����
`�z3���W�i	�ۣر3>Pᔿ��H���F�GA8-p40�"�`�����fפ�eC�@�	_d�g�3�R��~D��F��᯺d�(���k�+��T�(*kߣo��O����m�
+jn��|�'@�1W�'�[A��:�c��cu$���च�|E�;�x�Hw�Ǣ+��x]y�\�J���w_­�$�q~���7��iMaG'��=�S"Y)��neH˳!^�UH�u�&��-��+NH�a��-���Dqc��#��^^����wV�LᎾ���ȗѨ!�C4_��n�[�;�ZD��_]�,��G�W��<�Q=`w+�11��[rf��}}�k(%��2�hX1��ÇH'���d�+G!�q�s	_��.g��O+G�<� �����饌F�ɰ�t+��x1l�R�1�0x�!��7�; �IpS���d�3�[+/�'�#b��kj�W���/9{9!wԣq��`�q������ї1��y���m�J\�:/�\���A�*@�<x�司�(����r=��ƌBR��(����ŭi��|�7B3�j^��*EJ�	��l���)�p�d�'���k̛�e*՟u����!�@0��+���y>� �"�c���)�R��q�
�
V$�Z $2���|x�(/bp�ı&����q��Q�U�����������ơ��j��(�t����� ��ޱ\�U�X�����e�t� �˫�e���%�*�� �Y��-Ğ�F-�I奜CT�K�a�#_�I�Vw��)�eBPsx����T���o����$?�倍�t�u/6`�Q6���L<j���
c`J/<O��0�&�_�+'8F�����L�c|�Z9��`��P����p��[���?��x��u��˘'CQ5��
T�8EeoE�����)DýIl�R�RE"�L76��n��n��4oh��]�r��a�W�~�T�f�d~���w�F:�2��eTyC��tC���)�h�����SLղ���=��b���~�B�����3}kN���nn;�Gga���s�!��ٻY@��&����w�����u2�:��U!��|E7	��%&D,�޼��ڝ��烌�L㛑t�vWn��	�V�YS4I�lX��
��<���'����P�Ĥ���.k��/��1��Vx�`�@s���!P���z$e������]
g�@�2/��:j�k��t��-��ˮW��ƈ8��ҕ Q颫b��5�- õ&����w�^)o?n�m��1�V'LEཧ���`+���g��pp�ջ�� ���SkRG�y�/Nrz�lc�������k��Pw�zaa$�K6)�m�f]mv&���f��w�ܐ���n4�6���*)+�Mh9��l!�/؜U8���'�}=>�������g}�\��0��T�l@׋|B���bM���"Z�sbR���u��8���?�1rőQ3�3_�M���4�J�i�;��Y��v�F�H�11mP���uCs�i�x�*c:�"WFg��q/��J�Ḫc�5�H���Ȳ���
��:���+Nb�B9q�%f�HU��woq%��Pm@_0�|E�TN������ys+������~�k)�Hܜ���]��d+ݝU�Gg��U����N0��^|(�Q�Os�����Bm���X@�&�%V�����}���+<����b9��a੩���Lw�w5��`��d���e$'���B�k�=D[��z��kogĞlk7��=4�^��Q"��E$vQ>�U1C�WOMͫ��sy��NMݩ�?�%�e �"c����}�܆Km�
��%o�M9,'s�������8LW�h�nɑ�@{q'J59�j�d���p��k��R�V
�妅ҟ%��\$M���]s�X�G��S0e�		DL� U���x^��`��K���U[u�;^̟�]�\�ܿm����i��w����qL��Y�Gٙ2D����3�{fH�`����%�3p2��#�ˀ��e����:�(?��!��_շ�W��dr�:9�� jEɰC_ײ�$a��@�.�"@�_�rB�����rX
�����j����r;���I�2�J��NR�B���U���5dnv�I�SP�Z�|�g�8?�7_&"�Ti.\���;�05p��0y�fY��ZpQ�z	�^x͜=�ćhQ`\�x��~-��b�8��w���>�a�]?��pd��c��\f� �-d[b
�$�W��̄�Q
L���V�F٘��*����5N�&>�[EѾ)Vϻ��)�n�L�-�La�V���������jT�;�T���V���q��yY�aB�M����&.y WQ��ǅ��%�h9�R3��%����c�ߪ��&4�"\f�T���k�E�}�^�9h�li�Q��5i��}ƪAP;�)d�/X:���,[��:V�oyb�&��`~q�\sψ`��}�M0�� �����q��=KH˃����e[�Ԉ������Ѹ�Lw[�U��A"J�����^�~#�$,-׆���H�\]���x?�b**�5ƸG��a���������\sޢ����IW��!�p��3�i��g����G��{	уJ��>Ĕ���͊7p�,���2�w.|�nN�5������y���o�.�.u��F���C���L~W���@\��s�s�8N�_�xr��� 	m%�g�X8�Q<�let��Zy�\�W����� �����Hֹ�>zl�n��V�����A�,����;�,��e��,��.�~�����A��{�K�m���$c�aG:��Cu�������35���^�|ըω��9�Iiǐ�nڕ��q�b��g�;���.��/}g_�8���RB����rQ��B������e���*k}�G<�<�a��%�dEMI{�#����2S�*�Bq���ԧ��b�+�Pj��'��Z�]�%�x�C\<�a�5*P�O�@6��7��Ce,���NG�Jf�k����	���U y�
a}D�V-J�bRL�#<���pr�x��2q�M����N�T,QL�Q�Z�\���D8�lw�vq��lz4�tRKw�[�-��uEB�>i�4��f����"#Se�T?���\\�T~
�I����z��.c����d�ܽ���4��.�_��ӎU�ň,��������t��$!N�;��4b0�SV�yYUu�^�;��Z��T7�m�}��p{*�g/�ȓ}K�7�!�����̈́)1�o�	��#�IAq37�*>$d��,�:;���<Ƣ@Z5��a��1��uc�A��!h��_�X ֒�/���o�L�y.3nw��{�V�]Oە�;�E�:��y ��0��J%}��yy�@�S��؎�4GWtۡ�v�*� X�q&ӹ�@,J.��1��%��L�)�Gy�Z)����q9��rׂ���r��j�0�=g�ֵ��d�찵 C�u��-�N��Т,�F*���]�n)��?���N9��{08��C�y�4z�����'Py��-,d�l@�׍X��֍|��'���)��J�T�o���7K�o˩7��e��K��h1I>���L(&�ƴ�)�,Mo��&䐕��z�s%4n�#����o��U����p���c�7b
1nVb���޵ǏE�t�X�,�η>L�G��D����>�j�|Gz�jk�EQ/���9d���VzN�@!�+��J�+�3�G��҃�����%�3*n���s�k;�tF��j�ϵcd�����Z�^`l�(�* J���G6 ۊ���ޟ�d9�Fڅ�ȷ�Ĭ�$+r4z�my5���%�K��D�WI�5	���^.EL��	�yu�k�L�Ŕ:��8�9�.�V�'|�Ux͒AهN5�XǝB��C�##'[�<n�S�"_xe���b�m��j���H���|6K]�z�ՙ��6;s�����b�؞��a����oP���2-���� ��=bWoE�%�+���VN�"F�Xщ��M��V�©�l ��K���	���D���/ށ3�������zN�}����
�Y�	|�!	m�a�d躵Ӱ�ҁu�l�D�vɆ��=��oh7oy���V!FR�����q��JOj�w��J�]�k�b�.at�:������&� ڬ�r9�wKx�/dɂ������2Y�T7a�����wVq$��F������T�6#4�/�'᯺nO��.��v�P����\׻$Ҟq���3�:Wn1�2߮���ԎA�[྘ȯn��#(\~�&T,���j��h��P�i8����������3��Co���rՠ\ׅ�ٹ���%��^6	��Sb/$$�������m��ċ+�J��N����0@����b����t�[�HS�oQ(�m��rg�����9�b��.t��IA&U$����KM�!�z��# 1�h�߯��i���15�WV*��铟�Y��"�+�lc5�v󷛁��G���\�B-P智&\�Vd��-ۮF���c�k�%�j�91]`���u�"�3Ï~N��M�+�s�/HHL8���]�/�X�<�GD��l�7H"!��1o$�A�[[��uG� l<�pf���(���WAZ#j� �E�i��S��5�gă��T�|�}���ـ↟�BD��R�e�P%WŴ�Ż$8�n��b�KZ�%��Y�Ł�k�.��l�}�}s�U���D^��6^wGD�`[���8T�`ͨh��DY�E���E�Û�;!���\���	�B8�: �Q���;^�����7C/�[��Yл���7R����#�T@Q�)�Uc�·J��UԞ���e<r��[���t��&��4�M/�� ���\k� ���#FZE���L�������]��:�)D�Q� {y[�F�\������ު�O,*&��j;���z?�DA
��n��}4)alַ4����IG��L�BulE-�Xv�~�ѥ.yk1�7y���(��C�3&���V����
ܦ2NOpV��6])E��)�(5�3�.?�`���t�vZ�79Y��ρ��2ݥɏ��B?���2"�o�ƿ+���`BQ�#:&Q)���6����n�i����^hw��%&�^&���Y����c����IH����#��0"
��؄Tb���A���7GHz�������[��6Ǳ$xgor�7��8�n��E���tAb�/)+3�Ę�,�}e�fj�= r� �"��R�����}���ȵ�pw�0�P�1x����`(�:�C5c� ����TIN($)�����^���%Y\K$3� ���o{j�Y��J�6h�;WWQ��ns>�}_����1�j�V��T�����.t�K��?
^\��R��rl?3!r��C��Y�R>ȩ�bg� :�=[6����q���̛�o����d����)9��[��\�e�g�=��U������, �[49T`�P��
���ʡOO~�;�ͳz����o�y?k7��Q��#�/���3�����>���;�>_a�72�)�k&x��'16�:�8T.G"b��F'�u��0H���[ )�`D�9���.|t��̟�vȘ�s���.L�~��!�߶S�ZtnqP��`��_Aږ�w��p����|��TbE�a����UwnU�I��{$r��aD��~V�ҍB�0l쪯3]5�k���n�Y}3�{.M�*}����k�I�/gq�/T�&�Gt���W�CNA.���)�gȴz�C�p&� �*@�@}��Ɲ�'~p��Z3<�-�
�0HV��R/��4b�
���"�:�AS?����?�NB�qs�� S v���	K�7)�e�h#�r��Ŋu�X$�lC�6)c�p6���k�Yp$�Æ����7�(��Ɵj:<Q�PHq��m�/U?��q�\�����#�A�qf$t%�{�ö=��u�t�g60ͭ�l��^��T$�M
�)��̪�a��T����nxە�7�Χ��9����K��wGTe��E���
S����֝�Ю
v"�3�>��Rd��{�CC���Q���ş�U��T�9n�>�^����y
��01=N�yc�T^]�E��	��Y���	M�[��y.b���^W,e@$�Z]�(Щ���RZ���E*q�{���Xz��LO.W��BCcr��Yv��X��UzR�*"��,#K9�f�$6�WŒ8�
6��r���{�.�&.a�j>�
t)��S��LF'2�B�'�x�$h���m\�Z�"�v@����
?ִibz/��L�Vcݹ�h6ȳ�����V3��A����d����@<��>������]uuTzsZ��Q�炫��Q*"�x���T�tsY@�f$�{g�(���d�,����*
P�K��,E�������1V{3�� ��c&��[IWv��|��[X)%��k��M�ri�:�u;�Ҭ>�˨��s[�[�3��#�5##%��y���bO�^hi��͕���!����Z�:��EX!t#�M���1���Z��b3�sS�x�J���Lm�?b�ߩ�]T
.��tv9k��FO�tD��<�����K����*j�������CU&"��i��������S��#�4_��?-ee=j���8^
��c'M���9��,���<x*/�����$����([��En`��������<"��w�*��h[�l�=�&F	��{����Ř�ZJ_�0���}PS.�Lp�x��W�j��O4��&����%�i��6�@��wT��B$�W�I�l�.m7��>._�D"k:�,O=�Ѳ��2,�I?-���:�	~jx�M��4�7����VY�熾����w��B=9��XT��q�'�A��I��,As�i,���·+�|{�
:(���\��=Zݱ������͗���ct��Y@��>h��2�M,������zL�%�h�:�.��@��2���&��(����R?*���J��7�u+B�^9U���t�*xٓZN(5>y�u��*�:�N��	$S�����I'�����9wgw�����J���|�e�v"@4�	��M�����
�?T'F�G���==L�jXǋ�2Ł�NV��,t��ê#@��)v�Y�	�S�gE۔�&�r���B�Ö��/Q$z�=P�6bEu}C�sk������%vds~���Pb~O�z0-�p��Rt9X��P^����::�b�%�'���eA�b�F�c���+@�'B%�ϑ8l1�}яY������6�>p��^���t���Ks@b�-�����Q]�xx��D7�h�����k?��N(�H��#��6��R~��P~�s�͐F���� �c�h��D�rϵ��D���ȗF^(5���#�K��!ثYM�.��<r�2ӜP!�)���c=^���K�͸j�{ȃT9XV�]U��k��<���o/u�u���܍Y+�sx�p%P����V������y����79�g�Ԉۓk欲�;[h7.?����X��~0�H�r���"O��KC�?J
�� 9������$w��=���#Aŗ֯��Kpx+�����Woo�sw4����B2�ǩX[s�5�p�y�q���z�q���e�M�9�DA�,��+�.҂g�P(~�K�� �Q"j8(��=�1��~s^�ƍy��N;�!=�%E]��xݲ����0�t~�|�7�{h�O��1�Y(
����!Z�	����ġ}߾��:5ŋ����
�:L��G?*�ט<�:<�73>�ʿ@E�zj�]m���;"��l��A������������C�6w��OӐ:/w�#�#"�2�d�z�*]m�pĳWτ���F�O�|�R_�b\����т%VإQ��"�L��;���"tʕ��/d�90%���<Q����m��J1�5-l��VXw���R���ҍX�n��wS'a�ݼZ��������8��[4��4�
�PI��R62��~�6X�R���Ph��vB��^P=�}����k���@`F�L�����_)��]6W���jOT.�8���c�B�F�T<9*%�}5O}��ڎ��J���;��O�%�+�p�p�KV�=�i�Sp��#:��!��c��%�H���/��tn$e�% ��6��  i,� �@v��pSU-����m�NIYMaQ2l��ޭ��43ug��$�ِ3hhuG{���ʉ�!m6�A�&�7}���k�3ï�vx���#���Ku���*O�,,ݵ��h2j�oJ��/K�Y��Y�#�A"ͽȇe0�<'�(%�U�t�M�����HgV m���V�5*a1XC(k��/ �� Zb*�_�U��(_��w�QY���=����!����TQ�^.�D(��Lr�?���*�J2h�����D^Q�q���]D�3>�
:��Y-�Mx�P�jA��Z���7x��>��l�@(H붎zѢ��NGz7�ѐ�s~p�n�|�$�$(�w2dq0�a>�/QZ,���6���zb?�l瓮C +�	b�~1�*~^�%��s�#Y�(U<��'!��rp��z1F�����ZYk˟��}�0�Fb�z7�Y*>Q�4�A� |O���]�Ν����߾�����z\��_�I��juTT_�*:E�N�et�k���y=(������}DD�G����Z��[��k�Ў�Gs#!�Mn�7C��^�w��#!�ǰW$�%������"����W2�Q�\�JЇ2�q������c�=�O�����<Iw�]/̬�x&y���n�4=R���3꪿
�5n�?k�)��߹��GȈ#�-'�4t�1Qo"Ĭ��W����O��a�]�*#��� :��ڱ�ώ�]��; ����Ү$�r�T�#F��)l�$ه�yd�(��t�U�\�
JE���E�����ao����P�ߪ���l�w��x�(�_v�[Ì�&����_s3�1צ���^�ebcjJ�`��^v�M
 t |�=�4$�lV�ߌ}�����p;*@�tx�@��2ʀKcP�����i�R7���?\*�����
 �a#Җz��/x�x4�M %Ø����v�bQ�X��\x�G~T���c�{������2�j� QBv���'�Ơ����P���,�1H�}j�h�O���>^� ��0��r_}`�Y�n?�B=bTt���0�P !^1���\�-'��#g���/P�'�#���i1�.��6�#4ΨWR��ς�(�!O�W�u���ߗܗ�(�Q��w�g�$Ҕ��g[������|��<�l'�C�%�F���O_O5б�)	dA�.���D��c/�kC�*��#S�&3]��1�|��,�v����I$'���ɞ�������Ķ"GV�?�tHj�)��In�!�	��(ds瑘����!��4^ءwh!rL-������iW@!�6Q����\^t%Va�!���^�dI�x2����x݇�����f�����k��|�v�|���[-#T�W��������H��,3���Y�!�3<i|��tʧyS��tH"|s�ˬRz8k�d�q��Ӯ���0��lcC�Ek�}5O�r���C��G����R>]��zBg�$���M5ۄw@�m��I0Hq|����hp�Y/+_஀��yo�H����B���B(� �*��:�����m���$��|j�i�_�-W�%�9���Zi����D
o�Eh ���?y��v���&w���떈R@?}��L���)�y�!4eՖ�ج
���tE��������֜3 N�-Sc�,Aq���Q��:��X�cc��)�#�N�O��IGt}��UU[g�_?0�6F�c~:�$t�XH�U�Ꮧ�#�������
��0�S��be��z8�N��LM�@2N���88�j��>�q�*��?������'���F[��BcLw��kl4�غ�P��k�k�t��h)��흻cϐ��F�l�9�A9m��O��]e�S��6��<څ�����,|�O���}�����!��R���������6��7m�Z��� ��u��0�#I��.jl�$!�������{��Xp�5��.Z�{�����ĩJM��G^밧�n@�"f�l�cm���rN����y`�IE|�P��������~��ᩕ��������'�囼lX�2�F�i��MT\���=��qrd�t�K2���JӗƏ���[;�����K�W̽�/��#�=���S��m����i�ڴCe��k�&6�N�M�nOO#�&p";9ʆv���h�t&(���a-;��{�fDX��S�ZH�kq�j�#�O��I�|�ahq����5�I{>�
��uy�Eς�o���Q��uh��iҸ�3t�˚_+�ߝ H_^���r����K*���W(��H�cg
�?��	;l�"�QG]6�	�U�P=	���BE�vk��
db�5�'��d-*�l�?4u�m뻀=gs��MOx�ɔ4le8������V�u=����g����F�GVP��7b�8<Gő��Q0�"iY���;�eߢ�gy�=� 0����"~i>$�;�X�񈳅����N��Ǟ�q [Ɀ�5�� �������/���Ɉ}2�6c�]cB+�!ƥ�9ĭ���)���v����R2�5 �w���h
�ud���	ڔ�$  �����O;1�D���5�;�9~���k�d3�E���Qm��#ІNF���ډ�dCQ���(������EK��"�i甴��rP�������kb����EȗG4������7r�ᱻ邛&�{]g���.���E>��l5!�D�m�JS���I|���g^UB�+�c�Z�a��Oh`P�T����jGDa�z�J���x�%z����`ɣDC���b8�)s�8F��m��({�JQ��Ԏ�W�]����q|˖1 ��K���h�h� �ȓܼ��f�#�[��E��ڡ2�������e�5jQ\����}��$!*�)���s�-~�\��6m����T�$?M�I-u�ŉBs%m�ًV:���:7��On�ؕ�݆~�� �{+�k�w��h�@�]�zȕIR�<����cD�QB��9�U�M � p���07y��(>9�Jn�P��j!oӢ��X��1\�H��!�ha�=4�lt�X0F�'X1�rd.��L �p.�v��,�#����ۄg"��	���/�d4�p�N��hcbp�kK��.�����iLv "g�։Ѳg���d����J��lEꨜ�,�|�c5dg�e@�	 ��2��7.~gF�"��s��}��]�i�!d�DA]�,K����B�ӒF�S󴡈����=�bN4:P����5�����X*��U��y�	��4��vesV/����+��)�Z?-j �r�����s/�H����P������0��|BB��8���S����������m$�������H;�X���dͥ!؝ӗ#!_�G�XG%�,7C>6�g�wk�Q���hk�p��c,N�4�Q�sb(ӧF΅��m���q۫&�-奨��04�s�3��*٣�&%bB�@��]�1t>���Ĭ�9���`T��-N�G�ږ6�U*9�K�m^�gyݖ�I��C��h����3����Ő�W����W-��O���A���'b�#R�R�M\�
2\��r/�o���tʍ4���!���˵1��ˑ�.�G��Ih��#���a��1��X� �`:a���0z���+��5��˯`��8i�ܯ��[)ǉą�m�� ӯ{"�)O4{�EK�7=��m��@E	�}�?��n2��T�L�%^/$�
�E���A�2���f���2Y�/K1/Z����;���㞊-h�m)��� ��XXb�xn�R9&G��y�L�^�m�=����#Xα\��'��
ې�i(��o;W���3f93m��s8�>�@tAD��W�����6��j0;u��tG�#����l��7�C��HX0x�6�<$�x%� ���+���YuR�'OWַ�y#���Փ�8CA8b :g�@4X62��d�YGZ�Lv��^�g��މ	���	���k�E��gE��{�i������`�l���X�~�+Y��a8��C���'|6 �}���8K��Ar	�s����Z)���(Uyt��B���8y�q���yE?Z�M�Cq/�����'ʖ�',L�_Cr����Z+;d0��u�?�$����v1|Q.?#�H�4�)���>��*������ʞC���^��P�K%:��������f�-lU�9 =�a��@eŶ� �4#I����ZĊ�VvO�y��k-�t%���ڑ�N>�DK0<�w��`���{�M�4نB�m<��-��%QE��Y���s��G�m�U˶�"����
֜�r���-Zh��V�㿹w�p&EP�v�BB{��m6��O�@��$��[�?�d�e����]��^�������D�I�[㱚�~qH��a�>KAk�Z��}�0��4(&�P~b]��Ċ[Z�eh�z��ٕH�T~#)+th�g��3)!�[�:�W,>�8�+~仭�n��Q���ܚ3ń%D�u0y�3�*���]��{f).�f�:����-�ԅ\9o�sχ��/�8ٸ�Aߤ��kXQ�,�s����k�œ�G8�U�I�m���	�.�Ʃ`ԝ��P-�H	������w
� l��cZU[T��v�-N�T���l>�� U�g��֗4�j5w��|�����fX.�����F�gAڍ���sK�θ�Q�Ы����N\/6�Ǆ+ֽ�g~�8�U�����?���-K[���L�F����5[�K{[�K�U�,hut5U�G�,Z.�JM������*����M�T�0�\�q�E �������d�T�%~�Mj	P@Y����އ�C��Ab�3 ��F�AMdA�)s�(_}(Wŭ���4I����*,{� dZA�'����M������t�5��qj.բ{�i�	C�����1oV�y^f7���Ӝ5�f���3i����)v�*�la^43��)�*��&�����=�Ww�&�C2ru;��F����kj �� QB��PR��/����0'3����f�_��we�d
�������s��S����G|�"Ft���)��������e$#B�h̞al�wK��G��斃׋Mb�ʉ��䦋���?i>��8�݄ܩNh��L�D�j��,B�ܤcE�+&�%�O;!fL�S2���E����;䠳�x�-V��<�[��� � �Ջ.�&C��SÏ���Jw GU��
&O�c�E����>��K�������)A+ܾ�n��]��r@b$|������>�A�H�L�*�g������ѯ9>$X����%4�qJ{��ve�=�p�9�A�e��Ӈ��HJ������zC�_]U���$"�<���za�Ҹ ��-�^�Z�b�!�D(-�'�����"C"�#a+�D���<��G!�y���f�F)�D�;:�Z���T������p���3���s���6:YYp)�P:n~��&Qr���ԁw�V���z��Pk�����uw^+RW�ͭ��}S�u��JAC�~����5�g\�O�5CF{��\0�+�=�����?�������)���`��0ё�=8ِ�BLH�]����2P ��00t�����r�7�.yg�Z��ɱ�{o̡#�粩 D���D�Z�A_��5U�a���|�9z�s��V4��-}O��1�5�3!�F�-�G�1؟ܧ���:�"%��i�����_ۘ�F\7�*>��q�C�K�q.R�K/],�9�3�Q���p���4�U*�LL/V�`e�ё�/w��/`����(�;	�%�U��T2��AI��b���?mo�u��.��'�ZG`i ����-P�P~U��3���]�Gt8.�@�峌愣j�nMB͍�;�f$�o�ox<��A�à�9�iX���$��?�]��}��~Qd�ؓ���� �*�:nR���ޏޡ[\8�&C�r�edR�rG-����XD��`{�B�u�Djh�o@U��;�:l�$A�|�w!�����}z��Mg{ЀR�d��)�vf�5}+��~�ᐫ}:�O�� "
*�{�4�Gx�Lc�I&�j�'�b���u������ݏ���:Vbݏ���	x4��E�(��"�@"�#�;|qdֲ�G�\�'{3n�M�AbF`�G��1����9Y�� ����W�9��w���}�J�0-lA<A��"j!�a���/c�����#l����CM�yO�fc���E�Ի��q'"7y>��aͮ�S	���Rl-�M������xr;��rݬ7r6���T?7 }�FG��D�Y�p��N"��J橬����Oa;�4�wLQ���NT�	EP9�F�Fxz�Ë7���Y~�	�tv5<h��x�]yz�$�l6G7�1�6�Ǆ"4
�p17�OΝ��=U0�}E�R��v�MrT�m��=���{�VL��S�vd��<�g�s��u����_-�*k�Q� ��Uq�mvV�5U�l7%2ݴ>--���i˓#3'��	ҷ�s%�[����EV�%֝��(m���N��*�ƃ���=v1#G$i�Gt^}��Y�"U��L(�?L1����q�G_���d�'�����5�9;�ˌńD���д�D$���oQN�~$�8qD����v䤔 �
�-��n���w�$9z5���!́`~˻x��i4��I��:\�(�[�?��R���D���^]��.�Ԣ��
J�~l�K":_�d;1�� �/�N~�¸.C���L%���!�;�k�U��N`2Չ�+�Tb�ڂ:�c��m)��6�4�<�hxi�/�T�$��8هl�O�c	NpQ݁~.���T�KL����, ��Z�Je<�e�����3�a+�K��i����
�oflc�V|0s�R��@{<��-�B#6��~C�π<N�&��@ջd��/��8�\|��iU`]Ȥqط���� y���֎�(vD|�f���E�^�B�l{����^nt,bT^���#E��Ǉ���rr-xg���u�+�����Ȑ�y��D�'g�ݦ�����"��{�Ŕw�^xû� �� �
ߖUeN7�Kiժ�\�O�Ϙ���,�a���0�a���LO6<����8�����������K��g����n]����(�Lϡ�h2��^��_�15)��4:ϝ|�p���.W�C������CS�Hq�A3"���ip,�x���^/�4 ���K���M_�����8[�D���B��Oh�=�|UL�Tu#��px����\����x/L��e�n~�� ��@���"Ϟ��V���H�,F��	���ix�:�؅>joɗ>8@���c9-��&�c�̈́��(v��WB��v�Ha�?�e��a9�J}����75HUM�� �Nb	CK���u�e=�^_#-R2%Z�)������nl! �/ }y��(��h1�*R�j�#�}�D�����M�E��Þy�(���X>_�	�����T'���J���fȴ�yxs�_����wZ)��+;#�{��o 
�FY&��p�M�P�f]��*����a����� ����R$�J���3�M��+`U����	���o���.�����%�N�v]�7��,R���3��a(s���g�ݻ$�����]Gu?v-A��0�.�5,mzs<f|O٬�Y���zƓ!�e�#(�F��p��X�ԗ�ae��4ot�;RnZ#��zX��*��1�Q�ac��L7�cw8�s��?< �l��l����J���/���O9c̷	cR��fY��V	p<)�0O&E���B�bX�q?�a��j�1��/*��O()ݳ��xFf��Bg��$�nC5�Y�QQ��lV?�����^�O
P��^���[�#��r��	����Q�1P*�����jJ{��XZ֧Ǘ�.�UVS��Hr����O��B�(�9��b)��z�䋜U}��`�S���+��b�&ʇ�M���_��NKD�9��h�ώz�ɚ@N!�D��k�Y!�$۷,>NC�>�
�hѻ�+���CÝ.�=��N�o|�gz?�mG٫�y�G�1�qT���?�Īĕ�M���u�����-��Z!=�i����8�G���/������]\^�^�
�e����S�����h�B��Gw��ƌą2�9���%}[�+�-�y��ڹR�k���8��cyi�OT���u̿G��+Y#���yF�ܼ�� ����c�lD:�� ��V��y����h��TZ��H3��
��g��&��d�KCb����)�+ۿ��]��
^�-G:�-��5�[&�Q6�8��-�y��WЋ����0�Ei#��+��jK'R��H��o��x ���"N��2�f �w�9pr��_�eg�y�e:4*LG�✼����E��������iv�w�8r�r��,���+.���h,�̰�P'M��h����[�[���K��|�U܎�7�6F�]�]�Z]�=�\jݟ,���&����Gҕ  ��� h-Lt@k��+�m��̙�_0P����	c1��%���vf��/���߰ô%u�U4�S�_�I��?������Zn�x�+}-ޯ��^��ߙ�U{��{S�x^ߜ�N�.n���+�@|'�'�i������*:������YAa�<Q�^ƹR�����󨖜L$��w����L�&- �q'�`�o�W6��4W�g'����w�h��1�Ɏ~\#��CU��G�n�獋g@�6�N	M�_^䬦�ծ}��:�Dnp[~����F2ʣ�H���:�܌�埧�k��$�D��[P��EL���5�NU��C*_�>���Ph��Av���t�3���r�b�(M�?����8��� �W�!�4��S�q��}ٳ��V�$9�G> �M�[�4?�+9:��X*��H�'4�p��g�����a�K�Mtm���EG�]0�1aT��/�ьY¾3����s���˫�jgӛ֯��[m&���r=1� H����B�#���y���G8l&�8������	�+�|a�9xJ�����<�y�Gt6o*\��:t^8e%�n2?�����:�#f���N��^Y.\v;z�ѹtޏ�hQ)�oL��m3��9y^&�
��	���v]T���#oʣ]&��$��.��������wz�e7�k�ԲQ����� ���a30�$�Q6v�2d�m���"a��`�џ����7y�����Ϧ׋ ot�
U������(P�w�5���ji�c�Bc~dE�=���*�)��ow?a�N�$Z�G���ȩ��N}�](����%vvL�Hn�m}y��͆��t���|^d�ʐy�<tYP�]�]n��GX�,����r�8�=���	�R��;�n�)��2�,�5oF�֑5��(�x���a�֏�y��#,��Y7�CO�C2�v�BMq8o��G���ڀzk�B�_k�(��d$Yg��j�.(�0�
!8�V�/��(����[����P����zjK��<Y�lM�w$�����7-�O��+=�������X�/*�l�WT��>�"��ZŤ��d���Ȩ| ��c�邯��A��2��I�nI͈PJ��da��3^8H���][#��D�KT����o��7'�䪬����u�v�T�V��Rj}7�F��[:h�.~�+]E�&\���:,��͖�r7�� ����*�ȧ�s�����!n6efW��gd7��S���i��C��`,�"�f��2�Hщ�ܟ ��c܏��:ׂ4�qj�/��v�f��1��;��~��rsԱ8�Ŋc�b�O��Dl+5HmaR�{��!i<�5
��A��i�Ɇ�V[�U��-z�E�~R�xJ&�����if�Ş�_�<�H�%PpE�3��ic}.�L��m��`@�M^~bI��T��k9e�3�Ql���I�s�#5��J�u�ݷ�`��Sü�X�]�@Y�[�2K��(��h��+���U�^_h�/���J���6V�`�q��R�|�#�A��x ̥
�%�5`��iL�u�nݜ-z3�oh���{�r�=i��p�{�v�{�wD	��X�a9a{��F��������2���W_4ʒ�s�媵yB�A���k}��P=@Do��?I�q�wF���kjÒN���RmX:.p��.J��i]�����@(��'��� Ң�Y��y_-��"��f/or���t!�������$ru�8W���A�ZSK��K;����)�?P�-u�-�/3��yX:�`6��W݊�J�a���g<?���� ��&�L�p񄂤	�z;uU�3����Mݷ�0'�]/ʪd������V���;�@ {ｮ��J!D�QQ@�R�u��.�Aq�؁��d�5���|(��M�D�,��}gV٣$��t�OU#�����v�v���jA�����U�7ォ.	*M@*~����;���$4������0� �
#�h�����(B�~�"3�+i�A�|���7aW4+�#�p�Cǥ�rl6OS�n������h��jԊ���"�S�C�㶕e�� T[p�w���hx:��ɒ!����K@.�iq���n��j,��T#}�������$���¡��{�,���o&KF����$���2���࿱��D#�5���ƙ|I�hɶ)(p\�.��K��G������C@#lJ���R�T#�����4�W�C)5I��V�|6���6�f,��A�R*2'�WlBd�k�^�~1�z�Y���טn��61LǼ�w�#R�:�j�����q���`��wX����W��О��n�UT�@R10e��]�m@�Po��xo0�1b�VV���3��%J<���F���,d�F�|<f����_�Qq�/�	��|��.�im}:&J��qAjĒL�_V:�h;@��q�u�&W�.��&���	;�n������s�LA�2�A̍w�57%BZq���M�N4����CP1���B�8)�v�}���+�b73�W��GWn�~��+����Dޱ`���Yׇ��*䍋��R��c&p���j���6;o^�%Q�댜̉[{�?�a��M5Ơ�:�]�*H"���"��1��.n�]�J��.��~�Q9��+x���0XzX�C��6�pf�#6��C�ar_��gh�  J^|���M��tv>�����pv%	��Y�6��4:aJ!Q)>��f�\%��[��&��N�"*�X������]��<t�y�=Q������p�b�C��$����;�"����dJ�A82+�%�u@F��m��x����P�B>Ы"ue�MÈ����~�������k�\�$F��К`!	]��J�#��d�>ˊ�5T�D�O�v�n��9��X}c;W�[a�QL黓�Ğ��c���u�uk�TF0�*=��G�,�ӡ��Hp�i�i~�-��>{�=w�=�}�M��1e�ˌ�;l����)�;@�C��H{C�J��dmA��N��3�l�~�v�~��~���SҐ�z��)��Yu{#1�a������� (h�4��
ݲ3���,�e_��E>x\�8�I߾��|6�خ��P��G\)�����Il��$��'�z�4o��$9��m`�wy�8v	ӡ��Gj^�jɻ���={F��c��*�).mO��?��2<gk�ѳyx!`�l���Ӈ�H�t���FM���M�����mmE���z.�̏$ԇwY@ :`�4Ȫ�[��B��k�p��3Ld��`HUs1ly��m�ůЗ�T�έa"�/���B�5Pi�I�~��D��"�ъj�G;�} ���B��E��-\�{���$����� �.�� �#r�1셚�W��6��C��ѣܙI⣾��suK���:�E�_�J�(���eQ�$�~��*�Q�hU�'r`��N�h�b�dZ��kV�	@��v�1���o�+1���B�q������p;bp�����-�&.:�:\�5.
61�y��\5Rl�T�"��aь�5�:��Bhu�=�����N�A������_L파�B��N'��;�Fj�H�v͉�[|s�\�����7:@̿)r��3bK����<�S1����~1�w��O��[�sL�������R�cJ�S᧱P+e8�t3i3H��t��ʸE'ˉ'�yY0,��������\Od�5th����Ջqτ�h��"��hn
��e^��7Ĺђ"m�J�&߼e�����FtQWI�]�n����.J�;n���8.��e�m0�˔�ݐ.7j��,ދ� :�?���RO�	�t��V�%�Ն�Gm����U;G�p�S��:�T$�0�:�v��� 2u��ʷ������d\82�?R�%{T��N,�6��`�Se �x���CrE�k]�t�O��-n%{ip
�((Yʁօ��A�/6X݈s����	N6�d��#p�#p�/�4L���3�~��/ߚAB�A&��
!�*z9H��q�H�#��W�O�m��i�͐���6�nn�x}�p�/����C����N�Dؠ�~7]�_R�:%I�� P�w����)���e�դ}�C=��W�ȍ�t��NΧ�7U��#�y�q|�2^�aU��mW5��B�7�7$�>�g;�O���ې��6�C�B�^>𭺓z�����L��`O["�dϺu�r��,c�F:]�J��F�/������������y@�*���N��v�|���`�3�G��X4��BsVZc�2�kE�ۚ�Ey��]5uK�yhGm/o��Y"�s�t�5�q�&���m.\�2��Ǚ�"Dk'��5=��>��D��^�S�Qf@3^�IZ� ������.2�YX�'��E� ������oBM�&K����Z�����n4����TX��gS�3l�������n�gCi%��Q(�����nZUS���8y�#�>m:R}i\�GK��<	N���~n�K�N�:������Rmi���a!k�btG�~
�3��#��+M�r��#ѧ��V_b��X���ZAQ#@h�+�H���A��O`N׷�yᐌ��4�s-�Z�Sl��HK>y��Gt�6�s�R��J`4���9����6�ʭιm��X��a�.��ĽW�l[�|1>ֈ����$�)*w�5K\��W\<Vu}�R�}
�w���i�,�2w1����x���d�I�ϊa�d��}�7qa�(:r��y���i��?����le�c����a]Dv%�lO��%��Wc����T�-�!���	�i�ӣˌN��e�A�$]�S=:~�%�D]�Vt��5L�������!�z����/L[G9B2f�ۉa.<+ʫ��X�l،��X�LcXz��d��`F���x4��N|{�Y&���;+��A����y��Ȫ����^���u���lV���"�2�P@WѠ-��
�����S$j�+̂E���e���W�~b���ݰQ���� ���=L°n�P�jE�y�s�����ʈ����Ԣ�����!�g^���ua���']�5�H�:-*n��`�v�N��[ ?Ub��Ŭ�Yc������-:�DS���Bs�p���C��cP*ZG#�c/ ���l����M��fQ��_�Pn�9X(y8�(a��'��<G�f>�K�F�A&ҕGk���R[���FU�a
L�^Icu�lݼ�1��cA�^ưx�'7,�$C�!S$3f T:���D�j)"��xC@� h��՗7G��x��A��K٤�Ւ5�[��B*�f>J�P2]��t���I3�h	�^����gøǸV��HZ�6�ɳ�]�KՆ�'&��vs�
Y���f\)dpO�E�0Aƨ�Qn�(Vݙ�B�o������y��Y����ǲɄ}kA��r׿��^�9��x*�P���"�_f T�3������+Q�A�ԃ�S�o��~��5���h� D���.�3�EQʆ�(�6�*�7�C��D�>�F���p`���vϲ��_f�@5����{L��:������۲�\m�u}���؞3�W7��s���0P�"N�q��:�+B�)!�뛮�qp@��>F����̝=(��$�x�	=ɍ2�"�	d�,����$f���]��a���,xm,T��y�#�zϘ��˱2L�����1}&I��Ѵ���Ҥp� �e�.��)h	�cN"�t0y׺���@�{N)�"� Yo�=	�4Mh%v�R2��㒡�T.�%��������g����5_�%#+<�>+�nc(�w��1�jw3L�Rz
�	| �K�����cK�ژˑm^V�����q��u�Gdb5j�,Bk�m���]�M�ho+�bé�
F[J���m��ߍ:�������!�����1��V6ks���!yڡ��|S��݉��7�'#]H^�Q?"�[Pi�nξ"���B�AX�ª�m��󁰉�[��3����s�K���9�y*���̺jg�:.qZe[�38��pbc\�0��=�](�4�a��7g^�y��ō�����]~�n(��6!���,��T�I<jF���1o�����������WJ5B\ ��y�~.Y(v�˃��}W�ň6�M���9�.҄�bC�N�{T��+��I�.56?%�`Ut�������~��G�����u|X,6����C�]����D�J��枪���
׈�MP4qa"��=(��0��?Dr�dl�FjZc/��e�d����Gd���m��Q�k�5�!�� ���sV��u(`!�贲Xi(�&���2f4��c�[��,q��-�.w�P�
�[I�}���l���|�zv^� I�]����2:�C��#��� HC&T��\ ،�-[�pMW\o��U]��v����F6cu���U�Ӎ<DM3?%o�����eM�Db��W�s-:,mNY,i������T�VW�����,�1�q�7�'��k)��Aa9�(�jn]h���*B-�&-�9�}��R�+����!d�K_���3%<����`+8���٠ŗ��l8�i(o7f<oW��|Ɣ�S�ȸ���I��J���19��U5a��Y���	5}�3��
��\�s��'�՗m��9e�o#�+&��i{-<�����(���U��2��."ӪI+�B �@� ��H<+�5J��ރj�}k�t��-�%�
:����̣{q�eB�*�)�Dc�ѵ�gLH����j��n�&&N-Im���1���)1�uHVz����L`�hؤ�����E��Ή���]J�Z���7/������|����c�u�%qSckl�8C��]��S�'��ʚu������ ��J\�vI�R�e��d7��a`w�tiB�]�~F$׵�#�]0|L��1�'~���TEM�IwD}v'Ɩ�J�6�>~�c|��*����>��?��6�*�'�bh
�η�r���Q�!����C���&��T��7k�����F��ř��:gb�yp��[��e��B��Kf��c��W�o������{�lQ�k�
�8�d�o�Q$� ���i��']5�w���R*4/�0�9�+͇6���[MG⭐x|!O3ҵ|�Wj@� ��V����cwg��A�d���Q�CXI���ssw).
�z�g�B׭.��f# �>v��qGES�I��[��U[jA�;�E�;��a�
����߬���ٜ�O�?�O�rm\X��^�>X1��oI��<���6$Lz	���J�z�g;�t8\ɳD�ˬ��hy`O��幥���8�;��[�k����_��#/�J(�C���ڗ�!�\��
b#+[�h-;�C��g[���91ױ��\`��2��&�qW�L��8f���F��/�!����ՙl(1�mX�����=��M����Tʒ8��cet�� ƺð_�+^?$_�J�� �NJ����X��"ԩ��/ҖȮ�>~�(�V	�6H�@ϥ}O��߸�0{T�$L�l����]~v���lU�5�m�
td0ю�ZXgl�#E4f+ �����]AJ��b[]2���h��j��Ӹ�.�\_;� 򣵉5fu>�!��im�a7,SF��B����^Co����d�&���;�����T��I*_7�c(�r�\���R�Rt�������q݋/t
�����M�F�wa%���k�=������7�
�𲦓�3e�q��6i}�i]4���!������U���5kM %D{Z �"E����ߴ��kG�m���@��*k�V]m�"��=�NHy�����"��a���x)S�7W,��a�����o����=����պ�*���svcW+�Cg���O�\f͗��s�����\$�4��
9䒰K���=��2�%�������9��=������t\�S���*�y�ڊ��`���yY�J�rc$jp�����jM�k���>�AE?���	�/M
��۬Q��vжEY�˿hVJ�Ȧ��x ���v��9i9�#�]X��"v\�-��%g<y�E9}֮���X+esYs�O��y�֞�ʕ�\��*0j�{؏�U�>a.���$=
E7�cJ��z眊��'%U
[Oͭ��s�	�-�;��Z�F�Lm'w#�Yߧ9����F�9�ŝ���"��T�r˞��Z�*��_e�7��\  ��d,�2&V�#�bWzC�i���xvq���p�͝[v�G�q�̰�r�.��gfm؄��A=�<����y�3���95��r����<��S��b�R-���?2���r�_�H9:�F�4��r��H��@��i�ߖj���`V���TYQn��� 8�f
��d��cW�d�b-2��L鸓&�a�`х�#I-m�4��Lo'nV���w%:�H����2�,;�!EY{��S���3���m�eA��y��6�Y;����(BKO*�������|��͈���=������;+4�����{u�w�n	�&hg�^�ߒmB=�~����@(�š��Pn���OG�gA@��t ��&�y�<���}�{���`���'�hA��=�Yc�1~�d�^�d=ڥ����U�˱�X?�A����B�O�'&�*C��4���:� �?7��t`�v-�	z�:.A���R�8Ix�T�4�<�$]������Έm�s�P*_�b�|��CԎdÊ�"�s%�A��(3r/�2���f"~Ԟ�B��lȵ� p�ҵG��-j������ʇ3���YMQ�u�l�%e����Ci]�=�����ҍ���)�I��j�HiE��D<TF�	�J��f�A�4 Ρ��HYO^�Ӏ�=E_ăfB�S��9�����U���!y�J3c��Oe�V+��<#g�FB�k��0�i�Gp�ztΝ�V&pk&oU_~>:�Q�� ��ف*X����%a��ɺ��I��&�3" ����V�#<�s���W��3$;}�G�B�q�����Mƈ��t�e�-x7�^��[���і{�����j>r����O�}�;[
�Ԓ_-���r�^L� �,\�x� ų�?JP�R$�N���+������\Rȼ`t��R�U�d�ŻCӸ�x.����:���xɞ.��R�{N�ۅUf��5�,���4����I��v��O,>�7���E/1�uzP'r��q�)���&��k���c�����	��˩<S���GW��`�޵�C��������+�6��#h?5��4��N0�t�,�`;���ډ�!PX�9�b���=�� �9W��ԖhX$��J���'ʳŇ=.Mqt�����L�S�θ���RyY�J-f\WF������S�]HnڭS�W��̜��Σ/�	dTZB�ܸ�*ŔPc9�t�ڄԳ���-FN7��J�.�;��[����P�
��'�7�J=�i�"p>�
�,1j����h���l!���Y)뉛5p���(���h����^�%�?�V������/�9����
��	@gN��������REP�W�8��^�����|jl?Ko�^g;|4/��Q�,LM�E$V�6e��	���jq�����Px��[ �1�Ym�7�]<���H�߃3Uy��7f�A��}�J#i%lފΨcx�x��0�h��g�P	�6�2=Hs���.u����m����>6^�k���I]�"|�lL��M/�,�8P�����;K�T�*�D�hn{��H� k�S��1�~BJ�=;#o���Pj�*��y�v���v���	v�%Y�Y 9�<�q4�tsi|��R���g�.��K؟[_(a [���.��3ЃX�y#�԰������Oi��bh�nE[u�o]��$�����rҞ{���\F�[m���xf�"����>HkE��~��:f�A��.��u��<�Ř���5��(�pI����1��f�c_�g������:ҳ)������=N����yX��.0M%M�>����9�}v�:3G�R�ے&����{�,=�Q��L�[�D�|��$ñ�d�̇�e5�O��͸��_d��?L1�Ls�jc�}*�	�������+��L����}G����mc���"���_�¥V���K�Fӷ�J��UPO�	�<G��N�.�a^�Y���Q�v�(�-NKc�-�k��;�]�?��2�����B��kq�����ѿ�C�o�Jܷ H�A[Opu�(��E������7N���i3�JҌ�K4���TO�U���V a�ɖ 1I�B�e$�7�]��h�L�o���v2��Yf�C35��,w�R���8O�!"g�� 6>>`t��仚��[=
c�ئ�W��R�@�:�H�I���X���{ :�n����\�"Tu�-��yo�-����r>������~ml;��6����MkX�k}ӛ�lh��]��?R�5�r��Mp�8].�o��P�c��ܡ�"l���q�x�ڡ_i��%n6</|�md9�u&P��z�C���]�/��1B/�ʧ B�b�߱�0!�����
/1@�v���:����*�me����jqX�b��S�ǜj�e���J���/+������^چ��ixz�dK�4�>�5���h������sl�N�H��!6p	�K
e� �����ZVh�	s�A�\Ϥ���G
?����A���{����kL�B�F7i�SB}�#�W�u|�_�f�ԅ��h�%�Z��:D�_��Ɵ|+�,�l��Rl�4�xtl�}͐��i��/fߧ��27�Q��7$�	-F�L`��&Г�:� ���
��Dņ}�(r!D;�|�8�J�3ks
`<)x�o�1�"~��G�Ԧ@�I�TH��ʹ�H89�F���7q�C~��s��"���f�e�
\�,<>��H���i }�8v\�pܭ墅�q��Y�Y<���%:!RW�s��;��U�}��`�E�Q�n/�	�'pm"���_e��`�^�q#Qz�)�;���r�i�4�]����ȯu�P1+���d�l�K8�0�˩�*�;��/����^j�U�E��}�+~"���������җ,4���L$�'�>��H/�$E��W�oӧ5Q(��3k��ˏ36���E���c�4��,�9� ʞ\�p��Y�!p*�Л'���|�'oD�����˨��o˅�x-�⣷ܨ9'6�;�~�3��� �Qi��0&�W7+y�z�"[A7�?�wJ|�ݦhlZ���(w#t��{:��s�Q7pY��J�l����r
��_ܽ+lJ�{��h��_p`o�A���Z��%�|�_h�Q��E-�MV�E�Ɨ�{���o,\nd�o���|ݯn��U�a}G�J�ڎJ��W^0}H�k���(���i_�+;���9k�WG��:G��?d��C��nb�v��߲�2�<�M�;G&ȃ2�91���hu�qيZo�;��冩\�Э~t�����O>�f���~��Uk�!dV�A޾��cѮ��W�$|	��5���y�sD��z渨�@�|M�H�}��@-���	!ԗb@Z�Z�Ţ�'�r��4/��Ý�\�y�b:�<B���z�ʨ-���麝qM��!����j&�-��J�����覇L�aÅ���j�/7n|��Rk�����޷w��"��+M-��L�E�TT*�!�>�� ��Y$���<K��4N�_O�^�^�Q61Km�����㻮������g��7�ѣ#L�V{0Ƶ��]��C2"2���:�p�?pګ����Q#n�~�:"��"hZZ|'L2O�����j�
�m�H�˰�b�W(�As�7��w%�2 �K�����O�T:	�����qL�Q��
��m�ݹ��w�`0b~�cvc���'�K��g�I��,?�㢡����r��7�LI����$�"N��y_<�d'c�"r$@��$���s����T����n��;hK�Nܝ;A�R�$3�*����<wi9ɦ����o��Z|k��}�Rh(��w0�b��]U��ZR|vc�ve�b�����T{���DB�,�H�	�����N�XUX
C��7W�zNH���<}Q�h�zXf#�J�]���bcgӤ������9�W��M<��W�����;���E�A���Vc5�1�9�s#0j��P0�LY�Q�7s-5$ǰZ%�C�8��Exl,��Jo���[+l)ඛ԰��,^g�u���[�F8&�e�ؤ`�����~:���W���|��	c��������K���;��u��O�@��[��x=D���4�m6��J�Qte��(��0k�>��6����!��H.S�=�9x�6�����Z�s�0��
��>�y���ym�~�d���auC���m(�U���C�<���,��A�E�б�3f����
PFl�����*�z��US� N�Ο�%��7�6$o�0����]s�CA�l��c,S;��$���@VW}vT]`�!kN����-C�k{�(������m��L���}��r�ܙ	���>}Po�J�E�2G�t��@��*�����@�i"�6T����f��R�o��w��s(�?(m=ŝt��ڞ�o�F�=�����P8<��E��Џ�"�{ �.��p` ЋŪ%�q�?����n;����h�X�+�oo���U�C��߲D��{�i@���dh�̝Y�zL�i^�5Zm�h����y�G�P�M�*v`��Y�2QWYP��yb,2�K�k���ڼQ�p����7w�¤��7ɶ񷭢K�X�2Ǿ#Q5�ض��>�ؚ���2�
"��8�呇=;�"-6A�鉩��gZ�Cd��9��t]�Iߖ��E��ݿ6������uW�ZP�n%0��I=�rE;T��\��z�Єu�	/�X�B���'��&�q�Y6q��Ԋ���" "��*7k)Wm�N�T����O�r��g�H5c�<���n����sQ����`�.x�����y�0U����SIօ7OϠE����/�[�Y�`/�=&پ���!����7�qW�m�4��?��*�j��XԄ�����e�qp��]3@�{ڇ$\J�2\|D@f���GE�c�w�}�V��mQ7�����x`Q�/�f2��I��*�v���\��~k����^�(��G+�n�`�����;����Zm���C����kŨ�������`(�r��t�<¤y�/UX���n���JM��}�&��PY��T���hn����O���^ނ� �Fò㓑<��88��Ʉ�R7 ��+wg�{�J��,��_��Xz�K���Jʃ���Q5��KG�]���[�
`�6���O������}�-�V�3�BO�MtI�r@�IlY:�dOB��b��)
N�(!��/F[?����a�,`���v���a�MX��* I��Vٯ�AQÏ� �SF�&-iܵ	)���Δ�m���ٹ����X,}�љS�藋��lZ�������H�Xw�<v��4bl�֡�<�ޤ�sWN�������b/h��C�-�B"�^3��a��{oy^(���O��F����F�`h�����G�ǧ]�,_\�#Z���G�j¤m�b�dxy� �����D���hF�A���ݨQ�b�o�[�4�pJ Tdm��uY�ڹCz��1$��,�?����P�W7M�]��*�`z�.!�N�1�-=����k�հ��np���>�?��M�/oЩ��i�U��AV��_�BG� ���w�7-��lnF�Ƞ���e�ױAb��X��{��b�l!��m��{94㺝Gxb�>�[A�`�l��9#�5�x���6$�E���#�2�8'n�/�_H6EF�3S��ل�hZݯ��3P���Z>�t�\i�aTn�{��u��`��ȩ��>��.�\9Y,OO���W����"]���tXe����s�<����l^1�u��s>�&��������(�'���5��f�+�ރ�F)�z�F!�D�$S���w��"�̎�wV��Di��C�������|
�X�tQ]�O���5����O�lm^���&�>b	Nw�0��׷�X�!-+ �~�$��1�jr���EaV�ekEM����9yS���@pyPO�r��o���u>fE���=}������u�^�%t��6Z�.���g#��8:��6���4K�X��Ҷ]�st�&��8�۬?B�&�,��R��D.�ˣ@�3�@I��\�@��3������4��(�
�X���?����6ƒX�8�j��LUP�.;���_ ́�>ya�h�Z�-��u�������
��`g�+����X���󌠕�	8�%}7��?=����!K����Y0/���gt{�{�/w�y��L�7��X䁹;8�x���j���`O���a�' 	~�%�n|A�pg�JV�w(��uܬ�Xg��b-]���ⲿ����7W�&�k�R$�ǈ,�;��Y�`0wga�KQ���\�̧���9X����OM`���@��S��VL=�WC?��T3r@y���h�s����,d0<�F��;_>�^�����-�t�!�ntI�E��?bl��=Yۗ��pVhE�d>J�����MZ�b&�U37ۂk�o��J��������P���;��%4�h�F%���4}��d�7]�̷uNqz�l5ߨ�����$�-G�(�!�����8�VMn��>���ȗ�7xVФ�1�a���6_��N�=aW�O���lȗ�GGur�8���:w�o��x�F�?��MA��s}G	J�A���9[�#
K~o���[���C]+�7,�{"i�:ڌ,6�� �ǜ��(&�P��'�D�@d�??I0�	ɺ67��?�U𮒘�W1�rW[#�
�!F;�������N��Œw�7��H����-e&S�%�ؾ+�	�����u xC�R�>Хi+rSy�B>ɓ���AG1�W�ҘH:���Ow|M�A 9}:����W�M��"j����
�����~-�7
@����#�#��%JOlRp�2��f���T�%�`S)q9`��l]F����#��^	����cP>7'p腁�N%��eu5���1�d%��k��[���Nξ�
�R�'D��y�<�+샷mv;��4נ]n;�&�WJe��]��=�E9���^5��H,�@���~�nHh��u&�5]�<\��!L�o8�S��:�	�~�Ń�c��aZ��$����g;O��赚W(��f���{xEh�8.�-�ͧ��N�5�L�V��J�J+\�~X�Ēa%y8l������V��:��^H30��B,�kS֥J���,���C��X5��/�Ml��9pW�5�Uy/��ů�\��=�a��j�g�����d��	���C�8jlz�?=4�ŔZ�&���N4)Kg�s�
�P�y �\�k��2��R\?�iz��1����q�^�sٖ�ح��� �0�L��V����A� ����z�򘩊!�P�*P���~v7�I����\��w�QrD��2�`�ҽ��r&�ہ����m�b$�iJ�nm�Ո��/
����e�`Rd�
��N&rU�g�-{� K���!.�#��O���B�ʋ���L�U�Cw����#��.2���0ܔ�+��VYI֭����Vʙ��7��5��46!�%��w	��j
]�bT����R���3���y:��U.��"p�+GeC!�)��̗����Cu��'�5�7�gizx��sJ_(}���N���J+�:nj
���k|a5���U-Ũ�M����L�II�nĮ&�n��e3	`�g�rpfA|�>�C���K�wo�uk��<��&0%�]9�ׁ��v�U&q��4p`Ez�{��8it:�+Ʊ��1m+�\��B�Ǎh�b�'��H+n{�ޱs2kC�]-��Z��֜`��Ki\��fF��Kr���zڮW�E��Ty��\j��(%mF����6��V� ���邧����t�is�d�=�h}�Z�ʷ	H蚔�o{?C�Q�τ�����kr�O-����ŉ�@�Bg`0�<���;�?e�K6�}��AR˅s�S�|Lz~�ku���$!S�X$���u������w��%m�ɲ<*���x�5�έH�!�i�}�\U�HKֿ��P�v����x�賅$���������M�+�H�����6n�����Q�&��n���/��I	|#��J��UnS���Z�*L=�������?Y�/89q⩉�\��Ax�G�ʄ�c�O��8P���::H29�|����izE��φ�CC��~K��1�VE|�lhg���<�n�FY���MJ7{�k�Ow�u�_�_>w�T��7�g��m=;*$��{�9�ܒ|�1q@�I�nSp�	�m��9�`������[2]\}胂�04tV@��*�l\�k��k޶���KH�͝��K2=��$�U�z�*�lj$�,�-�g�S�|��6�+�N�a��ϐ=W���3;k�v^���̓s����o���@pOdo�������F��Z�n������"�ok��U�=�I��9JP��1lP���n�1e�4�A��#�������T��[���*�gBs�j }z�S����Hm�/�t���Rk�t�/��,j��&� Ro��`��q'����&�7o����+%l}�A{��f@��%��>UG���mg^Ǣ<f��z�2�ԗ`���Z�A�בZ�xg���ނ�]W�cQ�=k
�h�S�"p�y.t�՘gyX1��9��%jZp�ʫ�[T�d(�?ǋ(t��Q������Z��'��%��]�&
�㌞�eJf"��d�ᶛ�ԽE.�?A�\]�y�g�I�14�ibF���X�=}ڿ n�Y����ر���K�I�{g���e<��Y�A�u��ad4��[E�P2�D���ߋx�K�6�V��9Cg����ш�Z<���J_΀��m.���_x�&�6��U=�ؖ�jȾe�mer�E��Z��u�/������)�Ms�Ue��$\L���C!���W�!��DLN��feU����	��fz�����(T�*W�w�~�6<���L�j|r�2��4�fT��W���5��*6�v�������\�Ўb4��/�|o^@P�PqI��]~���x -����=39W��tR�BQ���rz�6X����7�^�ν�PIT����˵�kj��w����g�..RCh>�hh�jm~�A�ғeE8܋�|y�ڳ����+�#Ԏ��f6OUA�����-��4ߓ� �W1#�x��݃�h:^��`��G���U��ozc9�X����pf�f�^�P��FH%���S�����eB,�R�v�� q\��G�1�,n_�����A�\y	=%bL{K��]���Y���y;/�j�3�<��+�񲲀�:�bRL l���Z���V_<��������x�����V7ڬ���]�֕_�v@Y��քyG'���,��� E�zW�'�j���W���yw�(�Fʵ�3�ޫ���u�����������i�5ꖼT5�0�}����_�d���^P�R����V�"��o��O�th@�u�<�����Ib2W��xό���,�z�1�$�L�~���������r���l&�j��3�y�J5��vF���k	���3I���5��~�	��	����K�?�G��x�Z��\%T�����I.�� �	D�&�����t`�\�'�7�	���\rt2=�F�bm\�^�-/��՟�</(pq�Ŭ�Hِ�Y_����"��!�'[H�k�����&@�W�"G�v�&�?r��5e0��,��	m�Y	��`VڕC?�ǲS�f�� 8��}C�/�����M�q�,މ������k�jv�a��}b{JI�V@�|,H������1wv��.OP���`VR����&���]j�m_+�p䋫��Y�3���2��L���W����=0�D �f��y��b�N�G�7#
[ɂ䯁,q ��M��K�NN�TDg���|�P"�����>���؝-=��d�l('[N�ho���̒�u^a�A^Xv���%bB]8||X�M��eFw7��\BV��Q�}gI��Zޞ69'	��*Ix�\���~��.wc8Z�?¢e'�k��A�6�>�/�cp���w�Ō��\�OiD46��K�S���N�2}bA�喽�j�6 �q?wyݩj�����{��z7��`ۧ�gQ��h(�_��1R�uw���(�eo_�B�̠|D?O��{�酷(X#����*�f�	&��0�fD?i�SiAɐ�s��!5c�#���A��ƃ���8���6�9(��i���.�����G|����k�SΟ���l$���iL�t�8��,�a�,}q�����Tp(��P���ܜ��gՍ���`�Y����l��E0Ah�/(k6�^.�����I�Hf��G��tp.���RRS}1�v2�� ���V����O-��@�B��u��&Z��-R���r�q���~D����-M	X	�\�m-,�)¿�_�N�?�yש�Ti�|��/hVc��ݚ�f�)�8��p֛�1�*����iX����Zޓ\��pȉ������< (�'`x	��4ߜы2`����C�Z�@�h�4?C�1��L̽T��l�AW��{o����ݩj]�8~�d2B���Q���u���{�5�st��ٳ���+@�z2hZ��C1섏�M�˅x��L���LTU����=�Y�N��;�K�F\̭�]W�1��'tw�o��YаG!���=��=d�_�O����$�п�S���:�Bܬ�VL��vlLO���r:R�Qk��c{�q��мF���i���~ �t}�
y
��6��~?�_�]�������X٨N�|՞QkǱ�qLnl�mL�͠����Y�D�����,�"�Ue����nb0
A#w��-ā�ք�PG]������Muz0�m&�Yl�`�(�g��ΙCj�k�G��Y���.J}��G[]+�J�L=�KT�(���$cd�L��=��mo�%���iu#t�URu��F�( Q�RU�'[�
@I��/�bO�D�0+}4���m��wFQcR�9_�SPw��S%��T����4��W�5������}4��|Yx�/E��ku`��3��r��<HI�R��%װ-U�iq�a�Wq����n��|J;��~O�>��_�l �$�6��T}�j�.u`"�&ﭏ�
��t���$���@%���iy�����'�y�&�|"lj�^ӱn��1V�"1�
J�#z\�d�~����&���g��^"���d2�&Y8�v��e��|�}�H�i�i��D�0�W�����+p��;ؤ;���[�c�f�l�zK����EG�a8>�_�xTt8���&*� B쎈S��lS���^%�OC���$�M�=�H��9���3�2{g-VU۰R�h��t#%�' .�B	�U���]	�"
�B$��Yc�`*���L�_�3��`����NZC߼]�<0Ţ���3��e�$���?��qoҬ��Q:9��g
�Ђ��6�:;ݦ+?�S����h�	�)�-�	i?:��ܢd�F2?'��Вf дD�|��)3���k4�>�8P�鐂�zy�Q	톌�ą7�¯�ع��i�Zn�=�f$�`��F�&H�QPT�df)��;�,���L��z����S@��[!�Mټ�a�m7���9�K��'1�^��YX/�F�Ȟb�  Q6�C��۞�ȪWn1 �����A-z�v5�c,�k	�ֻMh�jU���/�JBɈҏ�w�_?�2���c�����;N���m4{��n�q�X���rZ�3X��ݜ���E*���VG��F3`�ynJ����{E����~�C��*�3ڀ?���#����1Xzt;'������7(���#>�^ɋ�<��s�аR o��^�OW�B��P���2F�̵	{i���r��5e�"�W@����>tX�T	�&n��|�29��`�<d�.]d��9x�Y��xsŘְ���iW�� �]��1���_zk���B���Ǿ!+���U��1��N��\��&mWu�%#����k4�ұk'l�{�]�5c�C�t��U.���C��y�B��=���8�0.ID�:m�x>�+kEw��j��biC\IY��κ%�m㠍��N~3G��(g?ڹW+����zV1�җ4�\�]m����s7'���T��/Cx؞*��/no[6q{a�3kڦ�4�m���(tBT�ƈR���*4�y/�q�T��B	��7<�_Qi�%،8id�/Lv��$h�M8D�dI�N���U�&��az^?��y�тT�"Fso����k����PloJ�У� �0���a�
T}��6V� ݐ�M���P~����Er`�X�}�r��V�`}V���SaR�X����s.��}?t\�ȅ`�X�f���7[/��{���x���X��L+�� GE.#s���*B�F��F��k���G5]�hhzIuY�~��ia��]�,~��ہ���t�~x�꾭���e{k��*>����N�C ��e��������O[�-G�>
r�c���}��Ô9�t�*N�����L[��wl��bo���6?��M��{��{;@��S����0����y�+���?$�Td��I1SE���,�o���a���j䪊9�^&\`/�X-TBX��_�O��.�Jb"t�)8����n���V��G�yY^7�[n�M��mRT���s��1�^8�K���-܌��
u�������pO��:�&��`�5��b�՟	�4�w����V!�4N��%�7�0t�`By��<|8kL�"F(��S͔���iXIZ<�2�_tY�ϷY>zNU4��}�F�*[bF*������7�;�.����tӛL-��t6%m !��^f�^����T�v���;P9�5�f͔.q�'G͉�����ѧ����y��'?7g-��
-C[�%K��X�w!��h������Z�a��+se�9�ж��Cx�=%�r�|4�h���J�	]�h"��p̬ ���L�/%��o�6\��։�?��Ֆ}[;�% ԛ�L������w� L5�+�-�6�T����v�y�Y�<���-�5cQB3}d�k������	�w,˝����ʊ?��ǈ����zO1yS��0��q'��;����	�s�O���-���8},Fg�i�d�L�T��)o����o���u�n�'� �C��Z���Vy8�"�~� z'hS�ql�9�`7'/z%$݊b�O ��.�c�?�]�;XꈇTET�����n�Q��G����'ms������S.��Kn+^�>��a0){���q "bI�;�e�	UP��J[D��$�*]���#!f(�)#�Ҽ�ʻ)��t�y-����>�3+��yRWA��Tn׿W���{k��#楶��KJH�ല�m�	��C�6��]0�3ϲ��;�"���¯p-��ZU�:����h?��	���Y{\��"U����A�	�DD󎀵��u�2S�I�~����f�����9���"�*���;�Vf�C\N�>%�tW�a�d�L���H���[��6��'Lx;�i�^����Q���J�q(�`�n��`n�"�k*����|�"�F��u��iq�s����=�h��(�p�t���-ȁ$x�4|�e<X��Ȍ��F����vK�[ɽL���a��o�X���jmD
�"���B����9M�y�	��c���"��=DCb�]?7�@=��.:G�o=�H��, �����UW�E��q��#�L�>�D�xx�d�Ɉ67��N�^�� +E�I����� ��5�r�O"5�*���k�\Ƿ�U
�k ����H��F�XNz��#i��8ֿl�T�I�zɶ��b����qMz6WtD�+X���Jo�#�"�_���c!��=�>zne�
��G	׾5����`(��I�X��Pzl���.��t���Ž6FKw�E����TF��@U�Op�[-��y�#N�r��JN�R��/��5��ɻ4p�7�Ѯ���?��.Z�q��q�~-�ĸ�M�������K=m�t�.���"F+5��F�{B�x��xX���;L1 ���!-��J_P�W>�` �Qm�2j����c� �"�/hA�F�qG��"�qs�|h23�@��S`�ÕN�*��ȑ� �����6ϋ������!m���8�;�p�h>�����m '�t	ʺ�V8̜�[Ǧ4�x�Y�֜|ظ`R�j�hy!��A{i��9�)��Vؑ��Ĉ�O@��'Nr}g�gx��R�|}�+mأ�n[�Th}�;4ff&��{�D����*�J;|��>����]ϗ;���[V�4S�*��_�S��Q�.�E+%��e�a��3N�Á>k�O�Br ����B?
�bo��#��D��Ӑ&��5B�������o��'��w�ٳZ�ٔ���/ �Ax�O;YQn�A��J<$�I,Y�Zl0*�����I;����I�k;�nΐ�b�GR�b^������ 9B�QQ����#� n�:2��;"�3��~�,�B[�|Q�ǁ���v��=h���Lu��rK�ߐ��hD�h�\B�&�����	8����f�9<.��8]*!,�,��� K�ъ� �^�������ם�d�w�/-2 �k�9�� ���j<��-[�d�A�~k��(��+?"�cbE=U3;�<�^/�ӑJ�y�z�ɛ�+����r�ۄ�S�ס�1uo�9�@�+C&#|)Q��q��C鼫$}g�����&6�� �i��x��] ܾ˿3�@P0��/1&�f7�<�&�(�����')�P��Z
�]�6�����Wɘ�^P����pOAy�TS�z}UZN,�AG�qOA�5�'���^��NK,C_؝L	y����-���d]��t�*;�.C ��G�\/k|���r�<xC5��"J��s?��͵c��	�
2IJK%T��
�b��1�}�R���z��bA��b���K'�ʥ��z˶��7nۖ|D��,~�Y:Y0��l�$`������]R��+�u!�V-/��L	U��Z:w��d����G�m#�W���[�V!�٬T�%�s�+��R!a	�\ n��)`#�O�4��Ya�3�m^�Шn�҄-k!sy��,~�"��u��)�G��}��\�
Ȣ���Us��0B���<�4_(W��a7Vu��94�[Uf بt���t�����b����8A��Y�o�u���2�s����:��:ߴK?���+���$��z��e��V���Y��8A��4c!��L�_XD��T=��/P�
,�l���1��&&＃ x��!���>|����m����f`�&ok�%���+���M�r�$A��3d���à�����I���#ց>̩�C�����t9(h����.if`��po�X�J1��aAa�N�ן�����U�e�Zz�Z!����������Y�L�r�H1$�@�`�VZ�,�j �wWK�b�kS�@8���d�92Tw}�r5�k�ߗo����"����mm��K�Q�2�+	X�o��zG�/%_�;�ɧ�����wҙ�]�~/�K�~��[���[i��zk�/�m� �,6L��n�h������E���;�������n��H*n+�W���eJt�ӓ�w�%��GB�<3��M�n��}������#G0���TI����hO�6��Fʭ}k�T��HH����	�D$E��쐢L�co	e������*�#�:��g��G�����G�$��t��!����h��{	����\,�1o}���w�d������^wx>0RzN�(1)XHU��@��]�������
T�1�1a���%J���w�Ǵ�/Q����M��J�jr��
,�5ȗ����SM�������uu� ��I�a91+\E�\'p��e�~�Λ�G�$�h��;R��X��Tr�	�X(S(��tC����c!3��Y/�}����w��kNK�i���	�bOTJ ��M|��6�̷arQF-�u�w�|����X������M*r4{�JA4ˆ"%�6�yZ��IH��o�2	*:����=>;]E�G:`��s�-]��o��9�"��)x:�����&�N���k児���	�(IA[Du�AR}n$�|�������IT&��C���\%G�n�4��&aJ��m��=g�;��~Ќ�|�ծ��O��g�<A9�FcJ$�"N�W��U���A�/J��S���D�>7��2E�־�|$�&Y'iLόsE�#�o	[o�G�h��&*����?�%�F=�׆.�gG�d�\�j��H��R:��A��C�0V�IN�_�v�׊<�>������iw~d�(�lޭ�b�h=�<6Ѿ��'3<���&��������������Wn�]8�e�U�j�[^$^@�@8rZ�?��'wW��yS~[��+-B!�<��EA�V����.�N�#�n�8oL�V��P6�>����@���Zf_��k�Sooڈ�E:Kyl�O���e��Pi�^�Q�\�Y3ʍ\K�i���愒H�zc)�`4�ւE���5OT��m�M�g�4�E�aEʬ��AS���Sn�ȁ�xҥ�L�B����D�Ud��Y��ڵ/��.�l�pa���O��� -��Nbgb�{�i�]%�N��Lx����7���ʤB����FV�Ϥ���b�5���褽��7B�(�5������X.%=�2�S�5v*����a�$���N��H�	L�p���QV����h鐉�i&}�y= ��Α@[|���e<�-�d8�L�F�|Xм�mc!�ׁ0�UaMYg�1�kDM�����4�y����F�+��k�V�2�)��h�7z��YF�\��N,����x�;F�#���o������� &�
m�C�ΰ�|6�%�ʛ
'�ގ�d�����* 7|b�V�x +� �u�'�1�_���K��G�G^�U͊+�����B�p$����&m�lw� %l4zٴ��E�HeK1ާz�!(��]
)��n�� ��hHƕ`�r�)��BV����d�k\�'ØPٝ��������O-k�?\܄�H�6l�Qyޘ��y8�aNU*H�����*�tu`��@
��x�}��GȞ7��|e�Inqc5#�Y��}��޼�k���o��F
G���H��)�ιD�&��h]wJ�6�@篑�o.�����,#|!K���jKS�W�`��GN/���~�j)��r�&S������gZB�>�t�~���r_��#�n܂�@�����/|�B�M�7-�=�1�h\��	�o�cI��;��(n�Z[�pw�׹XULp�u�����x��n*���j^�o���XH2�bxǇ��)�����դ�i<ܶ��L��3!0cp���ƈļQ!�g]%��NXt�Fʄs���[���9Jﳍ�D>G乢_���#;D�%����<h}aͭ����,*ϊd�R��w�M����h��B�j��T�Å~����C��9�|���C�@!`? ,LZk����Ȑ٢6��Ҧr�k=m}�yy�F���J��p3�7hΦ�����d�xZ���	��q����s>D�	],�7 �Z��r��*�CK�6��e	x"Ur*3G�j`LN��-j{�ЍyN���TV�[�I+��8�KJ��p%ʄ ~��Yl1p"eQ�F�M푨�|f�d�$��7$r�vh`���J�Z�Sj�w	���8��$z���d|�����ۥ��L�S[��i+'��h�'0v�v��@�[^#�.O���,����M�S'���i��F��NJ�x��s?���yN�3��K�+�<�Y��!���������T}w�hCApI@m��?�J0�K�:���q6&��<dBQ�>��}�w����;��b�P�l�����9��M�0;Qd\O�A������xK����d��2���eu�=� ��
V�đ�����#�no��CZ�&#H{
5�b򣙌��ޢ����Q1��pz`���XW}?`�t�@������F�R:,�F�e";�T�!5gv:�4g�� knV����_�y����b� �S,vE��pLr��e�ة��Q��@�V����K��zO��kQ;�Ik:�d)b���:@c\{�h7qՇ���Y��'���!��3�wl����ÿ"�)�^'�f_ݡ��W�"W�H\Hl�H�#�q"����5��o�C̃�s�H��|\�}�؁���e@��]E��W�%��.�|�L���XT��'�y;_��<��`���5�'��K�GN9Q3&�v��h p��L�Ȇu/U3���F+\0e0���;ܟ"��R�Z�7�q
f��T|(uƬ�i�F���*���\��O�`�d1D���B��N𑃟�3��Gi{���R��h	���fv{��k.�}����lYP�V���{��i�g���/�N����Td���35��x�t�1��Ņ�o�ř�fb�S�9X�x�--�H�4m`�bGn��Cx���R�d~��s�9HfI��]���N&W��_*R�ϗ@Ș,0�ʌ��R�M2� �$�h����be'�FGJ���h-���_������b�I��ۣk߈�[M���W:��/��fW��'�.UV%��*]Ѧ��I5�Pz�R7�����6����Xg�ys]>J
�L�j�x͠�닆��"�L!;�c*^/����Pg�Q}p�|�Л�%Xl	�FR���>9�5�N�q����0a�=�!��x������ 1L�)m��<?�E�*��I���ǩ���i��)�����A��� ��_�	��<�`Ϭd�=W�<"���$�a���"`�q�L��c|N-3�%"g�����]/�/�Pn���5oCt�ТV��1P�X��>*�J��{;�r�㢛���h�NR��٪U���4XI�Mu6�X��f�9���)��X���58�:1-�s-Qi�%���$�3�W�W	F������m&tX��>�:zH����S���~i�ec�9 �b�n�i�k����_(��-y��O���s:�}`�œi'��4��A&�P
ig��]!�z_�#�t����a��i)�~ifw��*�yt�J��*��k�^c�P#�N��
�Ǭ{=�Ό����(�#Ir�lύ��8�-���3����c�\;����x:J�c� �J��o��'x��[1Pア�&{�AڭP�?#lo���(��������|�S�63�F$~�����,�[�¶�s�� ��:����.뢼��|���ԀVM�Y���$�k^�,����WGJ�R��z����>{����[�c�WJ�ԇw��`��.�&����ھM;�pӆf0�-��hծsL�ɠ��2b��}
��\>oc��~�
+���%*j�$JQ��5����]�=w㛔>
�80��$��V��ڊh^�Zx����L\DP.���sBV��6*���mA�lf|���+�S���+:��~o�Վ��`�,��b���٪E��?oL�@@_ny)KѽIF�s�	���4���|�;�'�A	���_؛�?��9�������H8�R0?.0|�
$���F�M��f!P������2v2�"~�u,�A`H��7���	�Lv+1v�y��q&0\s�B��D���j�N��Ē��k
���u�3i_6~�c�{h��^���-I��&*$4�I4Nʅ�,��2(-Xq�saF�����n�����|2���U������%��x�(�:�[7��[�Z�Og��Z�3��x;��-4��J��0�d�X8�J����e���:2�@�|�]1b֨A�G�[����SH.lG�2��38Z��d���|
)�����(�1,=�*��+���P��	�_F����wV*%�=����1���Pj�x|���.��s6�!�ݕ����٥��2�E�Ļh8V�,����.!��ӪΫ�7{��Zw5�H:���_�[�&+U� �U�G�%���Q��ʰ�52WpMS��8�f��&4� u�!~��dHԚ޳�f}}��;[�+K �nB�B��V��~6������i�Xp+=
��X���k=>�k�ٔ"�tT;h����C�D��zJv��}F�Xjm��潤�Z��/Tw���߁{Qf��l븫��+�%�M�&n$�:�����8��d،J����%�f����Ǡ�6�sK@���+��&�]�Y�{:o��мƏN��h�8�OA��'{_��s�.�<��Ly���uU�ߖ�	��S�jP���41�zt
�۽��G�T�N�H���gQʢ�����!�`�0��{����M��� ���W�??��{�R�$<9'�Kohz�ax��и�.��)a*zX����W��4;%'�rHC����B�d.�` IW����kǎ7u�eB������Z��0�Qgԙ��W~��8�۾�,��D������r��BW�D���(�ʽF�թR]PkN74���*W�:��6j�R�x)������#H�6���������<%h����ȑc��m�f0֗����b��6���2IAٗ6Ba ��h��FS��l�������E���fs���Ё���N'�)����-Jp�B���1�Q�9]��,(���'�H+Kq�6l?M��;��ntl~���A�	%��g�ҏ7�%1��}�i���l�~aON:v�5V"�̀^��ԖnaN��f���a�U������̺c��"��a�Z�Upc S̽}�~ʁ�m[��,��V���aϗ�W�0�K����\�`��5������e.E��
BC���DV�J�6�	�+Q��O�ܘ�)�}y�"Q��C�@���^�\������_)�x�
Of�fe2t��2�9�6��J_K���=)��+Q?S(|�0A2\�DbVY�����X�ƽ� ҽR}?昢��KXYE�h�:qB�c�]\��8W�U(�,����d�;K�V[���᭽z��A�ɠ
cDRG+�.1hd.N�4������%��c���L7W��l�NO����GNȣI��{�+�jȠcuWS�59Aq{���T�)���ٛ^����M��B2c׻��r$U1��EU;q7<~��lVQػ2׭��4���e}j���pYM0ܵ��^,} "��xk�؞�¨�"D�:�8*�3�<p�L6�T��,�0�۠c�q������5 .��ī07�]H���@�aa5��RU#�N��S>���ۯ��+Ch�٩���@$1�8� �$ֈ�]�ז���(Z �M�pr�~�W*�F��_�j�z)҂�Dl06c=ਰ�:D��"�-�!R�#H�fi��b�V�/�	F	! �I{�yǲFA�J����%Z��� �!�gh�	ɻ0�W�i3\	��/D��>����0�w�&������ɻOl���U�w_BXb�jPib�
 ��de�t��t(>�Z��a�q导o��}Iz6^��l	���9r���8�����ј�P�'I�����}.�ʸ�+a�
x{:7�0�Oo��.�R�kR��@:Q��ć1�ST��5R9P���{�O��Kd�@@:�]J|��f���)�x�n���U�,.��ee�F|�W����.B��g��^L�����s�w�V&K��@Lr��^I�0f` ��KT��=�Gqh�,>�X���![�f�7�I[����	�4K��$�t���CŠe���Ж�� &Q���ѐ�Q��/�	�u���u\���XS���䳇��P�v�)reT�%w��(Ss��[H��vYYa'���3R^�j����jqt���⋗�����`���o���:'�;�{,�`��D���4%�U	��n����܇�C y�� E�˞aZGX�Ց(�z�O�vS�-jC?�� ��~�n?:�`�d��*~)*p�0����4��e��HSO��S������r�g��v� ����w_�}�Ú��<gP�ݠ���v������?W���t���;��6O�8�{&���/����Z'��w�6�v��~x* �igd_,3�X�z5OS%� kY�ڻM�ՠ�k����l���i�H�}V�WL*�ǟ�[��Ǣ��M˩�n�̤*m��PD���T�b:
ڠ��3��]��D����
��^���BJz�I�*�I�:7���z7�D�EO~����<c�5��{�BD�3�GǸ.���n��������vȣF0[g�}����M\eO!�[��nY��f�ŐBۯ�!�Un��C��7�r�)]q�^��2��3H��v�Cs���V����w�x�j���`G����cį�.��o��`���Y���O僯�C��v.[�
�A���^V�����6�s<�Ta̱����R{Ti�5b%#����x�R����-�R������K ���Z�I���J3�K�Т���'�Ðu#��g^��o���z�@�g��ʎ�����?���kzB����o�P1,�3��7���N`����:��ƶRl�`�2:��`y�k�Z�iv��3���!���@���_�94QDƾQQ܃���w]��B[z����<O���no1�[�MM��+J�k挭��A��u�j�x���i�@�v�=��D�;�7l��X�c����������>jp�b
�P�x�G�H�gY� 7�K�m.�N9���9<����Y  �`����M���{�A�Q
�$B"�ǃ���(�5��
�鐇}W��箑�����r��&�F^P�p>R/_���΀����y
{'�C��emX�
���jɮ�����;$����W�r?�p���V�\h��
�?@������i����z�(IZ��ѳU���to���&�i��#���;X�E�����{O�T�2�C���'w8��A@��)�b`�/�u�kw���$<"Ͽ<=@�X�iD�|�x�e5/� ��PΕ�@��2��'��z�SO"�&�����S'T�2D���,�_�Y�|�{[�6Ig8|̿M c�Ax�{��sI����Qtb���M�c�0�b�]+v�$@�_�m���J4�3���	�6ǟ�6����6��1]%u\� �#�Y%�j�h=��6-h���v���^�̳g5�p�����uGVF�۱�l�f�zGД?��Od�C�r�k*d�=B�
z���`�f�S�&�U�+[<_��Z���K��k Hs��[��5�V4���H���a)+��.�$��X���e����N��A�����k�R}2��F,Z�P��:���&�@����՘D���� k�����s7)<�v�w������,��ѵs�Y� 'VM��8�KV{_�R��Q���p*����U�It3�i���.��O�Iqo��m%P�M�j����<�w�Z�S@�乽�hރ^�Da���!x��+��^k���$��k�OT5M����wFs4m�c6G��s�/G���=h������p���e

��J��S�&�҈���l��WUز58�ڴ2�Uؠ��f�f�B�f�?���׋D�֚ �U�p~���������Ӌ=���c�=���}�
MKJ�����'WT=��'|����}�6L+�o�E�'� �K�Pt��S�������~�����m�؜Q�HT�����j����m���6��Z>6�G
=�M��}�/M�{������Jh�q6]���@��c�<�g���~�} ��d�#��e`-���f�N�0��('��T�]�`�s	'ug۟��ks�`�wG9�T����z(�����X)��Ѽ���Wz4۷���|��F�&���2ϕ�6Ba/�K���a&;F�.���r�yW~?��$���"����ɋR���e����"�|�� E��;V�)�8�a���B}�L����_4C/��	8;���,⫒�K�2�<!7!�3:ѓtJ��;�"�e���h!���&љ��xf:G:)��c�N��NT����s�J0�6�?R$�gj{��[�Xu�fj�yS��vV_1���M9����u�,�K����K0�����n�{TZ��2���~��c�:�T1�+�<�D�*��t@v�M�e?�e��%+�-��YK�w�"E��?�%b���-�M��sփ쟑�.�'�
��:r�EJP+��-ah���	���e�R�A�X��+~��DP�r�f��%v������U�.@�ڏ~��҄[Ӱ޵����0:���̀��̬��\ )�"o4�*�S��B��s o o��N+�l�}�(��vÌM�* �����Q�)$�0�BF+S�Պ���E�J깧u��,W���H�G��e���M�������)��63 ~q��
߻_5�5����x�^��|RFd�<�*p�:_Jm�D��K�	hg�������x�m��k@J'G���K��%�����8�w�c��D�y���qTi_)~P��b�f���iP��֢�x�lQ1��&���d�N�x�W�a����CiC*��v�2y��*�kXfY�v����a����b�U)�a���_2��-�Rɕ�5�!\-��m�m�<��/��z]��|GGA�����g�}`$�]��۩!�8���S�6���Z@���t��2e��%�:�	�6��G^#�hChP�r�4�C$	����z�Q�&� ��F��Y�&mC�F�n5�	hC^�i�Q�=>�^���'�\L��J4�W����U��A�>���9���U^���|��Z��I.E��68z���~�������V� 
6�aC9��a���HȢ���v�����c9�~W5G%�0���2��1U������X{x^A
r����->��b�γ> ��t���th��Z�]�Cm�̰m���dFҜ �b�p�˘�gs�2��ˍ�����.�,��>��	�:�8;��N��)^ׂ�#8��{�܊��b<ŗW�9FV��N"{������1�w�i�k`Ӌ�!��x�'Z�L�!Q�Ӝ`#]�(໐�ΓQ-���'4��u�G�ݟD;��D�c,���K�ɭ�XE�ݦ���
��͕z�D�'�}�/�9q8	0�+M�S��_P_P���E�7Z�Tf������DT� .����
k\�xu�s�l��>fg�z�t�Vd/d}f�{���)٘/�x�
y��+�,l��f����x,�8T������b�Z���-�]0�.�l�>�W���w����9�Q�^��`
#�(�.���c���sG �Q�/O�U��@���C�X`�bF�D�w{���$��x�O�
lwP=\�6.Kk��U$O���+�wN�������2u�m	s���p�?��s��'c�{�@�vV$q�������]j��qP�O�����̧��]є�[ߍ3�y�/�=k4	g��2�-��7�D�(A�I A�9d9��4�I�.�s����b����i0��;�*��2ѥ[Q[m�Wg�;/p3��@���$�8�o�Cj��d$;�E�ᇵ8�����ֶ�9vr�&����^p�YEk�}8�0�ǽ�o��LjVH3� ��d# <3\�X�B���F͢H^{Ea:�h;nj�w�e3�`9G;o�@�>��	y��P5%�w��8H5�`N�p����H�"��ˈ՚���2<R�ɖE$���=!���m�)g"qrCf{
I�|�t͠e��U٧��*�pN^	����e�F����C���ޣ����j=�QTK�k��� �V����o����n��[�О�~�Ē�(������g��y!����F�N�N� :gn���&qK��D�4<3^V���G�|�ۺf؈g�lצHi�ԉz�R�Z����(kDlC�G�Of�h\��'���>��fR � r���Q�A�x*��OP{�ӧ���@ h�=����<����iU�~V%<\��#��)_0�&�Mrn�&]��w1>5f��p��y��UsJ���m�^н�`O��GY_Xs-���grI!#�oz�:���A5�|5�>��J��C>����a�����y$�.虓�tM{��wͧ:�N��w� e��E�Ni���;ܳaf��}"�������!DԷ���e?j�Q�ԇ���v�"ʟ���y�Oy���O%�$h6��p���R�)/�b%�y�R-֞v��Hj�r5����f�H貕��)���>J�j�I-o9m}���F��K���0�,/�#3���-ՇF��\5��*F3`4vh���r�1i�����^j���Nu��1(���S�'<"��a�f�3ܿl�ߡn���w2S�|^�Zʻ3�XS"U$�>a��w`W^p�L��E���F��̌V^���⽼����Q��y6��P��AX���>-,��an���*��Z���� �s3�|��T��F����dTN�ǚR�ۙFP����g^Ȅ;�WK�o	%no.�X9�E���R1~�s��Y	��R ����բ �搐�y=<b[�ɸ�"��<V��n���uW¤~���z�=
�c|nc�ZE��rF�jCn��ai��[�wȋΉ�~�rOO�τp�uE��C��au�P`�4[����~�|��%r�����/�=ˠ�BT�β�5�<Qݲ7@+�J�]$IJ@$|g�U:�ߪ�gO��P7Y7Y&{����I%��*w��ӫ���u���7��oE�㼧8�ec|��Y7� �E%{�tZ��),�x&�y8�����G���<b#JG�]Rl��Ƿu�K�2�#��=m�3�W!obI��é�~�Ze�x�.jИ�F@����/�J(���ݜ�=]!s0�jf�0e��1xi�:�[��v�qoЬ��`�Y6�УxDI�̉;�ء�1gc*B����3"���C�)����<-}��h/�8G6Q�,�(�~��v�>��Y�}H��Ls g���������)R>;�B���qh�*?��F����@���P�D-���� ��G���&�N��hpx'���s�[������N*��p��df�>��l�� Ψ����?��[�Dh���R��E�4��S��)�ѾT��j
�h�h�-�������b,�졸(�[	@����=�	f�P�!8���M��]c�vLTf�Ճ�6��=���B�-���&KQqw�.�D����&�\�P��+,�{�������MDq�g4ix��Y�\�Av�����S�����Mm��o� &������].碕�_�/D�������^����~�����5��D�r7������9��q�瓒�6QN��Xj�ꢢ*���Dg�/�C���#�{�1g\~�w���:!tRrj�Ծ8���c������� �.
 �E��+���51�b��h�+��&�PI��ԭ���3��_3ڧѿ|?n����)A�[��85��<g��TQK��Ѽ�r�-��2z!Ԉ+v�J�q�8�Q�"�O��Xp�=�,��4�TY{0qm�٘|������"�S��-�2J�(���ƴ�n��Y-��q�s�� �����ě�:�(�^�
k��X��s2��R��VT�[�L��q���Cn�ڑ���,�������d J��q ���*A��j�� 3�d��ߋ��	�$��m���4��~��+\���B�q���?Io�5���F:+%E`���\Jx#�s�
���O����H�{%q�Q�E�t�پ�F]ͪ���� U"-,���y�A�lS�8*{7W>a�S�I�oA�$��ϣ�|R86���4��P����_�1�-T�;B�ƭr���v��s�B��
c^��6�Ti��r������c�2t�V|%$�S�e7` b%5���GԜ��٠zȄ��U�dw��sp�@|�;(K6�u'�7^�N^L�yW���	��vMV�O_;	%��[��ٴ��P�l����lZ�]���6(҅7cVzU���$c[L�c��הY�0l����.�	|t4��8�P�T9�i�[�2	%A���bN�
4��3�{�vW�����Z��@.�c���E+�/
T��@[�v
��dw�%����cc#ާ���8�T_r#	�GO?�Al��`��#/���H�ʤ��9j����t������oKj���f�=� �r������mI����*� ����Ȟ-�� ���"h�I�|ҲQ���|ɝ��x�m��*gщy<V�͏5nC �O��ݡ���F!�E��,�l��� :���s A�a�0;���4�w�ÅZ�4�o���'�����4D�@���⡪�.�e=���#�0�H�p"���_n�7���jx�mR>�(E��+z��������8+d�/2�]G�g=V���X�?�Q�8J�]'h�X6t�5W�o6��Ѹ듨���u�a�
� ����O�I�S,��ι�.(�澲{/�呜̫�{#&��v�^�4��	<����?�S۬�BYTMR�:���Yi&a룈�7�<�gO�Ub�Ry�"���uF�AY�x�2�Z3Λ"-c�,��i���6J���
>�f��nK 9ZZ{��}D�>̇���s���pD'�ý���W<-����#�0	��Y}"n8P�����_������'Co�^�	���*���%활��"� ��z��)����������$#�����Z�_ԫ�e�4u�����"3�9�XVXH7.;)�y�a���˸�֠ƚNp�>�2�dq��\��ġ�b 1�I��`��ւ���J֠���Ф�t�
����<頴���k�C��Zb{�.�g���<��f�Xx�%������ra��:yo��2���Z>������]Ƞh?{�f�tk3?��;B�#�s��s!� ��Ƽ�	�#��GVx>%����2]�?j�ٵH�`�:�q�.�n.R�DY(�jd�����D�ma��gW8�?n�pҠ�s��t�ۮB�[R43(4D��+���o��t���*��9Ȳ��Y�]�J�=�̴!���я��ɡq�W^�*F�~M�ߖ�������ۮ�c�*t�Z�p���̬���=� I�7�� 9s`(�l7����I�r3�[�[�j��)����~��Dl��+@�?�vD�e�
�:\���]1[��ib5r}e^fq��Ǥ��3 �+�����<�%�;;����d�����u��Ym�W�B?�u����6�A��e!��ހ}�H��YX�~��)��~����v��x�j�8�%�F�*�WM��\%�?��Y3YwKj1J��X�V�>�t"K��T��D�(\1#�aLq�~B��}�c2���FD�y
�Kf�q�كy[sFHt�k���2	�q�*{�oPE�Lؓs����e�P�/�L��o���Eam%���c��o{��{���V�*#5tԙS}Y��5i,L:�-[$zBx0�M������z8_�sYZ=�a�NL���d6��zo�[Q��*�*Ez�M���ko������K���5ߪ��%�`�p����"�Q�ǻa[a6�8ُ�j�J�x�2l+<�����6��C�:�z}�+���nP���$B\<�ur��5bm/�������g�����%��~�x���2��fVE{�uz�^�z���=�b~N�R��\���V�g~#�s�O���nt���}��G�t4K~�܎@ �O!nU��S����1��Q�tp0�,��k�1v!\ϱ���.�f*��G�;85�sR2�n��Xi���`N�%-Z�@��E"�'S��>m&�aZ;��_���fQY�yY	�f[8W�B����GhW�1���a�#�J	
��*!��E@9b5A��2[�r'=��8PNթ�����8����{�XC�%&�ۓm#c�%+`���K� Bn:��Ǣ+!��u6����s#842�a��j�]ĄSy��pc�"���կ�R&��X8���.����j��@��߳L����������ǩt_��*�F����t=~Tl�@KĞ�5]I]��ȌRC-f�񌧪D��E��1��
0�m�����X�2؃��{�,DS��]�An9��jC���s�\���kR���m�z��4姎��u�(	[5\c����:�6|��@_bBI�������+W)���5���G{�Њ���h?Q=����7��<Tŏƽ����i���xX1ʧS��^��b[u3�7�\̼����m�)��{� ��&�,>8$E�Gk|�t�|��B��t�m�Bq��X]`5��ih(f� �>`��Pz_��Y�Jy�$ztE��H)I��D�JD�ɭr]/&F�0�h�g���|����\��IKZ��]E=.�.,���"���?�;<�S\oR-�m�(�&F��6t�����F������MT�`�/*p�`.���Z:����XxJ�72��b�v��n$`�ތ0��S�5��z����2���r�Ӯ��$Cj���g���^�>pK8gz~��ԃ}"�`���s �$x�_�� Z�iS���0��"��c=���%C��ǬJx�i��2c������ɝ���C�OU�e�j��4�U�C�֜o�>u'���X1�.�u�Н��B�߻J�J��d�#��n	�|C�P�����ߵ}����8Mj�q������]$�``��'�Xus>��J����{/�����sY�Ű4=n �T�2=��yOj�	p��tA�X~3"i�(�(C��e5Y��!v�"Jm�y�k�a2�7 �j��,�}�=.�`�]y;!����=��yX��qV���f�w*�Cq��E�nq.����T��jMR�%Gu�S=��"���Ax��T*Z� n����C�!����G�a��S�k�d��7(�8Gq
,8��,�penI�ic��.� � �"t�MS���1�����m��5�J�4W��້���$BQ��S��ꦁ�3ŗrp�A�����jM�.3�E/�FT���9�3��b���Q�\mTO-�`5D��6�=�!Y�6��*+~,Ŧ�;���* :�EzY���72I����W3���@^�q9��`�Y5��j�A5쨲���Hо׀aXI~�>�[���U�P�B$����A����9��^��-$!�5�ʁsx���Lq��E�]c&т�Ic�#�v=�ը�	�X��}��B�q�±�}��,�z-8GU��2��dR�f�_`"� w��/�(��t�»��ߪ=���\�d�rK�я�V���nW�������<�{��YBA�)YN� {a��
���G�����`�����yo�KWO������5�����(�yì$�U���w(#@ZlH�M�?���L}��#:^�r��W�(�| IE�N�颚#��H\ie���oϜ@|d�~\r����&� ���<�M��FI}1̯9s��:�%uy�Rf;��UfJ����/��]�խ���Y��}n��H�Q'\	��Ki �0����uP[=�K#9���˥�aD��_N���p��"E,��f�x8��j�q)lN�x	���!~~��0�̳�c���3�9���#�BCB�0svH�����s���{�2�<M�'s�W�P�������v}�y_O^O=�d���s[��ô-�bA.	��f��!���� ����$�z*(��Be��Ǯ1"�'��'�XZvԝ��W#�Q*�N���֠���)ĺu�ث�U$>�W���O)�x�[zr�J둶(_vۂ�04Ux��j8�\t�9�d�Xb/j��"
v�����Y��������	MB\Mw����5��11�/-ו0C�w�@ɷP!�14/���ö�S<f����"��c�����YiJC�8?���c�au>�'��IS��M�����Z4���% ��KC�Y�g��d	�X�7%� G)7�̉c�j}��v��~����H8S`9e������o�2�Г�;�>�<h�}uf���$?je�� 
�ɨ3rV���3.�\�T��L�*h�Ne��$f�"@l�⅚�!u���&�R`�<�ɱ�	o��Xe�����䚥��l�+�/��1
l�v*�=�>B�aJ��Pc�_�c[$,��hS�"d���0u!>J#��cf� �C�A�l-�m̃�G��_.,{q1�z%�*>�.Eѐ֏�OvAJ������U)/u�Qr��D�9۫�䞠m@w�ң��"��5�V[�uW-��@r�a¡*�eX����3΁%�ߧe
ZM���WcB��t����2�f,�Im.�t���Hd�8�_��2�L�����QQR�V	���`�'S:<��t�]Y~/�$�!�۳���B��AQ�/����+��70ҹ\�k�B8<�K��w8K$��Ϣ����n�+��e�IH�za��[s��K�(ոT���2.�"O�����HJv�|��]�|L���]��5Z`	�O.&f��U/�eY1
llBɿ���?��:^CVPg+@Uv���Jk�Ht7�)A ,�A�o��(��t�s>�=r�"���kpԛϏ{G��J$}\S\anv�T��j��v5"�
��Jƽf��M�m�Q5�Q�۾Du��������x�ڥ�hQCn�?B�^��^j�Q��;t�[��2��Lz�=q% ��58@�漄%�F��"��%�k�#��G�Sv�g��2W�?h#��Ew��AQ �?X�V_#0��hI� A٬9n�����ڼ��7i4�wl*�$p��ǩ���a�W��aT�ڏS������o�GL�ɒAD������<�'��:��s�����I�;7�L�l�@o�i�>�_�d��y.�׏1۞I ���
�99�`xiS,�)��T���L��o�A!��/Um����y&#��a��ak')��%;OF1��������6���ɵ �R%\{�3%V����x�~8��[�iC��&��Җ�m-S�F�]iD���*�1:����s��!���֛�.�3���"T1�Jʢ������׸�֌i�v�!�(���Z��8_�4��H����D�V:w�A���Y�h�xs���+�&f>>,bs|2�j:��.��l�6���#�/���Ñ�R�G䎡�I^G���g5)�Q��d��wԎ�˪���#�-w�|���\�gL���L��^���_���,��-�>Q�xez�߇0?������u-1a=�e�sV���S�R���x��::fr���k�D��j��7��!��p��O>fi�299�������au�9Q4y��&����c���L��@�� �:lS��Q��"�h8t�T�\�'��<(:���m���E�Y`T	�K���ѧ"���F�x����J����$�քB��B
�h�+h����y��PS��L�РG-0�����8'�pSh��pN��ifO6�U2C���+`�{�^��x�A�orཻ���+�Dr�r��ڶ�{O3��2d4�0ձ�ط|�����X�wus�/�I~v���H�'�k7 SLl$�6S!�b�ت>KЛ�6\{�\%�J~�����?�ۜ��F�&?��č�[.A�މ�f�}F���]�)�/��n����}ݵ�^D}��� "qM챬�;����Ґ,_]��@���[*��/���A�:6*�c�&i��ߥ:eU����8Jԛ��V�p�}��T�Y���5��.�zQ%���>�|'l������)�y�L@�l�՝�h7�����'K���;~̳���7� ��I;�"of���@2��$���8��Pl
F�9�ݟ^���������R]������!a�p`}�v�~��`~+3M�Wb'��3w�dF�:� �����
/ʥ�z�Kܹ5����'��q:�
O;���2oie�}�:}^]��)�'���e��󮋀}]�;	�jy����@���$a�'C�%W�(����!��jz}>&M�� D,��$�P�_�\]T\۪��$n;�x�
����PX��7aن$ٸ��`oM�v&	:�HMWLk\w����8W^r�X���p[AwY&KK5������G�}t��!�����B*lt��(��)���V�������P�=��$$k2�
1���}hq$��dN&��D�f��L\�8L�a���eF�{`�$!�=�sE<	�q!�_�f6�^ �/�5�-.}M�T����وߣ�(O�s��%��\*��e��#��<���Y-��`�:}��H@�g����|��R7�L�#j�����.l��ᐌ�-�u��2߉��׽�4�Ě\�Q�B�n-]P�N��6~ �k�.���ze��%�K=��T��Us�g
iIޙ-�j,5�i9/����bu�EЇ�u>L�U���+V�i���{�<C����\D���}`���A��C4m�_yLN�O�&]K��H�~���R��;�R�V]�(�<�#5Mʿ,̽� =�r��j���C�8�A�+
0�2������"��E�PP��'ׅ��/h�z��MW��be$��w<������Ay�a֙�0p��J�'�E��T�����_�4C�"�%��Gs\�����js`�,(��r�c�����W���/�۫�z�q�6��St�RQ��w�X��a	������c@��o��M�x������k5
�깇70cj�Ď��!4��7Y�^'.�Y��{�P���x$��K��3�HXy�7����K$e��^%98�7C�U#��	@'8Ұi��S�Mk({3�Oh����PYͅ>qo��||��B>�G��mnBs���<Om�م0���	"B$G5�x)|3l��2�J��"�D��ə�ֳ#��;25s���]����MC^,���:ы��6�o�n&2?��b'Pr"{���_��D����G�2c�Š�a�X���/з�*�.�N�5���:�uT�zY���9��ܺ=�¾�W��� p.*�,�aU��g��^17z<��(��ñ�\��t���:R���� �f����:l�$�KJ��Nf*p��!
6�MM:R����3?�|���)��+@H7���
6<4��-3׃��P�g�qȯ%?T��^S�����a_�G��7���o^}�����́�D�4A֍������"O����ʺ����F[E�(�ڀju�n�ri�߈3<&Ҵ���J?������U�-]�h@G�f����K��V�I��Ym�r�"9E7S�T�kJ��բ��{�X�>z��(�Ȭ���2��-C�	�5��7~�Rᶉ�d��^Kj�rxi!;��Q������a���Y<�� ���y�]Ͽ���)���n���T'����_��$"�h��j��=�:����p�|� �䤔p�����"�}��r�;��%#�O��b�"����.��Ǜ��N2�f�����$j8��ج.����\���-3D���!�BBny�O�g��E\$�}�\�1T��Ǿa�x��?麑w��u�ЎV	��Ӹ�v���"$��M|�oCY5A����>P���TYb�ZL-��o��ޖ�»_)P����+�\�U����q�T�7����4��K�"���p[�W$t�bG^h�j48�-҃7zv
��Cd!ا�^�T}�ܳ��%�έ:*?N�b�����ӆ�C���� W��.���7���օ�N�����x��ݗ�����
�[���I�m���x	���xj��f�H�Ƶ|,݀�J����귾#��i��S��܉���XX*���u�To^�7otQ����q��A+F�H�}�d!eG|��C$��Yp����o1 �^Ȭ�e��k?���\%�����44*�F��p���۷P�
������4����I1\m&���bh�Y��R��b���A�e���ةQ��R�aîbd������At5�N�ƈf8���'^�� �Մ���&�O�c���AM}~�hZk@���/:�$�Oc�Z������a��/��i~�2�J<�,�&M��T�����*�	�\9�%���W�WL�Ѭ�uV!kAr�x4B�tJq��0.o7&���ť0�9�l�69oq��O����INx��z�`>���C-�Z�'�vQ�f��hϏ�р�}@jT˖Rz��I-6/�d�rSYP&z�_
)fO._+�`o�mC��!��;i�m��|��d�v_��M�?������(�b𫱷��������¯���BP�eܒw���#'d�#z��!�}~��ϣ��4cI�� ���A{�Z��/)��r� ����ҿ`�
�$�$���[��B;��o�2C�%�B�f�-�Dj�o��C(�ς�v.�C�<����Ě<����}-�T���z�'�r��2�C�#�d��PH�*2�q��+x
��6�R**��� �����2Dj��>�Ǘ��RN��M�;�����҈;�r�ze��u�����O"|X8��/�g� ��j�Gd�`_�����'�Y2#�������>�'�W�����(%�l�-~�DT�-����kV�7��|F���,Z���^�̈�@����ҫ K��?�����:��㇋w��^��#`�0F|��}|�)g�+Z0��<X�1fP���=[=39��1��&s��J`J<"4�
)`��uV��ЩA���[��­�gr�|S��&�I[z�7+ ��'�-Y<��S���$�Ğ�@���Uk�;�s�ჹ�ym�7܊��A�4
���k���fH"��Ӻ��h����n��3ޔ_�*�	o&7����5O>/���WM�H6��~ݭ���E�O(��Zwܚ�GN0D��<���J/�5����M�,�k��Y��)ƿ(0�M9��ڿ,ҽ���2^gB������$�	q��(����Z�w�������y�Yx5���E��j�[�FbuQ��X��u���/o+���#lo�6t�a��n-�x�oFİ�L�b�)�(���~�#ឳ�+7.��.H�J��B��p�����,h�R�:��u%�DF���,M�دS��3��.I}�K촴F�.���u���Dw��jnާ��>h������8�}�m��)�oF�������U�~dz��C׳��`g�J�=m��8�(��R0�)ۺ�B�o<Am��gfA2�Z*���=�@N��_����
�y�Y��=ٿD
񡇞�8�n.�!Q'�J�0(���;�P;)�Jj
CD����]������E���f��o�.�A��"��M#�T�M���}�k��}Ԩ=o�Ry���v�^��n���G=�0�9O�>9�kѥ�je�0@�W���pL��}l�����%Ix�����v��>��m�/�_玦�	D��/�Wj�#�0V�C�k�W�H1*˛�d7��B^��R��q���ޖ�R�3|$�<�ق�a��M���(�n2̜�t��,J��w��g�\�dے�2˒����h�����W�ױ�� ��*��i��+:��� ��)N�K�h��0i�  81��Ғ�E�亱d�%G��LT�N҂�v��9�o��I=�Ӥ���2{^�b�r�>�B+c����.V�3kf�	��c���^��`���~�)gߛ���|v�9���ێ�|��~}���P96g.���6������� y-wJ���%���v��1X���vK��e�V��#Y-d�5 ��7�C<Z�,�1�����PTLL�6��c�w��dT�� m7Mz8�N�3>�N�d��^����o�$m1�8c�i����7(g����
���2����>�X��N�7��>�e&���8��4��ݧ��x0�B�n�N��r'���g+x�᷏����OۉX)K�T>El�5�!��`B��;}*�b-"���|޸x���L}��mP3��?t)w�2��t0��]���K	B S-#ӐH������٘9�	B�����H2y���Ď-��'�[/PA�lH�D�� |]�m�U)k�<���JY�t����`L�r5���^&y'���>��Ng=A3Ԝ��a�����R�*S1��������Ϣ����i��+x�7O�̺փ�I""���ʱ�d�����`}�;�3^��]��d�"�}w]	���Kg�G�b�:�����z�O�i�������=��4�]h�1����\�Yq��N���v��l�6;�2�,�r�9J�!���`�e�Œ��I7�w��>j�;�Wvp�ò�q���5}�Us�*F@�je��G���
��1��C�;"3c�y+CY���;�h����+;��#�$��q�|ɲ���{\��ZQl�v�������B�K�s
��T%Ŝ��d>�a�y�
��gF:�L5�<WzLs��U�1K]�UM�c�W��U��[��2��/���m����A��>���޳��%�Rwf@���J8��.�1d8��!���!����"�:#�e���>]�%�9`��Q���2Y��S`ss�4���6o+�����a�u�u����:#�F.�ٞᚬ�p�G_�������
�/ў��ihVZ�$Ǧ�/�Χ[E,�_��N����?.��n���
hu�_����~�e���r0!���Du�Z.��/���I"f5�"{��g��F�����&o3��F��,~z�6��p�$rې�u��R�E�]7��/����#IbG����q�ƥcr��	�k������y�To�����B�|�E����	l"�y<;�:`֎���P)[,�`	gaꐽMPmmϑݑo����`G.�'�B�'�:�
���Eϣ�"Y�C��o2�	*A��;Y`N@�5�8�lH���k�m�s���*��<*�\��|<�,(��Y���1 EOf�F�y4:�̗`��n~H��H�T%�G!�;c�~���z��f��3Zy�:���m��~{�p\�N���T
4Ь����Ve)��G֒&��xR�ަ��w��ۥ���<X��|� sA�p�b\�����r��i�~�\\CI��]j�}<$�E�F��O䋳�!�~'Ð�mj�_�R�uɸ�/�t��R]gy~����.�N��#A���
K&�CG��^��[�@���߾~�����l��3�r��z[~X�)�">+nM��s�f��_�"�uzS0�W�b�����������"-��Lܴ�Ե�[+�k�"3�;3�>T;��Uu-�JB��d��|�L"FN����W�>�5�+8����r�6�dav�=z�oD�&��?���0�����P���q��v�TF���RF��5���=Uc�VNo��+jL�z_k)�5���Oʪۻ����$��@}�t~�㤑��@u��e���e,U;�
dBR4�� �4�b˫��7���H���#T��	Js�H�~�-҆k��C#�mch�a����5�L�6�O��c���Ġ�壺S��@|e1������2�®lb�S�/���� �ᨄJ,�����s�VP����D��_�a8:Ҋ>�ׅ3L�}3|����sr2�|`�k��g@�mb�Q��'��u��J�Ay��#. �S�����Ft���������>�Y	N�e's�[�hLKKB�Tz�X��7A<�~��g�,�$`��5)����c��c�>5ľr��n�%�SA;�&���4�zh�Y��V��q��i.N?=|G~	 8"��u�"`�J�(wf��I�fM���p'��ƌ2�Y<_|���x5V����l4ɥʕ�j3i��I���uԧ��6�@E>���ˮ8���^��b�G�I��I�C�+��#�t�̷ݟ���-� �|�'�W�r5��,�{�R���H��R'˦�^+���H�������ޙTQ���E: tޥ����B$�������ӟf� U�.�����:^!��p�>E��iKA��X�G�<�L�C?��F�Il \e�d�������aSxa_�x�8���sG�v��
V��~i�!2!]��lr�85���'���f||y����ᶁ䡯N7��7��O�{@t�˫��5�ܻob+�y��"U���hpBR������C��\Nt��D��ֳ�H�4[Ɵu91�1��Oޢ��Le���5�c����Rd moN�^�9}�4f�ѹ�*�4�(���YRa������*���b�i��5��X�Ş�;�>9[%��,~d������)m ��W�8�O%�ή��>��:ݚ{d�$���?�e�K�%��,�,w�Qb�N�]�P��z���6�m�K^��[s���c�]�{a�j�������u$��	YH*�Y����S V{�i��~�1Ȃ�>��bt]v���a6d sUX4#��t[4�N�âO�eC�{VVIR^̸,S��EWngq*z���g7�[���F����e�{{�	)Xam�V�05�	b�F�Ȼ�î�8Z���+\���<�P�]$�U9s���p`7j*�"3�o����"CV��bo�I���xz����f�T�hW��E�aR8<�d�9c(�lg�J2	 ��Vʭ�bd�i8L����͖��o#�E��'`�-p�s<oI�]$8ڐ�6w�|A�/cy��
o�M��� k��n�Kr��8�� [�����4]�	��\v�����IWd6
6�h�'�-���1�r�����>[�
�L��ȶ�B<?K�8Ś�펔g��j�,���"�ʹ?�)\��S
�j�֑�C��'�f$����"Zm��Z��s��U��q)F�����J�r;-��!
X&{ۖ�=��|�۟}
T�s/8���'�k͎�6��Af� M;�	$A�+9�6��2��J�����d��%���9�qX���Ć27n�Ę�;\��K4�(F�&Wo���Чi)��2�KA��-n���{J�>��;O�F��a]Zz�0\�V���|�+��52=ߞÈ	Z,�K>#���A�`��]��@�"h�p�s#L�~�J�@�A4N�&�9�f��iͽ7�[���a�Π��r4$�� �R?��$��_�.����q�m�@�:@hv��r�Y6w\"�I<���'L��pCf_)L��G�'�V
��Ck��wL�sjews��t���+�_H9|� �?�K����E�}ɮ>���| I��}�g���p�yl-F�{���u�D�pvW�j�����ӯ/���,�MAd�j����;�R���cf��)���l��7��TB��hƫ֣0Z4��J$��"�����K�A骝����i�>7�㸆�mAy�V�8��I�s}��~�L�V�3�ƂF2��FU��"�c��Bkp�-0�:miRSt�bD�ʠAX�cU��İ��%7�$j�oR�	���#uN��-��UҤjic�C�-r�����1kϾ��az��ey"���XDX=]�K�����ۑ��MO��'�|��7��#v����Me�Qn/E����R	���(Kh��O����hH[���jyN�(@�=��hq���}�l��[#1e�<'��@���I�d����F�%����)v�W&�
_�/�w�(�G�y#��NyG*-�^!f�|`���>@���d(%�Y"Y;c�L��Z� �^�HyT�߬�βѷ`���Ñ� �tF��'�b3L��7�����Y�e�:�Z�{��b�̩ͱ,���N`��U,����O\�^��i�
#���0̤�[�o�o��:JGBA�ܤ~�1���%�Vt��S9D�rA�����S�}��}UV��1��3J�'��Ҏ�J�I�G�l�k���v�hF=@�i�wא>�u.��%��˂N�;�6�[�8��ٳ��r�Y���|���	g��si��j�b:XE(@w�Z2������GCf����ke���2��=m�)'>3��A�)�\No+Гy��8t�aS�
���4}��D?Ck��惝����)U��N'!"�,��5�Y���l#kS��2Rq�8+X&E�@���yV�z�����qk�X������$K����!�
4���J�ֳ�_���V*�b�8� �A
`v �kƑ1�V�Z��;���z[�H����Y�
�!ߕ;��]��DZ�^�6	�,97�G���Q+P)j��@e��ؼ �[��[u� �Ot��ڳ�)���JvA��)��X}������e�+�3�"��c����$�@^?#���3d���UpJ�96]��h��%0Ґ���pS�
_�4:����<� B����ܥ��[�4��o v�f"U$�Qڳ]�ɫ�e�X]�<o�>��tG%���1Ó	�M�����L��3sƈ����t22)�HG��w�u��b��$+!R&ܐg�u�E#�.	�`�O�zBo�-P�U�������ڢ8AZBsC���<�G�3w{v�hxq�]���Ш��Bi����"�/�ܰ�"�qt~��J݆R�fL�����q�A� obJ�J���of��\�B���M8�1���	����\UB������������D�����l���ZU
�ϊ�d� a�P�V��QK{���|�Zki;u��W����
7�B�w#�̵q�P�����Q�dJ����ޔ�rH�CS�B�� �=*'�<�*�dĬ��`ސ�p�+`֓iQ(��S���B��5&\�d���Y��vA�it|Z��f&��RCJ�xo�d�Ã��2w��B�N��&,}0R���)���q�XԭAi}v%c_�V ��X��_ !�!5 ����Ѽvq��1{�/?YdW-�18<`^+����N�WCA����HcEC�5��h�+��e�Q��}���OnL�0�m3�6�+��+a:ሉ��%���1���5^L���6O$Dį��L� -!5��玌����i� � ��Q�w��c�O��_������#�����Rs�_�5�[A5�?��z���'>�1���Ϛ<��9�1LT�"���H� U��Xن��3���|k?��P�)�r��]�5�1���=L�Q�B�$Y"v7�$6&�=���NphZ�L�d�J�pB��+��	�%�/!x�dL��r�* ��zY`�~+ ����(z�����2"��s"�P�}�Hd�K�Y�K����$����F�w}pꃲ�c����&:N��F}>{���o�C�G�|���Z��̀�l
-c�󮊬P[�<�y�δ��GF�4��à�QM�@�/SLwSj��F���V��91PXi�H��:�����0_)*�׀�(d��$�W�N筩��d H
@� BbL�enW������n.�+4S��(�@s98L���b�$�xW��v���6��}�:Ɉ��
��١m�Ӂ��p�6��\>������i��^'[5�M��w�yASo��V��;~����Zrf7����@��Fy������V
(���T��8l���K�-����Ͻ�б|�����O@k��MT�v�HЌ�!M��qEI���	b
9�}��ڴՍȘ��&�����y�`-E���g` �,RAm���Th�&��*+ODF2��Q�,��"XN+5m�U��
P(XU�bV�[�V���n7�r����#��[/�2k���o�T����γ>�ч7{x���h�!�#�9k��~�n�R��NpƢz��Z�w3Z���c�穂]Q�'[�_�dLaШ��dU�E<��a<�GH�)���6
uG�.3���2�T��b�Q01'�O��)
��X�����=�5
�!����2RT'``�´K����n��0������7���az­�(;��`[����y��0��,�K��VG���,�{��ܨ̄۳��7�&;	�n�>_�6����a�k�2��m�������Ĵ�{)�=$���T�}�}�����*@�@�����$��P@��(9���*|	�S0���1H�{樧�,+X�=4Đ[��c�/��1��=��b��Ž�!�]MZ�'�
ӳk��UA/��	'�$~ؒ�ә�=�"t|FU�_�xy� ^�G2	G���G�7�X�>��T���u|Ga�3��z��2bo��,*�g�{���	L�?�"�W�P������j���o��d����E�i�j6�f������=��'�i���@�U0��;��h�\5Ͷ; J��E<3C��{�d������:#3A㚏�yk?Y��c�0��/�o$����O��0Ġ �������Ȱ�R	�1�Q°3���kd|兪�J�|��5@�O��!c%��%�Ew��S�I.W�\���M6�j����z���w��9g���0�����'�{��x�q���[�H9v�����$́�c�����T`����=�O��T�:�~�,�
:� |�[/$= Ե��*a8�� ?��Z�\ЎW)6vf�À$05��Gv��u�� >m�D���Ip�Y��t��Zyĝ�>�����~��[Y�V?W4�㷫]�F��rJ�d�^�$8����?{��#����r|n��7�J;���~5��A=!ݹ��@�I�lU���	�"��HX��ٺbe�P�2olB�gWd��)�/�g��RE@h?'������;`��O%{��3��dM�􆟈�m�R������g��Iv�4�K�y z�8��=
m6�V�E���W�5׵e׃?L�t9�B���ul��5��LX):����eư�~�8Vw`*X����eG���ޡkU0,�k�@���,�����/���c'MK �R�{��Y��h��ɧh��)��:������rq��=�������4i�|�B�_�ԝ��|�����A�UPBgP{�C�P<�P�FBQh��:�}�Ӣg�'��+���������;!$<F���������_�Y���w��G��ơ ��DE{��Q����+`��YR>_B���?Xդך����w؂1{��N��6�O �t>
���X�\��,�Fjĉ4T�����e��3!���No�Z���EӈW4��n�T�-Pʞوy|I+��:I����ge�lO3tm��:���������\>:�3�ck�Ӑ�����C�+s���ԇ�L׳��,����%ph�$8��ღ�JG��J=Xn�1em�d�I��э�X�g��ћ^��Y�颥�o�s���}3��l�'��١0�)�k���vv�b6�~�a��ܶ�;������q�s���c��_���#G��c���P�FlӥD�l��n&�t�j5�7�`��<c�l������{	։�C�N;�P�iO|�u�f�-rO�O$R�>!<�����t���B��>H?��h�� f{�6~
͘ɦ��!������K,]�x�n15)�
`��� Nϛ��'\ �pv�U��V��B�/ɩ�~�"T����~����6Ǫ�zĽV�`��A0Z	���x���DF-I�|b'�4Y)Sܼjy�Z�/���E�Fq�Fq%_������z9���p�����Y6c+�~�>�y�%V�J�0i-
㾢�`O��HL6��f4��K�KǃZ8�y��F���v������8���?���$؉�e=���X��}���r�#�	Nx����p!~�1�gL��bĦɀ���%�M�q�XCl�
_,��Vqy��a��0lz�pK*�/	]D�b{��M$²=���,,�������,����һ�:�#�l��VC0�յM ���N�u/��=��l`��3<�v\�7�1��2���PT�93Y�w��˾49� �Z�Ӆ���}IfWB�z���kE?U���-G<��W�J�"g~׵�T;|��T?F�!�/�D��6�y)e�z��<�#iO��C�'�&x��ͥ�.��1݁�ܨ�u�jh���;�ɀ!-@+��u]'�s�|�[c�'�(��g�|��qXY�S�_�PnN}%�s6�5"�� ��~��O����C�=P��8A�#a�hޞ-���_6	�w�}J�k��LWrX�?C p-&��m���;�C�{�>��ov�\�pw���2n�P*��z�b�	x?�y��,���򂓬|�p�O[��ʷ���1+��4`R�7{��U(>I!h�)5�cf)�zA��a4/(P����09]�����gٕ�:�W�uל�q7�6�kH����鎀I�L�_y��#`�h�&���#�r}�<���;��Q-Wd�i��Kn���|���ELD��IgE|y���w�-�t��O5*�Ad�@"UK���m�ұ/ʱ>�2����Ǣ�<�O���ܯ16O�����.�%�Ʌ=�4i��CF�����:9u�4m|͊]��9w�V�̩����X2�j#D�Yπ
;��P�9�pZ���F[	C�'�6�n��d�b9�&i��aǛ�(͟�J~J �e4Nc4������y��C��=Z��#`�S\�N(Q�?լY��5��@ƏE+���OhO���y��1�����;�lPL�E-Z*�-R@�*M2&߉
�h�L�[�;��ݒD��h=�� P�����SK ���1�8�E֜"7H~J�+rd��s��$&�G���cm��ҖA���1��^��uC`i���X+Z^�ۢ��m`Kt@���n��t��Y"(���pu׉�J _\��F�g��'�M�27v�]6�i����'�����KBH�Y ��>��y�\�}���]UBo�E�7#4�eS�W�2�Ecנ�K����N3s�w���d��s9��^�W�"�Hk�"K��wqմ���Uh���ҹ̚����gщެ�?���6�2f��J|8��!���JS��V���n�'��Ɓ��g�lOOl��?`(�k�8R�M|&��TX��%q�E�oNS����y���6�S5���G��uX���͋�T�^��}��g��S�H+��^�������s�i��1������OI[ۙ7��X£�N
�����[
R}ë�'���;�uE���q��$�rb����%�"��yE�`ҋI�fA0n�&��o�6Ⱥ�q��l�?T��͌��dE���$)�����q�Z������<}�s�q���,��U�$f��b�n|'����m�����J��|jC������g�_$���|,�At"'.��@�\��T\�YiGLp�v8d�!�Μ��B܅��Mi�zH�f(�Ґj�F*�����HZ/�/-|X�iQD��Zg�n8��i���-�.���>ܢ�V&���op�.n�MDƂ���%țٕ�ʛ�ۛU&�Qym�º��o/
��H���aLW�H$F�p~G)�k4��B_�p$"V��F�
��&�F}ϐ�BL�O 0M��%"�9i��6�|�Ő2��y���?̮?z�U�e�(�SG���2�8)8�/Y^^S��O^R�%+*yy,�������C��r��`��rhD.ܳm
^��@���)�H�쫵���q*Ň�}�&�e(��iĉ0�5=iC��d�Ҭ��,%�$�M�2����`�Kj�u���ª���W�`��{����V��?�
����K^<�;��[A������A�@�v��*B�~?4���j��b�ԟ��2�^cx�1�r��zغq�6o=[�6Wuz�F���4��D,!�q8ž��
N1tC�\�w�sp��j���ϱ4�@����G^���"ZP :��ϸ����&��}�x�paW-�M>���=�����O�J~Q�.�މܯ���@1ʎ%�E�y�Cy9��w��_��˫ۻ�d�+b�O��Lcu�[���Rk�5�OP���ߩ�6u���roe��>r�]�E\S�.�|�78�i�C��ꁝ,w#װJ}�*��C��K��D=44����+,�rZ�?ߌ��?���Z���Ê(#���u���!�Z���
~xF[Ԙ}���(��Fd<�X�3��e�-�T�K�q}>s�Z8�5%[�	��[|��+��O/2��R?^ U�ԡX��R(Q��Ef����5�_S��bN��.0�8ԏ�����cE�/��-x���UHə���J(�����?<T-H�Qm���tr$6uxmWa��Yه��H�gTRRYw�)O�"�h�����ĵ���k�����I��Y�ȍ��k
�5��l}���-PtA��4Ukn��F�D�	!i>�z�B���$X�'�q�5�ꡎwHm1R!I�&�{\�+}���� @��}�7��jTd���mu�m�t> \��D�dITΙm�Wl�@%����r��!w��#��}eǍ��<��>�TZ�c�'D�6+��SO�U/N�*�27�����ӳ�1\2�����Z�Ɨ�f��*/���� h���2��d�0)	�⵼cw�<bV�?>?�Eh��lS����I�U�'�ޛ�U�B~�B��;e����
wCJ�"��/Mu6kKG�=�r�ӽD
�K0ܵU#@�6;�g|�U���7~�(>�=���x�M�Yͧ�m��"�>vr�|D����lŪ�/�Z.��*��A<kD�CP�?d�}�D,�m����Q�o�Ě,�Z��[��	���X���?GI�k4d�:��}ٲ/��6��ޠ½�R�Q3�5�?-<`���c�M,�[������1���%�o �6/8�z8�S�n���F�P˛'4&�J*5���i���S���ѫ�3\e��y��`b�퇐�>�Щ���a8箤��v�.�Mn'��A��)���.XS�TV�i�
��mpeo������q'Q�O8}j���E���,���nܮ��=��c�lZ���[U&KZ��{�Ì�6L�8�����cY5j��������24%l���k��&�xjHl&{v;ٛE�ue	���]�U�bӨ^~D!���4��%�E&��?�����6Y�ge�%��w1��r�#�ĳ�8s��d�~o����A	h'����>LǢ/�dۣ�HNXMbrz�O�Y:fu�֦nhS>�h����P$<Rm}��O��:CX;ZL�W!���M���k,��:Jk��iL����m����#.E�o?�^}t��~����Sh�$�b}H��s�Pk��M��$�SL��k�}�VфA�\��a��iѼ��6ch�=8NXj��f��A�Iz�r���(���ߔ.	V�)ɣ�zOXQ�j�"f`Lz���qm���6hXj|�����?w�Um�����ʩ3@���Յ!A 0���foN���	䥪��p�pxX�R닂�����0A��Y��j���0:���y�9U0�`<w���I,��ĕf����Z�(��N�ߓR���h�jޅ��
��2��19�~���]����t-h� �v<	K�U�͕����RwzM�~�G��Jp �Ƈo�/�I��D�5� �����z�b�~��-^�_Y5���f:H��<ɼ^x��H�J�^6��"_��� ��y5��n�ш-[^���`<��9O�wd�$�^�L�D���E��qf/����ͥ	c���������do)捘L��W��`'�/ɝ����ϣ�h�aP�L�����1���c�-��lA�����{GpD��;�EK�hL$�S"F��#����q��ؓ��=Jp�������QeдZ%zXI4%򑇶�����$I�pj+]([�����L��ĝ���Oy����I�Uq�2�&c����H
����S�bf & #:�ڎuu;.��s�Y�L)m��@��Z��k�$��m���tB�_�E_��N���Y�X�G��7A�S߫�*쯫�x�'�f�H�	�.�VW����_r��>��bg��IK��5G#��0����с4r ��N?F���[ȋ�/S�e���S �⮌���d�aW��"l^�_21�����gJ�'�q�5qv�
�Q'�!X�����f`*��%a��9\#�/в 	�UAŒj���DJ`�E����{$Ph�=�v𴡢�����\���E���2u��z�f:K�L��SJ�n�m�q�Z��k:>W_C���u��Hk�*�K�/�՚�����rx.90C�W�������WCT��Z�1��B��j�2@�V��d;$�7��	�w��H�o���}}�d�uW�JV#�Í��'�����p��L���?*���G-o���;�tX\�wY�ȟ�~�'��r%K��Y7�̭ʑ�v7F*��Q�Y�i��1�1� PK髒��]SI�#�����`	xX��A�Iǔ���;��mhd�J�Wb���]6��՛����n.rш8�+�=35�Hb����$,Q���C���Ov�D���e���/V$q�?!1�p�T'>g`Ɗ<x��r��N�&� ���<\�]/��t��~��<J�C2�>�hR�x4yNW)�A��@d̂����&b��M�� VHh��U�0�:��曱���Ӯ
��O@�D�AU�Jl�u �S���+z b�0������-��ރx:.g�>.Vkd��Q�>ix�g����1x
���q)%����[�/꺒�kCV!��Lb��͏��)o+��o�Kk�3�~��i�#��}IR�.�?�8��8l碪�	�����G�晿*�2�U���BO/�c�5��C+�� &y����qa �kP�Al�guGJU��aT���ْVuBt�-��ّ�NH(���0�(�<쨂\ՖG�W���U����I�aٛYg��Š�DmI�)sh��kԫ��(t�6�@���MKWi�>�^���Ѝ4�?�v�a��G�t׏�Oh|I�u)�����9\<���3�o@Z��`�p�1���4�ꤑ��^s��RY���)6p��`M��iP�+ؗT�.�
���"��m�Ujt�j�M�S�'�
��~���7�	D��~N!@�29� ���u �����>� �H��/2���k��k�n�8|���͢P0����|&�q-�Z���Y`��V�a8E-�J^�LݿIH��G��;�f������ul~����y�e�_��ORk&�+jK�<��<�-ʹ�^��jH:6h�=uZ3Q�@���U��R0��i&O��v"����qQ���1��Z���L���I�L�� �h���������M��ϰZX����:��F��S,>�8� Y��$��o�������eKl�7�7�/�����3 5Ic���.�_P��u%���aW��4� \��KfӘ/��ʥ��4m�h��`�����7^l5tA�t��yϙF(���'f��1�B���KWI��|���2�#����&�ԅ�{�ۏ���rOic�Gy�I�:��f�CFEM%*'/}*B��� ��R"?�p�r�ǍdT���������&U����Pb�r'����Z,ΠӪ�
y�����&&yO�|�L+0 ~=�j�|j&�����g��Z{iC`KYIߓL�m+�u���OO�bUMY�H7�"HyS�c�@�  ;�6��n�@Iu����� �L,�X���aSK�or�_�!�Y�#��n����r�y�%+M��3��P�K�trT*�r^�F�J'���W��_�+oh{�����3~�c���	�=d�F�r��y8�>]�~��|��,{�]Y^XN�������e��ꎑ ���Ֆ'����# A˰4"�������#���$�ϓ��z�K�kLy���AVh�8�j!�y�Gf[Q��]�3�~>�J���>��شJ�7����8U�*���2�7��e"�;��B��2Hu���\21m�:�t�:��v���� E|�FR9ש@f����-�0���ך<1Pir�*6��~��\��Q�+�g���?<�v��̄������-��(�2�A�1-!�QŌ�>�T�-.�5
ܮ���wʁ|a�� 	�f	�Ͻ@��	Smr<�G�KG'G�S�<�#����D�bK
f ��'Ȃg٣O)��N�V��<$����sK�ګl�߽�v����r@�|��UCbN��Wa��b�!�>kr��ޏX�ɇ��G7���s%R-�gBL؟����աѨP/�-tY�Z8��a�[q�7��?}1q�z?�vȜ�+H'aK�\�fP��\��N��~����
�4��w-13���d�aKbC��4��A�q5v���}A�/ݮĺ�C��� �@c��B�52��h��Z�/��nC^,Q $��/v0(j�*��Z͟Jyp;J��?U�<c&��
 �_i��Yz�\'�:����LF���g�rW>���/|e�r� Ќ��:h������e�k����?ّ����CJ��M�Q621KF���0h�7U>Se�w�/lr��>��L]�A�n]cI�hp�m�Na:��/�P�I0�Z�䷦l��������{����~�H���&W�1�[�BJ�.F��7\`��Hכ�@Mm �x�^V���(����� !���욗{�FśK�� d�h��~��5@������}M�<��IV��O>��YF��Q����8�V�S#-Z�$=��E���Ye�EP�Jx��C�$}�yɺ����86���Q��<A�H��>['(R�|"K `��,o��䕃��4G��U�Y$�c� �Y�kY�arK��,��4�򃵊1R��c��ӅGg�������&jU�{���˻B^%.�{��!_�zgL�]z�ͱ��5 #��<4 m*Q,�m/��!+W���s�9�b�Gj�-�.|I�ly#�LN(0!lD���G��>�K���'�:�O�e3���� ^���,��L�Ԑ�T˴!�zG�Gd���G�F9�FyG��2�]�x���J��-Ev~c���-`D����'(�d���ctOa�r��/�-�D�7�^WZxstHu���7$}�ƇKH�j�Y�+��B���~Ќz��*�4��k�}JO�6�
����ݯ�]�4$��G�!��L���ث���b8ff������D��@����EȡJ{� rh_p��dO��P�r��@���?97S�p�`
7�w�A�D�U�v���\F#���?E�gr'�v�!;�b�r�3��1N^���t�t}���������&8�^v�j�'��oڪ��gT��j��s0��*}��@��"A��O9%?�w�]�&��O�%w�b��%�۝�_�ɒ�3:Cʖ)K1�Y�!Yk�w+��-	�;��o~ݍ �K|���$��eL�ҏ8��ͨP0�E��	�s��>��"�9�s��؎�	'48���݁��G���C'�H���px�¾�S��*�e��J�k#ǧ��o���,멡Jy�E�����(gD�p"�����=�٫i��{+vN����u��ֿqw<���{~q��.�&�?R�^o ���L|����/Q�lu`y�����^�-��2���8�`Q\�D2���eY���o����Iؽd�>f��	����s>5p�!+pۿDb������o���Nv'3J�:D�2n�]�vV�ꥵ�\Sv��-yP���%���[ꥄ�Aޙ7���zA���C�<
:��0�.�K�?;�/�uY{�ٞ�i�z4f���Ubo�	�_�URy0�ڠ)I�a�φ�ܥ1��?�3��{�Ҿ���˄Lf:Mߥ&5����T;�9�-"Y�gY���s�6 ��ή�Jd�:����`:�R��du{��8|�[�
�(�ٰ@�oM�Yǁ�4�a��+��g#��O�v�
����F�A�!5��H���*����"$B��sqT�l_��[c���4��IB0�Czv^��i	'&-䰻�� �5�S�:���z���-R��\Q�G�L|�����B�']m�CM��]�#�!�u�>���]x���K�r6/�h���K�Ǻ�$��<{���&����ݢ�Z _���!E�V�(tz�^B������gtr��B::�T+�;\y-	U��!���|��/��R����f�֮`�#�<J�W�]n��X���R��g=A��=�?B� r!��o�|8d/���Z.A�T~U
�<���_+�MK��2����؎�!�m+�v�O��iwr�ӕ���e�p�<�qo���ۼ�a̚���GHu-��=퓠!��k\���z�`�)��Z���I���zUg/�.yjm�h{���nZDȾ�A�s��!C�X'��D��գ�߫F�$��0���aS:�p�@X*���
	kcCgU8Ʀӌ�xB�ڨ�"�9�n
)��,7�8Hb��S*�V�>��>>�+>+��)���t��,X����xj3ƌ�K4'���,��ðX��PW���n b��@� -{��X}�#������ki*m��I��K�K��n,�+n6�Zc+}-�y�:U�h�bѽ����cl+�s�ʌlq����0܃;�t�����&嗞��.QbH�����;���G��Ӥ��̰ͦ�(H�%�0�	���*X{n���H�F��Η'P(	���̕ߺ#e�p{�X2W��
������D�����r}Sj]$���� ��j�MAy_q�_Z�=�Q�M	t!��BQ�BB��btߨ�A��ψv��d �
�]�ӟ�Ɏ���~��Έ�'ZO�RV+%�,�=��d����'�J������QuT�@V��u�v����T'�M��WL&ȂI��l�1\�`�=/�����^Ս�f�V��ꡳ�Q=�U��?���%_��Yj�f�"C`�!�Χ�!ō��D�Bn�u^���ZS�p�am���WI�NC��Wj� DoEbG�4���r�d������y�;T���{������������~n��8<�|T��1�}Ơ-���o�A�bK�? �,��g��Vmg�͵i���ΕM��gf` Wh������s�d�<������~��a��#���i�����2J)p\���������@>J��M��	Q�9���ʷ692C��W��m� *z��C�4�w��# p˗�RmP��C�S���_��\c%}Ce<Ū����5�JkSf<}٫���1�Iyng��%Ϫ�7��nZ��.���D�F���Dr�x��b�8>�*
I��Nv��BZ�7����J[r�?,�N���c�D����H�v�!�[s�ۨ���;�y��C||҄�g�Q��I�,Ў�f6yWrIbp��'����A{o)/�!���E�_Bq�[_�#HJո��R!�eIN�[�R����ҽ��+� �(Oy
O���\/Q��z�Re�,F�>��_Z/�v]W�	�{hq?��ȕ��� �?�j̕e��]ҝد�5B�\�ۼm���J{{�;c?�l'��A0��/�K�"��ND �.>��w!��=���y�a��o����אN�G2���;�,�C�����9�˷U�^siT_�2��̬-��:�b�X�Uh	;T��KN����xZjR��=C����(IA�/�M�>PG��s��mwޚ��#���C��by�G�@L�OX!j��s7b߼�G�m�R�x�z��F��e�J�g�?:!�������&g��x���U8�]�E���ݖ0�:�������$~��_��e�	'�j��H�s��w��cp��\j�1/�T	���� =��~l��I�7��L0��B�mpn5C��H;��IS�]2�'��@�Εp�};�w�gT�BH[vt5L�)����A���Z	g�rң��,�N�B6E� ������Y������J�
��?�@Le�@1��K�3��"ߕ��Td���%�՛�Rl]Z�}�`b7��*���O2���w���6h��b;�T|s;����T�����6�Ԭ�ov�W>��-�hJږ��!���3N$rrn����j(@r<���U��M((�W�%^]v��ﻂ��U,����n�X����ߏ�J�ft�ي�-�c+����9�̰atCȥ�)=R��=&%`�	^�#���A��f�D��+]E����͵�.��&�7U��.�AgD�K�"�~���msx\��q	��a��̓�A=�����|<�u;1uA�	2J��w����!�W�R��^Ll�~�͛�ު�*��KY�U|K����V�X�We�*���ϲ�7���&赑Īu��#��W ��`��\U�$_�}��4R�H(�E�[�������s��v��qg���K5���UT"�DV|j��t=ă0]�Y�`�$T��[�d���ŕn����t�gD�M�J�;�����7�����Z#�J0m%��(�^����&$�H{Q��bb�X��� Q"^bTÞl���������LI��$��\ȯ�&�z��4�����qtc�|)��^�_��I���['$�1()�<�[�X^�A�����yvQ�Ti������l�d @T�s�tc����Ũ{'�N�zw��p �+����-����smu���=��,0>�w��:�ښٗ���-�Y�2��,���w����A�9�!^���no��J�zrGӃc�� �M���,Zmy�ر[Hئ��V�I6� �O5{�>��~F^�'�6䎁ńl�$�@�0����iZg�S�o��; F���x����	��,Q-��Ƅ��y��h�Gz]y��G�o'N�,-�����/OaO/U�迗92�i$��l����xD�.&�Cə������
t������냲8�E��|�%Tz�U�t��'tx茔}�Tѕ�SՈN���U���/I������/�kq�(�e�Vd�ŮE)�����f��V�[0������;c�c�J6(��\���f���7�yw��d��N����\� |v*Gr����&^y�\x���*����xg����K�e�ܞo6��00��N,�2�es�:�ڔ��M�B�N'4XU�nz�j�_�^ )��2�{��6�7�wwQ�@��!>�y���֓��k&��>'�Eh���H�Il,@.�?{
Z���'�3�T�L��SHD�x)U<��i48��gK��n��FE�JA���2��I�����F3��R���b���x���&�^����O�@�`@������@��ɯ؝�-8�G1!5lᥕ~���T�l��Ɵp6�<e�D��y��M�>�_����:~Z�"I�3�*�H@-k�ß��e؀��mn�$�1\4E��9X���n�῿7�'��|��6��x�3��T�ky�`]���Y���d�`��9��(�}sT�������CwJ�Vr�.��&�_9;4�N� PϘ~�n@,o�P_�3�P&�5�Cɪ��Lz�Қ�a��p��>]�ѭI09Dd�󪶠:�F�b�}*�d���yL�5�ƜO#�[S�f�D�\� F�`����ȿ�6V_m�mҦl����"Y�W�fvԟM+"�ǈZ����Q���b��+�%-�Ɂ��$���� ׫���u�y}B��!��#�=$�w������e�j2݁��d����V��L�c��0�L�=����~i�P�p�	����	K��~�g�a)��U�R�,dkv��gJN>q��XP�h}�@	F_*����Jj��h+���x�7l�uu7��)�Mö.���J��v��E>�΁�Au��<*���n��2�w��,��(�v��J�w,�JF� 31Jtv>�㍿�a�~7��πR.i�Rv����٢�`��E�Mi)�"Ѕ�LC�4mOt2��\ƞP��uT ��P�og����I9V�d���N����h��Gͯ'�bBO���y�.)	,ޣC�/��S��za6~z�5���jx�QP;�����)*��Ϙ	����������.B�"t�46�9[�3C���|�x�+���9C��3��\��\���
���9=_���������hj�I��ܦV]y�@��2lZA�i
��������	�o1ZG�P�d�"��駦h�N�ӳ(EH�E��OI�ā��)
��������!������\P�wuꤍ�G�=�w��l?���*o�Ba [�������m�=& E�h,�7� NЉS�-�DKuN����u#\ի���_A�-�}yxZ��yd�[c�ű�>v�g"��#r�y�Qke��[B�8d�����7+�G�n��6����/lQ�1j�$p6����H���n<�K�@��Ͳ�[�vpL��6�im~��;↉N�X�C1���0@�:� �H`Xh�m��<κOL-���[A�#����eX��~�s_��7#�˃��N��V0|S��E�V���a�j�\�3�O�_����`�ձ^cG��>�Ͼ9�n�i^D�B�a<j������Jh��>J��2X�o�JPV{%QP�V�5
�U*"vt��%:%{ʘv'���� 4J���̗3���[�k��y֨��Ui�^'�i���VB���3�0��X�L���!6&a�/�r��cȟ�$L%���e�F���FH��$	ˀ�s�Jx C#�V��F3c�7m�3�YX����K��6��ʙ`��B�2Gx��@' �T�C$�a�3*�=����
�U(�S�s��l+�8�(�.V�oF�~]��zJ�{@I�6{��+-j���:y2
���1���7��B��4��U{�)�Ȭ@]�N�P�6�O���c+��%��̶��f����ŻFy�
1Ae�O.C�k*	��ѝ9��'� ��:�#�N|����>�V�N>ߤx&�A8_^� �{fX��7^3
�('�(�wB˻�5} ���2P�z;]���]F4T7H���q1�WM�g!K8��~��.%�(�':׈�7�Ʌ=�c��;&��n��z������m6���� S����t'7�S:=�Gsf~�f�ﾎl���������p�;幞uF���j�i>�����uU�]�_�4��zBPMSqw �h�w@�̇%���酚��^�1W�����X���[�Թ+�2��AכM�(�=>��'�&՗<5��&�qFEB"J��LU@兗��XG3W��]�H#F�p���+vr&?�u�*�'X�!&|�xXK-g�`�G�
�!O"�V� �q��4j��9�߇}P�o��`��▎����>�T�_���>�w(���Z�M�I�c��qS}
�a�p� �w������
b�QS;��^i2\qƥ�D��!�{8j������=�r����ǖ֎2d ���i��,+�!ہ�e�M~���Ņ��|��أ�"�`"���F�h^d=�����i#j�.g߫��SỏOQ�H�� ����j�N}ʳ�EJ<��m�p�a;��k0��CD��\��a�0H�����F&�0��vPG�<φ�=80�1+N&�oTErP���U\���*Y}���}�n\�<���sn�kSD.���}��ſ<+T�����w^�$�N��IƉ�T�ӈ]�����(�z� ?��&�}�[!]trb��wk'�1�V���kO�b[KK-��t�롬Y?�W��y`W���T��e/��[(�g�7��}k���5��K�OŊ�Jx�|b8��a^5�6��z.���3��v��ҷ/{U�/�~w��*��P�~<�*~}�RY�)Vw��OU?e������|�|�����W�U��8��}�'��"a�����/9��M���y���+]&��?�ܯch����2��	ٻ���H��}|�����׉rdDu#H؏��C�M&��u�&r�ft��8Ʒ#���
2Xl�	��5��2�GM��N����fЃ��o�un|��"��e1���~����u��J����,�	�'�a)��SJU�4<I�����JGi�Z�s��	�" �"�@*��#�x�p|��i9-v�i���RS3���E�AC��#�bx�+��\.S�����JnQ�mυ�� �<�>����;����r��f���|�DDԾ�Nd�����S���.=<x�+���'+�G�֑J�A�:�Kի	�Z�H�6��L�~���;?�ؐ
�}*��E2��\��M-.3�����`��C����_qg��`ި-ztt��DG����e�HeiN�d&c�d��|��E-^��m'��p�SZ$n�~'Ҥ҃�da�/S���M0��a�:c篇S�Ḿi���ǳ��8��轴�'B&�\��LT���(8,�FL@W}�7!�Ιq_hz؞+���n�I��!��<�dr��l��mNV�~�k��w|guCI���VN�^�k\��ڳJt+&r�^Q7C�O$�B,!�h��'�F��m�H�!I4�oZ��vd#��d<~ӥ��䥟��8=��(]U044�`��
�$K�S����}�?ATe[�R�=�τ8����C��m,9�`�_�����l�3k����-u����7n\X���9�NK���tX��څ r�)m����y�)�c�;�)�h��mMs�J��<���L8�I���0�J+��^ �@6�Ȋ\I�ָ�<��,c�!Hm,E�-�bnژS-ڼ�&�f��I��V7���S��B�V�"W��'_o��Q1�9����	���ج��L)��I�9X:g� �ĝc,%Z����V�
t���4)���hKX�Z3?I�'��~\"z��}]�kfX�{.)����E����/(�c����|\!��]7��06�6BH1~��=b��(���n�[ڰU�1�,����5� ���zk9Z�'>��med�Dm<�3[�(�������f>�e��ڍ�خ�bW���!����	Ĵ�@8:<ׂ�A(�#�'��:U�(F�|܅���wAT��O�����	�PW`	��)��xTVZ#�`��1����s�1(O@<R���m��X�:25d��8xJV)���At��Y4��y*�맋&׵8ѽ����[�Qz�vgi��(��P�g"a��(��2��u�U�>#�˸'�R�!�e��ȁ��K�{׆��9���̹@�.8$e6���#�8+�P9�q�/p���l���z"P'%�O��F����ԍ��R4�����M��X̃i�?�^���d�gzQ�uQDޤt�\PUa���YH�sf�v��*7�2D�(= A�����f�%#�p�s!�=�7��� �2P:�2$������E���������]���,��a)P�4b$� m�P�'�\����?/q�ԩXa�H������?���q��|��
�u7ZU�:��W(!5��K��`7��l!����p�)9AG ]N�;�����Er���A�n���\_�F?��U�q��T�Γ�dU��G��`�<=�T�����|�Hz���4Z�v����������|`G-ph�V̿���ik��!�Fa�BF�h�NFm|ʭVL@ ��h*:��J�Nsm�dx:�Y��}	qSk�x�@+lm�$=Sv����ʛ��Vd
�_i	:;��,�,!{@�5o�+`=7�W��Զ�d��5R��"�#�h�Ǳ�0�_j�ݭ�Ws�zl"�O��#>���q��}�%4��ً�N}�ߙx{����7�%���3yߞj��0!�#�H'�8�Q�x-�֭�$d�y�(��r8�C�1���%u��(& |�M]�{�^����{�,�?>�\�A��`V��Q�8^@`�w��7�*Im�~�wd�D��<�����3(�3�A�3�w�p�ə���RP��-�ޗ���ș37�]/<`@\�a�
6ҵ�7���co".(|-��!�C��F�!������Js	���=߾��L��r�G+8��@�0� �����*SZ�)��v�>\������r�F��em:#�j8��L�_.�Z# ϸ�ą�������һJMEv�����f�D�U�&x����K�vN�Q��A0#bry���L�&�c ��|2�qU����J?}��X�/w�Z��f+��͑�k�Ì6[k�S*��ٱ+� ��%��q�#��w �.��6���庘�f��9~*y���5Q�?�[�ۖȊ����N�X�e"�$3��q�Ⱥ�:%�������@��'���hB!Y��%Zz:��d4	���`ϟ�k6[�;-�A߽ޖ�f%Q���d�?�{[���ؕ������z�2�O�>ٱȡ$��C6'��33���wh>)��A��ŮZt0 ��Lq��#�� 5���[ow���C�D�_����J�)����fOt�W<x�,�9N����q�?imk'�|�v7��-7�uլb�Ƶ�\�ez����K���:��H���l�\DK$���d�:~hg)�[���5�� �^/3�{��g.��륉gh��lb�-;�Iܬ�}ް� Pi� �q"P�GI��>��<L%��/������gƅ���*{v5�x�n#��/������ٽ�y���^w�XS���N5G����=�fZ�i�+��ݳ��^������芆F�D?sы�o�t�UB�D�i��[�)g]�f���B=��#Q@��`�.O8���#��yHh���2;�����:�F+I*����O��]���[QV)�ֵK����)�%̜b�<b�sq~Z���z�EHճv5i��'�/���{ͯ.ֵ�� wī�b���g���T��Z4G(���r��jS�y���z�����;�L��zw�t�--�=�1X��K&��k#0 gs$��]*0z)ϑ*�B �}0h��,2p5�_+uN�9bܑK��b9:������Z��Y�󹯕��:��}�1�@�Ǒ�K($qac��iņ!qRmb�dY��6��&����g�с���*�E4�NEV��F��Z�GZ��՟3Ӻ���n^�+�m=��A,��~��~��
���l]�ר�*۷u��2Yp����*<�`pYfg߷���w:����# p�}1�ID�z2j�W����,%)��	��c��|On�f)E�li�BKrH���P ��f�	�[r�<�U�C$O��^�I��Ծtweb&�Z	�W���o����v8�o�ُ	�4#��n䥑�#|�s?�Y����E�kb������dD0<{t��U�=��q
�[n���ʄҙ���|�7M��Izэ��3�v�"�эg�՜B�D�������|����(%��n2�T㋒��\�T�h�$��=����A�$���na���Ł�0�Slz�ii�__�ؾ]������r��|�R�w���s:��d8 �{�~K���1i=5���n�`��{TɳCfŉw2�d��8$�oT��E��Ճ��Oz�}�t�O|gl`�+�j/D�ҍh�nH�O�^9۰����/�
a���0_�|�"v�P��?=p���3L��7{�2xq=��״�2b��y]�xOY}�q�	.�5
��!*��K�n���(�~N���s�9�����vɥV&��k��C�c rN[zh��1v����ʙ:ST$\ٷ�f�K���(ZS��x���N@�LQ�e� .�I�X�@6;���/,���[c7�fE�-I�!I�t����LC���v��xx3��sa�I`b��� 1�B�}=�;xmvKo!�V�{1X���l�Q%�a�f�q	��by���x�A�4�,;\C������0����čڔ������k��Og�,O�f�kE��&kLhp��έ��s�E�(�6�I 搴�O�h\�A�V�����;@�i����s�խ������u$��TP��;|�<L�����TU~"7���B��b��=ȣ.��ǡȖ�놠����Y�������p$�X���sސB.~2�FJ�g��\���s�'$��Zf�>z��GqP�����m��g��H�J ����^;U�h=����a��>n�^�GM��kJ�%v�ۼ�nk�M�;FJ1����^M"��aT��nXĿ�А�F�ko���}����c<�(�!#��W�/���>(6 3���ɜ+��"]���$Nf-K�e��&�e�Q�Y@dwq�"��!�Rʱg�>&�E!���Z�����IkEC��PJ���H�E�tv�U!�B�����Q-υ�N?K����H�0��֋NRE{#q�oWS�-�_��M;�����K
#��f��WM�h���<���9��w�=5�u�v!��]�����!�/���xT4�\��������tC�������;煐b�U�9�B���ie`W3D�Ԏ+���ݙA*F@�VT�]�������ѥ��#�(�M��ۧF�`i�'/��&�TUd[{��g�/�G���(3O��+Z�	yj�3��8ƒ����5����K�C�oM�,W�9lN��ӊ+�ϟ+&Cۦ�kim�^�~��^�/Eゝq��q0ە�w���"�@p�E+T������̝5J�La�vT����������`��t�&�f~�д�n�׷z� �_�1�Y/-G,]?F����'�>��l���a�+��K��K�	��4睙_`rA�ޡ��	5:�_�J3�X���2�j�D���ٻp�utT�_I��ߴJ�66�9	41%t#�Q�	��p�e��<Ƙ�GВ�9��ȼ��[U�w�pR[5Æ�PBIe�Z�M�]�_�X�,��2���S���ԓ�t�B!��ļ/����G'��-󏰜��?��U�K�}����8�q�l	��ya@����ï@)��Kf\rOo�s긦S�s�j^̄�J��(���i�Zy洳���v��uE��gH�Ȇ_M��d��q����f���,�����B� 
�=`��4U�p��gw�C�F�#�2��t�gup9���R�Ҟ^eo�(-��ð�[W�jE���`ܱ����x_hw�m�T���/��Lgx=��cH�9+s��/@a�q�c-{1҂6kOz���)����buWB�+�{�/;rߪu�)}O����lFc#+���Z��킜=���g%�X}ݯttX����
7 �%�U���$�c`�1��&d�3@k
!�S��|��\��|:P����۬�k�N�`BTT��Q�;^r~�v��5����eaX�)&�л�j�H0�JH�P����ġe+�%����������b���3撹nW!bȷ�X�(;��l�U�庠����!.�C������c�#�V`�h`�$�d� � 7_�6ܠ&j�ֽeg+JQlȿ۳-��˱��Ň+lR��0ʖ�_�6�����+��ֳR����A	�b�g(xt9T��#Rv��Pưc��&��*��d�8E ��Ҥ��S���Cy��\�F�j��+�/��ռ���1Al4���n�mA��.kY�x@=O ��N4�ٚM�m�D�H#<�����R��6RjtT����I)���#S��5B��=�ŹN��{�+7^����	�Q�kKL8�"_'3�d}Uc�����r���`��!���P�������[��c"��g����N^���!�����n�\A�{l�!��fW���E����n�~�P�C�]A)/_z��U��<;L��rGH:��@�<��h�v�u��y��\# �����J#�]��CU޻u��,g�R�\��E��ץ,�_^+ni}��EԼ����Ȅ�"*2��<�,�_�}A�p�s�����Wڠ���zlB�Au�>ʞ�q0;0r�����='��O�|�3?����=6ޫB�C����-���Ͽ, c����Yu�z߰��I�<4����av��ۖ.�bg�̑~ۏ�۲3;r	��*1֥���l��q��2Q$���N�P�v)�HX3���~Ӳ�G�K].@I�N�����?���Z��>{����Q�k����}ϥ�g�O"��_Xs�ON<8�x��x�i�+
G��Ӝ������]D~E�x���:��n��*��_��/12�/�m��cF���&��Y��5��W�h!��������-��
�;��9�ۺ�>�;jq$�i���鉧x.ۅ�G���Z%3�N'}�	�]��!�FK�1�Þ����/�q�G�S���T�%`A%����5��o�~�����7�^۪0.���71Vm�pL�	I.����D(�f۪�T��V]����~n����0+�kw�7mjP�ZTJ���At ���$�A!I_�jst�!3b����e�r�[��֢�r����֢Ɩ�R$�%6���0\���8&_i�:�ܽ��6O]��Z�Qe��gg�����PJ_٦�҅�e��Ό�38�$�g��VB�H$Yz_W����5"���%�4�h��6�JBƷn3)/L�-ǲQ�J�vQ�>^w��p��<L�%��c��#M6J>��ńͳ��<�����Ad�H��"��ƛ^DR�\>/Cw�$s���@J��(�ؓ �ڭ�N�gx-�����+\�xq1G�\4Z�Y��ͩ�)������j`�B�=	�.+�U�Ƞ�n�q�����H��kg��ۇᲳ�pQR������z�x��wCŭ�=�YF�yj�Z�������>#�� �i�D\ȓK�������r��}V.k��	u�Jse�_��רe�Ջ�͑���$�����Q�'��*!�((=V�3���kt���ŻaD55^q��L
��kt��ϯ5l�S-9>{��r��k��A�7��*�_�J��p�\�"��*F�V?w[Ԟ�C�!A��mOn�Gl6�\~�������*9���X�u	(~�l�R`6��ݶ��(E��bm�I����O���q)���ӗv��U�s���[��c~��)&��C8�i�[NJ��N���O-|�S�g����̏i��%���l���/?~Ĥ9��s�6�cn����Cw���ESq�V��g�;���[��x�=w㲖�R`Md±V�
i�/�Zl���H予����"���X�
�_��l�0[e;MȴP���R�y2<���`��,���H�,��h�x7~��6��X��j�w>���>�VR��=6�.$Fm�N� S���q�%WЈ�xSޗxNI��kY�Xd-��]�նvO�w��_���y�&oO%��0�B�W�N5�o��#@3[yL�Qt8��y�KYi�Z��Ò�oL�۵M���v0H�!`��X��}�L�<G�7��rFA,�Q�2�a49��-)�����:Q��"�c1����(�'k3��S��e�X��g+l\�k��(h�� �ArQ�I�J���s��%((���T��2�"h�q|��[��!l���ZZ4p�S��`b<?>�C� �4O!} ��Jy���1g������U� �U���t�k�Y�Zh���~���xT3�ȶhO
~�J����Z�E��	�&U!�y���㣜Q�j�u��Gz�;M8��@?/N��z<��(=F��Xbl�����B6��6��gw�?A_; �7]?���Q��
J�cت�&I��Լx?�����򒿩�>a����g9kA������g��j���s E�m��*TԨ���%ZI���	K���,9$��I�ΰ8ք�s)�̖���u?o�ꊋy3��U},`�M��ج(OS�0q�:g2���m��v��W2ݾ�S��(��<8"�Ǝ6����<R;��n��k�He�b�5i���ϱ��#��O�5<���bG����k��Hw2#��&��h�R)WuUci�:�{�3��,;�B��#�ʾ�ڸ��dG��d-/�=�h�(��H�k��rLV�kg��� 5�ϛ'e&���Guyc�Ǯ��[�+]{J��SI�Y�t��P7n�vN��ĶG�/c�d~i���`�I5�x� \^4��@wys�;�_��ވi�o��S���Gf���"2���$�f�tu�t��sŌm�A�2�7���~5�M�d&�r,��	��ݨ��~bw���$5O���ɱ	w,E,���l�e��$�(������L:��f=��g�lB����\ܐDx|��;P�Pz�S��gL�sO[0�/\/F�W��)HL��"*y˜[��"��=�����3i ���56��؋~(��s���o4��olL�%{� f��Lx��$g�qK�{��ĸ��)�3l-��a�lf �*��ٍ�-mXKU0	��>�����jz=Wj��v=l �@���GH6E�ꈭ�D��oe�
���{�g�m�֢z�7�6�6`��HG�`� �P_���6�E��8�n"�`�+w$�-2��{�|�6�GZ��f�����C�
Ƽ/��>C��X11VD��{�:/1M���E��q
<���^��舁�F�3�������N��*�rM�6�dc��Wp.��������>(I3�p+��(���0�j8����7�~�m]��h9�����?����v�
�ϑY��%Sg��S���}���iܢ	��Su��,�6��q��g,��B��� ����}ۯd�/-t�|��ڧ���kl��a#ݾU��7��H�0���u���N-�\��g [5ʹTQ�D{�cl���bm0��T�&cy$yw��
�ё���|ϩY��=I��Ge
�ȩ2�78�ղ���/�!��Y@gұ��li�Ah�ÑP*cP�{�Iu�����+��恌�з-�ɗ �q���C�̌T����@1�<�<�D
]���FV��ĹO�V�+�V���+qu�h?{Қ8�ٚY�ի`2ts-j��M4�]���ki��Ƣ�8n5zA���������;�u��f�����s��?���n��!@E�{�=�ߥeh/�BH�:�(���y9��̲���D��o���Z���S�U�T*�a�>��
ʊ{um`��,�-C�HHc7��&�`r%��D�����Jf�U"-d��|�A��g�=��%M�\LSB�\V�.�:��}�>�Wl�m��U{��|
�u57E�9,�	6ꨜ��oC��������b��VkeS0�s����呟�2�C#DLG?��T�A�ceBp�{��y2Osd(Y�k�L0fd�DG��o/BЕ8Yb���s����+ſ�>�j[�Z]�N{�<\��3p�����JЇ�h������Z�6�$F7KS�>��@f3x��g�;�щ	%�G�>n����@d���x;GL$�;�*������u>n���'mva��u��W��,�Fe7��HKZ���P�����*A�Xϫ�eKg�Xғ��q�Tرg³�o��(�k1r�a�)�X�U�FbFY��Q��=�y�Rr����	�K��Sw�d���D�l0.G��w� iO�*V�s�V~S�|�D�P2���)L��*�&
z���y�r鼬ñ>�uy�`�e���үנ���إJI�rJ��)m���E�A�6��¿���
cN����ed4�]P*�`�י?��,�K�G芕KJHF�@��]�.e��{(˞G�\�ۀ$��ߣ6��z��of�.�G��,��Bg�lw����5�a���[m*�{QZ��>2��&:��s�ۗ��nĒfs5u(��NI+�tˮRxgvW����/U��F�����?�4�� �Q�kF�4��uJ��+ݭ�����.6��d��tA��6¨r��-�\�X�5�s���o^!�e7S�����;C��K��p2��&)Vkt�a'P��&,�W���^��֫6*�>�LC�W;n}1��n�(%��D3�@�*3~������%`��P[�P��?'�$5�(cGzC��",��Y�@JLQ~v�I��
'62�h]3XUM"�ƾVt���%
%u.=��+,��M���E�h����� ���ŷ�9t��E[��6��K�^-�$���dx�dO^���:Ia	n
�[��ohRh��Ϲ�3�ڽ"�P��b�Ϗ���%�EU9e���Oy�vb#̶
r�)�w��w9@��+i;3O)
?b�c��cC������V�|>}�?���9C�ܨ7Ns��	�fe��q���&=���ü��j��]�:�i�%U�8~Q"�O��Ό���&��+a�^��~�L��*�>}����	�藫m�=��r����x�p��즸vQ>4�ys'�4�ˢ�'h�q��:�����D�e0�N��+��X����x0�=�si;H�e�n����~��S��yݶ��j{�Һ������4F�zY[���^����	��0�M����f\���VO�y���.89W	غJ$�����%R���Ŋ�����݆�J�!v��#��hVCM?9 >�FT՗Un�45&��������P�(��W������|��'+=�x�θ��kU�cZϡ��@o���A|8�v%���ղ@��ێ<���΀))�LZ4�^WӝOk�p�m�#~��眥�O2T+YL�����'YJɀ���K�6����������[BM�i\$��.�����u�5S���	���X4�őВ9u-��3N�x��h��x.^$��ؚx�?;˦'����B���;M2���4������\��t펂)�l�4	s۽���PU�m\'�ƉJ��P�_�����̄��Ǿ�����-��I�4�#M��5��U��7���#\3{�����Ī{�s)��O���j9Xfѻ�S(P�E-Æ`�<0n�+zg��	I�M���W-㲅Y.?��;يT��k��Ϣcy�N��vn�oVR@��ã��,��sYY��4|n��pT%�u�$ ��d���M�B��N��%���D�&��e:J3�'p3����ƞ91���ؘ���� oW�[�#�}�C7��+�vb֧`��p^�`����nD'Ҡ�XZ������3�+�6-�O+٢ٗE��3[��
>�y�O�=�+�J{��	�_��`!߶Hjv{)�!�C�����aŇ�"�d(E�洮5���k��ޮi-��P���!�X���$1|��#���EF������q@����'��Y� :̮��mei}�-���:c=bM9���Y�6�?h�h�VB�x�m�[Y
�9��z�{�(~�sD��N�k?�E2�i3T@6s&��U �UVl���3|~�U!���cvc;RŖT�rP�6���^��1�����%�0�_�S,��e�LX�oƱ���C0p,i��C%:�DnYB}�D�z�+�#� �r��Eܼ{�\���&���a�hI�tfu�(���C�.%C�w/%���׹.N@�=�w�3��ʈj��v	-b�$��n���;��J���W�Ш���L���A;T���������p�!���YDO�0�8J�������oX�5P'vVBj����3vN�ϭ��}��U����
6S�(��H��Đ�ϔo�o���T�؋��]�{��7�,���v��z��Ti�!�K�{�f��1�3� b������Ζ"0$�p�vH��m|�y���|���� �%���y�����WU���l#���6�"�\H��8!��?�%I7�5��#�$Y�bh�T� ���'�z��\����1�6�CuP��k-�̈́1Ɣ&d�-�(-���W��S��wd��e�0P��%Z�t����v+Q+����>����"z��USъ�sp��3�"�?v���'�Q��;yb���"gh�J�/����=1?ݙ�e�7����k��$�Ud6
HpR�b�$}Y���׭�}܇�l�/��c��8����`���J�p3ZM�r��Mw�%�70���H��[;ډ�7�������ϕ��z_,�b�7�9���! ��k�4���h�0��\@NN���٬2@kܯ|n�.���X?/��xX$�h�\?�iY>
�m�G�}xyCD�$+͛��߱�:�M,�4�p)�֤o��c+�Y&���O���LE�	{��#����nڵ#�M�F�/E��C� �l�ϡ�Y�c����{�Y��Ŧt ��J��8���,&�e4�chu�K�1��"��s�S�;�$gG����}�0���ek��x��|�]ɐ���'oR�qGz����/���R��ǫ����p��<e�A����A�8�$��S!X	h�g��׮
�� ��2=�_�����E ;�si;�%&Z�7hͧ���8c�âjk{�^�4xS�4���2�E.��FP��sLch�	��?6c����
b#�]A�U�9Č�#���g�[� ��i�6�������z�E�7g�BЎ��ǰKH[a$B6��ހ��⟶�F���Dgc�i�Y)�1����l2KQ����,�Ϧ<�Xd*�Z�>
��Λ{<����3S��UYY�#����([�ؽ�٤]���@��p%����dьp�ⳢqY�/nc�I>T\D�1x����I�c��f�n�rz� 	}K����:adhB<��>�=#P��o��#7F7��B�ƪ��hĕw��f�ګ�G_w�;���=�6_���Nܛ�����:�a@��,1x���N���D����<��K���P�>�] �\O�����]��+� ���o�t (D��l��A�-�3f�>>�F��0^�`�S/y��X�'ُHF�M2�j��f�? t!)�J��F�dA�MLc�c���cyLt%4��X���Qk.�I�"|vx���C�^�,���ɚ�k�i,8D��<>~چr������g����.�&����Z_�t��1��M-�
B5�����l'3&��w�5�WhC�Y�S��r_+=D5f����[�����ޚ�Jc�|CW����v�k@��~��ur��C��xOsS.�.k)ǴLK��\������՚!���;����G�8 gj ��1z4���q5q�CK�&�b��=��H%Y߳�0�H��!̶��L�U��?�}�xn	�{��`��)����� �e�@���2��%(SH�b׬�iũ�o`���sFOu/�����#ȳFx�S��}<x���XA�������Nx��2,�����n���|d4���V�e�p���$k�z˘Cұ v�?��,(M�L �Q�o�i���b����K�P�E�Jid��^To�7^��|��t�~�k����6��&�m;#D^�f�D����rO��1R�{I�䎭+Z���y�R!QVp����?S��;ӳ[�Y9���U�Ɛ�c�����7]kNV\&��3������l��KMA���kP���"c(�Т�_��cU���{��.?�j��t ߶@~N��\�eZ��P����ևW��&Y��R�o潀�~j�Y/uW)T�>��:�5�A��E���c�p��:��K��wuf�V�K���.�	�?��������+���g�P���kb�o@���������q���B�K�;�i�]����2=��.=�a5f����Al|�C^W��Iv��`Y�ÑaLfW�̷�uL�����	ઁm���}�&�Ed06��97w�0bT������@�It�M5ʫ�q��
��:7���5��UDK>��P���J�Y}m�Vо����ħ�@W���l���'�צ��9n"`�d��q�#nN���x`���z��w�j��	+AEv��w)�4�l�s;JCZ�������nS� �>�X�����*�*'A-��xqe�1��pr��.6��˦dt|�Ѩ��u�5���h�dA���b��h��t�J�H�����'=)9/v�踔��.2�Sg��&��T��g���>��t�{ORm�6�D�-?[U�-�x\�mU���!Ci��P�~	�Cd�T�C�h,�ъɑqd��/5t��ɼ�t-]��l���K`���3����cZ=��W3ZE��F8Uk�0��j�c���W,2$��G"�$�d��W����m��y;56�xSZ�Hdj]�� ک�i*�#�{,�i��3�T��o��-P�9���ϊV�����Q�j���B�2rǉ�N������Z3I�@��\�)/�>@�Z{6���!�x��b�2}�8Q`2�w�qj ���F~:Ml�d�o"��[m�u�5;�g��R�j�:�Z�,p5�$�se+��.'h$�+��4�٠��wE"?��W`g��r����f�M@7��#�~M�?3TlMg�.��+��a�����-�p�b�e/��A�Xd�asI�*ٞU�П��2���t�+�a��vKPh�+�o\���
Sy*3�����m�i��$�C��QQ^��
љ�u�Q�^�c[-ēZ���4�v�����s0;���wn���L"�p�b �&�D�-���?�}�ei��/	�C+HM��+-����ܭ�śq_x�Ҷ�6͠,������\���^0�~�垁m�>����B�^�çFބ^�
�,�x�(N,�ȲXVxlR��y�K�����`��t�4C;iU�k��6{�Jf!tԚA�>�u@	A8��l�KN�v6]�aS�)�Q:no��cD��ֱO�E�4&���ԾҜ3	��3�5�("g8���{=����;��&֫�OX`}�K8T�^p;�f払Z!���?��;�!���18�����}c��GP)jD�PZߒ�飮So-����}V�?�(2�ӕ���ۘ9�u�tG(j��d?T
�H��Q,��a��dlf0!r��9p���w���Biӻ�a��B{�3 l�ú.^f��u֭z{�^�xe6���a!��vGc܀�v�N%�-SXZ}�������,�\\�K~ ���J♧���˹!�d7e>�	�xCgUPuXs+����B���CM��&ܑA��w*�U��io\���Y�}2�%�=c/Me4���a��U���_Di�g�
����z�k3'-\E�P$�����\�"y#�I��8hUd}Ms�����so�7]2����H�ݕP}5XȘ`<@����N��`���3�(��!ԳR �*��F�ߔ~3�w�`8L��9y�G��?��������3�D��
��?�'uH�G	��nvΐhZ1L��~?�$Iץ{�	\%� 2[�jg{ǫ0k�K��ԹDʷ��N_�R�2�q�g>������k���*��
F��L�Gaz2CS��[K�;�4�%5�_���o{�\�ځ$STM�A1��W(+Pa	���|F�[G��:�L�Ŷ��3��	��F�H�ou_.��j�|2���+s:�E����m�����?����g��d�A7m�9t�p��(�>��p\ߞƑm0#�cuS��1rvϭo�����)�u٦$b�Q���*���/�G�D#�h1 ��B]Ƹ,�Q%��q�.i�s������EL밦��X�8@}�+�I0���qQP<d,�S��AZ"o���p&�=utg��әi@ �6�X���xW�Ę����ܡ�)��]i��/k�_��0d/EV�rZg�ad&H&��U�92[#�#��t@�MM����<��&�yKU{	�����#T���. SV�<9�#>YF��9�~:�$x��d� p�K�
ǨT@W`UH�!7�a�KlgGbF`��
f��y$�(�>�
ȰV�Ε� Xuk���*qdAa�Lo����ih;S�
�S�!�Sat�ԑ6��_�s�e9�����W#����'
�>[.�>Q�Qu�G�w��حd*����Kϔ.��m��J�����D�?��(�k�Mꐥy�R_�c���P:˸xGI�DVb�;��L��Z@ͪ�{[��5�9q�6�l��E=Gp1�ݯ)?�e�	��*�������+n��{K8�U-`U�݀XS��6���:����n�9�';V�e��6|O!'����.����Q}���Y7�����T/�=��zF�o6v�A}_Y_d���q9:D��6 ����&e}R�e�L�GT����I�{D�p_��%|���5��m�����}e��B"}��#)�w&��$^���%�����j~1B�Pc hh�#u|b�Hd[L�����r΅=�x0H�1���_�%��J�Ώ!��"@ŀ��'ټ�,���C�2��p�]���Y�����Z���Hm�ES���� Ģ��hT���.DӦ �f�r#�[zw4~����)�t��v���R�*y6������[� ��rï����ޔPڣ����u��m��s��J DPz��������DP{#��:k��z,.c&!�ѯ���&D�R�'�Y��Hu� ��e�%�:��6f�p���j�bݣV� ?���B?�V}_��U8�����5�E�<4�k��(�u�V����~hM@����'��]�8�dP�@��7֏�4J�O�����Aޤ?ԁu�>f#�2�O��2��թK[)���Ҧ�!;I�V�gz(-��}��9#�����q�����/B,�+�cթ~�>�>m��9[�!KR(P� Q����.��µ���eQ��D�
�Ŷ�
0hS��C�fVɀ�Ԥ\��^a���ܺ��2�c>�#c��{�k����J;�V��\��nj%�"0����h<:�D�@!�%��$g��[-���A+�z���t �(�ْ�2��]�r�������J�=��o�P�����]rJ)FЁ0�Е/!�*d��rn2�'�x�/P�Ohbv�r_<	� �\� *O��x��EC$M����91�{�G�.ʸ+�B�s_�Q����w�?� '�;�j�9B��2��a<�&��HT��Z�ٟ��L�'2��ƌ��kCM�̓qf����^&	Ұj	�\c��Ш��-&8	����]��º�|	��r��g:�4J� ����L��, ��R�݋�g�.�%�#?��!�s��ώN��8Օ���zGMJ7��3׃��S��;�9��s]���t'��G���lkS�.��ZȨ����j�%jyf��W�^*Ny��@J[	wyd ;i��<�L>��Τ�D������hR[f����+�?G���eg����к�t~���	oĴ�+Q�q�g�zU�B�I�V*o���Wo�`�&�t"�	_���k!����Wv";Sد�=�����nnv;��(�J�`Rt�`����1C6�C@�7"��7�q�"��@�2q)��cW�+=���ݔ�'�߬R
�~���m��_P�	P9δ�j�>�#N V�U�J��H����$�e�6�C��)w�pjz26�-��j��׍�����������u~h�����d�����c:e��P�&X���vM���>�9#���Q�G�����ʆ�\à��A69�35�L�0B��R���F�	�����=��}���Z���@�rNd̩�r�"���[eQ<B^�Im�_shv��J�[�Y�W���%*gV�� �Ĕ�M��/Q\�X�ͻ?�u�ٙ�,f�Eh���ϥT�٧~����]łG<��k�q�w��]�����d$N��r��V�	#�o�����a�1t��9��8��yRF�p�� ���.f)�g�뒛w��V��!�"�I���v��`C�lc�j2�_��8h�d�(��*�jB +G�E2�u��N��P�Ϟȟ��q{8��(��9��{�l;QQ��J�����O���>Z}	���A� ��j����9BҭB�%�3������Y��M��5m�<�`y�IƼFa'����D���ފ�\~�I&���z Aͺ_  ��/ʽ0�}E�ns���Jx9-��p�5Ci�q=8L�����d�Z�[��)�A�����˝f}�\����)����HeH|ѱ�hF9�_��!f�����n��F�zL_� �U�V�a($i`���7�Y\�BΠ�O�G��"���{P���\K�?\����%E�U%�ǜI�h�poȷ���?�f����X�l&��L��D��d)c{B%�����j���@�n��ύ��L�j��UQb��,��w�`)���\��*�d��ޞ����^y�:�e�M��x�U.�h�;��.MޅA�`��`�i�]����@��2����R�5ΉUNϋ��-��ԗ���+�'6C@H��%�vb�i������U�r>(Ǿ$Up�C�u	%�1��H��4+(�qd=Lw�i��"������q@f}$�X��W��!�fJ\�Z����S
:��4��6~S��LiȚ<�$w��`�HX�y2���Z3aT"x�'o0۩�w2�2�����r���(�t�#:�7�;�b�R>2�KR
MVo�:2$t|KG��{�����}ڳN0�s'�� �VFmkTMp�����]��|�)w�i����	&�>O:Dۢ��٤�i,|��o����?�K�i�=��a����{V+[lA�����;�˥t>��:	�OY���0xέ�7ⴈ�d�䫆��\����d��wwQ_��D/ �BO��{��9�e��_`]�׼
^���Y(��˕�%�5ē�~��v�i�a�.u�@UE�7\��Ԙ1X�ص��ܼ�~��U�������hd=-�!
:�� t��i;�N���8����Y�Z?K�}w2	Z""��#
��$x9�H�"�j%fkD�����٩(�-5�̲��+.���-8�:�
��	�S�U�ʹ�d8C�5c��Y��d�4ǵ�|xz�*?��C��؛}f��� �@Q)���B��|������z�ͼ]\5����z��֝"u6�b�i����|�BOzu��#�݊%A���xc(]ՔB���r�3��$P�)#�V'��$@4e�D^���� M��`�MۅV�D4��o��/���<�7��xIסE��#�П�Hhq�u��~P6���:�f"�r2��gJ~v ��[�r���Q�Pow:s�7�5��Ax��Nv�?��-$-��yr4��q�~�EJə/�=Dsh������|<Pf�,�]�#��sNϧ�B<]��:�CH\�,�@w��:�g=چg��#]�������}��gy�8������
�i|��-��*=�|2��Oif��Dzk*;������{[E�I%=Ĩ�� ɃR��]�䘘2Y�n�/=�o�����1U,�P�뗵BUJS	^�9]��#�s��L��������߅�!p2�&��*s0Ȗ��ܱ>pxR�k˭]�9sAU-��b���@�Ů�Vc���c2i�-�*����i�d��$�M/��)�c%��]ck~�c�%O�u�Ժ��}�'w8�e!�(�2xځ��L!b\s��mJB�)�!��+�^�΋�A|Ɔq�_8��S�R�X�6+z��ܔ�j�m��\,�n�eM�?�g�7�6$���_żNY?Z���1�����m��ݎ[�z|(����t��W����˶�f�b�,�158V#T����)����~�Q�_d��:����w#+@L�a?Wp}��,��qu�'C/��3kZ-����%Ω%�	�gb8qTP���FcގdpcE����U�$�#R�S�r�����nvʢ��Nl�lPv1]��D����aw�������yPcy��qU5�[hZ�u��U
}b�����fT�kXAr��\��E���1�IL��%ѳ�Vj��m�z*%�X=�VF��3Z]KEӒ�ڬ��R���*'��E����N�.c���T��|��L���̪��i�󳨮B�O�zr�o�<{��>(ȓ`���a�,*Ɔltğ�ӝE�U+iqD
v�v��T��ތ$�.��Z����q0�mR�ߩ���#��.�|��/�@��̈́�i�*�G;�3�M�5<�4vo�է�3dW�t�N�A��+�[cۦ�!��Fh� .�CN�=���+�@���e����X٩:�F��C�~[��`���K�h~��Hx�儗J��p�6}�l5�?��j�������`1R^���.��68�����GI'����X6���Mݻ�9k�ͮ�lExޔ�:�Ucn�3���4��de0x��$i��d5�(�Y�<^V*
���W�6y^�8����>va�	�L`�#���C<����'�;��`�Quu4K�I����~�[��g��R~f5Ո��\��(é$�)㬯	��m#�s��v0�4�)t����hE{ߘ��{�Q�bH�g��uMr������4��#5g��c�j2/ �J�!�s~h7�4* �f�dV4�I?�Wm	�Y�S
���?$4���q�_󊵚��:�~0e��(�Jm+O
��g�e�
��y�i{�~7�?ڽM�³�#���}��a�?�����o�^�Z�A�x�����1)�li�h+5#-�?���|�0'��s䴷BT������:D��4vk��<Mh��k�meu��Sl���~���ʑ+���Fn@6j��'�+Lx�c��M��EX$�`�����0T O:c��̉�C�#K~��ˑuL+�3�M����Ҿ0���JDN��23� ��*Au}�}]��{�y�}w-�tizt�9�[�tߔN���.��l�,��y���3<	"���Υ3T���&���>i���v�7���ε��?P��۪G|
�����oayқ�+�G�ԃk�� E^��̕=܌rJ{+�)�`��{s�v����b��Q�XMB��U��� (��UvY19��J�j$��SRHd"�'�s��Ǳ%�=Aa%��8�8�W�Vn��!	p�t�Yi�(큎>lsW��u�>��x�x�,)���M����k��`*��wŞ�gk"� �c�i��欚�ڏ�:�(��PPyqK4���ݶ-�ua-�ܦ��p豬VP�Hn���J�Yy}� ��A��}�*�0'���c�$�%��4��/����%�TQ8��/�o�;f������0���u|(Ԡ�b��<j����`e���YW �_�u����0���ã�6&^�ry�q�P;��W��J	�6�7x�����)3�*�����2{��Ь1!���yFn1��roj�!K%�Z�NV��,A�(�X�I]	�P��4p����O�DN�U_#�"���%+�fbb���L`aD$�ֈ�W�/�82*���l�6��A�DΨ����ػ 란9�j�N��!t ��
�j0��~�\�[9�j�ޑ�����ɬbM,�H5h��s����KeOҦ*��3�|�{rC|x`۾1��T�����+Yb��(6%���"���w8�����-�X{�h���!�O����Q)�)�>�v��?A���ACD���qnr��!�xr�ҁ��~���- j���Pg(k �-�xٌ�у��@v�c�M��!(c��y	d�d�{�d4��"�N�}(����'4b���Ye��;Y%ɈM��-<�PN���V�+G���,�5��mz~�{������liK�չ*rɹō��}�7���K9�&�ql��>jG"C@��	~-Lk|�U���jڐ�Rh�mEj���U8B������7�'~�P�|��e�+�xX:���u����ݠ7&Gw��iz������ C��Y$����� ��C��
n7�0�B�
 k
j6��ϥ e��<��D�F��Wʘ�ĩVf��ue�� +�`�4RFh^I�-6���b��	�+�-4�+O`�ܥ<N��tj�r� {Ǯ�Jt�M�뮫�z` *��e9�t&�N�쩽���N�[/�oR�1-�E>�O;�?�AS�Qm�f���0�?��.8��RA��X���Gv�<4�P7�-å�SޗZ��(�yeOB��D�,�����4��W7OFlW6�9/޲@+j��l�ʉ;�3�Q�]��r���Q5�A�]��D����nx �]��Vk[�V��뾽N,v��g��u�#����@�$L,��_���栗J�e�֢�B=$HmO�Ş�ڇ�	m�.0��H`_$�g�^�?�Ɠ�[o'Z�O��Ej�jM�5��r��r�/6	�{Q�)�O ����+NG��3D��"Q�P��bW��o��e��)9K;:����"��2�z~*��x/�vF�C�l�nK�	��SfG�I��NӰ���kJ` ��D�LXCb/w}oc�R�*��O��W��U����=Y��X�PvO�s�����HZ�Ff�E�
���k�L?&�l�*���<k��3�h�e�����R��i_c�����hk�:]���P&�$_|�߁���U��{�ڐ���gc$��/�sQ�!�1i��*�,}�۰6"�g������FA��`�հ�<�E�(��hž���/���b#�HW�u���I�*��)�
�Ր�8�;'���:�q["��E8 !ƥHMå��9���}���e���o1�jA� 㿐p���Z�]����%�� �:��	Ǝ�`�����Ǜ�X=qsG�6	cV��-j���B����@4���IQ�݊�فKU�W�C]�5�l�`EoN��g ��^�m9���܇܂��i� s�6UC�4I�`+�$ұ�����翄�h�Ls�e��KމL�eYgz�R��,�!���@��ϣ��d�R����?���̀��-�Y`^U\�]����=s� �Ou�7.@6}4��XwN�7;��4���\T��3�o�%���t�M���G���S�S�W��|����j���1�6�>�m�	f7�dUwг<��n�:Q\���01G�L�J�?�� �+|گj��wq�u�4�����h��?�2��R�s���&���!�4�Q�v�f���\	άd�r�����7�����,�Ί%�>|sU5�"]�O�P�@B�w�F������[R�+����c�wH9'�	8)���x$��8&wA���fO���t�ǣ��lu��3�+�>���\5���h�P؉	L��\���;�j���
�J	S�=�2��v~tٮ�d����˺������AKq��,���xI}�v�	�0�"aALI�tH>M�^Jlט��ku�>�nqy���X0�5#X�67xfA9����Q���9�: $����Ъ_Kq���MTn���9����s�V����(�U�P*n��|����#��(��M��Z^��«�Q����2���h�G{��l?����A���{�Y���؜��hݖ���=�7�:�[��^����;3��{�����kQ�Ͼ`&$&�]�W ru��+m�������&���o5�2s��?����n���Y���B}��q�jJ��(
)��$ʰ6K���4겗����'x��df�B������N�^�g�U&��&����WN�価%|��*H�"^d^�"s`ZD�4���5��o&xp��9��
`}�s)i���]Ż�;�{��sw�Iat���{E�41�
楉P~�4��\��^F��d����wC;8˂C�&��e�i�6��k��N�.�hE�_{_ՑYe�J� 7��(�P�]J΂�a;9�&+r����j�������54�1-��#�ޏ���+����6���P�ߛIc䎾u3k���T��[M��ع2+�r�[�A�:�Ѻ�����,�n6J*����2����.7�tE���}�/d���.�.�l��nO�<�������o�$p`��q��hX�`N��΄x�>�)���GqY��+s�5���`|;i��ڣ��F�����_?�R�0A��c�G���.�͏f�2!��;��d��(h��6�Ծ������	���Ӻj֪9����t=g�����'k��F��D,@ՑDB���g)�?g:;,p��#ߧC��� _4���Rs�ꎦ��p�,]}TtD�v(�y>+�Ll3��Q��� S/����\ٍވ�}[�]\� ��)h'1Ѷ��1����%�_�6�qA2�)87�_�&�%�e���/2X%���Y�Q+�42�IM`�s_.O�v=}R2��IR�׻�2�[�>`M�o��(�83X��O��͕rE�a��������`���6��XKp�fϦ%p�'#�'�_.m�A�����B�~�R)��w�O]��'��(�p��?6��x6����S^vMzӦ��6�G�D,|�$��	��(v��
�UKc�W�%���D�q�������@�5�rr���#I�(R��2� {f!�{Y�oi_Z��qM�!'�躪�ƞm���<V\K8����@ z*���j�p�6�,v}�f"��j{�R_Q�uh�ꠟZ�>Љ����� +����&��2�O}��m�{f��e�n"h�)W2���i��XDy�6%����' ���O{���=w`����]��y��c�z�v�B5��Z�L�A*w�ik3��	��knt��Kp '��#��/��!|Gޚ�Z���!ΝfÑ7�7�+��p����ևj@��J1��S.Ũ�+�5^�5~4)_{��E�Pۮ9����I��tEo��|]8Q6���[���UW�޹��Q��tտ- �c�pmv�z��̄Y���:ni�߶���5����h��2�ƹ9��l��_Gd�G����6J>�E���׌��k�{/"�O*�
�&�c����3k�Z���'��N Ra�A�LjƱ|���E*���	��/��֘�M5�¶S�6S���\} ��/�'�>0�-%�~}@4��~� 6oh��*=	Q�ͪRebZ�_����q9�P��yC����K4�d���enn^��wѪ�%Lʗ�}j�^�HO�z`���YB���a4��	*�8E��j� Rm���p�Bֵǚ����0���.�|�Jow��8CB�tz?'ј�m�D}X&�>��׸\���3�٩x.Gő7�B��ه����U&�^���O��J�-�Jp`����#[���o)��>Ll�o2^�+*Ғ>o�0.����p�I�9�p:T�����)��a���ۺN�W��٣gʔH!�YF� ��e]���7���(�}Q��3�u����E!�6"p����&�;"
.M0#`�-�͘�&��A'r���WR�y�Uw��MQf���G��V�����W�����h��SΙ�'��)!����?�͉�a{>��Ϳ#񂺔��1��!�Pr���A�'�F�NP[��G�l�Q���D�ָ���<O{�(և�r��vh�.���Ω��w%p�����u��8Ntҕ��OZf��8Ӥ@�3��:��7b-C|�];��>/^M�@A��}M#� ���}�k�,=��/{6o��t��`�����XJ����Ұ�־ҔRG@�:���!iv��}>���*�]�n?���@��G��l���S�0�k;Ƀ"��إM3f�8CJs(�z%�bF�^���o�D�[�Qb�\�]�L�6e�|T��Oum<Z���1u�@ΰ���ـ���Z����x�M��^_;�|�'��8o$�v����հj�u��㻷��J�Ҕ3e'����@V���zF~)F�D�� \&�W��#>�H*����LN��s��Ҙ1]TP������Y	{�� a���B���vWZ;T���n�p���0J�A���ֻ���@�V5;`@�����i-��I+�8��XV���N!5Pu2�^ykۤI�*�gnp�J�����
�TԸ7��NR���o��8^
}�ȵ���v�C�F ���tI���p�.:�`���Oކ���[�P���k�	���kɹ�`E�S��z:_� �yؖ�?�j�}O�荴ǘ/W�_�m�UvNT��u��BG����ž{��fr���of�h@��F�O%
X47`�(�N�0��P�=	��������wԙρ~���;�80�$�uW�tC�V���������+B�*#���&3���Ew���^��߄7wɐh*T�گ{�F#
U.���r����йi.ޕv��������f#7�27���$Z��S=]�8�u���
5�-������W�	�sP�x.i6�p���D���@A�`��G���wܻ�Y��Ƌ���ɐX���S&���3������d\л��w싹y�׭�4<	ۉp���x%.:6�� �nQ��o�b��o3�CZ*W���IZN�Р��x���IC���b|���2>�]6X�ǭ�J) ���V��I�ط��|j"I[���>�ʯ������u5��Df0si�%�Y���^"'e�F@�X��+��٦Hgs��rǙWC����"�c�+�L�P:�=$��rq�G��}F��ZᏥO�l�NA����
"I$��y�Z���jfs���eyN����G`P���;`�l�,Tj�i]�lQч/0z���E��S�%v�mE�N�E"q7�`*(}��
��`�6��g�R�����5�
��Y�ۢWqw0́���'i d�r�)�\���M}�����";|pv˷��V��L��N�=�*d�n�|z���b���9�ۣB!�w���Wq.��%:��k!h�|G�Ⱦ�'� ai�KHb�����>�[�S���n<$I��V��Q,��mD��E�]��������ľ�I�y�
'6��)m�)mq��3���:�H��Wlu��\5E*c�N����n:T.K��*�6uX;#�('�?�_���u:�6�šk�Pg�e,�7�E	Os1��%<�&?��'b �v_�ÿ�K9P�!�@3^ch=��ذ�R�h��2'R�������������'x���`���~!�|h��ʖ!mX դ�s%�Ѳվdq'�\
6�z���_�n��9c�(_v���jxS��"ϓ3�L�3J�`q�>9���Rz5���������Ҥy]t��3�꠻�g"��>j�b�>o]J�/O��8<������i%�Wͱ�M���
\�T6#�0��QmD8J�����2$�m0K��*��� �����7YU{9}��kP����I��P�)&z����;)G�1��ޑ���Մ��u������ZFaNI�e$MdO�i��Ppf 5�5��6�1��Q�;FTC��������ꇍR��lF=��NO������~����y�$k���u�@������I���ӡM���d�yˬ_<Z�
Zk_��-T�/i�~ R����M�g��$�m�m�)�R�g9�zA�������-ӗ����b:!X���IQ%�sa^����ƾv˜þ:3q������f�AJ��0Y|�}�s�]�+*���Lg�o�n�<�ϢE��zƄ�1U�@6����8�F��i9�I�$-�<��˅���s�-������!�_�&�o�a�>�Q�"�ɏz3YZŃ3}�jm~ˍ�D��!�R�,C33�'�S�4p�cDS4���Ā:E������l�Z����Qҟ�n�xx�`2VNܷ��U��H�o���iV�����#ABXm�Ǘ�8�Dv`S�'� 9?aw�|��]��)d������H5�/��,�a�RUjF��pܒx
=��H��bf�{�P�W�b��y:�9�Z�b�:��0^m��BEј�G�n��x�5&�6uߍ��f�Fpe�2�
p������_)���:+	����Q��������sT���ܘ��j8�0������4G��۟0���n�c�ޞP����"� �n��J�B9�f֦X*T�ר��5[��:��UJ,�o�@���e��)�0&��t�bi�xɗgZ��Q���QI�/z��0L3��F�z�\�K����g~��%`�g0�֖�h��z�7�H�����wg?��t�F"a�ك?pI��E-��raQH�;��4���IA���us�5�����̏�uX@��Õh��f��? ����5�50c ���j�{��[� ��>dW�=ő�]""�6�D��>�plJ/�0��j�#?��1���+?�^`f��;��C]5���6UƔ�/׹���Q~��L�J�rD**�M�����B�`�j����$`��5�(F��CS����yE3}T!א�j�g���d	�;de]�
A�Ӆi��e��ƅA7��')
�����1|K/Mc��ߝ�t�i���}F�8P7������ �nv��\�@�/tKG:����ᠪ�It>��3��EĮ��T��~�>><Dw�b���K2$�W a�G{����S�M��]����B��A"�NVQ*DL Н������𓄩>�tl�oG�#������4B]9&D�0�s�uݢg2�Y0� ����9ۍ\�b=��M�M����]��P���ZQ��F6a}c�����>�Ei�ޣ	�U�*c�NQ���� #����D��&�orS�6��oaGI�Z��5������[��Κb���n���l7���l���h,�LҒ�6T�E:2v-Q:�1Y�M�#�+a��r�<ݏ]
~�H�2�4��zOh"$X�
������eèL�#t���4�3���)֬�^G���덄/��ٍ�~�sYM��.E�i\�=�C�?�0���\��[��؎)@u�}�3����'~���%A�r�B$�u&$|A���s��Ԏ�8�5v�R�a���2�$��Z�Z��~߈:v/m��o��,E���#,-���:�p��1���ƆG��2�ft��}��͔_e0�SHZb��;�>9�Q� Φ��f��&l���p�����aˈ͹e� ��\��[�y q���@�]ˏ8��:��f��ݛ����ڼ��o��?�����'\�@��ĈըH)�CDC���[$���{)�u5�й(���������&;I�^d�K���9	���#�-�ա��z@��A&/2�H����4����TP<�!.v`�&�ur�v��Ԧ�:+Ecฬ�A\:T8�ƕ5�n���N��%"�
�XJy�G��mH���#ۉ��o()!z*�'hb ~�Y�@���]J4��9���	n�:�
6n&�k�X2Y�q�M�S�H �i�����I��N���~vQ��q�*�;j��	�YT�p�X���[5\I:!q Q{N
�D �sp%�XM�(���b}?��jZ��hv����J�d����Y����]��zg� ڳ��	!5�-{��p>���S=��Ck?�W4<�1!�";�RZ_ �s# ���4�շ�.������,�$�/�oYA�4m�u�ԛXW�>^I��'�J�]f��}c�auѰ�s!�|[8��."����H߄o|=+��XT�CD��K(����e�c8`��CQW�8�~KY^���?�����X�UEJ)��[U�Y�/��ф��� ���<*F�6L��Fp���B��ࣟ���l3�*?�1�Yt�w��>y[Da�S���Յw��#K���Z1�uv��O�.��X�[ѯ �0��BH��gv��1�\����a����`w�S$ �q}Kn��6�R��y_��Q^�N�R$���S�g� �(UV��@�TˬY�r��SԢZf�q��>ϸ�Z��+�S9����ɚ���i&�00L���%��|�KQ{���s#P(H`���^֑~91�e�ƶ��*'�,U��j��Q%��_>�a�;����w��Q���|�����R�d��Ѿ��_G�W�J��G!�d�2��UD1߹+�4�F�]�@>�f�R��!�]������&J�0���/Sl֫��G��������;C��'?m�b�W�i�v>�N؊�"s��)�|Ѳ�Bj� ��=���iμ
b�m*�7T�_��=���8CW�f�bs�а{�i�.�y=�x�������b���%b=�B���aE[���OTjx@�T�ٚ�y#����u/�M\12�߬^s�2?��!$5zV��Ρй�D�2��φ�U��t9i�q5���:�4|9��7���ú�|��׶Q���\�F[0W@�Pv��_��� ˡ�vs?�`y!�/N/������p{}s6>}bSpAp����@��[r���S���^��W�w�j�y	wK|v��@2��f-�P�Z�3��mpQR7(^H����Y^�T[��y�0"�
��t���E�׳��m�+�qF7�#BH�9D2H�����KcO[�p���(��0|9��z�RM��:�^}7$un'R�	�b����)]�x|3�5Q�b,��C+�k�	��P����N����d�Ȇ�.eޏ���tXO�Rͱ���H-*b��e���7�9��X�8mzߤ��]�⠖}��h/�Vv����=9k�򂇙�-��QH�� �Rx]y�+,@M�WB��B��vO��>(�Zi��K	70���u�����0�Tb9>���j^�s)K�Xf����sdxk#�X���)g����`uT�A�&�vm�w�Nnp6U�7��Uf"�����Ô�A�����հ�U����E���{`-a��+�&��,2cBG_I�{�==-K%TD����U�H�2�{Y��~��?��u�Y!�KlE1�%Xj��/d��N�m}�$:�4�,\ �]�`��C�MW��$r�l�n�_^��Gh* �]�ɇ�Z��������ĂG��!C��T��kޒ����)�[~�>X(�&���c�<@t�O[4v��R��p�l=�
=g� T�rx!��2p�	Wn���X<"W9K��ɫ�����;<�永lԚg�X��-�F��S�k�:�l��0�ږEDUn{ǞVJ0؛�R/\�M��%!7toLk֖�j5J�z�޸Q!��n�(�z���kM	c��oh����bN�k��Lqw�rr�$����֡K��|\�˥5a�4�h�I��^A6�9���tF�L����+�!�1/P�(��,�o@��9��#�p�(��*�?�+\'�G��X~�{T��ћI��Ҧ���
̫2-�cwt�U!OX,fi�D�F��H����k �!E��Gy�Sz�;�,�fN+GJ���>�R�ǫ����7��L�i|`�F�G4p�f��V/��h2Y��Q],��JK��3��1 ~�n����{̞��p��ah���	�ؚ�`�#q|.��q!�&��cɽ$�7k{�Q��]Ip���|���J�o|���~��r��׏%%�l�6�
�Ox�3
��6A��f�̩��v���f�0�N��Z��iW0\�t��U��L�q�1|��C1��z���{̕�B&ަw�R4j��ˋ�_��������4�wrmF� 9Xk��̈́}z��Q�}�݇�s[����^�p�æ/dQ��̔���*�~n�������$�6�o2�[��D�TC�z~��*�d6Q{���;;������+/�� Z������)���i"'�1wl��iB#&V�cK���GU�h���83�z��Zi˝�܍s����>5=0~��Ď��DB�i^9�4���q+�MJ�I�r�,��|K����g#=�l%OuHRI�����@vL~ɔl׫tJ�ִ�˩�����Na.C��r�� 78v��y�i�/�L��EOTX��T	ƈnA̬����:��{��p�ɤ���3_����zǜ����X핁gw$8b+��T*B�ұ��y�ʾFm{1V�dX��Y��L�\��+�;�eR���'�u8�Ԁ猂<����LO��'=�UlQ]�r�ԣ� 6�G�I�$�s�;SU�=(�s�s��͒:��U���I��<hY�����[c4A|E��s�uUj��1�����d�I+Yu�3�Y�'^��>�r���Ł2I�lXZi�!'أy�*���ng�������1�
��������Ν;r<_}��olt	բfz�c2m��-�ĳ��d��-������Y�S㵧ed��R�p��=�A�����c"
�g;yS��W�X�ĺ둴��H�	�Y�⣢��ϮFC��� ;v�ƇẨ_ƚ=�qǗ��$��ǧg]A�o
&���
4�Ӹ�x�Ԧ�q��S1=�
�Ҩ�pV�{pT����`�$, �����C�?�b�f��o=D�u2p�1,kb�)O�Y�b{���)?Ɋ�A�(	��������׉|�y��πA�;g�dg
<��n�S#�����B�վ	�݁/K�����a�o�����x|�^}G���3���N
#���*"Ģl�/6�\�m�#�赚���zO/�yWY~FC��� {2�{��ڭ3Jez봨b�ĞI뗸�#$M2%�����Ȉ{}��X©D�CC`(6���).��}�(ƅ�7���@`����W蔼�4���"'%� ������O�M�SX��a����!��4���CfU`N�M�Dk���XG��l���`���p�� mL[��2����.h�^���a.c�t�/b�]�8��E�����}+�M�~%UЗ£���i(d�A��O� 'մ��}��F�tU?6����Ɩ�s_!�CÅ2���:���)��i��֠��u��TxncN�Ӕ�>6h�?��oU�� �S���楄�帉2_�,��rt��Л���>ҏ��@�n_���N��&4�3���S=gw#�Q;�s]\����P]�h@�)d��j�ڢV���)c2t�*E�~�ۜ9h�p�W�˒��SL��O|^Ӹx4����/iE"ڦ����2�����j	�L�M�Y\Am��3[�X��B<ڶ��+(	r�oq����?���\��Ɣ��R�ՎI���衒�u�]r�������ڷ���Z0����a5����(������N�
�#�]9�*Y1Ԧ�X@p-��Lqǎ(m���F��,w����
I��=�V�U�k8�H��k<"���쉬<uԵ�/�I�KY�2!��o�S�O������/�:K�W_�;�q Q4����s�L�����0�kk���L�F��S�}>�T�WJ&H|����[�=c����e̥�F»L)&D����a�lE���:��pVg\)8C#t&��oDHD����;Jj�r�ďꯗvS'��)M��87�<��Su:�k��3�P�ʹ.��S���fD�=�q*�Ct���e��7���k� �P5�.����{�(������k�%��#��= -5M�����yV�7�`H�C����;����p�*+	��.� /�����u9���{ț����%�.�Q��)u�*u?�\f���"/�s=��Y��@�_̣$��E��Ă�BMR.a�%0�@|��R�i�������;u�9G��Go˕� �u6�_s�My|V}¬{�����T�@;��,m(v���ŕރ�b��
�ҁ�+e*
O�MY��
A��7��UC�B�
W�?�n<���ä[�)�z�NH�b���29��[�C� ��,w�ti&�cO�k��,����ݵ�˲�lP[ �kBԸ�?��BEdsx�&��q*~�	�
ĖYߒ����g�Ue��<slv���<��$Q}���q{�rQLu�Ǘ�P���>����2n��@2�S�c�´^ �}(���ǽx�z�䮰�2i�B�'�.��P�Tc3x/K_ư�\�6�{f���Q��{�MAn)�r���:%��h�r���e1��/�ea!9�Mw���:d�"v�������~Gb\�-"�L.���!%w���[�Jwj ��&;�����MH*x���(�⯮�H����	�D��s
��#\R�}������|�;�4=o@%Ӆ5�7�� 	.w ,���t{�#Z��N��X�C ���x�p�G�6����|�Ԑ�{��O�)��\&`os��buI�OȆ�Eq<(�u�;A #�ۿP2��g;<�z���$"��US�ĵ}Kgh�q���,;�%�w�����R��p��U�~ ��43τ1 ϯ�������N�Ms2��it��X�ILs?��\86&,��*��Uz%��v��&M`��*T�x&jG1HIs�O�N�^�ee����s�����:]:���W�0'd�$�
��)����*2�t��N�����ªス�z$�tz[��m�a����Zñ���o��$�Iu��j�<>И�_9�E*��w�pO�Y��=e](B�f;�e\PC/�L]�_��H�/a~�M�]��ƌ�l]v�IXh_:cL<�ɛ�OeȜ�U'^��j{lOR-���&�&��qgå�s�u�����H�|������ϕ%Hx��������A��s�l|U��4�íI���h��vKڏ6'T����$P��a_\��O�0���ﮗ���K����&0�(�U��;��.��A�9%����l�׫ k�����=�����G����0Ҽ���ື�z�P�G��Ed��"��l�1N����'Ǝ_�Ui2��p�6��9am�.�������dr�3�&K���T3'�% &�v��}�59�Y�,���uY���GY6i_o�nۈ3&�'�Y�1�oI�����V]�ה�E�LUّ���@ڗ�mŠAIkHu�r�y�c:G܍�tq����~z����vrm����\�Q�C�a�`��}BE�s�\���w�U�Ļh����/.@���܌&;���%gK�^��F��he:OE��#�!KXx�:�$���[Aڥ�/.�ZM,�
fXiB}��[:p^�uy7đJ�'����M�t�B4ZH!��s��% �M�ŉT��)��?@_{����V���BX�Eq�5�7��|!_6dr�[�M�e��?FТoA��iP��PZ����d�2�7���Bg�Sj�CFK�*�m~j"}�[ؑ@}�Y*�R�C#7)���j>J�:�F<W�ž:�����ۮ�~��k��f��3@���'!Η�Ȼ^n0pkѧ�i�_^do����wMZa�|�ߥG�M���8&�S�����v���$�����3E��~���xg�C �o��().���ۛkJ�2���C[:��W���Wc@��R�A�L������g��m=]P�q�($bD��]�b��3B�Z���Ǎ�fYEo��R௉	�5�͗[��ۨo8���vg|g���7pesAף�<���lNk��S��. mD��`�'d=D%d@�f��Ž�s�L��T;�t�P�wK�g'0$��x,��䲿y82�-<��dHCW����Z�=UI��9���νA�s&�����V8J��	���ڿQ���_3;aC0㉛���\6��bR�x����|Ua).u�2��|O�͉�8"EOV�(t��j�@���P~h�٤�j�f%�#���e�b~3� G�y�|^ O+�*���eDuc�m�7�'��hX�fà������9�Y��{u��p�eҾs�E�;vZ�\w�!!Y;���Z�N*�Ҽ�������. X��ˌ�m>��	d��4�?�`y^2-lArjaw�p���wJu��R��u�dc�e�!���Ɍ���ւ���Y$	^m{x�E����X�fos>:��ꐯ$ ���5�e��A߁�}��ַ@4kQ�K?/�4w����m�c�l��C���$�T��gy��	N��[37J'J.q�,K����Z}`P� I15�N�w����퓈�o͒"�`-{�*Y�p-">�e'N����8��1��M�f����_I!}���k쬺�0Q������w��B;���/ʁG����_�"V�=>4�׻I|�윑\6Ќ�1t(2��7؅R%��m�<���D�L4�-�6���m�&�Ӎ���/�0��b��Y���s��N,R�� -O��f6��#py�ڵ��?�g%�����rΎ۰Zfa�xE�a��k����M�2G��=�;x�w� �ӢG7�Zqc�i?`���C�G�D�T;3�^-)��[o����!��o�W!��Vz ����wig6.�ݯ9���b�a�F��6������`s��+g ���m['.����S�oJ�u�e'�,x&D]\�nʡ�@�-���W�s��+6��}��W�d���j1'����+��'�3�#�B;#`-	���ĥ�TNE�ft{b���)iV�QN�9�������
*�� ϶����c.��K!�d�ٟ^��ϝ���ͬ��dê��_��>��r���1hwN,�>E+�}�jf�K�Oi��Ӷ݉�R��8]�į$���J�8S�2��R��]c:�&�r:��}���,��7+e�V�jy�ɾ/3�B��_[&����j��i����m�[�Tv�t�T�kG��.3Ѩ�G�c?��e�����4�^I+2GW���8�ҕY�4&���r��`wV	�+��4��v��h&��4�D�:� �ڰK
��0��H��2�9ax�U�`t_��J�����½q"]�Sb�O\d�N�yI��n�bգphL��	�5_H����7�6�u�k�f�OX�>;)#����>�ڜ`�w����CCI
6.x�ͤk�6�&�Do/��)��U$yjp�
���-�>��B8'�5^���F:.�2�I6�<?�Rhs���]���x�_X������9�h������]������A|�sh���2�4N3vz��$#�z^�l$'�T�6P��e	&xl���on�ag��x.������-��	��s��-a*��ѺR��{*�ׇ��r����TS;� ��_�`-�� �v�F?��qzk�Mk��G!v,�ir���*/�����|.6��\�T9x�H��B�?�VK)�X��r6-��4���
�����p�7��h+J%d�N=T�1c)��S_�s�L����NJw��L��N���%l�^m�ղ�E���s��j�!��q���H{F-�A�ȣ�1���ʘ<���C���:�0~?| ���܆n�`���+�5����$�>���/G(;�o��9`�ͬ�7{�Χr�x-�ȼ��$�JC�ҫ�8��U���p�%�`��`>��*$*]O�ҭ�2Q�eb�b WFږ0�I����?=�F86��p0��+>5���^I���4r��G�bڃ2��;��S���*	{�?�\�WpDbnn�\j�v�42�ؔ�th8�@V�H6�X��a�A��f���>�w�c�·s�B���[�/HIfw��6g��:͹I���=:�~s� ��6�Y��숒��<�jFj��,�ĸ�d�!ƐH�E��=�]"�u�n�Ɓ�fΚn�.�xN��Q�� y��0�1?d��FZ������UҐV�E�%�#>&�s^�-��}O�*��Tc��\*\ȉvU`'���&�ȪI��82f��b|��	����hb�2�":R�{�7o>-��L[iVM��Nl#lp+wn��Ť3���w{ğ��P^�i�����oq'�&W(H������Xx�	���DyP�}P���}i2d0(A-S�� ��X�Z�r���:��e�����p~d�N���l�#퇭�c�g2.R-�fM4?Wq]G�s<�� v:�A8����,�0P��zq5=XX�I~ϣ��>�=��伒w���&,����͗U~935=� �Mo�
���}�(x����!e�K#��٪��UTP�r�D�B���a�E�^F4ɫ!� �����	
�#���y���4���f�f�x��ʬ.�|N�j[�c�|�l �Qj����;�����-��P������RA{����h��ƒ��
�	�������z��>�25mY�I�|�T�D�}��^
�}Y�c+�<���U#���6�M5���_H�YUd)1�CJ�����+�h�G�����D�ٿ&�|�����y��8g9gk�HTd67cF�$O��z���'Wŉ��=95ߟ�k��;���G��~o�\����Gx���>f�5<^��#�{�,J�������eQV����Ŷ����Ӆ�$'T�W���rug�	R}�>��OYF�����.	/�y��/��شS>�ڿC����[6�萄�v�ڿ��U�=����EZd��A��c۹>f�Y�CQ<��i71�ȇ���U��X~�Պ#e�+��{���;k�Ô�D�f�8��'ò����#E3�Z���+<�h�9X��)�p4�+� FX�e����&��X�/���cJ��5%]�7@#ϙ��CnT7�9�E�?�ĸLU	���?�`�����)X{�}��5ya]�֕���5q����>�:3JY�l��*lQ��D�l�(r���p���8O�P��)��f���6��?۽4M+�C����[
�t�e�iw�!���&�!�1���s/��.��c����-#�����m.�<���>��$�$�V��*sn{�RrIR!�&�^0�'{��Ǔ���N�֡�y�8���҉d�L���_���v�A��N�C������B�7la�gS�~��VG0F&��Tv�X|b��⇲��q�Q"��j������ |��d�?<�STC%�ټ<���9���,���_ң_�?I��<�0kV�8S[�Zd�R��7�����)կG;����yϩ*{Hчֽ�F`1/ \��a���� ���S��NO�w��Dq�9�N𰅪�t���eQU�@�-����bŅ�-�V[q�,p�HU�w��.Ni�#��Y�O���0����B	r5��qU9�ˡڼ�+�6��Tq݀u�H�J��/3�%�J
�"l��1��O��&�%��<��0t�T����������:�&:�c4W���X���p�2�o_� �U��[�A�/n�1Qڱ.'D����	�CZ�ʿ������
�7_�7W����a~?�J���s�+~j��:}}���x1X�j�X���
T �k�0Z����@lj��e�T +�7~W=��į$)�K�1D����� 1�tu@��������,|�RKP{�̌0��4��p��?�-5�#j-��a]�J�x^�_�v���7C�B5���#�u����0
��W[�ۤ]C ��辦�Efl+�ԛ��� �/��I(��:#��R��Oe�]p�O:�V�=�0%�ۧ(��;��'U�_؋��7!c�E�PiM�Ka��{^� �F����$�ac����bX�}v�{>��M��5 v�ˤ���_w-e��ca�)����QVa�Nʃ�
3iyl;d�1�.f��E�a�x'�9�L�$���ii���B�D9�I�s�wN��!�hX�Pm)�!�?�-Bya}�z��iF�Gr]��ku��q��������@>�RD"*���pڱ��Q4��]����2_X�m�F�,ܬ�����b� @��E ��\n}a�ɩ�S��\�;yy��6�PвS��I�H%l �a�Tc�����f�Z����1�b�DS�d����m�G�[����h�k���:V������� ���Vx�[{h@d"Q�I������
e�{EW��U`��`�C@S���ǔf�w .�g��B^��t˾z�Ļ��I:g�E�w:L�ߵ�̧e;�N��q+���=�������x����	S�^�xl���\44>
jV$�1����s�q-�%�*�b������a��S��B Z+f�p�H�|t��f�0�uV���A�pNqD0���F��r>�,�g���uǣ!J*��6�>���T�n��E���Ǡ7�t&e�����e�Lq	���@���=D��x�0�G�k����j(���9�����H�؞/�_n������4_�����X�)7הq>x�EY2�\D�5�$>��GM�c�$DZ�:jXO�y<�W>jݽsr�L���r����4�w��F�M��ݳ/��Sc䨨$��ї��S~�${$��(�8���E��lg����u��V4h͝@9��|��/��5x�K��j)y�Ab��Ҟ�n'���N�����
����y�#��-�l;'Z��ދ��k�[�tX[�	q��o�V��ӂ¤��ec.gt��dK+�@��,%�a���3,��~��W�Pmd���4F.�����v��a�aD��C.��%껵������@���I�%�H�ng��P�O���zn�g���:�[��״�z@� ��[{��*����������Ռ�#b��D�K�I��ҁG�?�f��� �e�*�	�z�K�J�3�	wE��0HbF�c�K[Qv:��1�K�׬��8�B]�Kgb"�U�|e��<m���n�5Un��<�}^�3��&,���|jI8�_�`�I_�6כ׫!޻/�����:C��>�O�jS�h��D��	#硠��V~|�|�.�t:�¬A�&�L^��A 0)��I��7��>7�����5<3p����Q0�H�9~xpwx��h	^��,2�{P�\-����R�X�dK��6{c��<���<��}-�4��`���/\���i�
��l��|�!�7ڻ8��ߐ5 ���� !����<����0}�-�&ʳJ(>xBע��=�����S
�GPN~Է��Z}������ �+������ ��X��!�G���$���.6JG ������?���5v>2���ּa2�>U�-YJ+�.z���9��$(�(d(���]cx|3U��h�B�I�&�8�i��8�yR�*g6,yqE�������}�^^�h�N2���yA�ܐBDR1�d�|Br�<�T{�c�Ϗ�t�Y�v�K��D��k�%?c��!���臲�wV����E���$C�`��j����Z��O�@�6�뚡��7�J��6
�A����*v�(���b�sۏ'�v���c�؈��?�y\�l�C'!�LE%�.�Kۅ�o��ihE}L���B��jN��x$������$=�Qi��8d��"}���-X9F�Iզĵָn^��{���]�r�좎H�����Ϳ�8ni8�ç�18Ijh��s�L}}�^�25��|���,��Y���n�d<�� .�c(���q��w�� ��J�<5�=/f��m��z�yI1_Ȅ\�H�A���	#�]�2�
�\��3�;&4�X(.\�>���G�oG uL��P�M�VS�k�E����eƈ>t4l�t3��~o��,@2\y��1�`׼r�DRb�5 �4�wh�����f���)j,�JRv��mVqfJ7�@���x����9���F\��e'3A"�`��sCM��u�����/�r^b�����A�JB�'u�u��.V�h4���۴�A�\�?!�� B"�ϲ�F��� o�C�b8�0GR1X��uVuG���q�p��_�~��>* }�d�����~��:�KMEG��i����6¤-��?���n��#��~�MR�=v������$ Z��{���[H���^��&�ÏS]�5�CW�)�zc@�5���1�������[�I�e��v��fL�~���Xr��R�tm������yLs�/E>8�6ڂ�4��]�p;:�= -���bO���j��"�BN7(ܧ����氷�6U	
FS��]Z��'7������r�w��.kr����n�4�'���s��ʉ�2�� �f��Չ�
�:��2���8��BԼ<Ǎln���
%���z0�$5�U>N=&� *��R�Tv"�����&���n|u��7���C����ڸű���S	�zZ3)#�z2po���l���Ρ�/�H�@k����N�t�S�s�g��S���m��S#H���CWf&@����N��#,�=�p�K�f9P�P}��d��XV4~�*��`��ǎ��o������p!H��n��#�N5��ox�J���E�hW�����j��Jo��U��E$��=V�!���;�L�Ɵ�j/�$Ҫ�O�b̲|X�]�G�υ2����(��F)'�6�0�n���x�C���)�+}V�����bZۖx�v�/�g�,��v�ݜKB��y���R�=@�tI"+@{�X
k�3m�V�8i:~y�0Is,|���uGZ@)ye�]�\���&��V�{��
�Ҝݦ��e�[�ba�)PԖ��S7��I�<PDcyx�Z��>�+�Rz�}DT}H�E!���/����L�g,��痐�Wa�akݥ���� ��U��� ���%P��*<�s��;���W�hh�m���f� A�c��J��صa\��G�����p��nM�Z4ؼU�ٮ��	벡�|����K�M�Q�o�7�Y#�I�áD����3�Iߛ�Ą8��f��89�;5t��`͊M�5t�wo�"�s��Qy�NW�a�<JI/-U�:$U^��H��h-���D,�m5��e"ovI�K~MK�#��I��B[f��c@`%�h"p](�=lX�2�[��G?� O�H��f��T��
��ձ�2�M��n����%-�� ��B1�~�y�C[�ywk�
�?c��'�4c��'�d0���f���3�@@�*�IO$��/W��$��2�A��R���7���]d���Z���|z��zc}�I�U�HI��"UQU���G>�ѽ�}��� ���=�5%W>�e�Zѡ�i�����7�� d"�<8�X��V4��闗j�}�F$W�>#��d����hDdc��&,�"���ڡ�ت��a$�h�_�&H=��t��CAF�cȏ��9u"�\�F��-�����5KgJ�e"F�u ���1Yb��.������	5=�����_��q��إ��f@������D7B�I��p�G��&���B�7�h��9eB0	��X�#�΄EP�p�����M��/>�AKw~�"��F�� �z�2뿶��0b�^?v�\�c�޼���O�7i�%��)�~Gt�I������P�b�Շ��~�h����	gm'e�W�m�s�3�Q�tQ����C�yS+��NO����l��7��G�_`����: h���#��^�d���BSF96#4x��vc�i���8��q!<e)h�p�,ؠ5��&;њ@�ށu�N������}��%Q�:�� �zs��â𺵌�Y�/gn�^Q~�������?v
@�?�u����B깎U�1	F,��m)A�R4�(����!� 0(�ڴG>'PvH�ap����qS@�|�ϭ*�l��xq���k�l���do����Z�v�N�J��TDO�g��-}!^�VYk�k�eq[���fI`Eel�ud�-�F^HH-1q�͵H+	Pox���+%W�
����q�����8���#�����]�d�l1�
�]fd�s{c�G#�y�ߙsbp&��ಾ�r�55�W��R��f|��i�W���ksLK����FIc���2���������Qd)p�m9�/-�U$ǀN/Xh��_�C��S�F��s:ht��0���&#1.�W��`)��?��E5�V�"m�1�X����UG���8_d�N7�e/�f�`v
�Ϋ�sK�%�	Ň���l�����q�<�?�U�W)y?�nPB��;�#8��g}X�	�|�n� ��a��P8B����w(�Y��Ӿ}܅�D�����K!W�.hU�XR��ڿ>�C�-�X�!���!@���Ё˩����5z��3��Y�JU�~==�w.5�V�G�NO���\�!�F�,=�(�
��MH+2j7�q(|�-�\�0L�>0��4Cl@��8ѥCL+�h!h{�a�0��#Yt���d���Ƥ6��� 
���$~*PO������	��2��J¬�:]&@������,�y�D��?}tG����8\�u�@ �u�?G�-u��"�9c�ˢ��iE�1*���{��ms��[+�k-�����E )L9�g��ħ]�} �¹�P )�L꩘������y�p���}�P�3��O�P������_� ?Gl£���/z��6����É��2�]��2��cN���4�t;F=.��M�C�4(w�ͱǅ��:�IF������*g3�"��Sa�X�SRJY��%��|��ƨ��*���%޵@q3)2�cQ��#ˡ�E����s�����I%֋�c;e$���g�|'�蕹ҷ�!�'4�A��q��~e� (w��U�/B���wq����'Mc#�̔���V���Q�=ætQ9�e9?����et��>�9��HC�z
Φ���󥢄�بLs��<ޮ��;��/_8�k_>�Ϭ��W���p�ѿh��I��֗�p�*�+�S(&D�Ym�G������'r{;9�a�$=�p�%����^n� )����2h�[X ^O!ENAN��$1El��y�E�!H
a��B����(L�0�D�v� sV�ƚJQa���������x؈P�@�!lw�2���t[ԍ�vp�h�x���_�jU������M��;_�7% |Z�ǊQ���ܬ�P��P���dX����X�"�����NB"@�Q�*�u��J��+EoO��Y��|�s�4��G*����Q�5����~m����C�A��'a�{h�~�X�FNe!��=Id��=W"{&������O+n�+M���z�mƛq�	H]��ЈL9��d� ���/2�}�ĚR�-��0fu�!�	bc�G$�j �H;N[fU2㹕�1��8����� .�7�$����D�F�㕜 ���Ý2q�sI�`�-�0{��X�1,I@�F�Ł8��盙����b��d�aml).`)u�vY�$;3v�bp����RZez^L�jC}ƽ_g�8ϚT��2%�D�&D��mL���I�[u=�3Ԩ��2#)m��i�Ijʕ�L��qa� 2�kp�q��H�Zc���&6b�vt�)������4�C�8D����E�Ʊz�	�FC�i���� �	E�Z���&b��D��mJ�H���1X/\#d�(C밂�=�L�@���2>7�v^z�2�fO�t���V��ͧ��qi���9����È�� �uV`�;M	��p�;�� k����sac�̳�_u�$̧�_'�Y�9#��v���:!@t>��$ί��Z�J*z�)����/ߝמp��1&�l@��n��s�0!Ҷux"I|�T�i<t1 !����0�U|%���(� @m�å���t9v�	�v	i��=��j�hv�>����SYX������W2����^�\���+l�ks^U��I���ZD7	8�X������q�/Y`pu@j�ޙ�u��:%3�T�ۦ�]-X�gh$�h4�n�R�\�+K�~��KA�����Ȑ^���ע��[�!&#CqK;;�Fӱ�T9�R�!	��^}��y^�"�`V��E����zZ�|#$����\j�
�kkK��<�l]#Y3��ZY15�8������f�����Rя|^?v��or��8�_�H[�E��9��n{�7c�^�6��%w�Je�eVr�`՚���ߣ"Œ�c����\I��V�E�&Ug5'=5�{TnnxdQ��H�-.�Es��g�;.��~��p�C�^+o^rƻ�#�� �q�M�П�����j�ت���d���5�Ԟ;:�%7X� ��Q�&-��1@V��
Mi�����__��x��)�E�.s��H�U����eC9Q��݉p�_TR��Ͻ�e�z&�[��|���׬������N.� B���;0�S�s��Vi�9eo�����^8/LЛ�6yw�.3�)*`��._��YN@r��	�`�Fa����% �P�
�`�9�]�MX4w }���(/Q�/�N��%���V�xf]T4/�K~��CG�/��\l�0/��k�²-�qF�&A����P��
�o���k���7��@�|�>0��ޠ�ų����w�L����ѵ��}�o�(�y�2q.�Y�[�1y�΍'˒S2��Py� ~�F����L*&<Z����m��[��t�C��U�.�	ސ�~���|hE-ɹ��Jx)�s�KU��C�A�)���r�(g��+^R[�cό@�y�D�4B��H��2�(���s輪Mv�����+�^�-
8��)���X�'5&�BePNlqaQEG6���o|.��n�v6�*'j��1��_5T����Ut&D���A@�/�I����,k\�{���T��N����Xd�~Q$�~M��e�B@��u���!pa���O����P����"�K�#X�0n�@�>f��+��_��'��Dݸ.������>Δ�R�*-�R�7�������{����p}{Ͳ.�T�d�O"��8�v��(/:k:�p�����ޮ�lا�xa��<�WiO��L�8���s�פ�D�_�z���_�6��vQ��E�Qޠ��]�⊅n��o�̛:���/j�>�p��'h����<�2Q�4_�j��"�u݀o�{�ϡ�0�n�q۳�Դ"�^Y#C��L�z1j������(��]����lC����/�e/ը+�(���	'��Z��owY��\�0����W�5��ݟ䣪�'��!���?�/����&��x��Ԓ���\f �-pb�=$2/���K���3jG���5(�%9,�ɩ��Vǡw��U};�_oc�ę̽���J��݈/ے�SJQ�8r�gx	ɠ/��7%?_Gt?{5 ���X.}�$kK<&r���it��-�s!"�����.7�c�����h���=g����R>��V+�<I��J��	8	��]\l�bu#���ޫ7:�*ʝ�y��B ���W�)Nb���'�?5����_a7��h���$�Ͻ��2]��/��jBsI85\T+/i�����j���!�� �}��}�,������y8�����^<ʒN:�m��|��0a���Q�ɖ�(�u���S��$XM�Z�}ͤ�3xdG�If���^�$�'�Y )��Il�Pg� �ս�>c�4�f�h�M����V�;[j~�t��m�����Y� ���R�A�0Ȫj	��R�mn��K�4N+j�F��y��H�O�(�ė��wu���2|�G�8�8i&&��+�&po�K��+��ٝgA�f՟]�[ ��$�"�㫞FJe��m��_zˇ�Z��R�.�Cq��Z4���S./v��GfHoc��И�/��ظ�K�28�����rķ.�\,ٕ�s٬&|&�5Z�VI����y}^� �𵞵J����G�ń�����L����y�W�8>0G�"D��[D`LD�,S���� P��/\�w~~���;h��g2�f!3У�^=�0����s����=�� /�*>$ņĜ��I�C����:���Yj�Q�����wn ��J:�o�<mWLaoco��o�����Zv -`��aMb���_	=<�5�4_���!��dq��'����w�qK���U��f[�]p	&}XX-�b>	�K
����-��r��,�I��@���z���^�9m��&S)$�&o�2D��GK�R���v�d�����p�Xf}/�����gm��n��6���fy�R�����Ç�%���j��e�Y�C��?�v"J�D�����b�BZ�﹣Y��]%�/��*��0�K����N�uO������=�����[dnd���I���l]ph)�Ԝ4���JSQ��B����d1������_���������ۋ�Wƞ-`Z5^7��۳Q�"�i�@��`�qN��BQb����	*���Q�V���֏�X�q����h�Ի�@'C�i_/*Ƕf�*sv�&(���|��_��쵋_f催����$'�����e!J�>_j6`te"��k����7XST����7�����{	Ŷ�\��G(GP{L1Ua��-�Ħi��ɛ���a޴�m�Ԟ^���z�L[?*z`@np�Y�(�;Bj�n����4	?���������J�P֥ou���	�ѭ6�r��]S䌣�p&� v��L��]��{��g�᧓��.����F��m�vW������{����8���3ۄ�T�F[6�F����;nO������Ezt|�)�O��6uE��+�@���#`�Z�S�3��~O��>9��R�����t�*i8i�yҾ%�v��>e�,#쿽��;ͣ�GQ�$��sh�O���&�f�����n�Ej;	�7S"�9�֑�W;�P -�Y���V�!�VHx�ľ-���i�_L���O���C]g��N���69N<i h�{�X�{܌����?�A<�x�8�hw�΍w���ft�F[�dn�����
q�Z{��Qa+6@�M^�d&��{P���z�
�**X�SRņL�W\b�G�pv�*�{n��A�3�
�{��܅�c'e���Z_B�7�v&$�+YI�Q���6�o�+��9R�����<�$�z�ƾ�����ڀ��g� �������9;*�reƑ6)��S�~��7���T��wkL���&2�3��U�K�FE��B*xS�K@k�G&�����X�$qS5�K���l��!�[��[o&��R�7���m���hВ��D�ur:���ߒl�Õ�+��2��?k�
I��Ttd�Q��s�Fde�j�T��N�^����-{����]��cu<������sPV�me�s��u5�s!#c��@B�-�
�O���wev�!V$����y��;<S��,+DҌ5&�cӂ�_Ξ����Y��Tn:���R$1� *5��K3��*i��g36�{���Jp`���"�̀w���MaN�ű��3��y�����>o�l^>��c!�.t !>�`fa�>�8y�윷��}O�hߕP7k��AqE3��=��D{��������ƼQS�|�Y����1$����������G��|��-�SP0yP~:W*M���F�\�\|n/�3QP��F��-���v����4i@��'�G>'�2S1��#R<pH�������܃!�F��� ����_��hk��|QzH���V��'���N�}v�H�G�SӪ�IRՎ�۩�{�y������/��T�,�B����>�p�[�]�dmu;M��Jp\�/�@�׊`o�摎[��`��	MR�J�vE�i����2K+z���>�ݹ��� ����]Ǜ��'�"����S�.��<��S�z���
�8���:Q"�+S�7m�5�%Qu�7�:�m؄kX��*�ݕ�o7t����B��½��ۆ�ͺ�FYfG<�l u�����9'_�{ �;{���@f����r�
�f9�np�M�.�r�`��}T���8�ʸu�G6!�s����Jۆ�g{�+9%�Eϵ�������E�b����{��
#Լ��l�S�����-y�ŏ�̧6�W�˦�/�[툊�SM����՝Y)��g�����/M�!sP����D�~l^�'�0L��w����NB�j!�U�~@mdQ�
F����/ܽ5
�Z��;wEӁ�`0۬v�ݨ���#ʑ�a5�0��:�X��Gь����=�K���M�K� A
qc:��������0y�L�eN#~9���,՘��>P^�7�������!� mg�O���B8�>��W�����BʣE���PãlWxF}*RE���'n��Cn{^�Ě��;!����ڈ��M�&��]SLh=���]���§����Kb�o>�r�� ��������I�B���B%bo��]���WE�K
�FdVnϏTh����h�)?qh��w.c���O38|�'��B5�����Qs�"����RM�1-.��`.��R>���&�z�I)�:��R(4��j��`��Ch�>؞��R�����ck�IfÒ�?y{:�F�����T�|a� ��w[S���6�ܹ)�+��G���n}[�ԅb�v��f��7�ww����ml"t�fw�P�n���� ��$�S�g�g�:2��{co���a�T��"�#���c	z�I�(El4a\W�vܛIO&ų���a��z�ߑ�G��}	|f�{�{�$x/��7ꗼ�<��|;�o�v4	@�*#;��x^\Lu$Wo�z!變�Vvf�}���qĕ8 .f��<�����sȕ&iPu��S��T�J9��z��DҪ�D`?��c�J:O�a�g���>���xI�=R)����Ȥ�^]�0�zak)��4�\ :3E��*L/�_D��g�fߏ,�r~���gp�`ڋQjϽ(�ObT��Ϟ�Z�5C�/�Ig��.��:�w*P�7e�}�c�E�hc��ENNä�z��Ink~���ճ�ӳG��穊�<w/[�\
����h�)�ߏ����A-��*�5��A��T^�巍e�������z[=#Ì��^��(?�ʭ�s��;TqC�����>��>���	�""��N�:��al8��DMz24�������b;��ypP�'�BK+��jq�B0B��(��i��s�����ч�h�@f��C���X}\��}�'��$=��sg{��=�1��#o�z�DS�M��TEٔ�Y�6YTʁj$P}ŦZ���"�D���=ߣ��d0�=}�N`4�]���O�m'��^�V��o�@��9ҝl�c�f`E�=��ig�8�8L���c�Aҭ��
������8 ����yG���P@� ��ʬ���9��������8���G�@�$z�Ϛv͈ؓ�{��]�ϻ�Q���(�0MP	|����?n9��2�z��i�)��b�ϸF~-$�������H#�{�]}N�js!�S�58a��p$C��6���|�Ո�I{��"2ߣ��ޅ	��ti�+P9�c��Y
���7����4�z
1�E�����}i�e��g�0B�"�H�,�����z=��v��M�b���f
�y�A��^R�iRe������3�D:|�	-�1<��d}�h��� �E�v�C���7*�P���髖9v�.u5WI��T�-5{q����=jF,�����n�eH�0Qol��yN��J�������Ss�[p�V�sfH���j�_�.b�=jLr��y]O}�� :�K�o �X͝�<'�9L����6\p���.u.���l�+��r�:�L�Gvhs�[�c8�n��T[l��X�7I�l�T�]͋�d3PP�-
��ҧD���7�^��8�I����b���_����Ѿޛ�p2���x�ff�J���9Ց}�DTaRl���a��&a�A�S�խ.��/t�*	s�F�wʙ��Y�y�Ld.$U"�z%-���,���#��kHG���c�n�Q-稸_�8�G�\y�&�L���_i �H�D��߫�q�kY.:�,W�V�C�^ra�ߢ�rn�/<9{89���	Z�E�d�ћ���$�x�w$Q�;����o�XǨ#�}	�x�@�s���1��m�+'6D>�5�tQ���6<�s��C�\�5�o�/*:�İ�c��|��/눶T�c���N҂.�
�9}M-�7���1�ֆj�-a��g�m�����&�*���}B��M����iq�
��\��I��	w�vr�(��'�ꅬt쑲�5�φq��F��y�D��/�(�j�x\
VG��c�����*����&�P�ޫJ\�Q���$�)�d�|�=ι�-˄bl;�|� �\ܐr�`�1�k���#��QF��DԨ�pj#Kl���'әZ�N�˼�s��r�9�vPB�&nbt��?�8n/#Zq�a�f�O!Qg��~]X�!�3(��Ϧ1���,lƽ>�G�o\RK�wD���U�Q���2��XP�����9i'��]��M��5�O�6�k)S����ؼ�}�~q6�F?�r�W(�5�h���@d�j*S�7Ό�S�����zIfh�t��4��:>	�X'��i��5�.��Z=$��M�} ���^EӮ�d��� ��6D��01F{!.� �	�&ei�f���kK/I��h�ض��oc�&VT��3|��~=s�:�ݓ��I��W�|u��KA��{��z�8�{ȸ��d2���IR/ux4m]�����z�%�m�lR0_�W@/L��y���ԀV�����0@�";Y�jbBvyG���O���|+(b_�<�aތ<8�H�ֹ�z�Z����*�F��x���YPX���M����$G�t�}�A���Ե�p��m�W�oӁ�:"ki����:㋕�}���N�0�C�b+�2��)8\Ku:q_'m��m��R!q��H��͍�{g���z
���i[��E�l���PYM�w�ȶ����c�1o\e�ݱ[�o��+�#A E�����v�t�����kqyr��:C������G� �/z���Ӆչ<j�>�;��� ��L���a�T�����j,L�@���"�s_*�]*����Xc��F @d���`xa*� o�`+�a�s��p����%��҂����1Gxg*%���b�]�U����c�1b�$���Lq��	��l����'i��1��Ar���*|�P���fO;v��JG�&��3-�	M���D��O�� �dPO�U�S�1!���
[�B륰ܽ�}YCav @g�)��tH�B8&O�e�2�%�x`�����F�0��o�疕U;�W�@ �}s�ڷW�F�K�qs)/�Ĩ�,-��c���4d�{6\��r�>	�m��l��F�pc��_Y��X�k���wV6[0m��O���ؘi�a��\��1iF�Kڹ$8�U&R�:^�Q�ӝ�J�$��P��|����%�Pp�}=q�ǔ����;D�!Kशj��H�Y�d�;F��w���ߟ��L��p�ƹK���F���݉�[�gC�Ý�H����9���V��������a������y�V��ݘ��5�3;P�:��-�#��T��?�%]�l���z�S�)ʹĸ�Z�
�욖��.ab<N�E1M/�YzGSk0�\ƕ�1���IL�1$�W;w��M�ǁS�G����->/
����"(9 �����Z����a0nN�ED
@�HS-�9���p̈́�!z�g
M��k���]8s�&�?��׮�#O"���Fￛ�"�����B�cV-��"Q�8,Yl�)���@�W��"�u���F��֖u����J���c������X9 �9�>��d�E��Ff�%��Y\҇�%�WD�1r����2��X
�N�N�ЏtV�=p����9��S���q����옏"�c7�P]��f����/	��H�7U�hH�1��%��2�US��+B��^p�a �#����V+��}/�*�/���:�ݒ�S�k(�w�H�@7~���.b��1�.��Ɵ/2����.o�ms�l@��K1�G p��E����n&�������Fq],���Z�㱄���3�*��IiV8N$��µ�s
�6����^��_�,�e87|�ri���(?�.录�L�>�=�T���z�D�	@+�+�8]��1���D�1{�n.�ӉdG�s��&��|�E˶jast���ܐ�V����I���ь+z�����&x�.+���p�ZD���Qi~JPpM���T�XF�
}���w/D���կ��:|���v�L�"krF����0��mZ�{;S������i�A���uDۿ+�j-�m~�4���F�������H��
�I���C,>գ�Х��-����b���Wa0."�@�hߨd?#��N�����>9���N	=�8������u���?�@"jT<~St
��!��K<̿0�����i��~ �[(��	�T�� �n2�'B�(��قB�J�T1�+�V��ͨ��j^��V�e�ʆP��n
x$u�n����K�ia���1~�R"�\��7����6�#�\I�G�=XV3-8Y���P�T�/^��9�=:e�T0$�qI��U�+<[��'4$��M|3>����i�pg"[&h|b�;�e�ht�jI�?b���-l��PJ��3)�~�Y�[!�3��BX�����\�gL�iss�R����`Y�da%���������,�`�ȼ���zE�����ά�"CÐw"g��"���v����T�V�|8U��C����p���jR�(-'��j<2bn�<����LL�{�� �e��O�0��y_"�ɒ�_�C�y)%���a7��wW|^T9���-婽��1�w<����5�,� � Ch���\�53��Is����#q{1J���+I�a�"��Y���'�,�M�Ժ�Y=��� 4�i���o�&jFqJ>��"}4yx2��"ߪ�7JO6���v��R�S�~���2>�)��	�R��
�	Op����2���㓌��c��=F�
Z�2��|g{-"Y���<�D�k�S��\�*i�^�O(�03�m)��I�?_�X��e��f/xSqԛ�M����JF9�[ S��]�᫖��6��j�d�eZw��'hȽ}�w�m޻4x�5M"��٨��ҟa(ܔAI}M��!��T���kQ̬�(i\j�K�W��Ji"����
w%��Ň���oW�$k�
f��u�v��_ ��9��Kc�>P�p�6��4���W�C3yݍϒQ��ss#:���Y㴯w�C\�;��5I��1�4�{�ɉ����� r�S�{�>�_��]p��L�ː�[&*�UD�$��ͷxI���p��p�䟐?���H��@�Иж??c~*V�)F-Ng�3�&�O�)�]�-�o`�&�fe;kK^w�t� ��L.ŽᦲhC�"����-�&��*#�:�]�v�y̋�ob����l
SK�"y;6�)b��wX��r�uE�k{p�h�� bY-ò5}�B��k�ę<���s�萎^󷣰E4��������>���,Sd=���\<+���I��8���3�{Z�0*�v#���'��ȨK���ǵ�&8j��/�[#׮��7+D_�zP0r6O��`�7�]:T�#Bؠ �$de�s��{ii;m�h�Y�P�8wv|	�L�ӽ�r�cDS{�~%����m�%"AP�Cݮ�kLU�Aد��c�^����9Q�v䛗Z��6씡&�n%� g��Q+�=�-�C�}6���������0��ǽ�	�1y��E�6�4�Lb���$��4����˜���7%��;O�TlO��� ą�g��Kx�|8�k��`~�D����!�_�)挏�u�B���bo��FI�0�(�=���e8<��`�6�'���� !��J9��<b�,����g5�dzR15.s��ȉ��ۘU�� 7OYk�'jn��"_�#oݫ]���}Dc�j���,;��~���K+�H��{���1A) �$@󩼨�#k7(.��,���xqU��vj���o�HzB!�H~��_*g{��V+��@�(~����DH�|�4�ŧo����P+�G-��
E��n��\{^�n�_/�^�\M+SQd~dK�lw��hǩv��>4�u#6�KZ�]��A�wH�R�H�ޓ":Ñ��h
r]�N�qke��E�
�Z|�#ŚG�N��я��H���DzU&hJ����bsY�n�Q��hs�(=�l�����%��̀Xj@�b�u����+0%Ԫxô1nj����_-�2�����i��ðF#���;��� 2,K��#s��
X�
�L�Q��º�@�p��V*Zҝ��K
����q9_��{|� 
J�#[%F��g�P��!2��Db*������"�?IʷV��^�v�DH8��R߂7ٝn��D$8��-՗\l�<���(�%1��{%7y����w�=���{����F	�q
k�D�x����F����L��-��L��h+��R�,��aP%>�$k� 1p�#�e��͞��X�M�Q]K��xl糵�h]QK�r�a�qQ^3C^�ʉ@msCa_u�Y��;��9Y���v_<��]~ W*��H1�`9'�Ы$*wI�L�vU�@x�u/�yb�N{o�����WE�k��U��G���F����w�A|�d�1V1��'��"��>L[�dPY�r�`f�q���Y������Bl��b��a�(����>���=�Z��5`)�',��ަ��#��I0�������Pӟ{�hI� vh4���\J 6�)9�
�f�&:��#ۡ֕�Dm_�0[&Ӡ��F
z4�p>�qt����{��.IDv�D��8?�G���-�.��*~���IW��opG����BΛ������"'��qj.վ��?��"�C�*��Bj)�(���s�cƙ��hH�qRY��z��A������Ef6��_K�0Q����sp#4��t=1�dg��h�`u6��Y��v��	�L�X�k�A}Ә-�<�Z�Z�RO�C��Z�%�e�h@�F������f�[C��=�!'��P���ڇ,Fu~�mlxĂ
�#ߥ+��3�	�N�wmm ������S2�b��@E�%O�=u<D�pM�[��)A���l��و��t��u��<��g �֞ۧ��T�?�M�C4�f�2���}�Ccn���Z���"�R�-�s��Ї�n����q�ۥ�'	���*��sP�^��3��s,����(�OVq]̾�}r���Oķ�_M[�t<+E����^�xNB��,̔�
y�v���I�����f���΅I�S�d�8 ��9�0�>�oPYw?K�mVRV�������d�|4����c@"�Hj9HՕre�#N9b��B��cj��p�
>�ئ8�,+�%,ߪ(��gl�ӻ�	�BY���1qUM�ΘL����z��#��tV��(8Z>�O���+��>��z�J���	!P�l��+�Nm�	Vl�wn��n�	b��ތ����x���^��"ߞ���Ŷ�R
,�#	��^�����+�a�>�nV*���x@쩄zv�2N����r�0="�����@�6��B��qG����!�a��oO���Ђb=��v��L_�%�����2d�CX�9_�Z#gZҫ��_��4�b|.�c}ч�xXE��fwO����3sS���(�j_}�?�r����]��y���2�E�4,��B���U�D��hv����yJ�y4yU��5l0��&�A��-��-��Y'��?�ӻG�SQ_\���a<RJC�e;@�gDЈ�)��e�R��6�F@e8,��c��>+ݙ��Z���jS�bTW��u
���^���	E�Dm:�۸\1�=�dB�ߢ���0ȫBoZ�9��뎮��}J���� "F�R�(��R|��(�� h �W�G��.P��w1ޗ��9�^��bX�W�u�#�x�x�XjD�<��A}�!$�B�`��D(C�uCFbE���k5M��U.f�'	�HNm�B[ޙ�Ux� ����E�j���Sz!��4��y�c+�Nova>���]��9���a]��?�H�޽�z�4#=E�X�{�B�z7��4���~]>�ى��Ͷ�S�Gh��.wzW�&�`F[���✫�>�ԥ��nȗ�������ڳO�-F���̭*��&�g�l�6C3^�B��X.�X/�h�+([�����gb��OQ*��%N�O,S����$��5�F� f<eYʰb{עY_�M8<�&.�t`y�2��-�]��Ļj�myZ�3���t�����r2��ٽ�\I�X4}Y�x��Z�<:���w_R����{�u-:P��@��93Y� XGUC�v�貀�oe���sT/e7�ϸ윌ps��&�o��х���hL��uD�h���ysb*M2wY����:�V'&�Q�eb���H�'��ݢ������@Zn-+��D��/��4��LPo�o�30ƶs�[��z���^��d����A���Hj�N�z��K����ƞ4�F��3"�d���U*�mz�YZ��(�v�F�S���"�'�-f�׆�*���k]Zz�@h���U#��2����1S���qf���4h�͚��b����"��<�?6��>n!{I$�+����s��	�w�&�����f;l�q���}��$./Ջ�/�±ew	\��a�*��+��N���q�~��M���(��i�camf��I�["*?���.���#������D��E2"䫠'��M64��GK�S$7�����N�N�Z/���ޟ[��5�Χ�����������w��y�7���ݚ�H�$�C�J|:���DZQH��
j��E$�2�����e��%������M}���1�j�G!̂�#�Cc��sײ<R;P�J��d���� d�`��no�uμf�C��	;��\�?%X�8m����/�l�4Q�u����s�E6���ys��m��Jz�dB�< "6���5t���������̱�_��A�O�������e���Y��~�R�9\]&| ����c�WcV��j��
�����[L�B���9��ҔF�|E�P��.�`+��u�H�I`Iw>��F-�5�d��N=rY����`D��LT76���e��n�K���L <�c���P�4�]�V�@.Eӗ��o�I"gy-)�93ǘL����<Z�l�?`|��I(�e��?�lA{�@6%a��ZQ�DsX ��4K���;U8u͌�p���@^H`x&�$��öY�*�T̜�ʟ��$�H���a�9�m�T{��nb6�����4��2c�Fx6��ܖ�^[�,"?���"�Nx�m�t���i�̊�D���5Gm�u`�Om�|mU̇�a�uj�]���AuyY��:\-���y��D��.}v{>�a��
J=�Z`x�z"q�h� �`2��IS����f۷��Fo�kmHr�ӳ���1��(!'cOI]�PW����]�#�)��L�i�l���*��<j�"�N���ճo�-���Ug?/��
T-$9;6ӛ�vf(�?��&�H�k��~� sj�d�]���3�Ṻf�M�{�N$;������->8�o*E�^R_,�,�zy�f�
��՗J��<���,�g���P��͝�ͼP2{�Y�5`���C/�ګ�L�N���� �����ۄ,w��5_�r�	�'t���?b�E��|���
!\gT ��k�M�� �MY���s��+Κ�Z4��%uC8+�"E@	Y�r��,@���K#��}sZc���Ǖ�3p��0�9\V��v,���0o���#C��-|l�E��l�u"��V�X�z�"lX�����jx0�}��9�\>�;�����jJ�f��������ID?��#�+��T4�К�?��Y��=���53W�#0�W��ِ�2�3m��%
:D��abæUd��/�Б�����^O�Ug�D\8R�.x����K��T�7�Ƙ���*�Ư9W�~Ng������ds�<2M%��z���s��cBANj�GFZ�s�_<�VbO��z���C� ]{}8~���Y�@|�h�hѣU���Ad]9<ڼ}�Z�=Ϸs3������̤T[�!�G��}��R�E�#�A��g�~��R�-L��|p����#��0��ӥ����������?�EyV���	e�Q�ST�,j��z���ʻ1��:t��ܻ��uQ=#!_���q�.�Biɨ���K,,����ɠ�/�:��AoH��K�x��W����Z?x��';0���L�Hb�6���0�Ƨ)�y�a�1F;9��iPB�C�d�ːV�
�C �D��&�.��I��ҴG7ј�����䎃T���� �1��i�?��N�����V��/�"[<�)�XpW���J@��|���`~�b�l����=>V ��|�h���ⴟ�Bݴ����<u��ٴL�UT�Vr�J���-O�oPҼ����b��V��RX�@k���(#�j zy��{9S,���K|�(X��^ڵ��w�}d�G?��5l 1��=i���h��IGu�l���y:$�\�_�G|ᚆh��\ߡ;P}$<�]�ƿ�ͪ'��qf�$u�9�m��"#bB_!�A��yv筺�����L7�J#w�3�v�Iai�t�f��i��1�� 2��Ps2���Tx��J�z�k��ti)�'q��.��LKǢ�Ļy����!Q�R��%_�&�LH~�{�Hѝ؟��B������]z 1��_��OΉ�g�e1��9OP'�=ߋGȹ@����#��1�e@�:����٠ۏ�U簐���r$m�Ǘ>õ�N����gК�a$ոZ�b���_3�۫�z�3�)36�j��g�xj�=7`)��d��ָ���~���2�~�[bfb���mC��s�Q��j��<��j�$��{����Ln8�u]�� k}�4�(L��ǌ�����/͓��]�R�k����ū"x��0`�S�'X�!��Á˕ޜ�?4Eo{W���λ���hB?{�cJ���X7�*n����XZI|�ls;S�%��R��e�d��&�餧��c��Ü�UᭃU?�%��n�#Hv�w�']��2�:��y��]}xy
ɵZ;��o9�OT.�ͽ%>�$�M>���C���0�kR�4��v񤊰�A�/a��T/�2S��9���kB��'a�����ǹ�B �D�l������	�K�����4l����br:��	
����8ڤ��#=4t�>��(�G10�^J������?>v��1��uZe��C��!�N`ǩ�mɦ�o����/��� ��8��n3�|^�(0˝�9�'//r�nY>r^�%֏')<a~��<���8Ǧq��L��9��~��>#k5_�2��f��e"ȇ�a��X)�@�I����"�)v���|���[x�'�!������*�I�ti��������1�k��I��ܜ�9g��lM��&�]+�'��Ⱦ��b��Z�WzP���R�[��ad~U����"�'pvFo�0lu]O����0��)�}J�5��sl�e�ڎ��d�.((��*#q�������pOMfMc��a�"Q]��X9��tө/�b�|��!��O�[#��:m���p��%�c*��D
=�HH���+���Z@��&�ʻ�"�-��I�ro����S�	�dN|:�?����;?b���F���5I|eZ��D����ܶ�� ���|�^<Q�@���N���mu`�:��1���l6�f	�&ـ�kiqP%'}�Cew�}�)�HQR2E+aj��mQ��ȟ��8�}�$��E����-�C�0�&[agG�����I�L��)w,w;�\ú�rq�ۛ�aD��_�V\���Ջ���/��>%܁��SG���n�Zn_�� w;.zZ�v��p�����gj��Q�by�I|P�����1IH���,_�L
�搐�^%��%p4��XBF����ڸ/.��R��zCg�4??ז����2:���B��O��-uͦ s&�z��'!��ዦ:�����^1�
ֲ�Yٙ�Jp;P���ƴ�ԸWX�(�L��e���E[b�b���8��㊺���¤�|�� ��l7����Q��˅t�Z�˻�(��m`p�3��@EҰL�sӃ7z��*U��o����_I�Wg�Vq�5��TT�X�8s@Ol�*?~%�Pl2�>�T���$��`�G�;"E�߱/�]��d��k�m�d�3���*�ams��q~��ꈅ��w٩[b�$6����0�9#1�.�0�Rc�ZPɕY���?.�"t�����I:5�-�)�e�j���;	�ѷW&�*!F����hI��a^*�5XikX�^�6OwQ]mJ\���&�]�Fq��m���:j��>4P0G>:�~!W|��pA������e�w�<8(�e"݂��?g4�}LG��8싐L�z�]�>��kRK>���#a&�m�����3rp����mo�?��5R��u��@��1�-���t%���Mu����� v�op�ȳ��{�`�qx����-�R��?�Lo�RnU�(���:8�	�ϻ�>��cՖ^�X���ue�iµ�Hǉ�;8�q�Ȝev�&�ɘv�叾t$�z}�"M�����&3P'oR��-�� ���l�����>"�2�lc�2ZU���f��=�?�"螓�cU~������I�OޖۏE.�Ql�{M��O���`ᖰUph�{��"J���n���4���F�v��d�)�g���-&�v`���nP������a�-�:���p�A@����g�9��G 5�T�2=�Υ5�*h2-��<�X�qxЇ%�E�/D��/��¾Lƀl���o�r��ʤ����9��e���V�79o^dt'3�k��62�i���h�ʽݰ�B��.�`�}�I�BCh�sðPIkf*,{l��/��y!Eu��#��z�.N���ؼu�����,�=C`�<%*ې����3}��Uj�����"!��?��Qb+c�
�fs�%�����V5��'"�g݄�s*(j�d����@�uV\�,4Զ}���;�P�(�lk��n�5�Ԯ��%�h�i[C*Z���3�@sRijI)�Y%�9��2��m�_r-�y�b�\5�9��4�Ȃ���9pg�ԡ�*d�.��	b�tB����<�カ(�<��"�>D.�;��XB� �U~�E�����E?�I�n��<x�-8��3Iʳm��L5?��0?�,)�*��}92������~:�i���r�%���Cw�P[�{��b��h��T�4��خtN9���<h~�9M�������s��:sbN]L�l/��7�U��j�vv��@UvG����,�č���Ms�Ϲ�ų�{	�[a�{��P��ckF蹡K>�`d���|c��ER�o��\7'20�|��Q�XU{��IhHU�8z��C���Y��8���`�S|o�?+c�t��h��c���诡vz�;��0��劒� �Š��S�d���"1��Y6y�a�:��^͈� �m�/�
E�ʗ.+�%Q�%��U�R����2��D; ���LV������
�:�g�6�$�������Fƀ�z<Y�@���bVo��M���z#���� ĺ-���QnT}%�ҷz�n	fk���������O� ��$,�Ԉ���Զ�e�@�;����`�2��F2�7J�.7�z��������8��7�!���j�wrA.���7׺r�v�z�V3@m��$mx�7*K�����Ã�W�"��پ�EpD�i�U9�a�է&2`��^`"�]�*1~H��Lm�>a�|��	�z����1�"�ݑ<(�����o�^�\�\O��:k��:��g�e���<�PF�t.��{��X՛�G��ap���W�!��F�V7���({^���߆�۷���Ij��Js��Bk�Y�+�w������۷E�}����g�9�rnc��]��Z��S�x�h�5��sq�ZAj�J&)�Q��m9լbf�~�+�N�n���(3�P���%c0���2���d���T��)�KĨ_���*w-�C�u�rr���t��Ys]�5M/|@.��P�ͽ������������`�ik�Ù������4�R~1J~�'�� %��gk���cB�aK��m�^G:G��ҿ����e������1f�mU;ۃ&�%��ޜ�7�"�\^�"^/~�7\����WԞ=~F�@�a���J�t��7��,K����O@�|���L�'BE�Wl?
S�p����"��6��s�5��LI{z����b��{��覹Fi惴;G�sFZ�����O�	)��U�m `���+�#"�0����z�]d8ce^I@�w�{���;�A�In��N�-4�Dlٱ:ØE�A�wS��l��������G�B�7�̓K�zѫ�)��­"�@4�X�@+YR���]�TL]�ơbOFaSs�,�FB����W�X��s����_���Ӥ�P?�JC�Tf��J�o2�ʽk��*�L"8����~͇)�̪L�.x�n����7�W������Ĝ��E�]���w�M�0ԓ���
I���=��U+N��-Z�z�f\,f$8S�������4�����Ⅲ왌O�%�5�:�n[�07r�<+`�����-��y��ۙ��͢�4�'dFܻ��`mv@[�i���šf'Y-��{��i3�:R���죙LG�T�1F<s�b�W;N#�͊ny?�KJ���v�5��{��9�k�Ee�|a 6B���K��6��/(�B�o��D�W
Y��a}������i��H)���(���d�����m��i
)-��.�ʏ���Ӊ[�7�>>�k-�=�@x�/��*e��}����*��d��JQ��S�y8��P{d|��"?A�d�?��c/u
���7ʍC�^H����w���xy�;��Z '�=8�=(�©6�D~;�H���Χ����α�f�@�<�źI�^\C�p�E���V޳������- õr[�}Q���_��J�\o�f��'���+,
e��xH±jm������.*n�[f�QPB)�!���.�����Y��b`*����}=�_���,�tVuO�<(Y�Qj�oW�Y�mԟ�m��z�6ߣ��사ZTW��n���M/�ɶ�Q:�b%_�_�Gst����qN�F����5s+B�؉���`s�H�4��p�)Eԣ�9l}�(\��Ҷ� I!\!1j����F������-�JT#�Q�ņ���;o��g ���7	
�ä`����ʓ8�fQ��U�s��c�{���N��pBJF����~�����3.�;�	�r���>Kf�m�~O~_gxs�`_iE���}�*��{�V�9)���^��̓��Ր	��z\�\�`�|c
\� �wv:e��r�[e�l(}���� 諭HY��~O^��/Jg�e����]%��暕��X��"�@�G�]|B�?�®٦NHN���ch� c�a�'�*��g��q8ku�l!\�(�A�t|?�j��P�i7vn[��Ch?����y��}��-w!�Rmֳ\s�� ����:&FXY59O�Kڮ�j/'t�-|���K�u�0�_D�����l��
 �V��N)�X����F��hbX9l���1t뤥4"/��c��D�QƾP!"eJ�xE�vyx^�\��j����d�����c��&n�֩��޳��ݦ3��X7�� �B��r;fDa�*M>!wVJ�[.\�v�XnCo;�2.ڑ���� rQ
:�ʹ�%>a�f��#>�� 4��أ��g�� �Cƙ�1_�?Z\�W�N�5Ho���+
�=���Ȇ��׋k�c'*DD}�����[1x,hEK��!�el�e3�1�t�PH�E��t�t���х��9�J�� �굼Tбg t��i^��H����T�'�Hd "W,)q���ȷ�A)�����Z�� &z7�К�z��k 	�?��f)����˧_S�~!�+����+HZ}��dV8���ڻ��k\ΊS�,��_cF��Gp 80�c�.�m��u��ǥlQ�_��}q!x�Cz�S����(�Q��ÿ��9�L����u����M^�}L����u��ZP)#[.Cy|���<�p��5��6�So�f��MлQx�r�id�&�ꏌ�n�8�-g�J� �C��D���k���dC���:�O��p��;�+$�\�����-X١��a��"���3- c�]�I�Ů̘D��==�q��|sL��>�sY���\<�n�	[��X1�N̄lY�dE�*�G1��gu~�Nt�A��e>�� ��Un��fΟ�л>%�\F��61{��\(8.C�F�����x�j\r�5z-$q�2gff�H����	��_ЀD����c�uWk1����t�}Ċ����N�sn�Z��1���-�Tb׿�����ν9�Æ�J8#��������_Ȟ���	T�2��k52z�����u'H���O��FU���� g�E$Ȋ�6#�t�~�b,Ή>�i]{�z����DJ'9r2��q�]Z�M蘿a+X��e�(�YO�S��V/ ���.�ѹC�6��W��	���l��}�����eB��ֱ-3���A���v١<N	�
p�����kΛ�7֗`~��34^m�M�`�r&C��
S _��28�s�Wr��K��/��A����,����W��:�&E�-����n.���d'c!)�8�����>�fǐ����A����E�2{�F��4��߲X"z |87�Q�p�"s�P�sg�q����p-�-���k�J�+p���15��:�� �6+����Z�3(7ȿ�}�C���X���5�~�̡WQ��a�x�&�7qB�6Q�̗BtP~ECʁC���"��ͤ=p;/E��)�k�Q��U�,C����!'u[�a�"*�S�m���j�γ�|Kί��cXRp͸ٺ�2}���M��ُgI�r�S�Ꝟ����s� �pc���Ռ�71���`"������m�����j�ԯB4l��v�BW�x��K���o�R���K}�~䲾_	:H�ā�!p���5%�\��sU)o��Fh��G˔>�8K��>LG�tg��{����֛��<�=
]�J�)\&?�~�����gRa�� 9�K�@�F��ᄡW����}�s����O�	�N��"�q�M���6Ԙ ��*\��gR���?0�{�E>��$�a^'�t�ɝ�����k�� �#JT�j�F��8�����SZ�9I��LL�]c�[-���f�`0I��4{>��|*m����. 8]N�9��8љ����45P�45�b���������V|�
%~� �F�L#��Z������#t�x�f�p\C}�ؙ�޸|S�$pZ8I�N�&壔��%,�Gyj��v��ظK��H
΁�����<�mV�C8l�c�.�fPQ� ��6b7�e_4��H��d�/���0'e�-*͟�$���@�����k&��1/ʲRp�x�r�|��O`�*�R����@���;���'4k�%#z��]�����xÕVL�+ge)�z77I��H<H�p �_p�Ԏ*wW?JGm=ɀ������=���ׄ��[_��-��-�IoMΫ�Т@$y+ۉɧ�$,�N�Ҕ��m���N�����z����" ��ꐥ$�9����7N�6��Ųc)^�ƨ���Ϡ��1h�x�	@�l��?;r�oз�Z����0��Ze4��#�����ժ���/��K�a�OOn���J��d�6�|*[���lʁy}u��3��ૄ�"ҭ����v�.��CUġ �{[��+���A'V��I�����	g�j� ���KO}>�smN��rH�/lW	����u@,^|���$`S�8��K]vP����/)wi[%&��]/Q쪐0H�F$xP���В1aU��.��k��3��j���4UuNL��jn/�����Q�(Y��W�z����̌�Z)��Ap9�t��NS,(5��PQ����'��l��>���EL-��I߬g ϘQ}����Mp�hA��9
�ε7z�Tۿ�����?������y���gб�4N� a�}#q�r��G� ��|I���<q���z݁_­��x=hg},�c#x�u��p��7%8����y���
&�U�(c�i��!L1G��#��H|A)��h������F�p~�o�墫�g`�/���r�a&�q_X�N�y»�(��`:�&m>�[�)�oF�jL�t�04z���hq���X�|1��.F7��iQ�d�ƍQma=�|�ۖU؟(������������}���xA5�R�sx������qxwLE#k\��;�Ĉ#�UUm|���`�=[��!��+f����V������xy` ���m.K���p�Y��[`��æ�m�tC��tg�K��6/������=�fm�cB��/F6O1��j|�e�%������:� V�?Y�g�$����gjfo�퍠��y2��]hD�U�t�?F��b.�Sq2��be^�fZ*b�����7�/���5��1�l}��B�����T�\u;����)_wf�������p5Օ��֕���7m<���ʚ��&�?����C�h�O#ע�S�'���g�ý���;�N��|)]����
�"8p+��]�U��?ѵP._v� j53�t��e��d-o���?��Qf'Ф&l$�����hZ��U�������DNJ����|M��{�$ޞHk��t��,��鬧��sr��;=�f+��ӷ{N�'�]�Tk��I|��mF��F���[��6��j�S���A�1���.�7d�vv��?]�0�^u���@Y�t�us����=8�P�γ���zQY�氦��g�7�r?1��՜���]&�M��ѷЙq�薲ծyl��ӓ��k��寍[�_��Int��)i2�?~�u�=%�S����D�/�s�p�[m�D?<�f��t>������1��
<Y~vbs$Q��v���T��ч��UH�7Ƕݯ-�RQ�LXk�a�x��N��9�ǳ2�E� �"i�R����h��)Q- �d1�)����E��:�VڞM'T��,P��͇�Ч+b���˩�V���9�<��|3!�r���
����z�c�d��d��8�Qg���P�E �TŊ��,�Usp�qGb[���?��N��C��ڥF�����"P����A��5�h0�S{�eƬ�7�$���e┸�+{���qN&!�Cfbn���m�+���Z����H���
���{�"V���b�XL5vٸ�p��E���K�mUz҂�y|�!�&�+X,��>�E�W�7���C`U ��K����ic�#BO[R&k@2�h��c�~�oǮt�+�O�s�&Nq[�EdD5�Y�mxβW[�z۵��>~�R=�'�i o��� i�3��C��s_����[��YT�R����z8�
���T6��e�nVC�ۄ;�D�"e� ��w�ȗ��������ݖ�,
���ԓ�Ǔط�ʁ�r5Q.�QH-��� ��M�~a����M��5�m~�'�gd��CVK:���<�xT�Իܻ�����I,X�!�|k{��՘�1���9S9w�.l%�a�l7��[а��
&��cc���~�������w��]U �z����K�?��.�������V��%�Q�G�����{%�XG�]��TMY#
���>҂)��QtB.t<)'������hf�#�6d��QrD�{z#�;f��-�������؃*��a[R8��G�o�`��lཎ [��&3�,�'��q���k�}�[�O
>�S���>���R�y����-��;�I��'��Q�k �$���fDSbM�c� 0G3��$f|-Z�4�v���Sy���<%&P�t厦ܙ��ו��@5;�;��u��Z��g�I�Z$��H<�#�gE^]o`�lkI�9�y�=����Dl��������}�$��I����ӭ�F�{}��n��	��Õ�����Cn�>�8٥���/Gfe��'j6zEvy�� Whd�|�m�����q�Xp�Wh��?���t����I�Ha��g[�8��9M�{�|k�|"
b��J���g�ȓ�^_3��H	F�|�7�,i�-U��Fv"O�v�*{�K��[�d(.�OV�=�l��
���~t_�^�`�"�Ы��=���,��f7НƧ�����KU$^}�I��<�q\�0�	q��V&!�		���`�?d��ָ �I5��+7)R~_�RS|����`���F�����J?��Iu�+[[�1CյI��AW�r�)R+��SeO��όjw�W"3�N���G�O��D����	.�^���\�����3���ˊ;{�����#; ��#�� ��HTU�M����@�2�hI|%�~(V"y�E[y� ������CJ��S{�p�)�f��O���"T/c�;��O�U"35:7�V*�)��;H�,6nc���I7?|�-�+�*ir~�l6�\ϋE�[_�X9�oD���M���Y���/MX���}�"_�y�-��a��������͑8���_*��I%s�l��|֍��;���h�b�:#�Z{6x�9<�x�a��,~��A|���H��A��KT䟦�Q����j�ӺI(����YU������e�B��[>A�N�ڤ�Ik���T��z��(��[�^�	���L�&$+,�vi̻}�	���>��aQ��E����^u���9b�����(Ւ�4���������T*!Y�Uw�Y�]B�u/tP�@<��U;8w%�te6��|MqtP�'���BdR�'�`��\!���iF�UE��d��*�����n�sh���P9��fh���؅F19�ث`�=	�DAo�w���z��ֱ W�r��oԪ�[8�>�>���î�����K�.��.ʘ1����&�Z������O�L���0k�u����&1=3��v2�84��Y�����ķ&��S��F;�~a�9I4n#}��ڛ�U���O��w��j�#�p��0��$�u��f��5�#������w��E�n�;k�X�\B����b�PM߽`���r�����`�Y	Z�� J4���7�����v"O73$ �I���1�s6[#`�LX�;�/��Gir����2ОGC�YW���N?A0N��F����
bN��5�5-i�FS��_��;�P���1Q�o�6uf��ݘ��K�1��� �Qˁ��a�Z �^L�J�5Ʃ=%>�z��g��챰��h�ֺ�/�����N�$m�lR\�-�L%�r���j��Ҁ�S� �Bi�3j��fofLh� HN���\�Z)W�-����lf��h���+�ԋx6���Ri�'co(�	�	��J�5�	_���b%{��i�����M�h������+ x"^9:�|�B�x�� �z��p����'��d��T%�K�A.O��5�YWB��w�����Y�|س{��p�{��JO��*�K�2f��a��-�d_x�*�K�~���Yx�Z��r���3Ff��d�Ȏ'}��辗3�K��P��Θ�
}�B"T�%��K���~]q ���V���I���Ǧ]*�ʟ �}P��Y]�����%�l��|��SP��K�N]��^Jp�H7%5��A0�r��L�0�1��)������5x�Ϧ#I�"MZ����3J���T����0�D*-����82{�9?�� s��9\�ˎ��%����t�R�FE%���*����y�b���tZ�w�
�bKT0:|Pr�Yj�X�T���*l��x���3)�K�콛�߁,<A�s�V�3�7�"R��4V���c	*m�Y�<��$�<6��\34��<5$��=u�������pGH�w�L�&L��&��/$��	��c,����}ڶ�ݝ��ubp&�Xf
>��f���o��0P�)� ^Gn��an:���+V��i����jիG�0�^�6���Y���
�ٟ��l��
�]Z`����j�M�����^���U��)��9%S��C��_�x�#�Z~r��@���s)�;�JEs
�tl0<͵98XdN��Է��RT��|�~��ġ�s�x�c��R�c��l�w�c���Ko]�tܿ��=i������gK�^L����g���f�?�ϊ��0���m��nҀ��oYM���|&�_�O ~%!9��Be���UL����z��u-_5���<ݑ2KiJ]����R�e�"��^x�w��1��j�D��N�&���Y}E��搄i��o�-�+�����-��Swi���9���\;͛�*/5. �!��у�ή�@H{ǀ��[��
�A��U@���LӨs��)��e���~`�A��O��@6γ�N�|\�)�Fqc7Cx�I��V��&W<�~n�9t�*o\U��Q�4���?	نUF����́�a�[�w4�	��%�,�e�F>��{��V�`�I�G�I������?�p�T%Og*.t���:�I냛��4ZZ8׵m��a�����*g��8^ ����Z�W�ĉ�>si��Dx&D��z_������+w�����X"�P�.RL�=erJ��5�]ao�j#.\�f�"W��ٴ2������}���������i��x��/�yA11T"3�[#S�W�Ni�߀����5���Ƿ�D�PV[8b�������	k��������]�I�
�A�3��g��g�G�i@`	*�S��q��&�^���e6îs�h���`�X�w��Qj���Df}ސa�Pz��B~�@y�m�!�v$D'����+8r�<�
���Mc�U4����K"o�J"�@�Pj���c��q0�O�M��q|��s,:,d�� �T%l�Y5)H ҬS.�c�h�%�l?�G�	Y��We�~�XZ����tϩ��qr�h��e����uF�[������� T�ރ�r�2�}3P'mN��N��^]�{mjD
�2�~����}���P�P$_0ͪ�m��l�=t�chA`�L�i{�yhx��
PP������n���& �oe9/ue�n԰^g�WR
�
~&%%;fnBq��X�R��%
i�޻[��>�&����T$�#?ԋ%�3dH����	���d@���?��J����k�b��]&�e���k$����1m�dT^��dBM;��t�O<aa*6	�2���ށ����Z�2�C[vTp�ʗ5]K_h6P�Md~����-u7�w`P�qw4�z? 7�������׃er��;�����q��rSd�hܫ5iE�:����s�o,	V]յ-�'���]��a�J�#��W�>��¿Vl���w[]���T F�dH���8�C�1߲2
����ԕv�����5k9�Il�6�k�ڛ���}����M�����Ӂ�:z^�P�^�x:�ۉ�qz^����MW�x��Ƅ��5G�-���^��cSg�K1s���@� ޾;�b�a�솎cd#����<	�B�ف��o��y3}Cր�l����=]O"�,`^��)�1I	Xڿ��()�D�(��)j&�BS��n���گ����~&)M�C�i)�^��p%\�Q�O�U��m����"��>�[�1�ދ��
�e}N�v��A�ɭ=�JK� �/�iվj�R��.���M�S]�q�uc,[���K�Y�'�kPؽDqdM�<��ߢ0֞����^�z��7.2�`+
C"�L�_�h���\�8���lh\񨔐ӳ5����@v�HT�����^!x�CrD|�A
`��%
��ń�٢�R���) �XY������ԢB<ֻ�c�����>�Cl��ݳ*)&4	&����G���p�hH9�f8k���6�#=���u ���*���+D]��D��X�#�|��s�?U)W�SC\ 3vףO	�>��4?r���嚮G��j�1p��{nmƀ�G���I�t"x{N#.�u )�]�R��I1�z���<���R��E�)�4��oA�x� }�/!D����e�t&�8Y��*�/C��Tpx��A��%6��*u�Ú�`���p����c�,�� V	B>�;��%�ʔ�-��8�l2w)�y��bcn8�yJ���N>NdBu�� | T��*�`�/Т���ǈ�̞=���Z�����xc*ߺ�iXD18ա(Lo3V��Q��t���,�0qg��}������U�YŰƅJd�,2�[F�9��dѺ�Dr�|�8^�y*4�?5!��fz����kc=l2�����y���Mj���tY���`�\嫦���x�I߃-�����w���쇸Qǫf���9�d��4�6'�!@i�`{ ���rw�~��t�1g�Q�	�.!���L��5aB^���E�&�b��Q�S)��N�o\:��Ͻ(-�Ws�Je��&�81�؋]��v�z��Y(5�Ϳ�)G�
�Ȝ�q;�y�����$�ݯ�)]ܘsv��33�r;���j1 ��E5U��TV�k�eI}�<�[������3��:�'>�@O?ψ�S�r�-8����*�8������>L�S�F1<}L~��ɮC�p���*:��jq���v�\�B�U�����	MK���SX�VPŹF��x%t?�Pj��m,�O�"K�. ,�7�L1*��b)�n�`<pf+RŹ���sP�F�����Y�49��A���ó6}?3����i��a�^O�5Ŧ�Y+���\1�p�{���xW����W��Yh�d�D7�.�,?Z�^��)U������7w-��wO��G�.b��*��������(��r<s�b|O-����"��Ʈ��}ץw!8�g����Rs��}���2+�7�S�w�e�X��]��RM����6�̭R�4���� �"��!���eHq���^�M�.�s'��3�Լ�.�*�g����!���a��S��0]�D��9G���۴�x�R��3�d��aշ���_	Pd�R���ߟ�ې��*g%��A-D�e�?5�s@-�����,.�{Pj�Q��<�oʿ�BXI�����C}��/]��
���:��B�+ז^�>��+��u����+�y���~�53q�l*D�WC% Q!p0|tI���پ~G�sE%���9p�S��[�[�#z��G{T¹��B�;�o�SR�����P=GIT�����������S���%,i=���`�jB��uUZr����R ӻ~��=�,��E���s;�`�*���;����~X���o��))O��[�4�����ڋU�B��M�1�q���S����̎�����D��3��|�M�"�34�Υ��U��K��HO�3����6>�n���x��V������_Y�"`8��xK�y]�'\C�O�]��|gn��"Qd��g�{�+�	��x`�-�+I�n��i$�d�v�����#�=m0u�~*í��	D���~'σ�h~-�s~lm�ݙsw��Q+x����9��ܲ���v�.�����x�Y�by��(��!���K��%�Rɩ��	}�����P��1n�=>�'��`�H�P^�����[�� ���D?�ax��1��;/�vi��i� �EG�2���6�
D F��e P~Ps�8������Ů�!��a�P�
��c1��B��?��y""���Jy�Z�9u�_�ܗئJ E�|�����K��>WMF�#M��O�����ۓ���veNY:�����%��g�kg���" T����vIY<���X�"��Lט�!:��e�4�f]��z�p�k�Il����{���=��P�8<nZ�s����1�H40�$Do��}A2�#U�����դ�H *��6?�M[b�$Zt��%�鎆�f���Β�!��b���삏K�CY�!f�=#M:�1���Նlk-<���@�"p�Z���<�-zb 8��wҨA~��dˆ�4�(� }�[Á;�x+��&�������/�k�K�R���swOE�ڣ��+.�*�����Z7��Q�TZ��>���o=+���Ŝ���u���Y��V-Ine
������=b���|�y�%{aC�L7��c*��ci,��K�	�yzrv��
�×��d������-���2��ޙ�[漀#��_��>��iq��4���[e^LW�,�:���� T߉պ�(����T$H�>y1@hr�:��Y�W�6�����Х�k�'���S�V��0�x��5�zZ��O�L/�;.��H:�n�JW���i�Y��A]������>A}��5rb5u����'�JRI�b��ຖy7hˑt�;F�X΃��y �[��2��dY�V��eC1x~�5 �X�ÕZ�*�[�i-�ƞk��t�����M�f�Z*&&�<j2�nPc�n��c�`ɹ-��DM��?M�/�Z����&�k�ݹvnVI�^����+e/����Þ�$��b4���Qk��=�=���c���(��J�+~�Pxhx���xG�s:�6%ҁֿ
��a�ڿ9�֢8+��Rc��|�6�%Je��ހ�a,�ԉ[����dٓAs���Ε<SJ�Y�I��Ny��M3�2:Rw�з�4ս�t9εE��b�#�,=2��hM�'����	���������k���^���3ݻ��IIJ��O�	���R��8N��3Y�XYd�Ys/Lf[Q��d���Z:��*/^�8��+I�́�۹'�`5u��߽M!#���*F�[\nP�>72~��e��̳�O� ?~�⽕κz�)��.x�	�2f�r����<�d�n��zl��̞j�%�#b���	��>=/�!�7��Io��9t�>�Hq7φ~gz��·ؕ�i��R*����{���=6b���t?:�	S�쾿b�]bW1yg����=�ǧ%��b&ޠ��4g�eO���VG�%�V)���{���]�@`L��
�{Œ��;�CcfCX�x��Q���	�W�H��(�]�P,j�����*e�8~qY/b�t�u~��
L�(���!�B�n��K�6����^�����v�!��{�X-�q�a·�,L	f���j���8v`��,��%i����H� ~ض�̬�����y��1�;�J�YS��v�N�R'�C����/��Q�*Y����n;s�7÷��s.ձ]m]� �G20t���C��Z+V�T@��
�ֲl&a{�'D�Me连F��`�OC_�s�qC�I2_J��*���]�v��q wO��Ƹ����5�n���
�ʨ�dC����Nd���$��ǵ��P���h�B�J�B�@x�����T��y��t�EIuF�Ώ5�W5ޗ����l?nK�qŀl���N��mL��_���a\`J����o�9��G9͘���Pv5�hty6�Z�D����D8��
�j��/J����-8��%\�ӽQmvG���0���G�O�4�DY|�q��|㴲���ұ֜�6�i�k���?�`����X��i���WT�`&"`Ks�Ѐִ�8��l"t�hkG���΢�}�9���V^:vu�)�$�}��6j ��.]Y(<ٳ������QI�[���s�)�KC�ūㇷ�HRFN8|sL7�w)E�"�T�V��� �ffj:�{�ꀞ)�j�3-|����K��Bg�G�ǌr��\�O���{�ɗ���3��G}��e
�ԇ��K���4}w���H���;�_ң�(���x����T,`\�&�;�� B�^r�-���}������%9i��3�k�l0�+}�q���aġ�]\3�%�R��hd'�v�
>�I�{�	��KD0.�/&��ʲ{`�dC�=� v�
�4�S��]ULA�rw�!���Aޤ)�O鬊a�ק��2!C�3��ᓰ�:�밉�S�`E�;w�D�����w�����䝂�V�g3�d�����"��_`x4����T���Ďpz����)���+t�e=f�A�����C����w���_F3΀�\�SD�ʌJ��	.��ԉφY#f���X���{TBnL�o��Pr��Eo1��*�uS�����~fp�� ��i�@I,�_�G�d�ҟ��`�gy��\�aښ�X�A ���F_X�r^��%��u6���h�������ʥ2c���:_l5+ghN 	���� ���ۻ���Th��ͫ��F��	c����:�y0��q�r#M΍���n�O�:Dk]�i���4p+�{���(ܟ<d��X��f���<�B����p+�C!eBq��I¤�?W�G�{p�	����;��v�
�e�g���^�@#抌�O3�WշJ��M��6Ⱥ&�I��qE,�y)��=��V��z��v��V_fZ���I|�\�l�s^��c�\�M��#�Y����z^�ko���Z���Տ@�D�تj	��w0 �*�zxWm��p�����`IP��#h�C��.*L`��^�:���Afd��5����r̙|nG��ʻ�D�Y���\ ������7l��;p���1���	��V��J��� �o��*N1�:��v�Wj�D�{l��3�i���0{q��1u7��r�3��a`'#�?g��u>`ͷ��N��$�{�� �	�+\I��^��-��g|5�H:��AN�}�s#�d'U�`�Q!��RF��^ec��JMY���
Q�J�L���rnߣ��lG%UC�?��,�����"����*���E��t]�$���
��&�z�^�T2۔�r$�+T�*��rSg�:Q��>��f���V�R䪡1Q� �A�1	G^>�v��ve?.9Mk	��K��N"��Ke��������w0�0���A���gп�Z�iże�ٔ`�33bc�J��
�T|��}�� K�f�#�5�4v=��eⱳN��S̃"<}UT��gZT���\a�W���|X�	[}{�Ed@�����nj�}��n͗d���pS�m��9!��� ���|ڠ�O��̮��9_O�ľ"zk��l �þ?�4�T�׵�����i�Ł?e��(.�p�������H�h�N�ۺ���yt	^��������g[�9r���K��'w�~�/������e_�`��-	K�Ǩ���u�Bt�4��u9P0�e#������h�nLcg+��𸾁�����ֻQ'�ڨڹcϣ�v�ȸ�6���� ]�4OknK�E�锇&�*��N�a,NkWdaC�0��M��M�= ar��0H��U��Yh&K����3`�0��@&x���u^=�!���)���?���N������A�zR�9E;�mCC��ȟ0
-ꉃ���U����mlR�l%��tݣ�f9�t18��Ο�j���&��p5�o��93��_I����_�U��/��[J_0�VD�[$�"7�<��F�]��j���'}̨�"�!���'�,�I0�Jg����M�ƃE�03�u��H��N$.,�7�M�Z�����@��֭���m�G��s���g&G����C�8�t�� ���-��?�ƫ��@�����͵��8X��V�=]���"�t{��!��&m�fvlZG"��$�!�wb��Gi�
�ע�X�RU<����1�fy��$T%�SV��T�&2{^ͥߑ��ضJqHG�^�8�������;��hɒm���iy�w�%���G�#� �au����d���&��W�fo��4)����_��Ӭ�=`�<�u�9����p�yB&��}����L�.�{�����pzH���='�C�ʰ$�W?Pf��ÿƏ�c�����$"�D�骇�̜�Ј̛K�]j����f3O��B��C�-��?\CN�Z�y�_�gy��]���/���Q"�Y�r�MsN����T�fUz&a�E�o\�J���P�-gq"da/��U'Ό��O<0�+��`2L���	��u��1U쨄�GSN��W�LM�x�9Fr�uYqk����|䅰��m����7K�ω.������	�! �&�*�*24����u_~���I���l�*\2�K�"ꭎ�q���^��Γeo�U��9C��^�s��e��{r�K�gZ��N�!Gi=؈��=Q�acyW,�b!r�j��Z�1�p�i����4"����uIW���t�D�my�8����Rr�۔�w�
j�_�P�tVN;�h@�?@Q:�L��l�+M�2���#�ޭ`�y��)]��Q�i��n���h���n��p9<耣�[�2�}�����jB�خM�����t�Ï��M;z?S�}��7F�P��*=bd��nL�5<C�Hk�xzc��{&�r��ƾC�v�yé�ȦU]��tx���/�G���}�h�`p���
%�&�Sqׇd�J���)�P��{s��.V�Vq;gg��L�Np��֍g��FN�n)�G�<��7�}�����1�5!��I/.��HH�b��כ�I,at��*�R
��yF�a>�Y���	C~݁&�ݦ�9���LL���1B�L�6%hm��q �+�͆��`/�
��V��?����W�h=�2D7\ ��&��Ճ��<��C�.43um�������9�[�a�!6Y01Aࣨ
�� �ͺbp�:��`�W�n/�@v�a7a܉���op���,�.�ӌh)A@{n��^�P�@n>�_�
NN�V*8�C�kӫ?��� peӓ���ʎ�3��
�(�nnK,~��%�*�� f�Y,���!͇��v�8{��u[���E���غ.�6Ң0�HFb�xáD�(l-��-���b@���n���jA��S�������jlDs�]f�9��!�D$�l��e�f����ǮS���M�����in�m��n�����'�#�R�_������I���ďXv���bo>��W�[;�8�"���~)�VHgu�)$���N��W��}�(u�[���`��N��=���K�TҖ��L�2Z��#Ed�qL�����?A�+�PLJU!l���(r�^^�}�é8�x���	����s�mp�"��Ƨ��e��q?�^����d�<�+��2xX��5�f�Ȇ	��쒪5!AY���@����-��<ԍC��d��<���i�M�8A�0�#=���is�����;�E4K�وFP	appw���l,Fr�sQ�� �Y�1��Xݗ�PO$ka���58�1���	\/������YR�IM+h�3�k�輽�A����U���b_P����N����Ѭ���DR*`�kE���\�������8�0���z�lu��e=�B�⨰��Q� �8����h�<���t��Ta�p'
����5ݎ�ؕ��V��p-^�~��bR?=����R���yj}��[�� +��ɐԸ��gX�Ts�����ץ\�J���~��*�D]���.���?�z��[����:5:�`/�s8K����r�z��/�O�ʁ���m\�G�cAT�[�2G֦7�9`k[���W*EQ�ȁ���vfn�W������V&����|��Ղo�m��n=t��^�@0���w �y�p!�yhd��+Ǯ��W�����|@?�� �|I��U��+��R�:=�#]�|>��#Ns���e<
�@h,AY
�}���7��ew�q�����PҦ�t�z�3pC[�&V��n4�=�(����BTw�F�2�Hެ�s�YEF�(�0/�I;/,O�)nHĞ�¥�q^�FlW!�ʒo�lP��­F�tޓ��y�8p)S՛�(���g����3�7�#I�TI~���NfX�cR^�Fv%�I�'�#�rh����������"�<�@ws�,�<4L���Kϴ.��(N��2�\�^=<<��*����e0���h:����%5�w���u�i�m��1�S�K���A�Q��Fu��5u�R�#��mn�oT�c�ĝ2ű�ӸT�ղ�VX�����#fG��ꐱ�-�i�j�::j=�et
�NR�n>`|Dtc���Wcr�P l|�꿐�8��3��[y'/&'�XV�#u�Iб��th2<@��&`�����k�;A������k��c��*n�-n��H�/�m��3LP�8�Ğ�eiPi�?�ZDr&�rZx�:\�pܸ\�K&H�z4J��kt'�)y��wPqH`7��ޡ�c?ζW�~�����;���6ט ꋞ�nd�>����I�"��%�3Sȡ���_��C���!�͜��G�cl�ɟ�<�ZC��¹x��������=��&U�)�<��?�ɕ��/Ё!�����T=�:c+Շ	FB�wh���i�i�<�͞o���ӯƞW5�m�a����h���P^i�Z�X9��Ծ�#�	`�lǡ�96.�M킒G��)_`M_ã�`�z�,t���!5K�&�D�O�qO	ٺ��9�ck<2p�?a��U?�^Kd�`�-Ö��aRM)`cE����.��#jt���L��eS4����Xc��FI������h�y>���_�8r��]�������k����]0T����u$�V&�T���W�wa�Y�'а�������A�P/���u'ϋ��6��6)x|�����il�ZP�cɕŞ�n��t!�ן|e�E.D�v��I�w�f��mRe����l��Af�'�t�y��^��h�C~,0)�ff�H�&4�#]�Q4	�b�Iu~I����E,]�˱��N�!P�q�]����c�n�m����F6�$��\1���cq+8Nz 7ˡ,���3����n� `�т\���ŔwK�0�s8���-A��ة�8 �D�b�y\��H�ê�G�=�0���vd�ߛܩF������m*�wepg�������yQ��ui�Re���#5���X�6IE�
�Z����^�����ٌfOZd��4Bύ�)����B�dAwt�.�}���An0,��ˀ\:����˥]��y�$����ظ��1���y���E�7�����EkS�)�{��#�њB�8��LK�l��d1����y�6��t�D� ֧J���6d6���h)����,H�5fr�N⣉��v4���k ��K�:�ˑH��?�γ�*��6�O�� I�䪃��|�2l������H�GpM�{�fVE��G���5��`�����N���E8���.=�;���&$G��1��O�M��d ����X	�CU�����-��J%����u�i��n}om�?���߾�E~6*'o=c�^34��[kp�N���	";y��Yy9ͰE�Į�*��(`O�������4(�r��\�ۛ��{2�Rr���"��o\�"�#������i�ⶶ�BW6����-�%����E�jN청{ᱞ��G8;_��w���&�л��>+��$���63%�b�T��~]#�bT�^R^��f�A��6d��\�9/�/�t��חޑ��u5�O��N��%��})��@XA��qf��V�˭��+���!`�$Â���^�-��!�C���4,L�yX�g6X((����!y+G��9��Bo��r��(}XH)��#�lJ�bn�"�����Cj�ne�k�.B�G��|�jI�.�{ul乇Cl�&�M����p�0T�w�\��N���4��=H���K*���CW��2����D����R��*�W�X�ښd�Tg#�]�5T 0�(U߰)��ȤL`�����p��S�/�nIh7���<���j�C^�tqU��2,�v�)8@u�t�D,]JAJgc��$��ҥ�û4�T� �;�ej9��"c�oMOP��nBqB��v�n��*��pj�>w���&�:n)&���XT�t�&M�2�ZpDrCV�-��v� hh2V6������|�)o��(�2�,J��",�%�^LW;� C����M'�o>cU��4��Y��نz� �hFqܰ��_Z��D��/��fj͆E�V1�<h{>,�P�������h7�3�ټ��]�#hL_w`�Ŕ���bƚ��-bY�5Ir�"EC\Z5��1����K^w�FQPijpd���M���s�bu��$.�n�g��Z�s7@cN%�x�����>ௌ5T�°&�z�L-�{v�g��x��4�LGߢ6g��K4!D�P�f{3�)�`�������D�v,
��E5UI9�B�	�X�|9L,�Ym�^���,g�КUp��o"�C�Kn��Ɗc���v����)��flΙ��ڟoB�P(�lQ7X�O�^i+�{9�͐���~N�����Z�?�՞լ�\�wNh�|@��Sd�;��Ţ�\�Y�ZSA�5�z��P,��BZe;�=,I��wd���Od|t�+Ɛ�^ ��g��ͨC�9��G����~G?�L�U���A*ܕM �m�fyE�J������T���ns��Jt^��! `��Ͷ�g-�i:�4!֌	D@(e#0*�-W�i�}k����-��5N��H�3�d7�Ψ9aڪU�o�$Z}�x����]
>:7������-�7�!��G�T�l0��������Oܚޞh��#]�<�v�4�oڂ�Z]����%P�Q�E��>����QEG�,�uƭ���`l��lh=F�m4�ܰm-NNN�F}�@�0	��r�q�ӳ�(��n�2��z3@����IcW@A`H�55&�"�4�.�_Ƣ]��9�0��"b����&=�M������1����5����Ʉ/�Of�ڍ �n6�ݭh*f�����_}[v�`��5�'��
�$�6�>��S�����G�=}|�9�
�_蕷�ʌ���׬ll�x� ;-���Z��M��Q���8o{��z������c[��5yL�P�����ϴ����urH)i-|=�~mu�wk�O�w�삨�\�zd�,w}"d�M�!�m��W6�gr `�v�^�r�g�x~�w��/��U��Y� nZԏ}\3
��겦�����Z��Qr�"=u#���� �r8q��̆s�μ�R��]��!�:&O���HEs�<QC�t|��`�,/�8��|�T���1cE��P̣��>��|�̌5��n�jK���p&hR����#+g/�-���5:NK�nrM�r��#_bO�	����{?�3k��+��������+gUS�U��p��9��Hb�V���(K��=yNr�]`n�1�ȣ�[<�vܷ���Bj��m�z�W��6��G�I���P�0���^��� 7�Q
�;����κ�9���H��
V�8�G��O��j�*c�M��$HC�5�YO�! E�
p}������H�z��D>������%�3����[�����>����GyH��a8��ٯ��h�.w�NE��m�%�Qk�VN������|��	;��d1v눕jg�������W.&�$`�v)ۤ����ߖEs";�k��O���_%�\��T��ы��s�E�^�Z��y���QJ[��I�Z�c�Sm��E���y�U�;��a�b��PS��g�F�7���U\�2��mH%���d	�Oi�*�7�)l����� �:)a���"x�)�]��n?���=*x
LM+��鎪r6�0R/;�MY1	�ԡʋ�4��1N��qST���B}����{v��1��k+j�K�3��$֠�n|(.�5��֊���*]W�Qe��~
3߮�W�f�,Q�ǎ��Mt6������R�,�C���T�J�Iڷ�NLO/���M�-^D�v��x�0�,�;��gA��/��D��4��7����+�d�Rn�ɱ�3�
�.�j9?�Ē�A�cT�B��v���}�׀��R)��
�vr?� |ҨPV���(���4v��y�U�JD��JA�A���>�"؋I��X�|�o^4U��3%�x����e/�ſ%�.�_ϸ�k����6viњ��_�Vn߻�T��T΍q�n�.���@�)�K�Kϫ�#/�o?�yn��"-�:�/��>8���
�we4��E�p)#[�P�1����E_!�-�p�����\v��K	!@�����O����ՠ9z��	^vkdԈP���{WR���p᡹��~�'����F!��;�QOW!2�C���Fb�C>@b�Ϝc�K��O����-XA�\����k�g�	??��zj�Q5�؀R8����*��bev[d2���RX��뚛��d&�7���}�	�h��y������{Z�Ԥ__�0:�X�r��$mٓDΣ�蔱�V?-M�D�[#�F.���֩�!\�l��C�����3�.WS�(�N�W�������@���@�ׁv �@X�̹Ѿq�����٭�6�q���{'y�C� ���eW��C�]��U&�A-ࣈr1����a�I��c��g"2���ΓNR;�W�x���U+�4x��<�����X k_���Bƈ���pf�X�ǡ�@6�5���>]'�lybΈ��bwL��>0)0x-�Ԡ�GD�j����_w(�f5���n5K�ьk�@}ᑒX���``k�����B���˸�'v��SO�Q�`���
�+�9��D!Y&�'��\�����@�.�Ob�E�A�	��M�E:Tf^�;49��9�ÅXA�k�J�׺�~�B�n?�'��! ��59$�����ߡ��E�
��o�9A/E��[��6?v�h�ӽ����R*J��B_g\�j�
�ϭ,��r�?�A���1��aB��5ہ�Ē1�oc(�-�56�G�jE�����?Wx����w��zA�d���L�g-Q��KNR=r~U���Jʲ|K̸P寀H�D��L����L&_�b�H�O�7g��Q��F�k-��sEW�u�0yՙ��JG�Sm�^[���<��E=�f������ �̪���E����E�����2�^Щ�����آRC���-�����&SkN����%�6�W,f�gL�Tnm��E|z�E������(��/�f�Ƽݺ�F�-�p�9��F_<����~!����q�V��>R'�:� �ݖX#����^��2$��}��_���	W��������ș��;�a��
鯯������2�J�r�$����$8��{�'��T��\�n��뛫25V��Jl<?]Q�qw����|�b�f��T��k�kH�����Zڻg$���8}��'ڙ�N,/Eh���g������@�'dLgD��	]@�'uR`|����ֶc���E��:D)�����l�c��D]����"�q.�SUku�Y]��ҁfj�t�����Fڒ�Kd��뎪0���`�AD��M�qn�z�_ԋ�g%��N�R�k���ZO���Df̬1�0��� ����D�Y�gZ�n��[��V��g�(.�+���%	28�)\B���ja)�t4�����i�����g��:�O��t�V0T{���t�+B�u�m��x�5��:����}�('�	Μ#%�6�v]�y���P`���z��Ϝf"X� N�uʥ�P���UC�̨����˙�������v�8�I�!p"2-�L�ݘ�]2!k��1NW�l��G+E�F�9��R�����V���B��!(/#+@wd}�Bg�')�U��&�W��6�%��{=� 1޴%5"�cM_�RI�,PVǠ]&����&�@����5�ǓE�aH%�Y)����V�Y�]H�]}��4��BT~n�]�,��¿�u�Vj�wY�L��tɫa[K���&��|�r�L����$�#l�μ,B+:����c�c��3´�\R��g��գ煭=e��Jt�������d�	�O�0-C����7+�4_R���Q�:sb'%zj?��&�.��?��H�_����i?�0���-YEz2gˢ\K��ZB��~ ��Bg��rF������Gט��hb��� �,d��ۘ�Sf�+����fs���������"��|�f�1�6@%m<v1v�R�W���>���Z]Gj��bDC����T8�iΑ����NC��?�G�W�Ғ��6q$(Q9�VF6m���H��/��2��<JY/4YwlD
��s�S�ɞBg�"a��V�?�	���KAt�L�g�9ج5��gn3��=u���%,S>(at�L�h,]g�9"���P{��C�O�ؤ�B5C�>)��[G��uw\d?6��{U�.��ᗌ(��d�P ƒ���R�ZNd��f��r~��u��(�КT7�{8 �;��y�YJ�)�^�o�gɑLWs�*�X|�	�e�8,������t�6Ĭ܈;R�E9�:b:��/;����o��)�H��]�ײ�������{�d��u8i
�hlH��@��7j?�Tr��{�����Fy7}H�()S%7o��V�ܸq�l��w�}���k{�:����gO�[�����WB�=���2�Dj0���3���	.�P@�z@�����f:��%�B�n�ơTa���;�U�L_��U(?�g�˔��!�����h���A���Q�4�F�nf7�2��e�$'��|�pz$�MG�o�M����%ط��:���Bf�]�ٗ�3dx�,�J�#[6i���0F欞ᰇA���+B��2�jh�$��Q��ZC��Z���)l$<4�p��Ũ�M��	�P��kA��5�f��^FK)C����m��E�~�7	��n��H5\\�l���zV��l�	0]j����xL��]��@sMr���m�h>8ô�,��l�S����E"�-��I�\��5����f�L2�P��~ˬ��1�e�J���8��������������-O�x��ݴ$�|�}��n����OW���OO,��Ed�D���l�g�]�!��Q �k�#/�_�.ߧ�!*7D���@����-2/:/�M':�{�na�8tn�-��"&k�r���n�[������}������ ��F�}�#in�qb�L�	���āG�Bf2�.����������R�ڼ�XM��⺐x#+�F��pJ���^P�ͺ�~���d��h5�������4��o;Vg>�MB������;:Q��y�O(�>�m�h��q���8��	���c,(�_� /�S�g'"`�"���/\�c8Q��J�4��"JE�+�`����+��]��Z���:�fBl�Z` 5�bo;MÛ�t�W	sN���������E�>4�B���/S��gawqsف���w&�	5���c���1�n��2��P_t#��Y����\8	�����B�w�%_xg?p��i�/چn=�,��H�~i����i)lw_O�g Uһm���k������|jO�:܍�7�����3X�u騬3RQӮ**s��}�6K����F!��v�DX��e?ʒ-/���]�	�Y �f{]�M���>��^6-׳�\��ǟ
!�ܠ��`���[�#=��z>ٳ�*Q���ԕ\�����ƹ��q�[>~���m]� Q�N��;(�5|o���2��D-���+gc�'XS_�����f�`2Ul�����pK��U�]��[y��')���p`6gl��4�IV�\�&�a�	������`49��}ЫJ�ˊ8ظ+�?��ј*�tGt���E.�W�B���$�� ��Y�K �|��n�g$�@��"m=Xm��E��ꄟN�nB���K�� k�G<�S�	�D�?��,u�8�UP����ȴ�6�2�k2�
Dcl`�oS��HBvH�`h�Z̀��s �w���rv��0u��R��g]���K�0a�z`��m�ަ?�@&���P�˓'u�x����@;� ۙ���%���em�]�
������!i��y��Z�҈��q�8���S��J��fSy�SDD����ǫ(������/\lԵ��Īgۛ�~=߶pe��5v,�Zr^��8Pε �x�L]��U< a���a�;<�/���� �<���Ǉ�H Ĉ��?���ݼI!�T}�S�24/��eZu3�s�Щ���ǥ�9��l� �7w��b�Lc���5��"�|򊎵��L��3y{�����-D��{�|8����|N�-�Ҷ+���)�e6�dlA���b�a��kG-ܩ��j�u �B=��i�ps�Y�+'��&�4�d�}��n�%���eTo��!� �S�F��'m8��b����޴2����Ӻ���$56����^�����&u��Q��.��6u#	$��`��"�1ƴ�Ɇ8Vq��+y>��,OD�N�7V��c���IQ!�Lk��P��i�γ�*����m��,��"^�sT���oD�@^^I�E6�9�a��y+���a��X����$=��dI�Q�0J��bt?���5���L�O|����æ�E�D�SW;I�pC��`(
�A�n�����݄!H��H������)K�U�~��+H��%�눳��RT�6}��~�o�0�+�x��	q_�&�����q ����fFW[r���c�g^�$�m���M/7�I�zrq�p��yգ����N
}�A2�J%#.�2�^GǭmӐ!
�&�/�'m~�e�W�N\�o�B-C��G'>�i%���J��u`䬴��)|�&.l�ڋx�h}�J��)E��1����������g�P�K����vh!f���QN�?\��ƕ�$G�A��'���0�[�WD��t��x��`۝s���^�^�����X�[����OvH�폂�+j��=ߣN�����=(�I��V6�;\	ѯ�� _��|$�����QSb �R��[�%�]sB�C=�qM�7�r�f�l�*ȵ���U�C�a��Iy�@c�lמ��$!<S�;��;���x����8�I7��y�#��_ě���wc��Z��>�Ez-��cmYY֌:�Dr/,�t�*�Z�:��XF�F����o:�bkPo�A/�E�W���{F��3�����Q��Ӳl!��VrA����b�2��ͧ	WLҤ��E*�u�;+��Q�\؍�Ulf��l��A���oC�d쓳h%m�������}��K�w����/iq��Ψx	 �X�\��Z]P��6�J�3!�v!l��3y��~w��;c�H�6D'�$�n�4Sa��IW�rx��U�Y�-k>G���޲�����;J4>��m1�̓�.}�JBB��/�3s�}�Fip���z�hzX��3��_�$��^66�þu<z�����U,��R���:�Zk���Z�n����C!�1�4�(��d���z1&��@�Q\x��AyH]PNe����@�PVZ[�uĘ!���R��aM�Cr��q��hEo8���=�{g,��%����@����Q@�g(�Ӈ�id���d!��������y�M�ے:�e<�N�Ք�<6\��J�=�o�g]H/Q-[��>������G�Z�(sO��[V�۳�%�,���	��n��i�D^{��*�u$�F�n�bv�.�֑��a'�D�E׆$S�z��"�{F߻�7�/Hv�^mߛ]��Y�&S���T�9�����#��ي��Cԣ<'� 4�Og?���2޷`>�]���eF��ڢ?~�T���xdi��$����V-sRz�f:����D?:/^�zvi���~��5Mr(>��o�dD-cz8���q��\&3e��6C�MU@��J�ʔ��R�+1��������)�)�a���n�?9�FF��>���9��>k�>�3��Pd��d���E#��a���{���'vP��ƻd���XT(�b�P��҇�7���K^oV}	o�G����[/��_ʫI�yK��)��D�|�'^��
�.w5��?$�{wd�x��G����(�Ӕ��u{#�!�"�U���x�~��ז�"tZ6�+U%g����5�6��P�`�@-l�w�n��b�m>
�3r`��-�
f*��r�#f1F�齺ۼR>�#���mȐ��ę�/A��Q��2
�cuz�Ik�cVq��Ţ�U42�x�ً��d���+eA=�[��u�k�`��H�U?Xj5,�5t�k����+hH|�ܠS�z/j�\�����)�Kc�:�S\�D�i�y���#��\zY�q�fY߷CM֏�f�y�ሀ�.�
��)0��0冀�"T��I�$U2�m k�*q'�d�\<>2�`l�d�	�Li�]J}�]B`�x���O�8��9"��`�,��B�if�O �Q�7	zn/_�y��������>�1����q���4�� S��`.d�W��� &6B�M6P��R���9[���E%��LfƖ皧ʯ?C�J]��3���%eN،��Ùy�o��q0�Q�J���ʖ)l%���)|t��R ���Yِ=����z�L>�Ҝ״԰:U�H���f��z��g�w�5��X8�?��k���l�Z����8M�?m��%#H��+�϶�ZB�)ފ�Y��CC��jj=�����:dU�a�Q2C�Fv-�,I:��rhﬞ��T��)�4;�|1��ӏ�ݩ�4<��;
��^���X.�ě�DxPT��'D�}L������ ���ݩ�`>rSp�L���a�S*&U���=�M֦TC��L��(!ǬHH=�c��Α�jU{4�Ѓ�s`�T
,U���#:Z����Nh�	*[P��x����p������
Jg�*|�\,qH�w�U�>���=��+�����?A���CVF�[��W��_,f�@r�͂{��,��1��j".��J�)b����:�.A�,����-�2�e5����f�H�T�[��4Z��� pR���[�L�x�l��b���P"����<1�q����y�rG9]�����
Ꙋ�|i�k��2|�ӽ����4�!Wy��w|��� �����uoR��h��^�X�P]uG�M�Zo�)��^b��j�;;>~s��!�p�p����tU�.�0��+����C���óR_�<F�L*wi4y�nώ8b�@i�̈́B#>p�	�B㚣��ڑ�N��6�R��8�{N��5�/E_?1�v�8ޮ��j��a,�^�,@�}_.-8����ר"����H��N/䕵�~<0�biHn���T9B�k�\00=���=��.q���m�t�g�-�����&�{Q!�RV�k�0��C/�[�v+w�>+��yk�1����	ȿê�S�bd�:	��_�y�&,J\-�J=�b���T�]{���O]+�YFa����U�	�4HA�N8�{.�DR��M/{@���%@	u�q�/	���T��W3L�~��w�X���"��4û���P߀ɇ��J���k��Hː�=|��!S!Ǎ//A�% G�IiL]vʐ��.gxם�E�T�Y�ct��t����sz�C�#te�D9��~�	g���
kU"ב�{ �	V{ ��k18v��ݼ9}σu� �<Y*��ǐ�
���StPeN|�`�S�ʧ�m1Ǹ�:���f�u��j�Gv|�(�}���w1���{f�g(�C��C��##c÷pje����<v�8�&f}�S�ں�~�tBH�jy�Z�Ū�:�,��
a���p5i��%�M�a�/i%�7��g��u�����v�w��p�'����+���9)@=�[D���b`[~�]��ة|�
q#r�Jn��j��d%5���4�*�5N\��t$cQ���x[-Jc$�V���5X�����i����iʋ�h��>+�Fo��;��kVF����U�[�QIu�����F�T�,��q]��^r���]��դ�y����Jd�����
qieg�f{i�(M�y�C5g���j��W��'�ς�U&��Ȣn jW�A���MvB>&J�$/��E���E:�J�6.�X��F��_����j��$
xk�wo�=��5�| ���"6�뜹�6,dnd	�����tT�#-+BQy���15�;�F<��\���H�09�ü>lB�i�����\�(k�;��&�q���� ��]�yx�4��Km���|�N��bs琙��ӹAx�9�ٚ�7�)�Ճ�����d@͕�H�x��IV�/q����M���VU$��!?0�.������W��y$�Yt��oT���������'�Gǿw�J��n��-kCFM:�q�pD|�*��\��Ҏ�Dpk���>*N��Ƌ�6�xqI�Ԛ���Q�����(�Jee �ځ����O[�4)z�\�h�jg��Ǩކ ��+��U �d}�7�p��n��ӉZi�W,�<�ěc�>�X�QuD>^>��񬌏�*r�N���e3�����U m�����;�r`@k�J$���0���tM��jj:y�~|�2��OB�,{}Kt��צ4���Sr��Q�2*���{�>eMe