-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I1AaTrwVKVXqVrz5hSeuLxUOZzfmjcmBTAI6zU2Mog9JoKyuD1Qv0wMtjsruf38CrIUUo0vB73b6
cW8vxtGWabpX8VNuYKbEL6fS0/qAik1l9ig2SUjnGnCUnQhtnypEbWqj6PHX8epUTuNrR0UTCnt2
hrOG02CcDFwrhtpVZ6EYDd7VMFwckqU5rwvUOQUnaQ+McyI70FvBvDaMTLQuU1PUwVsHjE9sL/k0
YLCLxgz7xuXvB49+pVssnwL2Vix3Caww5kNqx7A5K4DGFINrFT4HyN+dOE2GFprzCA4Q8kFuwKEo
Ed6Ahdi/c0gncK+fQANMVBUJx5UxVc71coAa5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
RG8yPISAH77YhMyFe24UvKBz2qpysNEzy2d8NsdE7QilmelDwJzDv9OmimYGco/1PQpq02FcIFQ4
o4F5a8kdMhMsNnvccdxc7d7vhv2NRgQFg89dFIa4lSCgAYxVtlQHaCXiWluY+z+VV0j0eWddNc6T
B2jrqY9f6ArNMUCYTorVm8baqlOUQ+YR3SMvrA6uX2K5gKf/mxa3W3gDLvJPq8BlaFk+lLfq7Inj
H7Q00snUKFscgJIHw7KQq6t07c6GhPbc0zjSLLwOluf1NDeiubzJ8p1XXaPbUsx8bvmmuO9nzklc
4QKO2gdlb1ROuvGkULPh9Ulx+cRdx5oJn/5gwzIHtTmkXblodF1iWx+VEXzX+Dj+X4gYVMXFi+dp
YOtY6XJT39lQ/u4ANy9uJo9ZOAnoA7GLGtjjVYq49jYsOQSZNz5hbcV0xgs5p5glPFnnTSB+ZxNs
fOedFIkfg8ENJ61J72+qOf3wjo9MpvWPdu8ifqBIp7/NasRX3la967xTlF5R2WGHPogfkovY4+mI
uxmk3NPm0t2udt3mxAP5Dd74Qm9SYMsgosDsxyJzVd9BL67Qv5aS5sWO4+ul4xivilk0IftDX7i7
wTcvyKZ82nrPzOfAQ9lgrGLbzug9Jk4q2QJQAD+gm7puWX1QGHplYNvEWUasEAwlbNjNMuCcpCGx
SifhgD0XpzHFG7NeZBi6LiJ1B7+mAWbx3aWIuHyIquE6kT6SV280gU//3cSqpjPxnwduSVjOzMU1
JaNu3enqqMByb9J2AKi+vbxWsRwtZt47g8A9oB3OKmMN7b6mVDgdY4cT3GSaEyyLy6xES//5lGUU
7RR23n3AY/ssCwEBXLD0vo4VJaekmNtfa2tReaRsfXyYPawEHTvp5/dKzFj2y/LKNpjUpD4RnewU
75xt/e6wF4LwWlAlvoltv5U5KdqZlqocc59KZ0orzGm32aiToIxnzyE76D3B7Z7Xyl+ANukC3IDz
AbEPMJj8yWLEHPygYAnTKgeFWQW6OdRvu6cWqIGnzOEC/I3gkOcDa1v2Y+WI/NA7WBjDFhA5q101
euBlDVByebLyvOJSKcG/9LFHk6SYSBvKSZ/50QJuwLRzKkArZWC+AFl02tyQCjYRtPXa0dc/p3og
EHMIUSg9HQLCQ+vQ7szf56LaUHQxzyHEMS5xP9/NsToXN9xJyMEqE9huLXeIICKqgXQCb9DjRWLJ
GyVHANLyyOrnyHK8e2+lbnwSafCXnowo7MWjAF8bbzVKD+pvddmO/tIWc/4rdmwEQTDI00q67Sh8
Qb3hBDnj67wnEYDBaE8d0aWYr/Pbw6YuUcXRWC8Bm4F3znQGUa/eriLIUOqi7Q3oM3jPyhzORfkN
kMzLElnDWFgDPS0HV8T0s6mhKTIONjKhe5rfSRHzR/50V4WqZlvyT5mK2tDSAj2PkgSR5vmManZK
So1xizL4nGv9swd64FwibIY4CYBLkwEyCzsSgnZhe76775w+Ax3dnqKUESN7hq39P2d/Mxahy0on
8qkqOSC2qSmKOwMekc84EgNydzBQMLByKO/vQLOYzeGo5uBFFs+3IXmFyy+bfkRylfUZrCfNYXD/
EhTPzrBGvHDEqcZtX0LSlZQKgSApvbMpoAwR62eLPAi1WN8tEVI9gzUm2JyPI6cWxEL90kKmNpF2
Y4fQzhmIgvvln4BC6YhbA2L7YoEx2WDx0N+LGitSHGHWF5xejhvbooNGM0WrrleM7EbUHJJ0GDEx
rrfRZYX7QLLpnsEVbN+ZOPFDjqRywAPHoFM+croLSIVn+rTTvJ6/TEJTqMirZoDSBOLGoPHqht78
kOQhpl7bsNvdVBSwd9sfxbclGEFftN49P2atvqm0d5+NLZOZrhleJjVtdazL+GHnJLFwppDWMysr
yLoksw9C4uNIswGirfFZkvw0NqxyZ9XeFF32AiaMk7235Q2fNAAT/q1QzFazmi0FypLX1CJ0Udar
Rl4GII96rMP8bYfd6GfZYGRzjamsGoBEeIisnzWTNnwZ4GRtnhcQKtqFAW3l3yvN4PaMg5ImMjME
/X6Q9e76tFj5Sn74UPz9e78348ZCugW5Yn2Y3tXdsHY/H1uz+fcKkNQHvcF+tyOW0KW2AwZRbmnG
UDyG3rGyjHdH4gRCU1Cg9OHFKpuVA5tRkjnSsm11c1grei2eFXX5AG1GLMOK2hfZKpyPRgui+a/Y
jrf7meOCwnCM/HjXT1J0E7neAObUINjtNGRfJPemXX1UGwsYHB0WTJoIfEdCVGpd16/XMlOR/sst
87Zxo0xwKI50MoIt4IktXZ2PPniQm2Kdl6sR/nIGcs+W9IoxYYSjW1/ue5c6zj32SumOrTB7MEEU
PcgMtpJKmxQ5gpiqKRC4GsBviEbTndqsG04xX3z3kdW8tJ/54X19DJBD1/HzPlWet4bTcBYmO3D3
SOyZECHnjmy87YnjKLmdEWoUUTRZ2e1R+g1uPZ2MbdXjnyLFSfu9rdw812BuWOiews9PA2CO76YQ
ts/kxdBjQapEGYUk1bVy+qunodSMTuoUnCKzwJ/BmQhNTCKZhvGObdwlIqKvo5amNMXBjkT6mdFt
xZTnGsr1CbJy4Yq7qmSJMDMQ71Uvu9FQZkVaaV71RegS6fR/PttsM6X6tprf/nzlfw6E97vUYBpa
n56NGOlqXFBhLk1Jn07qp2mhpvpmRzg2m0Y8JdLpzjQVUJXCA5UI6ATZX8LcOrz9M1yZJ5EO/TBV
x1qBmcbU/PX1TV8kPMmxuhZzUxvltDKMKYiq+jsg1fg3sNFnvtldyiRpptzPZYmpYorwvQsETsvV
Rh3jPY55lFVcd2zwfxpQK/5Kjr42svHn6GThN8Ug0uI8TJl2I18IwHDF5ieiBpYxmIxY94bLXZDV
jMxv7XF9yyLdQ1tXCZG8MgZptwT0wM+IBWVtcgVlErN/YntxlFSy9PPd7Bus3OF0pMVZFUXMDLCt
ZkSzkgKSr4fbMkp3f60Rm9keoxej78wBrBbopLL+J85z1Fv0nAsnl2F4TJoqtqiq3Zut5rDvsQOy
lLen/i7wVuW44N81ZDuOFAi37TEFRXxPyDEZPruIZJFFy1p5heEtlnzcEAs5bOXWT79P683EgZMA
2Y/wc4aLCIpqJ+IjyTQaTdmJQ+T58YwZNy1op84C17NSy0r0aytHbydOW1dsUz3QbffOD0JIlHVM
MjTqsvg3X4q7xL95O4UAIE+Tvfj2lrzORIY1Ef32OZKyXae/zrT+YA0/8PxjUYjUpEMjwaIlMlco
IVVmqbhdPa9ngSQTIkSBaGrC2NxM7JfgMLsDT6DZkBayH4UQ7D0SiDAJy/IpdD1c2S1Wuxm8r0it
AwLuLkBCEzV+4wJNkSkCGD8sjUq/1Qo0H8jixRJmkwUPdHlnklTQFoDVpP/7RyiyJF1opI3WgynX
M9vOjDLx5s6RXO/s5fgiHLJPcuEjBl/5aXET3aCCBpij3Ysy6U5pp812x5kae2YB9eO0ASTpEgtY
jPmJfZ9W6bj2ID/odUAqL4geh3meX9/UyVceDPSlW/KoarIkk5kFRllcUXurfiMpb07/rciEN5mm
fG7ci4AO4HUOdqaE/+vdmMOhivedqJXvdo+N7q8VfpqXhU1zJ3HkuiXPdu6NJkNiRWtMZP71X8ex
q8bYBXldQo93Ej/ppy2cB0jH7tAn/+A2Uhk68sK0Ons3M0h5PE4feWz5xGUtKqvTw8XQtPGUEyug
XLRMTBOHoTRBGDrsdOKRM6OzAqs60rvstrJsoSOMfTHdvQaBUG25a7V3gzRqNUfKjYD2XY8D5vkf
dMlf7//YVt+PqfFPYu+jWUW0Gey61QUunkpfiCNXKyHDBxVrBgcGKzDGFlDQluJc80SeRhXyCKxB
6Mj480sxWq1iCDRY9tf9Pj0nUqpj3cqHjVB8oHToqMiI9zL+bJTkCU5QY5PsNH7Ag2/VmoCk2hEf
y3M34uq8tp4rM2dgu9SvRykcQZz+oixgEKIdr4Ddt6roWZi2PY8NnN1MO+HaooUBzhFw/a8qK/w9
W9s+gYsqDj1o8H0APR5Fg17Mj1D5/E0O7KtJzYqHVOvTPpsEtQFBWdhoD7g0WunPfQSEc/zzO96b
D6dTdbntfaowkrdvNFBvAKfGv20JP7ySHockcrN4Ptr3iXIr9JeQVRolJigef2ENyIE5I0fzAg02
8RuheBo9rI69QuDq0ak1rq7NZlOaU5/yF6vhJd++YKgf1/I/0owVVTfrmNXrS5uYqVrqkR7TPZjj
0aA83aUOfq4bWRhvXy4JZzIxcRhlenf4NAdmzlOtxNIFRL+j3K/ARg6IWXqCsDBIIck1HYJbk000
AkT4zyFedNdiR9a/R6F/ioGV8XrkUuMyshw9P+NiQ9fwMcTzBdBeI4NH1iaADfNAcZbwx7JxtIPV
Y8pD2K6KwBoKgsLUPjrIL8Z1DZRgk8ClEvSv0SOw8CT/R155mn0yc3ESSaETyhChyZirjLexVkYf
hvPa1jqskwtgVnbroektJts00iXRIjZpmnl0IXUuisKQ2oow/mMLnGgCKOdbPr8lhaR4bir8tSTG
eAW5cbrT+wC1FWrg3KKh/ugvkzhoo6uH76Mx9nNDhYeSYKSdIbwC7O5VtFHSY7mFohcV0psB+ERx
ATgvvKuWhyWLWH6QgBX15hjfnQoGve+NDy9P/ZaNLpjeCfRjKgfHrTE5twm7hii7x0/bR5eqn7Fd
W5wAKM6uanaEYWSxIvWulEoDTGoLKgc+IRa0EwOg6nmF02K+C4PsG0n/SohKc1aBEF5g5aC4ozrL
UJq7BueDD4tJ+OE/5sP0FKw2Rd1SOKxF7xmJNYDo+Yn5RcgQvjKdJDkqnJT4dNmSchRpe8esJ/PB
QQk4PMUJVBWpxItB/SQfL2Y6x+yITuGG5k/ypdLgG2sitx4Iv/nNf1OcdQlop5fN+hYjIeOhAkIB
LsYdntjwujBkbL8wB90FfIFbipoHdXVy9uUSndVgWsWiB0+VHWTPk+z3WNH6vX9OSpEcO4qcvU1o
m2GKuyZHdr2VvmlS92E1yBpxRiYMUhVhKzfR9AeSRM8+DRkRRFsOCiIzLI3z+8DnYYub4g0Z3QW8
UqTyRH2Ksg6lJr1DoxgfnsgdKi5m2gDzkxQw7ifKhE3dZIpxg3Q3k5ndCL4mtghQ20MedSIVSa0s
sdjgv5KPYEzPdx8B7lNE7LBhqAFthOqJx3wUZ5McA1eGu4RT9xX4urs0sCzQoQ1V8WNrtTuCt5vb
1vgpQxDpybSobO9q5Ay8NY5brG0FkM4UEYxigHd9kDxz+MkJHmehSx+IBhwM+xsjjLd+9IX/rtId
3woRdPMge8i07S5lgDtlL+2jLCkUB5Uhu9WcNjderg0b0gdXG4Zu0Q2btpzYUWFCe9LW5qflMYOm
UfScYJxpSmctWe99c830wym8dhCGjz0MGUjB8yECtkg8kzvAcruMqRNAVYPk+XoWQIVZkka+Hpq2
SzJe2aVPZiV2wh3OwV6iaouRf161JjBB8IyKFWFTJ/nqxbvTxhg9prAP61fxKYWK8Hi5qnYwmP2D
FNm6MhMn31YPspAynLgNSszyX6+N54tm0ckfKIABmgmz9PjGeEv36+qoTx6ZDCKNCLo6gwFG2rU1
v4BwPyi198iLGUEV5ytZitHWs7WCkiEZ1RfbkG3mzUqYuarv02ZeAYLnpMSMJ4GWBDWZjiY9AAnC
34M4BzsvjNnur1AjNkokdhA/tRSQgE+7BDhQcXf4rLzzF9nWUEybbx4HxJknNpNr2A9fVNfbDYCI
OkY4DoM4V+MfuxhN0lZrQzylyZ5ei8QlqFUe9wpRUB3z5sG+YYHHWDH8psLfXtbP982HaC41TMo6
herU2WQCocqJwuwg6A9IaERLaFdkNLMg4z5ZxjMhrLLBfFOP2gCzKasF6d9Il71nv6pOHl6uGqoa
lITwWn6K8zsKU/ga3UpahBLF9TUtU6Ew2MuvWtDEmu+KeMKN7e2iLQTYaDgjdITPuaSQkpH8swbg
w2f3UYVsh3LRz8lPDZQfH8JMqtfCeGk8uTDytxBC8NnD8JSAGy8QFuhHvrUFbkIn4+WYC+tgV0NH
TkQthojGkE6WjhnjmbYJ9AK9lY24j5g9es5M1x7zUq8anW+/M1D+m2cgxqefFy8Zqh32PtN7JjzF
3pGdyAMp06tqfILupHwQl2uyeToHyqO385Zh/70V2GustPkzgLWm38xrLUio80tj9eoX6ppvN8Rl
2iugSY5U/MxapEEhkIIKje9Dp8h5on5eF4Pty+UzPpkyhh4+ckrncFrZq2xIXa+F4DkcM0CYOLuD
RvTZylhNFOfadqTFRtMN9OvGWuZKS/wSWPPtiwPO+SgNr0Q9GddTgYhoy+CZA1nQSg6igZFVaMl3
jkWIq2LEEZXgCfxYurrNVtt3xduuQNtUzdCUDVDBky7gM1xn9PV/1fYcHyyU0szQMNennAfjX7/l
F1GwxEy/TIn35HriH8fiiP3smUertsQvYOdg6VJj60eGKullSdG9G4CUnLaRGkTAaAebTZl5Sol5
Ze14jZ6S4lynYLDE4+QoahNPbb7lmqFZMyj0gwv9mukAsMzcLM7BRaqTJ0aEkgsTAL/1r9mLGAkN
buQQCV19W+Pu4QWml74RaKrDInIkh01ynVhFD0gK8eZEYhEOgIxmglEAw70T3q5iSwJofUoYv19O
CiakJDR1XKsseSP/4tv0gWPRxynZZVyNpifLKUGS0z3VcpnpKBrRj3SNy357fU5GfF1sIlA8G0Wh
TACXlTKtFSrf3FkfPUWMoDa6mQvTxM1OiBSEvLoJd7uZRBsR86obxz0V7zWAANgAJ89TrXPSTDG+
IZH8rVOni24VEvPZuSDrPgYP01FZibNRTz1kEuWOyow0ghDOunJzxwFxqR0QKGIa6c2qDL8UKPA2
MRtrssa6GzHvkZMul84EeI1f+vPWK6NkjUaXHZ3UE1Un/I1G5LwAUUpypCzG7U99nZglAtJdVmzZ
WkNQZMjQqnWp1kHAr4J8vBVQyC2Qq4q3hnxOCjYI7cjNNVlDOXLaSklqrEDjjjqf8NvWTlNqp6iS
5y2Z6UnWZnLnnXoypEa/5wC+eFMSYuJ9WMM/6GQra33p5yMzfz8+VYEU7r3zuNO5lRwoeu1tK3Pv
K6m78TFGCfRBKCSkobAyqVzaEn/bJ+LCBRAQYedZYxph7sh8WDKQWXguJEjy/YYOjE96/ua36XWs
aK9B9OM/hJ3kHpavEn7br8Geg54U4i9sbRlEg1nDQHaD1JjBAZ7i+Xf/064vo8CL4yFogVfP+8X+
IkaU3aH5a2hHlpYiHyTOJF4we2xhHH6UpGiT+rpGaLrKokkd2CvaNmX7eNZ2VMdJeFMpQgAWFP+L
OTdBDXVfH6gIAiIOGsGG1yoXBG4e2QMtYF5uCAOXeWXOK8/go+X37z7ynsbH7vAlbSocVlunyUAw
rEYq3pixExnY3/7RRL9UoMuU3Ql6ee6PLP/3mttKeUjGdO5jUoBkaG6k8zpjIXxs0Zul6UKMXuHd
XNQCqM2lBfpf0N9/BXrubRzshd2CBUC8v3alqJN3T+jw6rFW5YIhG7sa9RXMllQ7XMJslLRIxSpE
+sWcyK1M8dtGJ78TrfCFQQsT2gtD/wfip31VEApyCKXvBFz9PFE8/57XapwY9S4w5MOKS68qY6qq
gVlmCXcQrap0DB1lZ3U1SiAqjGZJfHhXa6ZsAm+HKbhLY2V9Jla99Sfhm+zwZ+9Ew6jDF5swzwL/
2ttp2/4+LTQgKwbdJZOjeX63RLDgwf37GCkKLsZJ2irWp1cul8ykeIdgfrCRStdfA1Ih8AZhlfd5
fk4m04LYOP4/NtCaT/1EHnbB1uZXWX3XEyrMzPqaWqQF2iAOPY+7GEa6wy3C3fMXOIzpk528VjnV
T9jdtEH0gW+zcP9P6tKjCFBFhVPyWtewSkrB+krVDqoOFJXSBxEyn0t6xl4Rn3RoF3Qjj5Nau0hy
P5Qr8cSGI87V6dsk7NImtDrVrgQCdnNzogHZp9BJd12LRepEqGbtpqsXu7d6gi1IM/92QUU6Ok8a
ayEM3LptDUFLBLZXbkzGMBxgq3otMMvIp0NcMoBUuf972DudhxTKLki64uRJhNvou+Jglo0OeJMD
z630Qo8dvGHcTH9/zRIPu1uyGgltj3gGcFBknktxDBqdkz04HxN48nZOn9aDv5NNzhgPfsMfsYAy
mZnI2CYoV4UMZz3uVGvdUpnJzowL9we4MYZ29m5wcx/yug/16V2L/yIkHokzJUKR9X24bL4RDs33
BkKxPxhgokE7B+nCdl+n3yVFg3OjibhM+F80ICYbHj3fzUBtqHZw6qjANRdZweq1msU7USjtMbsz
ciaujmHXLR0ToterQbgHHnTSd4RImfOA87OkY5wSo/8WYMSciOaCAKUchG/0nMa1rXBuGFuRVBbE
JY8Kf4DC7LzokRrz0r11NfP+RfSMsf9+bwp+fOjgNqCVNuwbxc4FeCMF5fc1NQBR4KUDn+Y503g+
7Bm5Yi1z0X5bRZQrJpksmA7gTQYCfBKVaAxfcqBsDixpU2pp2iVLh2P7kPC0Nwy5jot27WircpuG
3M52Dy/4C9T4Nzre6xL+tOlDJxgRdXXu3nWQLHwdQ3nfBGJPH0VqO63K7/XL89m2/WBRL/TWK/26
H1v7s+9E6cHNp+gGP5I38XVO87wZsQy7F9jDv5K0VnR0yUx8Asr3opeKaStWIwxh6R15a33yEEUx
VhAJepK7nQf10kx10m30x6AEHji61FDcwsoZtDxA4cX2jQ07EQnQxXVObO+eHLaH5a6BJHtmYrya
opmAt9cYGfiMGJ2pzb3spZH6rs5XcBnCyt9DBY/ChV/AnnrqTPEBXb1e4r6pSGYKsQFvIlgriHXJ
FLWOU6F6bxh1GS7OaGYcqLWZZjHxmsyGBgqa/PidU4CxI/q5BXDRJagK1zIszuADSf9SBlpqBcNP
5Pu68GjX+YF+xPc7ATu4oLfgAsv2pPkKSS/3JjTqiHWgi/scXlvKZ3+bZxHpkAoe0mie9+ygCx0R
gOIr9ZmdF11QAHiQ61cCd/9Q111rwXREQoUtcsrZmeAY0Z7Z9oLsspUrVucpbAcbKfu+UgsqTDkL
RQV3rFPACQtlttp/2G3OdAGsjV5sUvf18a6DfjNy7WUPoeqYau0ljyVIXDrO8uv7Ls6q0fr9KjVs
1zkSnyaXYWy0/yZzkNMVCF6QjgXrXE4cbafYyrhruoQRlM4WWz2ZCJKDjf3MO/9xqxdmwyQ28S4E
jeawIXoleMbGYmVwl1rDIjI/bZhFiRePrcY9MNUdNuSTXxOzcDjUcTLRE8BDdLLAp+vDDcGVc00H
EaxpXmw5ekBSkix+lzy4wgk6h7e9HWJ71p3PldtjXdWHCMtMMklmrsnBn5WTyNN0uaogAcmK762k
UJ3kjFf/xjTj6h/5+YKCmHLTYluOSkTGbNHR++OuPj+5VW6ssFBmzZs78VXQOFr+6diwGOKRYYEd
Y3AuFoaETrBbvxOs1eGCoxffqVlap941a3xXT2Jm55mapjdqh+sqBlZqLmwIdPJdWhZXzUE4J+cs
rHGepQwFgz23ObGmAElQaQwsHnhRedWxrf51taO4EHN4suGzReT+vWYTI3tPHjV4hJXwZqGzSXnn
Av9pRr8uFPxsD9ew+fhKrxVjRfArn1bqvlnosSFrOXM/Sv4pFAnofpvj4eAidfhhJLK7WlrPWz2h
fxVnLBQL5Kf29ORyeNuvpxpJIm46QFr4Qa38BaZCPM+HylQ7QCbySLTAnHdduIeGHT+zZ8qFWbl6
5179fZzkuW9s6o1sJ5jfJR0eS05JYO2aBjdzW30LSYyUoYPViB94lGMWlN1OTm2nx4GmFF8kK7tl
swgbK4k0xuLenzG6d7+qwjK1vMvX1pAlwoJy+LZE3LXSuCqyaKFAmOkNeKuLob6SsVaeRHZI0v7O
Lvfn0xLsa7kg/VZOl9SGqgZQGAp1HNr5m31RjtPPXoIjfG8QHvHrS7xYzl4qCroy540X2wpblGAn
ViDPLOvJGA+da5xLeRB8cFOI8vkJnPB244gaw0z+jiD5hko82lM7ckwJfGn4xi70Byn3/+qijjVl
HP2pzFZXzWoYwtupJKAJyO4a/BmtVQj7ayZqsRwD2gzAx6RWXsS8xk2EPwSzqiWosQtS3CMKaO8p
pTJEhtcK1/yqYRbDbHfskEvL5tWkucU9TpyZWJXapCTeIC74yFzSVgwsnWBW7R6JtXlBbsscYuxm
EQUNaPj5XFTAgRv4vUmpY3lHPa58TNrJnWsv5jXeMcVONyg3mx7YWlFCJywAMnfGbpLZrnrvNdJH
ab5x1Gn7Dyh5qk1UfqrjbwyFAsBfpbAFpHkfZ8nigVy8pLpJoequwwxiDx5w34dp4BoS9uwM81n8
l0ACyPdgJ6w283AJuT0FNxb9brA4qnAYw5n0I2wLDHeQe52DMr+xFpl5iGV5wxVBM3/Y/G7hXq3c
rTFDrc2Jav5IdERpoMTk7UPD3lIEJTtCKbpDHTcvRt+jKMzkip95nPcVFi/VHUnVtW907Ey7+hHj
Kip8DqheAtRGgUtSC91KSqz2WqUAPo0kqk4oZVTP6NY1aCtXWBD/4ZRxdAjCvxKXoPRUJkzxqdMu
wgR/8IqoIENVW1V6PAqkP53VEQD1cKdXYFip3meSADedex4SKvfEvAdZLOAGhRS3OKGeyWy4Q22R
xVCo+wiYVrtCne23Tuen+k7OAwc+RBFBNQ0SQe9uRj7/UkRrH7QKuTemEXUJ1aljxjXxLfEe6l9c
2QKz1sn1L9qeTwqNIB7q9iKW9aiH0qnDn/ZMSxoMNkW+Nt1iCGrAdyabDiUEThf4LOJvKbR9OIXC
g0riSKEbbFIPF3XywW/AN7G4dKh9MJRTcSSBkklJpYE2pfv0yh4CbfiBjmUQ3QvJvAYenpVhZwFw
T4c2Hb31ja6qR+auc7RSF88ZCFc1KQcTjWYipsslKZWOMaPZO3v3y/8eFblne1LHv94iFASOjp5y
tw6K3W4UJvSm3RwtbgXoCThdjoVBtwpwhtKNFvW5gBgFPZGSHQKfZjP64kIi8V3KM8EUvsy/uzja
hQNk/Ztl4A000GMBk85MjKOu29qJjADznf87UUneutG2T80grlCuqchg3Cs3K93vMlqfPde5nnNN
8/WjIh2GIA9HwKKc4n/0RX/apUVoggKakZI6Dm+7ZFUPCS0upaWWa80cRCx0HKZWB/YORifqzhFP
9Pu2ADmzuiQxA4uNQxAjAYaRqCzhP3PkScKEPEDkQS50OjIwTOLOa2X5vwijAqRB7AU9jL6cwhz0
ZmakH8vWpqD2Ek0IakjwINVE5HNsfvnsJydQdfL6PB1A4OWNabTzN1SAO5q+rhZZ2TXGXpxLB6lb
DCp7YdrTHpHflAK95AqO4syMJ8MQASXDKWVuzmWhJayjL+oHAv5zQTPcU0zlC5JfU2ZIBkwnA+wQ
KHzLjWtGOkUCeilBYeLZuSUJzRUL16HMP2GSSN/cf9UD5P2SagB0kB3ljLHDfW5V1yzF9Eumjl0s
g7fsxGUW9jl/VjmUdcW42VtOn6env8nfMFKlpAzbqLsChsGSClmR4887Trjkt3NWcsHAbAEJIA6w
Wd1B8o6bUL5U5FlH2IxJgqXpjHoX/Y0x44XVTG4ewU2k2nSik+WJJXTNHiQcNVYsSpO2fqHD0Gq7
sQe9nK30e1Y2TzSd/XGTOVLnRr2r40Bn0Qw/UboAeEvzKcQYKpVd5AzICRXMn/AARQQWCIhJCuXx
tp5eWpvl4AHpXf6KzV44O4RaH3bBMK5oLdCbkc2i/L9tfLunk+YlwKxO5glSn35ZkfSXPrU37uvi
Y79kzoGJLwSow4LnqT9g4nVvoVuegi417EEzUuIx253nZ4WpmSjpmUHNVNhd5pms6X6KRfklaGzq
9y6EKQ7gfNKyKx6tKNduDm2eY677iMF3iBsTEpFrAz96VwbIwXReupYete3Wqh95klAELMmvfN/C
BctzFSfA8ikMxWXMnyNPVKywXOpPYT4f+hZbshGpVXZBFlhbf7K18PtkS7y+HhysOA/iF8exMBe+
GjHFJMXQH37/bLFRvJX5dy2fa+XEMusBwyh68u3bOJzNW7f/SVHA0NwkwugPyoUhN9eyOtcC7OjZ
IIBeTDc6Tluz49jR54tEsSpdFYDzWPMjU4e4K4m3IZhsrOenNRYpziAGa08zfoxmItilajochSNw
J2Vo04ba76O37OdEH0T2JostqnGPG6eSbHIAwzC4UWRulnHPzQzmHGJ3WnF3gZi5ArhSlallT6Lj
O3QGPQXAAo4mf1608EzLJhJg70eHM21bHpfa57kGFwBdox/qiwDWHpbKspReQ/M8ntSrsX2otVQO
oUoaOUkxmXsIAUAXlttMDP43JCwWY2+VMy7cHlzMifE4WJjnA/6BcywI9bRm9uLYQvTdNvt3dRvv
moMif/TmeT23q5jF9rQCe7yWlTIKL/OBZeJw4U2hBhjHEXQW0X3vJCVVJAdGwv0Y8OYk6GTicQVZ
KdBQoNj0PLfG7a/uYxrIEv5TM4I8zkTla4deHqc13Ouq2GZEPMvxylYincmAvXn/BsfDQVugZZGk
KDwTgJKiGysAeKaUHaex88JmOaarTxs1rVd05Lk31hnfnXp0k5JR+X4F5OF6+2Gv/uuT/XMUjHFW
9zZdGJVYjFKtm+ugWh5zu38fjZlu1QS9f1U3m2EmQF0w59f+Io158rJNkeE5i1d9pNR7hzO2ZW83
LZ3lo45QV9m8ACm7ck91uRZzRAknjMrhNQ04g9zklA9z4Wco9AroIUUVsPusuCh0TCrI/MTs8yZW
EePmP9H08TrDn9M+Tj2/Rvwhj8aqHGEzDCMhAVggTSFaw5N2596v69+SHA1P9pTPp22mGWyFBa5v
OgdeXxq94fv/tYmIAhJtLDyTd1Xti60GEs98BF3qwP/VDwXHbsoMiqqr/7aqFe5CZgrNClI/1dM9
SidndwHwrJggQ+RWXjb5Xb4nvipojmgbGUmFErE8NDszkBYB7us2fi631EOKim8dK0B8pX5tAxxE
zhZpKLbioQhAYEzUa9ZpsTNjCHwQRhgvJgwzbvy8BThlqWf6fq3IOCOzDVtVkRWZdehWMOjts3dn
qebSCo7LaWq03EJyHfEjAFf1E7jDd7hT281Nmk1/lueFqUgfAkrLIFeIjW78ToNDKHs3dtnHr5Rf
lOrNAU4uKoQTmdJSUSzIDqfXmc5H8JQRjwiHB1F3c3BErMgm/3JPyZSs/ZTaiQ93fWvnJMz7VOhp
+brfaOaHxmRYEJ/eVtNV7wwmkWxoKS6Kg60nnxM3lpdCU8SdRTWILir3vDESg2BDC5jh6aQIDt0k
d5poqiZAIcZ+EAX0qlYL0e6rc6wb0pTXaoJx8R99wctB7gr9xuRxKidi0XOerYgIdEm4MgAN8EOc
pWMfJkobhkrzzlc+GRzxybjgHaV9sK7Po+DTMv/0X8TrRmlpm1+6qdLKS3TBMztoVGOH27OPIJwP
usshnT9tI4F/8BrkBFt6HbASsuCVyUS6be/x4i5hW2fNGeNrmj8UZ1f1kzbaXnJXpvUawPw8s/zD
K3FMB/wAviLZN0dkGSsj5qVsXGHauVmkdHv0qhwXDny6m+0XL5EJ1xMWh5TWXxDh+FZSEoNxnY1R
FRfNq7HS6frmvKWwYZBJtT10jcZtULOFx5ckgrgIfIaariTGbV1sZI7KULL0bVelPb0YGUjJFh+N
Tg3bZUWBe+PBhgDIA2mIraxEW8Px5vLVhwATz9RVBXpnEix2aG/Ovzs+tiXtLnqz1IjpWAV+SSTK
4TPfZD3NuK2pYEwvfXLd1X+MuDXIAncQuDv7vkkZH7hllyATes1oqAnYKNpE/bYgYbIAVOyFRFz0
uHh6uJJgVc3/GjAQpFfxsVCl6zAUHw1DNO6xryacmvQ2AVDtE6Ig66q/UyzHWJWEhjvbCMMueLbQ
LkZwDImrmw2D8k8UbupEAPorMUYpUfmAhUbNbzdB0SU/6p3khF0i3pdheLhzM/9HIVH75YJM4/BY
tFG+rrXlQD7ehbZ8gSGz0FH+OHuDkw1n0vBljiBLUGzaOrquxz2h+Kx4jLw6N1yMdebvbkUaER4Q
2R1B0tJfBOTe9M/ElRrg57fspqrL/gh/5AUb46Fae3VyOAEepc8zrFC5o6vjGkvqIXixUzmCFpSF
n+1KhADt8nILLf+om1rBLx4I1Z8xpxaeF7SFewj6kI/ZZJX1yHw+bLOm7G2dpOlqmyZKR1kpQ/GK
uKQ4nytaR8UJ27eg+9NyIXsXV9bWF6gonud1ivNOEu2G9kH7Y0DkhowSecqajocWBIrwuVrLaf8v
srIOPd400QcTceyq/ooJFFOgwwN7pj17IFzOrLA3YJ3SDb1XBkFz0F5P2rjtIiexmB2ApxOtZSPl
OaEibYbg4TT8TT2nooobYkIJyU0I/B4GcN62pRw05i3DQhWwCCSkB1KDB/yylpHbzq5/B2wDyQX9
s8Ds94PRXPtVyDQP+Dwx/BJY++Yy2oynCQD6IyJQRKxz0nVhmyZccNrNu4doTOymbG1RW10iiL+D
ahkJ8k0aLhDxiNrM7+GplmXag7hPp2LdwpHy8fldee30jujiXFtJsExA4eouum/zKvQGZ5oK92ps
tPRSS7XPNbm9Tl7EgH6IhZ/pUpl7G9Hap1b0OBKMNZY0D/XxeKkeLw+/EKBOPYgBAbvMnVCH8hnW
KPJHPkWd/1PQGtqZcXonmW8zchRYArkrn2iPtMgkZ5QGrTYfy1kRl+OVH+i939bDTi/pq6KU87f8
1z9ZmCM3sPaiyG3wzqUwdV8A5O6IZwG2diYSlL8qbeHs1E1+bNIvKrvrUQZkoQyJjs+d7t6460cF
Q+ordx86WCy3/PMs8Tse+WDrHKp+sCbXVABmT4c49utLQ8+q+RwE21lwa4bSI82U7M27olOqK4gN
HAE3R3noT2fIw2+kpLbKT8RwFuYee1blvgkkNSUsTN6bexe75oC13IdflARWL302cKO13a8h8Gsx
sUJGeMXBUrIGqjTovdBxBlYmP6Am7uBHbP1y7I8xzNB9BofuqADOInTzAptRv8iKZq2OAmKlAPUd
KDo20zXzlqU1UV2BXXncDT0cwzIYb9IaGSg3afScWvWS/HXU1wuFKYoDje9gyHKv6eMMYSWkHp8S
cAr/PLUZxpp8NbV8gDTmb5yfiUb4j4mq3EyjbR5Aa1wEOjLepYHItQXMzICr1RWN6a4SWp8p/IBK
QfvHLhl+7dAw06+ChzAgtfRqT4wRwejrwZyDfLGwZyhnE/OexDmepcVHXEvJJ0pNR8zZcNC9oALB
YC+B7HV+syfByCXf8vMdB6n3ItKBr1/0yCsoMEtUjX/Wi47h0cING0hIQ0O+aPsKpVfXWREJXG2h
F6RLXVeE5rdItuK46YiJKFqDpcB13kZUTThkMednUPCJN0s+6j7ViFtHo4vq1vop8X8fAEFFARlL
afMVLTzGw+6ekFiwRj64+yCCpzKK/QwSTWln+DK6pPzbnn0t75iyO/Px2ysqL7ITLHCKGcwn7HJU
aaBWA79sOQ/lY3SKSabUbGhixbyVCpuWFT7CVZ1xLLFuV+86b6GjowUHWF2V/jcmNGWIofPscmxC
cqKMFCQs+axEDAKJzGjDQscSA5uDIBCKosCo3haQDWZR6vTQrs38aBjqxNaywVRY4PHQwkQ0rh8u
2Ih/3TWvlGJT0mJwtSOFSr8V11nYoLzaGdLuFPYqRXKxTBjWDBsrDCtFw2CrNCrmbv/U5StNo/nY
hSz7bAzrHu5+fIf2TOFyenBMRc8Bjtwx05x/4afYzstDTGvxrwkHWzrcaSpuQ1RrsKeHDpOz9S8y
319oIrnyQc/UOejGCkz8LIwyMuHFrCz9fOj3k7KEf986GoV7jVc3GNJrJQw9y0YC1NtYIjBIv18E
XIpLKQBxlAAkUuIdkJkrvnDHF/XVTz8v3nNx5w2T+YDrzREDdwGu42XiXCY5M411kkTMADAp+6Ik
b8AABviUh9urVLyT7QaGMewZUCMBk+H9nqcnSTtkusmXnc2cqy1sGC3vbnCTDb9xCEbWciPQcZ9K
WpQ3MX1o3vQFRblNRRzJKxkVCXM8GOIMfXn8x23te62Nr4uuUgb8r0iYdABByUkjddqM5C3nQGJi
9RiHkBUPUmJG0tFpIBe/26jLw765cPAU8JFA93FVPJXbO5w5w+0Bxgi8m+Chk2mY4LEDQcM56U95
8fhrFF9vWweDcobqNSZR/zx7LoJXgRiYRCEDueWZ86Id9jRZcgC/VQrC9c4koz71MKSsJ0PoXOrS
XgqU3uZ2U3bCmaqCytU7zxesU6gqbzuf5jwvlImuQxf3ci8+1ZV1F8TWIp6gPZoYLZkcZnw+Jxsn
Oo5JutBR2sSujmhk1OrBAj09at5wYRIhZikWrVG7HSezGaChINmAeXWFgpOCCB5nXohrPYVxf2fz
IEY6gSj/QtALCy8Zp2catohBlup1nDj0MfAgj0XYGIfD+4j10ZHdfIiVLe3HKNULJWukhCqaKFSz
yoF3AWBwg+AhWlc9lXSgZ0AU1KX5QV9lrYca+O5tSDrn8DpgMLkMZFCm/htoJ7S0vFB73LL7sCU7
nXg3I/BeYotW+e3nxcn9dKJIIL+PzjkkRfiZaExF+W7KD1FLgejT/AmKpbLF38deuHRM89tKTYXW
+/i3mVU3IFbVtC2Tg432xep3DxuU3AyCh2tfIZZnpHODPFL0wwqRY/G455xaceichgIsg8REfLlv
el8gcO+wpt+kfHtN+xZ9P9VOLz3ieW2vAF3LLxEJ+TKaMAI+SV6eKOrPkGHdthgirlYIo2ZbshjE
NH28JWkmF4oEBwn50nE6lyx5Y6R2ylMSfsVn1Ga8kHirMGVZf6WFFaGkQQ/+yppYQ48qbV3YWukL
TxuelKvS6JvzboftlsWtXgwujwnOopXbcoZv572eErDz5BzGYEtKI9ChvuWNnXabacsvsjNsYwD4
wtf78VGPFpv8rS6zHHaGdcVx8w4LpKMWo3p9zKOamSZyb6BoHST7JEMu/br+QhtNY06qheYHdgoV
A+V/6HxDz7qw5YSXNzAaV5/rj72qBfUJELiLpPil3SCMLdzZnpuaO9k4tw+zjLLAdiAXn38k65jq
3a2EnuLJxVyB6pF1DMKdBCC3kAYp4l5BPFMZPwkN2lOuDSxJsczq+vl5d1lajznygD8OT1kZ5p4a
jarwDZUjow81TolWJ/k1ErGhmcTFaxNZ0vG3lbvA4Fg/7m7ZF7npGCYr4naBvL9fi5JEuMyAPzhK
t+CBraR8Wr6Prz2yz8+fEXswP/cUmEmAn/yUnVhvvlMUJnY0LrV0/CHvWATOOV0bXSSYxAnAWEPQ
M6SxdwlUMHH4/VNS5fsKGvEb06TutxTaJK9byDcjsREMADOXuplp2M3MCkzFpCnKJ7oyCXdCPgso
xVTSucKlKcrIBf4MuohMud0bJCsQQDr0Hgu5ZNDqXMUZjoKbm9ZyTg2ZbKRFGCwhMCoxIJjwTP7q
oV9SauAB40CQF0DQFbPwr/4rMMIokEExAp4/VhdVZGceFbQBC5vYXYx05muEpvPml3OpE/abMW6N
NmJTv6XtgRviQ6lGb5UMp7/jDLSvwuZlDWdUCEyIvW+2lTeGeJ6uuOolTWPdamre1cttkr0idMiM
eofYHOKDskwEU+zBuFgSGqyMkobSkwgc3sc+uMesDdBwWPGHdXfH0lhNpUV2JFtclsIrj2oZ34SN
dGJr9S+XIhAqzKOF82A3L5K9nhnhLY1yw2puZAUYfvWdwdMf9hWYkXWnFzKPkWfNAbWSrUFOz5ZA
rEClCtxjtq9ep+hcFuYtoA6fovaSspg21q7DqzVVXJ54ttNlH7LHYEqCSrGq3NtTbT4rjNz9jtlt
93pmxJQ94TpB9PEVmnF+3YKcLTbypkRqZ83aYyTERRYCg+jduEVZCp62kO+aZG+SEBfg4zLJoldK
su/m6lqoknZ6HW4OGlF1ZZxzmGbrL74FAZ5vZM+LqpgxmJ9a3zG6e7QNyTdohO30V35UCAbdmTiz
+ULE4JGATnEEe2FwfYcR/BqGYBY2U9NPfHiNtHcJFm2PXlB7t4NO0RlsdkYnxInNqz7Dd3q1QWST
0Wbcn8BlxaVZoeeGUXeOlmDLpMNHGYf7Mcp0/ZKojLG1UQj/aGWfY2QkGt+h2VaFir68eVtkAExX
8PGGUR3/41m4raDq+Sdn2/6t7jyY0/VI7sfC9I97iy8TxIFnnGeVzkkws8FI31KTUuwFDtmriW5N
nif9E5Snn5hh0lR6g3CB4oq9LqhU6n1pQh5p8dAlKcdKX7DY8YdcN8Tf329CUzGEFdNf7mfo3npj
2EY7waSP9wAAuCDcLOVLhr59VjcdQ/cTFiaPA9OpIBKHRPpcOQdhF9RFMmKiaWSmvN1jTOPsJjwa
clOzLA5ywGZUM0f5F91I3ZC1BBLDbAu2haOhyexdR2KAnqTLtK4zV3nGA+EmcvUYXlFRcdCsEbQV
8AZ43hBvk5JGiFOafyEBkJ+9E4t9+Ebm77sGK+Dzkpe2KWmTFW7TOeexeW2CV9KU98mTWVUQVJBf
zbH0N8laUYo7gJ9viCXZpFpKMmPdFVUEom1T6gpIaurPwc3v9s7jpJTU7JO93NP8SvWDsAg6oxCO
jF1iYecX3t5p8brBMmCFMFU1M1mDAKZ1o+xwDpAF+bftLwcwKZxH/GVy6xP2Uwa9aZ4A1H+DJIlE
EgTWbfDmnLJpQ9cmXkaNBEwsCi4eBhRdm+X1iUL6djQ41LE2tPGImRrrhpEW78kkrbmsiE6apOJc
OcQmwKWkdp8GvWTKOoC/7tQl9130CzbjlpzYgEQgjBr+0owIiMgPLv+tvJgrX2JzOKPvzbwmjiSA
uMRDB0TG/s3r2TuTy0dISi67h+JsmntvZZFxjdtwepN1r6X23xrDmrs0LP249mL5gE7FKm4YJCOc
JO93MUG/+I+/C4vNEyu4aLmI2qqCA5TbR4rjc5rTJufuKZPVOFV6W5ITrDpHucca0K8JaVvNrp7e
ILB3fnKdsRn3b8y2+kC2Qsj0LD6c9PPozPbd/CeleSUq8fY62vouNKHdCaYRodDVyADtCxKQ0RjF
Wi0zG83osT+fseERy6i1GAFXRRD8noxElUksDuT1CDSVEvEqUobHMBZ2EYQdk9HOcfIl8ir5Lkba
m3yhBeTMQ+os1xegi/uH7/b3ZyTrbpQ/qASamhLNtz3ogk5/s32IFZHvVwmMLk5X9zW41syE0FXQ
SLyR+1STqVqpSgpqflXGYHG8wSE1TW91sB04bkj1r3mxkds9Ib9+LAjVx9uHhHX7vlMIB6fg7O/H
eb3AFL+uSfBmTQlXRivwkff8sAaOHoDH1vmGVI77naTzUs2zOkhOpFVonGHuHo7tafbFTs7uVkJN
Y2meC0l3qfGHxLdh9GcEm5j9oaFiC1y+9XKYkxwbyubWrCVXTmliS3baM7RpdbKYfLJ76yTzIwjE
ARKksBX8mTE20nsuxWlr0um8RVELrSP2LqufmyoIgJDUeHGKn/MFCVn9iV77+OtZOlVowlWsQ9Ya
Bm/JhCEIb/IL5FjwiirQyHjCBBiBjF6MIupM3lpapQsQUyA4EmVLor4YUYCLPliMRcjyWky8f+7s
o1IgZDXDXUO2mM7JzAEX+J4iiatasBVue9FNZ07Bd6YtISWOSFq3WV+9qxwVLceTuzVT+laReQJk
y74+RDvSSOKobhMk3gNOdV3PCw+NebIU0F/uo5tRvhWfM+h7frrN2OPmp8gC4HsrJQTBbTVNeI8C
X4S1Mcrkpl935m6kqU3T6VzRVk13BbKMlEypUZOgRblZNs4Ex2FxRbvKGhAoqRyADeH2CqDxJsH6
oFidZjDH+cOdp6a43rh3fgLyMmMDKxUJbv7Z4eaxwylRfYUHZA4xixcasjTMDjqjrwBo+O3yeCjQ
bCwyV/EeeEgTcrU5ohk4WUoCRx5iIJeWiT/zicdgBMtwOQWgi8ihWiNkHnNs/xDfjwnMktmbcGTq
/lxqMVpZo6RQkFD9nByzlVa1l8tZ7X3q5Go7Bw6VKJV8UGhLQY+kcwvTv2zXdAbbru29HoizNPBT
fNO+FelsU4hsBQ6FgjwNv+34V3s2PutyvsLx8muL6hYnlpOJJfPrhYjceUOQBwHkhs26YGkSB6dt
pnuPekj838sF6goj9ZFPdAv1YGKT4k8dMazdkGTGrzvyrwZ+lZ8CtvLXToLDl0BpB9Yr02MXUI47
U0EfcYdaLwHuPWSisD7LIZWG3R3KYPbR5hdmucTOqpOyJ584J5q9Q7n1GfO3DzbpdEAAdZJKCKpi
fZME82mLQTJzbZ5y+he1gswqzxkd4vcjSjw6LcPo+aO6q9xhMeVnl6z+Uydbvvnx17kHuS/grUo9
IU4YvnIQdD9AVzILEw/1f1TERg26AYWibMXGVZf30jsw4/RvLleomvqS5gVUHFhtHFjg/iODkn2o
TzHuLddgD0HcwmmY5s36PCwaekDr3+u0YICls/NxNdrruKzEHULuDgyK8SGh0j/Imgh9I8YDgbu3
07D+nLAWDCUAOU7//nw1qPF5mXLqJ7YskBzCp+jdX737ac7BdIhK8AplB7rwG1muSYFF0QXtbjP3
Y/slXy6PU8kjRMz72ekGnyYBH4s1mgcGiZbDGM/Y9nSyMckZNzOdXoQTzrqwIjoo1s3PnYlh2ytt
wApQx5F/dF0EH8TaqHLGkEhmrRdRNFXbYQLQGGo3rkbzerg4vlYsk1ZnHtll7XNCvqtjUd6tckyR
zFEEBHWIuqDQBtuR+IX7hyIgkXyOv3FpKbNKVe94peJdkofwIPZwjMPGupvsA47uic8jsPZXbtQ/
apf9d2T43Hwuo5oNdviCiSO0X8vb1zqIzP3dKLQi3WKbSkwCWhgJydXNH5dwYOC9oQeGV0bcnwsT
BgkxzX4jrQrS5LG1su8oaW785cVtCptkXoXzMa+MynZrnTC5U+tVV8H/iB0GDfUG1Tl9cAZoKlGW
mRRPDGVUqOtHGQbUB8PD9E7CF7WioMRXpChsSybJCOAS8gQp0KB+ypJAbGnjyKHOLmrTuwnB5MxZ
zixfcGMmuIFKGAF94ydBe7mI4wtFkdfz+HvOoHoC2mtRKsa1Z1r7bRW7PqkO1lLMMLTlS6t6NYZc
FyQHLDk2XIiPG/qrne0YBVj9Pp12uJxVzg+Q6idYIWLDc4YMxzjG72X013A7fSlPkYNuTsMLfN8e
maRijRhm0henGrFBnHWsjhbNU0ONGQn5gWoApgQzVmfqusYzSnGJsqNRyXDpjg2LAwBvbtbRJeV5
pUjB6US6BUj1Y/2XS+SBEjIXxikm5gTRR8SbS9RjrhTFofj7XK8iecCvsc1PUqoJcXEM9E4u/0Pf
1capXPTSwQVcaMgAf11qWodTK5mvDNYns+SA598fCzs3DgXwzMm0UBPe9NFwYmZwN6cw2wSTc09+
71GhwrkACUiFZvwAjCRYxdrrtQc2nDk67jHV3D6p2Z6+X7delkRK6qYWmzWHanrS8GobqjI4ATsx
3q9IvbdUkIpNB/opT+dl0VurPEKVYgFf7Jf0SmWmPFpe3BiiIYD6mZ/z+CWD0z/47CcbaiF3sHDY
p3uXGn2/eq0MvLgoLyfg5oZTsGSYnh39cdpOzpFMJnAESjRYBwQ2WmLv6tiqNtQR7UaXVqH1Rfd/
bHaGWkBhMGs+LjrHNSXUR8qhko3LeLy8qAB/gJBtHFbnpSdKFLudNI8DVswMyZPuv/e6Zz7RFcnQ
80lqfJB9dkacyWvkK6bWXNfVMcrvlA76UuFGSt4k92wBYZ6dpADGN1Mujk24cmXVKVNszmejDRIz
GKdPctTP/bEYrWP4P5X344MJ3zz50SSRtxmyhlRWmlmq+fcdDDn1029AnroUpu1pe/yLQgrv6V/q
6FVVXv0stDQfE20lE8McogzDGrC5nq4jtIIZrSY2/Yh4+n9IcVhBP6xmvK13vbQMBhYbUacCxAhD
jIqKDdpGDm9mtm9qxhPDgVWcQUBg2jA4/grxM2JGTZACtKk0X5KsDsuCCesZMvaVWdjmaE7muoW4
S3iAFMiCz9Gf1kPHRpwqy0DT+fn2XwXIYpE7kSxp/GTRlS5kiCIG3TzlYGDUBwSj3Ql8W4NTGQI4
of0Rh+0YJu2J7zQTpIMyG8Y5Uz2fxSWMu3cTp2xsBLezPltsvrVtApQeQqdAB8liyjvpioBTfR3F
0+zDuCFxeEv6xK2d5AdYRQKjhigsV2Z7pmjYLL52OtSBptDsvywMDQ710dki2Imn05d5eC282j/j
1RC7a/JTN5URNC0JQjNHoF5GlfFJKCr7rP24B/7NPdQiZSXJBMB7wmbGKz3zZSVnun6P8jdep+xn
1l4iiahngQ0crg4rwfA5Pdf9WG2iXklLDiRwanVT4tLv889ySePdY4I3FOZU7SLwmURqhnXreKXV
z07y0Edf3XTAtjPyACskmfdkriJQFLYY2ru3DpkiDHONtK0HXb12R4YsPQKrCWRdgatcn3oV4Mzh
3oENteIcThxzlo57lImHFvVwcOGgN+XApQLbjApBdXR6k/WIElhvkuXjPdZCObIQs4RXKLoFe5Fv
LDDvPDslQ91pS7HMdrHU2A6WiGi2/uqdXV+aVH5gDIbPyJbKCrwB00LUG8J6dF9uQZz3W2pLbgpv
4tYgxCgOnbr1TVnPVoKCqe3KMrosqBYlNsbEQnotIFuPCQCicmptLQ0kH/IGy39ovgh+mvCNBxKQ
kCe31Zu1nZ2u8BlhQ753+HlokreP2vIFMYUV/1WIRs8D3OQ4NTT62kv+8OlGJchmNvLUHjfbdCUP
60UqpuqGReAo5mZeKnkWHJjoKiWXJNlUTJYTPdTlkBwOD3WGpIabyXLXgF9E1SbcmBhlIHcT2Qu3
BPeV224VTo8t4liLz8nt+kOBCNWxgPAwm2ShvaSYY1Dw/yqFcqcrvVhvKEqRe07rTHkQRSwMPaDG
LFRQrutTlEFnGrZui74HZuwayjeH15e2CMkECGrtQWWtW/PKJXDB6jaLCMyI+VsfvlaWEjgcRXg4
Ib2EvVXX2zjNBEK/TOivJOP5XG4io8aP3LnYUC3RsScufgiqNjKf5k0l8ANewKFwlYG7QJkbycOW
QDGLAsrwgwZPCLlgDU/BN8Z8ZOeokqzbcYCUB/m5e1wWOpyDMFUi89oj3DvzyTTby2UoldAtoOTS
XRuVwRaDcpflUpTdxcgX4qx0GI23VMOkmxRmC1Br6fF4p29LqZdKrLZrjz1d6hbQ5RNGK7+p0i3a
Sfa9cQ2s1LJwUPajLegmjDiXsb8qx5T1MXLGqyXKRSHUJ5WdOlxi1jWzXMD5DczmQq5cALsr8GHR
3Y+yq6p+5TAYH7whBbobtCZqQUVGswmBrEI+kKfGs80iGw2vqk9et8BC+6bakW5Y8iIPpjd8teAh
WiIfr65o5uoCI9goRQfqlFbL8lFVb1kXf9yXeNSsgVlJwENZkh4lEbX4L72h0Lze7IPb72eGYGae
Bif35y6leblXtjx7SZJDCRgqWFo43W27pbv1k8OLBYQd/n24oDEKkPjzhn3qzPKGcZUsS/lDhEeR
REaS0cLUSiNqGlCgaXzBUuDAC20cjr/8ZZGoUXtUwN5R8UW39aJuQriEo8cmUfQ3KMB7Q1CmpToq
eY1M1UKAStAHe5E/jej1bwzPkFZlB1EUAshOzQNz6oJqDebvJ3SUr5BWNfWe8dIm1sLWdaCseOR5
9neeymamJSzodCb77GlwkYmPsuU8DpdIWQZW/jPK3roHuxtIAmaN1pK8MMW35DiYr8UpIUZmmup9
tm9jJtxRHSqNKUkErWszIW4VdHZYcPG9sb0j06JdPtO5oZrVz7mTpTOhZXDayI8Bxtqqrui5NtYS
h5x2MkJ4pX0fe5MzEEeBm4uM2+gGe7KSZ2a7FVQWqAuU1QMEAsvTzfMyw0FeZKjbrhu7QkXZAklb
tCb8yNjWXwkWZE9B+Z/yWySFC81BInhm7bY5AFauQyWrMtDMP9+tBqZFU5HyGG+bB65nhsSfM12e
p73OsxQA2+pt1HLJVSnTavKOkZfPO8rNddrlKGqyBfUw8CaJvGHsmuFqzpJ40lt5Hg3N1w4W9yxc
bO3ZATspG5hvUyBFmbZ8H/vOMYgpk71npCUE9EPbkcbrv5Nkc8k3PHDDQpGvyaa21QQ8N6/PGtDx
GVaWl8wTZryFZoT0NLZRetfpkmbrgdxrmDOqktdEOuZKHiJc/u7v6RC4m51vRbxnTFmBrjJsOYVo
vBzKMbmdchHa4t5Yd2JsNCPgKZOsJDiUZB0NSPU/NYWqiSVdtfTiagJ59tIudOjZAjWX7YzNbCaS
OkoMgPKfbLr+kUhrP03tnwfXmbJZ0XPh+tr1J4C/0Pk+7Ky50kq/Bdoo9QQ21T0ZxywtxuJEO1jx
Z9r7xnASK/Zkke3TiIOhEyBI5N8Gx0GqIRjcNXbJ6Qk/18BbRSe1i2EXVrraJfjSAAVRUrTkUgPW
FdNeA50WFD5w8r1mwFzvkdKLWhegBxQIyOaaIad6cdpUyVVYQXb1e6eBRyUZ5C2zYMm1LeznBnNf
fq55+cNBPHoj+NZv5xalMn1pIJRM3dRT3xfR+HC/yBnpt9M75+ysJiSPtG2oYdjlZV3hVz58Bpaj
7n1w8zyHSiDzVe3CZ+wpHOLnPnkbDLyS7O90JmrVaxyAo5cqxqo6qpwFuBTWci+zayXAPlbaCdNz
eVIX8SLUJB2+1TGJD9jO8cNaoQ29GjcqSZO7xsE/9huQSmXoCCeqQqizNqiQ6nptjm1QTwWWdhNG
Jg+624D4aQtev/FSIz+XWtV80AjE/IaE/6yrxUitEgEp2ziPfl9o1YdhXsQ8tYJu1Z5qtu1Kkt3m
8hYukoFop0H+CNIPe5ZMqE7IH0u+oYtqjjK5g04Mx8mXSI5UdUBcehp4UGzZ3vv6cp2+MkMjj0bt
JFGJUUodnVS8F/R6tXFslQthhljEaOZ8Tc//gxpQZzky6JorKj1USqsXMnH13UUl8sXOZDLtjzlc
ihr2rmtrnu5wJAUaeduvIcgHT28Gdj8TxYhH/3i/q+o+rga3uKBtgIXcvWCs0vxNGOwmNTFhlL3B
+gAzuoDDsJj2j8YSgVbFkFpK+jVH7GIiZiPqdn4c58GQQDPv0frfkITRjcCAtWvo/xt3h1waw9+B
+Pv+SRpB+1r0dTBTq0ZDsI9+LP3sa3ovOLLyJtxilVpfMDdgONXLMTdZJPMpiNAt8IsR5ehka0EC
MhxyzDrktaT05Z13JRCo4aNmoJTq4ot8FK7e6Bz9elgajBKpxnGRhBlnbHLFJegosv5k9FUHL3ko
iS721GY9wGTbe/11PoUqJBDYfDepoGrJ47/u6uIw8lJAVkzSXmVYCBUpGbM1nhJdREeF16Y8Z3PM
6nUigu6SNZ42Zt3HwXyg+iw6NmgL8BcWVBrzB1efvXv1TTojUeOHBMdztePZFxl/mj3McUzoUOMo
yzeeTiS4tcKz25u+ky2hlu4i27OxxGHHFPrDGSPM6RqRNp3V6ZyKKO3JtVeEXPYPWri46t/YFIJu
BzHAIU2eP9Wx/ZnfoZdatOGqFJIwGPwozuo8/PsaXQESpxUoxIL8BSYH7hhF08jI0EAVabj/K1Z1
3WqoJAvcILRG5G26odAO0xyASLq98Rx0C/Mgss9qhdc2U61b4NLpT/DBTltYD8bmNzKEBoKpQ126
lf5z/EnbdZ91hAIDop1g3RgMJ9ea8yOOhEj0vhdLRc1ZE/+SaKuk+kMcmmTN729R6obV7kon0ycr
bFbdb8HTOH9cQaDu3ZnGCvx7xPVt7Mj2n2ktZF8HIsISXNzkQWsLM17OWuiJHmstkd4lGJZS/aun
eWuHfNDn13o6uTwfsd3zsA8WcvihakZIUw/OH42bTrdDnv7yYJpe6kTVn872yTNANCos0cMCzEVE
iXSu5u9zNevZVWziKGfh84D4M5bkwSankMTYYAAmqaAvE/c9Tl+MigWqBiUy+3ViUhIw72kCtbFt
UJCM26p4pjcT9qwAIgD59gPKuQ8MgI2XY3z59eGLyP4/JCrYSbm2kf5Oip7/ODaBeklfkua0h9re
h6oZO/Sr5nK6VQGJlmPmWaSa6m9xysOR7rOyGGt5LsdC9wA8CinK/8/PaMOzIeuEaS8/cv6oz/e0
YHnA/j0EwRLGyE6rGxCkxK2/jVonRx38ZGz2bkW3G0asDivlsw/QWcS5pV6dkyfg83O8vDMRBDfJ
EDVELINApLILh7ZaeXdEwDh45LKnfYqhthoVnML6gENhKRttjwi4zdW9WwDxrsICbhm9jQUpssPz
N8NpXS9yGdv5MG4JLm1LxcHhjYzbofGPfhzNVMSwWB/c7zb3U5TneHg0wqAkHPmEttg1IkeTEraw
Xg8AqiBoZKOGjZafWrNQLve1I6FreWw2Du+sJCfAOWIYadzeVDbFEikjwp04fbzueOPheVfn9mBp
R0IwBXo+19Sc/yYtAWKkBlv2iHbvTb8SHvotvilovlqetwqZOHmUDzdCc7HEUlWvsYIUKQijIt/Q
3SHB2G/6Z00p9EEMQTVEnyWYDRAGuweKgHdEeZOgZ1JEDWkdUExOaALji+rsB5YweFO+YEEQPSAo
GX7FBwbzAP5KsX3SVXhUIAoH/z8Lkk7PwgFcdPR6r5GlviN7woC1a22IaAWcfwpgnGhCShbFwAFG
iYbTvPYRLH/CYJSi1sLY4NbltHjJCF8rbSwRBKavgUNA1MIT4pvZrBNW7H3HhBlXcNO6Yo0UaWp1
14D7oUuE3fK1ny8L0odAaaXz3C2xxnMTCQmaf6BTZ7FUFcggtT/TYrZjWv4kcmFynQMsKtMafEDR
ZKNpbLi0tvl2gWtsQp7ZMZCIZiFvrZzdGnIVkUFATjBxSblH0yImwns7wa1BPrLT6A1WWxlXpZdZ
Kwi0NU+HLCBTfM3oQmFaYFnnR3hJkrjw/sp+VSHXESGKbrEMXMTbDcJJhcKHzbuSzBCvt5Raej78
F5MCrvWxkmjXU/97Bz5NzjLU0VzMgQKlflWw9S8plIgFjj444bg5bUKcr4Gv7HpbN/PfDpJlHPzN
M/hNnJ0yNZB6wVYyS9klv+i/T3MDjmY+Qc5Z7C9pLaCfedyyKN5Y8TDmRD6BZJ4r1dvVWUaevaci
k6PNbrAkyLzvHKgc+Fgh9S5gON93QRqpNUdHuu0H/WUaIkPDp5jlRVVeyQwB2fLhlipWaVKSjVrP
BEA3Pu0uP3QKC9CCJh9mE9PB5zzTmZQU6aaonbXJdo520VBN5zGvxU6leflxkZ3vsp029G/s6RPS
XveLlZWzGNS0YEJxu2CI6io5Q7fHR7PLn5ciYT+ljE6Q1zVjcmtuiz3E1MD//lniRnddDMVwguDc
9IUnFvYPx/os3PdCFgqK5fnG/w8zOMZycAyjb7JB9w2WxTFddLeyJ+apt4DrIWnK+lrTRj3h725X
YFwbObo0S58qJ1HC9C2b4lTIO4pzGRoic4myU//PQukrO17WeQOybUVrplv+bK/XC2dpIIuu8CfL
D1jW0Fi1fmWS7IIoxZDiPwJ3EVIt3AVFswLR7OOHWGHeqpI/ay239oEOU3MKITFfKw2zcwXV8ZUL
bdzC5vET8TVhM+W/IOXCZXKHZz6GJnnn6tpOb/Cw4mSskVOA6cHPyuvsJo1OBlGfBhOdEeJ5Hwtg
gkkLOIGfQEVmEem5ihwLVrFy1h3edk5QSZolcG4nqFoYEF8bMr5rv0UVn/RDN/LXU74jrmfl/wCb
V09+03H5rhgDb+E1n75hAWBUiIm3AuUqrxARpbbu4SW++0teBGgoGKDyY20l26BQfDhpAmZUfWvh
+RayV/mnY0X7cKZcDB9+qjaIPGemg1tmR4vYY5CmSDsYu+XFtmSX7HAl0H2Bn8iUof0TQcSTlhjf
2znf7Ynng8SvfZzpcK33HqVkmqmS8BweZQu5LNPcX/M3JdMUc/Z+hWU1wuxvkBpt53iZv4KAJ+Jx
2dlratPbzsFvJPp1FWV9WzA8i8Jks8uT5dnkSq1vQfvPFy6SV9RfYhxiBV1z7MHa9EyAko/4XPfn
BGn2jG0pLVW1l819MKF2JiyyNJJBsmoCf9Q3MNgnSCNGURLuH/rfeyyORqtqsltSgNA69SRvja8b
/s94wZrDSht//VZ+RPPP1ArSW9sA5XN7SCt/G6NCinoyyBufiQ4jUCJ51Clacvpp40/tOV6ygGtI
/VOYA6yuxYDJyX6eibCOt6Mb8+RUMmAn1HvqNmZEXqrM2bl8DsL95UUHw8G9xUXNQ8qEB1uNgvkr
Ivpm/96iTxvgb4Q50sDxMY5VDBIEuBuEqANLYrYrTFmGu5ZCA3l6AWbWdZgTxcnlrLcr9L+fOYp5
RjuNaHsbLjrdmWnSj4IJcLGQ791dbcJRfcle5HeftoUSeKPoEpYcrw8P2KHsybqw9soeQFpvsFCF
eOTltiXg5Js09Urqe2NN/OuFS7HxAxRHyVjWYx/ecZU8iglUj2pWggDAaCxlbUgQus+f3Tf1bdAs
6UaUl00BpV8Z2Ghka0uPP7h3J10uXf5k3vomSIV7wx17SfkSWVXuIh9GFpVA/MA4HRpwqzVLvmkt
DbkEdZ23394JnO/ouEc5T76m7atjEg5Q6miwenUUwkkkX3FXfUMTltAvc6eu/md7ZX4ME8jQOriI
zf6H+f3CdjZY1tFs9Bo0OgnseQJupXFKwooUDBLL185LR+ObzU2D1haIV5Rpc4DUnqrpAabxMhKa
mQau61u/ZQ84hXOv5Jj8hDr6wJO2m4BgqdFUE/HTEMnuDH+GVzsLJCEfliulhECi18QQj0QzoU4T
NLdidDPdasC+69oi4K6tO+jEnIO7eHMR5uqTDw8/kJq0qnR+lM9VXW3aIUXFahDmX4FaZMs0X1KZ
CgyZJIQANdwKaBMln4iewJb9XTYL6TnruHs2UzaEMhMkLD5IPG2Y6+X2gsRMIctra/RgvbLln5zl
DDT2FsvQUOsp1pJdlKUBydFgAnRtHLKaayln7F4ERk8eZSa2q54cLoJXYUL5MTSYrmwmT1n1iJon
o/Rly6WkPw1FOvgR7jXF2huClqKnQR9usVKpYfABXIszcS7TbYCbzFSS2S7Qu4U6baqY/HNu9/xT
TixU1MGrcp4iQiBF/Gn1Ea9AMzFr3Uzw96RJ4/M1HC8eqkF9k1VVaIpV0UDwTt/uYez20pjRWhWl
UzYT7On/68XCnRA2IVq2hvFuPX8x28S0NC/VY/UUYkVa40k1h4UqzowE74S/mSiI5wttI6IJQjnr
FtozsmY88dqM3otGvbI++Y9gd6GxKb4FaJp83xYJBkYoUrckRfz3H4HNtdoOBG+VCLZnz7Hw+blg
4/PI32/mR5gat+UHq4hXIECFsQOb/GtLPVtOMWENiqup0SDZqHn2B91ymKzUNS0D+LBYgHWEnBvi
8Z5UxOqbfBBjCbp49/GtWh0jGB6yzgAYY23PkEGC2Aq40AKLXMylSYWQODMoaDfKE2h7o2jBemIY
8IDiDR+tIwYaZkSlOBRA7D26OwHurNZUxz+JJm9uKzO2uoyUQED/dDEE/BGq51iYOMb4q+0kKmHY
Vg0Ad1hJiNEmdBQwoDhGakcO0dqAshh90TmOThSycy53aj3w9n4dOFk0zagAcDLVbDLygjfkaTP7
EU0KGuyt9kgcTwBfXSz11vDE/REe74BGX2ajObUA6n94MrLzDsM2Aa5tsSdTC3w7ECLvRgEv8T4Z
mRTuEAanZd0/W2eLpIuEe1fk4f4fnJaGbISSNoQ7veqxQXg5kvxM7KcOkGO1oHzrJVnhxBpOerWi
zm80qgOeZhPTFespXI080nil6gRU/TixXI0w+mY4EaYMiek+pLDoEMxyJ+tOykBAq8LJOH5Yx+Fl
TJIgV6SOVw7LVHOwR3qjPP1jG637SflHhdW+WdASgef3YDcddDF75A9LvyEreDVDwsItU0Nt1ViG
fQOohJFafXUvoLr/tIgDOtTbQEZi3k37OOU6imLSqJSQm/OD6IrFrqv0t1b69bhAK+xQGrGhzYbd
8A6ye69I2PQ6xSOg/Hqn/2OLIa6UR3PbyykfEkkRhgwROHcAJ8M0iuCeHoS6FV9nZacExRQWWHMU
Kl/2TWGrX8VLMfkS2OF3QfCfGtgczr3JXeAztekILFsIWdcAL9FWm8ZFrVDac5feLXciH4FmnRdZ
qIesyqOk/gID8dsjSJ0niDfm+HBufHsgHfvfLnkik9Vu7KU7q9D+WxqV+P3akLxCktZnF0+D/OTN
TmS+Kf97KDx1VB3FObSS8u5+/448n9hxn+bqXgyb1g4xpXCe1ACeZ6zR+4WEdFrMqEumh6jZu1sm
+GXAX6/y480MwpQf6Kklbejxl5H79E2giDWkzKz0FKN08eOH1dRH4W9gkAWBNeH/9G9tpgZFb3mS
KDJ8MkKuRARTHTaP9gbE+W3UfzO5txWJkVYDAfa1hNSSjrpU8ucE6/lcuuIaB5xGwSUbJT/bmnNQ
ou99XTAl1yvmS7u4svAUtsfNe2mXJqRCRUDAbv/r8PNxviV7xULCIZWdIXQhU0bc9ge2KK21aJUN
VxNwIGfhccQ4nkpnibuGrms2hKwU5wsX4uS2/5aXOpg38grL/rpcCrqZ1N1XsAo2A2zQQeLR1ddg
gTsYni3oYSE3UgN8HTuhK348R778k0Yc43/wRWT2MPYgl9PLLyVc7uEZfHtQdATC0uu6bdtSXdHc
veGiFHgCxlK+oPruJIX1e0FXYOZnzQR/f2nzBB4L44mxnUHEyJqpUBKO393Roaw05FTFczV8T9cF
ikGgCfiu3BR9GP1COM7ID9JnByFEuZK3PU+wOOq+drEbPvBirLI2uqas7tOt4bukNRdTdFVkKf5o
cYPeDe2XfY5y0y9kqfceA9VSLpHDz1lO5fBvcVtbXyIXmNY2NUZAjjoJ7/dPLknYe7mcj6aQ4z3q
rujS5wtKRh08VT7I/HxIkwccGaVVovVT3y0J2mgy62WmvHk9/IDFPjPjC6YMW6r6M5UtsQTOF+XI
boTbHx2gcdK4O2S3nXFtpp/F7vHLWONmtg04QdrpsiR3uiPrxTOVK9ntJP9muoCvPdUsXrO6s5EO
uYKQnM3Y71NxB0RFUcZDORBxL5BSWNYIODSSAD7atHMk09F9DZ7Nkf4Q10pYboOE9eulcTItyk22
+n2zS2W0MfVuLulmW3g4ta0RJPCo7kD+L8z8dh3MiID5VJI25TcmP3dBk43uTJIUEnJ203pB7Rr6
ng4DbZE4/PHhU3xD/Ayo9JiV5Jv1pFkMrUdgMkHGT+T3tr5skp75qAXhzbLVodjKWyf1ox2o56O4
AWFXTvpneMieLylYq3OxXzJcddAV63lmLkWsiddO8QMEHfGLCPW00cOIgk/8SCKkgDy9VzDykYNQ
uzt8hIZBiKcYXTfgCBMUr895yX9PDTwzcDzmWVh6CorPytO4AVSXH/3/JYFzZWiqffVV2KVu7rvl
FmCYuMExLK6qpDaWS/gIjZNe9GyL1yND6zsVdICp1VLi3FR8h3+wqXIIrswbhrWALKWYcFA24Qhh
Dg7+6qnliZhPndAQXqmn0VsZSvcAL9Hw1qrrBl6cGX/y1d66j9uTOHq2Iojap2j9U2qSJTAJHSth
0FlYao35CQCYpLVtA3DSkWgvLhXQdMNC4AJuPZGQljjbZPe6Bc4JS/4kUtHrNF5USSj77GByRCl9
m86KQ0hq0OojQEUm5LvQQ3MJGwXwYCB5o61ecWcFE5zqvKnqCaM4znMtwdbrpT/UroV03JPVJn7x
VwvSD/xgLkjVPGLKu26xzwit/IuuknZ0P1I1LGsq55XvQFMupzQ/mKO62grV7/Nmq2W7sK46sFoE
pq766IqRv98vCbLsxTbLqnczQuhkURtZVyc+wFz254+6/B/+p8Bx1ucfKq+LWJMr80mkDQv1P4z1
oucX9klkrOfwzYD2ylWf/zgWrYTYY1agsQabmZZeBKtJag9ilrXWhM1BER35VqF1tYkQ9ZyJ79WP
DFdfEbocuJKm7LKKgPeyPmpiatjAzOUuO6vBfLHBRrXEVduoDFMEhSn36JtL9n5HSBypIfx1VdtC
PynYsA37d3bEmvcdYNjriCm63nOv+ml7YrT5kgCQGwr24+hFzF2wqiMfBfLRfH0Xgo+RirUVKXwi
1bBUQa6a8unwi+Vf7yQw9rPuH7KVrB8XzOav+f7bOYaXfQ/1EeVNTrdVkRWnHC1in1NGxPKXLvdE
gMW25y1l8iJOllO1/LpNs7BS5ex6Q/urSwcGqPBkoKgC3joH8W0Wja2NL/IEAwWRh6Ts8dsrHi0g
ZKCQa31/RfWF+kCypTKbhwltSAWY6Q9r48TFlT1hQNUP6m+umS8XdDGYypfEpzXBxxkcrNqO4Qa/
oArZSZt3Y/8OyJb4KYmrh9DJHwjwAejNOM7hM3TJ126UIyQ1w0oWRC+KBKxm7GjG2cB8h7pLAJ+D
aaSZyKsSkxFw91QeQCVxTzhMbuRfMZT1BVZ5PNqsaP7ufALWErMlJPG8AphkRCyYcU2eYgb0FJuU
2bKpfvnLbBHx13M9H1FqeTSagcduGk1/cc9NRy8Pw6TzAoCjZAP+ThIv+MutS3+DUngbIVsfQi1o
rjx1tb5y00/twD5nPcWe8Np2XGRdcmyfDIjSHZNwYLnKMTxO52+5VnQAcd1cbAK69ISacko3uiiB
oamkNwlD2eGFZJFLa2mZtkjtwqxaZB09NM+mnrrbC/p49nVMJ/PdIG5oudpgisGkjnD61ORIrwcB
c1ZWwkZZBkvEeJV/4njRTKZGpGW9wvhHc8LQXB+Zdx41NWp2oqfVHKoFa2Dysc/O5zzFCgzUOPlz
aj8MY4aAKvglh8LmKiYfNe4ZUHvhGrrDCtJlLWoUfyWUb9XFEwXf0Zw5HXaSkiAOIe6z/Xyzth67
uo0RxE6gGJ9j9cbrrYsgtosw1lkT9b3mq+m2zj6h7ztlStIn24qUn7bJHAya+Jdbtgn3H65ZlI0U
15KUA6xe52vplmtK+27d015gNcyNQi/u3Vvr6Ho0ZndEnR1rvW8bCCSCgTfBn6bVIh8xe4Bxj3Kj
WmF1Bxi8WtundCrelBjWOR/y5Yvvfx67cNkqM3pYNCP5Ha/AssK1hrMvbMId0S1u1PMh24HZvM7P
B72Yh+XdZLi66zp3jumBNE/0Db27wNj1sLTmHZsXJc73PLHQly0Ru5F8LGijUyKwA1ME8kSw9SPY
F1jUTypciApqv9KELPmiAI5Gdr6Wt4YQaBn6jT7XqsH9VrbVHSD+gevflgP3n5/ESEDTEBWcrFDP
bIro5b+XbkTPKMjKkgk1ci6oCTU9eNUHBEX+fy3BQLnXvrcJME+OYtF2SpXeJqjAjyOFjFllU5NE
mSm1GBfi0aRCvbQquD+1e1XfrklkWZ5oAHasGO4Amxps4JIiNtilgT4pBFNGbiwKvV3V70QpJV5T
C6aeDoMH9EOccw7nVO/wdnFSxWPs42S0A4h6lZFGU85Bg0j+7yItfUvpS5QOOiN0aD0b/bWUVxGU
CRMdFKABHK/Vh8QzKkjNIUEzS3G7hBV2bHnBgtaG2rlmQqxq+uyMQpTfwzmsvHyGhaWiMy/9q/O7
g5ppWKtJaSf9+SavtSKM+iI7wDuEmt86Aag/c7YRgT9eC/9cNbS67WVofi2JIImt800wu6VmcKbS
T6IqNTIExy2Z7ITghCApKehrEwjcfOOKtnGHNg0ZaSvUYB9iEl4QJfUaC5fYl0bw3o+RMlbdj2cp
fl1JPVvZ9blLKb5Td0JTKKpJPZjRFY8Uuslq5+cnmUjXI02HSgFKWGv4Apceu6Zi9ipz80tN6wFm
TKJPe8IXkB/09/eMHLqFQhVCyOZM0ekruQXdCmQ9uABh1dC50TqfaKUT8poBtBo4boJswaEpOcxV
XAtJ+QRwy1qDpMAjIYBDX6WzejjvhUi+YTYFeA5bYNDVKrz49lJM/UcXJjsc8ejGubH+L7ieMKLC
7mOmd1dkLbfeF8HuZFhBK48agjLSCtUEAF7iKk0jQdhN7A+Hnx41E3ZJlHLJ9AmBg77gEhoihptA
1z3zH4QC+PE9WCvziTEPIC58WFo7iu9TC4RT2oLUq6GVRewO2rZwnnQy4GGiqEo4rSmk6WdJlUUr
Jpiv6uzQK+FYjAwcSH7vHrhkXa368Lgp5zxA26fyDMewsFfNHp4Ftw8tjyiyqTaG1kyTJYRbPrvE
x9MXUad4yYhDdC1FRG9klNiVdw84E4orLuUToFrg0X7PEBu26YFCoXyDlgBSFxyTliyoo1Qcf4w3
2SCRqAMF4IZSPTLoKtCgow+2nSu1m7DL0ktDXVSFv/4STldnt/2DHt9FoSXMAwaH0KP9lMQWRRHn
U+Y2J2RoeF26tHLKX8TjroLbvIV8XyR0/Uoad5DddcsHYdW/Ddlgybi8dJeBng3GtZg5AOvpBjnf
Zy6zpDYZGmIfjzYvRXH23Si/wNbSGhFM3WV5d67NfJqWve2q17wutZtaD8UpmWWWZFgwo1ggbeT4
JWERnhqe2ub/6VEDeUhxU976kT1+/z744n7qpm4KWTB3KISvFuDaszEAsJgOPDL4awzkih8A/bQG
3BuFd13PRQkdlG0jXZ/Pq5TpVq/qzt70OXIxxTB1JpFeBrCF8EjWhYmNsjLnViBDkiD6nUlOoDAS
TM+BXQVrIVbR38Kr7ZL7L3mfSPM26pCmV7CMTb6rjE7IUcdIj2T9m0+97TGaeL7cDvqkWUdGi/Sy
L5bScYEZRoEi5/kztBm0smfHcEJ/4Tq4amFq4pc3Ab6btrT+qyW+YgybFoEULkrykxQZAZH8EBK8
ZhkfQb4ZECfTBDrUt5ky61t6L1WgSkRfV04bLP58GJQ9r/YJN5erJb04wZNlF5fPOj/M1/q4q8BG
Bjnqn7rHIPRVj6zXRTfq+TmHEZmLDvwI+5EHAkFsBGcDsyVQvcWMgPsL0it7SUmM1azhClpgSNes
r/aSzYuTW5fg2XFpKrrUobVEHkstZWEl/6RN8JLLXFxUSrKzO17qW+YcYiL53rBGtei/P0XP0MC3
g788871F9vPja3vaQn2/o2wOZGK1M/yLUKnIr1q1bVrxbZDrEZXQSQRYsN1s84xv7+OEvuJnBKuv
29cG3mNfjXDxr5aofUgI2NGP+9cVPCAUPS15hx28jtM9Ba/KuOC+T5+19mDHIJLwypyIQcVEnDms
t105kBMbaf36atXxaBXHWVRSx93R9RE9xX7IOYDkVajbErUPfGpUbw+zWrcwRG4i27ZD/Y2vRKUl
RdhXfQLbmqltyd0NuLgTFmMY/vnvRTY+zRlxpol3hyjOMz8mqrq2Lg8Ikd2AeWa7LMiSMLUQNR3W
MExxX+949KhW44W2cvzdH6IJe3tfL1caDL/QcBrHIFdjQJTpBGJwEhw5FCi3kytjLQQDHl0qExpa
BiqwvY7N/w5FdBw+ltf2rqKCMyOPl+KcQ0aveCI3sJ1deDgJ3udk4FqMP3TWzJVSQcCUPKqRBkUp
G1Qjp7aLom9S0UzKWepNTYOKxIe3U2tXy9gozdOp1cZ8I58w22lSr5I5Zfmj2rgGaJVsQJkDxy/w
TE9CAdGvM9HKZsP8OorDSt1fpMtGPCNAm2rrDxB0fZxj2tolj0FIh9Lh5csOlKxAmlt9n45Asw9+
UuKtMCyxyqdihed9pIc/ByxfnQYKu2USn2EtJFiegb9U9JV3GGnlyRI1X5M/4z5cvu449fzReQhc
Et/wxVIBT8uDScUI65BLVF2gtZmIvz62qxz9b4CH8ous9Z4JKGOhjtS35j0XaZ3Y/pSUZWz/ta2m
6wrNBsp2tf8eNnH7J7SPuFhg+kIhHlzyuyPu3b8HzDBo7RPQT9IxZ01VMQN6g8F+yf/M7mW+BMkb
gbSdmQ+PMk2pNdS9pWAKubAlyHc1QiPvIWl8Yp4TXIQyhu6sTs+tRoCnTQcUvpFGqr7pSqgptsZO
VfhBJEC3B8IPaJcbrM+J8rrCTw3BZlmBMp9tSFqWuTrAumOpUbgZ56LBl68AKtIc0/HMkDjFV3pP
LSpVzvGmutM0jJ8pT30FILo1b73NhLZIcVjhOneBSZi3vlUVsGtCVgeJb8bdxr0o41kWW2hUK6kH
08qnzdb9cxfXb9BHGpcqIYSh/SmDmbi3PHcYPFkj+QvScjUSbHGI4w1wRz0I3/IKnn0aG0LNeDKR
tyF2i1d9iVk0Io9sPYGqB8I1WhzYlc7Efdup36Ysa0XX9I8pt8GVOa07sBNkc+e+zMGQ7mRu3AVy
I9Yn95qjJ6pzEkIVRVuQDXg1JmE0dzNr6K8Cz5ZDwKEiKcCia7u5OI8AEXqXCSA/1OrvbL/Myrdy
u+f8DqStewPUBNQWVorrcWsCV3oJBQbLwumj3H/Eh6QMhQQiaZIQWfO9hZRWndPq8T8LoYQ+yuIs
HXnpxAnwnkAxJZWAfBvagYpa7IcCmdrcmc2y06m2E/7vUYFvF3Wc6sycO7G2fEUp47nRgHifpcfG
djyJF6uHYP8U8yBFCob9ZEQ02jsHjd/zLJau1NayNbjcJPAeOKHWla9TLQmpj5kfizNS99btlT5d
7Icy9/oxKJQpREFQh0hT6YLCMgeW1NZDLz2KJX/0eBjzxuJnTbG+Yp5iro1fFROhKLTghP+igMEs
c8DwOMVZ0IgQPxpZm156zLdtSN/hGGuEDe7ju6pQ9kPiotgY3OB8DChb6BrXFkqYnm7HHStDgBMu
dgY8NLZQzS3o13fvXq+5jqJOvGVycSQK9HYskCeVZOpcJvM/TlgZh0FicYpe8iyrS21ITeNuHSbx
9Yy+E2BBkRovoE91ZyunaIjCon6UlwsAMfzXWUqRyVzqcqK6Zkg5rJ9nlbXHjj40UbzJt367f/bY
WF6RnCNBXwvNYTadZd+eB5VMKKXjCYMmGHit2+KXk0B1PgYRV4DBgstPoba+QnILUHUFHM2WGY1i
2ffEBMTm+7kkfucRzorRR26PDL/VuV+NExtxGzc5z/ii3G6etlg/cz3oR7hyh35/CRqsBm2GBjeW
OnWVOAZ9nUhEffSUelri6mG1FuWxotoqqHopQve9ppb6MrBxSYlhD+n6yh+Gx9O5wnry3s+1ZO3A
3rXkTo+iZNgPEfJq24+9VkJmJJosdDHRr1c4sgoEV8HjS2Jzv08MGvFfCoXZlguddE20SGVbOrpY
dyT++I+VeV8fq0wwKZ/GB6b0C9OcCpLtiAM2Vk9i7fqGyRlpFS5blc91M7vus1laLkawrt2w3iby
aWKPxtAAWyvLT5ZiXS/WoAvDzjJmNKIZhjv2NCjzTM1Q8XEsNHkiFMkRH+Zz7gG5UxVyK8Sw3DDW
gjlBSQLYcYuLPv7hcRD/m8ef1iKHa/fMKuZZYQjlvBJZgNHQicov+Dj0Wz6uC+lFqJ+eOpoFo7KC
uShgh82LKr77hxKiUNGV7gyy2c/NnQtdOON/9dYEFvQvWH9Ffk5Tm7IugxbxhSUK8RiwZUSxPe7e
KoNzA8OrVvovtHM/fDb8JZD/ZaCVfkN4a+JeaxX6Dvz3fLY9N0CQ/+GLhcIQRAaVjJEWhmBGnzek
Lz1CgmYJbmyj0wJWEGk2XatDfm9e0Xn+vVmUVH8LMM9wsWynrnrSBl5I+H/cENSfCH6YC6d8dFo6
eQ4XsDWKCi+/RVIPhVJVPdlZic0sQCoW3lxZtSMC8YX8s9btc7KohBo0ycu6r6lHHoOQ6YWCIaH2
Rnc12OgaGUyjUFDztHMvhh4ybD19gjt5hYRJPbH24qCOwls5RjdDARp1B6abO2aK1WaUGI6fu4gl
0NzW0lzSJmVgpHRpbwtGxrs5J4M0xyKCE+e4OhDTu70YYdgNHd6orJKGyF6iC31snaCCFit4KBh4
TVhXNLXrbgeJEMRdoRGp1FZY0BVsoAZ1W6MQYcD6GzIyMPoAiJa8s1cIdLRi0CRFW25Kn1IBnUaV
tdcXc8wChp/Rle9CWlP/12fOcHSQMWKBXs7I9h/hav6YV5whMCgxBOpDzNZ2i81Q5ad702+eLVRO
l7ANIipmJENuZBTlDksomLXwOn7I9DF7FFk35P7Le54gntObGlc/Vpb8ooERE3Phjw4I+i247ROp
dvKLajoZ++u0KSAu3aM/R5yT7QrySeARIwz3TKMDBM4HOYQzpCWHoTzimX0pv+VraEEP2KYnQHfc
NT5lmux+yTUJV1PmyqOjZYWy9aBnBMaZMVBVDIiqZ0YqwoS4LCSFe64y3oTrx2NQOt7o1JZUelKM
Kq+TgPCoPS+dY80ThAowSIZ9QuA2JSYtNdTCqLpdr8bPKGKyCoGMD3UlULv+pJgVTfeR9WG+3WKI
pFyFDoU13mVF3NdWXn8XAuqh4mloII55l/hR9RJ71sjGBjIt+Ta7dg9vslxSzIgVT2vgNpmWboXh
rbO6C0iVak6wWct2bizu2X5qg2g2iJZ2VMs3lQwrakfzUlVudNe/IUmLzUBaKU8W1Mo7v9FVYib8
PQtt48wUvSUDMeklNNOwxJprK3AvrovDVYCYr5JugfM1h+DR8fQGczCH1yz7tjqdBtNb6yzorfc2
tKz07WK38bG2q5T8ZGrK7DyCoKmXYKjWtkInUJdBeS7rgAmlBwU5G3m5ZHUquHj8kjKfn+R5uuLw
INB0FwEagVADbQ2lAEtvSgiEaBqoednn/EHa1VJrRLuGNRlf28kRi/cciIBgVDUcbFvj1wmo3efF
1AEFB0WjDftil+PU9jwh/TlC0kb8suRF1CEC2BZEwhmYrl4JPnE/TY35CeIOCmbrk7nIyb2PU8ws
Rb1eRjsOo4+SrLD1WP0TuHFvubHXr1r7Wc4X1D51nXfQ1v/XPjFatEpqQeS8fEuHVAdqwH/fZiIh
oOf6SQFR0MI5IBJFzUrGBlGWvl9Q8i9O9wRXz7soG0H+AILqG5iGEMhe50MXDf+tZnBKifsEIBlo
TCYojGEpv2ZKzzHgA7uF1045WUHRmz9NS29cMV51h2lDvTLjh+F9hDlgn4HKjR3gDKt397iI/5C/
2ky5Iw49Pn6lXLUvkeTn1BoaukVIS48ncBFt3hnp8XKB0w/P/F/Q8w+AHK7fRpiG5lvD6y2zf+/e
/FoCobUwJ2lAdpDYqLQD6aPMxgoDFunwciSZeujMxMWy/pFcHJksQ6YCnsW2mucuIbzAiYaxr2ir
9zmzmIUf94MnSvN9hBME5bF9Q7I67xwMPZYcXH+S9lq9D9hzwxBjGICuAP8BMihsiewPTZooNeLk
Kxk4yYZstYwNWkwAJjrHsYXEg98paWPtUylRH/6e/ZKDnatCGol7GOBJPAZNF94ubTIrXnGDwqxo
s30bu0HyV74gcn14iDCvAxh1ND+j+hrLay2AtRBu7FesxITe/zaoxxU1jzyCaige4qnf4kTVVlXh
eDsQpbeuIlGiNhMLJA/qPzm8SngcnLzPoLr87Qu5bgClqSGjdT71E2zq3D5ioJCcyoAFv0KjdO2S
pTwRZeb03oehQUXwz7jzeYKDzZbyrgMuEGlf0z+v9yskA78zGV5c/gZPuU2nfGZp7E62geGiKMte
60pWQyBVwoDILG6MzORVVpJghJZNNrDV2qb7Z5dJlhsNhrzEBJnsKYdt6PFQBLThyL0lisO0f/lT
EiolUsBS6nJ31UPFCyzD7Er8JUJCzTMwnLLisdoeDnJwNlXFWB7Uiny+ZrnXQsMjA5qCCH/wBlHm
Vun0nStSgurxmN2LMvyyl62JQw5yGzj8fKrxLPhpeP5Y4xBL5xMVkDl8pWncuqpIETdvpskk0wrj
lDUsXgFvNELeOa70QeLIwxqTR/lLEWeiymP/yjwGzW+OKAZBIJYldVWhCBFz2hb6bPSYOituT6rq
XzAigyQkJPkwQj3JGMbz4PkTjfKJjaSdiDkaxmLWOAffzufLzfoEfgBle6P6PVHKnt0o1EePwJ1b
MsS/c0w1QUWmdoLBPxendBNtkYQJRgDl5o2IZqq/vIWg4HX75BkviChwa3UTncn6pIr+Gh55255s
PFOGQcI15lGpul2HJ1sPEbV0RkU+PfLDbrW/8J+eNuhLw5jG2PzP+IVebnEggigZSayxxdBGE4c9
ScCYIoUkEn82EIiMm/YYwX/zvu5lNpVlEk1HfBZ7kMGISHNEy/SHpV3nSlTX7Wu5pbgRZVL+g01R
q1p/lDCZsq4Pol29qMA1bDFKGcQxhjmADInLSlntpiOs9YMREEDtI0hloQuyMkOmUQkKAoVgLyD7
GQm7LvBJmGbdQpIRjxHGMvX/jZyZ0gtUlr8fWWRFwRZt9IWBVYfrXEe2artUZKvjMeuep+la4qlh
8pPIIslvzi8H/kZ4oRkV923VYQn4gUVBxacs+g4OFH/G58y7RYTdUcMI4oOmQ7JS/N8x/bKmdiE2
cD6D0KqmIoG0soAEv4yIN09kBrJ45l8lND33kY7c1fz/OtgS9ibD1zui5EDV9IRkeZy+XYx5ye2e
d4doTyAGl3SIbxseKn2qi24pd00KxsMjmz0z3CAriqQjYEHQbBODjx1eMkLdhnFH65wb/0SkWmMl
HgZOK7BBL2VJ/m+SDjuvDTvryhun0OKFigw+GQCToL+6BvSFgZneY/xV/d58X4hypeo9vB+PUlRV
er9nELrozsYM4EAPVF59+PZGbiQUl2/qnKf4qCzJQLZ2LnHBkor1jiuOvbBJNhFiKa5i4jjCLoZl
GGnoYa3RSRWz28M31UON3iYS7lLkhXmcSTwntfSn3iSLgkeftHdJryMRqvfKyYvbwRQEJmvcVxLD
jH8sNXhvAZP8eiYkQRmln026nnOo/VO5aiRzajkoKoP2EvacWzQ4cAEmX9vTrUPKQivluC4gUHwf
9QvtwRV/0cE1gURO0fYQY2zRv2mFcNO8aVeXqkrFxWWaqyupf05FUeXO6UgeiavDjsvgS1K7gUmh
to7SCv9McPq8hVKKH8sLX92t70QtpHj11FO1jvrFBIC4sE6wdT4gLVTfbJtoE1hbR0Xpp+nHWbAt
8wxVck4CCbkCgNu1Y9i7ZRBeeIjRq+gYtIDb0+PXuG/GHPv8g+Onu9a7Q9HDTLUOW6DPG1eQfiR8
cUCBppnEAX43Rs+CXGaiMyjxuSZEjRGOqHShQSkADWgcaxr5I0IXqoYDcK6Ey81khUqztJ6jpsTA
pGyCvEzPG0YGZcUqCvTjyB7R6H2NhxKQCrsk5byV4ou8hW7olYpGXaDhzH5tYWR/izUeWRaypAXT
+JonvESkQ9MVFEHIpCcQIiw99FQeY55v3jg+TJKgHMAEM7RMwz1qfJGiaPXFqr6q8zgg3GySV65S
11icb5LCquvZIwYPmq/ZI51kbptGh+UY6yADcjCupOIs3BMK2s/UcER0Tj0ehk/CylWp6g1bPkmD
OVpZz3sGsnXaO6rOclHJ4RQBxuI7JyWrasoQlsXLctwXLqnTZhQ92OiX5HhI3sqiA4On9fIX5G9Z
aN1EF0NVWQoqa8BMYAgpOLn9pQy3or001xutQZVDaKwqznahPnorgp9x7MvRDu3FeBmQdKL13KjH
0Fg/NNK4y+MHm62e+SWjpARzA+R3cbE2HDEHqr7DXFnA/6XVUhV+s8hEKDf269rGUL/SN90DbPWA
XWVw/fYPdSN1IXDrtcafQDucrPXGfsmF0rbHByYegWs9DWKjVdFzcNqU+PgWvxlbLhLbeOqZD3SF
0mSiRLtIr5gv7k0N0xQP37jC6sHfqPKaNhh6gD2vMEwVQG785Kdl/lR6Moy4XHgmZKcYUxTrmaHi
ygSe5XoOYUPIZJF596TEjvXvf/cvGxwRn0cQGoyPrwigmggKTWrajW9OJs9raNmX8Y+ObXi7NhVq
LOfv8l51EHZAzE0RbAxI7ArJXSkVFCXs14FJzQoejMfi/FA2VZXQwDDi9r+Zi92U3p4HcDyLiiCD
4e4U/j8agPsSmFA3UBhQPUa3ZB26Nt6DoL0G4arhiP5AvWYKo6fmKVlcVmuWS2ujEljVSuq2kwZp
OGuTuGpkIj7dc6ZjU9heMc2MXXahbzhUf79e6Kj5+W+y5+0cC9aSsiSiChPVENlXTpaXNw4sH6F7
tANkawMAAPIaOrN+DsPxhfgJq9XhoWeBrFM9agT0dxNWJIoQ8SawN+VYGi7cii6FyZhvTKY8HAfQ
G86dW2D+OtPH/6FfD2KXR8by9GC6SdPYxqsj+CzpjRd8xAA9Ku/bQOncsRT4eoWcbZ+ArXz0zkMV
ta689ks41rxZY1zTONkPCvaNgRNkX/ICYgYTJAaP5Tkkv49vXMFQweYra+FO9w5adjlbwUi+z5Vm
3tTG10OzSg6NTfVZchq7afVvhec01Y5ofvdxREiy2Kqoa6QR3p+6HbSrVpjQdNhZXDE/IaWwkXE0
vUdz/1BG/ETvKyC0hQ5joKWMb+i/H6nukMxNJWR2NTFyq4CFa6hxGo+Dg6F43N0izCteREnfvAMc
TtAZgt9vj9FKGJ90wvbmVUejDWYcaXruKr9QagRL75HYoSJF77g3NOzIZ3Ap3761r3QJZNz0zMvn
pMlO7kx2YE+F/h8gezOG/TDTQhECSL2lodoFnL/WjE4Nyl2eG73xfOPnlx35JHdHJmffdcIzaDln
Ox8ZZp6Esm11q+/4kV4RQeI1WWk3VkiwA72/20vis9R/pFPqFA6fk/8aALXQtIpBzU7osPTd94BF
t2EfqGasAS+eOJo6TKwnvH3wTL5dgAqqUpVwqz5V32DEiIbLp45OXM8p0420O/hZ9rftr5zgxp1q
2nlfsaHU24nnCMpCEOK3CKzTCgufmQ6hz/YL12EwbbyhkHjm9Y6Ko70XgfZn37LFKLoVkYAn68NI
5JKwrN4Shwycir1h3m3a6eNMo2Yed8mpVa3iLyPtwPUlhuVSutMx9ix96PAF3garnrPCMDYTOv0C
AMtr67J081VllRMjGmsGo5hk0gmoYu99xgFR5zdOAle8F/hE+cSzNBs/J9Y+HDJBJYwncsIh1e3e
rOOOcMkFIOqwkThHjv0Pm+WIP/8D0yy7Qbt4LTIjPq4BYviM4i0bLXXz5tCIXA3gXrQSvbz4/jM2
7ae7rZj3G3F27kJv26t7oGyvMfpqD9xqvCYDf+NUt6lNEO3lO+NYHpBsiDgBQpcslwU2ud1Hnn1h
M/YamMu8vl4vnu+CVs2/VqF2oC6yE5+ayWLFZpqGit1yoG70dNodLQ+0yd6ORTEnpYP/vg+pf5ex
h8hzpUYfLdTqfr6YyBPILC8CI6P7y5A/9r+pS4zQz5b6Xq8SR+ur+XH+8895npIwXyVHHu3Mrp1Z
CcZK3/r9KGOFANjhHD4J3Nn054g+hBzEPAlfUHPXJeT9l+omt+2OT0D4SFLxd4WvI1FnbjzGjBDQ
QTf5JZ2eUnyUOXNmVi5fT2lqldbd1j3TrVs/ZSlzlVlXAxOOZ1YcOzKGf5jXC3T+bH0Lgn3TQwLZ
c8LLguzkUuOyAoCG5kjB2NS9QYosEZprjMjUePGm7JdCZrydDurUP9Ln1sgiC4yabUHRxvdwefuN
NWeMGKAICrG1BERG41OxXB/aVr14WxWtchwgJKPhTtbbvQF+sr6HDsMiujxVIFry0JKhFJ0tRt5S
aFJfiuMCVkQbmlFQ8T14Uqf/8hgvvw8LfvvBwlPRGXomXu7h3kdNtBVpn+uLvLjDwFymo3SfM09Q
58kss/k3n82xzs690QohS3ApFhuQfen4Cb14VdO1a2xBHyiLsmz18zXZIIqghinTaNxYqtRecIAG
Qzx214cueI7zXaO2koaq3HH4dtzWqTNU0V+oeTTjiUv1wbcUTfSaryDZbgIqpUIUMWP8WVaE1JPh
717rbe9v6Rb183umAiT0ad5+lyHuvrH1Y+hCnBzVV1twiM2w6Xz0xGffKLKyyM8Y+pH7RrFlyMET
l99cT2u7MZp1czZ/Vg3azbDAhNRDSwPZTiKfQnoKhnBy9slGdqkF25xKbsoIvnyuT3Qn7NNUeQce
2IqElSJmLIVAxhkPuScxMcthRKleQG5/1ExdB4PNkSAoE749MoF98BjywGoZuT3L+BrQk4aMcnx1
vnVjyZm5F3RmoicPIfQ/Z3531Z9rebPwQEOdjP2gAT2CSM8ju+SEIfc1BNyYtO1y332KiCtthv5B
+BXuj4cX7mMH5gORNlIgJAj/i0iG9Jt0zu+TDU7B7sdOYYjRRlIaPQtyfBqaGSBLtEE9hvxgQE4n
x3Hy/ZzGH1ubCKuL+b95N1FZdCsekPO1cqOgpdSH4uRG8PMdMyMpY+sv01sYX6GsYVteLGLdhWLs
o5D7iGcnyDr/CH5BZtZuSPAXMcCqQub6bXd4Jlp7frErDDza9z33/YdahVJ1FuPiFlsEROWi4Z7j
eGRgvFO0dPkZh+DH88BIAtYibsw07naAf9lvL91Uau4PbexMH8+xYjtw9zd6/1LTs43G+n41nWwc
J9YBSHg9soqo24L/PfpTfmQuPNztvIUngSNZ4cBmYK07j0P0YJaRgH6He6CHJlDAxWURNXWc73dC
AdGR0xYht1nYd9Eh8oha+hhxEjShIah8VOAjIzXhKkOS0Gl1a3cHceL87KTFc731RJpfxWVM3Kxg
IZHNpBtVS7kwrW6LycIkRYShV1/gW7MWm2NmNbxjrejndP4ytMzS5c3Ts9kOoPEwUnwRaGf143SY
Z/fd7tbP+OvK0+jBEmypkchjZ27taiT2sfGn0BgBah9RdKptz0ved2mItMLnXYtbBgXPUL2MBV9W
skvi+Q7aa0LeH9vjS2NoiUxW2AIKyte3BEpZPM5+8wr23ArdpkXxrqHH2bcLXGD+7nY/ZCMtJ35Z
qpLZCtoYZCwymWft4tx1y0bHJd2GAYbBwWcZ4cxjoNrUlgYR7CxzujmC+DqmbOPfTXQMCdXK1iWO
Deon1z5Ur8IWkKkPaCRrFwufZjs6xF/LKPpcCWQneyqUrb1ekCBe1TM3f67uqrfKPBsVOoz+GqWJ
GJO/bIn3ePFetV7LcpED16HbwTGeS8JJAj8BQqzmmr7oaLm4wF0JKftTLw8ArJ+HhY/uMBH9uA3M
ZikVyH503A2wJ9/E6N0S8CoH9UiQW7Pql8CrJMGxW1ES5VaCbAhTA0FWA6J+3qsMS6bI23D6HekT
HsHzKFD1kLv/IIZJZJQojkOo0WA81MeDhtezYWApS34RwOcPUeYi9dm1Yk2MjwjZdI68U6QdPfoG
7hlvL4kHv1/vckzzHVfTE7oNzhhPgT+4veOS7HwuF0oAbE62ZDQ6jEGRMppi9B2Q+dhQ5yGc9tC2
367Hmv9w8R/KoM3mKJq74W3YEkfv1uGoc5fOfSvuXvSX9I7Aa5w3b4c6L7o/VmM2SBpHUpi8Hko7
zobJ8AwiW3TidyP7cq61RqPBEjxUljapecuJ5wqRgnsqLF6GlKl9ThdhRheweMMCzheBN5ui9tu8
w0BpdQ3x3iLy/mb92PAXeGZ/Cxr/31PBD6zjQ8HKmx+d3VYuKo63EjUAgxCubEp0Mzwuamj0WPj7
trdIakiEaLiF2SFGIRsIZtc+h70/2iFCmFsXs/EpbeHNxfBp1jhEMTO3kXSz1N/l5qmFRSa4jVNJ
GEA0+jzSathgxIX7LngHInVzFysXY7D2gnxvVGOweSmVu53qZnYC84+8CAc3NqkPLP1uA61YZOrH
oESAFgjdFBwIQYnlAhFMK5XsnawKXhXz6+GkiyqgV5/4TN3hCvXLJLUdoJ+GYYFqGvjGx36akjp9
UQmqSFVXSdu4eizI0Pnxeiw6r2Y8ByQnlA7vdVtfWDeBxNkH8UGBKYEjO/mviFvOazgCnxZu0fSE
2W8/83LwZwO1OsMtbZUndfdKJx+OI8u84u3sKmer0Yuolgt8Ydy/YjEnaFxrV9S/s7FY51x4mmKr
GCRSzN+QoGF6/v/jXtEALVQ32J77+tXV3xjJxlnHfEjX3JFih70H3cCvaVhre83KtBb7fL/ZNhLh
8kPUhIevP7DTr5ioORfuaA2Jnj4Him5aZU5yrdCC6fwwBk2AM3wc5uQpvcg1r5bkppYAa4C2l8aP
2upSBhOdw57Iojx9glWbQCoDye/TzS/cYFElqDGvwboFYNrUA5nJIVbIn/qnMtgKnyi4185f9WNB
eKbP0E49vSiA1UcDHH/T9+l5EVATch6q6JEeWQV9DegSNL1DK05sTDs9k8kAHO7UExVkhFjY4lHD
ugppWM4pBPndSPA0EsVqJzAj8qWfdxrnIbCM9UWTb89wQC9KSkX2ei/IxKWHzaytE3kT2H77WFvD
4ecIgehDXRWGdZ4H/YUCS0tk22zi4FZTUhvK8WqR1cq4Ux9WUy41jw0MhRmmSMo3Fz1ML4eh53k4
nVN0vSi6qqQHxHzDZF/4T/NuZN5ehKpF7X8ODuCcuA1e0pZmFhKXGqex6MreRPWMNTZ7N+gsz98M
GLR/xsLwiAFoUrhXO3OmMbTRIkc/aTXg/CFaVLCjSaSDeMQoO1LJwBTogJ9qjYfTuV9qjhhMKNIR
JOLBI7TpgBxyPOFXy+xWi2pMJn8td9nt2FRQWU3Od0X0ahmb7875bKz5AO1n47+tRKalDViAE0aw
IIosBnRiOQfPyLLnNV4EXbFnzqCndpyQbzxu8IlUkIZP/hSLZGdHM2Hx05EAFBDlpjIhk+hubtUL
wQDDGDKOelyE8IU5QgLFTikGIgbprAWxy3oGkz27iI1nkZhHV1ld8NCIMkqslWjqx/GEFZ/kR7WT
jW1lASbTo2H4oacR1HlLCWqYuxRVjDlkRmf0DrhuyX+sgFIemy25104a2/9kuqBGoqNEY0iRFwXm
SAg1t/uS4CXl69WY9AxF4tRaVBM0mjYxDoB/KX8JJpezmU1nUJFcotSh3RpDoEbMO0W1Tw2unoiP
Ie0tgN2YzNSwTxcW77560DJt2wcFZJmtsh/iTyRM50Xg9EHNoN6NFeG1nFFmAUOb1auUidf5lIh1
8t14b389DXGhbzIY9avW9bzFkS1a/lnuyIKI9yU93S0JPUR7BubOwxXdpc7Hvz0aOdanFM6yC6r3
qfjeAI63s+Wc+doOdCsNa2YndrDNpG+hxN+VKnS2LesFPik+kXmTcbhZEWrZZu8Lixuzn+jg8pKG
iqO0NxtQUyYQjkFHtxqnBaNblmZf83ExtcRQdLODr7VlYW+2lV7jvKPszGCNE2F5f9OBuBW3+w+K
bAHr6kCeY+YBepQOVp2LxClxtaz0dekFHQJvn5o4DWStF4DoW20tl36X8YbAcTVgQIW6ACNJN0kE
cgtazTlrTYS8rLAMjqEZelSNwcsvTDd77TLovoeH5l8AqhtA64TUqTe6feXESPWN9QTTJmh80hGc
6uJ70cuGVo35nQ4PpbgyB0/QZ4v3X4EU+rmtNcpeAhfam2DY2B086VK50wr9rKOOjGPprf/m4h78
FCVMtM4cTO+yDBlMMqbdG6LUJU6WNJYcb53yZr/oZRhBvsJG3oKOP+fKBC55mEQYFb9B5cn2XAYb
mNJbFdZPFVE5wPXzZMY6Yde/yCedTnAElfEiLzZ0Prhc97uGjcqmnkYhOcgF1h1Ngh6ShlLUh/1b
ZX9S76Vqp0cK+pnR1dW1u8znIbiTiz6eZAZHb0dpjc3tLSXRhXyClcJvJoNzcIH+ai5ui7471x7U
Lqz4LsiGMMjtjpRaLj2jl7f1eWoCVW+tXzYXKFAr8/J5aBHPllKXreAhL1kyXOncq2f9WuMkuVhN
tqr3CtmvECOe+sLwGGrACWtpGroL/ASZxYfRFKSE23p2e0qinWfwkIn9MopjqeJ2jdD9J7CLreiQ
gNzifd4vyGeoZnmG5qt4T5XbGhFyDr9GyZkqjHSMen0MgMjJk4IAA5xoa9MR6dZHo/oPTUvPs66l
wwdU/q5ExARAfeubl6SfFMhp/vuj9g4VU1/SFVlEDB4zIpZ2a6NDS4JSO8pmiRY4m+5bGunPaAvt
4eSp+28ge1HcZQDb1DE7u8EVrOHPiDJ7Bne7q45po8qdRg0FdY6QkmMtm1fr07u8wZT9napCf4Ur
SuDNOFhbxConDiAtB1awz+ksR4PJMWvk6m+QOIf2QeKKV9p0aCRxR/hQi66iun9rTSzjC/utp5HL
o0wyR4lykxcGqMd1oI5n3xE6ShQNFfs9kpboZRAkHD0//awBUOrjnCLjQUQ7dDLsigGGVvUQ6diH
XlW8Kg9jXMx4QnjBvSnaMSvr/fZkZmRerZe55zFhGt1giBUbMadfff+m5sv7KD8qXFgbNJRLPVDF
KGLC4AdXIo0Rk85PiKn7+Zy7lzTuLOZcv07xihudRQlTJfHtgqs55laUxDP6CtFhh5owepuEUeZ0
y3+m/vK6ge8hED2NGdybtY1gcy/8LvFyWeiawaAk7YKLJ9em9tMHxXte5/cOBevn5N5PqTu039Kk
gCc70Tx/o7TgTbi5bLjF+w1ncWSThokS/YIeCfjZhq69GqzLnBBiF6b5EgT2Oa++uK6h2o18jhw/
WF+a6gfAB+DqV9fnjRdSQpPAdiSEg2FZzXeodqlF9fjccHeSOztQ1yBI4rpGhVOuRU+/1kFf7DIt
FXh1FxLG9T3BV/8b3W+Z3VPCYBY1f5o23/uowIc7W2IgPZem+C8Zz4qOhKvurLUeIQynuZT125z0
3W03nl3j2z+kOonOHvSvNGYeOAsbVcA3b4sZRG1G2VOE5+U1Xmr9c+VhtmOE4AlnVaGifFdaAkXH
G4Vhae+VkFnaAY0VmiYYO72NLaZ6+GvdsMhCbkmfy0bWxdJDs9qxxdvpeFQ+i7Y4LtxXX9ADdQsU
F70ELYXed7CbF5Iuj8qqFsAOoHKI4cp5aw0yNFQL50PR0VonoxM7eRrv9VWXs4Lcuqs7t88ZH4vW
qzaFsoDL+Xj0pHvRz280tvEd8k+eA27Y23MoZSmE2hUPOu/Ji0TtYoWUjkeII7Nx02VSBF4x5VLK
2Fn3QZokc4zoxvUwk9vrrHz3HXwgFjm06asSHe2Faefaw+jZNkXvnDFEpX2O9l07zQtcXOmykSzP
MAw6tGRtPCdm5GkFhE7OhcZIC5CNi1z0xfSXD9n4l+tNromq8MH7E/FaPP6WXP/SLcyBl94BZcjt
uzM+EhJ0Uh+cP58tpixwXGmhS8LzymRdzsRDo7Iz72ppVvQDfozNoWrM9noP3iK0FHZwKBpGp0HN
b3nlA/arFRw7we+srGKQ+PUh959406ytL9fLEAz7mWeSvXsBycjSRlm29gqLp3VViiZa6/PZiOkd
UQNvXOhGBI5OHpRCtrH5ZA5djyv2URZsYFN59dGnyohW1oGGEqS2GzV68+8T0SHGJwY2+XIKTZFf
N20MaOA+BNqqIm3oewgIAqShdPcYr6tzRuPQwfwMOMEfOLuZ56xP4UOwFq8OMLblvMJrhkvEXYDk
gNO6bqqVT97rNnA145ajun+th+DuiFVZ0fa/MHbU/cH3fqTXb4JCPJqpZkpgQVcBWQTpx2fbdg3W
Djh05lIBBK37eXZZHyDOw7EmyAI3/7Hawuh20MTAYeP8qmy6L/dX9KaV9aZVRlic8UPiLLwYvCJG
u99wfLwOL9PYDJOTlpU/cpfU4CCF6ymPCnqCC8nlYyCBPXzcIECGt9wiAHfNU2CbpQ7KYF10f02g
U/lL1VHaq+InlNG7uOjL4dks/FyoLqhO0ZmnEBW1X261Xb7THaPVKeRVwIHDxEUvwoB3n9q3/YMK
idO+IgoPN3sgQ40Tpsv7j3iWc+0AoA50NKOD1NEUzLequg9gnwyFss2RKMJaUacsyi+BtAjB8U12
G3S/yTskbkh6INynDLP9TCcBXRczTAi3r/LlCHNNTFpwVKenFcLx4kjrOmSD+x84H+6t/5GHPtry
nGJgpytr+41dzS0voDoCCgXnzUpCzseEJy4tg4xvajiLoqxU3KlyFAeLaPE2prhQ89NQfcAtAfZO
rW2uypn/kV83EgF963S7NRuPcg86wFvPS2YURTrnz2fvzEhjWIsRZHO8w7NjcwJDUN/N1YaQP7Ao
IWC/sIX9LcnrefuoTAnceHgS3pFmRHS+C0WTgZ9CqgUtfQVXH6qtviLtr2NbmWLSLfMmT40Gjzj8
6SqnwiskYW+TwnOBdcQLxZ4W6Qd10IiimtbN1uSIspE661BXlPQBdmeVWejGe0/o7EPw9swBEfzI
rpCiGDe52Kmw3aDDaZSMdGEZSbmmNnSIs0au17kOw7piUuvb3Cenw/eev5acDzSYmZet45GDNSTe
SPam3zhQ6KJ0hqf70ZUZyQfkbpxyRrBAOyITXb/uhw/eWY+LwstjNN0G9cX4C6eRs9wgkTTiyJtY
6JuO6VIPRR+2V1EB9pcStpUVqO9+YIBdVQsuQLlp3abPnULe080DrXuH3ET+vZEaY1NXrjhnEg35
hLT4KVhsaIVbk6iXZJr//tv2qeHEEKnn5zN4URyexPqTVh/3thmOxWol3F35QzfgO3AbqNEe5oxE
KVIpFb0IxmYOy2WjIH4bPQ9O0FnEBnBk2BCjhpoTo0u9asTw/hIHJidmVeY5r50p94K3z5W9Y277
x0kaA9onov2aExkhVWZ7EPqWPxtX0bQapGVIjKstAK9DRdSmwKiRLKB8r12jowLoYXeHOjEVIULM
G2SiYADMji4w2ePuLpnKuFfmK3JknEkT4/lafjI9OAuCrj8jL3iQdrkaWxKOJ1xZOhBN+zJwu2GK
OmikO7A9ROFwgZa1pvEnzDx0FGKGRPU3iVtxVgQr0atSv67YhuCLFGmotqtlOBr5Fwxi0Q2TY1h5
1lDGoN6YnO5SSPLjxI9kQ7bRTm0FtTBBgvUrwQUjRXZEHSukD++UcpusZo+OmcKwlIhRxZmrkZOK
nW94hcFXCJrFWzJkznn81zmgcwrF/3b/IC3nT2XkT+VA3XGCTfdQRgvRsBJ8OUttxrBwRJG+FsqE
Jjav0DaCOW5CnMI5wvbY6mHT9RaY+1z3Jve7llavj38DUVPtqyP4r8IKOUZMatzSXDwYprFzdUv4
gMP9wzMgfX3rygIMTT0JfdF49DxW2C6FrXmCgvrsog6GAVU8ufwBRfvWTiM1GJaRh7s+21z11orm
NZdCIUu9TjGFuO8Ilt5fj6FSxGdDFHqubfTpUYLe0aINLCxsKcPC9DUz42sfpFBu6OMGVhPwaVPV
Rn2RvHIXDPTcYWPH6x4B4x0eXxxDYmHHjbNiscYquxWslbhZCihPwWCLWcKhcGe2FmYVSxaHM9ez
anm3CK+k6H4RjPJEnvIBTbplsaHyS9nqQs3xPtmcgDXmS17h6L1gQS7iPXQR5lisWIEVwm8JZnhU
bX8I0R682HQS5+Tx1fvMsroYvPgwmW5a9DnSIQaZBV6kaIQobbo4+8griofFkeqCcrCmtRBx16Xo
cUXxM8GbSgy+QXRYuOCpfQ8/r9GFWpJ1rbwz4BtV34Xot61pCeFBKK02jWk5BV5MpGOdG3bstoJb
3TmpaKIq7F33AjyqFsTS1O/mEpe+1sBIOgnN21QifQgWcWnNyrmofYRwUza8PYck6w5cWiluP0lu
id/rcXBdSFdwCLfIUCXOvoJD6IzqdFyIkldrCgg3jr2zVA0lVYm+BYQKXXf8CKfeE/iVOIgPBGwZ
1JKpDWxz3X/b7q8ada5N1vE5zRiVKdQf3a8SafOD5tCJCElv7pyc9DeNx4diCbFiUqpUfeKYtmuU
iAYPUZump6XXgO6NurrwyS4Z2cWL/AzuhHaPf9MH+molWExajEUcuJFCAZXMFqDP7nxt4CGJgOR/
d0pu/URl164oSX0EMAqMit9hhr3wHDOfY5FZpvGBs4/MxNQbYSNTfljJ7ZGtFOAqfNDw4X0gfgid
xMnHkGBX2hogo35yktlfO9iwahmPd0xrzfq6S94ObQq90EvnvssPz92S6E/mVOCXa4emmPGhFHSo
CBCFn5Eo6u0jFmzfNza0w/JH7EOjaaJ2IuwuMMdf6AqgTEbN0n0vCPIFAOFp37oPbjOojgi00+ox
3JZhXkBeKSFaojNnFoCtiVV/zN8FQzNTRIdvFq2lkFY3Kq4pTVnsfsxXY/5+XyOlhkVqKy9nJqQ6
8OlTvI7yr/1g66s5MaIVCi92wGIcbLFj8DDQnTwSNWkuuwrSbmkhY+HjqR4NQQwnJfZL5KdxR2CI
h01rWoCtwTG6O90wkcWccMtfBuA39jE04kgor/fl/yf29i8OtwTMph9NqTzJB0+yPABFNfc0Hm8o
GZrg8UgHmTRJFbpSgH51sZCw4DUSgAPI/1ceptN7bFbaFPTUzgywAr0FsDwbkCrsAyWwWVPwrF9k
NQcmlOKLB4qDEYNTEqfpDsajfBeTQ/EUbXjSYlIsiYK8PsJNgLfOu5mLQtOTvjZoZzC6AUqqvRXg
IRnyoZFNcmbnDtH3vUybq3oizywc0wBCOWmZYXZ4gTBpfjEvVV8uYYZlWcJyq4xwwY49px2mHCri
kWEboRQ4roOBqSsMuupAITxMCJnijatTzsjc1vTjN3JR+u3lfyuppG1XlWw2jV0yx/fWp7LxpW93
XYQkD+H5Ncr291TRdGZ733AVQKR1RNDFb1lGuBPSVBMPcJu09kLmh7TFdszO04/lrY5Pb3beRZKp
R9/iKFIhlwaULkpwvKetGbUNvK0Rs/wD1oZXpknziorc7lmU/15bFOvfEpNPRJwOmDXBJ53HxW9j
rKiSYjrhuvjZemXq0ARndcM7USHYeWm1751MzEK6pUtNDb38TpEwmamfpXrU3HQNEp6NSSiMrT3A
8TV4md+SMNLUpHweFeF+qmGV6uWyaTGs1z3PUEUIdkW3vr6WSx1u4ecGbU0djTEZRGpYdOSda7ba
AtJ/9uXDg4gR733fZ9Dp9dKA5I0yULgOuFP52jL+0BAu0TqPv+Sx9VVWkwHOH2xvjy8SRUiVAf/c
XpjZ4u6CfeQM4qlg9Nbtq0A9LNCUPu2a1tsqTm31hUJNn4rbFPgFCBFfWyIT3VII2hhzFgJIXf0C
dkkOvAYxC04ywDdE6vrOeZEOXH9GNjpJ+sFDYtEH4JTMAv6pvzqjN30dPEBnFIPnMCns9D1cqFNs
McdOShp8kuAjrBJRArArz8LoWLFgUWnT5/kyXP54D5vzY/Har0KPwej2V8Tyvep1MftnInoxUzQN
JlP1TxlamFlubDNbbUQ6L/WAvTA38T+eplAZPypqe1ZXo2m/UPKhNYDm1Bfg3wKIY4h/yirdtiLo
97d/GzuQfzFrgpENzteBbjc9T5++kuifId8UD6JHT/OPDvmaa3Td0i2W3yKFBlQcbgFMtyk4ZG30
m8eiFfoqMZD4aE/1oz4GU8DkbscVp1wA8gvDMk72eZvXdrYgrrnMDKBBhaKKmB5xG/OyTymaiNM5
UJBu3tNI9l9gMjGcbgfTroImQuhh3eed4IyojEHXIAmW6hM9vlIV96MDmz0LBatdlgO+CyQsrzCG
iLXnR1bObmsSv7SVNbQ3c6S0pmXb7mJx9DivT7QyjwqqoJgzd5MbBG+yh3kIksL8j5PIAq94zEi6
n3B56b2S1s0MmViorVXqb/AfRVNgagMMgZKESGPkMO4PlA+2ycmMC7MysUlkmKeWAgQdYsWyqiu5
2flEwdONh4ksNwiw3mSKHmpwev0QuhTnoIWtZhB2emjg8088GBntVbAzfLjAxkipdJ38RUhlqngY
DY0dCFD0Oub95YnGHof5xi2/ThEk14ubnSZ74NVIbWb6TBAtbGvoh9OIZOe3HWD/J3UGxxpLebh0
WQ5l4UfjPTFAvwbfsNKHbeGTec5sHQVJDixt8Aoq/h9yU72aM5xUkmuVPXxTijV1uK4z6yo9Y+36
AScgHW6x4B9CATwP8TA4VNrUnfvZDKCygNwbG3ksST+occSOYoqxzywth73drWSlIcLdn2x5VqAJ
hI/1AX9Pu719oODqg4PGyY+qAAecceIpy/nacmggIrJqDwaVMi78actvu1un6ZGnc2JGl+ExKSmN
3y3Sms7WKHiOvtDrUGn5uRG8Z2D/4P8BQfCkPkg38fzEkPQgIhzAzeLIYYXohEQKlK9IqnpWLLk9
KBmSSyiYAU/nfdSNyfEuz+7BZi5kkISlNgppqoI1Jk7cQLkZvQ5OiqbnO+08GSEeAyf6lr1zgokq
1bp6iDCroaA+WsG6XNk52unTtuiL8KuxuIoNJQycPviYi2jMQVYYaNIbjtLy1yLJnUTtX8vaRcYc
tDNWhrm2lp0zgqLgrNWxkdyMrYZ5+WRUFKwnngMCN4zAE6RdnNd3UpJwQwhmBEN4WxAeLwXlYa57
FUswu7yk+c/6AwhvAHAIlxjI+i40sd5/EXNtKjwKiGrQ/y1FZzA3Wd4NkgfjobQLJYi3xZQV43N0
4o6bT+Gu8xFthH0hnMJxYgr2K2bO8QMYirY0LWU4/ciFX/iDlKGZ+6j22j83NO4qqbu8JwxDNpr9
M2VU3dwRYi/DdWGCsjaHudjQyKgmYnvj1Xw1XEe9TFSm1FYI94fTEa4bPo8PvumksgnGL0A/RBEL
mI9RNnjewgL9CdQHWXmGp0r65X3W6Ii8NQUbKVkGoFbkfkKPilQ2RIbIBnh/eLOyc30xdqjlWCN9
RljI2A7Jnh2atBaNPip9Pb0EgzsMQRbKq7Tbff0FAKFmb36wVv+pwH5Li1mTouAbag/lSd8Qo0Xa
C1nhlVMOCe4qKHVsw7KXnk31k5bVxCDQj9JQk0D48rXW6cV8nb2tWpfBV9DZlOnUKlAGWWayuU25
/2HEWUJ6QCjymbmHQwSVDkhjkDIhD8fL0EsYzHDsKIwzVwBDyKTAYoIW96ExC126Yvz2jN3xLnEr
xSUa/mLg0yCC1zG1KQ4ib6720wGcpIfcqt+o3ZIZB/BuKStcj+NSnovWpyG2+7SgFmzRJhN7eUJo
RVH8+2bjs/PFTtvzIk2YPtMDGOBt2OcEAcgxYy2uJbwwad9Lsxi6nyz3HsMnVNA6CSUSMErh9X3/
kFYRdJwCTMi+Tp8WixoLDDqtxfEsWgSV4ZwlZ7K4m4YlJjphD8SM6nxNwLrA5YGD6Jf3wZ0/K8nm
q/2pH3kKhBAQW9jQrw33deWnFfpV8hGBI8E7CQ9W5f858YaKeYBlQm6uP2l9rkstNen02aSTb+64
XBLopbt0uNeH/LrLZVxSASIlZsIWthGVKeFqezrog+/JpZTf4DOYNGxqRDKmT0x808T6TGWAulSY
aMG+bsfKXlq27HOq+QNEsgUJrZx7DjnSyT6RMqYaqi1Ch/ryM77k1KAady66FmGacUvyqhAVFpne
nsN6dR7Xhe4XJy7Y1G+/kDPszRvlc9ByoAvGNb1MlKM6q1jQxQBn4DvEDpaE6gepQ5iUPxvLizoO
iAjxXlveExczucEhzG0SplaOQn/a7WzXrLTLRc6cGwTfhBCcxpFIpxH/62GPffgooETOcnJpAKzq
v+x0ytfLNOz820XTaaQhi4D5vYeLDO6kEh4lHSgO0oAwwVya0o4KKFIgnYVwBc7QerlHh9n04ubH
zo/Dq9Jy35sh4JYpJZOi6UV//08qKcQ83AREbYDc/Z/8iQUyOkw4OBNcg3ul8Bv1nPDCs73JxDy/
tEhs8DBIKiTiErH06gJJN2Sj7h/mhGDkw1Dp3DRBNYxa8u7YtKhWSrlxCTbeJHwjDYG8PfPjiksC
nFEAkDudol2E41kz5MRq46ujWxbCXMZ9GD5nLSaVMc9wWyGTypmzKYgk0A6R2CVbo24y69xrAZJu
VRu1c7/1zS9ag6mNbqQIFGafe2nCmBfHe8gF+I+q7x8D6/xl9AMzH/MPxrxhitcRw3HyuyLgDOpS
P1OtUIdq6rtyAoFUMJjDm1zPA/R5ycFPikbYTSVwEBtK07IfrDjKaCdIqi4W42vZV7fwJai5CzOb
hsFAcfhNXW0ECOQnY7Y4DcmfkJLMtjWnUxDH/nqI1lqlxyMDf0pGlW6I0tF/YqunZkhneGq7uOX0
fIQdPYu7IGzF1kJBdpKGK1kt5ta2CCnfnZXueYOzlytXK4LvRSLB5BRMIreNv6fL5wG5yp3OnoXX
tY7g9rIqTFOqqrA9vOrFSL5/bACrjxj7ggCsGcbQMrqPQ1ndkyc9QqwN568NMJ29iFd3jyL0a68B
d1Ye/HQUOJwoNNh/u70g88GuO8TwGQPvDqkyAKmxw20MGYs3wHYhGe+BF31ULkHnatcv+tCPkRbE
aG1kcp/qELPA159NwpYCAQ2sDSdBkO4z7zq0Yqpfp6/MFNqtcCUrkaTK/aioPMQBHq+zvfRyU/n7
D2eXD7HPPJ4gFBUfzA0GTkIpGCxbWcswazg7KGmXl8AHcw8J8ulxmKgC3REB8agSXVbJyDLtaYkM
IfGXiLHDNpK0ZCXh9mPXyyKKhBmK3bEC4fT9lgorcoL57SzKmNx2mnidekkBkUBoBN/cxn6CaptV
lyA8Fr+J7/I3diCUWmwAN6G1LUZoGF2lhdqKqAgabjSCft7K90ZT0hmvaljKyiz0tAMRh5nGhFxw
kskXbUQjjQSDeTZQfzu6iUjHMh7UbuFE/ozTg6wuSC9M1lYFOoUi/0ADufkGnyH1eMH84Ht0CmWk
a/IPLx0p6UO9mS3+lJbfry9BJdVlUi3ab31beO/Mf3ydY5aMDSnjBlYeOoWP3Bqx/pfF6PlUdJje
k25lJdDlAScQIbkWN+oIfY1na6bl+3hVRzfnO1aC7hB2UEXgT8606cfrN4aRHqiduU26fkf79+wi
o5vADwkvFSuBTXtZe6FY+yyK4xi58OuN6ZfVpptxF1QFZuIdtIWlhFsze/6+Id2zzBU2IDQTmLyM
9B6zsp9u0ZUfyDBkElHEFZRdR2uOfgSORNzsY6BHEBdadEaihpNdj0H3Puc6VvS6Vig7pMXv+pBA
JahG+SzrgFehP10WgF6JZ2QLdSjFl4ihKLRay9cmr4893Dx+ElhTqJSIJ1YyKKL9IqCGEHRfD0SM
4eelqdOel8jvuYI5WSLGJILSL2sCNHaZWuStJMnexbxZNc9Y5H6AL02QAeImH6dwYT0xdIabEeMp
1fl8j06GcK6KME3uS84w1dSstIe4q66bf1WRipOLpFJ1TwNcmyMBo9sgy0poVSLnQwSymti9078Z
cQSj52zDdN6ZzHU4WrnMtgYIr6hiYBXlQRU6SJRfmMFwRvGHhS1aN08aUqLKGM3gVlvaCH3uZOXd
UBUm/UHd/DUxT2zH9Vhm7dass3jmOx3ZN7WcDZMAEuW5Z+ohMwpdrYMYZEUGP6Kqtrkvr8Y+VjsB
8UkYPDYMmffY8PCAmHCAKAcQUIZ0lk9mZL3u9RFcY+U8qzod+8sfkLbsaQvNS3YKjgeh59AQ5Vk/
VGf4c/NCiEfELVhVV1TgSzTga6/PPNMOyC2xwVO6ePFZdIqWOJGOgKHlQR3ilE4cpH8lKOBi4XNi
5ECUK/Tov4NXKvKCobsrveyddtbQVyqSFOg9sGV9Mclo10IAy3ptPzgiTzebcX/Hg+jATQsxddqr
SbLGye3cGg3WwSL9RKYQL0lZZZ29WvPELmKcBLU6QDAoIZxp6G7dTt+ti+dr3faK5sV+upSMAQZc
eglZTZrlTG3eEhpU74MYYdo5fC6/VWk53o71ze321t/oxdWJUDF2hQ6Os6wduXjO7niJz3yHioOm
1ScbYx1iJ3ngUOKhB+hiET76NFy0isxWO3fi1/sViIUge8iqsaB2ksgwou0rKOgQu6Hw2KLQeOVN
37+VDtjcoWgOqsL7ME5Ny8G1HH8kTLqfOT2i1vxB0F0qNbJdIXazJSSjUebv6AudOynLVw+CENMJ
aTwkVOFEpx4QDV4FZh7fww6iW/kUG29cnEDgrMqgqPR6tcOKg9I3nsG4lGoVJ4J+LNK+TQfM2zTN
oLtwYS3o5c03iQumJrEY2cwWrAbw8RSUaILgMQiawoidprLnTH2JhG29Ely8+7QpBr3NioKyRMKY
5ziVTn4mPjoQGgFBqJIDmcl8AMz1gXCfECgkjDGmmpikV/EK5M33Y+qA6IJbNlzqeaJdC/sGIpoK
wZfDDM4zp4MK0KAvBD9bWOq0aMk1XvLqNDGM6+NxP60bLrbLy4GoqioUygL3fVIod6QJ9wavG53s
Ajbr4cOM0qLSR2n32rf3IVqv6re8Oaovh/Sr0kwK8rt0r5j1L5+mx54OWs6YOl35YoD7lyXj7Lft
gq2Jg6QYPJ+DgN4onzNoobCY4Xx2hJiVm9zfhyJIulffYyfSjboOK+T058I/8g/7rcmvXxIDW/su
1MKf6KgztsrPK3qJFLFSzVehj3/7i9Astvjs0g3btb6CvmE8/tIdO7kUaNOLMeTnwR5v5LxyIR7f
NwVmENYY1ImByedHdgW9m8mg+NTNjRysuicUP11IhfTvlhhAq6g+jyXtYXfiw3ssVR6na+O5r2iD
/1Wk4b/gedKpmLhZkino94qbLGTyS2hAHvImbbfqTdDUPGruc2dqj2OwprIpcygvGu/CQFNRIwnR
622F21a4gqcdJVF8U50WmL/4GFyrPPVFHfJ4r8WB7iuhRxD7yzrO7ouwYt3/0dtMuVmE2ihrdSMr
N6TLn2sF/5WZhM1Ev9IVoeme0BvJ5anRkhuzwnOy1lhN76qY1OtL2ND0T9HmDUqriB9TmAYZhDOE
rq2KNBuvgO5ylXyHKc6Pf0ScghB0DHbAAs5v8yDBx732xyzKDVh7sJ4lBG+q4vkhshB3+16HLoxs
WpcMJjlS0vBI+l5xrpwvtecmW1pA/0I3RZDgDJAmDg8DFIPDbIvw1p/+784z6AbLTU8drIlNJeQu
uCEvU+2Z2C8qC5rVOsjXpoq+EaOXaq8lJ1QXWBKroRVwK1m+/EEIJ5RI+aZ/pGLwOxW6E3+vwd9K
FGtWKiDwPfkj25w9rPBHoyPazrugcuu/Air59Vu2ekQVQTGgcYJH73dOB7DOXs8zy5RD5nZfZAi+
mhCpedk9lxdUQaPjl2E4yhZZRLb3C0rtf9rtLQOgyghhte9wVO7RvsEa6vc9wOrm60mgRzNLROck
hAyYfNkNs7GraanDK+piqrj1j8/YRNSNMX2sHaDh0QRzOTUdID15oG4qR6u643esux6dV/NIhJ/d
vviep87cCwQPu6+ZYAnLmLFasWvewt5TAIT8TSfi5Hr1kurN/Puhcj1b+6JEml1M4BcbS00wqBWg
KGgyBHakO7FtBFfj14TpZ5KzAtapHT5MmSVbyzT1U3n8Vm4waAE4Cp/uA9Seij0LzKhm7KlEEbDH
gAb2L+QUMNa/qpHFfvv0YGagVnfvw8OWwnCRs5hE8yp35gGPuHXlAUBQBAH/FjXAJu/DoNE4U5T5
VZ8eYRubBfAAA0FVC3S4zplj+eST2JVHitc+g1WkrqICB1c6OxX17wFav91uD18O2Nh3P+MRTwz+
jK9ze/pqkK+H8yBxQXpc6R0ZfJeItXl6NQQ2w6p7PEbX3SBID88OCsqngcquLJBxsb/tmwP06gls
TJ6lZNsp85KyBJrW43LZEMqNvsSavDuhGRuf1LlKr0d+5EaTHFUkN+vYFzcKKhZJAVwBt/9pL271
ZFQnXFEqa5mKAWKpF1TSRGf/DKyFYeW0jjJxY59YR5NJys2VkgpDPNCbK73MrRaPLTj5J9ReZJVw
mdAzQ3zskiHCsxR76IO048Sh8BWPNT6e4C0wnFgS/BbqlRgTzHk+PvMNgQF7zm/oMZEO/c/kB2Ey
m9ksRlEH8oiGPo9rKCMu3hOwdfVWkI4dX55WqOnOVAXJjysv8PtFSDkow0a+VSm1SUhw1vFvdC5E
0ZZPIjf6lIgwM3FiGWI1EJ0VUEAvCx1/5KRrgoAIZWO/uimYL8I2gwIq2LLEplnnwQIERudYo3sN
P0Lk0s+QIbKzivC1JhuiH6JQc8JHlN8gCZmJ61o96uuHZY1767UXDbPu4JLp92wdn3wGs6odgDzj
KTa7FCWzbcf1ncO91IJs1f29ENXiW2A76I3G7vPPjnoPWQ3ATPQNQZJYiij2WqoBzMeKSjoFwdz5
v/82wx0LC0DYUgZnTyrhEbtvn+fC5m9vh+mNshAatF76K6tff0dKalE/F9saDmo0uyWw1sqVLRwt
rpiekPrMaxkklXq2suHunFqAoSWACljJ3xYFI9x05Ica6J//M/MxQIzpvCa9oOTWJZblKUuX3Li4
gC7kVwxUNLxnN5ygfmUnEro95yKP0Xds/9AirYzqyesLR2+1f4NWD0t6kdwnpC9C+xytWluvIsUe
N+iECrfTTV52cW/KAcH/cqWO+9+9Gh6acJxovJc0wtmEYCQ0Lrn+Jm8i78hWiulV5hSQjuzWwwsG
jUaR+1PLB0YXnUTKdz9EWppXwS4M7COpL05Hq7zjlKviWbxerlSijYobwtDoDKNaqE6AX7iqwYeH
P0dloM0ZQKpFZePZNrqOMG3PgRff9unywzagd+9FbDU5IT0u8wsUcf9+C65dAquiaVbh/QTHmRiU
Dgulg9ScP8qZPvxrTZs52Y+zXL3lj80dVtoRiIGFCzO7QNvqK+ehI1IcfnlXBvizMKQeV6O/RJHW
1uA0EZLKHxXFAYSbSZtwpGWmhF1RLk7ypbsqRJooYEuzpTajw9g6sRnCRgBqICpq++0MH7ckfNjL
uJxHvnw/2+CGKUAwKAcIv6Yb7P1N81x6eG5tvTWJGOEKc3ovLt96mZqA3I6Vp82R8iQTdltefpcg
/E/mm7ztONxEPH00K/Li2VkX3LWMtEuceggmelSW6yhNqmSpcA5kNgJ5giHY2dbr+B7t4yPF45LA
p8iIjINimpsso44rQXXp4CtBfTiqaGMwd7H8KuP8TVF+00+KEl45TgWUilrF24BZig4gX0FU6o69
eCKCWieSPffZMB4oILD5xDXUqBy8LMO4PsRBtlE77qX4s7lvwfM5MthrLh+ZtOOXubJrVkDS8VtX
ifZvuJkd+GTkGNgvxIr7yjjYUucldQ/EarIi5VSGBXT1Sl3pj7nwhbOqrDpqPfIUMMIyBQNsQuAj
FHfeHH4maCv0ocUITxMQtuactCNgrRc1ocf5FMfygpl7s8CGL7uDux73ZK+QuAHLdp9tkwX5QK0B
SBZMnuiNMXObDMmP14zb66H6kK7i8Oh9BOd3mnDjx0uBOVoW8W2dqg0xyqPyBoy64t0PM11odxCv
8VvS6fXSq0z6sIT8SCnhC4mpExwEsKS2qG4lP3B+Cykk5lZgdxbGTSun0hJ9M5pO1S3VfNJdNN42
Qd31NrakuZxN1QIfpeEvmxDhdCN4e9blDNRCkX2kGm00B/NUMpIcStEMF1qnp3GtrByjeA9xo4UM
1CwLGuuv1cAWAnElUNOiHbCD6FlVdhQ//+Z4TQwJZUIlUlqszq7KFj7SneBKh27bjst/qiI/9ROI
tGpH2Mqkla7P2d2U2ZIMjTnvYFyx9QiDQb59zazmaDxtYu5pSLHIAoLcwkOB7G7vTbMTjdtoyK8n
7mgIn/QJ1HSIOZLEoGcQ3dh+znqTlxlYR13CtfjjzNs6qu+fcY3cN44BHdEn8ohmbLftc9vC7kpw
3Pvv08bL2dR0M/p8wU2KdSbdCa4BwTXHXWrTGBQJpiGsqCX8qhDQFU7UfImqj4gv92jMBKq6wjuU
uzV/Cld0dhjZLxuVjwkfZDQFvxuycNxctTAVMZHvyxDb3Xk7jRZb91cX9uK3xnuIGyfCVzvQQ9G/
nLtZ/uAdXFDIhi54qt1N8DhhFWNK7xRyj4JYZ2nhWUilfQrEzce9AqBnwlX75WaYqnqp2rqPs548
/E98cBvHCbKEofDIMv69oMjeGGCwePFAj4YGPtVE7St1NJmeSMAdb+l0zLHU/am8VkRWAHujsAXC
Xcf5a1Zf4mXAKB//oypr0fuegTcYVW44TGLPoPJhjeaPLByiWBm0eurguOW16BH5Of2cfD5k3Vl6
aAoIQlIz4Bw+M1hz/SFsHrdWtC+43/VTAmBOWI6P7WUgnJbwdcdl6b5MFY9Zj4nsS8bNIOkoO8aM
281eOC4bmEMP3pTAdQQSlBAsQTrVQXkY1iyxEFU/cFXcL9mx6Zyv/maLHagZM5vSdprOELT+7zLs
G2hd50D0cfvw5uLj9vJ+00hE/Hz7396K8RKM4ava2gxvWV71E9yNRI+JP2WEjASHWz9LW0gXcJVK
M2KyOCceIeub+uWa4tHXH+5OSX/krn4WOMEabyT1zwpxpqnRuX7FAEexPMommv5YmD/SvIcpmdLT
bwHFYMz9HoqgQgBVfIo0t0PGxRcDxIlC09JM0YOnQhoq40VNilR9Sx5kpNlIlAkSSj4e5v+PZUZU
kkvEgqmcUEUW2D0dgL4N4EwePeUlkaTzLj5jpWO5I9x/c+PdEpBeNS8t6hMRSDkuiSLVxx05mKYQ
j2Yiyd5kgs9vTHz9AsqNR51XxScQUaqhvCQjFEQLkMAnRrUDHZAbkZZUqGFVckooOyAamj8nODPD
FyXB4WUQwA1b0EeleIOKRN/yVTP9nrd5Qe5Ai5LV1G0mUA+29kMuM2MWeix19uzus7jatws1MDYH
YeJIOpcxdrgWAK30l8BUAceO6HQ6S2ULV7R7Q6mcqXh/ogB1Tw/Sin/2VQQ1lbnmH+ffXsuLLH0k
ZKGiu1Us/qHmUs87FCCm6dgOtwfzBtolctoF01jOH9kO3kZC3/XGg1IrALeU0U0rz4xQ4TcmYq33
1S6U3f+cym3d1Mmw8D1Xs4wd0spax3ILWFnABvFQyEXonBLQMZt9/fbfdiBUbZy3RkogXRUbEg3+
TcO2F/7H2xuYJ6buP/G7yVjR/7QW8fNioczEyWULA4giDPw8YaWAYyOX/HfMCgM5p2PDxfKnD5nN
omZ4q9y1aTO4XZDwv7s1tSJlgCSVxeWSLJEkDqHPeioLNS5YEA128mEl1LSu3HDDXpClSxygOA6A
wzVEWno9UY6G2Q6ey2b9wlMX2Ssd8LZ1ItttBqZAT353oOfkJxxfySy46fZR7LtZMzmbxN/2RvC3
7QHnwKqgLba4C0iMEQ+tSpB11BsJfM+yv1UDcl3MBrdYtVlGpoWRmjzpLcmO23Tn7gryTHOLJGCo
NCo60+gwzCt/PdkcvjrHaRUL9l7EpdPxPqW9HzOTQmy3HvzXk/h2+ex6LpFdUD+9YmX2lQVoZKD/
aFaqwMKPq0Ym5NKCv5lHzjcxAgO/jt41/3nniTYol4VtFhjnX1DoNIb5KBmMb52AvZ0XrbsmdeJp
HK2E7tATGwH0JDJYVMq0fiRU0yy/JKnbHa8iWwOIaxgH3kbKD71mvRt53O+Ru5/Q1yno0iPdrZ4Z
K6kCmHPp1E+TsXFJqwEMBoh2pLan+PuGgBwQ9irXjZhLeBl+b6j2Vz0MiswydPWIYTieB54Zku8A
SQ0/BblbA7k7KOa+4TaMy33xDPzf1z6AlOlFqYkrOoeO/CdZ4dlZOSZeKoGrhf2yUgVdz/Whf0C5
dS9WIy05EJ97+APOGgxgco06nK/1JmI6weLOupRLM4TLENyxfWIj0FjsklSR4RK7KhccRfs6mLDL
PwbLhslKivSAgV3fbxg1zhRzJvqUHq+niN14+B1lbLyJSWJPP6abg/tmLRU9skfeiV682GczVS9q
mxlAjlq89NbZKlSw8kKDlWG9z9FzXCpZz1aQkHrjb93PewliApibxm5zdPRTE2vq6y4n2IVhwcHC
PPfnCdOdc7RdiOehrLVgd/QHd+g0YagVLjKYvHhskeydfGXwaj47b6EVN7vcgzAvy5gQKMgHwV6J
JbGQ/wRPPp3voTjtH5JYCB2xRFOO5OM5zkTSU2pI0J4gbWblKQgEJRIyCQHqB7ESKTvnvrNqOmOk
dGbtWkbDRpG9IRmDtdMEEyHDr5+OakczMt9dMXs8zGv9EdPk/Tjb4PX7b7GyQe2C1pkPes3dPftZ
uwjMwSe4rs6Y9eEUi4OdM2P/qoGTBCgvbLN3UoZF0Z3xLIdsxzqHvM464ibz8io0i87y/ygw9JvS
KtUOuK4trSuSuB8Lk+jaTmJsJ0JXqFpLG+if/vAiBuX4Uxku3PxPbUdvnRMjpyT0W2mCq4OPbfgC
q39OSs9wIjpvzpM3PSE+KRM0xA5hguLcLGk1EJ8QxefyoHAo/NodU3Bq3aZxor7rPwDYhAiHBYb0
8yZeOIpzmbUgWWSmsObA07JOCGza2CyC+e5ReMU7rdkMRjqWaJtnwC9Z9slFGjn1ow7upXJUzMWs
of0eVYa4ju/3fSwGjWFEaU1tor3cvmHEDhZDmzwitYmQgeQHJgUHr7Bou5g0IV/2cYDdXhI2swfU
4bpuLfWXYxcdSpGuTCUBrFL0Fk7h6wjgkjM5iLAX3E3jd46mXHxcber2QBbyZWqdWk/feXia2sg4
4Ajk1gTGthfP89P9j9wTbRpT3bdGyRer79ZRDJhguqO2TovwsXl4X8HJs9T/Z/a1HPftRombnnZY
plObhzZP/M2uZmdKDBvHhtTQYtAV+xDN94xiMfZnIpOyMXtFhOI5CvJ0JKkQx6l6Tq2dAfPUbqmu
M4ZQWRuhTHsi+xizsU0AHwxcRfSXMHqa7YkeeA7nEtXM4YdtQfsmBXonIKiVC31feKL092lzipTH
wX35i27kiLLgh+C5GHB0k39APhgBiCG1HWmXxjIwTjQdUIOi019H/47pSuVU4x5nDS/Lx4njmFG7
tzktL/RPwa0/PvvmjKjtd/ypa6NXZ/BpHEnejhg7nX9lHiwnXlbKoSOiho3uL6k6Yok4wOYG3zJS
kXGRLHTvCyB1q7ufAcfv28dMkUciYaDRu5rKt5VlM7hNUbVoLl5HGKxoY0aFC/sMPEioEN4+Fd1u
33tbg/6+jM5EfDxwz5e2+5MvFOS/UaL0+eJM53Mo2CegmgD2Ez5pw/0C444o/2+J9VF2PtWhVvvm
xV2A53uNSbMPB4KpC5oyJU9TiOEu679BTEkTC9rflL7klXTwfbPILhdw/92ZKRH2r0dgIowK39za
SK7mRiTHMcDFhlzpTPgjNAmoU3IvyjRLTER1KFBgtce3kDzU9zEqZFruF1ozWUShHSVZlmZj97He
IHn6qwKQAT8rHHKFiGuMBQ5G73B/VsbVFzMCLpqqlgI2R0tt5HnfhFqb4gudGHditShQm8ymXRpb
UFjFwxsfFYY6M2/r4Tpzm8pLbQFsSkNEgEhurZDG32ngVir+KeESv4v9RQFH8DkCfRuEBV+ZUD59
9K4sxB0ArzHjWhu6pJbPx8VwkX5NPP1NSzxBFw5aOP8ygxhIxrQxlVcFGKjemlxNO0h3n2mVbFPo
TLLXF38+BF+QWn+iEb+Xso6Ke4HsDVC6vEbkaPNeNOfRDbcZZo6/hi0amJ/xYKDgmU6hLiIKmQvo
nj1+YSdbVxLjiEEUg+RyCKWjRP7HUsIq+0YEJNCKww+xRb9SHkqvmvuHZ4SnG5Bwd9ZDA/K3tEal
+ag88h+yJABXWRQml4G7DarGcNJuYzdx1pev5/nti/uukO0t8cFhGGRQiYl1DHk8bW8CEpkHZn+s
TA6EjAn8yYBHp9JQt3HgpPheOhwFiukllHD3oSupQZ+Dje+YmM78jvQaXrqpgxY/VIRzUtjr9Iga
cqCX8i7catTpQ54pcobvEyI5ZYJmdFw636CNfQxwBAd3LwQOvNIG2sNkigJf5/zPKeVUH6VRsez5
Rq1cil/u882nBMGDPUoZS4vpqGLDfFX9qftvdJE1PF+Gk9z99+XDucjRwj0YYOluVdUuYLg3xgpe
n4W3Z9eVCG0dYnGvdOnFfnj5jfvG9H9V7ObbFERbMPsEIkfPn/0o0z+Bp2AjuxyJfGvVcHLNYmoC
27wNbr42IZWYCRmyJ2RH9ga5+lyOzSOLZxj0bIw8h4sI1QyQE5l8YWekHZsR5//kaHnXldVbIhI3
z6MAwh+gK6DMOhco9CidIGam3csiL9k1lzu9upiEH5iibumqjWF2ZCZZbD/tpwFM6he9jBb4eAxu
9iNF2dH9nZoWt6pXqJx+8C6lt1TB68iXDNsN7dIVjS7K2DmPtn24H6EXTogYNmFRRBmo+75Q4W9S
lapXKTlFbo1FHY5xAvL/FHshDlBkD/bgfP5aaZb7N2ywz3so50rI3DwQWzbpklNM7FtKLBHv4B29
J3u65BPIvNS/5J9m3WCZuopHOJ7p2YJYSaT7UjxskXF7hbv8KZ8uVnNFAWPKuCmyVRua2I/hleND
n4AXpS2VCvN7QGuzSNxLLEbAakfgEjPWDHVGifnHk9E3UIfpuaIbYnZ1r8U8xl5LJCdUKeJPyCrM
6S0uPv4lVUalVCrPJiMrBVLhiT29+OMD/SLPK/2ZyV9kwO3yaQgr7Z4vg0sMWzK+ZfWvxzsKVxbF
AiJzrBy2xHYSauE0d+l7fJxX5AgsSpXJ7GUUklaJv+YrYxczeGWOyjmItN9PfLzS8jMXg9BrJcP9
g16HTDidx80MEO7fn+u3B10goZfj04FTdL6AXJHajP5BtmJQwLizknd6hTMVn4RBUGs1RDCShB9H
zxJa2qrczq5Y2dglqSC59xqv69Hn14xsIusuz8kwa2L3jNJaprRBggnbB7S3kQ8ZbrFU9OJsPwcK
XmxLYoI0MvuXP2tKLtV3mz3CNWbcSzvefobuWIlj1cEx4CbJcCSxRPTWXOc7u07gIghyi9cwQQWs
AP4YoSqR9gO4ewap2Jb2c0VhVLv8lP2x9mnT1sVvQKrKr8D7gqFWMX6ujvHrj9AtjPCtawYRtDRf
6CkQyKfmh5q/fzU/SSgAgI7W5uuDdn3WiGuMC/I0f89RNy75+0In/dFao1IEnXxIws993vBpMZjx
qcFf44by2RZ3fKX9Srcmn/rLeT/cow2WyT1V+fwB2Qo5hAS1OIOsO4FZpzu3HYCW5D5lXZPJT5vg
cU9nXCW1OHBpkmihuI3Ph+IUpEGi9Quq5i74cArUM786k7zj9pTsIsAN3UhQRKMlGx8VRpMNsckI
rhm4wpt5UN0feW6L63aNHaFcCEQ7MLrpsncImZ9Sp3VNWvpCFCUDO53VHpqi0hh5Fsf0fplzq87W
NDAP8vL9UNR3KW/f8oOl+DmPkFmj7TIaXe8PvCL04LrPNEvRjkKVCYDX+k3aV0r4hJ2qH3VlRvxN
Pa6nVd6fFkaC6D9NeG/kVj0aSzqzga29K0v8/nZMy3Au8xfX8X+deMW/iNzxjmCudgLDYIV3L2Ll
HU03RCXt/7pU8qSnaMb74/BGWgfsaP9hGKKi1sg1/YgBh95VU0cWXPaQJ7cyv+BsjUXdj5j/j5dI
qErFlFvD3iAHNMHUkwHkPpcv/HfU/rSKw8OUeSGpSMvv9x2LsPg9+zaesDyxmzbP5FDYmlnRBBYb
1yhG0SPuW0M/8r4V8ytE9qoDmXJkwu09sR3mc7Seb9zGHeDwsgmMsxWGICp1sxtgdNJ5Jxdo3vrt
qeyT756zV8ITPMq/Cbse677oixkfZaElhpduZcB/5YkbIiEl/PcS9s/FRarQp6s+oPcGz9vlwta/
QycyPNjavwYF5pvAFUfx5eltkf/XbaADlls8qJ8TVtR0XkT1eEj/R0/IOYIxixhuGfc0KfpBr1RE
PxPHsYWc/GHXy7iY0jx8LO8Gc03zfZMpor67BHDikyKZaeD3zBuryAKrNysMOJWoJ345PjJOpSdj
qDUo/PZ30/sLoa/cFXXpYjm0CauFbuVFQ0rr739wGqonSZuQGEGjR47CMplEsItp4RSNV2XZ+4dM
sm5l0hHiaPW2AjD6DAfXSsiIBMMsxm8S9XNuIs4U8VoQmQq5FfbZHX4RT7VAqK3/vAao45XdzV5y
K2MrooVPceDo18gH97CzY/ieuZmc8wi9X8m7SmwlgCGaMDvA7V/rywySvND3MviEFxYnxhutsvhN
sSD0trMeyiMHrxq1747oWbx2Ickx/u47tfqiKytpwW+8zd6FLKven3hZoGnmUpJ3xrsbUSkJFnFR
hkmq6uwnNxhLoycVw++GTvl9RBqVHr/obWNGi/SGJ395UybHSO+rnn5+EHpsZl6vGWBNj5RkShjX
jiSQ+xtM2hEfIc908jLyl9Ca4WdmSGj8S5j1+BYN9Tb+V0VyAVS6/GBRCFbhE+pxfoBHwtDei164
7HOI33DqOs3jW9Meyi75hAWVLpIfCzyIqQ5cqA87qRvYm1129HP/mihu5/bNdacZHSFBr/3Q9iJv
7hcfVodEDyofRmyddryfR7AfFwnZ4U2GprwOLWyjyQhYwyxWUMcEEBbgG/x9jPsoNfikBl9V48KP
ZIRvc2IThxTs/JZ0UZRpVYibn/iJQ1rqapcKBK2JKpMz7FGaYbWTgwcaXp06TZs2VTzlyB1BW8Iq
gXFnYlKzqWSziH0OI/kLdPFt39Ef2UDJ+0wJ2ndhNuByEphBx9Ewlsqnaj3x6iPfmezx1oGsa7Tn
xQMUKL6mzWY8wf2w82R3mkwm6wXjxV59o9HxBHbO9RwCpz1XICtHLUvZ0006+hEgEMV9/g2U+m7K
9Wlj1mCyX83JzjrI7ZtILe5J668xiMxalQ+1Dyrz8HB2v72n8abJ7YClhfKakTpMyd6vm9JhSuZ9
6xH4IJXmlTmlydTDIhWdg64VuHHCtb6dI21Sb6e/clUMad/RK4wghwdO5PfFGzEiMDuIwWm3Kf3U
eCYmyminEklszIcCJF0fFDmA3iGc6eSk0lDpd39Cy07yHOh7BtIBaHto/A0bjzMk++eCX2GB/wBh
sKFYdryMvuMzCSlBlRNwkWW73vuF0Crx9ZfNEgQEN2vLEeDG5kfMNqUFq6lvJCAv+TipAxAI8VF7
ygocBA8RQKVjNW22++AFkhXUIdGMKpvk7+NWG5E2kYNOzOrtzBm7HfOs87+n0VqJjziGq6SYLy/5
ZB5sehQbB48T6G0M3Pvd99Pm0/X3OMiuApU48am0s7xDrooVcPTEs3D84upwBYczU+5F5JAO1xCd
gJt/bruHk+PuLiy7+lvozf5/2QEzYT8C+6XkcrSsQSG9xLsSqtb8iCcFdFWd0slQ6JoNV2bXsfFv
EcGeoZEsyualoHqDuQxq7tGjgPjwhxf4ZR02CrzosOuvovVTvvlrxF8AvPw3G/rXdNoVv/I2FGMf
i17PtIT/XONCTimK0qcGUZhbrT7OfTSO9fmmDtVKYgDKyjkDznnrJacxQhtWbnLRTecMDoGRqnQc
6BZJEpt84EcWYBaeDPzdjldKmjR8UD8CFVRopo+QezG7Xst9SpHDirYFx51jKT9GIu7v8uLkgvG9
OK5ZsBJq372zsxDLT2N5YRakZsA9nkDt0MplB1evdFYcB7ipRgPLDFLlEc/Xto2TBljbfWa1oJqj
yuuMBhtZh3194F66bUNFSuZ1dWWC4xQ3638wXynxnqASk/XrGzPwowRVvioPCxYS7nr/+0Zge+5V
Q9wgkLOWDL6rQRWvg9+Kez2d4njho0KYXgGPQAa/1o3ztlZwjXvWx2OQTidObJvpcKC0vDWr0HgM
B7kLiw55StPvov3rVtLibGJ5M50uTzFncQ13j2lHo1p/XbSl528hMbUu0KWVXT/WpkrXeJFpBr5s
6+jrUlORuB0sxEXhCOcB1h4Xy+G3MxRKr05hrccATGZeYDlQYiZYghsxWWxRPG2D2dyVmVuC6wkJ
7KxZxkNNk7x/HjaDfyCyQRNbT+YA0Kks6zoGb192iHGaRMUCSyNoL2EzZEJgkRbmAG7tc+VaAV8n
pu1s++X3eZvMI5sb8CBRQ49+VuuAazkzC3JEGdKPULOstAeSXzX/Di4g0UORaG6XUiK2gCTblEpj
ctjgTI1VBFA24hdFdoCz+LvZVj9QWnzL1VWLv0DhVBa79MJaswrFSRXV4Z8Xc14n7PPB5mQzFkRQ
0/48p75J29SzNqs+PQfwZkn6I1bMfKJfAGI4fixo4ht2HChF2bzgH7D699NojwUHmUtTP29+2ZBu
GS5/zXqywIKczRazaA9fWN6B1iMsBVCQpcJ7ajcmfH3lSww1AY3LU/5u+DvfWff3PHm/hbGQQIJs
jbpBsIxrTd7Rb3CnH4+uF/ll/z4zagnx/CS2w4FbHedSDwJjEXAkfefJGcvWKxGW9JkokRneeHYV
Cj6MIPnBXvLmWfIo+Eynfloi1aBgK9vOs8Tsi8YRcQfXuYZslFEU27ZqUcy1OT/70rAToaeoeIc0
pqMTZgBJ2H3ckvvUHrUk4HNd+gJHeALZjQgdikDJRuCpQfh4+tMPEK1zI5UfnIalbfVleh083x7U
cltSNhDdnKLFVXlQh3MVplbSE0Xz/ivg23QfUDm1sjB333u7IM8W86muMI0PAoZ67ql8fotT4k2L
PRW1t2gYXBmJZ3V1M1WevijSHzXQmawGnbuEnI0uXOirVmgfMIXmATJGEPB33K4u9f6QCOQCM7LA
26CnGwMhAJ7uYvMfu0Jw9w6WpcbZcPHLZSP/iS0hm4D/Q/mnpG1dPa8rX4Egzggqj2ODjfLXZuB8
aUwZ0/WiVpByWgsQwRGeneoYu6cIYsDlpW3vzHUcj4ejoJU5machf/ctubTyqTBikBFF4j0wByjc
iqupbq7zcbL0+MEOjDTe42igxHMRICdtE4Shdjk10SdpWvpSK/rB7wxjdQJOq9F54DfKIicC3uRx
qJE3nzi/g5FJlcsgMoU4SagLV5WnqKPNANYVmRHnXPFOOVYJIoASQB7jUhRnnMi1w7rhT6hbSntD
wxcaV9q7U6IORqqs3WzZS0Vfxq5lCpFrYScXalS8830wQCLhJHT57tm3j7+MI2l658073Xlhatiw
XFO0jSWuEv8qeflEWPrJASfZ4iJvLBHjYuCqhZFQ/sx3uImJwTHEk85jOin/JRL0NXCMbX+qjaja
8rAxreSBVZldFILQzdGYPPaNxhhy64THS5jt10LhGI12UZLp+ErQ0yrPtI50kEhF/Ze0Ss1dGOET
RfZkJSKR34QMtwOp7dwW5Yng5pt34c6QNvu4X5nYShw5+eKdidCtk+KcNZesogEKoscyuZEBY7lm
HMw7Fy//PTKiAopWTSHhtmhyiYOWEPv8Bh1QPbnOPoUqFjWNhOaYXgMeFlZ6+8tgYxBl7u/kwvlu
R12X6VcjI2qMshvBUihCFelt9KjvbIoeif7ZFFj4/e0uNbBP6L5aAGN7iv5SpVNdiEgTTFQDxQyK
TzB0V/btqgkef6D4SdGHnrlxZHrXzbcZ49WOZTRu5CP8IN/S8lRzyKfl3JsDiD1OadLVxMgmehwH
6fNJl2wGnRzHL2Dr7fRrCI2KDHLumFaX
`protect end_protected
