-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ollq1+Lde/Eg4sBiAclYC0ZeDSGvbTIx7pcebgBuFLcBgQr0c9EuNhobBJFWQ61fXZPRZJAuBgfv
ZFdXXxIi1pfdFo53+xdWPT/ZlLBS6a/GTibRG1LkGo6ah3yxOTivY4Z/dmJIbHQyeVfubEMALsgy
/+N5T2furQG3sZ3uHHbdSE5Lt9k3mjTMaLzrdEgJrTnsJEtPGrVrCq12U9/NqH/WWmHn5nfGjCL0
sNnxm9S2t0+a4TTjbKNZHcL6Hb6jm2LREucA/dPVZCEB5Hd5Ue8luhHXgn/5fCO3A0hlXWB9CDyy
7jecPMsnCU2qT6kyjDz5Gqw9PsuKLSyM6bk5vQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
YfUDqgyno7mDMqq3sURk8mjFiSLHG476RqxYoQY9iZmFSYU+mYu0QLEdSpZuGXlneERVyNBxygov
sVMu5UVWaMGWVoRMC+N8qVnP1ONwrw3QWTAoTOCE6L/wEwJddxyCm9N2j8UqMrZ2f8nCE8GZKsbv
Zyh5MXDVav2hQmYENFeUU4ZWjO0hbWhHvC9/Wgz4p4snZWW/xp8fYk7H7rTtsmMjAiPXzH3uM3tM
boUr9NkwdoI773qSejKb0iAYe+rdc+jhHvnQ8DDgM5s4C+jyykCSd7eZdi2DSLnkBV5fN2RQ6bqa
qAnPE99vxpthljyjiNcM5a5831h3GPeFic+VMTMKxkztd8nMjg90A7S3rBk6A9Uz2MByv6+EoBLo
0Y/5DD33EJ8Zoc7zZghrqoR1fjfhZOi11LPwdGC1ypXYP2moDGrK2Pv/X5iRgOj2OLnZz0rDSvsf
YwNu2AHPDaYlyIzh+uCtDNU6Aeq1vKQpY1U0or8p+mldBOtJkAT8PeBm4MkaDKw6jgEpCNUiYDaQ
rLQzcbaH/NBjvI8Fo/S4j4wIE38aTiFWVUbm9qLv1gNVJcEW2C2B91AJiiWhT7ScNKLQMefypP9S
IpQ6IdUrlb7EarX9BUz1Iz7211MPEMKgwCuI12R2im7UUGEFExXn2QyfqbHdkd0JGZPM7JI0EcHM
NU0SsN0zyTX9Vl6ZfG4QJ6vQlKFCaJPiy3pBHc+i28gXkIo2NaC7CqnFGJ5EPZeYBXZaGlvadAnY
8s85Thko6W3xL1JSzCcqI3bv2g9YNWd+jfN5+hYiKLqIiNtlgQEUbhwkeuKJCVeGLHf1m36eQCF3
01G9TMR99q0EkDhtQxyUi1FfI6Y3f/pRnL3lTn2GBj5refx75b+ZpfZpF1jpT0U2W5cvp+SMe5M6
ur7Yu10pPo6Xp/JCO6SMTkf2x70i17X8GNTlpEwQFfv8uPtRSHLedG0Tg9z1hfQKQZlatjE/if+f
YQRgzZvEzwxp5anjnC7fhmyL2iWT2wBuKjvMVj8usr+8PBS2zbaDv9bLK38YHl3F/B/37NFrOkz4
WRzDFb1SWevntIHv0g8a0MR/sNCwNInU5n/NOQWkQKFbfDu8/WQQ3eSJD7F3zvEuoPWzd7lOGtxO
hbHPIo79aRQG7dnDjWnO1rSqZpdIOMMOvcmaAR1V2egT+6AXuZlfyyUkGmhp6gPGReUsY+mvodYr
Yb29eudteot4g2yZGSuS4jMLeEVI4XckIRarP6oBBMOrUvJxuar8LcH7UTGY/g7tj65nzGjvRjqp
foOEd2zcy7XTxxGhkbELLRjJT13kM4SrKLUSPJrKb093oc7C8MBPJ5YdrEO88VGJIfoBgLvuCrQI
YfSaGIjUXB/CYhi9B18y9oFJXnkQe5iA35dglzzxvlgEbwt4xVVTueU2vSiI13ESmuUtfhcNydfU
AsvqlI1eY7x8fauydhHH8Whk/qEwFzfQjQF8wwrG0I5Rd1g48pCwlCcBcspuYwh4yxKr+W2bs9SM
W4GzZthpOEOsxe/DSzhuY0T/WIA4xxoR9U7liSNJ7O/b6radZ5bCK/q7kxiBHXOy7xTIJLluEO20
4RdYuSyOX7mMG5gODSoop2SGMoHstrSo9eFKUsiHKhbw90/MXsa0TdoN7/7cl1kjiMXuByDXKyjs
qir8iOFAL8vyyh7+2YmSjj9Rv9HUvSDidcoOqZGZqiQbRfrZ2tR3ZbWVlPn7KKXj0liPzpaqlZHj
axBUr27ppTrV9ysnVJVXFHYQMnSMR7ob6JoKf/8kFda6f8PycrjH3SkGsPeXyj6PHbggcifnh3md
Yc+7Uj9jbG6GwMslKi4kRSKM1nCQYKGFneknjGifkxCSA2gpr40FdWnZa/zORjwLMvu1HJqchG1t
t8vD5YoNZkqtt2htXJyK7hx16eQcB+MuO4P06XU37DUztYnn9k+rkqDUbgMtJbAYMxzgZlHG5VEL
uIuArC6ylNuUHyVzKpwOq3CN4fIfW6CDg/6WsvZTOGVD6TMMTeRnkUGo8cwYWrLPN6dWYtYF9miM
lek2I90Jq2yOeyUJc3ZkIea/z227NlDqACDbadvh4SFFmAawCOhlo7r0U4uin6ir2TE7OjUkBtbd
DbTQQ2b+dhDyQR0toPXeg8bZcYH6Q334SiDLY4xLuX3rJZhVLsGbRMCudKm2czPc7QpWJeEyN3vI
mR98izhWQV/j8zJnY3VR90t1O7Wh3tBJtvFmjc6nnUdZxeoIcILX/dG7nXE9vjGhDvjAnLuE64X7
Z4CdpbY25Ii7zKV09w5odN9COlDLouZykEyfwJ5BltiU53lwwHPWeaHIhHBvOGI+xNFu3ZB9drTv
JUyDqE5jZ4ydMC5R2E9cLvTBYVhj0IyTwowV0Lyve+mPZRYfkapxcytUQyIHsRngP4uXZ4y84lua
wnsrC7T5G+ckvH0L4iLKdhxpOGrRdGV7tGSs2MTw27sd6KnJJM7JtojnT+tt9N0GTrBYCfdzvITa
8CeJaQxUJJ0qxh57IMEhEu/LczaUC8019Y3yFDpvAqmjllnjcrLzfnKzEX44gLs77mLaU9M/UgW/
NMZ0uEZXmJ6xIOWuqUSwE7pYv4VxHfczKrOBp92JFmQQkHyZyNGmIbQoaoX3g269DOgOmSTN7CBt
kKhuC6Dfl3xcOK0SALQ4yN+tONNFLtWs3kawlMXiuvXK594aS+XytE/q4t1uVcHkrSQKQLeuDlA+
Fn41EYeVNgXT7c3vvx1Zzc+42LRvWOTTwE1w5QZyVCJO8Y4RzSd4+zlQkwRdapdCZgzndpwKRGDm
xIZ9ZGBR+/R9uFxw3UHsjPmVsbsvILHQdHFoY9szWsTVMrUL0N+6/3PU9qqGtvL6r98GjD8fEDNx
aXsx8zwzBV0nPo528Y/NuxKp9yMCAcU1aBdYxEhwOrFpBWE97l20tvOs1h0XHYNf7eWXyb9PM0zR
rT1Dg66m1JuLWDAIi2oKBu5C3VAkYcriCIlp1wV4Ri5bDKXghqZclW4gsx+GvakUB46CHaB59wLN
G30/80WzmtRtKEJTYm8XfYGSPWGdD0p6Zbs95twDfBeXrUwvlqRZ1MLrjxJ2xcpMv1j49AmxyrQq
ebhrKWNd8OEUmtp7Wd4jmx1ix38PLx2au8zAaKJNRlmI/bc1CvRIV+RIRGBB6bZPz5Tw/Cbgquf5
7aycL2FPyFxLk4ISNtYejKusKgtqtspfA10JcQraNX3rafT499q9vZ0PTHuPgSRUMnwkmemHIwf6
0saCIxWCBv+YrivqM6GrkRSvDCyh6dsV/2KjcgVZz/7DtNYH7cwFsxh3Jns/6gIGSWSIKzNukbb3
4caxDMEhS57haLzSg27L93F+BF1z2o5cNTfUdsVc9UQ5C7MTh902BHweNOcra8nPWDy5Xq4B8m+A
Z8xpiJBlG+I0DLmVrXG4tzX0ktg9eSSayIsIbfhCuoyvR8sOmZQtzzcMssCbZfB5j/LTgSBxpgzr
lLZ78FIJz1rgnAEq2v6BMSv61+gJhPe+orRenVRUH0j+eLRC6keewO9pvJXskh+jOhEnfW7SDESN
9wi5DGHjkLQqIBC7CAIcI7GFm7UO6a5lg3FfD9yeFPzPovh1hCTKcIEYb6FvH40GLYWms2uLWkf1
zerC+ED64ICSCyoB+aKQbOgTRZ2LpLoVjkh+nWlx+V4HmJavC0LBNKG/7SubT6AvC5MUMOmwTURY
GzepqlbJIKyOOqBqckYFeUdQLREes8aqtKNR5Us3OteqrMDABpmyh5kfevETd4euAjUHCC0H15c/
+kClDHX0rUcvhw/v+J/nToSFt1EsaXEkWRgJHyNHuTF0W5R531IyQd3MTFegDS4YqxkUyODGixCX
lw3t9yrGiehKxkcRbMDytrZWXnbEMRKDaJH5pgPTEyz5DW0hMilCMYO89T4vqwgvGBcq2F8S2U2J
nhx7Ppg+NhL5tt+B+5NygxLl56kYEBZ9OF8+zTibgXlRBiAs382MlXOOWj454qDUqOipDQ+3XjJa
izLd7xeERbd1MtfAH2m38g30ZITUbb6XeeLzGfodqIPNTd/sS5OjVw7PbeA6eOHOevH6LRKw4nA0
69lFJhHF953iXWXw6YugyC5DkTrpKJU7T5RUcfTYlMPmJuKd3vvIv5j58NBmFVhGEGDzzaa2LPvi
SQa/gSwU7Cni4INoNjA5x7TctVNNjTNgIavz2L4vrLvVtkXFqZVJ/izHZSbJNWz0G/LLUsAZGXVq
nDcO7QqtRi7h/LKl7Esvbo4UinSXCw1eCjfI/RDkDorT8IOsaq3vSvfuXd3iDo5cc78EUyIjRwFT
k3dRu1zHE6ajfPj4IUjjWa14wTL4JeDzXTUEmkd+LkZ+Fz463okieyiukSXyH5rHPHgzbTkHuwaB
vCN4M4FRCeLAQfKtiVnJY1ZcDAPICD+kJQ+iV/c14MF3SoJAqOmCAK10ROGEiJZKePxgLCwRzniC
LDAjNflIfgb7yc3PqdeoPelCccNiTl+xZ65hOZE8M2q94zkqFoKONrU4nASvJBT4tWgOs0VkDtH7
5JM1dmf0Ug4ZPCX13Bv1sbQFTuMM7Og/FiC9cIPENoRgT6vsyrkr5+oIKsbTCMu0VLm51vnnuZL8
HD6zvZGI5c+dvPkbwCS79qP2qVvvAXHNHdvebhadeZv5mib//5y+ycQvYWVmLe2i8dMJcVCsyI/E
sKC1keJTzf50joHgjhPBpwqQ2Yc4YaBt5OEW8DlL9nTaNN6cNKmlKzDNVpzF4IOGc6PQDoVOZrZ6
Rf3M6FgkNcrWmpbR5y9465zUKxCuVvkS5R1NZC2j4EG92ikoq0fkDyBbJIiQERN4a0updWsX2yED
UUh/VlsXzK8n3k2/lVhPd18kldbLksXDvNk2K8loPZzqc0IekGa3bkGO6WIJdCn0pv/zGluNiuGy
3XsQKJ+itt3mXxOqrLxD4wjA9OOCA1UX85e1t4i1gfYHyzB+YIz88Nkg8SnC6Q7Z9ZWB4dDfhkAL
/fQzp/HtCjsNMZPfTG+gn1Y9FDT6aZsUb+oUlrqHIzTDlHkq88MuOCycFXEO1d21wzCT/Y5X9uMP
9RVHy0MkmUDaBdYKtPhnoQq0EDCr7sDWQYkkIKmiIkLynJZzYNco1YKRVcsvdBa39NgZTkQIZoou
HWwQVzID1b3iQSe+VGlamdSJOSWWzXktvLrytUcKtLA88Qorbz3JEprxjIb+Tmjxw+Kkq1VMUrl3
iqcyJxQPC5mpC0dafX2KA/ciI1oEpddYSGHYOXqPtxY9antsBMzsUymJXrpYADXsV+KsNx+zBiQv
t5zzhSEGQsXJaVprvGjcnQQAVzdL05X/S6RzVN7obkQAhHHHF09ZygCt9m52DMkAogayvIDH7F9Y
HlEo8H/CjaX96EbZ6ZO4UnnbKhYiPww3aZQlwcOvlHO51boQblVu9oQbo3vPVscZWot5Z8hXQDou
jg8Hv/fNoGwHobo8UiMmVz6wBCXCKUq1d7yo6kxvy0RnXnrJLC/cxi+iM7QkLgPtxCcMSLZsLbSD
RWIX6yVAxN9goHrNoyJfkTc9hz8pqHn2VmsVeLYHGKcY/qCFAhr36RlvFMfl1IJAEQfbf1n/LUSP
9nm8MucX5nyU9s9cjZ/7bjFG8wBg8ygJfXjiFRxVOI6qKCRlNl3nt/sHJIIM6+0cNvpgFtXhoucI
CLe7P2+DAAL/OGv97TyQftFlxPEzw/2XvG3SV8dscKhfa2s1qcV0Msi+5whlFtc8dHLb17lS1HVD
BLGeVM1rub1/+NsyGeJlKLeVx9G3EmpIdgG44G51ak6lvFuZDF+VLm9mQutRv6XR8hX3TE1ixnaW
Knbw9k/H87C8uwQy3goU8A0GFdG9rwb63ycOiV3KvQ48bSZ1IxTl6M+q2c0ir7tPnyewwPLDDGKj
Rd6POZnI+6m/FwccJlTTniO2a+pPaU5MJ5nMf50ZqAhwO3NmJVivTsFiOrn+YnZBW4+H27LjnOD8
F4W4wO3TZWgCV6QsGoeDeQaTtrfyyNv/XlEYYA/u6+G9lyNlA6jK0E06qsXQfC+1ymo9vyotzjHG
BHEgNfMUR2N0LqtugNPF7LPS+4E/ghbkmxgikNxKNXlN4kCqk+/SVCIhCgLheRTlH4LD9ZfMUGQs
K4+uMyAbPMmm+4TJYUNobnusbEPE9YxDvBPlR69xxgwlzeFdYDYAEaNcJ/0VW2nzkEdONjzSn6YH
uxjKxwo1aJaoe6vo4zXrR/uAyXJjbBZkPvMIRCTcexAghl52tz4/CNOsgZHuDSACB2vzpX/TKNz+
rsd7EA7foOzIc2bnlVZj01i3DZT2yrmlgwIoS90a1wSGQPaZXzNGaUf1/FxKRcjRbM+WzTS3Qmxf
HGqohBfBpQHRuZGuqiASkAfgqePyUrjXOwNQzfFpHgNwu5mNVPvKIz1OmlHld11DxpejdlGYFads
h7B0/HsF+LyJDuoDaHF9AVeBmCzpofoj7fYnwl9se44h+pBV7elhXUlTxsv71tlHVeNqKCIQ6t37
Ji96fGOof1HRxl5TLUW7URu5mRFamas/3kRwlUXpzojiTFU7ejK1/f/cEY5jy2n/L5M1Mrbvrryo
JcTI42DkdJkgcM9Uo2fx/QN4HkL3SYtESitqTCOj6JcLOmJEfShqk5pY/UmykqXkwIbkPRG6zS8d
0tp4Y+S5R6slHT/epikcbcvIq0I9c1UejIqitBbNIyVInxTWnAp0U8PAXY2D5mmWVuHVm9+vaIoM
GGQTwUXIfUYUa1PF+SA7iW358qvWq+cXksbjm/yDj1xGue5nAR6RBsGAqjVbOWxIHhEVUZzlMXEH
bOB5jVHNinknmXetf1s9t0860lnNDVsUViIDel5QQaUEffTolpgxUrvhECXN6rfgTonFO5Aia0y+
tpno3LW+eWLKSLlmAqo8x4euvN5u97D6as67Zl9V+VmTcCad+nh5fmsLg7TUPeLS1BRh3UUDGACM
0gujFtZOhR6hUQBefzzE7TbPTX+CrCFTorBy03+bPufWjbON
`protect end_protected
