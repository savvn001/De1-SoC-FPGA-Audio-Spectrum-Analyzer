��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjH��mR�L�J8���`	774���%�<���/�0+�XP��1?��=bC���xk�J���7���[�P�8��h�_�$�[0�^�"��f�����"wd��`�{�ʛ�"F����8�U#�S�|{2�a�[v��RhE�Ý�;"9�9������<[Sh'�/8��%�(�A'���-���^����H[]�3$i�T}<�zo�+����8��������x�H��#ʕJ�@ҽ�ipP�r�G���w,�RS"*����SB6 )9X�Pr������ �[�d8כ��
Ng)�&c�RO�<�p�� n��V���Dm�G
>��8Vgk��~`̦��
I��^����Y\�\A�k'M��\/Py 
ҕ����{_!}§U�Kp�3��X�1���g���<!�^0���1)8�Þ�� �-���$ �r����H�6q5ۍH��lcC�.:��i���J�q�p'�A��)s0��'�w�Qh��|T�Ɩ
�:;��xN(�U���>⁺��{�Bk��BE4�\L�����z3�䑵�-�}r�����>3��Y8w��\d�V@���/p��ɻ�7������,!�!��;m^qg���M��C�t���'��_H�I���p(ֱ�,�:%\�>"�C��J*
�q��!�MDVGmCO�R���t]&�G	h~��H �n��H!�!�}�S�;f��;���������fh��r�=ޕ-ҏ��I;{�%�wz���/ȷV(���#N�(*rc�;�Rk��p��wT�;eS���M�h�l���`Ϫǔ�0��w�U�[%F$ol3�іv�]�B�	��N�	�(D�*""��-���͝��Ν}t�5g��V�Q��ua��d�., �����>��E�>SCA)ɞk��j�������j�E*{_Tk�/b�o��ݟJѻ&`����h<_A����c����V6�M޳r�[C7��;���v@��(�^xl(�%�;{\��	�Ɉ,�8�2N_�������KP.��a��|wT�d���+ٶ�(�GIh�*�d��1E��a�S��Yp���P�����en�[3�3L��.Q�%]����� �-���{�����r�J�_@�u���k��J�>6��ܒ�j`9`?Ʒ�C�����<C�a9[|@��!i�:���[ɰ��k�ͽ9fƦ�v �ZW;�^�Te4���Fu�A���f��G]����kQ�#��|�D�H���>��祓���>&t�">7-.����þ���bJe=/��u1{����gDԛ��MR++�<�V�2�e!yP��+�D7Q<�c(�S��X�w��r�l��E"�h(�|���r�^C��b��Xy"]t&���a�ͳ�1��(b��Ym�e6
˴$���LL�aO3hm�RA�J���{l�w��
J?�o�3m���������'������ݍd��8��+~�b�
���������H��A���R��m�/q��r����7�^��HꂨO$C�k���L�6��c=rg���Y�ߥ�0��Ѫj�2`�9���|��[�:�/��d0���浨n�u�H[ӰE��Ů���zz��J�/g�e8m�Jz�3�V�x!�-l��F
QU�;GEK(]��"�j��w�����tT����k���(qԄ֣�9��?���cCB��.�}��q��G�3�d�ͱ�|�eH+�`nFy��8ï�?�;��5�����=أl�������E枭�ͼ�!��F����Ƒ{On�Ѡ񳡙�lz�1n���I��o,� �t��9K�mӢ-G8c��ab�9+'hRƪkO�3a���W,^���v��֔�I^���_�b�::N�����.�5Lu��%��3��j�^�>ǯR��|�D�>mvP�E��A�H��Q��0ᥓ���Ԏ��ڑ�m��D�9���O��S���r�)�ɦ�a*atz�@%�z�ۙV���-�(S�}9�zԸ����1@�נ��L�l���T��jr�r�n���ކ(�J��R:c�՜�.��ܲ�@?̶41���&87�9J'l�6���5��4E�� T듟
�^W�#A���d��U��$ �@��"h� Z�MY��(z?��`]�R���b��WZ��"K�=a�m^f��Qg��r�S��Q!��v!�y�zW����aN])�8��T	L�_ �p��Mz�u��9�JD�y_����k�H�z5��T�A��6�fH,Kp3����p�����I�I�DfrL���9��ØA�*�fb-��_�j��+9+���)9�	��	�\#����8S_�m[����.Ӝ���~>=jR�Ax��#��2����Ԥv/T��ZǛ���;OB�Y����/�v�Pf4���4�7i��e� �$O
�*|[/P����q��q
+��6������}�;}��O{*V�H��kD���=��ևhbXX�9�CPU�Z��������P�~|I0�����H�@��d��Ә�ǹ	��q�/\Fެ����_=�žּ�P��Z�GZTvv�2�%	�[=0�#�����9�'�ٟ����UK���\d��BVV�����=ݧ�n��ڨ+~�N��J�Nu쑶�#:��-د�i_������m��(�,ۍ� c#`N�����>�ܠK�p=��{΃*Z���2��t�|t�K2��l�K{A�0���|^��\����jZ���W�4C`�e��l�2���~��l_M�c���:��m����c��6�>��}~cKЇ�z������� �w/h�|��\���.��������z��Ø0eB���" :����m�Z�U5���/����p������d�߮����A��'1��(V;;b�+YF��]S����޴*�����eg1Ae�eH����FJV��m��	��(�t��4�;�g��W�f��z(�z�R��Q��E�\'�����[J�J��l6��Sn�5�nJ,F����hbIG�Q 8���;c\����*�=���� c�_AA�P*8�n�뱾�k�vBU��3�[�>�T~r�.�(\���"\��<�����m�6M4`�WW�0�Tx �j�����w�6T�G�yޟ�j`���rs��Ǉ1��
*
9:@��>�ZZ����)� Ӵ�9\TҖ�k�U,��@���{���M�L��ik"�J��Q�0&�fߒ�P/�L/����2�� @.�����yw1�/Hќj[.�dP�P�a����XNHY������K��LD��1�PU�s4��}Q:6�����=.�/�{�㧐ב�{�X���%J!�M�-��V�߸���S�����ߋ���/�D��J֔��WA�d7�<�wt`��6��ѼwJ���?T=��OO���]����K6��NZ`�;*ݔ��U��(���F㶳�-�dj9_g��m�6������>b�]� �B�vXЅ8P
����v�[�{��������9�!�i��iØ��h�j���1H�J,���8]xq�4ѢS��`�����b/�a�j;���� �~�o�נ!B��'���T����a:�ig��Sah����?=k��)+���	$�\ �{%t��hM�i�T>��Z���a��N0�����VҒ�/��:�Ys��k�Mw=2AH�xS��PM�����r}���{���'+��_� �2�#@ݥў��\�J$z��C𡷨��1�c�L'z�g��Nɕ�`1�č#�� �v����W{zvȘP��A�2H�{�����]:�{�����J��n��*��5����ɤ4�#=�k�M
�q;��C�m���`3>���Ϯ5l�F�LZ�����AG(R����,'3莪T�OS�p3�&aF�f������.Q��2��������WC���u���A��,T�(�y}������8�f6t�}�O� F�Fm~V��-%5p����pD^�6��j��Ȫ��Z�+R����C6�8�@�.��c��=�拚�Z��$')!�A��H�h ����mܔ�ĳ�;�{�@ j���M�	�G�c�'y�n�I��?/9���sR��c0��`>�����z���a,��_L!ݳ���/n��U`TFesc2�������R�Xw�z�JW���lEs���՝����a�O���&��V��~*�v�=E0`O���;�hv��)J�3��/���ݽ#K�'n�I:�z��Đ�S#!�!}����-	[gͮ�:�3Sz�F�C�܀���eN4}�5�|���Z�Ց��)F!�l&~)L�!�l$!w��R'�'D��8��rF��|�����MQ��U���[�5�������m�;@R�wD����
��t킺KJ�jPSC����w_�:����㯂I�e�sǣ��Ҍ�`��+��<O���rx~p�����Qx�u�TU�ѠBRKe�J���E���U�K�1!s}�F͂?�ݽ���	���44����¶qm��!�Đ��u7-w���f�p�-�.����\��!�
!��:��c�H<���ڎ������J�< ǰ��+�o�B���҃�kB����V,pxtPz��z�-,��It��Ó��f�������^�|�xN����	xX�{��^o�_'�����ë��g@��q7nG>�N���%�Lb0ѽ�'����s]�=q�\y��A@#|�U�I��9+"&��+�Qi��x���(��7�s�;���ky�J��V��26���jV"3j�T/,Rp ЀJ�/�����������C�;�!�"n>ԮI�(.*�]�_�����;y��=�~Bv��+��{
k�o�aP���^Wy�Y�M�N��^�v~��uG�գ8 �_07ߵ�P�Φy���6��>����J/~^�4�0���8�P�-��4u�2O��,�9���ݹO��{�j�CEϴ_��s�y�����3UQ�U�h�^Ȓ	�Шd3vR�k��W+̸����iH�
/���
���u&��~����@[��\n/�u�.yR�x=�$�����C��b��\ ��;r����ڴ�/;QV"��"[0r���c�o󁻓�8G��i3�!<8��}
R�/���b�?v�p�Ƙ(#+K͵�����U~ȵ/:h�_�(ڻf�j���a�;�'�N�h�8^���`�,G���[�&�@�_�&�'8�����+ZV�D*{U�v����6DW�c�J��-dR1%�I��wD	�N��HH9.}Ex��[�׺��3��-�v�%�
�i6�(���M�s��E>�ŭd�������6��թ+˒�j_2DJ���\���8��#�R�/jB�t�I_���E����$6qL �-�6��V�j�n)������2�J��4����6���0��qD�	��:�A�`d#x{�H]�w\0ۼ��F�$��,������h��Q�Ъ'�I�2�U�i�nMʺ��̎S����sm�'�יִ���2`څ����(C�@��pNc}���	v3�-,��2/IO������_��~-�*�w�~��ӺQ���p"�n�_8��p*hYw#���P�O�Ӡ㖾�þ6��䍕����N��'v����:a��<�*V7`�(�ʂ�j�����2-�m�QR�~�m��q�F�h~�2
����;ӷ^5�c�?U(qZ> *��Nu+gT�޷�Q���{<�)�n�Z	�tZ�g�����UMR��%�*��{[G7�r!��T�8��ũO�ʵ����r,|�9����f ����� ���ot*	��h���@������;c\�"�9?�^}?}|�7��J���8]��Q�2�Վ���R�̺T�}�3�+������-c_R(�i �����z�[���+"�+,���Mk�n.��=�;�����_S��-��=x�+�Cz���Z4��-=�{��e��8U���#�������)���wN}��MR��*�!<��3C�<"����Y��=7�mvT��'�r�$�n#·Jr8�&�p2 �+�Z7F���<��rH�=��j�x��v3OD�`�o.$�ל��Z2�_8�#�w�O�σ��K279Fod?Q�f��Y�B���O1����8WLHu��15΄�0�!:sɶ��Г�Ԇ�V�U�Y� ]���3>�r��/f@+?�VN>�_$
�ŕ#6{iUo�#T�0��g�M��q��C��O����"���/����,�����U���#�w��c�@���0i�6krK�%j>r�N��C�f�V5�F�<�	��}��4��@�$�σ�4�v!���z���D��	6�w�׿h{����K���"�4�1X.<qÑ��Y���(�$K��k&Iشie�/�ZC���RC]��u�O��1�̐��%~5�ϟo;BJ�p���QI*v��}��Ƙ����ť4��m^���ѕ�&�c
"���v[�0"a��z��.3q�0r�"�\(t�����X�z"�yg�9�wJ��j���q��xМ^y���w�7�J綄��!syJ|ʠn�-�����ȨVcż�?���,���d;��Y����p(����p����Z����;҃��I���v�[�I�:�q�#��_J���ൾ�d�n;�D8#��}P3�^R=�#�U�P���6���3RӍ^�[6�0�4������h��B�}hu�qD�am�,H����	�z�1ё�HE��r�(����^��5g�ϝ�i�b�!�W11gt�*��~]R7�7yS�ܬ�Ƶ}�P^�d
���vU'ʿLWK�	N���lQj/�����\Gj{��C*F�ًGC����g�/CI83�Bu����5}���9�ډ����k���B�����PE�t
�Id;�W f|5gʳ��OYn�g����^�rꔄ��$t���~�ͼgFϑ-�[�V[eFдD�6'`�ya�x�H] ����V\��K:��L�ߏ�`�J���w�$�nBr�3S�mmڑwQ��V)�Y9��p��w��W�+<(/ۋ�����c���
�.���`�����Y	S&�JMRh�me:��"O��Tc��{d�5`D�\^ JYx8R��ͧ2< �M���I�9)�z��%�?F��U��s��H����y��,î<�6�1q��~G�ZW��-�CpQ�!T$��(�u�O>����g��8����6�VSDQŀ������A��c}(u)3�4�r�ܙR��b/�m�@\o�]~����U���Du����&4D��Ǘ�{o����zFN��/���p#��j�u�Ґn}��_�rw��3�<��.��<�����0� ����f�5edU��\{`>��Gt/�r�$9&(��uMm6C�e�5"���b�#g��|�Y��-��e(����~��Sv�5S�D/S|9�,��������X��;����2[�藭C�6�?�V>�3*��˷�)��tU�o]tBѮto���(E�4�?��8��?���D�wԬ��<��`f���v�r�!I',$������V�E��l����`�\�v�������\�.��v�6�6��ݼ��t�C�:����:�%{$[����E�P�.S�����r�����֘QA憐��p��e�޹b�bE`��ElP��n�+5����D[p5[�4�죄V7H�u���|5Z���۴$�1,'P53��S|<�%b-������c��J��V�>���t��Q%��Rd�`�$ۛ�W�i)��pr��0��a�I�ߟ� ��K�ڍqʖ��EJk���p;�#X $5A���!���8��C��ݠ�Nt�Zjqԧ"C6�d}�D*�ve��%|p������f3Z�F���U��N���jO�/T���3�r�{2����6��-��@�$[��S^�)6��tl=Q<	\�M�>T�+ZD_�Lu ��X[�.�x]�g�y1$�J*��H��&Սmq2�j
��qO�W�y�Z�4�ɶ;���r4�D�Z��i��p��Iy/ώI7���V��;��gȐ���[�XӃV5�^�?
G|:������זR��h���H�x���Vl���e�1��v��(q�yD���t00IM�&I,<z4c��Ӳ�[_����Y�Ĭ��aۇ�$g�.�W������Oݫk$��Hf+m���3b<��/�4���!9�F��,�P�(�o��޿�I�R�X\�X�-/W��P�A
�@�I�S4�1�>�x%,n�M��Ǐ�4�80�i�x>!�Qɿl��?@y
H�}��̳,&�;=���n�w��K��n��R��ӌ��8m�v�Bx�)���ˤ��C���~�P�1��U�32�P�/��|�ͨ\I{�tx�!i�)z���.xv#<	c���*�k[�]��`<LH�n}�w��3�{P/��<R�a�ջ�ʔG����i�$��v؇{�lށ�ZujՕ9,���R7��w��Or�׵;��j[*f@��9�a��٪��_�
DެX�-v1Cĩ%/V�Γ���̞���=�G��D¸�C�G�z������	[�gL�n%"{*,���É5�[R�u�J��6�D�XoX��
�e���O¯��ɚ�6�#n�E�r��;����iX�%�$��:C���J�3�~�p�#G�q�%MT���[�� .�N�Fl���r�4,�<�K���А�#16�&����)�rrGE�Z�]%e"��%�R�N�28������=�c�(2���S��5�Jj8��66�
��r�a]�Y%2����d�'��hb����PN2�SY�o&�lC���;�������'���h�yA����	��c;eL#@T��o8��Ǥ0�~8�_�i_�f�N�5]�"��vv������i���)W��[��g��#<\���V����w�2�j�rN1��I*��Mp�ap�lX�{ƹv̈́w���i�ZD�3�#��f/��Y�o����qC�;�x������|؟\�(�\�	Ia�<�U�i�LM��ӣ�(��aN��}P�D Ĩ��a=�R�S��F�.0���X�?5���h�����)4٪!����݋�W�Ҍ��6as��-�\h�`�`����R�JR�.����JH�G`�O��`�,@����et����JgQ��\��|͢����cK�)��6�ь^!�p�u�OC��ǩƌ���ă~�-D��w�@|���?�\��1�J|S~�C$�>�P����;ł�x����&�t�fIOF�9�,5��|���O�^p�A��ԛ��[
/}���|q0H}�aU�T2K���jH�l)���Uҧ�4�����W���h���Wx>ܞ�� ���o$�+����[8�l{���<H��.�Y��YGZT	D��&���d'k]��CbA�����<�������N�#��&���}c�L���$<"y>��n���@\i����`6��6����m�M�9W{&�W�X��X���*���?�<��8a@����	�/��:x�F�}8�l���!�i����R�{s��Kg�˶G.�.��3f��Dko�`�~�Ќ�,�8�%!{̻u[�r]MV��W�`���;��t��I�M �6N�e�ח$����DW�Y�8 �I˭'�8��G�.Z�rW*ױ����@���E�=�`9��S~xdc�D�m��6����ZG�}�}�$�&��<���ҥ���m,){R�i��E�_M[w�")�B���r�'Q��v���0*sR��V(Ƴd�p?|�۾�Z�?`FX��ޝ"'^P2ZZ҂��D!I�o5�fB�c������#�e�&b5�@|<��p�feWh�7{���x��8Q���<]��-Za,c��.!]��Z�'��=K^�v}� ߳�:�M9'g����������&�G��QiҠ$���<�BTc����rd�*�^R�L����%��?OkD{ �R�4_/��W�ۏ��"���f��q�Ss7�I��0�57P{?�s�sX�fb�7���j4����zL���4�����Ēg#�����ڒ�\�qg��D!Do0<� �)�e.J��/�E�\`�*������{șXX��Q=D�77���a�bطs�r'�'c���ɫMb�r(�nE�|t� 
 >�"�Õ8�I,&KQxO��E����������d��4t�oMȌ�kk�fO>�|Y�]$̄��H�Myum�-���})i,rz
�!�Z{*�֘���H
�yA�����.$�����P�U���P�dm��&(C��[\ret���z��#a��6S�a$핹���� %Ђ��Q�bm�w��ar��) �j}����͘q�B����"|?�Թ.Ȗ0W�e��	Dk��z�B'�7y�H���bJR[� K�E���Lb�-�:k���!ӯ�Q��	�R*_�(��;��I�-�B,�(�X�o#���9X�;���E�f2'n�j�
Ӡ�9��ˢ��i>�)@��|���K�B�0��}`yXMEQ��6�Gc��ֻ���&�Ӿ�^Y�.}�n����_N�W����E�L^����/�`W�R������D�+hi�|q���a��df=`�T���xy6 �'����q.���K]�!I��-5��r�zp[�Z)�:���$��ϧ�~��;�9"�E/�h,���x�k����\�Ë��ql����fd�b���kv��|��V'Yh�J��,ߵ��t�[U�Ĥ�=צ+��FqZ�]��ױU'��['�b$G��%R��_:H�$J~ɜJ;'�<���$$Z�s�>(��v�n�#?[FU=�M-&m���rb��g®�g��D���4ݛ.�,LI'USE��Z�QWjC�����ԟ�%� 6�x�!��(ȸwVv�_�`A�ǯ<s���R���%ƫ�QŢ�JA��5�M�z_5`�+B�桬�ڲXt�-8nB�ܚ��`e��t-���96��vG!sg/7�Z�,PP8�<��Dy� {��	5���Ժ��>�k?MX}�ӗ-p�׵���D? �5@X�2_���'����Vі��s|�L�i�1���m���Ւ�j<f�bY�@N&���6���7Y?lS��p�(h`�s�%�zU�w57���	���2&�4)�\))���@���<�ń����̆`TUd$P&؎8B���j����,mAX�=
�i�.�Ξ@b�^we6�@]�b�x�����e����	,�5�}'RV������wQf>�[�{���b~��[�^9/�2���O�����Lh�g4�e�(��FvsIU�A	�#��E��Q�\/E"O@����&l�[8���K��C�����gHgẂȍ���V$�PJM�]�g��z٤v�ȿ�?��[�d7{�����V\&��y�c�`l#l_��K�d�*�+�}�!�R)<�:LE8qi)�
�T��j��h��k�S�/�jLg��#������A���y��y�G$u*���lzk�+9=Z\�d@˹h?%YȜ�{�Q
�x|M�C@���lWF��餸JԈ����<���_�Q�L2�Pi��g��s�|�*���Y>�\�	�j&P2rY{���L��{��;�1�p�lA��$|� Kt/�!A͎�=u���N�� ���O9�����7�
X�����w�=/Z�+�`�1ϻ����E�rKj�r�����I��4�Ľ��Xqո��>DMxY,Ǡ��Nw�?��&��0���!��~�"�z���I΢��4[����W��`��󴐺��