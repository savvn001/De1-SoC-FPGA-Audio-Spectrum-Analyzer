-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IW491pAmGTIsXzDaFc4Ew8kTuIHse+zMJ06fba+fTNQlDItQhVzwOJ4BgDHGmvKG9zpGV/HxByvB
/nBbu2Se7HFv09FSqURYkAZbo5aJsViS8IN/ZXzzqzj2N69gXAwT8NRmllzr2sV/9byieFitVnZL
+CMEjPUZi6Kv+7dg4UGKWYOOU/4i0vRuIamp3fBJtnB4jskAJbLmI3T99yTm0vECUO3KtMIIY6SP
3uanjz6X4vL8WQCjizrx/Gmw3Hrv3wVtgi6BT1trepqKWAPgsoMrEnhI7N5dn8sOEML6hAHno2e7
qvT7tBM04blBX+d9WsjoAf1kxHQvpNJEa24PRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9600)
`protect data_block
wEIjLzWs+d0TMyTrUHsJd7ERJug+lhVGlgEHMjr0oyfvwSRGTmWdLGxesFomy6lhJhacvSAriEfx
f6JxzRr3dk2r09KACufacl8Qn92LMCjJR1xdP/ooUrjOlIVBjytuUSf4ic8wp17u4sgDH/06a0bv
Xu5CzIBkiXpNyfO8oCsMHDOEghFz1vRZ5PAHBvFpiZXMzaS1DSqDG1miRphaC6rv1WctDllZU8b6
GzIf2fdY55AC2vtMxyOwS/tBixjdc9WHZPw2r2e4sl1rChvlRt3KSzEprfNBLpDPVlZm5bzwkFnD
fSbwOUsBujte2aU9FOprpoRFxN3Jiy1kvCK0GhDFctnqU0TJmzHQL7rlfJSaJ0gPoIS9/WJKqWXJ
gm5J8yWhIXBhisswOnMhuU2Kw1q61xTNjiHi2DViSsbTNn9HQOvHiTGMwDhS4pu//pos6qgCBcRP
QFwcGqInoYheGRr3hbNAlIstzxalNgNbGrOYOyMZ98xMmXjZr0xMljPzklHG4bxB5R5gzhz9zHxv
nXNlqDS3oISEnC2mcwpICcHK/W0OSHVK+Q3SoS43UGPt3xBO1Z+k01FZJOdFPC53PRe2seknwGTv
oKbn90Vz9BiHWH1ExIEjl4cZF5RTNjPII11vxVwsfV4G7fO/Yen2OD+7ekAK487ilfLRK3Ca7wAz
FjvZzPjzpfiWugYJYAWgCDkKuTIJYVP0f0rU/okijmnPCEFUFWcU1elxunl/mYERqBQ8dEpU12uO
0CcL6frTBWoDw4HhG9oDu+2HYG4OIeI8b84PDslsXrdqvs72qaLsOuAY+/DTvUhXbQbzX6sTa9MZ
LXswUCT7iX1bNvNE9Ck5NZaS+MLPHPHUkJExrGEYd9YNLU5uH/lBJIDCWK/5ksfa1sKhF0HEDUy5
up+jOxDB+NTrxz4Df5d57xSB7zvGctdy42MhBDWpwGNad4pjhceZtFXSTqRfUvb74wlMEoduhk8L
GF756GsjzZH13z1qPCuBcAD6rPIo1rr+tMva6n9WwdwaIjFKR2QBn7fdEaWE5T5eWRADmN2MqH8L
WbQaY13ydlCAm2sBTzg6x9LRrSDE/t89AxjuB95NX7wiW+XMm3H1KYUusgS1Cm1Fh9LE2NGb6kfP
Hgq+JtBkeCc6K8IzjlVNmFJRTsCZXvgNiAnOAubYsiIdMkDZzMjbhZ7rNDoi+f1J0CSSHVzJ9GwF
xyH+8I7m42/9ULFOn5pKjZzAhzHQMbDAdCNbq5eWAvEN4ZG1UJka+I7KYZzQm+bCgpivHtOdgt+K
bmahScvh2RyjveRuUWXLlrPtGfE7nmiNSpUuctQXp0OcSUnQ0eBH+VXY/tFMWyoO/XpiCvOZY7FU
kqZaiXKovTjuPtLPVL2wZO4h/JRr+WsDlEx1kuOMnCSPZfXalodi+1eDT7xMZZ78cy0DYsPwKSoK
ac34LficPvTV2Fx6CMx7QJx9N5Hyg8hP5Ca9meJfXZPxrVg+HufKSLxtmIY18nbiXJDshBQcB08M
/8e6JSpr74b/qb53/S69vne3DsrHVUbwu3MHwXQU0FlsgNHAWXwTvlf6GxfZze/kN7JQ8+6Go/sb
FpRpguhukjXS2zq8J6PaWJ3fS3EQaf3v3zAeA6F14ascT+WoQtqGMhWKD+3k27sFMEBDXPSTcjit
BlwLwTNM2KCcppHI01BjjuaKI+5zoJUwTCwqe2dtkc/xHpo0YNoKNgcV0sD6PGPoiha9qw2iIOdT
hwDav3ny0tejl3Iou0llbtAQ2k5PrDIgWo70igjAD48so2GVK4mtZWQ5p8lXnr2hKD0nx3/WAw4D
kC3W+4+193DNLcPk0VJ9lpi2pfqp8KY9TaNSrNZXzIc7bYpOg7KS7R1eQtL2ofMkh6CC5YVlTFHv
zAB+cwuynoJNiQr/NBxCeK0h70+uBu7HVtDaCPJi5GCcYdLDDZ+nhWGoisHxrDeiUd6LUgeqjwR5
RHFjzHbON+s6QQByTM0fRS9C7naaViD3DGhYosNPwE6vwX0H66XNpYO8KJk9hCB5C6w7TqcrJEDE
/KArzT+ADkIMH2/4mItCljpQf1rnOTUtFs02B35bAEuBwzsCNfbuhHRwHtGmDUAWfF6fnND6LqMx
PEeDh0NWBV48Sy3GrTugjgkb7VRikvT2H88J2X4IhDi0N1mmx8RyXd5wlaaLQxrt6DX0BdBDauet
r5jcH2zglN+5GS0KfsA6GpJ7ayAWh9XblelnGDq+/VZeiOozpLdk35Ea8lHnBzxxlCYRy1rQqC1M
kAz6nPho6+k4lq9c7iZd/cZK983um3yGc2sBQ/+VoDl6z2czG4KPuYIFslOgdZohx5MBXwIvaVbx
Xg6eH9e6ZJyZbU7Az9UEvc2BVlime/AOVK0CV561sLRU/8d/4cNaNA4bvEkiKM4yGym86+4moyMx
nk5CYAqHT1CER1YVLp5edxdKnvcCZvLm7EfeQXj2wzF2dNaSBB4OFhcI63YSZGBPCBt1vE0jx4Tl
drk/6JBNm2z/VYQBwslU+HImSVCBRWz1KwtOm71iP5kf4eA+E8Zlc4KRtaytl2qd1EWyAqpUemtv
XjbVRRZFKKxGAuUq44w816CXRXKRr8uoy0LpCb9bNsCHaVk+l6QcmMx3dHmxpAY09HU/xP3SmSYn
u/doAJlI6F725nsHtausVuq5au00gFoSoMgJbES784/Fk1PFDxCLlSg8KLykQ5+ffSuU4pXFo6H6
leJBy24wusu+tXHDhd0RTT5a7y0tBDp7c8zOrZZnCJc/OSzdum6DaBMW3ZU5g+5A38Ll+bjovJMW
94rqqIoQ5vyOuIbN3DrpQNpLS1HZR8mkPZH8SZM6CDBA/JwItKZcuQTW840xxXKuTrBAj9XtlKVo
KfOPpBSVjm6u+jgC6Ak8ZUTCduRh+P0h27NkIlcfGdVGXbkkdVmViwnOXnE9bdXa+KqwONfAzibP
pybJ1iJpm5oDSo4S1QxrYoCWe6GYXqYBMEi/2h8mfckL2Z/Db1cWFg2P0ZuFHW+pvrkenP5+keKa
k8wrGQV/Y/B9z5gtOokJzD99fSKxavDH2/Y5/j/MjhOOalMfxVkZOusCRCcBLb/9XnjCXHG6J2xp
kNA3FJE93bw+ctzPpiJaDVpE0XW3IndJnhPIk02qkNpORV7MiMxdHR0PMyVBTfGcbZDcK5Pur3AL
ahzlGIi/2E6oO02kiESAL5qN2ZNMBJ7jT+P6qK1qC/ywkb1BlTZh1sJmgQ7HVbYoFeSitWJ5C+Ur
Jfyf8TvW7pBaR29XQeiF1OfIyGVFCh3/N57hb0l5iwKYxOsVz+X8o6tsH1ZlYtJGcsF8vZWaxQIg
scIisuZcQBbZmYUjt8uB5+0TB2da0+CW+HBGYE/ECHaE1Kjy2tstGyzPXsOGvq5jRZ7qz7Fs/ReE
T2Pt7FegTkNO7ZRBMIQmV/fmcnCiZFJQnqqftML+OIfrb3K5e96goMNic8HiAyhzt7gSAUTGzCkX
fNxQIEzKg0S0gW+Kf2Xx01vOumI4kzaldRvgIwiJxAa+qXFNxHL97+hyYl89e9ZliXvIAtwkZZgS
c2aBQCAezBhCZFyN6CJof2aHIkeOp1KzxrkhXV7Q7QGhqNd5cCifkQI6PGk5wcGKsTm7eh7t2+6a
w4Sl2JqsGqQJrPIiwQrMS+9QwwT3r4v9zFrjvyl00BqJjYw4+ZaIEjUNgv5nvNf39xD/OdhLZ8OJ
FkcO3YhMws6oMbiGTxHskBOjzA64KWC7CesLOMIMEe5rCrMkqdHiAho8Fw4jMay+UiUnWVV/qLe6
oOqBNWYzXH8sw4Jdl8M6QyRM46RFGOyejalvWZx7++I7iY6zaog0Mf704mY4Kn0aC4dMLdefC7bA
DRpNY+mmU5YZN92zyhZ+78acsSTiVdAhNiZpLGe/zX4YKXnVjdAMvAAp6bGT2iAYZrYvs1fsG1xS
I2a0dSPI6Iaw3zlGd88fhCJ4ZMS2d9xxqjObOE5jIUhajr0cRKqx2IAbpPsl8lmrLHtIgUNtaSHt
sL6ZSibgH4SupXeU9GlbfRH3+qO+TUEQKBuWGSg7al6O2zTd931Oia1l+bmQ7fMqTsPc4XlwMabA
jNE5nMM4sTm3J1soiVUYwtSgal3ePstEewMd9Ozs/jABEKfHtWUxBurPKPR2Hnw08/PVIm9fqkCH
9U33XjC6YFZnxLWdUHaUdnoTnxHuxTDl+pMQrCaafFOVXWUzWHcEf7/sglKVzahxPG4ymQ7ro/Gl
nl8k5i+ljFbv0Khu+EIBJezI6IMbWGXywMq/ICp4+FdJBTKU77iySjYePb239cvvGCdU44fewDKm
3x3Bl+d236bg8zejHIoDT89jF7dnQraYjkOKHyPjjyFuczQBOIJHG+Vp4q+MIE1lFu1k/l0sJoCB
cg4g9qUIQyES6k1CuWCtSv5OFpU8xf9roSJxjZQ/mUpCnrxJRoWn9Fl+MhgcCxb24blrS5Sfde1I
HRlqGcKS8wYurlvDDqIM+A1LpZ2zwhOTaym4ZlwaYk6rQ0pqdN2qJR+8n8vCPEPE5Q4tyBvxx/vn
LJwN6FPQq9z5qL1zuJthzHnLPG4e6tA5fqeaCkHZvVDc7uNvXU/FnYQw/9bGkPG4OH8eKqPqJ0nt
ZeSWXykFUnQ0Dosq6Qp6pXJ8dHT6VFlsjoEmDxL7nEvLRNC5ushjvGgzLrV3ZK4sw9w8qYnkvHh2
fjFhrlkG+pljM6qeacTcjpJk/etGaY2Ls0wGZwA6RYB2BZ8fF5aNWh3Jrd+GHtc4VDHF0qjlbpUR
95kl/lGYr7eVXJsYkL/wgqs1reJUOc7LaZpiSWUjJh0D0yRtoKbopEuHvxvsr+piZFcFNvcGBC5j
6lzy4YTJIx8Rj4d1dJpjy63qiaNkL1CRF0Ovq689pi6yywU+qXH8HYRpRr46T0shg8a7xCKr9125
yUcWf2o7CdOEg016sDLT9OUE78AADxfPvvva0ysWFMbt+9jT8esyoCMUzPH+vjk5+0B0Mf5wbuCY
JcZi3HJlOJy5nLEWjcUe3NFdJ1s7C2OHEb6i4RWPKzZN4vp5UUslUjz+FXAGQMDFYmUzptyB/2du
J7984BSATj+NyE6TlGjXd4aQrTpI68i35Tl7ggA8tLXftVfEKNDjrnekU3cHuxVFYbXYiPuCJYLD
ZMkhId9buj7VJE8bD+pAR456Z6u0OAlnBw9rnSaQ+jrp9xX1jdDlTbMgHlQJCddw3lRCFEyTIPyQ
v+ne5ATcocuXzrc590DTSijI4MH8I/0znAsuRd1dmgbBTOsKHAZuao7wMLExLnsC6b34dst1bvjH
5j/u8q9Ifyys0TEms/0EyEXoHDSKrh8TWCVNnCfo7+D7ir6wJk4Okys8UM4oaRBVxCvTI/G5qvzk
bodyw5v+uev6SPd6WKbykfbzRmRHE/SZ8R6CChjC0lPb9fvEK1iXmHInHao1oIr1MD/SHpDEmMoU
HTyaRO0lm4KSZlCev1XBzfh03/CuTLFBsvvtYKrIHaZTZKm60zJdb6/xKv4KdyEaqsA0UUD9f782
1nlWffZuJx3ZaZkMV/Pc4E/TIAcEaYbnW/e3LEpCiW0Z4uHxIGdTIP0iR0eWd8H/b0uDW564YMdq
HMvd8Cc4EPP2Bh4Q6/SofKKQ8Ffc864pf9YVhYM1sDhULc58qS7fg0q0JyGG30wJGKgtj9jYDvxO
cOB4/iMhq1sRBLTl9LRJfjcoSdF4EUSUWupUn50ue4/QJT31FlUncAAUOgp89ULl6j9yVvK3thj/
J7F2Zs4vMeNDaWwRkWQI7HNzTVX8BbYv3jsqh0DSaiqe0L408tThJAyE0SFUwOS7HiLUor6GId67
hwV8Yvx9k+ZhQMIy/mQ/+0Sg6+M/7orMvXBCu/3p2sJqL/X601ITf+VRZ55H68KQMBWNOkjXm1Lx
aeQnBmAAgXvFrE61JsEFvNxOzoJnEEuDQCh1s7OHV6sOiK6LAa6JbvgDTy34K67WlNukP3dsIY0w
vByhkiF9Xwaa7yeLZ9ICtCeWaHYNtnRMZD1zQ9wNht91KxEIi8B7FLw3ODwObBMpzXSqyJymgl43
nciKy5GuwNGjL6N0qjQp8GDHS+r7AszrY7uH11DbebUNZk6C8uiIIxU4PFEcGfDuPqheRW8U7+40
vjOgk01Udqr3R/xh3A6bRtTkTCf9zcb9RTNfbmZQ9iDrZtNMaF6ELoa4O/7UdNu72Cf5qR3itbsX
0APvMeOr132hcwXesILNQ4NbmZ5/SsmRZtt9bsdRTMMp30MOs/fSzSUa7GtGPGJ5TSKsX1BGmRpd
jpkCo0Ck8DwAMW5tiVDG4KjZUJIDb75jG50ZxqzesWB92t22sbQzgQqWYsF76jBx/FOOJQuobnXj
TZQdyvdrK1wKjkg7DrTL3iMlIluWDzfHJWqgIrWwG8iS6gQu7dc5ROQLJJVT2ldeiZOHTbAXssFi
jbNo3ZcAsoYG7YhV700lKMExrXacf9uerr4J8xopM93yoeK89vo2LDRtpPctc1zmBvXKXjvhNAka
ldd3ikNKoHWgnnyDzHFEyRBIbpY5/Dmh1kH85pwReu3xZCDGtRJuFMRzMveIWHGaxqLe0A0Fv72L
rv2vfUh3G3K+DDW3NYE/Rmqc4TG0XmxdpZuynim7qM0FQ9IJ0OlK4/Jyeb4z/dqV0Huxh3Uvrpdb
YTw/OK7wQVMiiAJsjaZqDsgiQIV8xpaqCUBVJpOo/Ld/UGeRZOpaKk+OEKlEpjFqfFUPr5swJ8bo
NjC7/P/MEjAq31lRTAgVniQZYK1uSLtubbo9kJnLt287G07qxxwzxoUdEPUROdCtECXW6j23xqfa
YNd9jG0ZnS5PqOggw6Z5B3ogNJH19kjROCBXlZsejJng4ykVHo/lp1HOsuuX8c4gVK3GmcNcb36f
e27jOgyGXIqFOIQAZxJD+hKRWdxLyBtXdTb+FkZVCq+9PWZIrf2u6Za4Q4xpncM3Cv8J7atXRODA
aYwCU6IwzSaj0VGrQh2LtveV2wkwuCuVXwkbDG+LyJGOqFfxeweRRqXHRGFqHRzUwBVYdkLpkmO5
Pai7yLUvJiloeywMVs6wOI/KGXbdLz+dAUP7y3br03j1o6jUEwW+A7AzXolv+8PwcnCifGQ7zCTn
Gvol1UtfPWfXdryRMguejIsiLgA7OkqfIpB3oVwTNQOz5vIfLZ4ynBAwTr0WRgbs6yx2XtTASfBf
qiCjVCY8wzd0cLVL4Nqgw3Nz6YJA+SiBca1UGxoiXqVQTFlYTo1x4vV72uBdSuODOjxGrMZXZ1c/
H5XzGhCEmHKFXsGXyUBTqYXEEBM5heizEPJoWXHJdrKXxbTyTajWo7TeTZ6Dmd6uTA6RlnZXIBCg
NolaxHCghvNWljjlDEr17rmmgBZn43qiGiijbCPnTW23q9oap0H6/bk/IC12FBIa5kMMc8ychDeY
cCjJSMiJiFuzsefRNJXfBkAHDPlA+/FhdUM2l7grkdIn8+Qrorj3Aw/FShAj8Ek0K+OMcO8YFHIi
GB0D6qwpd8QSIOMYMQrjb5HDmGbc9cFMIrUUa7N1vqZPZTj1zz3pKf42YJTo3XBE5gJnlQAcfeC8
DkvS+Xwq6yyIuhf6n9JqKhs465tdzLksVWhjFeDbNTBioB4WKyaRGWBH3V06+14Dv3SOEaVAr5br
KsecWvDXXoTR1Y0tBwRWfKnVO4rcGRo7Nnsjqk6K6f8ZHAdBa8PzpLRjJB666QTDkyoRpeL6GKcW
mDZ6s24Geq2UonW3pGUuFirUtYl6okUva2zSudLHsxK4buAV/Qn4kuFE0bZh1SLwN/5lnX0a6CLq
UBwnimy3edwTCgC3uYM0BHkio9SLaevIOosnABZOEpp9WhowScChJCA9jCu2Q5e7R/3NxP/j1OcQ
XL/jOg3SOlU+NJIsMQVCQFNqcykePCAZd3/x1r5CA6ndKFEc6tyL3kGN6fOMe12eOpLy3emG15Cq
NlSKUXSA4nO1UC+YW/dPd19otYGflI/Y6EeYLpCV7hwwYQcHnMZJEUi8lBHzENLi4eqhsxIOc8JC
X7WByAIOuahcpMaFGw9HoiPMiRwCzo83NTacW/ESiKojlLCrpB5QHkU+gBuM5QqpBaN85lPf8RME
czoaCIvD1CAusxN69VEiVZLaKb+p8zWfwpXLau/UFBvFDbEeddVi7rBXmZEUgNQ0j78EhccdvdyG
V5nUUq2yNHJZiDtzHHDP4u7NX+TgccmAY6v4Uai+zQOYW6joy2S9QoELWqwaRlA2Edjh9NtYLWao
fyEAbm4l16jTzV2NvyULd7sWfMyWgtqUe7d5sYBh7UiyinItzqfRtYopMia9vaIgVb7/GNRT+bb8
DiQeAsgj3PXWAIEKGKIplz8kVLD3vXvN4agX0F7+whbyHnL9vzgash1CoT+iOXCay1fAtXt8k17I
kNWYFjRna86yw6tqBvw6DN7tgi6wN8OxKut8g+U3lTLINe7icGpm49uoCIe6O9KkRPhFGXNUmE7j
zRwTUEI4/eEdtFpxGQd8fGQXgeeklO1xI4r5XTxUmqxK2Z5pYn8Nhurs4npsHy8MqiiBqbl7i1jR
lh+nweAcw+WTY1ZMBFUuT28RV5SFfEu0hgn1QUpRf3KE2XIcMTcRQGTYAWshDo+oaTvwdIa50YPr
UJx1Del3SMEW61LeJHqUHmSGc8TkNJ5e3jAtKN+vw9wI1I0t6jhbLaBKn0ZX3hLGy3gUJjCwLlPC
aEn+r4R9hG7iuJ0L+Eh4YsriJMGpaVB5t6wO/AZfOTMIHka28MV+Ak2Dv8BrDkkniAuLTk/FzImA
j6na2+d9tOLjIgx62bordtWeCrKOGN6Wu1Fv3Exr/9xup9EkpVg2MJaFA0hxaSQio+7kpZcP7fd1
x/0/iNCX2Mku9VE8t4a9bsu0y8QxadU0SwjWRiJXEIREuikrXKOo6pKd3UNtYB1xmhvtaJJ732tI
dm5mLn5lw7LInnMILmV06WPTyKy74JWcmCSfzlurIvje//6SByuqufBFslctVHJS6AAVKRJe/5wY
Kz2AMVRlAEBnRAWFLSqkuPW5s1YH2zi+cNX6MMBiUzSe9FJb7qYAvi2mcUg5vY84MpFSMVQxWMQf
JokszVA60HuIB3S4mmiSAslR726badJbM2DYX6cMImS7xsKFxSk+rn77WL6pVYn5V5KoNMv/RXq5
04rnDz8hMf3PtVV9d2y5TRgEXbJb7wTPyvlcjzLE5lRHNCyRU4DdGKtw8uPjf5b+cwkYH3FNHZvn
ayLP6EH0DRyUFt8AfGEoOmYm3sP+t1U5TEM+iI7zMkQCvTyO1lfSXcZ3D1P6+469tdg2rbWixnvk
FmVJ73NfIBRwG5yEX7T2lKsIwtMkojcxCxnT3xkf6F2ghqcfSvGzmG5iy4eaI4hRpusEcKPqhgI+
uwAxWEEyKyW1f4O8bl5iOcMnFQIS6tZMjLPREl9Xb2S3mHpTVPpTj7kn/khkbHx6Iflduo0lKTFd
56aCdfxIZiWkjEhdYyQvqDag7S2T2vlLJWglW5CiZypti+bX7bS+S5bygvh1OR9RecUUMGRnsk/l
YNRRqVW1IJ1GfZUOBW2+e2mmp23JrqyuepZ6qE9KqBhus/8bGk4wPS/u2hZk7dHHCuj08E9hLpUZ
YTHGHZi1HgBk0ggQULm5zWfq9A+Eb/I0A+L2tI0nJhDUuTdXuK7/XQZJIc4579L0pGz9LxlTsTDO
BIDzO7lX0SQXPUafFDzFhjFeTh4AiCnKCRKhOmZE/g75xEH95kVQVnfTFWD0tI4MTR2/fSQsTtqo
2XmPHdYjxCFfB6coIyL0qzqEaJg4aL8ZaeYy3gMUWNtOVhkOe8MilI8dAasRMXL5qRSt2fIW7nPZ
8vHRTdulbUYaunB14VVsbLb725tOEY39Znq+3yXcyQTV9wh0euyZY04BNBirJAWmRzg381UrUViE
vgjRU4nOUrFRVkNLG84v4VGfLfrF11SIqRn6flev2He+eOAJ0M2MxRI2z6o0iJltPulaKqjjgr2g
Fq5kH3L05t4Y5Gn3QIWAsU99uW803lsExoEWr/kgQ5Apc1C81MQV+QIf80KwlSMkYv/DTM6BiE0J
tJCX0z61giqHWk5QF9Pl6qO5ocrZzTKxrch9jT3Iv+WILrKRSNkSIO9B7pmRZN0mspfDxRE/us5J
Yw+7zmQdHT2F/YDqCqWKlBiwGRtJqUmxUbnWKkH99CyCAUEDU8KBJGwKxObEemRIl0579aBdwhP1
/mbZuYstWdKEAf1Gp+CZOwqpckGvob6sp56W1ZSlscU9+KsK6C71Sm3ckNmBrG/sMaD/RII4dNey
WQebd92ldF4i5cMEoCBwBb4cchk5ozVwCEAqGi5QcbXzBn/MOhKnGFGok1TFuKyUChGbpwVEfcF4
rsZzPaJQgbum7rQLkyLiJreh6d9Pg4lpbqznq1PEdda9UpmRgCTLJPcVOd0jcNnB1i1mAw8AYhRL
ew61rsK/Ydz1b7+iGzOPeXZEAcOWabNs/IuBWb7uYQS4rW/bc+4Coke8E7+8C4lybZAEjbgVClds
udgWeLB/MeTfBLgx4nMXbCGJEjg2W6lnYfyWkZP2w9vmstDeatkTmhCcrv/h2oYgjqheipohVGkt
ad9QFX3bqKx1Co6HrvbbyKpv3JLEPRZm6BMmUi0TPkynxG8++FVyadWn6tKLD4hwrUyJsYRcqymI
X19WlfQ4hkiixmLkemjkokUiLdUgaVlEirmBMJ9nkOHOyaIqupUMvPPpRwb17H3aXiMJjwunuANA
ekttnrFx3uoQ92OaqVz5NLOlvPOFyTUFrtzalNKpuKATkL0fG5vTgu3R2N3cb2D1P6jNTVuoLWJn
UELLyf/lLhIBZgPdNYbUjcGmQmdAQ7XVJNfa4+L2AcGoZWy/HVwGJDEDByXyyx3Ai3mGbYCrIGqB
sD+8yUk49tYvgz5GlBcZDwh9x8vQFEQo2FPokq3ekM1zx82NVCPHckEiaxB+Zr6MXpYeXMUu3Eea
BxxDHf/Lj6W+oyHa95kTKPEoRWqV8Xb3riNNJUEsgANtcMwYfhdJkigbNih5RiQwnG0SEvPpbPc+
tTxdlmrEtkJJNnCzq+61AB+GqlEcNvYI5xl2HR9rLuIKcdNetBLxjhz/g2J1WCdcNYpOzo3NQdJ9
ykTXsdXFmSbnAXrCuEbBXK6jzqjmc8zU4d3iCCpIIgR03rU9umls8kW5XpjekDfqiDLGuHIbE25c
+vp/UIZ9ckn3EDCNlZ7GH7Q7FOH52LkI8PNX4DoDPBFXNswn4ntue6mrgCJaI7foLGJpYv8+WAsm
i13yrrOMJPNp/oxV90gzfTbvF5KUHee88ea5PI7hgkEJRQJE1UCiJl5E54sGA3ZU7ExIz8tbgqsB
K6GUGoyx16fNEdo/R4RmRBSbQl1MaL1dOepesjbfryncQecwg+V2ix5f9YzJYF2Sk2MJMU8gIQUg
c/IBgPOCFe75+WqW2FEXVk7afFT9Crl93HQGhjx9vlS2zSqbBUmd8NM1bGBPjylZZeH7x9mUJbem
kf6nTXSzYsmy1zEmrfqUet3Ps5pTrtI7lgKVPoMg6DLFBoLLTT5rrwTTE9Jwp5CGTH5Lo9706VLI
BwXZbvOUK2+TdD36eKsfDSO50zZC2+ZcLDfMZWea+kF4JDEF6eCXMjhK28DoQILff9sH6fhoAAJQ
uSsVyL4VKxMNLM4YvBbJJkOeIGTOM3vwbmGA0LCLd/IMUPlUta0moW+5bz6S+6QTEI7SaOuFkg0q
1ISrxIUPK7ELRCdaGRkBmME6YWLCwHOrGdNAsLb2vIQz4CKe4PgLNGskr64wnmP+Ywmov3rLuMLi
sHgidKb9MFvZDGInEWe/49rhE9i9PVzXtkjCEqNUkovK1JPnUSqyVUf0pzoiD7roxC6UrBIYjPM8
oooudY4fMNxCOdhgE/zpeGCQFUugw5b7iZ+qEsh6QCT3ZiZ9ZPl3w2OKCch+6q1HJxr9csbFJqWy
tpV/2t3SuOhDCudeegSg1pNrPRfXTyV9CB0GpLPPzBpHqkwbG4nLZnLJFMuWHg/94m3jOd4+KYoH
7mZR1rOIbnRns6Qv5pcjOX/USGXiPhaSY7AqCleDgk0dDDQt4Hglh4e2yx7p+KOc8VbbgqCaw4NK
Now1bivoplWiPdP2day3nlcdUNuYTtBMUX7HdQe6eP0r4XXub7JCTm73NU5FbUPlZngTxvykKvl1
lHWyWpWY8xFCSO61Fax1xJz4P6Cr535i4P9TKbLjW5FRJSJwSZZaoSOhpbLfK4Bb0lx3m8Kp7HHx
mgcM1q2jqweGFOicxTpaNE15RoV8vqZCLfY+xSduvEQYsNd0djNLBWDNudTKpmfEJaBj5sU2cp6E
TVVVQXwuCSOns3k6b9XOOvwWAQyj4tK7yGW/TtQmwccJYhFQdUiuw8QvUT38MO9ahS2dXolmcu3N
ZboacBwzXBzkcdGRaLJxHnnXyPo2chhVLzfxS1SJXAOYgdkXe6foey13POm22PMRybUzgJWDGEMr
2q+0p2Z0nmXWh1mlJSzes+sZKTKWVv1xEZs+vHnNO1NxdWmLn6ycFLfaeD6kby2iziW/JBptFH2d
luO3CMwcqJsmaSuiMVd1BNXrNRIAkjW2yrcntg3TyXRvf+5IR0U6kaoPmMSDiQxVIqGMjqIHoEZb
46sQZjVpU+UA4zkv1XGTK+33ty0/mlA7Gil73/vA6PU+uYyN7+mHfE6Huc7wFShiuIQCVvDAtFvK
cGkTYev7g6xNJFpdd3EK3Wt9vHs7w/p5
`protect end_protected
