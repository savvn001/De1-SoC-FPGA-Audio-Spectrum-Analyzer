��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	���)R"�A,ֈO�`�Fk�Q�D®��'�� {��5N��Yz�־�v("�>��g~��p�$#���$�/"�cl�eR��*&V[��窳	��B�g>�x
��>�峽��v�D����{]�Į�_>f��Ɇ�$Er9'L���T�ѐ��Q�T-����m����bf ���J��O�f��q��+�xeb+P��^|B���'��h�vՁ�n ]S��Ċm¾qm�̴{�lᥚ�����w �R�L�ܐ�P5I1	�p?�ݿ��\ `��d�^ɇ�Kt@'������d�"����
�0�)���;�����`�����I�7�+g(�I�C2Sj_Ɋ���>�c�caC?��U�,@�zn3+�/X�J�F꼔<D�sa��I�#0���,��&l�R�!̳��`���ͦ�3���G�I�����BJb�K"�?�&���?�w,������E�[o�_��0�&0D�v��ʽ_�H���6q�+�����E$Oߞ �����I}W������>�8���x�cUR�w)IF�3:߅Ԩ��T�Uj��d�k��xD�)x1�n�nL���4�ܬ(ta@%��$�5y��	�䋾 �1���G#R����<����6���i+Ԙg���V�yH�|J'������MC���+�[�0<\��bY��<[V��x�fr�}&��8�i諸��̸v�_����f�εS	ZX��tQ��<�|��:�^ �z%k�%��J�R�t[��H\���p���,Lƒ�����$����b2�tt��G���}�Q�S���nf�A�)jE�f�ƌ>8H��o��6E&�T˚#����Ba�ZT�E��<wOuSKh��a.�`�>�T^]���S���'����w������|�3>��J
-p��RK?G����;擬���%��f�5E>����Ɍ�J�nz���t�nJ`���!yx�A]g��]b���H`�h*�U�[^A�%����,V���Ö}�����@	[�I�2�[�'�qWc>���I���Q4�\j�3�Ex#����%z;�ْy�����ط�s��V��LW���^�+��f�-��c"@�P�ޡJ��z�.�,HM���2���ܱ;�)���NeRu�	L���C�٦+��ޠ�V�f��hh��i@k횫����Y�@�����9�p?K�yc�K��R7� �üո��p��~&Q2����_�UA��a�2[�k67Y]L�V�%-��`'��!9t!��J�17Wۖ�QH�qk&�P��]���n'��-Y|/�2���� ۊ���5'��:4O��܈4S������"�QӞ�b�ϐ�Ŕ�F�H���!)�m� e��ϭN������ǔ$�#���.�����U�km�?%�T|��R�K�`��7�&G��W���{[Ɵ8B�ԩ���߿q^��9�#)��f\����p�s��nڞ��L޵�G�@��R��S��=���/�
��� +7��,n�Կ�kdx��)vP���㭸.���3��ܠ�����hu� ~�ķt�����m���V�1\��u��<�� @�v֡)���S�4�+�Z����,��k.f�l'�7�����LC����&���E���._�����Y]\6nu^8R��	�Z�Uܻ�^"�hC��DB��=۹���xG�	@���*�흨��A39��<�3~&157D��ԙ�sjJ�i�Q�Q'̵<S�G2/)7����K���|K�[dW8��l1!��+�1�Q"f7�D��:����0�bj}�m"}%)J�n9:���^����)邪�*;����O�}W�:���
��)�L��5Xr��b,맯��ѥ���odOMf��X�����Oq�6��Y��	�B?���ː<�FT����^5@M�`p�b��D��1��Nq�I_d�yJ�����*'���i�:є���<]�;�?�_}�o�@�K��g�������ڳN���=�Y�f�L+��^ْ���ʹ8��tR�k�s;J.�J��p�t�cZ����L(�L������+\��]���1���&�GN����.�)�o%$�<�G��o!��9���A?�mf����5 �W[���6�B�lSu
�Q�O�����V��`Cp��a��W���f�g�35�M|��%X{4j��W���/>yEn��_+�`
r� ����"c���� ����wM�x8�$��P�'eL��/�;�r�>Cеt�Z҅����)Y�2�m&20�i��fNon��l�q���x��+�	��ŵ4kc�m��,4�(3���x�k	S�}���_�A���:�>%��0��#i��QuKsޓur��8�c�Nס�Np�|*��&��'�^bpp�V��!C'�a1in�,�VĨH���1�8?:,,^C`A�=B&Q@T�;���[��3����.[�/}'�kJ������}�됖�֬���,�s���c�S�ډ��~�Rn|��s]��ߧw�����8������Z~��P>��t3ʛ��R�����>�+��^�e�S�p]Mg����*\�.Vh����ĸ�B�,��;�|I;�A�K��/]�4�X�:c2��|�K��Dvb���h6 P��٨n��q�'�.Z�����R���f"����0��F�M������H���w>�2��v�`�7�&馤�K1'�G��M���;ǝ*+d�^"��{_*���{�䐝���6����v�U�-SE'd�7�|rwn�"�����1Năm�B_�sI���kv�<u��O|3�^A�E3!�&�gϱ��[�r���V�u��hN�TPѯ��T<cP�C�z�����@�Q������	�&�Z��m޺��'�ؗ0Ŗ�M�ߘs���2�/�����"���շ����	#�;1�ʹ��6&=�k��ų`|!�W�#����ʌ�!���M�h�����T1�`	�_��N���\u,Ͷ3��	B~rS7���S��"AE��]("�y�NP��i�ѳW:]�Vƌi�U��=H��$�o��	g�n��"��M^n<�Y�~��>Rzj���@X����,��U�-@����ȢY���w���覌ܔ���4���I���0<hv�'�������ƍfD���u�p����U:�X<�	!	M���0�9_V0�����|,��Dc>\6&�^���\��%F�R�8Wz�,7����j�RNA��_Ӡ49��Ͱ��� ��
�fƐxJ�=2{�P�L��@o�*)NQ����5�xM�e��7�p1;����F�����5�x`6�tq���l���w	M�Jy�b��?�s���E:����W�J���ufV�[@�tL� �^����|$���0�$��L임q�tt��L�zG,'*��,��������%ûǻ��Q|2�a����A��X��Mc@�!������V��#\i�����9Ѳ_�&���u� a2�7H�l�Y�]ʱ�A��x%�
�k!Q��@㆔���S��
�i���xI�͂{�}I� ю�2(�ᗔk�y��^��= ������"p�zظ���b	(�!a�"��}*���GJ�yɡ�0��-m�+3+!.܋�!U�}� �0�]� Z[%��k'Ubh���l0�%5_�^���
=�n�.�q)s�3��5K���PzXDW렭6�K��S�{d$sZ2$k\1粲z��>$g����?�O�]^���
��������8$����L�YʋMt��s��������7R���^5l�����I2a�_�B6L�+CɐM��k��&�F�D�&��_A=��U����M��(;^!v�F:�lݣj`/sa��������}�����lZ�ӏA��ϱڈ���?�h�b.��w��M�%����9 b�|��g$�EG����NP�I�G��m�3����%>Ɛ���Do�au�m5�;�G�/>1^�=�]��h���G���E����]un%{��D|�[Ԕ��آ���\���O���x��P��W����:��r@,�K�קf�t{�x+֠F�!�S�]]��q+;cū/��
V�����{Z����zl�"�L}�6��P�rTc打J�'�RxG$;�c�����k����"�I�g�Q\���g#�n)M�	��ϔI=疭+h��3�z�(4-N��!���uQ��R���-ZEP����5���)����@�!��g�L���zG�0��9�P��B)<�q��Vm��-��A�Z��;�)ǈ�2�$�3|��%�L�w$G(�	U"v�d�n� ����K��FP�K�񩲼-,�2[t��<��+#����f��d6a��M5�1[��e�R�nvP�k`,�]�p�ӽ�����9�<����� �K��S���5�.�TJ��Xf��͗ hM���+������	���LDel#4n?�g>z-���8������[��QMF&0����j>Fr�������Ja>���x��&Qx(�ի�^nS��^�5�x�.]��g}��RjC���x<���L\��|��e���+gJ������/���[�3�kx�UxW�l��>�0��r��d��a����~@]ѥ;�GΫN�{�ʄ��U�i+�D�@�bg��vZ��R�~2�Yǖ����8C�/���]��7D2�{���.�$'[�P2s1)U1ʾug'�7SJYL<�F��*�-��!!U�sX˴�4��~�1m�O�~GyC��@��oe�M�󋝝�ʒ-�h�+�=Y��o��
d���AF˪#W�"�����9X��=�aa<�M6�P!��D�1S��4�Q��M|AHv��2�Kk2���bN78���%OJ�ӭKSI�����)���^�G��{L�q�f�����9z0�h����v�5�&'�+��hB\��O �!M��B,Re�SE4�]�f��@�	�r+�[R��4��E�",�%L x�섮�YS�����b�Q�QX==f2�bX��;j��cG��mI3/楝9��ڮ���+��R��D�t~i�r�0�>ɋ��\����)������sJ:(,�g2�||���n�mn��� ^�HxL+�&�$��ȼD��A�wBB2/����w�%�hiJ B�1gr�����*�X<>M��:���P�v�v�e"�D�h����L���`B �\�