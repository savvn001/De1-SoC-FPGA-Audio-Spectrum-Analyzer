��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl8��M@�A�ZxzG��8��,ٯ�S�y��dTbR���9�w�M>&hvjvw�@���C/w��F1�Io�S�̈́D� ��e\cB<�����k�RzǪ>�׮��-�D}������dV�Mp���wrᔺ�~��.�klXRz�~`�@�ߚ��BK��E�p��ބd/Hxv�}!�-,�^#�N[�¾����N��Ә��o���.�S|kl�%̧L{�H�ESg髯2���>��(�C�p@=�;�qv�h�$���w/�`WT��69��
�(t�Enę+_���#�yV
���|x?ط\�6p�%[1�1Gh f㒫jcʁA��qFwKD��quB ���.���2�2ܷ&#u�������|�o��~�K���Z�������/q�:Ex#��r������'IQ��8>����}J�H�{���#�q6��leٛ�=�&K_����H���Z"����#D����$W�/��gV(]��g�U�����e;YcR6fb�h�X n�#��{�B�HӸ���@�0[�Y(Z�@~�4E��9R+��o:���:ȸ�H�9��ݫ�0�f�7��iR?C��o� ~r��Ç��d��.�ߠ�Ƞ=�췭���,���,i,�m� 4�duzR���}\A ��z�g5��Ғ����m	��N��~(�2�j�*��l���|���+s�]F�F;����Hu{�%��$>1M"_�J)\����Q��O[����7�~�	����������n���I��B�[��2���$��,q����v�/�:L��<�U�Z��a����`N&u8����?7Z�z��,Em�%E�E�ilo��y׆a'�����_�&��r��H��M�	0��啶�E .����_?3�*���Ư��6Jid�K��x�;�¡���<���L�u�̵(L$�!?�B���ˊ �e�'�z.�D�lPT$��������<�o2CHT\\�'C�Z��-��,i<C19S!�b�_kFx)��в��+0��/�bw��𜊂y����_��X���E
Ԓ���1���Ͻ�8U[����Mcw}���TH���K;�s2FB�FP,�e�3��CgB��S;B� ����L��E�,6�W�����\&��2/�Y*y��=2ƺV��(���{�����H��U�wx%sF�� �ML�9>�W�|HS/�����xB����Qkw�� �b^7�>S~7*M3B��y���G�*�O �_O%+i-�@!��4SL� `��:~~��@��K���8VBuj�T�z�V��v�Yz�Q�D���� ^����?,�P�>L�ߩE�z/�k�����u����6�����jyl'�/g���W�	�Ht�C�+�)�Юg��@}�vYa��i���JL����T{*�?=�^��c�1�w�&����t���1'�bB�˿�v�p2-��аt0��'&��>�C�*z{|��R�?bN<�߆���r(��ځ��wľ:�+�Z��%� [�4��G��`J��3>@
l��C��Y��ʄ�Z���S�J�<����!����t�ߒZ�J�e���ړ&�з}8��'Z�x�\�>㞕X��������(@�GE-W���aw�|1�3�٨a�b�=�hg�w}���4ʾ)�jq�M�PH��R��e@f,�ig�t��)���L��Dع�����@È
�]LC�	�:�BA�m��$&�ߩ�D*�W�d/9�Cl'��t��K��c�H�B�m_1����L�NuH�zU+�>U}#�|H��H�Q�w���/K�u�m�@-���#�I���Y�FL]
�ب�S|�iqY�����;������=�~suh��r�.���v��Y��5͝�{�����[���ͨ/h��dp��N+��߶.�_^����\-r��(���y`���B{+O��nΟʠ�k'Ŀ|�ɧR$.�ظ���oɘ�	�o�Nc<�0�#R��MR`-�nuO�-��Eg�#ޭ,��c���18zjؿV\%��iQ����Fi�oKh&K�R�������8��g�:�^�c�@���v������wx��RӮ{���w��X�������$���[J�hN�αOb�3oJ�J�GH*y���O�6kM6� 9�FХ �ѽ��ߨ*�G!����?�l�ʾ�i�M��m�B�2���T��o3`>�,��L�cL��g�����{B���y���T;�V>��~��[�7�c�K�0VSgu^͆���o�hasK\tX?��%h���hh�WGk-Q�Y!,4�2��9"2�^4Ҕ*E�~r�� �B�.�ᴻ�� M�B�zO�vf?�:�*�]��w��N^Z�� �oh�����%+��/%ܺͷĹ�_A�Ȭ���<��;�t�HF��6a����\&k�"cP5Y�̹�����s��~�ʚ�@(�^�vyT�V��pm���vYH���鮴�3���$^o�)x���<�� �I�~(� g"�?M�,%�����jA� 7��cR�����[�Q������.���zn�	u@�5���b$f���m��A2t
%�#���7AsF?����MfF��%�=�kx����`�7%��6A�49�>*ڭ�]�O?�H<�I>6�@#�H�`�H0U兗W���"J=���s z�J_���Gi�/)B=�C`�7�»֗��γ�8p�6������t�>`61��W��B�Y���*�aΒ� ]���r��.��0��;�h��;$����F��x�\΄�&&�����iL�Cr5�u�`�*����X�SY'�
�,	߻�l��DR��1�:gx��084B�k	���,�ؽ���/�*�^��[)=+���Ljj���?2L��;FO*���ɀ��,�&aQ-�X*q�]Ϩ�_|G�����ք�(��8���U�p�IB���y��R���*��1Y �Y ����k5���������F~�����eN���Z6i<I%,���@U-)ñ摊�B�����ދCl���f���=`_���W$c�b�5�#K��O�FJ��/��6�" �å�,b��J�[/B�l�����p���p�2���V~��s:H�=8Gv��P H�@2���@�h��VcH����k���"��`�=Hw�@a�ˆ�o�>6A+����TΤ���6�P&��K:d0�����`Sv�;�0]J�ܥ�N]BJ��Ҏ)z'�ۜ��p��!GwN���e�9�)Ț Ns�	zD#������ָ�l�y��B��8���X�$I������ji��
��"��}I��z\��%��3r��<��ӟ![A�&�A鳨f��s���J�\ V��
�V�Q!��l���ޞ��#���L����0�/�7����^�
o���f �j�ׯ���|��vsl�\f�M���4����Ʈ5���8k���9�����&�ty�lb�_�mdWh� �?4#?[ ��x�����3�.�V��љO�Y�X�ɴ�E�!J-�=O���4��P0��f�I��i��3W�ZV�}�ҩ��˶� ���5�T�ߝ�6�S��B	9�h���~'��LԎ���7�u�c~r��-ϥ��y���GQ+��u�"u鱃d�/U�h�W��`� (�*_��8�����s.�G!r@a�Lz���y�5u�<�N��].X��6�����ސc�ڔ?Q#��䦿�]��p!}9�w�2(*a�[��ISK�W/��t��riG�����O(���<��n%r	�~S`�%�qH�������Sh;�����n���#v;�`�	
T	�Sjy�d�f��Eu��J�D�Ƽ6�B ��挢�<�^���.�����z���f��h��4�����9?�<Ƒ�픨�h�u��|��n�U�o/����(jjrU���zGϫy'[wInu'��QNP�����
Z'����n_ ���<���c�FENNʶ�?�O$n�	'�5�{@�����J,�Qwk�¾S��"� %_��OC��\���.�3�m��E!�b6����!���G�2�l��{�\%���O���TOC��M����[D�
�gd��_�VW�W
�{��4?��4�����f��ۡS&<�*�ݚDP�?�өM;(⢯V�P����I�h�"��0�yB��E��0\�ب�+wa>�SCI�'2^Zl�]S���$�[������s�� ��?q��؀E�N^:y�I	�=Vn{���"w;�0h߬��'g
����+XȦ	�K�T��Z�$G�K���O�uH��W����� �.��@�˓°7���f�L��$5.l�*�tL���g��fO��L.��q�\0�)�fY��Тp�xa};z=��>� <SYy��_�Mi���#�el�`�� #�w�\A
,�^�"��a�'��������:��k޲��|�ꊭ�:l2����2���b���`�y�٩}��b�u������v�{��o9��M��� ���IA�m�B���d��H*/;�+t�葝ݶ��y�D���9IV`�����e��nK��ee��e0�lt�^�u$!Sk#Q�q�S5J���9��ㄸΏ{��tC�Ӕ�������Oԫ�M����@m�_2G���iM uc���̌7����ǩ�Iq�u���ȭ�=��)������M��eG�H����0�5���C_�v�
KN�kR�/�R9��qc��#t��Ůo��Fu?��+&���+Z����0���U��R�܍�z�����������=��hE���	�����沊H�ن���G:��*��k�ǝS�ڀ�75)X+���ta|��'b%Xkw�������T���U��⦎rg)⪰�r�!�$�r��4��*[�3����pW��[}ѬE���P��TMujrw��p�*iA�D�c� �P�M4:�;�������f�$F���D���q�����>��@T�ē��v�k�5��v��Ę�K�Sq�V
u�P{�Z�\ß&�t�4Ɓ���W�cF������_���~Zz�혿<M�İ���O�]���Ie�K�nF6p9�rfy�9��~)>�����乁F���}�wAl
����x���}�yR/^.�S8άw\���R+̓�}--9	z\�[Y�FS��aR��ԹM�{#|{��~9)3j�v���\O%��&*���t�I�����b�u�����TkXxI�}/ϛH	��YQ�VZf�H\���&���z��{%"ASI�0�v�*"
�>��b�-�D]����P>��SJ�С�q�	$��ɣ)�F��NE�D�$�b70����N�7��w��!�u�so�l�S���X�Z_f߉CW�;��U�,�CDn�Q�6���H˛��2��Z�T�Z�s�P�ړ�v��,&'�4i
��Q:��YG7*�GRqg�f9[�!Ա�p���[S��������p���B!_&�;��{��4�������H���D���$�w{ʂz4yf.��Rδ�'�n��Z?=�D��d� u���W�^Z��N�&ڹ�Z|���x݆*�@F��������nO��bE,�ms+���i���X�L^*��'��2�+^�s��{�����K�Y�U|�uʻ����05�?R:(���U�w塻�-���S|�ZI_�k��o��#Q}�7�-��F�UG��=�1�b��g���T��%W�G""����i��KY]������L�b�A捅]��d�}{wK{��5Ǉ�Kv�u�pG:2�����8����6Jg� �5�faa9�U��(!hJ�T�l���%�O³@=�\�2�fzY�q�P��N��;�FI�A���^�_�U���X�6/�\�&�&	�7�#��I͝�IW����]���V~Ή2N1���,d�
��B�_(��dU�H��Vh�B��r*�u�g��zY�W�T��G��ovn�]����gɓ�x�s
�Z;��_�������n���7�#�*�Р���}l)�̗�z�md�����.~�S��$��xE�FgT��q�U@U���F�]Gw���փts],�� �$L��o�zB�k���[��#��>(gwX,7!��.��f>h���)x�h�c��T}tvtZ��9����y�m�]w'�L�)]�+{��;i����G���]�лq?���Y��g���Kw��Ǉn�����<G	4�ܛ >S��In��w\w�����脣u��~��N����\e�A�q�~�x�M�qo7W�����Ɠ���ƶ�3aBX��(V�bFdPA�)��-W�~��Z���$L�Bٸ�y�]�:�r����T5g��>s�l8����#���a�<1��_�]�4mZ���&�O� d���=f��3w��:����(��o�Z�'���߹����ܸ ��9N7j쭘��愙.i8FC�$Ibϭv�P����@�ph�"�U�/m��j���4m����N�*��%f�'� �qKDYhW�aao�丯�>(�C/������GfǴ]��zA�$�Z㯶��=w�>��f�1����-�}K���(���Ӈ������<���jW�}��*���|���q� �{�j��+ob�]d��#��%3�|JC:3�P��	yX���8l�7|�.�.X��,&���1����߈c�q)Yf9c��]�gN���-��G(�R^`�txL����4�����O�P�`e�Z����=}���pF[���`���I^TI2?P�^!�3IB�(`J�6���q�쑭!p>��k����������ņ{��'������J��&��dQ6{�����2л�J���`ґ۬J�[E���űU�����}���k�h�q�9'��6ZL&Ē�o�������g�5I@Ei�\��ޏX�G:a]T*/���o�.QǴ2�����,zu�eQ�Ӵgfk2Ӂb\�yek���Z���8��W�$~�֎�J,*�`�mt7��r���q� t~CG��C<h���1�	0�L|5Q=ȧ��>��HV��i���Z�]r�cM��dZ���+��~���/6>�`�;'���2/�=�:��(�3�S�>���c�P$�c:L��v�՞������b�h	ֆg���8D�����-<�]��A�Rg8k�W�W5���_;Rop�����Y�g���/����:H