��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	߳vg�32��WL���|$�%�,~��Oq�GJ�JUI��1Q^/�f7��zܴ���*��d��j��D�5K"~�[%�U�^�ʫ����3D�p�}-��T����WS�w�#��ΎĄ��T�_�̳s�/�G۟=���m7^����z8?@B�H�GA���Ɉ���J5��Q-�XR��"t���?�=m�f�c�%�#E@fZ*a�_�\�����f��ڝ����.�Cdg{3�П�8�⁰ۅHq*wP+�spL�����LpO�ȉ̴B%�����O�+U���>��$h��t��(�X���$o裥L����*�Gxqs�ݴ��܊���ߵk�_9�o�2|A�����P2�ʈ���G3:�.y�(�=[[Gom'������]L��c>�1����4t��.@�2V/˖�.yc�Kd\*�
�2�ĒW�v�^���Ga�e9-L̝\B?�'P�Fw��F0S��n g�"�9�����F�D����կYHN�m�8)��s
�����AAf���"H��m����bE9Fg&�P�ĲR,�gQ�H�g�XjZB��������[`y���E�l��W�����z#��R��A�k;!#���=�3�:�q��cx���e�#���������}{-�hr�"�!����,� #ʮFMɳ��d�h��1;�iW %�\t99k=�t=1+e�r��9����F���!}I�E>?�'n�V�Jtxo�x��KH����.��]˻����[֎?�8]>�<�?�\�'��f�j(�f"��������T"~�TNm��㪤rB{�V;
���Y,,��P1t>%	�����$�|d�u��U5�pGO�asj��A�@� Ќ&k���ƹ��ɟ�d�	�e0�:�Əg���9M�X�&[����2UUF�[���n��S�{��(�J?S���se��7��b��M@�l�����A�t��h
���f;�T����w�[o �B�E�U# �m�ut���;�X��B�^�����՜~j0n��b�*��LE��p��̩�L��l�MӋx�;Ŭy���?��^��Qa���䳸cd̂	� ����C������a�=i�a����\O)n�.A�F�/���=��%�L���l�(K<���a�M��G���iO�&DX�l،�{lOW�6�;�\�BH��v��>/����U��LV���� ��ِ}�X_�ݍ;�d�����G>Pe<S9r�.�� ���E�C�h�7�H��{"橁WPs8�ˀV��W���~~W��#��Rr Msr��Q�0�Z�|�±�DmFd�7%�"u�����N�uGt�˚�,Gķ+,'�u����}_]?��b�U�wҷ�4XÀ�q�_� ����j����{�4��*`v�|��%R�"I8�j��1�zr�\m�
�b��1�u�-�;����W�L�Cɐ�����9B
Hw0��o����bv*H�C8�\\�W�,���*^�Kt�H2�C���.̛�qC��{�?a�oƹ�&�Y�|��8�oԥ��wPq��{��3%�)�������~�M����P�:�V�C���	J�Q͉KW~8�TQ�\p6�w���o�s�co
#���In���P��$7�G����u������N��A�V::�м�w�%e�ze��9���3]��_��jL'ѡ�$�y��7���m2"��c�>�4BK��p,���D�v~7!����B�T܇mN��cQ��0� ��3���:�¡S@�D,��pJ�&���]�>Ѹ����@��������9�D�M����k$��\M��Ь}F�z��y4���|���r��1���T��R�C|�����b2����ԃ��l��6���_�VC��2��7�ɾF������V�Wm�g�ƨ�!�3�B��z��0�kA)=��#'�3]�T$t��f���{~�hv;��&��X������+�ƶ�4�/�iQ!��_��ː��l:iC�s��I/u^y5L���3u��9������s��<�|����ds.
u	�m�
���2Q�\�9�I��U���kTsc. �o[�$~삷"vl�hY�iy�T���,Kk��X��D~�l(��z�(nM?��_�pyO�r���t%�WX��R���B���������k������+�1����8�h�w+ŅJ��)��,\_�3s��(�(��?q)�=�70V���P�FW�^�����<q���Kp'Љ��Qe�a�v.$�M�\$Ϳe�
R�%�ٚl����:C�H�^���%;7/ɍ�-�aȪS�lz�N��	����z�tn��oΛܛ�u�w=_
���um4+����O�"r����1������O�C󂿱H�zi�
jg�%ɔ�˲8��L��'}��B���v���:�)O=�h������4��U)��X�N��,��\�tq��o��`��X���b)�.-��h��z�����wW*�gkB+��Fڷ�-,g��˖~�Cn�;�뱊E�R��mql��9�<�g�g�:.���Ŋ�b@ծ55�@lҒK��V`S�� *Ss�͟���1�����_%V��j��P�w�C�g�k �d(�*��os�KGZi���N1��C#]e!�]6M� h04)2q���/7��;c7⳼�d�M�;k�(n�����	��a�cTM��b�/ �1R���V��K�4s��V+�&vI�gr��Sm��b�9�D�ꯑ�ǀ�	-"eXX���"l"dX���N�h�=��LgH9��rhBu��DS&��\V����[m��`V�!���s��u �� F�wU�\�gp
_��$x��5�Z�$AG�C[�wfDT{����S���
�1���2!=M�k㐬��d�z�����)�[U���y:�%r����S���tsȒ�1���k�nl�Ӟ�I��3�qIcC�Q��s
~�q�Z��\o�̅��h=|��3Z��1�͙�y���N� X1
&�,�Yl��̫�80Jto�>JlNO<�E�]١��݃�y�L�Ǽ*��G��EЕ��KH~���k��QZ�5Aѵ֚t��hm�R����ڍ
!�H"��c������B
�{ߋ�[��F����%Nc����7T����k����L��5��I�#�價˗i�%�����c� 6�/C��Ѯ�i��U����ԫ�������/Owyݭ^���l�*;鰫�\�]6�|��I%T��l�dd�c2B�� e�4�<&H�x���l�Wv�t�#)p⡏��V-�*��l$�_�N�(�.���/' ��B�vL�	ӯ��@ R���1�l)�2���-�fo�ļ�q�$���s8�|��`�Ɩ�JkT���s�9�c7fS�n���ys��,�Z�3m1�g�ܗ�r��$S�"�b��Rd�]�ť�u�Wg'��C�� 	���ZY�9�T�v*���^BȢ�����@73=�[4��o�|5*'���g6 Xl臶����Pq@�i��~��Cp�s���mA	�GQ��Ό11�Z�&5?y)d��IH�ͨF�g�Ka&�P�Ȍ��5d��#.���%�'�% 'dԖ�?�	�d7�4D��)$>�-�!�|r�tb3@X���(�k�:�v	g9�2Y��~t�1��w�xbힳt�e���4�=,��FY�p���u�v+~ޅ�T9�B���툉�\�ED�B���؁ũ������=ҙ������Qn�`�6�i����*Y�b��p �}��e�r N7\o�F�jp<j���O�=�K�5�N_��'�"!	����/���&;��߲qS|<��;-c@ß�ol#��ț���?/�}���³@�S̚˧�o 8�>���32^�j��M�T�V��?	u(��ߔ������Ա���
���9��C�ܗ3��+Pmۡ;/�w+�������r½:�k[*�bE��)r��k*h,X���>����>JX!i�J�X}�z<�p	K||]�ӂ~�B��>T��9���Oy�QF�%�R\2�`�������'�d5�آ�'{�n�2��˘@�_W_�^�ӥ��?�, �C�:�|����ԲG�W��K<~���&�_I;j�(�Sa�L�֓�S Ҧ^׵��V۟eo��*���q󵐓L�'K�P��Wɲn�Ar-�w�_A�S�=�`�t�n�&,���FnS�d�BX�Z����; ���'�����ە>�����Y�7<(�L���Uv�2�Ntt��(:���_b�y����0	��d>���J��3�A?'y�+���儆5~R�;4��a��4+pzSsJD�&�D@�<��x�*u���I��J�0>��$���oȃH��	!cK*,a&�Ƶ�cD�N_~�'����}���c���0;Ű�K����ul�s%����"�oSx�| {���x��ba@�y�M
��ԡ?"���6zK�&�	P��5��wh��f2A�\z��y�dP��T&�)������j��I�N�j\��K�� �%������������$<�7S|��<��5�f�&頶F�`�z<ӊ�
 :��6����m�������dŻ�<�.)	�U8�����Ã�k؉�":��-c�ԫ�r�w/�]����c��em�r�O��)�F^4AQ�{���cv�vd�����]�ղ�T[��s`q���@r���cjn��1�KM!"�`a�nw�E�-2	J�W����)���#�Zq�&�T|ɋ�s�}|tA�'���{X��q�t�"�׳y��R��k/:��Yp�ʰ���XO�Y��|y�[�*�T�	qB�I�@����::��{u"{��T��#տ+��:gK���k����1�6<OG}��w�sR�B6%�5�G�o��x�cS�8� ���T�)߿�v(�����Pg���ig�<� �����a�YO�~���Ȧy����h#jm������i�0�Y�����ш�RG�Y�%����a�+�Gƪ3��:y)~�A"�l�HB�Q�s�	�t�8�t</�U�	�5 q�����-��$҄�:j>T[�j�U���켻���k>�̓I���~�Τx4r��Ie2�$n�ld�9�[qyf�W�	-������
ڔ<W	��YxY������D���ߺW@���]�}B�V��
�R��K;Bqk0FV�$�`�Q������$zn�R\��S
/HL�e��,)a�Y������Y��Uh�V���Wl�,�a��1�ek�Bm0�!���n��u�I�-���6>
$v"��C�W���-BP�9a��B�FL�R��s�	�YzT`���� X�e]t_��:˅|�<l$0�{m)]N;� �t�>L�.h1AZ"��xl�j�2a�0 dǟ��M|3�M2��r	�uC��=��Y{�g�y��b�����[U��7b�D[)IR�ɵSH�[�9xۭ�fl�R�H�5�~吿]��N�y?��k�2� ��`��D��3�b\��LuW� ��P�G�t׸�c�IlsFJ�9�k����;u�Q9<�W"��HX�j�S��ř�9�3��-�\]�weH�v���@��l�j��"5�i�ฅ�r�Gz�fB�-^�dG4f��a�H���L���R/�=�E7r׫8����"�7�j@+�J�=g������XA~N���Ie@E�[Gp�՛�D�T��]"g.�DO
e�U��3U/���l%s��VC^���_^�؃к���Y��"�b�W\���p�=�Ij���<).]a+�1��g�t�e�A�WFa���*PS���`ScB�{k8���"��E}0����G�d�f�sK7�,�]�1OL���N6���1u���j�o`��IN^�-����l��Tmd+�p�I�C��=��߯�5���?r��!��h����#�x1A��X�!uBZ��݌j� �~��;bw��b������ �>�����?�_���ٞW��-Aρ�,�b�ڢ1����1`�-lC���_�`gz�'���K_$�o��Df��w�[8��3(Cc��Y��JfU#�i���1~� ���R@L#X4�U�h����T�
��~��2Ps]�x�6��e�B`O���;�h�b3td8~p�O�i�PĿ�I��B�t�>j&]�G@�X�:����`
&�N�E��R�.8:;�J���� qM��pIuY@�w�GT2u�Y�-r{�d&<f��~6xJ�R)��f���;g��5�Kݘ;��#�D�^K�-U2�݈;�&�
 ��ֺ�Gu8K -!�7�Xَ�jOS1�<��r�8Y~;ؼ-xU�wVΒ��Y�h0m��)��~qZ�����#1뻍��U-���Lq�*?�!X��Z�$|`�=�����G��e/b���q����C�&���3vA��O�
k�i�+rf*�X.�f�g�Aj�/ 	C�$
�]�{C:���������W3Z"�p��*��]�O�+��YZW�S�A�lZ��+Ӏ��?�5�	۱�;�Dc3'J��D�2��4�����^����@>O�W�8UƟ�0�R}9G"K��pC�S�E���WՏYY�Y)� �v�b�~�F�v�
�����d�[׽��(�O�t���y,��i���<�jv8{���Zxft?�p B}~H�Z� /Ǜf�ip\O���ϜQH"L���ƃ�=����K�"y:�"4p*�>�ڡ��/���@^UV�rTl���~j���])��p3Z	V�<)5vɊm��^p��ذ�%q�<�����0I����u�nt5��l�8>@�v������T�11!p��S;6�����5�-I��R{�j4� ��d�+eW��߿x8��`%�W�}� ��+z�	�>��U!/T��ܩ�yn�cq�>�<�{IB���)!OSi�]O��9CS�JB�9�t�����TՅZ��F����4���L��O\=(�7�OQC���r�~��S�~�85�bq�M:_�'u'c&�-��4ۮ\�ԯ-"	���.Z�u�w�P3N|G�lXR��/�墂�í����d9�X�Ӑ��ۣ�4�&�z�tX�U���O�P��y�"�!MX"��Q�����y��+�y�d�P�t��Tϵ����z�%M���b��1d �(�\h� ����WO�B����t��)�"����"}�=�
]J�E�����`���HDB�h�M����TU�.��j�D鰭vM[�S˲� � �Wi�U�ޜf监I�[�w��xgl���|�_{����D�etV��4v�2�S=��?CT̗�)\`䜋l��O�ܯ#�+ݳ1�|=\�T:���"�DɔMƢɺ�}oZYׁDpv?3�f��{���{8����׷���hꛟ(�uZo�9�'���0��N#�0�#�!\Q���Є�dm���A������i�����yN5�^�)�W���^���I�]e��X�H��$Z;f�C;����{�Qe)��Ķ����j�rʇ)���&^cTj1Q��޺��s�����W�`��|K��M�-��i��T�����t�{#�g�����0h�8��s��u��/��P�k�+y&&O%J`��$g��_���Q���p=�G�[IQ�媇�����'���Y.-$�*ڮG.�.��ME�^<�:�`�pA�nfh�iB��>��/!f:k�&
p� h��o����T����,�*�$���8�9{\��8�+�=�F�9��M���h����K��=#܍��~ݏ6���x�c��v�:�o��nj'���{p(�mn���~3gz��L|!T�>�����9h6�? ,|�l��c\��יi�Tr�����X�}��ϱ	gEcL��N	���dZ����R��e�k�b2�v;��