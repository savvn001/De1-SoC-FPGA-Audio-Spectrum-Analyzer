��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�~�O0���*1-n�89�������+�M��0���df�c��_ۤ ��LJ��������ss��הUk�����*]7j���U0�VX͊�����ֻ�Q�v:U2�����I��nm��h!zq7>��8�!H,��LV�`�������5H�:cb���w'#�~��S9"��ｭ�k�Ȱ�6��`�GM�I�����=��y�s�`����fGر̬"��Wַ��w5nܹ.y�`�>�� T�7�/]�Q��ڪW�s�XE����, *����m��]��o��u���Y/ �m�	���u��`��L�o�����Է��":��O��:���ס��<c��qs_dJ�Up,oq4�c�I��̬�� Qg���mCN�?����>Lϵ|%1�G��i�v�n��r���l�F��"K�lf]��}{�*7�Pv3�ł�2\&i*|g�(��pl�E �6f��$�Vޕ�%qۗa�`��*��MBOc|�E��$[�|N���Kb��R�̭uL�Jq�;�ռ����H�2�x�4>�㝣�u	�!�Į�A�b�� >�k��Y�� ���Wj���5�`��%0_ro�F���ǜ$�� �F{���$�>}�Y[�2ST���N$Sp�d�|�m{P��B!�wp?���+��������ހ��.�qp��8��s=.6�I�}��>�_]j��á�d�.5�:���	�6V��0��!�s+�;�f�pT�����-��o�������Чf'�����Ï|�y]�����g��=OZ���(fcx׿��3nWȪ�_�c1$PvL�
ż�&)��۟�eny
O)��e5F��W��[.���ډ%mc����{�AcDڗc��C�)���Yw���{��n�V�����G���<�r�?R2sM�j�+DF�"' s�p�^NB�§}��|�&��ɭ�q՘2��I�?#la�;[��oI�+}��0t��BN�c��-�
��k33��#b*m~�	��/�0Mr�Û��v3���[x�����Z,�
����=$L �{���Q�
�����qJ�8���j�Ę�%lɀ�X=VX/����f���f_d��~��'&�X�蒆��6"v��y���̞�+]2��e�ؤ!�,L����E��,J�kNa��6�g��j>���;����+�=(U�;jw\��&x��Р=!�Ō�:hPTFGL�>#�>ؑ�?��<|\�O�W����틔�`j
��OI��a��?�}��!���(��ׂZ=��dw����ld+�yG��m�@?ͫ�L1Q�NmV�oeQ�QO�������%��0a$4�"����f�3�
�t���7���6�D5�ǯ��^=���<S����]͠����"���tU_1
W�Ӣ���+2��yUY?�a5���j�kh��>0���rԂ���M�R.��_�@���<ֺ�������i�Vy�����duqd��A�5��� `�� K�8f5��z���%("�лM�*kes����!�Z�Q��g�Z���{	���yj'�9���#g�D+r�su:��c�C��q,*�3�y�R�a���S��R[�`e����&�~�T���ű�?���!ӞU�?*š��%��<���F����P�n`���T�O�@_">5_tw�F�a�L6!f�L!Y�9�Q<ϊQ6k@w�sw����R�"�<�E0�Y#�+ܬ`-�@�I�|��|�_M��W��b���s��Ɲ���1��K{��?����lfǴ ����JM_��l]�J3�=��{��Xr���b��v�jM]	l�7�l[��o�j̭P2�0�ܞж��;
�͍���
O�$Ҋ��Vc��U��.Wz��s������F�u��{4�~?�=���X�y�ӄ*�͒O��4;Ր�=���3��������Ʋ��YWlWN�2���e=1�6��M)y��bp������[�Q�3��*��ruplO�oK�P���с1���'z��ҵ�exV�u
��c3xO}�I�F3�,�}��e5����cr�$��@n�t��IΏ�),e���B�����F('��l�=e�p��半GWXq����3�''��Xُ�1�o��y⸣�u���0nv�fl������mh mѶ��o��OݝDa�����Cu�y13�iPK�:v�[�<Ș�F�-Ŧ�a >�l�K�?\i{�0����iW�g�//��+,S?�Z�nMbǗ/S�T�0�`��֗f�I	Cs;�cJ�<9ߗ���%��z�k�E��_�&��=C)qxR&�`��Z��J�l��eV:;i�`�q��ٯPP�!��$?0z4����y�l�N��'���Ҏ�	X���#�<�(���u^ރ��\hq�6������kE���|�£M���g��y`XQZ�(�>��]�t�ݲ��f�p�9Nws*KG�	��]�����)H��6w����/��;��S��3PSeM�����X~9qT� u	���"�책���q�I�z�����>��z�y��m�rKv�c/�������� 
:����d�P,4���(Z�Q�]X�D�q������	����s�JD���O����*�ҟ%!�(�<r�j�XC���b�.�@�_ݬ�p�*�(��Q��̪|��x�ǳf��T�X������ٿ�	$ҷK����L�6V��X���g Z�c��M���M���+�K7Gf�����H��O�?an�|���7�Ȗ+p��A�Ƒ&�L^Wt��3Ɓ�SMV��DP7��d[j�!���4���r&1�ɐ �"=�p�i�����v���ݕ��iӓ�ʣ,Y)n����)�"G�U�$�/��-T-q`Av�Fc<�,q���[�I*�������X�+����n��mMxQ����ḣ�P.�^ib�.�D�A��<�>���Nh~�(��n
�,뼌J�H����B�n}�(��Zܛ�� ���pǭ��}�lm�+[A�j�����g��`��F�*!��p�^���}��:�p��/v
�N�Ap�v�H-N8��Z�@t�.ג)��b����1����ݷ��H���|�S��4��Z��A<�#���b��ϊ?Z�,\��Jq�#s	i8����پ�!�7��m�?�o@��L�C�7�r,��PӦ�<N4근н���,m�zK7 ���T#^Cr�9�D쨱e���h�o�f^p+�&���J�Q��\zU�	�
�eTg|�
�ĳ�Y�ж {�2~䰰ô/���`zĳ@1�]���q�I���w5z�sk��@`#g(��#�>����w�wҭ���WG�#��}���z�7`��:�Fq`������`������
_�KkK`��2r�L�7¡P�B�^���I$�Sk�����Ӣ���`«U-�������;���
Qd�Q�$L�Q������{;\������eŹ9�2�� D��,@,n06"��-}`m�+漦����{E�=ש׌)(��W�n���}e}^���Z�6�	]a��|�g��;v����8�2c�g��z�=����f�{~��>�`��� {�A�u�-�y��]ݘ/���F�A��U?�Ì7�w�dq2$D��|��O /�=��j�^w�[d����ٲ�lD��x��Z�t!��PK��6=�p\�o��-W}��Z�9gx�S�������S$�&]�x73��q契�El�m�W'�t��ut3�|��m3^�m���gz̨紟<���;��а|��~f8Z� �g���	*�ZX�W�W�pY�Ȋ�2�ڤ՞��z]�M��iiBq���hj���O�����
V4� }�=��w�V�S��
�~+�S��s�om��g�:��h����2��\6É�Q���@i��&4".I��I���Z���F�������m6��\�+�Mh�{	@wB�x�Nx���h��H��=6�'�v�Q	���^��	�^e�e��ح5�U�?6�X��«i����	@If���2��2]W��� ��	�Z��ɑ�Ѿ_�h9<�6�i-^Rt.��A���`��_ʙE�M��T_9��Zɬ�jV^����8�^pE�*����d��0��w!�8yѣ��:@�+6�g}u�w>��rC��F�R�D�f��k̝�0j��^�)���El�e\G�$c:#���#��
d5E�e����%���!�,��R㻹��0�gW�$�Ћ/���q��P9P�\���᳨�f@��[�*=������ v��B7�Bn�<� 
��3'�\��I�ruNq�ǉ�}@�3�[�� ���vR�KMq��'�tZ�WY���.9^e�S����>hdFy�ͅ�������_�,:e){[��kt���~��AeiZ*�8�hU���]�iK����1A�tCW&�d��ǽ���zg��ȅ�3b�j#WԳRg2��s�}x���Q��D&�]K'v�B�LUP���-:����.G�?J#᠕ ���5�Zpo��3>���N)���Yq��O���@Ji���;��\��������G�u��#꡹�9��t��X4ВR'�	�E�H��%�!��ʦ�rj���TP��whG�k��aAы����ޱ"�P��H����~������WmY\��!+��D���x��# R�'�l�x#�hA���vd�uY�u�sj�X!��+�@ɇ
0��a"�оd�����zؤ��Ty�pI�A
-��e
����JZL��񳊈� Z��{n=}���6�>I�9}�S�Q߲�� ;�	 ��`;��Q�N���e�}W�+��Js/�h�M��G{���Z����{<�Dh�|��8�}!�Z}�@��v�]B�v)�K�
(Y4\l,j���d֥���5,02��:��+�1-��ݓċ������Wd90��#�և4�9��M�X4z�p���a�����:���q"���ڏ#WRZ�훫��m���b5��Q��QkH���(�[�(N��҃�O����a�{-�n�=�h���!�:�<՞�E��k���E�.D�e3؅�����P�z}'�gL��Rj�5��yM֥ �:�.��Y�`�Tle�ACl�^�������R�c�:-Ujpb^B��y�N��W������AE�!R�b!g�i�-��-��d`�����Cm'ǡ�����^+�G�&d=Z��MA��i6p���Ѩ�橏����e.�7?�� N��P�4�
��M$�[���D��i|�����.��̫�e�~�obΦ�}�� �����QS0))J��r�ӆQ����\�C�ĝ�ȝ�q�����SW�Zg�s� ����+��{l3��Ϯ.n�^��O�H*.�>���%KH�ak�{B���%f|�\�\�ڦc�V�!;�(�qf��9jZ�v~0�PK���(�<Te[��r?%n��X�"UH�b��oVl��m0hV� ��q�1��|.o2����
�r���J�OGR�E2W=�.�{����ic�oJu�ׇћ�c6����,�Z��E�{\O!g�8���v^[Ur�9DA�(;O^/?R����G7�J�ʼ�����X]72���Ӷ�F�ϛ2�0R��H�M���zıQ{�k����L9y٠=.
�)})�P%�-�t����H����	 d��t!&�q��ܽ_��V����������Q\���Yw�J�<�"BKC���8�1%e-�������������/���w�	���6e��V=4��TՀ� <���ǖ�U���%"ۀՑ�mC�	;V�L@��!#U�B|SM6Q�k_�|B<�D��O�U.oP`jT[�X�Ev2�[U;-N��]Xg���	�5\TJdۆp�7��.3�U��ã[p�
 �c�b�@G6Y�(��T1����߹ݞ�(Bo�Ȃ/6��,$ŕ=�}Ϲ �a�� �ĥb�ꪄ��8s��3�@����H��`ͤ�=���ɣ�>^�;T}��T��U�eI���_~邙A�en�SX��c��.���s,#?1�#UL�w_G�҇��i��ph?�����9xK��� �܆K��6��l�ߺ��SV0�|ot�b J��U�@��)V����;�a\���Z�� �'kj�����G�Gxy'�IE�]S�]�"m��6VF�UW�f��7��O��IM�5�h�j,��-�� �H���I6�i�RT8�EV�P����#[��~NH,�#�����S~�`
��T�~T+���_n�� �o���]�����]�'�����4A�zX����.Ӥ�W��9�W��3��V1�E$�o f�]nH;� �_��X!ʂa�$����+�a�
R;u3UwPU-=�ʣSŁ�B��3�t�������-���ԅ��#��GE/��S��ɾ�;����s�K��n��w�`������r�D����H�>C슖�fZ�sg�j�1w�H�Q�E�A���PҲT��ë�I�TRx%��e�W������R�!B�I2���;�u��V_�*�����y5L��Kg*���u��8��,#:�2����m�o�Rg�s/���C|�w��Y��*��˭���^ ���%���T���*�&�b���k;����.�F�H�6����f��#x�P�e<ON���
�����:-��Θ�����-����렌���1jq\zR���Ğ�B���a�k��Y��F�%!?� ��|�?��_\s"G����BƝ���d�Mv.�y</��ΕG��w��A�>���Ή\�&��$#����t4�v��=49 Ӟ���Y�Jtz��^ �.����;���ܑ����-�����9Ag���5F2ie��7f�$}�eB��3����,t�M-|�V����7�x��U<U�|�.
�v�(HL�2C�����_OBH��� �-��ܾdI�V������Ƕp�M.�sR���z�l�۞E�o�<�#G���|bF4G�7����PU�s�e�EL��%vk�f%���p;���Z�=JAN���G[��̒xO�p��N;�C��Se��}#
��F`��g�r�36l�UV���먳.�ũs���m�f������y�}�v���P֜\N�8�m�����[xL����@�ü�CSY$v<"��o�҆x	��1⁹A��P��q/v�bҨ��#�	:j�xF����rPx�c@f"�D{L�̨�n��|_�*����:�M&�kk�m5���|J�I����?A֍,g���H��U<Hg�93S��	~�gn�}z#������ q/,��KCͿ�\�h��P\��`;�p�
s���y�J�8�3v���H<�AtL?E��j@y{z�O5,�S�<�x�̝GN���X0V��o�D]bNr_E��P e������i�X��U'o(0�m/�����P��IK�����'�\]6��6t��M��C��̷m�d����Ў���4�.���+��g��+�Y ���/��Ch�P4�U�$�5\'�h6����
s���*�XS�d����ぁ�$y��H)zHY_�Q���z���{Vwˑ�q�ﮆ��~B�ts�����_��j����x^��<@�Ʋ��D@A��@AA�1�TO)*
�C�gA >�>�G�ɵ�����Qˈ�"w	i�%"j�� d��uR��Tm-,8�'B��>�i3 ���`���V<-�����>.f�S�s������+��3�M���f��3j���rl��H���'��g���g��N���'K�S����@�S[.�ؒ �3�J]���M��;�9jf���ᢵ��*�[P��dIA�|�Kb�J�S&��nn�4hQ��GN�:o$8g�h)�lm��B1έ����a�Pz����LCD8	�!p��P�1R��1�P�.�jM��X���s?�Xɦ�+F����/�Y`a��x�A��9�6F.�PN�� U���q�S�RhңI/�CQ�;v�����dr,���l(s�<�Lp`�=�!��hz	_`��[;q�&��R�k��&��0��5f��.��*��f�/��՞l�ۃ)-�i@v��.\i{������������z�i��d�����$6p���P��C�|��G pB�`(|q�F\o6T�7o��&�_�}.ϻl���j�g� R��}Z�����R��u(Էǀ���>�q�(~"J����3$��=�߹�#ʃ���&���1P��c������O����a��B�XbO큋$�i������P�����������@�g�s���ՙ������闺�u��� m�o#��K���,��!i�!��oE�����$nϹ��N�SnfBR�լ4*劅o&�ԹG���Oʷ���u�(%w���]e��Z�P@(7y��e��!I%w4�-<����/����ʰ�ԣ$��L�y��\��2{,�hY��E�{�߈����,�)P�j/P��� -j�
���_to/+Y�W�ת<0�fN���s7�ٴ	F1$��t�;�\���@�G��I���!M�u�RΈ5���T$���꜇�:�t�%�?����U�����M� ]>�i�m;�z�頾��-��<cU3z���ai ���O9���$3I ��Ƚ]ō�������و��+��et�Ĉ�~�ũ̷���
.��S.��z!`��)�^ ��J4��i��&�ǐ���j�@��.��r�+���a�VD�lAZm���|�U9�R"���L����7��ϓ$�ʀ3xL�����_�9���]�h�lA&�J�z��D�|�>��K��K����i�A�OE����]�l;����Gf������0������jw�$��l����P��nF��8�^��"���&��b�����ǅ�> V���͛}*lZ��Q������5_�3��!:�.y.f9u��w�@pX�Gs>#Z&$^��l�^���Ŝ�~�:�l���}E����g(N]��P/�7�.;�w�E�4�}�~�Rkdd��V9�84�����"�v���:/�i(��'�;;������vn1�~�4/�u�<�V��t�F����ύ��>X� ���֫5 �:���C�?4���� $�~0�:zL���(^eS��}d�X+� &֧���&t�E8�d��YwU��7eE2̍�Sz)1��Z�&Gy��&4<���݇�GN�*f��G��l7��F1,�X?�o����W�ӡ��x���(�=(77�߸X���P�e^A� ,�Zr��5$2�jx����x]����n��S���;���$�)�I�g~ >���60�z�0C��f'n�"%�/95�����xW�L,�_&�{;��j��z���t�
=۝�/�{��b�h����o8<��W��7)ĳ@z&P�ja���z��~� ��4�~���V��X3��ε�F���O�R�N���4���O�g<+�#��[��Q^�Q�9�;�il�H�L�u�0u���"� ~�%�Ph���r��W���X�c�3���ѓ���}�L�툎����B�?F���_�
�V�B�N�R�έ��l��#�x�S�2a�D��Bz�pe3/�O�4�W�$��M���V=ٛ�-��NR�-�f�4v~��fI&S;��&�������m��U ���C�� �ŋ��Qc�w���o��B+Z��	�3d��9�؆YQm����Vᓛ挦b�-M>��8/��O�p>�ː|Ȋ�]l��@�ON�\�q�ݳw�#	�$�Y��_~
KŨn�f;ɷ�Y��������6t4��g�8��ǚ��qA��V$@���ؔO��T�X<�6��G���#�v}���&B���Z�t��a�
4�۳ڄZ��(:�pe�u���2����OH�"��ͻ�8P���](���&=N�)�L�����{����	v0��ϡMU\;����t�{���#sQ˳��3�T�.�\@�A����=?���%�2���@��9ĉ��������	�J3�U���WP����ͱ9\U����3Z�u����+:��2�U�Q4Q�D��W�%6��}���$��H��G���ˎ,����"���]&���.!�/ �dK�$�U��zށ�Q�o�;ޮ��q�ga�+]/ŤucV�%6K�\ҺףH�0@8��նuC�����u �n��Xv����^��Q�M�f¤��	L�O� N�PJ9*�-{}|��*��8�2���c0��DK��F�w<�Kp�2��7H��sO�D�LIK��[}�_�\ܑ)�< ��=A���Q��Ѱ|� t��>p��"�4����:)\ �/�*_젾tR~qM^��J��]�hqAJس�Y��YK/@��,�2�st2�(��i���ۭ�Átim���zψQ�6�Z���Yp@,�;����QY�]i��`�ݚ_����ډ�#^�_XnҦBG�R�2�e��%6�JJPN+�\e2O�o��� #\�~n��ueҀ��v���
�]���}Ӟ���?9���m��<N�Pɸw���j����~����S�"��@T � [1���&�݅bӏ �9o8|!� ��(������Q�>(���hD��*=�����rYֳ�|��a��h�(t7S�2%���νx�D�K�n ��x���R��B4�i^-y�����/.�R�`ؐH�b��$�];
��$�����=�����>@�Wo��5�$,�!�GLI(�5�M��5 o@�f֠�(s=M^�p�wѝ�?�}���ve���.�/�B�p�0P���o�pځ����)����͋=X���Y��ݕfR0k0��[}?g%Gş�G?�\˳l��C�q�|�{�r=E�v��L������6�'�M��N�+*�QGb�;<J�C�s�h��ZCk�E�x��.`����kN_�9��g\�� ����g<��+l ����"�+�vgz�Ȕɗ �:VW*(��Vl��f��bW>)P��g瘊�+��6��t��%$"R�.��a��N i�f�+3��ۮu�wp����!��wd?i�&)k�JZ4�]1��.�Q�0d�����A��r��ՙ��s�P�1Ghie3Z�K�M����[c��}��tC�ckra��nNy��g?��=�?ŝ��#ⱷe�����m�E�+��M�����	,���}z�cqk�$8~oONe����l�z4��e/��`�d}1뺈��Ky�xfawķ��8/��	!��!ſ���LR6�! ��z�<��*�z�.����m������Y1�Qv��ݲ�nu�������eNE��6���f�%ǅJ����g��r���ֳ��_*zx�
gY�� ?�s��R��"��k�&�Cw	�����@?Z�M�g/����'�}`!��J�H;tel�Ϗ�:\�A���N���)��K5���li�~���T��7��	0�]q?D��g�r�T�w��z���L��� M,'����eց�$�	�S�a%EB�o�VAb�U2�"�^�jn�1!��5�f�ǲa
�,U��r���+l$�ע�}	|���X���%L���
E�'͹E������W�Ds��aU�~�1��n���k�[�W���n��{���8M���j���z̗�YZ>�s@�+�';�n��(�����N��*|`Ƕ���v7�C�ܯ���\gɜ�&��a�`�ՀBڷ{�>G�D��龭?�v/R�d]��M���h�Rξ�Ƿ!*�q�:���l|�.���걷u	�A܅�#�#g� �����\/N�����*�L�p�[�03�r%���WS��φ�k�ٸ%��7g(}������q#:��2�f*��t�<�N&�n�?'.]�M��(L3�	F���40�Z|n8T�<�oې�'#�`�j�:�S�W�
�,0ώ����;�Lj�8���1�c�{����$�%:(�W<wϼ[h�\�u����D�`z�E�t����Sob���D�`@x>��:�q���3�i�K]_x��9�-�٧���Z{�;���dF	��+�Js��B(�2QS��:α��І�#WK�&
Z����H�*��ɋӪ��:�]O4�+�G�`�>k���SS�d*\/�=�/"0q���C��v�� 4�F���J�f����ܠ%q_w�h�8v-���U��c-j�\�����~��x}���� |���|�"?�����.E�����d���;{$L�*�,i�ߴ�껂Q��6nɄ�����j�Vn���τ���D��Z�����S���#�\��*e�^��~Ф��ܙ�z�㕘m��.S���Δt��J���n��	�f_&��Y�=�'3����WW4-���?�Y��momL��-��`�l��p8���!r��|�և%H"$�������i�JiV&����V��|g���;��7j��ѻ!������/h��r���g1;|W�¼�ܑ}�1��ܝ;D���K�s���93ȏ˷��LZ��"�E�ڂI�|��DL���d���z��ք�	�t��.��1�>(�mi���"��[�F�ٷ��$����M�gL=aԨxn�߰t�kX�[��&�(���I�בy�� f+��$�GN�JO�"t�|��<����90���0x}�Z]K��!x
i�P��af��i��p�6>��-��}n�����ّ5�Bfv��ޖ�4"�`�6�2�+0{��>J_s�a����G�k0�[ݞ�ߡ s��Apt	ж��K��["}V���Q��#�#�٩ D�<�s���0��d՛T��ӕ�Z]�߆'���8�߸^��	�������)�M*��O�O�=#U��]U�tp& ��e˫;D���Tטg1~:����_C�,D�Vg��PoK%(�6�}�LG���7����!PLw�|?D�Ά*������{*��,�{}ԋ�<ܵ�tȧ���k��&7C���1M�L����^����;B2�4�Ù��6��S�o��(+�P�C ��i�?�k q��݆��p`5�A�_-��}���R�<(K�'�l��t�������`�67������ԯȬ�¢{�H;��8�9b*sr�|\&FRe$
��e
�PPJ�B�q]r�E+'~�j�nқ�����^�IX�k^'��N�y*�/$�nd5�>���}���9�L��Ɓ@B���1�D��]Ԗ�!��]�ӛ~��gg>;6|Aâ���I�:�7*i���Lʵ)�l��{T@B�-���<#�x��)��b��,	��������p��ۊ����S���:s�W�X(0���赃�܏���
>dW[�f^g�0]�B�@Z8�,��pZ[��W��d��,򵦴� 5?C.�`�uo���Mzc���#�A��+1T}�<�9˻4�D򤪓�Y�QOcsى��џ�N(o�<�{^��d_,�;�U2g.D�[E��q��@�r����c�-)͞�gO���"��ho�@예�:�}�D��Y�"�CY0F�K*�/q�a9B����r��-G��5��ݫ��<����k�2Q�����C�44Q�g�;�1%��Փ��?Ȯ�ւ�5˥�eusu)k{O��ls��/1�����]��ש����0ѓ'�C��I7eAM!���.����c�: �Ut�c}۟,�k���q�M���3[-��ׁ���w�A�}�1��q�?Ӟ�PNV�=:m0��Y�~�N���v���Q��^��q��]�99d������{Yݷ�n�A��Z�ä�:s�?���z�y7F���g�#�)����V���W+DTP��,�L��%z�#Qz0��u!�)T�4њ��ә)~Te°qrN�Mne��k��"T,�����-�n�v�9.kO)}�7�&��'��(0پ]bx�BͺR�4 [�x[?I�E��@�怶�rÏօ$7E�?5��X�U�cZ���ԓ�? ）7����dS��%�g��o�t7�Zy�hQ�WJ��y*+�c�|�ܵ�n�Kǽ�+����2D�T�-}�-6H=�}H�	=K�M��������+T	��X���ݕ��S�1$1��~ ��N^�t�\��A��5?(t��{��ph�,`	�3[ݵ��C�ĳ��Y�Q"�3'����w�L:�ǃoӨg������8�#�l�a�^@NRc�ŵ�Z��zQxk��yay���$Xy���2q�]�O�z��F��Qo��)���t��8�m�����E�Y�ۏ�y_}Ra����Ct���8y��ˍ���@����[��h������U�H��҃!��7jg��V�ov�ؐ�jwJi��$1����P]����&�����I���mE��T��8��V��=W�g�F�v�1�Vrs[k�L�o4d��ֹ��%�����dח��/wrD'AxP��`ߙ�V��ʨG��ŷĬ���aW2n�K�q� ������+880�#lX�>�O�y*^���BtXQU�n�e�j(�ǎ��=r7�m}K�3�#��.��*�:�t$'0�"��&�W[1�Tt���ggwuHŦ8aǢL!�C�}|���`�N�FZ��j�W���:�1 ����v�/\~���U�<{4�#yBv�Ӥ>@p~�F���k�ag��QYs��s�1n]�M��_�!�,?@:J-"$Ԧ<��2�\R]��+�z�J��jҡD����V;-Hcp5V�ν+�Z\�s�* ��,?��F�k+���/^�>�����:#��&�T�3P�9)N݊�l��t�� k�?����0{:b�&!�+��*v3���B�d%"_�3�[|�*�����4;	��TE��k �(M�����BR���)�R�A�_���|=�ڎ��k$EPQ(D8���4�Aϯ�Z�뇴�{TV"��7S"'�5��t,�};G�(������9r���er�M��kW�Xk2V� �5T*M��$M�2	6���f';��y˳5�UV�/U��S��T��n�BN���WB��wGd�nX�+�X�}Ʀ�67(�9���n�`t`��=����7@S0y �QR ݘ���0��}(%����d�ζ��c^De�ΐQ���j*Ԍh=h� Kbܷ�.�j��EBMy@a���ِ�lᬈE�a��� ���Dl�y�I�nv+�����h��Q��F�2Ȧ��j�|�e�!����V���yr�[�n��4ݝ[���xR��ݚ��+��5�� �5n5�?5���z�#���AޏW�qw��)�mq�ʕ/�&�ji"=iy�Y��Ɂqܯ>ҧ�����]N�8���&�F��P��L�Vl�4=��6Lf�#���yT���x՞�p
d���`%M��$`m��Ɗ)M� ������<�'�o�M M���69���G��M�*ļ�)A�c:7�j��Gbf�)�W@F�6vA�:���ŒT
�%��ל�>�
�,��P�!!kW�F�g.9���	���9p�|>�e �B�D\?���W��_�D�� ����
��Ҽ� d�;}XV3��j�@x���HsR��/��~�$��5�����T�Nd���5�J&��WB��j>�E�Ϯ�G5�wƵ%A=츸���<)
�}�SJV7L�ݔ�:	7jm�\1{N�;�+�F�
[��&�"�I�"�Q�B���c����<��%[׹%kb�-��$�7�܄!�3�z�kw����Ԟ� �B�ms��
��<��Ƞ����&���*�aI�A_�r��O�b|�y!r<���V�}}���Է!�5�D��q>#��MԄ@y�|6<t�9D�]���>��h��;�Ә�'�+�$��
�D�Z���1�ߕ!�hT������$�0f�rAk�b7��+��~'uIZf^� ���y���q��B��X���G�� �D����|-Z�SV9n׃�h�f��%Z��Pf$�z�Qe�P]�md��o�D[��od���C�`�d.>�&�Ed���b��F/�b�t���1OgtY!�{�kf�d7tL�izDe�5�9�/�|*?H&�C]B���c���LjY�19#I��f�/퉞Meo�����u�K,[r���x=��M6=6��hH���A/�;�FG�򦳢b���j�֗�Rkf����8q�h��=M� z��;�x�K�!"v��Ws=KR�̊T�k��LX�#��Mľ:����3�pp����uT5`p�5�|��E4���/��b)D�?V��p\
�񖊁��m.fB}Ĩ2�Bo�	�_a���l�`�b�S9���,�z����P�������]�f4`2\�_�k�=K�nQ� Sw�1U,�*�Dv[��1J���2q�!�9���h��F霼�����(4�_pR.0
��,�F��
O�m>Zщ���0�Ǌ	�?x~��d�m���ݞ@d�m o3x������{n�t�c���ౚ��01&$�*��nl��C�=�>��C&�o��5�<���g��$I���j��^~��*m�J�)_���$�'�k�B�u�2rm|N���٘���pI�e`v���6�f��1M����$�����ܣ���@����4��E��7��f���ixHF�Z��O{��m�M�*��h�S?�ڈy�Z�Υ3�L9̒9(�#�,�g" �f	ApA��-��l��]�?�s�	���p�������4n�Y��$�p�g ׏U�ZBG�{BY|^l��~�3@�G?~���!̄���S�ɗX��R�ϣ�����q���jw{�������q��`��b/�dxm���V�c�i=D�a'��� �e��wPp�2�b��wf�~�	?d
-��*lpP
<�"O�&��|Yd6�K@� m���T�+�JR�M21�x駬���:���!0EK-�}p�����Z��S�-�iT��(Do�{���-�]|�����1��T~P�N_3�j�^7v��w�x\�$�߶�Z2���O�_��4��'<����b|�P��b]�S\�փ���ߞ;�i�'n��^��k�!���?�{�q�����U��9��c:v}%���{ja�I�F�'c�}��o��Q��1���2N�+�B�0?P�yT�L�I�;�Tl��yZ:;�>/��F���9��H��B�.M���Ug�e��e�LB�d���{Bөm��rVR���w�{8��/�w�#Nf�(��˙$0_��{6
Mr��>H�V"�|]��!�5�j��r�F�F���\�~�ic���t`�7{"�n�����c?>�]�l��i�[����!��2����O���O汯�~l��s|0Bg�2SkԵ��kiʀf��~���R��x�լ74y����&>e#��k�b��O�&[�4;�7�'V)L�,���ΠDBESm�^I��kj�-n�3�!:Σ19�~>�s�k�I�3YQ{R_��~�`��""&��6�8P=U����🈔��or��V9?esgR�y�բ3
�� r�{�p�{�.I-Q�ݨ5e�D�&7�"&�"#,�N�b`f���� �T����xw��=N`
�(�==C��x+�Gk�iq���p�H�n�ݤt%,`�U羚�4\RGrg(QkY��-"�ס�{Q��	�`�#���N*��%����d}�m��_p�T�Nۿ���_�fdKꁒ��P�o@��q��T��ge�L&��zL�ov�|� h<���/lvLAt�}��'�s-Y�%$p��١ep�/�&PJ�Xމ0�|��H۟a`PX����}��LU^l�ݗ�6Q�d̤Լ'�+0MJ\bT|�I-��>&��W�P ;b�d\�$(���������\��Z27��*0d�!D���t�K���R���]��L��;����lr�YE�1kN;�L�����0_	0��b����� ���H��rG^Q=9���� �Ah�9�N�-�x縮��u��Zd��N�@�fM5A8��+�M��Y��/2a�I6�����Б�bѮ �]��L��$g�Hr�0�X�)A�c[��O��g�&S��_��fd_Q�B\tr�,�7�n� k9.��$���s%����q����d  ���W�OR���O�V�}�}/E����(�zռ�i���:M�S�N�]BVL�7&�So_�n�Q�C����O8aAg��ëO&2�j��50����I��qSfgDW�>X����f��`�[�9ϘG�C)���5��U�W�1:�A�)�r^&���F��Õu��dy�.ZEl�:BBE`��=��xL�7?u'HA^�����'���T�S�6�����Z�4�(l ��h;FpҐ!a����5{�v��a��fjx���=�	�tF�h�q^�~�d	]m��p� {a�uv����@�oƎzZ� @˄���
�W>#*�Y��a�Ta&	��}�@)���vI�ʰ�7�qȲ����dN,5�a�C豅t:�^�g�K�R볅M�9i�\M�Q����V"/����0%ڽSD��c�P�5vu���(�	��M��Wam�p�齄M�:�k�����L�����m�I6���߷�UTIm�Xf�Q�U��o0:S�n#<��<�-GY?��9��/+$`�#}T,o�	��<ֳ_yVw{�W	��
��~�$��:���)U��ܜiNG� ٘tm$�z|_Q���tD.$����r�f�q+\�L9	�蟂�F�BÁ]��	�re�W��2��
����kT-�p������J����>��U0��S����$P6�j`�:�KuWV*���+M(?{V�>)� �߾�!�}J��3�o�ld~�����A..k�%�P]�2. &���@_V�f�� S3�dj|!��J���a�ͤYm
�X"d]�߸R����c��E���� CUk�3=N��ෑ�
?x����Hv5k*:��\5�*�S>d��UlH�<kr=B��������^����Y�@�.�dr��
 �M�1��aGJxVe�|
�&+�²���x�����oX�4� �{f).���?op;85e��9���v�D<��;��Q ns�[�sY��:����:�����!�hwr����ؙ�|>�0��k�(��/Ս�!�I� k�N�S�R@{��G)85��\�a*����9�oƬ��6��E��J�#�Z��Q��YA�%��u5�^���f�p���~��a��V)cVX?ݪ����϶{	�3d#��="�!&�dPz�g��8���c��{���0x�b��I�Jb�9���u��� ۿ	Y8����ʲUDɉ!�`{w���H��nU+��WS��L�
��Ǎ�kY ��e5��S�V����ɮ�"����6�����|�s>^HDp"�ޡ�4	�o��O16�a�剄��Rt��4����^W��m�J�k��I^��4K3x��m�0��4�6Q����E��6|��Sy5���2/��y�!/�Y��p��>�Uaw�D��4��@%�K�Ҁ����	������u����K�]v����p?a�:�G����#ik��*|{�{����c��E��;HS:x@�����Tn�?¦�׶G�e�?�s���Z����4;�Qq&�,�<)��7�#��V1�9|�(�q!(je�'��@u-�����uM�Lucս+������)��g�W6g���J��"j�B��-�Q��3q�|�oz���1�J3]i/)��/�Q
��9���d;��[�{r�n6 �c粄������%�V��{�,�q�1~}����I���d�ԥ�;ty�l*�x��_(���O�4�\���Z�anי%L������ؒꛛ�}'�n{����G�.�7B��`���
e8����d���	9�$;ϴ����r�F���Z�@9�k)N>�K֜�`Ѕ�"���U=�-�b^�y�]E���컓�,CzqF�:@m��թ�(�k���ڹІ4�����C��w�?,���/�b�^�N�	�,zX�b浕�ZZ}��IYpŞ�S�)*H�q�5ٍ��(:@��0H>Y���0*uT�Vd�|���^H�.��@�uY8�b9���ܿp�hMQ�۲�TW#��U��NLXgpX���l�!yǘ��ȃ'+��b����0E�\��q�N1@�b���|�&�^W3?�I@I���uAIj6j���T�YX�[j��m�Tꦍ��}^l�Ov�-S=�U$㎟�]_{�`�g�ի;��	] t�Gj���σ,_s�=%F��
��k�.�֒��#h�}�AO3�"MtФ:��X�"��CDƷ{X��f��YOx&k�e)�	�߷p_� q"�tZ�i4v*�YnsaM�Nd7P1��6(�B�}9VU�E}�Tɠx�8��J�������?�d��g��}�j�ߎ�%�=p�4k�L�X��6C�j��u}B+�QȽ��9M-W�B��Mi����Wx��
^FeU�6w�R$�m��Xn�_AP4��9��x�
�m��� )Q�a���D�,�����}�Af��x�U˦9��z/Cc�m9 s{.�
�BA&�$B]�n wnS"�*���lw�#B�8ƈ�,��Z}Ǜ�P�,4#0�@���BQ`u%�E���24\H	��HV%��S^1x~�*T

�y��
��6��%�\<1��x�}��X �v��b�{�F3C���]Ȟ�P������������'�����*�O�Ѫl���c�L�PRy����P:Ur���s(9������6-ٴ�����r��So�;(���?���%j�����V��߀W �N UH��Ú�{	�#���Dr�|u��l���U���������9��J!� � 2^������i�Iu�)�_S�����{�yOUK>h-W$�o�	j�Rwݲ`��cqX�5��� �
ǽ��.${�5�v^.T�$ډfɵ+:?�φR�w���?�aU��\̋G�n�� �����(�f�K/�c^��f7��$aT�J0�[9>�*R�h�)`E��M��,����˅40ڥ�d��W�U(I\�~J	TIK�8��&�_����,S���o��G͕��ȿ�T�]1$o&UՍ��e��*6Y-�M��j�4�D� ������{��U����������5�Z���7X,D_c�B�j�k�� z8�����Nh�P�������`�eC�=�B����!��M<Z�H-n8� f]{���ԝ>�N�]#�7�ژh)�:-;|:����8`e�����ѝ4[����E:܄.{
i���R>-n��6R�M��j��TS�V�#���	A�F�?}��zgz��7��[�r|!;k��6�ػ�P�c�i��5��བྷ@p
d���_D<�z�T(�X����H�Ě���
�@��%�����)Vz��?��>W͵-��z�(��C�w�UEL͖�bF�tX؆�
��U�'"�/� wkw��х�H��>����&I$,�g�����K*�(�b~��7#����L\�G�E���SdN����v2�{uZ��tW��{q��k�>ȉK�dНZh��r%6����/�:o��� l]3�JG�h鯢/�	�A�g(��G�#�u�A���1����M\�G��jl�p���d����C�l**agY����l���.ƹ(�*+{i���ܰ|���/�T�p��S-~�.���-�j�����>!J\h��,G�dd�:��٩?4[��b�\娄|�z^��{�Jq�����,��n�ւK˯�LF	ĸcB��sW���[����`�<m�T��ԓK*yz�����1HkH���v��|"�z�9�+����1��Ĉ����Ƕ�����c5�<T�T�¬������Y����:m~	�G@@P���rL4h�˳@6��hm�5#�ژ��@��G���~Ml�%�R��Z^m�	r�macgT D8j�����\�^��Z�ӣY4:�%]���9� �U���"X�W��\�~��@�-�Dm�B��2�f��Hr>;q��,�O	2g��;g�%��(�)�J��	�j��Sa�Q�G�t�w��8O����0Y��LUEF'�wI��1Ï �,a(ˢ{�����.�M�S��3�S'4����K_f�mݟ~ʦ�,��l����j���b��4�&���g��l	/�7�x��23�aw|���)�Ĝ�RÀO��B��D��3��5��B{����?�4>�$!E�M�j(�-6�S����T�K����>���~ݹ��1�e������)�̘< �}O\j�3H�βD�^�h�:'4E(����T��.z����&���[�&%w�Z�G�A�ɼ�F���<߹ʕ�+A_<iOnx'K�$���"�$rO�����ۍ!�-h��8c]��^��m�|n�/���Kh���V\����.S I*��J(�1`��-�PH#7�	O֠I�m���k}6�T��/a��,𥉉2K�9��w�=l�:ǔ����?���9S�±u�$��UD�d3wxl}.��y�O�Y-ET4������z�^y��>7t3�1��h߂.2�j;����TkȟL������(T#I~"C�|Q�mV�;�K޻-{�k��3�KI
l��xU��YB�j�g$��!!���g��^k�m�B<s��4<��$��@�mI�w�� �H<�7QA�-���� Eb�Eb�䡟�R��`�j-Ɣ=�P���"�uo��UB��7N��O����pS�۹Y\Q�xF?L�It�3eN��&�����w���*��\F$��(��D��Ϭ��n�[�}�ު	�W���w�[ ��A3Z���'}pP�)G��S�o���@�jz����2^�*�Xe<AH�,�8�ެ�9;����$�+M�3�}�\�����!�0��v����X�/_�z���0!�YQ7:n^"��%@��s�b�v)���(ك���٪�A�n���o���f-�oB���3(0�7.���B�Y�����MoA���g�}��0�*��}�.4���=Fx��{>��������!?�	�R.��b���2��V�
;�'��cj��8%{�W����L2�a�γM�m�@�xG$Y���k��F�#8&b�<"��u"SD�F.\�Js�e��,��m�_��fa���n�Wl�\R~qaK�W��4�ϻ��m�T�D�/��`��\ �����W?����ZH�9�,w������ԧ�2|¶⋰k`��t�Y�T����y�ֆ�磑6���ԥ�Z�QϏ���I�8�7���ޛ�`-@�K��M��
1���]}��s
kBp�c���'α{v�7�I�U����Ci?��J��.u�ۻ���5O~8��&w��|v,�t��b���C"䢳����$�����љ��h�ʮ]ؐ,D)�6,�4�[�N��s��%���
;x?���GEE�1��Og$<@��~��F)�\��|�о/n����^{�,�!�s��4�~�e=&�h���)M�/$��LL��
�cx`O�2l��a��]T�U.�QB5��o���=��o����(y��
?�x�mvm�{O[�3t�W��B)=pR�-�4B�%>'!�u��g��>UF���x�g=gU<�/1W��r�M�,n�@G���ѱ��k��`�/%*@��q� K�(���sS�t+�Ρ.��:0�����H�τ,]��)9�X?��7>#�U��+d�	��^A��r�.�O�, ���%���a���$�+�.��uYO��k?���]�)��5t�	��*M6��:��s����;Diއ���l���d����;0>�+y�X��:�&Pu���ZC>��H�H!I�����X�/(��^��e��Bl�80Yp��x���^�|�p�+
_%"�$�9xpD����.��V?�%(.f��&u�c� ��n^����<8Zߺ��ދ�L��O�m�1�����D�ӄ7�e�qɃ��.��j�C�x�,��3�F;�l�8DW[�ڐ�Ue��h�u�aVi��dj�̹�=p���S%X֋g�r�{�l:�R�$��	�|8�#F��:	4��f��,��pƞ��MS��rd6}*��������0'��V`�����^�PSHZ�3�C�$�2��;�h��ʡtzV!�!�<+G��+��i����Oz�4E"x�6�EƤ#N�a;���&��)(�=���2��8�eRkl#wa?��Kݿ��1�c
�V�Ȉr���ÿ�y��{�j�o�HnIqk�B�`���h� �~4
1�K�ދ\Oy���vA�}��G�ڹG�B($��vg!',��aܙ�<n뛽�un�q! ��\�f<��� �k�PvU�k{Y��I��a��oK&����y9��A�6�05���?���������:/�C�Oʹ-��K+�½�&�^�q�[�~3����֋�f���%zc8!�����z�}���:�N��\/� ޴խ��X���[H����8��[�<_�ø%���Gg|g�T{^{���,������;��ᎃg~P=��TǾq���ic��+��F��1�����I�ȧ�Jl^�/���$����6K�D��,�%� "y����2y���