-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UeTFljlXeDsp++qmDQfUoY27mrzLAYjRCYlgTyqv5T64kHneA0v3AlkoxFUpGTzWkxPW/nGJo85f
VZQu1Rk0qw4WK/ZUCg1inIdwCx4nrlceBi5Xy7ULYHkkuPoNMUCyjE0yGaabFzmLUPhhJsuQziTG
G3S3GxFGTFzLVdu3qHqcq1lvzVyjLLvxYMXDN/ex8RzKDXKFsM5fzjSXdH7Gr1XqmXQMmEhr2V+Y
w4mhKUYOFIqa0+tz/YMF4HmnGSw4u0dVN3rE0v7uavJGGSHW0uxxJTBW8bGqDUoJFEq9g5QVQa87
DNPHkrRYAc9vkAzxA7dG84G68ETh4kJSKq8Baw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9408)
`protect data_block
iB30B2n3smqj3UZp0zg/i0m9HHlBuKQK1XAi7RA76tS8LJGzvfDYsJJ9jQgkg10NcDioIo4B3tbj
+fPI998TXpdplX8tB20usEdifL20+GSv0gKUNKlVbfmoIUv3t8lEtHvLM8C+diHG/385MXdG9ZCP
g9jSG+O1yw5oj4f+SAvEowxm01CG8wgyCMNC3xxAZ72q0Oo3bQ+rDIf3jLWfEtbvvsOt03h1TmQH
a8SVeFBdHPExcA2Ztnm5zD1C7Dsc0F1Rl4ns8sXkwgTEXq5R8PIuMfkeyBohCV1JIiscLI0MSFRO
OjXoN3DI6UvMWLPUnpkkmv8Y9LA9rOth+cq7ygJ4Tho3EAZHp1IxNnl0ar86k7dvcwEsvdFurKZq
FkQB9W2P8UcJJrBuQW2HACWcFK1sLaZWsqDYemqepIm0oajkva2LukMQim5LyhIXqd6c37XFiqM/
h3Vg4kEIM4X1xAItrHF0YTCHMBprxXOI+lnaE1CGmSinnjk+oOByoESBcRbDQQcRH9u8lusc45oW
y/b66G3n6duiFXEJp4R3pt7GfNQesEkn2jw+9nhAMcGTovvTr1bHQhLtO1EoklLcK4CrPzM9laIX
P2sXZp0+huOWEK6chN1w22xOxnbgU8qmQhRhRQdHoNBj78xcbYMGhGvAEwSTQmcYRg/70e1T3nXE
9qIidSerNDznMdNaO7bV5jfGO4c4yRZU1i7CQ0HtgyMNcjeSpPDEc92fAyi83dvDnQgZab+NspIz
KpvCPlHUGlsCRR0pBFEp4RMiJRrvftd4G/X0lI9PYTu2vTYszH2kQpmsH/gDZ8B3EWEcZNLXRuxD
iMnNI+KtWk8HR0dphTwpWJPkr9T6TO+Wvv+HJscUAHQUS0bbXqkML6bgOd5Ywer8d8+KwRPqrwyC
16/TtPBSZtKDl2SflM2tS9QNAXIl9Q5wspMg6MDg+CV7pPE6jMzlS3Z24GkZ56Vs2OT9EBsaYb6G
U6o6J9QAk4SmsfzdaLZn4YheZ8RxI3glqtIoJds6WpTa+8EO+1qKngsmHPegpKBuXJlzJsa6l9Xq
5t5e/17SOhg+DNlDJF+BXCszfIhnS5N2gdUpUElLFowzGwbPtuJzh7+LK/IBpL7xkGYw8revj76W
7P/iTY0zwFZzVto6XeZAAPDKRzkAtzZiImShooMKfpOmTEi8r4Gt+nVJC2E/TwR0xYZMGlfxr3oW
BmoF6Afa5z5MMPYsslyKdpc8EaM9Jce91KoaxlgKIdVeCNHyM9KC2rhJTeU1DWVfwLU2EeGWrT0g
vjQhfVrv9csZis0ehU6GbEQ0Q3godbfiY3E/n8+Vw6DFsGQa1b3sRUWG4S7G/2SY0XHVPPo1zjGU
W/jnmsSJ/NdjfYdqB3xuwNpHol4UAULb1eSvwMq4pc5aVrRfAkSub2Y5ZqdnSw6xFtLnC3xtS/Ae
u5OlrrgYwzJ84uv7l8zzWktyyf2qd7HFbPfKMDNS8wF+V7KgsQLnv4oDC0FyqqXWIbLqdKyxy2sK
zCWipzozSn9QHzB0IXWTxuVwqCAHXlVSfHPvS/jmLE1Xasmj7U5weOgeubEP2ox+HZ2Ib5kKZInb
7YvqQCgYgATF+X7R3r4MtMKi9T65s67363khO07t8kHlFgFTLE4mRazLe8qCleI9MSQdteAF+sS/
Ta6EUfph+456Bgfe3KpSoBpL9jjhEi0z3tzZnPpKW3LeiTCd0tGsSH4Wl+VJ0Mvivgrgc/DeB2P/
C/B5Ab/6CDp1Ge2FIIha3e3TTR2s3kSBjrrjbPb8TEk85LhHn4H67tAgieFvYMoFCqIBv6MnOJph
AN2pVhv6HYjW1+uM850vra+ENR1xhmm5P5+62ftBFMGjf0sb5ii6lZmUJHSGLKj06xOMiClVLI7e
6zTPERIFIsWiCRgahq8NV0b0RLEt0cB1FhGIboq5EJoccYQpTSZb/zVTi/xwsp4VOi2AV52Fb5TL
LwMDWTTDwAgIz9hdaQzYI0nuALjp6JpncjY3S6gfBhuodBo/al8x6k+MWwyGaRtGrmZ+Fgm1JMiE
ddLf0lcB/mP2MeSU7WHBZOXdoJEQCAh3Pm0RB5wl/iYa9d4ob+4TZTfjs46JCAb4ylCRf1Nmzxsi
f4i7TBj8UNlxN/4plT2G6K4HVk0XZ+XYQ8A0Vvzzpt1ITHoz87TrP3A9GU4rtnb11cGXpypOowcg
Jyxh+GZvnsNcB8ZbjN64Wh4Mx/U1CPDXQItvsxlqs4K0gZDrtoNgcvM8whUHwTSl7WNH0/DZrMQL
EHz+h9JPIlu/xT7reXzvOZnbFNSa/yoy7KcuJ5Gb0P0B1spljjmtvR5P1iK9eNELxpTqUZjbHwPW
QJtwfy0j8m+ZKrlmzFqAtLJKBEOKfz7UrRfV5Zfsw5zIrs3X3C+KtzPvMBg7kU/lHNlZM0VsMBti
s3qSzXh7MsL5ajiqqKpLptj9+ezu89n9f7Hcbep6LXgqVghVlNtVuGXUzqfKiR5SN6XslsxgZ9Mq
DMEdEhFL4TLWJ5cGZqXIb7mXbGNe5YTnmm8eHbCrhDQFIitcMU0NJcO7gzes4X/aRJXaqm4ORI5x
p5XH+UCux531LKDm+UgnFxkrZnRHnbQfnLHfA+vrZhICgU+rzFXL4jsD/A/3SD0o7nofygrNyeKK
/G4S01PNr9xXUBS5yZiig5Fzf/jQXtmC8c/r2IUNT5jIMr0IitXTlz3cDXu429dv1JcdkY47pTZS
g54DqwRYkRoUX3ylVjNREl3qr0tZk2xrGMQViocSDrdvMR3L+NkQWcJi+fvQ9S3AeGPv2Dk2O6Bi
M5L+NudxKDv970z/UInACYyPZqykl5Tw40iq/HDy8VCEYPO3Xj0+Fu5Vp75XW4zdafT4K61OjsEV
V5hL1+BFEPnABYWsFcu5V4KWJ+BNHOuTBvc+3BoVgRWiIFxPJ9HPM2em0P0B7lG7OxCLZZ804DY3
87nW3aNqSX8ND2tDO/CsxHxcFbzh41rLnNVUcRIF6uuKcFzTsmLZr0yqqB0EfG+RkvBO4m3XW7xc
BnpTRJ0HwTU1bm2cRtaJwFD7MuuWvGV8MKHf4FrByc2nzxcrKtScKfmZCQNcdnW1bdt/Bh/PsyqM
875nriqySgpZz07o1inVqEtSupNS0JgrAbOJYelLBByilPc7+5Na4ShHLNuvOLKLuhna5B3vQss9
utwDTOp6L9gfxebRCDY6fbIwJwGFvt+6qsVMj0OWibG3dqTfQLxciWXpvlKshD8g34qBScf68WFM
0TTKXYwCqV7JOqmL9XDHrBBTknyQjAd3fLMzdoHpMEI5er85//TcMDgr44Fzmq1Qi8QFTZQA2OPI
YaICBvjq9ArLRox2NUGWidCvIuSnR+EFNseHmK8vG+RHn0aZXUa2Bma0DUav9B7cUoL+PU8EV7+B
T4z/G/hXdeIPaeHapDHaPnAo8DDl1hiGPsn9SHExT9Mkv7XNAo9xJOeuWkNji4k1QGwceZI3iD6H
gZvW0bOeSu8RZsMKtnjsjqXeVDmlUx6mNSARdPNqFZpymEQU61SbZXNjcowqOZl5gIi9eevb/QEz
QtmvjApzzmc1ng1sADjvkKO3/2+99wd7Y5SF7ruGTG6WM/6CqCfQT2b12DvhRj9ClrCB5SXvZtHS
+iEZ2ef+vxlxHHVJYJMyBQQCUgG5KiH187LbAANtFnYxlLNtwEGZM2ILyLQ9BERhWc/xFBDxkyrd
zCjjrkd10A9OzzyPiEPAlkbcUqYuVtI0CbyIrxUICeNsy4Xr6xFD5YcLOQZkfakRtcOqDrZJ+oIZ
ecTCnRwtYM2kfdelzeYHvSRcAH10MKARJ8B0wpzgbaH0SNYwgBpvhtbnkTekyqSAwDnoZ1h7m5WU
Om3W763N9C9L3/dv0xa6uONLIwNhqSXRco49kZL++whSb1BsUhIR8xFy3YXNX+kMY6DGMKpv6NXw
uda6hszkhQvuK4hWPckV0gPDHAdB2L91Ab9M9lzsQ2x05vohNRfT+vWgZGuK8bwple16+JervskG
POR6RBGgIc0GQWdVvFwZXNimU8xotqrbY1gl4jFug7bLkyqIF5jN12MZJXfT0DxS9v4hQ1lyZpZO
PdUXiGO2LlJ35M6YeKztjKDqc9GJTIEEaPH7I8sI0L1xZsFk0mhFZ0eIRU97ClnBEYD//1AZSOsO
08n+4/PyX36aZ548zHkGuiHqoyCUdEWYiQJUQ0Ej3TsEJJYvj7i0/61WlEtGLXFRQg/ASs4lmmwS
afu2SQfenRhxqqZ2fA/8ffhjegdtzoZmp2UIVDSZgK+fdp553Ouwa1zjomm4DI1Fz9V5noqfD1Tk
7NX//umJODiNEgkB2h0vSGNV3YE/3YhARVmB4ypcplQpDxFS9S0ERQxtj/33/92//xZykLeOiJL6
riQ+e/2f2l4hZrCoekyCAlH22KofU0+sk4MR1K6v2DBZXsu8jZYVRfKUeEwkpPDRtnMPL7fkVnJj
aZLQTHfm3J9pH8vlfAvKnQ3vPkhwiysCVOVMJjq8ilcguJKT2GFS52toFDmELaMX2cItvYYmVVz2
EZJQIezfoZ5lM7pNuD+qQlmQxfAbu+yku9hKrYzKgpVu8iRl/B5nc8piNG8QDnx/FcPkcaMSlRZI
IwPjaVBI76znK4Suym0VTPAxP4dB61HS2btaAU92KYHCm40beXsItlTgoFAOJ9aBshDT3QU6GtHE
AeklzZY+kEcEbcFAGH9Be0NN6SIiJkiWJv/rinsn7DwvV9HD+sMC20SPi4dV9UgtqSi+DjcZMvEi
vsESeGxT5L5L/siLTNx7Gz4cwPFFPsPwNOmTpJE8JJzNMYflTn/CePjpxMvv8mgU/oBk1G/QtRPF
aUXmMR5snIHoNVlpwT65wFcBJVzF0h3z0NU0C+naxa9i3xYeCfzAJgwk+AMp1HV7yRxucK6w4EXm
kZR8DxjtRj4CJqPVVr2AxYIwY01k+Adcbon2Ue/9IPu0B96gbMjUe6OnixW6uwSlS1p1bGTH7eis
lKxgweHVnUPNrHukcvMDk6IkjNJXfQVYV5+ye3giGR4F+tHprD1pZAMDfa3aLhw8JSqmdV1Dvtpa
JxcUJNHSls/eONNwuHWtTi3lPoBTPa4xw9pj0hY7bqYQSWTYqTRgAKtdCiVCOxs/aHf8UrNVNuMG
bBNCxITVDbv177xFerJ7ap/zqAy00jKQV6aOlmte23jtd8NtXfecrRy82zXhpJ+T0pkHiq+WEUZU
8v7hSoGF4VGGu+KySu2vmBSM2r30uBiLoIIn4bAiUJDd2TR/neGJgjIRNlUvH/HgiXyAnIiByXsn
BJ8ZDPU0Br647amiKtVlY7GaJZDTXshAhttr4HNOZ3D1v4Ju9FlHssd/DJRIT2+2HOcgdAQ4Etws
CFM5eAzKZNsiYBMo5a6DR8GschuLsi+xaiibvrO21eYaWmlwFg7oX8tcjgjQZSFh5jvYL7/TLnEz
SzTprHlZ3U9BwHIV1+z2CX0o/2UsmrxOlH4LPXCxdarF5IojAtwq3kv3Lg+sr/fTG0+xwM7epAK2
OHNd9/qfArHyqSRna3N9eoUD0vzXz7dGt2JJFwkIlpSgPG4FD6ihlKMN21HaK32JjEJJ/IrqFaqc
Uz1/XwipOP//lEyeUzapIlYky8zEcRJve+ws5/CTUVIf2ekjr3pe15oAzXb8O5lg+AsaJT5pHWUm
tBPP+oSz/VWJ/Nu46s/jEtFaDFTn55joTQPcnWulXW36hquGxDDl/cglVN1TIfxzwGSuqtiFBQiD
4XekvsrnxNKSRdjzpqNlmmIpxaaMZaJVirY3iSKujjsRZcukWZX3CVmbRHeh6YRwn9xoBOBTa8fh
oWTV1kPJBDVSY9Th4gyLyI7TgxhUqG+P8X0Im4qGKLd4FkAN6XHidLLmoQbHMlkp9cAE+5Ws/6SV
p1rN7Zx9fxWQFWLCsGpa8ARi3rL//CDE7Bv5bE/leSno5XXS6BWeLJtv3900O5MfObjH1UvVLF/x
nbBJY8O81iqcdS1dKouEof5N5ctJ5qMyeyOimCEUjZA3/JKY57UJTmYvppaocFPQE5C1/g2Gp+lS
sRliDf/jmIOYEHrwOgys57A3iDv6Rmgi4qFF962HehompMEzAaLpdr9bKc4LPUSp5A3hWg/WMdkx
J/wbvhJ+qC6OEdkEblwxBMpotxoU+cN9Lhq/dMki/fFh3suCsnZrpM3aN+FiblssuOkJr+C6CGot
zFBGnhKDUMtIjkRNHQEwViNFa4Aq0Wh/qWi1Z0vOZN/ZO6Ylc0ezN+WDwa7m0DP3KVC7y/5iLXaw
QMfMel4iahARHCFrqDEJoiTaAvCgZC3CHvF2WXRfbIpgneqJajHFnyGPNC1T6K9mG8nC9WGqK4Jq
R6HPwWdGX8cS3aPhfhQpIqz2cHHhfQNuj+fIg91inigVACkypZrO05kbf9oo45k7kCmgfJ3MaJZ9
HE/DwLQGSaRGjX6EcmnY0w9L8nW4mXR2/oRWS4SgYhY6u+72dLaI6DEKSvVJxGJHmTHow3CkwkiP
Fscs2gnxcZZgTqto2qNc6Fc28lp7EPFLgKx8EYsvRWY82HdPwyzEjI2GrCcN8qPNeq0lDY6kHCpQ
cgubD68oWVZFLc1+KYJv1oxNOMrDzetLJgxE+2/QMQzTV+1QYwAtCt8Hzx8dzouU598UEF97nvgz
7qhwD1jGNPXgHAIck9WRrMTLCnqLr1RH393VtMDoPdL9DABjlc73uzZO23s+T2TC5wcLjrtaOnc+
nWBvVSSraUd302pOS4RLZBmAkvDv8fCCJxY8/rCPJKx/lawlPGYYVFcGVzVvDzLel7PqEVOtgjqM
OTSZdtttXEdWVAdXxCFLkiXi7JHNhd4G9puT1hAc+0vxts91zJKehx7UwdXDHWP/2yR9vcMSr8xG
O/T6i20nke47p/vJBk6s3ZveP4Awr8zMUlKca4nNp+QSjg0yu3eO87BwXr/QMQPHNSqA1qHFPgfS
eXCGyXZc4jrmQy+iYfBcI1Isz7Yy4Y5KC4M9GO+x0AZvNutiFrT4AemkoJoQR/ExJSW5ki8twuq3
xft1cbY23UunliD5zXCl2zKRhItOVvYBT2OMZpNPI9guQrwYUkjNCmu2z+dgMG+4MuV5PQKY6YH+
XZBhMz7p8BQE7zN25C5Y9bt5XK909KE9oaOu83EXR1jx8zLdlXeHKHXI249QVoAyLB02AtDjdT0g
GToR1HmzyC8SU+2iRjEm1ThqGm6NRz9DFuPNTTu/cKnn7gRvTGRWr+B1sPXS94IVlJ3b1IH8EbMH
tH/jDREM61Poev7qak2S0T1lz5xKPdFsw/nHoJ3JQC32cxiANm9wrvzGEMh27dSmx44rBXw6sdC6
SyOrDUIXlp8dCzPs+z7T9KBeD5YD33yAHb4P204tUARU2G2kuDg7MvOdkbeB0jCdtBfrBoqZqwQ/
QiJI1TVTAYLF9EPbtuAa2/73S/5mvngBlLzTNot9aeYz/6oXoHlru44RHFi3Z+aEkPM25rAa/tGw
4n4LGcJiKnMVzrnD7nOfUO67bCSOJZHEFmrrc1s4H3NRhkAykQ9UrB8AyqaZ0r7flFdKxSjHzcwm
5uGDi3weFP8v2PrKS4OAz06DPtxs5VgMv4INPI7UrDlsLjWOF3FUlZMgBUCyHpmvPI2iJ0MhP3X3
qyqDHYlokEWEydOG3/VPRxpVOBnhsCCacgP4H6nOyPNaZKMDFiXxFTk5lqRKFvlOAa39sqQCE8Oa
/0rObIiwyxdZDlq5CmncIroak18T179Nq8spvOHfNBRecB7g/TR0kQ/0HO1WA38bXU0+E6qjLfuo
IXr/XrNEpZZFscuraU8JFsKtiCn3L93lYGz8s/fa2+SCjI6emGjfiSeFq216tovmr08qkoCErU/e
qzJsSqvDF4QhdQxgIEzBjTF2UiSuz1TfeutyFd1tU2+AjrZ0YrdzKKUMiHTyfG1KLFaSUmDi6b6t
QiCZj3cWQAgwgJobSvYcfxX4NFkkhfmkTZ+GmWos2Li1X2a5Igo3CvsXw9n1y8pb6I06YFC4IiTP
8VyLzFoylRk3K/vfxXJcvf+zHnOISpMpuo9DrPKm5f6AWRTzLYGXjhGJ/FbpzTeEpEtBUvn5LHBx
pYFvqs6Exaa+APplQAkgUYUx6kNDuZyaLA0PC1FcdRClAPocEX2Q++TZzLTm1Zteh38+5i9UMFK+
2RLI4Twe/8URrHJza3+QN6Ml0v5ZNfWUW3FaSkU9QnuY49J9oIU6SnMWDxLpJoUKfM3iwWfQ064x
t1mMZPEuSLYTx3oFUwfP/eO/DSoHkpRKx5q81Y2RTRm2I7kznFLRYaR+3gfHd3A2mGyZ+bsuqYxR
kJN3C5h2gWjeO7vXX20rpIpbtez9ZKU+TcB729E1h4j41pyl7OoVAHpiUh9ImvtA5bLORetFeEeg
lFQNK2H2xjbIQ5oQ9jYXayIrmTIXDOXrqAXyaEsrghk8qzo5bfagd87OE329WDo8CXVtMijei7W2
e5RFh5CJ6aFsD9pHbnyKrEa+AtLVGkRbUCAkIBpBIc/c7vfmmCDkwiP+2chCMKSz+ecEzd86Ynf0
bSs21zu2woO1N6213i9s7SGJdXSwM1Okb0vRAZpBWGBoyTcNjfgeenqVL230ZR3CD4it/7Dw8Kq1
cqcCdfntwvAWhrTQ3oHXJaFvPv1rP8Kd2ynp1nXvQS+BhNgq3u94KFOtUPY1kCq4t5MDmGE4s1CN
Fcmb0FkPBlrSgIFpb96tMDU99J8DvpXU4vLE3wm7uV0IZbZ4j6bck+ldLnakUYbvB/2kX0RsJN49
7UzPpEbDrsSm/Kt4lQDyxSvhuGXhWoyCGArtD1Wrk+gNJkT2+GaLnZQm4V9GS/lFspdLHMI2tbWo
2PFgzLSyACa0YXGV2b6WnyeC0OUCUWDM7mb8KbDeZ9PPN47mdavfZ21qb+D8kFbs13q8sKW71cvi
3jHOQtPUkhDUQcVk0yFSelfjgMmqlQKAW89GflNLD0KwI9F/dJJBZS1lL42oJajG5Ps4D1BpwXIg
k2KAub5d6uRToUUVSpLWtxZOj8TsTaIonRoX7UmKSKhDSWb9LnvUPh54inVs6kAS7L4wQLgm5V4W
AYI6Nea1yqLRuiqwHg/GPMq5DZ3oklTlN1m2zauWIiq2fyMPjqSGX8fy+/lwEejaLb7i6XnE+K9y
IOUTwLDwULE31wKHi5pjfbIpDLC3d5PyuTrMMG2ZbJ+2qeMsZsDqEaD6NOe2I/QwWQNzmnAEZRow
x4NCLK8WK/LsnCSReHNa2Z045qDpLADmRkBZEe6OW/6545Wh1tB2eO2PWtanBnKD/frirYjOgEHh
dDCat+GgQz7KEkm4+l2n7Y+LYEhLn8Wb2xn6+/nawaas5lT2e4JH6ynlls/xVcn7nTMIxsjcaL4o
Ir2O0OFYvZ8U8ycwclzN8mM0HI2s7f1FLMvXr9O9d1Ui9tsz5NjxkXE4SXkI1n2SxHVP1P7XfuEm
DxGsdeOic25Zo6Q+jQ95rwnQq8K59FTHKxrCvNxX50et8EqwsL9O49wpKw9v9j6nwmVpIMy+ZP+t
xy80hTOk1frGA/HjaguvT2pPglPetNt83nJcvV8Bq2GZWc6nvL5skooqsmoMUsTPEaC4hLo9SrPD
bC9NUHLEsAIszSJvN0Mw72bLQzmKnQTKNz4h6K/YsnREMSMkXTF3kcSigzpAJvODh2nwVqe3iN0w
3jmd+bamk7yrX1VugcgmWAFuC3C2I6Wc38io+Pq9g6lsZxOf8zwP65HJKwD+NzX1EKp50mipr3Tw
sfcgFqaWyyrLyPL9DHOhQ7F4p/ON/lAh+3XC9PdGVTu1eRyPJ/brMqIzB1l8dp1rpNPbEXOl2Cu4
l8/3ed6XyGOSxDwiByUgj14VxskpkSsGhGJmBUi+MUdUY8SyU1D2sZqwVOaBzP186DjotVDcFhCk
XytdZWE6xz3v70BQj0B6U7g5tJKHqWgfm8h5LRQxmO+hJDVHOVcmU4B6uUFf1fS7TIfxwLGctBph
VjA09WiHnb1Wddrqze1rtMgzVRyBGq93na21xNyvfV6kCTL/204bwjEdwSsoruWQRL0erQdCgeaZ
ebcrLImBds+8nkNLonRUNjjX2H7h7Vmio2JxegWDKe0BmxU0TlBdKLEhNHrIfqmjM4WY7R5gqrWI
u6mvikq8MunMIHY4DkesE6zxtQmTCLjD8/D86foJHFiFkctOWKyJ7AnHLnAok5mhfFTLC6YFrx+j
FzcKqeuOmDkHOyiEh0hvzfrKBBKsk8xx0KrRaetDKUc9uWJcDyzyHJ+NLJgVU5lTtMbyjr3ogfLa
tJx5r0lqav2m2PC1xt5kazmhkWNvY18s+gFU48G6Fo27Ib5jKaq5bHH2NKJAEiRi6RZ4j1moYByE
0U5LYtkZyt4N+YC0Sy/lbLGhjJksBHPv6Ad0VLYhCkQ4XRvwWu9AmB1r0ThEiXLkruvD21LfNO2T
E4qbS22MCy+hRSNiCawtgOMXyzlLnMkY9WIVVhEgHDqNSQiZGnxrbD0b7HC/w0SrbljyHQo02RLp
qwiUxWn68dez5RtjEJWQWV/dYINrYK/VQFDZeI7dNKzx55X55CtKos+x3Sn8Tc7tFDbFjkURrfCF
JbyoZ7cLALPk0qUpTucl/W+NL1WhdV0/FH+RqMRm2r/0l6iZap9AQeFHfX09KvuafH22JML/+d3q
6/krhuLQ9DGlqfBaPA1WE3amQWZxCzlDZWVJAhOmmN/gjVJT4YFJy9cGvKW6as5QxidhSJcZVLGu
m7L5gvMVYBms3oOnMiKiHW9DGgs5motgD27RVRt6gHucFjHqIy0tcJ7nIViVQRZRak80BJEdboOo
Z89Ui1lvCSDRTqZs/TP2ZZV//TOiqoutIrV0qS9si8TZE13UqSE9vmjI0zvKm5E2uLzjDeEFWHVA
hP7Nav3CaT3rseNoV3cHLt0cpVCkKKo1i2elxf4B01B8ethfOYx4OTa6oEHASf5wAX8fdJc4ZgQL
xGZrEVGRCu8u+uo4r1A7QTENZq9GGSXv5CT63zbv/Vo30X5c69K79IKQ5ZW+VtDnHaBUybC+zSZK
yDl5lfPSiZXjyhBGqkGCfZBbpRPGwwt2zMRe5mDGuZsScgEvU13E4wZIwho5/wMsgVmoGLOUmH3U
sQeKn2qImknl66r9kR4+a5NEKI8KEmy9fGFPS24A8zcys4j8qP4G6gtMghzN6z/I4wk/utpCesGI
cYs61dmaDh04hz1+AbnAxPwlCcTzjaTPv7sPRryPWQDm7DN/R0XCw3LfaoTSDqmuZ/Rj1nJ5VSeo
6OQNp+X8TkU2dL0hPKnpBkIs1ZWmqzb6YgLVguue8K35pw8I8ZbgWiEIXZLrgWD8Dwlu172vF/C/
3SpI39ylmJzhszg0vtS75ktvdgHkQQpuDnjJgX/rdiRzH+8SYZckTgdYVRwkeB01ClM3ynaqKdLe
JzkBQ+oZKn6C5X04u+KQtUjVyKcvqzqTHz7GGdlt1JXV8iG9t3cS3+p8KM5ku3CaGS4y9u+S3y+j
6gaspdRPJXE812woDvO2qRkJ/iZRTyuCk0X9du30ht34OS/g8PQ1Ah2TbRql9DYQxjrfYMvT2xlL
qCevXCchE+aKmK9eMRs6b/SbOTRJ5KiiIq0W5P9lcySPDFxnnQyWafn2dChDLDMvQ5QNTGifLTzh
cGyy3EicNQmXIM94Asp77L1iTE3mZ9bzcdqazMEqDHqycRiyR+epSxJngfMj9uUqvr/TGDO9u1p8
ggVWfSlE8C/fUHeGle25BSl+OMZGC6JBeTyujbQURIIkxAWMyZJgIVRSK7+praydJDbmJ4v7Y8nP
lp4ogEB7iYWffZsaqDzk9bxwJ3Izm0Kw6TBzf+qGSsYhrm8lNgXP2dpXgF2TRt4Cy2cfmG+1XkJX
qYCfJhTYLHeY6zuIlQdkSO4MA3ROtB8N2B3UVXD2QPxHOMcKb+Xjzu+ba+STtQt92xWKW7E0PC2l
ZHHhpqZ6ojG3V/yhK0wkO63xivhZAtMGNt/DDZFBINkefdVA1/VvWcVazN0K2bOlECEsc9AXnE1p
nhLKQkEiTnZoEVb//i99goHmRfYQhotzTn+8bwVO5PKTYQOCyuf6sbMWDHDU7CK2ODIrpSoF8KwH
dVP3Ab6JVyrjH/pYAg9ikdk5xfi3tNROBxIcQMWvyYSmTMXkKVkYpAEqhry5q0bakCBLHuJx6JON
AXRBSGrCVsRTpKPuFWurrL3cm8QZ+qS9SB0Ic7CrkBzUAmic9w4WCWLTioYEk8ZCvwgIohirzAas
l/y5IYzdQFLBW1oXC4V/aTJBtN+Bvdu7JAywiqHDvOTk9EQ08xq5gBjk6NHhN8M06YdxJd7p3Xp6
orwKNzRsOAXkbZ1/h4OrneY2wOZCjXwinxreemEYvGyZ73mcmaE77PIKqWqFg5+eQ8L2W/qC1j0a
REEultK0aFlzGnxb2Ty0He12z425WAizQUfEzej/lDUo/yXUh3c2Hh0O/3pAqByCIVr66eVPSdDJ
SW5L
`protect end_protected
