-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1tjCKj2Ygv0xlQ4M9WSEWHfx9w0v4PCfHU8wV/ZM46Ogfjf7w3exHD52SerDuYiSAcrBb9c8Bic1
85GEAM5IR56anxnTFj8unUYX5PFSQioNDcobjWQOB6kcSlM5M0ZDgJaWDTfN88b053C43phuTrb4
tcReJCJKuj6oXx4nMbsFFpNF1kv2a5kS1MUSeZeZS2ln1gvyJMDZUnRXo+vYdhinaL0hgIFOIuhm
eDY/wMVDkMFvaTPk4cez7W62k3zZT09h12TpF0RVulwAS7mFKy5PgHu4YtK1cm9bOYwHa0I9y2Bz
C4au8rAGJ0bnlrT5ivlYej3epESGg5CNgvxecw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30512)
`protect data_block
P2gQrsVoPqw20XSSiDjhBLVPWWrJy+yKADF3O10uIcsTS/xg31JSGsUQ9pGSaHgrNKvaT9UArloi
rxDB3QXevMI5IsJsz1TAMgxQJwQ4Z0m1rtFmJ/eDFzVI+dswcfekrf/7wl4ZLE6eYhSK1zq9yFrg
JLQy0oJlivmHnBYG4dp/UOsB5eP728gluX6Kld0MykGu3grcEHeIpt4w13XH6hrTqSEufl9IQSGq
FJdxgPO2ggq9yE2X1Kl476CMFSkuYaB9RCFsc0cXxKcAXvmAFvIB64kEvXR+vVFhZV0qRgm1DFDp
oBn1c9wPceg8zCwFPeHw5s5htrhGhn6rk7+pa/o4TwXeNPC25Mp58WsMEGqRZlXEGeeF/ak860qo
92yq4Ho8oP5grl0lkRgYhsVM8jATOMk/xmoHBNLL0RpDM3xMzqFMXX9T7Dx7BaauIihD4gfjuolQ
RSaG5sE8zHN+ymySsP75riDAthSJTWuA6YPRIywRomT5WRuiO4e9+gn62Kn1r1+oiLiYahMsQnZv
KPFOLX9duPkaqkmff7dkkx4sHEpWH4qdVjLToOO3mV8h27xjyhSIwkiuvsLPNHF1rDjvf7XRtCko
qDYjZ04jyPPD6Yq6XFsMpveoKouFB5C5oscXIHtuLtgAapN1uhcKcb/TNlH/yJLPIRMHAgvqCA5Z
qthPiUCbg6a17BzbH0GyW6h0no35TIlLyFwlbMFv9b9e3byPFSwGVxoVOn9PpLl4xubljlnDwzSR
OR7vFw66ug1lGnFzFTxDIHIlajQwE4DC+1dkNyvyBYpqrc1UgUDDwD9PPJFeQpG6+FKMpJHIVR0+
hVm6x1N3dvo/PAnE18kkMGQrNbk+dXz3EqhOyzMsi1WjecWl68PKZqupg5G+X5jxjB4XZLJHBo7I
m+g0YQn/nH6KidbvRzHdM4dz3BHAREYXc4jGxXoOCjMrMd148p7FY0/6RO2A8B54ExoAUM3VP/Md
SWxEL8JeuMX0f2Q6lFa/hUxOJuaxdVBeZxCcNB3bwbT9NHRJKXToNndEDCLovocVZymSC5wDtmMx
2bAZLWobfTUpg90iIb4m6QZjQ4VSCkPgV8mlq5xRcZ/Jhf0vQf5MqlCMNHTitUaHMSPrK/+9f/zi
4rPacGP4J/3YOH0BqE1yL3X0kq6Mh8lPUjc2Zjp01oWp4HX5BC/LZlQztx2AfP96x5y78pvlh6Dk
iw2k4K7SAlwuyC3eFJ+3WT0DIXcTW8vyMWvkxsrmGo4dferzMDnMyCJJA+D8s481Bkd2CS+Z+9sR
gdanC0K8IuTDOoGsOBdVAukrY6SF7SbBMxbFYG5RKKgmN46S77FO+E35h4XshZtPAXgIS1ayeXcK
nPeN4f7tm2uVd91AL7ndS9nRnWAl8nc9uwG+LyHX56++bGPuzTh3Bke5Gjn/KRxUqdfLLbAZJxod
wACwvtdE6t0qaa1h96X/Vn+yzDcd9dLkuGRt1LkwTnu6u4yQZ+Ha/TxW7dOo/+FwxG0KqGlGEKOs
ZcadCrL87H0yYQxfRB1OBJ7bgbBRsUaomRsx1Z7m23A4lnXZaN+dfKS4QAjuxdU5xqzdkdCY6jEd
En1yY8U1KW4XCr1u0RY1YBBED3GvRLR/esTx3l7KqTmJH1sbNATd9QFeLTqND0CIzTCNBTgZk+Rk
5M0OSFkzuII28s8afp9pyrWkCGER8/iHWT+a+ACQpL+5PU+LWG5vXweq62yPsHcPBTUAU2llg4At
8q2um/sZueBTbgw545lF7kSOb5TNF6GZylS+ZiqQUoz2pq1B17/B+d0wYmfj1cjJbv3+mcYMUPR7
w4E6BGw0fvPa2Yt8FySfX7LkmoEj0CWoANRS2HfXLkjLE0iJN+4MROBMYdOXmcU2TWhQg9RTkIyi
EkZk2PgsmE4gQOV8oz3Vkpy176Ap429E3/D39UvLcKg8+8CCBsij/3iM8EtrRVUreNl9NjIsh/F7
xOg/zfPdnqTNzY+xKFpjNGDzi/2RFE6N63hiOm7opmRO3gilYm1TFwHjYcVbqLs4hAJXCkqk3jyn
Z94AmVD3emOLRmWYO64ew/toZrNZvfcRM3QPfQJtEM89sU2JkrNmNGP4oZCOYyjdD291z2sJtWK8
G0bgV2MPCxUZGNGHOUFc5XtXt3eu/b+2CVWqiVTnEoVoLlzhzKK8t3nMLydqkzg7K/AsR9oizWWi
jm6361M1gWwYf8l/l5zfC2+d1ewHdVy5G2N2K0QgP1SjAdBwV4PtoQ6iAnMuTHwPUxKRbFjF1DbR
iyRNX6fntOCklmXB0yRUFWA7h7j0JLHU/+Db9n1hByDZZhFYEsWGBE16DAunW91QaJNkcQphth07
2bg1y5n3Vj+u6cPggmFkMAvxlhnViWwcSlNNtCAa16qXb06WdMyTuTd8kCGcrgyytTcBA+QqEOpI
g/uT+4aETNQBI3AOuFqDW98Rjjva94liRvZvXvTQkmueChefOtOvaTVMQAJiB7635NVXfsPXkabi
2n5xcxRDvqzHHptEhs/Ct4uqDd/Q0MnQDKboGCTfo1rDHHVKI1OJIVj8ud6teWZFZXyFcYuAZAZ5
io9pPDtnkMr93+G5U8NQzc5Aq/+AcFcmeq0JxoBjCc22PvS3sw4Bim4jx0MBcAVq37g1DJkBORPK
A9XR5ewqo00paNqqTrazEtOK8yvUwpOMFjpah7rH7gbZV3r5wYccsTmP2dUMrU9QjpB7O6ia6RXI
6ZWOMzPSSHQUzxuyRPLyl0xFsndr5dPFkORXQG5xDCr3iSk9UZwA7LEsScJVoRiyQxz0/UUQfbY8
wreI/43ovabAC/2ru9wtEhSQMzWf96EP05tHrhkBvAO7jgPp7pe80eSa0Lxr69tQkxXWCGzYzZ/D
I8kwn0NxaB7kXaME4QLlrwzRjN9F0mCQ48cl7UwvBvFY2h7EJDVpNsakyuvkgDtlweGPof//y1Eo
4m3hzT8eNqcOTg+qBVLwdre0MH87wMPZ0OPpUd/eirPysHOGRNaBb8YBr1zAPRUEugIdR9p/XErM
u7Ic1UZA9SCAswozKLZVEpn805UmoaQfdlXJOi3bROueVShhWMnaAYRWA2PwpHibJUGvdY/e7vOg
8MF2cGe1HNJVRs71lQWrmnS7qow3UFa3vAIkwnhL1ieWrbOq6tNVSKsXafRiFzaUfPs27TjbhG/S
j0zaDXP5SJ44MtkETFF5Lo7SdIUJeGECkvATWpqqqBfViCgQHZaKn4hAgLlutELBs0QusdzMA56+
9l1KZS/j8IZaFiFY87Ti0Arphse0I0wMgT4Gjgqcons7EASRAKaYJL93lsTbYszMUh0FnRWbYHh9
SNjyTDYYRC0PfMgzJO/MRVCwEKsprrr6Ntw8pAe2Ufcb4pMAkEdMH6UHvQPPsevjEwvq5m2Mi5kL
77KbxZIQN+2Gm6QkzyUYiYDgYNvLZ6socCw1xMzkWmHmG/Q9RjRSMEHYh9lFo7laxtNi4Y8led43
pa6S+mjlohyCm9qBqp6ieQ3Y0JjBFAz+vOfp2B0sY2JgZ3qQyiYKsdcj7VAfh6akm5pen03+tnLa
rcFkgPYyuMgZ1YfnacfgLi9u0Q5bjWcs7nUBtcaft7oGoP/sqDeMkmUihbd/Am6B33iA938aEu5C
uxICPtXS2v00w7HVlGXQaCRv5zGcGUwlNEnOAj6xtiYPGbRC5jBSwsds6YiuvK+deStt3AsfzWeY
upAwlccJPTXTSbb9TqixBsaojudKiaW2sjW5QxtPPOIcytW11NnDCmoV2cGrYEkjGANDiDvJG27c
LnpOMS5wCVadSS3yyC3wVXx684Ljkvx7mR9QcaLVvBrymaXBM6j1qCQ6NXzG57DBltJ8cVTwhyGG
KjaMxwOsfBNYB/IOHWkfe9GTZjehL9STkDuBID1n+PL7VmLMWaODKi0KZuBTmnZ47YFIl7pYuP81
NSLHIW07Bsv6bScV37HPMtMLbiOzMUp+yfXT1WqLyJkwSvzfBFsTzppnPc1wEomewME75W0gP3QI
yVmCnTFnHXixjVw4QrixMi28SD+eUT10KjZGvocqLXRXkX0TxHWHuHjViCM7ZPOE9hWGdXEwveFU
dO8+DnoVlpgiXQfEwXyeOVe9dBqvfByTEv2g/HPV8srMSOXf2bYEtE2TKChZ84rPDyDbH9RQDkAj
lzwhdjrqQjnrCnwZeVCaQU0Ha5gsAJcwf8KcJtQu4eN5lYBMAsdw0Hxfoa2HT1rO4kC8xVo9GcFt
8Z4229i2jJF0K+7ATOWaXJPUwDxcNmoofh3XyQMJMPldyBHBfu0L7Wg6wIrovfjoohSUFNB7VR9Y
a1K3g96nzMhS0ZuX8vzd6ZGHa00P+Qo+NFLaLd32bWLdsjS9DqRupMxbpdxWdgU5Au6OBgeZV3M3
TN6+ozsgvEEVLpt8+20YimmD20k6BIogfkvx7jmm2PNkAvLtWZN85w1pyMfVX9OqRHIEuHMoPnlN
kMaOd1rtg0J6l2EYnY7fqKI6LZJgKyem+z8vbd3zuHYoNPLYq57Jh/0+bFxrjBYNtz2+fbYcKX0q
1qAK57OFnPNOEbzv89O+RQueQv4RludI57xsFjS1EEX1p09yCCbVUj8PiM0CSyo9anKHlaALy60L
M8DxiKETJXLdE5cdDlPiGA08wqxkePbC9BVTWnMmcFitq3Z07EGnBfhXBRcx6G7wb/LplyGE5REe
Adc2IlSxXlT32R6CZJhZJGqEviLmg8mn6p+DEaDZ2Y+4JhNF+t+iu2lG3vi2R1cCr0MifyAP6wdo
eTW5ywC3A+v+ojMNXmkb2SezxNSeuAmT/sla04UTYeynYRrFyzV1q+pjss6vvY+LjqnzzWnCzHNk
g8htK2Wg7VOW74Gwfj6oHP2nFz3+kjJZtOWUHu0r/n/qBiOsxEwwwnVF34sEC94RURoC0baHTvpt
NzRlA4j9SQHjczZsfycDD6YUIcqnwdlpOraxjvi6EPWfSQePC6So3bVNxEIQ8r9De19VYG6pDoy/
HjNJeOvlxX67PzW8DqIFD9MQ9lccC23dXl5UtBu4WpifJV7kAjMXSuh43DlLe0xNKC+aLFkhI1jm
kfcJBdXutSdC4D1Gu3jP6oQKuXKP/gkju70l+EskzB67BObBlKW9Wc7lGoecSurkATnT8ar46YqP
1b/9xuJDBYH7obDPD7IUn/xUpuO60XyB7WiVvEJHcFFCuCApIYrVg7rF2O3vHTftAuqm6pzMx7Y6
9KKXwpCmV9Ji/UlzmQicTa1DVzQ8PwkAQ1eOIGfFzf0/FKSD7JtWyWNv8abBweLhnnsddcbNYIng
l6jmnPN4ZqqTeefv3qO2jpN+8KL60Cet1fGvCKdprKpYPaNxXWgakDI+kqb58UN+iTCOkVompRhx
/WgwGVE1ZwFHx/QquDFV/vFF0QTFQUz3vd3Tw75DmM+B/h0XfILtfDUO2gKA50Y3SM/HXvGuorbW
CBlcB5xYdsWN+dibOqi8Ur5G5Ius+1NDJEbMtbEN1VSDRDt4D0SwCFgpHvg8LiLdtQepqmlEsjWc
A47dxfkCfyTeONLJMC1MRkCUNoMb9m91s4xhTnrtQFg0+gX/c5tEyGyWhJE/Kyy4Dmw33LbO8V1X
rhXwDMsNnx00eoZ/yVr3mJnhuEGP4FUQrvOmy1l1jCSxQBUfx4I+Zw8VTgiNdkwN3M7fNSaW6/gP
VsKPyKNKs1E6fLcyW2vpbNt5SaoQ7lzeQAwW4wrg7cc3GoKAlEmx9CSYjsDfBCVIFaL274yfldsC
mW3p1kYFWqDgEIQv/ZN3k3HkTVRXWvdG0PJ0aSRW3IqFiznaezcvCkOJtRSgyMenklEYFOGJ46eh
DK0AOuCEwP1KkciYfkPR87FTevwbFtDC4vEUV5cQm20uE9+bS9BuQwEIfHRN6LoZ/t176vNOAWzS
alXMv354iUIoxurZrPTKFG+V9f6XiD9hPgXuAjRAx5s57H1qHJJ3YjZiXgkFQd0jg/QhCGR5CNVG
aiMRtBn94tuAHhUG27k/5y/MUs4O6Z8Artu3LVJjt0QIqLwmGjumRbBb2ceQi3fllt9al0+nisgX
ZkckEoXhWQSAh1KebyUZ3FtwaA9O9yPdFZhtdgssCGL456pCHujcPyf3LyT7EZZFyLXSg3l54K74
rhzHY8HeoZAawkeZgACw5kh66WA63ciE9F+L1sNBI0loBqkBG4mfK7YddeuwCECx/CdYwBYX1mAV
riYEiz8bOxyRiT0FiMoYZzpj4pBy9QpC3/stDD6+zNl/Ebi0oEt9rVEA2pmIBlVpeixC2nck1+zk
wImIenm0iyyCPbSBtvA4Q2GDDCg5FMSJbgrJkP2l1jRusK72xe1QW08f9WdbiyMxSpG2rgn21e7z
xSpMWSFfE32M1CuoQM/JkvidWEL6SdCiPpz9R7zB0c0ZUWJQmGqg7vkI0f6wOVgxc2DtZen2OZMV
hyHFakjaXMnXcpRNDWMqkDGhPXj/IJS+bSsvrF5hJ0iIe1DgfaR9xl4b0LDK8HkndgYU+Y5dgtlZ
d5xh93PsCLw9i6mWEx743jgWZO00VQt/fLg6zBc7uvbnM6WP9c903VKepbaWw9ZeinNn6/kkkmyu
77X/rNzH+WAhFTDWOHTL3OwZcLd/U7bwRBPD9XXC6AU3aKtKpNZ83i1WHWCwQrl07zYBk/jDe9fk
zCG6zmkzePGmlukR7c0xQF671FroayXCcKvnSa2ddxC/RCT/VOZ7ZuRwKs0tw0Kj9OgfUBh+49zN
gX38OZApwgaERLtQ+F+YICOvpzWuJ3+XqlsPOTVVZjS4B1BX91Gnp7lml1fZS8J3O8Yj0/3cZZn9
grCeNFrO4CSft8LYMFgHC5lzEIVzfhCskFIXsCRLaUUFfdl27GtKE2ykAtNd+lKyMgpkgBILKtsN
QR2+v9dbcBqGoIRx37YwuYHy6O5TCtUUMEtjfHnVsQbJzkKiH/YTllBKqIbpt/jmUEFOWI5G42Ty
JCkYzRiIB84tyLF59YHVB7pc1CTcOw72P7S7WJXSqwxCfPCK6yDSUc68ZpOJ5WJTTWWIGCcZLM/c
v9YRDjR/adVMRx8ETrqBsOySoLsonkt3JXo7mqxKNYREkoMYqRfSMI5XV8WMbf5fMYIxFwsgq0lV
TWgTV1OsHw/Fx6rHEaaxdzKynNW1+CLc3HFxrZGqFgPIsOkgB8pbjqSdJOm8UEiRexnHbFf8DJaW
0UIn60jqHW9yEEciSFBAh4bOY/Q4fgGXpmjnS0OtUUGlkU2Cc7WYTiwjzePnCm1to4q2UD0j7jTZ
/9BWSlROWXjuFto+BLCNpdcKPz//oXaKG6wD0aWG8g/Z9TNjrmv6vwLsW5RqHRGo9z7hZGa9WnIE
W4MkDR3DzQGKvUjklqVyy/vWjAfjg9RI05WNHXAoXBxGmQllHMnwT9iS3KwNY2KY4puH/EEy3A5a
rDPfL4USwr9Bg2lyzOFn7re4LgszFRil38llrYh2Hdj6pVKAvuxIjT65zPbKdW7M8kSSH0mdivd2
5s5eKvVEjjsccypCo2DWxrE5NducCR23taP9r0s/2nGFLH0E1gpUqPDxjxTrCZCfUeHI9YLTAtIb
K687giZ6I83ijIr29qUJdrF/yixfz+fd+P7Vs7lfR11TGe5jrxB/1vW9MlwpzXR8JMkjI0jBVedR
DSZ7oOj2J8k2De86g8myG4GlYohd2ZsytMFBWVt2w/22uCtCD6R/JjH2nOlcJNK1P6Ux6ie1DNcm
PpYtk/qi6jrK9xdO3+cUg04bInHK9qgDsRhisM+NbxUzBU2NHOddqh3Uo3pF6XeNCmvxcalcsqbn
ZDYkxxfj9xOYtAah2eXwUsPt+AFTxdfKRavankQfVT5Wx3bHh59yURh0vnoX6+C4qFN4TFlxfQrx
NFkBVDB6U87zcaNe0zcKmUXEqXEt6ErtzZH2JQUpyCicviYHtmOnnwwoacp+PubYg3+M1YTF6/82
hvngGUv4KDHXd8ovwf7pF+ZBqXWHBvjP1N9exiDrAGTRt0z0vcMimxD+gRJP2+pXfNoo1w3jgPBz
xokTDFpeeq4fU9aVtDYW40Jd1hDahE79W/j4mAp3D/goi9laLGqujhBNXaL89bBKZ0eA8l+y7DWN
F7HOOkJTyNPiCrH70Rpvsj5+DQMwN8Q2FBb3HndBpycIsu0SNeVHRzw3eZkm3ob5L6mlhhMCXgD5
xXPeFS4CuU5sDruRgGm8sGTmsENVlMorx6lLsT5Kkh7lpMjLzaPhcHsNuifPSoB8+08N2+UzP9Ll
gXQegKsH7xE9uTJwsPWl4K4nwwNu7lFkYCxA8AFxrZdPTBl7/MlOCJmgjXm+ABmsZYqNtZmDC0L8
k4HtqkuVG09JB34c6a4ZdL+yPcUEdByU1c0dK+KB//9Pp8tTjTmW3CY/oNnJwYeGfSyLhGQi3ZmF
gryNglQI8wlGB0wVgIgCXjxCeJeEcF75Is49hDlEZfwbhkIj/S0+l9Z9mY+NzOvoHOF3pa4cUR4E
6tt787/5+RQnwWrMwZjBe/oQvlGonYfEwLkOTKw5w7u2lL3pBEy2fgzkjvJ7wQilkjl/t7aN6s5p
QGXy3OY73OHsNQzI9jaomMHPsaivytwRF5FR6bAhKPgdjORkb6KAXF/nN3PbfCNlRMc4wiRCi/AQ
wYxwpFMOt4bHkcFpeXkwOkPoPDmFvGTPkz0SE3EY940FrCX0XS0UhSFFMoZXBApVwmUJ7NyBIEIL
GcVjB511PkFSQFytLH4S589T0tSwfkt0WXdUU/2/XhHMF77QT+swt4Q+GGWso5reR/WddZyiTA75
DjmJJZWfgMFinJ0aMCErIj7XTVFv137oM8ea2lzsrUdOwCU1kHERVpLnlu2pC8CE2wAbPUZzP/1S
FAD8VFErZZumCMjCf3l4ZNndD3V/Z25f/lI+bwh89h19HGmI4QdmE1C95zru+acOsMEruHprbTov
tTXkWSDztL+0t/StBUhDO8B9shInEdMvG++ufE5u9ZmTX+yWo+oIcii4SCFcmftq4JDKeVm1mAWD
FhMJTOuRehsuUo7U64M8r4C27TaCXsdqY2y3dggS751tatTgmSLtW8ghdA4j59cS6THa23xwpvyp
w9jb65F5pNzunfejubVrKD+vaS96GmsafA04GeGyUx1vswvMn807YP70jqyrUAL2PS8kYAUZviS8
PWVecr4Oh9+zF1rgkwn0H1KM0sqjvs2yVqc1js5blZEp+gTGOsLYAmshx3j8tdhsgJ+IFd0ignpl
rmeGqe6BBO8FTING93FiM5OFsMPgW8vr+xFfPW+gie4Jkr4CsdFDfV9p22fBJ6amUvVizJBvxT+U
jQmYLg7J9IYubuZJSbX/Zz/OBNYLV+0m+Xx1Q+0vU72aHV6BhPWxltEqkPTI3kmJVnuONqbyMC9Q
cQuaOAA79ryFxryxR2N7TLdri4SbRTlPQF6r8N1JPqjET7ZhKqkNzB5oYMBHMycYIKCl5Vm8Fq30
q6mVcBTYTVfHEMMtQBxEbB+AW4u0yMjhqadhr2A2PSuXADiqaRkyjfX+XQLpB8yBduEGFxHuf7pt
lECoKe/6ATCdP0wQ6byc1zZ3wBt8onk+CB3n6kaJrpv3pUQf69leg1ckoGeN7jEHBKGqRzsSsTq+
vV1jsNnY7KLJ+XTTmxPLOYZk8BF9fbejAp0JaUT5Pge+G0UZk+dh011GKXdtfDGWIGPpJ/ACcmDp
Z0JxUrOs3zf6vPI8RSxrXrBnynqAz4lRnp1MgVBTw08PZj5iTSz8nRqyMrdtRhwV3REX4RDaS+gn
UmhxX8olhmeKc/pFC7EtOcUIsaELfSwLCDM+2EEfqkFOUq0hoBhvOeNqiLI1edBNwXaKaDTempeo
nVYLPalhQ9e84u/HBLuqD8r8OgzgYLgPpZmN/FV8Fnj1fi3c/gN2bgqd5CuVDD9ztSlKN+tcWMPY
Mjhf3p367gPipYQLN7gcrQpxst3xi8qgniRSSVFuvDkMFw3X1fwBvk+Wil6gdRCZXTfHjH2YBzc/
Rf8nzIXA9W235mdKGxFORrcqCI//GSUa+BvR9cnMkv+2qFuGSjnwRLfDVMH0Bq0qcuE6VRb+LHZ7
tKUMg5fKqqXlsCr+JJx74XW55If+ys8sbsGcCoJc6uhZU52Btd1Y941Jz3dbtn2ONLcw9pHKce/z
jxupUgFjQZAn1/XTpLL4/nrhMEHAQJdswLURjNgH7OTQGHYxwmssGzLVeUVBogwcuvUznS+iE0I0
b7g1siIvcC49k59DvDkqJ73Pyi2Cg4JiG1R+hzZwmtUF/STXcQ9O0VDaSSEPEsC2JBBP1J2Tpdx4
4qcMaRVEdLlVuRTc1T7m4TfVRdd+WpL61zorIeBUKh6xGJ11Gf4P2oAczZSRvXb3trVKg3wFltpx
gq2dzVOmAOAszPSbh1L49xiRfNIdyi+Hl59vwqvjG8Nn36xQPgKdfiXXUToh4n7FXeGnp757D0R2
/Uhp655XNm/O8XYbEUBMGjsgMnPKqiUuoLJ6v4nyimiOlq7yuWnFX7sUIQtLtx+V+fJ4xFE6TpW5
QDgHniQeYkde1gcvK1JAkSBaqaCcycIjOpy6ArBa6/ADHfRQuRNyn4zvIN1QgWDuDL46t8/xa1lc
m0RfXTjo8LKk6aOmpWknKdBf0MXUfDlyiTC54j4FnkRUuI6mYhjeRnovBvftjiY3DkFgOUpgwOk9
34fXKLZxoc5OXUEOvs5332vzmusEv6btGU6aR9WkfZuQNVBAeMk8GOZUdryP9RedyXuICrewbI0B
8QfeNYWsvclszjodKPDMVJxweDWJ8jl4qdnQkIWAldbk5OJyZBxjrOInnvqFrSxrq3aU8Jd/+KKS
DKNdDigBC0ivh7Qul8mfJba93eK4ciFsutpZteS3uPDx0uL1d1q85GuAv6mKnsrCdR9Rp4mXFt/e
8RJRtVU6lp8KyUwLBGMxWe3TyRFP1s20P6yG1aawzLo10KKf0fmwbJeQA3sgZDVI5/8Y6mcrHA4E
RqxSY+A5HiRzFZtZRmDx6mlMwAIS5iIC84luisrGQ+sOz89WrPDZBzHGqmgk7TsBYbCqnr1xSCVq
k6DXEF0ULNEMo1L0QqRO1r5pz+O07jIZhnLu9NLFNY2NteGcAgWd7VXNcI3lABmfNDrHhZqVUDXn
ACA0/GM7n6WG6/5G3Ng7NsYoZ3GPuar89f/zhbptBrK8X4u4w2OfO2xQPqc87md/VJ45Q5fCTxsI
faEW3w8SxVPh2ym/V7xl9LIiHHlKBiZdvBOoMeomnztw3tcj1picNtujCOEdAlZ7larM6aTOVwmm
mFCbNVcdVrZ8Imq1eXQnBrZ9rrqWplcKgGk+R6yMoQDfDeIQ66FcaF+nZfjvDVkGnojGZb13mh9B
zBuZ1+uQ1ZzTJ0WhrXzfBZJ9awgcEByAbBWZLg5kFAd/xB1e+cUOYZ/wrtX+au5U+kV7Qq2+e1CA
qex50eLBlyUV+Vx8rtrpqiXse4+dS4xlBU0EGoXgiFBNRbj2pqdrYUyDoftWvMpMF5mo96xcx7F4
sM6XAge42wY/hDDvl6E9bpPIb49cHusxy3YH6v7hMz7eJ+XirvVGo4oTHDGMlZniaO5Bpp7Zyndp
bQA4Us6HbvfR1sZeT3abjtDmQoHTVd7fAj3IJ2nMKPFVV+CDu13Oe5S32RfsJH7n0/simkYMsZnS
AMrrJ0wFz+sdR9gOni+IOcohXH6eaXLstaMBQRoSj7xDrcfn8QsYM/PxKyMZvGWKKVyWIeMqQGyu
C5cuk3QVzG95uCHsf7ol1/dzGbgiXmrSUU/JHTk8zfPej4dPfuhVwUllH9XfAEZvP1Lr6+iA3/TR
kwBlo0tOk4KQVS00800AW4U8+FDKwYvy/I5Vzzh4LWuy+ecnTGO1lUFcv8idBBmLxZ41bO6gyqGW
Xec4oxqTh0xIiM21ySYvta58+sEEWVMI3IZQuKhZA0C05mPDEY5ooSeP/WHkojQsgvWi+lH/fnW6
6Y3Gmrulttnx4hHlT7KLnTQLjXoj7uGYdm6Kio3Djo3NskyfzhuZ81/nRWFIqHZlCpU0kixc2n6j
Ya66EkjCObVnZoYxZNG/vm25YZA5nyg+wet/8k2qEAtAAL4FFIUis/LBL62/CzL08qBvPqEsHe/5
BYkip3QXv+BJGPfBkH7otEDMosI/wkESryA7vWvrOmv0RakNsVFW4y6uIo8QbLtksw3E1e8/Db+7
50q2NcXG/KIaqYYXgXxct72CHXwy5oHJ7t66Z8fe/r3kzeuKcTcmGXVD+AgS7fL7dyaPMwdQpA9R
AjSKbRDr3tEhyztvbj/Af2UdLjiu03Umv4buiQhL0tcSKPiZTZGfnsO2q0Nk+OIUWRFG6nVbv2Zu
CEh8LW5HuwPwG5c9/s3rM8M1OyvpTbWbv7TXfuKsY6Z//j5vAME9Z7ynI8Q1g8kdWkn09PqXGjti
uAN7Ae0jc3hbkwV5Q0Y3IFpWjM7+bhLsBb3Q5YvxLCl4V18rcYkr7Oo1sxvKHQVywmG6Xrxeenz2
zrrboygBiGWO3+z4gAjWxYaEpOEmfPxvaFpWdt+Aowg0FFyhRdxOFJ3lcrGamh1iWaHD6VajEGh5
zeAXVG9cHhZciLsS+Gx0g0T13Vhce09Q8o7mk0BH/h72NXfBHtp/2Qa+Cb7LdunEeapataw/n4lo
GzlkGBcz7VgFdvYCHtcs4+njLsfBf3PiQ7H6vpEBV8pwb5xvjhjrY7KSMzFB4mHer3aDgpuPyzGJ
x3gZzgEY/OUPTIlaWp9WQjN1GhV9PXaqN7OWdLVSSuGQpqPESXpQ5/99Dng6ZZsRcUU5XiAgh112
W5awwf/U12nA2045PYQIENFpjQVVeVUYmIX+8Ijb5VKdF606N7fR/stqtAKGljBco0XoxUWcx2Wv
SjEVMmhWryZMUn2HbYM1gvlRW1SaDlvLfhUrvGJRRfJtoj3OG9/AFAw/aiU6zf6zis1SIpuQr3OD
uLZPOke7dtK8jtgvvfwQ7Hqqd2rZxt52MUS2VEbJO5/fji4wgdgygNhSyYuiq368LgD8zoeUn5Kp
l8cRBIgP9/2lVJ0RDRpLBuDN4yV4vMnjrRU5yTt467IhKwBHIlopOmZoFXCZVxGeANSMu0p9wNPM
6SHn9hutVD9zUCWnBgVng/BQ+Yh2t7sfPQ+Npw0fHv51HluvXNuLUQPBtuupMtFpRt7NHmEnuVJy
AA1eEJNU2JecCrDWQgkJX6028PsxQOyVaA246OdY+aCsZh8tP5rWc47PUfkAERTCe4KBKMX+diI3
P4Ds3jxziA64HtjYqbHQMJ9+cDcO8roc7ZyiqnwK2ePdEqYtm3qm7p/8lXneom/L6SfQ9p6m+qig
POB/RWPc2Quygt+GXYsIcH0Eh2QMRiTWnWkb1w3q3Xb7zGTkKqetjP1bg53WZy+r3wbTdWrDyMCg
JUhh5T1T07VevngCPMpkLZMcphZ76qNoy8EoG8wOU5c7tB5pAKTsARAvhyr6W6Y4Q/uK4lINRlAT
jdLnItEvDyyTrA7gnAQyeRhiqmeltcFaYBaB2xQypU/V7ISfmpuA3d6N0qeCiVoL10D1Ml3IV+y7
vSU6Vvs+22KHkDx7q7GD8+8LywDPxH22U+zQLixHfyxg0beqnvJFEKBKQbzsSX4o8BRiRItKsSY6
kZcTNsl5IDowJrM1evCwxM3Hvfw4d0LFEwXOasmSJZLcMDTi8kNClOAHxLdxRTZxwHW2mhxEEU6I
ngwL9MavFnEdS4iHWdKdby4PbEwYASkLQRacaezQeE4mJxFTnTK2sOyeAUOXakLIFyaqDxCIjRoP
/VM+ZTKNIa6I2RRw8L+tpP183DMoYsMSkf2HuTMCeTooSYH42PG+Zy0R0mIy2byg/5ASGpFYeJ75
C9tlbBKY9GvT0Qwg0m+IJILdT/84RF87SVu05ehwJCS/eBD2mqyiJhKK7owFTrlEGqYD1t5cOIxU
HL1dCPKmrZnmp5vw+2FmWZ0vZBReOO5vYbLK7KsjdMBo+z6wNvr2a9vS/cdAg6RdvzDvSOJuZx9d
n71/Yuo0Oa2E+HNTeSvoBYNTG7zqPL2B/Y+3RsOUxzXkrLOgfLIPaKJZqVKFlrigPM3c6qIGl2bN
8Es4ILrSmDUvmoaJymeFrvfWz+xvuyDgC7IStm5o+7PKRUUMOKECc8NJPTZeprTl8T+gOPlvAILW
2ekecWqJi56gn34XHqD3Ds3gpyZM7oiiaTXfF1XaacSi7vkCzdUFW1lmmRJKBCzWQ3JBtdicqaq/
fxckW45gO2BODMbmQbi+vI7TgcgqGtLo1NJY93xqKxQjU0x0tIvY/Sez9++WANKiUUiiCTtU3edd
uxFAM73SseGVEif6o8LPO3gFoawil0VP3z503j7CSmzIvKeUeVvm76sdM+GY9mr4vhMFtwGdR+qN
Nx9eWC711Qiv3OWI3+gE6n1jaEJ6xLWzN1PlPaPFOO4CGSSjI68hZ3d14XHK0L6kBp54fbm8sOxt
IySHIN0lFiCdyRzt4B2c2DiRnfFyl4De6E6cwV+FJqFnzoQ1tUUWfOJhcw/7aet4dj17+qc+1cR0
BjE+N7Hpvd0gx92lLqcZuUVCTCWuG+cNN0SwqIBrOWjSIDFgG17nE7XA1lxDfNNHuK44aL5l/RHg
McHdOKx+8GWAv72fgk9G3BIyFvTr1bFbOiyorP2NK1GFcHEj7Litjny3JabiD6wCS/AVnsImsvt8
x+Y/6+dtplbZ1EyCHRu9dfXOmX+COKsS+yOzkx71v0r9hLcr8wmvQ/F6IX1qhcqxCcv5J84Zz6l3
jKLY3FybTyDBn68H0W6a7VkAgyRb/te7gIWAplQO1qtP21yCfo2AvFepmjQDe36tLPwniQ5uTWCv
SBucbwLnyFysJOjMHgO06fukRFZmxfHBIyE89Vut7wAaUfuZp8gck/LfeOnK5vviXtLPEBu8m+Td
lD3l60JfOKsp6g6WnE4AXFed56Mrb5yhKXXNXOLmgfflSv+ivxtXZaAq1DlerLzVIblO33mRluVO
a6EzlgYd5D8tQ68JdVn0xuwu3W6tI0CHMdE3IKOfKg86agZ1olNwx4v4ywUbfg+11AtB/Unq3q18
ABLPwdZhJJUyaFZ8yz9lQK+wJZlMVbWDSbizJ6Ws+5vzhq87MLK1vmx10OQ0bRqmmkgNz3LxMdio
ypnxQ0Men3tQiJzjWEVsDCD1h5AMKd4bNcn+aZe01zv6oLI7dfVyJQtwQfHU1CURqT/gSV4WO/px
eD8VNECHM5sb2btsxJ4v9Dcajo22MZsPGnFhY5Vx2qyUP7oHQcPx9UXL+F9tUr3PWzq3y6m4Gy5K
N2AwRJc3gocDUULYgmUBqTurGGgszzoHQRnCs+9wO0evZzjdZwRt/fPjoq/rLWH0lJC48SEyLUtt
3IvyrydV0XSeQeNtj9MjgYuyDGrTFMo0WTEYNwHuIEDrjnp9D1h7b60HgCAKpTLbWggQfrOr0t6m
Vf7LaRknrNmI6CVfuJ/mixN8jmEsfaqHYmMKEYthNwTJrXccOqbBVJiP/QF/nKheJRspzNecbg2o
KNixONlI58jgF5MWwDhNpeKVHnv4ShzINV7SP5ac6Q8ZDhoClaQOE0b+4QiBfYxoWxZa6B1lMiOJ
5mSMeY/mPHV2KW/PNQS4anXGdV18HjgaLXoOPeIQseGYDCXXl7RL3rfqBHKH7e0RGFE/GaPJiqYe
vD+LfsKcC6e5Z+GZz2VdMQsukI0n2w6AAug2oLhWuxaCDMW/g8q1zw3NeShZPMotqz8fgx1xi8OM
4Uk1x1UKT5wpPDTTvGflox/YoEk/+nhfOHCA4h5J6Cv79pSjrols2iALmAnBeK9crDhFzZNCPoRh
5dSY26a0aR9rWuiAMtBf7GekUfQAMvoBUzJ6yW9I8xUVOSywUKNW1y0LN+aeEMyU1xVf1/Ynjbwv
p3+W0WnypbkCStoG6XgCtkOrM7UTHdOkQRRnW9CWwfUGClm59Kar6UW25hk0rDjK0tQ6DOOeK3YD
90hJksV/kcExzn6rNUB9qYmzO+DekbocCAsY4krK5GkymyzQC0Q0it6At1jB4PIU5e+BnzBnEXR3
xZNldy9wY6rk6oXTyBlOmdJW4sZZenZ4UknNb4N6uBlAYRp0OcV51N+nAzLyckcM58RL8w5qvQMH
dA+H8OZn5oA5afS+wgj3jlPjBn4M8kOEfY5ZTTnxhecmFAGQitDZe0u6N5/vx3C7n3EbsvH3pmUK
v07+mtEEZ3eyt7IF4/7ZYEBmbkJesP4JS3xAuXsqzEbpW3LsUy5vpXqchILj70XHLkMB5Enj7sHM
NuSaFpsxJXwG8TgZCFc/P0j+jhKlxmCjlNUyR8eeN7cnoEbWtuYjpqkF4IRHbCJnQnekZ91etcYS
rlSsmN0OirT9jBVdrJ2TY9l8vkbQ7V4s9F6f1AdjajdvJUI5P0xxlBNJllDhWtrgN4S8/VkOWn19
JrcYb/9E1IMeSV3sugRiT/NVF7hbDVQLh/AtpUXBURhI5Eag8PkTvZH80vkckx9uVV6rG0g9arNR
isQa0OfljYlrghdYWDrB4udNTKBv2/mJXICXe8QiWPnO8VEfLy7MzNHmFBWqVvenamlle//QS1IM
hGsr0Gm7UDR9p6TT0TQfaCsGTnTfiZz4R3rBOHM6bWI/xunulpP8GF+CVSLR5RMS26/iUpk5IgvD
GT/MIb9grfu3kfAGn20456/oiWBqhMGBaJVPJ+lTrnOPijo4WC3QHbIXIcMpIkOzzfVjhwisWqUZ
ub46OMcUnDjYL9LxHuYQirtWvgxMyMJh65U34pnSpR+rIRppiSkMBGUL0+InFxZMtanwVgL1e77o
brUG6jqW30hL7dmsjElCHHZ92CsC4WELU0BpcKK8wlxhbODcaKG4eKtmKXJuBAJ9LYudpGHpP/1f
ggzbK9czXknLmy+ubaV+r1UOTaJtLE9Erue54jVIDz6FYrYXmKAcy9ssUTWiduESxZZnvmtA31w+
9Iirg5ZzvS+S5t7TNOn9q+IKGUOSPRGXRNGa8I+9ngjpJP0VbF4z+iQDP1l2bwn39WsilSrebiAh
fRwhbiF8jDNOY+fVgAPcM6DbJhaPYi2/Fz60PWpxd7q6AuXfmoDfFnUzD9LW6g1vZyK0w7k/iCbN
N/zsjK78O9zya+qSfa6z3SNa7GJKXrVemWi68rNc3HGpSovR72kvnSX9FpmxarH4RNR9uLrXMd8j
4Jb5p7lymgV5IsepzEU8ydGiSQj+TTrqBNeTDPEQ3E6Nk7Z40/G8pPItIjqgBgYx3CG4pVDSfM/b
WhqL5EwbahF9am+9cTUrG/zcAuv0/xbRsy+z/tAvk0+Bg9586FgWC1BpyxyZLRxQqaMudwgIPxUC
UIJ0vRCD4+3HYH3d6jyI0pxwwNAp8aWaQxpUbph9z4+KPWz9eAevbY4E3UiCK+lUJ/HmYAr5M3fv
VYx2oLN9xqsOgyqUgFJfi8oKjd6LOLNFNoKgPrrR0f2Kr+ORnlGuzpG//ptDqB3T8cQy+ifwFiBM
fk82dtq8OQdXV7UB2lmo+RoVT2bRP9f1kIOSTB8RLzT3FDcROctqxIslVjt6r6mjp8/YfApMMd/6
YcIZIoW8JzIsvuWMN428BomV0VjSLLpgAW8tKJsi+2+eIavziG1tkCa1qcnkk2RrZgp34v3h8Co4
GE4R6wUSixFCuCsMRbPChDOgkrgpTz9F84oP554HzepeD93cdVE5RVvsrqsSKArFXeq5WGWMysYt
QfqlKs38JAlXpZDoLzI1K41O9Ir6kDeIKfRMEutH+kYKbgILB64ORX6uUoNW8cNWZ6L44cPwsPvD
4Kuk+oAYJNmMFHkv16wBjskcvgOyU2yKzPXlUfNGLk4D1bXWXcd/WnCKOd4quTP/e3ONAXnrptKH
1QQqUUlUY72r7JLKa0mthQ6dJG9gayww6zCJfFuAzoy+a/GMXVgMIWfC0KYnFt4YhLzteVOEQLJd
+2Vzg9aPwH+jfR8y7w9bGqexLq9pwZsUv/PTF38QInFasBwyi4g+qtdP2u9vt4luV0GFGyo5xE9b
b3nVBNiF3byU9/3gxQw0BCeRDwY7ZTT9a/1DZ40K9A9z95YBRafB205dRA/ho4FiO01nhKYw16tX
4aJbuFsJJHCk/qqXcs8yJsJ3Ez/XJzrV/BmTPX4Xd09gxphGoEmhvKarw907FDML/1j+bolFnQL3
+lZXJXY5S//Jw59FJM24CGSJ42C+Ws9z8/nEC0fZcS/vlSdoS885aSnWiD9jw4EmlPDV1SGmcre9
kFbu6Pyn9SgADwOfK/t2MRPGTbeyI6rw613lfdSrNm+3UgIuJX2twMiDV3WR3yiK1g5qxiVZbZkK
MPLPHoAJOjgLhyBArt9Fi5XoEhm3H1XNadkudDGxOI2+gnZfmcAi86zQcrHN/z6mIdLGjsBMrk5L
RwuBEFANH0BcrBGnAp75D/l8JQ/t3semGXO//71OLFieu2QlI4zq4YMYKMM0h5wzkzJO1K1NNZTX
gNlmjp6na1zzBrG8MOJ+R8G4xG4/Bw4x9UvPPpGUOExBkV7nQ6MVTcq4b4zVG3tczSC4EG4GbrWO
rRQj4/ldKe6e5GHqhJkhP9n9XFWM/I+3jQyWo7ZcfCO71gn2ZdZivo18My2ytZ4NuRq4pVaK/ib+
DqZXJhsih7rfEjsDhxjHy9yl2Kv6I/rp+GEdZhVciA4RFPtP5IWKm+oRkznCEqJODw9ne5xLqwP4
FAWhajWK0WiAjQ5kJ4fQKvgrRoHKxz+MKDVJSlFDiA+FkPPc6ltJ/n/Iq+H1RmBh1Tz7CZ5yDjrZ
OAwQy/S5tHyomrgMI3Pzdh/0ZLr1gpSLuemS3gUGoeYftiW2flakjhOy/tZDs5BqTmcLUZVToV+D
3k5+vRN5JvgKIF9FgkSuBV3u29JRLeky4PJC4p9+P2vG4HopVSXn4uPvZ8ADOwML/Ywj4beseCiL
KTLSe1xwnlYJ3VOr+W6paW2LTTx0iqG50KOdB0plsGKrpO7YcUKRDX4k+nbnA+hG+EDbUbUjZGIU
KksqIqsvU/ld/2xvSP9n6QDS55nliJAUzuzsBSr0113fXTL11XdWOX9JiXnnDXrPveDhVQQgKT7D
DMsetRvIwag7EsALCp2ulcOoo1Zn3s7LSITUrn5mTDFTcrGhepRHC3no+VGM+8sVClL94HVRXCyv
LnphZz6/T4ExX8TEwdnnqrBV89mAgn/YvReriaoYmYqOVaaNaEKarSZ2aA697YrqaGnqoUMcQyoM
B3gz0Jrxg7cgupO9bAykSZLzhsKAys1rBLI2q/hpX2ljDcXLWAgpImfGj1Jx2MCDxSCfXZCRaiZ5
u+q/l2/q4kHBCaAflTjd4znceGCg5+28vUr0vxxRfvQXPujxunwrAF4c3AK3MCKy+yN2+4JtiaAz
wNAU0a8wx3W7VOoxguwiBaXH+VF23tvS3v4G7XdrHZ1QioBOVF3bHPfrLxFC8L4dSJLpv/NxrPEK
4wyMogvY5JmIn8lf1HguhCGz530AVcU/6bGPrloeD5V+ypsXJ1wPAskW9xIO/IvyQOsHKmrw3XoZ
pWT74e82xzznXnMvCGD+R/ULl/GJ9EsINsRlt827DbVlxU9hcaE35sQpbFN2by2bhEqCZ+wa/CO9
Vo+NLyyXgDyfTF4Vp9KoEwgifdH4sdYZMjJjAVSj9NhAEA/J8JUbjikYbpfmXSfkFks89Siy+nXC
fYs+9dZKtLjsVg+XtrRI5U2EBCWA96FiwzzA097LqzWwE6c5fSqN6s90+fgKtHfDyoDZ4rESkOI7
G21uKCu8/pErDOgWOmrR7/R0W6PLDr3h+8l8wpKbo4Af2aItSCrj/4quAxmhsLSEG9NooxXhOr9L
89Zj8/O7YeS9IwF2z5mPYuOBtf8oaY5CoF1Xyd+d+5YA25Q/ExBkDErC1iCsmXznS9IzOpfK8Yne
QonKR921PNsM6OvVC2YcdKhjJJgTeHsSGJrWbjSWWq//fSZsPkUINjIYKHEgOcI6Cc7TfoyuwuIQ
hPVcGh87MnAG/6roruWDGxrhYwb9NqE+yfNfw48Xgv0rU4agREm95LYzveAyn8fKfMSuow1iAAXz
XmcQ/2woi3QhEFjdcmCkIufsS1ix2GdpCEAKie+GGCeXqL8Fmo/PyShsT40kRfi0VvQ5NnqgxHi0
bQ7Gdq1BxQC/+updvObUYFtOJUMY3QqQNzHpRuMxm/1zM+O34EwlqN16uNd82U1X7ylwkQSEmhVQ
T1M62XSb9B2fh+sVkHQwcERffsx1wG+T3UCaadIJOtG7ye5DBuDg+KJclWAU5plbSG72W24cgWNZ
l+spIsggz2MWxJB+4jQ/J5aDLUxSP+5gmGgqMxf6xPOQGHGo8KR+gTWkQNqPK1RkhluTP+7+PBPc
uY08pOHg1OTtw0q0WamZR4E8UI3jSNyOgHTRBVNFgbhCsZBJfluE+g5IBx9TL1GZmZ6yauN/V5/c
cT1pFPerbScTb378HhBL8DvCHr6mK64NCLWwt3q7qF/9n9Ja8J6fkC2qBdQfmdWj4JVtuqnumixo
JzNb7C/ortWrchNjna3N2+SaAbjaE3l3YhpOPM+6B9PtS+6rHM8qfu4GSN3BFZ8+APQniwJPtfVS
zyRvJeiSflxS8fOm27dutlZ8/wAV4pz66wW+K4ooASK7NFC1EptCKt9QSGO+M8fMw1pBjJVlG6xz
ZcZwtBjhOPdrpkRA0xNFOvCe1+Nq+bj2lCb8UdRLpd6em7RZHhjJQj90m6uWPEF5yQ2DOjnsRsxd
uG6OqedYs0NB/kIUy7GD7ywmr1pv8UWC0/YYhSQOn0htNCH54s0E0+ybcq2mADoPLudomQkuH8Bj
8ckX1uEEBy8y0LotJfsPnL23eNf8ogF3afgj30vcLcqvhIinFi555aqK9gxkKdHNRqo3UOMIdiOt
aB2HDlTqtCd5EbkYxUGlZtIK433cZdeaX+Ed0qEqWnE9Yfdqei/qVN+wq5bIaTkte7EPSVjowFwd
u9zZCVcxIZK2HslUrAkqVKiyT8jcr2nN1VriRZXu5bqvfij9p6ZXSMHEWyAUcjwXReT+5IH/9gr9
fiBgLHV6aTkvdcga2lE2ETN7nn968iEq0vvg02GcZ67V2Nlx9iowgfvNS5u9KDWeIaImXFAhvrEF
48EvF885VvYpVJdByyjW6OgtT8QFZ0UoEx3wH9pAM/+REb9WKLJNQnXvDObxBcI/gXaefZiIymxg
GwirWqCFOZW3Jo7ePNVXcuuJsGf2aGsTBerAPoK+/R/r+59uoEwkgCaSRxNnKG3vcDIAxFYvurTX
zoEHmNu99S8NtCciri2Zvg3lgqnTIiK9rQ4fn7JMD4K/+B2AOn4E2lpzFFeuxXLw4WKThPys5GL/
MPgyF7GQMoqkSDYI6XRbORGr+D1ymhsECpNLuRypSXc+d5qtERY02J2dJtauFqAw+p2nWw1nItXX
4/+pm7vvbRzi3z1AqUbXwP3v8gsd7R8kqKAuciY4wQEHGPxevCoGRj8R8vB5h8EBuetwFulPCC6M
ojPQBch1n3m4q8ukgtuU1tAGHbjO6I9pgwTNidcQrP8mAz441NtcuVYcPUQL2dpxKsXtE6A94irJ
09rQ0dvbUGDOPXZxUn+7mBRnwqC+R1Yrg4ZapWPvRg35Njk9K7rTQC96N42mrN1Hhczbj/VGGXCs
uY7imbJmo/F1xhEmMphXXFDkW3u80YX66BwrneF6He75nCmGENXPE/hOaxL+Pi4yHQE3xMhdNiNC
wUAswc3YJxeD2Gi++UeHHxYCyeV3IFvgdcf8L8TRJbR66vrVPKdYvoaBcUGRQLFp+UI7QlmoYFZN
+FqYsQQS2OJiKEwFnsYububcOlkIzkJ61XS/Hg5yzS/itl/V6jntuxJBhxArCwjFF8hyDUvc9jBq
tBFERwyYi06cPdkaZxKzvyrdtCVCdqZ5mg4X3l0Icq5p1V7HVt4BIUmufRiSWEFAwJeT/VJ1o68F
SxM6nbDtYDum/dxHpWAYPEORJNGpN1MzgInDDmotEclNMMgfJH2q097UsVM0StDlghrOdyoDkLgr
8paUelMqlnaeQyA9ylz9/CQL+glpiA3CHH3mioLku4aSgeOkYLMx4DK/dsSI5LuFJCQJP88ezEmQ
rqWV+BmQ6RV16G3kXLOcd8JiQ55PsIHADOkki8pPZWSlaqzgvnKy55j2kSIU7ja2HcmdTg1SVBol
IiCFfYf/2H4R4T23OWo43rOmy9H7TQ1YAj42tn//FfxeSpULBgUdL+h/Oi7k9tihT/uIKmcb8Xna
1FIMBIkpzAvObymiTTASeUerNablpgCubxhpuhKtFjkqKm8CKIRQQ14weC0dtvRMch8s7ONHAqdc
6dKXS9pmejH50lmrCotIaZMyHAH8c/J2/jdnuxBGOjeulp4LxTUog3J1hENsvPDfKmm0mcMRdCXF
SKkgftt7vKkoIfTNDvq49FXAWgbeCgDKVtr/Dy77XI5NZwfulf0nFiwC3DBElgOko2nyWFZ+tU9G
7nWEx2t9w5Qk9HNwN4gRLlenlF5gMqN/nZcZVfyqKsjXHjB1z/6/3RtVZcq9UXhKR4aeDeu0DKG6
sSIPRqbIqjsu5wCrY+Bo0OyxU3ZN3EC74sMFaLAQQj/vRP8i8SpsC5XqM/GRj8dqnJHuWfSvI1ds
nUaTWc6q5cH+50Vwlvb8PB2Y1QATzAb0eHfmFQ6S9RKCr4Pu2NZVmxXtx7HJMPL0yUUR2NpE7hLc
Ljwpvn0I8g+eDQr0a1nBO9VZWgklK67/qIjZUlbo57kUpZQHpnFNhFYd2MpeJAYaxUIeANvk5vJt
5AMZ4QTrgs9Wl38tOF4bgAYdzPILqaSTxLg0ewKxcFGunOu09igb2gr1JMMqEPUYWmuOEntBQL89
uKRtY/0/uhNY26dZAjUlPYszViJoVi2Ylj4/sD/Bukz/ev/ZtmXAlEMvGBEKARAcpJ5dAYYsW/6a
d5l9NzykypJDQ0InCP4QnpC75i4d0BvsaxnbCeZlm2OroDPVLxMPtAb+erNJVpLQGvyq1TC5fiT0
YkieM6OerwTaJA6IFGazj4N5IEEV23a1Kcl3mazSSuK1eQMZnvHGwVU9owJqkL3PsvLVxQJqk/wU
BXNZnFCLoUpoYcKZ3qTDyp4UyYEOhvX73jaugbrGsoK0vNLcn7sisgeF/To9CzgJMHOn2SF9m039
zKhnk6hz0ZlrUG6Wn+QRP00o68yUbdT6vDP/WmV6SbZPVPN7j4BUj7qdy7FKlNsQrivF38sZaPeY
jHqA38Vn9DTo58ZyaHgRgNaaU/HkdkzkqJksdVKzDC47Pm2GVzNy1nOUwQQ0FUwWVlZuFUTB/xeo
A6D83AQscUt15hWEhR0Wfr4dKYaXnn17m419YnWeqExpZeujGNHijcb0bgc9bUyT7G0qz2k1i+mZ
uVZzz4nNtVvABQGmg/mtLdwT4KrcB5yMyUvEbAHWXpR+HcarGi0WBEtL6yteXykoXmRwoTo8tnmL
fduJyM09L4nUlhkHbUFBNd3TYN5pujab0+3/N57mVLRFfs2+RaD8QMfTipvEvjWjzwY0UK+fRahR
vY1hWNKEuBCdyDVTVaQEDbnciBVDLQoRP9k4qhTuXUkuhTeYHb6r9WQCcUVFA2KL73/Q7oEWXAcJ
3r1zaGU4FxrniJSSQUMXqTBcvqp1wY16FzyH9UWF5m/ZP7D8aKjamd6BqMJtLR8LXH/OWPKDWsre
3wM35fOiT/03AvSf0oDE9VJL/Wl7GLc8oTl+ESLWxHvuCia6w3XCLY2zaEPwAwt+1yn84mhxvCR1
n91htzMBsXotuaHAeHEHD2qUkDISRAMU3baRqp6zi7xI7hs/V5IRsgsqZyK9M8vu9WopE7oac2y1
p3R4laJ0tRxfdULmlh8Gz46VJwoaeLNDgueJDc1Ag3WXBI7OPl2jY0Dgk6Nbq/QfPDZiN+LuIMkk
lXtd3utWHSAvyPS3fHrBPkVON/aBpGkfwHv0ikvffA8YtyQ769PaC0ofOzV2v4UwP+jm52wN3geA
N7zgm2MC/Fk9RswEqOxwmIbVC5lXSbGLZeHdot83EFT23HSEfOVUW47QmZXNsmOtg7GpzADoZ1z1
+uWkhH3q660a8z65Ekt2ZCSo68tbQB2Az05J+hX6tm0UDIsCm632K2w4hf3pugD0VvtTq6T+FAC2
1+o+v5g4zkf9GqIhS/6bPDH+L22h3WRNy65CkeQt6WFXY0UEmu3+LkVFWaYM0VuT6njdmVHa9XuM
w3AN3sdipblQY7JlUM/+RzC4Ze5jdsk4u8ukvlwzRgzInpi3+kRhC87s6hcNYNsEMC9HiWktNNMR
LDlXEs1xf52wqvkNGhPBTXur2YVJ3yKggKgJXGl5narcdktnaJ82VfxhhLeCn8J/jW9wpDVfi9cJ
caB1syni0nX9SxIMSMj3RSsbZXdOy3UsGULJjexBe7jfCrV2pCN5u50AYkGWXFV5K9Ffaw4z6Qyk
s16VJljEele7q6UxWuFF1a5if6Pac9UCP//9N3Xd8bLBg5XZDpcjkAvhg49Jv8Y6MOsUP2IqY+Ch
vmx4yBqFAkQZPwXr57lbe1xHdpFGt+Z79zqLmb0ilsSSRkthYwTpHSZWMBRi88iYD8pWC+xNrO2d
OE9ntdxtltCoGgblZBfUr9yYWNZ6RJzUZscffaw1lEluAaH0p5UEnQ8WC3m0cnjyYu+9iz/TmqkM
Xoeero/GM5csmXrgZueAp1mu+NC681Lk+S82jqBeSjZzj4hI5NAwIVrkkXZNAvn0VwMr/upwvA9Z
owfo36Xtcg/Nu3Ygro+3aELHnJEO8Y2DGaCiey38guIZspPRDfiD4bnBcWwueGOI88hjHdQ/nJvv
PbwqkDcY0HlE79dFMTTmkwxngzAThQOm3cxVrA4vFD8nAOXRKYRb3FXYNmEbz8811AiiUzj735Nk
y0M67/nTr19quQ1t/UH3lk9kzCSq1tylpnSH7OzE3+auyqcX6thftccWbFSnIAf5h1p19zcpc55+
oFpBBm7m7ifFDnDcWeUWTrnwWlI1qb/oHtDUf4wNPpW6FW/Nd5oEYIXQOPbC+HhI5+Vyr3YeWkuS
Wm/RohEfxEOstlj9uXybGMa9eDP0hafxVuknqvfJ43ciQhq9qTd8d1KiW5M21Y4YcXiU+pDgVMhV
1jFz6ulRn/D5TYHlnufDbvtvUeRSO+DlUZYDkM2W8+irTx1hlrdW0WrTs+AzCuB8Q8nGxCznGixg
rYIJOVcB6PhYYd2grXOmo0657ZqDYBYNvJQovjLAhiukF3mNaKVUp0EUQF/o/5znsWNDCL6z8ovH
PqoTeYbFPip6vSw/QUgrTYb1Yl5NXOMZUv+ppK3Lxcc2cPrI6+8xaKCP6P068i3l/iRBV/ymWvAb
PEDp7l6QTskH14f7SnYrq3GeexCac2f/kVwHUq6r29L3ppNMlJ8WBvMISTgWtgB8qSury/EHE6Ze
biIGY18TbfRfiIBOPv9erZdHi/7D8foZnIREJ2PqN1t8pwlQu8N0xDLrHFWj4xhH7353y/6nLylk
MVbp35nbcjc65msl390iQ/uWn+n8liZChNgxlz4ckvpjVLZKi4WMMhhiCv30XhwAHaFA3WRodMNC
qja4JzYxYoIrQ3IJLnD1AzKEcNYB5yu181Lw1NuJFeXTyqXcuybUXJvMFnncX4Xxby+kSIBfYxpR
BB5eCeFN5U0Jfh42BVL6MKl2QAfrBCaLCwH85PvSNLYctpFzKeHqNXESN0WdegajKpP5frH34ntv
aOcF5T9Hlsn4XBH7+BM2Db0c7r+Gq0mQmKfylShdnQrkYBOj/QgF/ELvDduVFmoz+ukhVxNydD3B
uihgTuayJGAwhTrdE39GyUaU35kpavNwTKW5dngPjQcWYB9zEe+vVEMxN4SntqfVXB5ME3J/mJCQ
+x3TKM+fQTqYOCdXpikIhspQJrrRp6ODTW4M52IUvnG6/+24XCfrc+TgzEZRcStwjTn0Swcg2mbK
oiwmTZDiETzyn93EW41eWGwju0NDjghb1ZxNNgJ5kx08Yq6QfrWUSw/MGug9v1R4/aUYw3ihFmKD
xLBpJAfUOTEfKUQyJe/9kLaqR4VRwcc/PboPMb9OGS1QRcb+EmLUKryKirtAuoIYA0yUf1+x6RU2
g3fsltjsRPm8zshT7E5VAhjSY+AkgG6vBxLyI8d8FOIOpidzIN1USAlrgGkloD2RlUsh5yhU1OXq
+sbUWj43dRzz8rzBCbr9XyjBQn16C4LfiDq3DGaaZqNvycoyXRgmyy5frB7HOWRZI7dQwMd8Deh4
bG+AP7Hf3r6a53IXOZ8fbr+yxinA7bNoilnyVRmr75ywyhHLr+yIkfBekOzrnZkyGe98/NpfkrgT
Kn/JuncBa9/HhpccXTRU/cSEEc8+GCgrOi46Kt4FVnTkHC2xWWscnJJgOxHNqpxYt7VpQHAbl/4H
7r37XlivkCOb45LqqZzglo/x/GQqZ4sQnQImKgYrZnQgkBiOu4vZfYd/IlSrPwx6wVmxEzd0kzFm
QDpEVXJrup8vs7Yzuy6kLuk31xg0Z0CjHTIS5F5LuHIdAh8aRbgHCXfXdVMUXn0jKy87HFyOwCYJ
uu/UjhG97h1IkgPx6C6EQy+CH5kJqHAS+U6PngcHFv046aq+eTB1nsllWruL6w/ERXLpoPnJtZ0W
T61V0Ucbevrz2pgCBCU6JMudL7UniIhFO5dGknRQ39LuLpQhxVLMMfaxJL63iRW4GLCiRG8e9WrO
m1BF3DpJ74yLs6V5nVrOq8HLv1V+Jf5raTCf7PJmF/OYMr3rN7fNonXceEuMU0Pjsy0zftJSmlxX
yfZZkHISUIBhlhcStO5QIa6I38IsQW/apZbi3otCTgDUi0tX3nlGlxUrchfHii/dMYiAw9GDUj2a
HeXkNj2B6q3M5NB71psOmNVSBU0Er/FYYjy3mcUoLHz6eMVuQwXGZjEb2mbaPn+K9AuumiB8lc4B
PSU4+GxZsENLk7c6kcZLc5Pli68A8AWguMvfj9uACe0gsFFEeDYOyQ5JXts7H+WkOzGxsXcJ2NQf
t66BYnWwa/s2RJaXOAmBz8yd15yt9lAaxCneFJkgO0W0DPwQVWQ4d2sM/1QKRbUizKD9e55ha5wX
kao3/bVlbE+elfusXn7GzIye2kWWB80Hptcsnw3ObwgKKyvITvfKKu62hJCPWt/v9D1bdVxZd3vy
ph76uDVFVACrFXqj8uX2N8NViLNYmZFpxhe5lZ3xTGBZnbO9l+b8W80aKkXuu36dgSxw14fjCNgv
RLF9K83xtIqsJmwKcf8XEY2OXalT8OQvszTQz4LbcKgQtRJHMDITqyKlxSZwObdtCqXBwvLQQ73a
iip1wF0CE1lIqc+MtvpiVbm4n6J+if3V91clJ/KIEcemCCzm6KySsljtgWYZJnMrkYkUs9L2aQ09
mTx1f0n29mAizLyHq3ybp8OQ5NlWRfRzwp4ho4GAOl5gHjbSVv/2mNCINKSpk6h5bnpCKgp/TXXF
7amCxHBBlEiDj3iBYZ6eRZh9236wBhr6PuTdBrR8HJlLtZbiMO3+5Y1Ry6yZebs0jn4bOlwmH128
UyH2SLdGYF0GmLbfLLTYDNW/DMbccLqvHRCwQfqehAea7wz1L70P3MER9qQXQEO6ZI8apHe7IkLr
hcjbQSazkfobzISGWW7VV02lEH/L8jbno88rhhVg2cU3iDsGOPFu2ne9eUSqKYLqB5Qn4NOYDfn0
n90WbVitB8KcKRUzS+oZFz5faogS/OSPETAH+3eNNRNR+Q3wjvpXn2NjwUCepnA520pnV1WCB41O
jdosmJBGM3Kx0WQzw0+OYpVA2gP72i/QhrI/MP/KVwk5Qdd2x4Z9sTvmlSpf+nLPVhnjQRpg2ghk
cnonnUV43j09qeb3INritohzrFiAipWU/A3ESx5uIlTotabTmYOfHLNOCGWhAvxDHKxDYe5Ipt8y
6a64fv34tg1UjMvzSgzxic3dek+EFFQeuNQ2Zpt9pX/hILRQjSyD1kASmGyj8WB9GOZ3QJD1SRT3
OyCDQL7Kw1ULDrqaIWBxH6j/kyRGCfPVEmwdEFSY6Bc2Brcb0EPXK+4ZijRkeEnqQJsq1hi5ymgr
ZVGhJPT5v0zpyNjkTG7Tw5T3FEHT7/9PJLtqCr8wWY4OJhonMd6tC45gWxf1p1M0JLv2qNzDqy93
727u1XzIKpxBXag1uelK7+8mX8IxQRDc3G1nxCs+x1ZYWle7T0ZPZWS4bTEEuAXIM4fkYrtEatm+
mifznJtAPmr0PhTEBSQ0IL2yWpP4opLVqwozSNfq07rciGCyFmcAhGwMpcFRjJh3TSxQsfdRjujp
IBPT5l5Neh0Pk+/KLbddVqtGvq9xWlDQsd9bi4UJlZrPHDoUVsV6i60UfjARhfpuDk6jYn/R8Yi4
5PJTI4/6hxtOjVAijSslNrbR1/9endTAxkjtoe9JZ0DDTSthnwyudfrfIUlStBEwtPFPjMjI1S3L
nZ8eXWfaJP/Qm36+vz2+U0rsOaqRW4geRsb9ieZkT805hxysPikhWR/QyWv3z8XeFgsc1omTF1BQ
E8E/N8jUxfmCBLQLNo6Z41cr4OL9uTq9vggA4Vcd8e0DgS+eIG4WKkbplSXAmc9+OpO2i2KXvV6k
p5Ms992xr9fjIXauIxfXSRASTkUMWp0PruzOshseK49hBPKTHqHeBH9h01vCT6RWN2leC6RyXyl4
tPg6YI7Lg+5po7puxyuFtnLoBMVO9sgCnunTpJHD6DiLHTtb/I3t4tobBbp+ypdMisTPz2Pb67C4
kNkhJilo8bUJvSye+VzsoPi69QU+25eaQRwQMpQpZSX8iEPu4A02SPbGg0C2QWQVfthIX7taGelJ
ZzdcA6P5OL7k9Byae5SpOl+pFy5Z7xHYUlLfpuf88enp52I8/6bfPQptSeJvepmkyhdIFOlhij0H
jfmQwrJHlK/Brav+TEfsQQj9gcJryD7HOqkXk/AM78f3wtNFO0BiAxmIDuJosLD5Edbj27+RsI+E
Hnc5yuGauopoDScoGAIMehopWPBwJGNu/nqIjJRXFh3+NvPKHm12VjnnlADweWzvo6Yg2B5KZj9I
B5B2Txs9eIBxbnOwcgUI6vA+5m1tSVbkgtnHaNCeaDDKI+rIDC3D0xscRxLghBW250MjHdW/Z+Wa
tCJzvwJ8BF48vDyrmYipQC9uXkY+8jHZFVIjSQqNQDVIic3/NyDRnuBWKALNOTivk9L5e+t1oNOU
zflabGlNCJFRwLcRnnIz4oXrgw9w13n0GulVdz32hlHXZ+G+I4s/hw1EprxNlv4GzFAIMOPPUu8w
n1uiiYsxIdKzcHmVtVt3rhSV/W49hF6Lmq7iD8YURska58w2vbF75+yCU6p0WTEWOsEFCFuLlTar
1aCnR8413RQUasSUiae5o2TN6C9WDvRxsPEU304bM6ou2xsxKFogMNshgI9bGCPnLuHHjzno1qjS
edadLuI1V1wMNXttWI/5NAQl+WWprq9tEWMAHYb4ImVYgfFxX8COfjyxLlv/4MUytiLj+kUOBL9+
/Q4gHxqhhfI09GMS2QPZXTNS8klFEWtB7AuoV4uQks4ZjQwggjS2mRD+f5gyxyHb/6vIwF8XHIta
muN9vlu81cci5EAJKUnFVJVmwGO3CeqCZT/rc2ozS4LuzkL+bGuUlnak0RlG3wCsryo7CXYJIzkl
CM3UfH+pLyExL+AURyaGPE5Lx/9rnL4P1voCd6P0Guf7CsGnrWeutoBuFoWdlPvXNCriWi+4aDRs
wGvvSeiZbLLJrhjgY741e+dfUWkJHjCKWHAZCoqdfNhkxLtLneXuyp5kFi1K7qnze0kNFm5xURtY
qe8hzOIHB9hqIN84Yl6Q0fE8ICivtz3ByaeghLYd2lPMBL6MxTKElG3CaKafzb4nYHZNs2z9qxiK
iAD+62Rd8LU5QuhsD+sghWx+Irj+QKlpw6dt495GUAaPgBjzx1Ckvg6HEIleNJxpXanYHL4BdlzL
FOPt26961mL1tyBgMbirp+YZpet5yr3xO4c3CRyFc5hCEor9YaC/aEazh7GB1NElDJmNi+vXjpS6
U/wR95/Icex30gwnK1R3wPf89hedcYbP0pOapYfQkxRZChPhfXmATltgQILw7nkxW/VbNa7qJ1uX
OJ/MxY9XVc9urbqQ++yJAuKi2XoLxJ20Wpb9Oolxnar+tL8DUHCdxZl2NSCzC0eWLhh+hhtceEnf
vkK+8fSviza6X1kizjrgUdPvWeavTI7s/YKPxW8Dz8TJxaTZvkBn9UMBAEDAGG+H7KIEz/E6Qb3+
L6i1D4/lu988w8DlnkV1VykGqiOzMNrgdXqhDQScNYnWOattnrXB1AZSs/heaXH7Ca64cYw3+42o
kSPF38Z5GuHFaidVVrRr244HhrqADTiNiiC3JCzRwphK3KsNZIoNCRgTJrd16X5r7QVfIRtimd+l
nx37lY92us76hpHT6POSxBTVWlYdzWR9WFRHqSLkRG/+QQLIHFe0JA7wRN6fSmwybNcSL9kGxvxr
SRWKQnPyn9aGxTo+h8XWhCkFbxFn+WPkcys1Ooch2meH02VpTm95/ddLkXz8/mGjEU+1+9iT2Dlr
NJTvEipAcT6Hy3AeTTzlWR0YxMoCfjNzVM+OZYfoGZVGnm2VCswFYK2jdFjdO3ThD70F2FdXTp/K
LondVLOvmWcuSjaL0pzT5Jw/Yd6IbgtzLcU5jdNzbRIueU+XNHsmJnlsXlXZ6ez73dv3gtlOyC5w
cu3hd1LMzWx4LbbpFco7/zvRHYDoxXeopsGRYTBzOndRljtGEfIQWZZeWlnFy0iuURlUR7TUrW6h
ec/kgOUbXFgmis6pK/atAfouO94EzEcf4xJQac0JTWc9vJ2O1SIKzBV3vS8bBFyZOqjd/0AJ/35e
cGuKB5BWXErwPMnWo10WZtA9kBE/bVR42fvGVpLeILBaVxstwJdNqcGjIglzsvpFrtaX4kuzT4Xs
AMOQYOMfsz1YDTLL9fjts0ywYqm3Y/vhkgmJfNMCFGyPktwdK8GieUCxCjWGlkfyfTkUIqVV+Iha
uXAkd5DzQOKBUq75T2x5vjNrG/NBcsZAUzwdCTGWTi5IVFH7i805De/AAAMPoKiMURSNstMjb+/l
B3l8NJRP82mkrSyP04L/mJ0dMJ4/mFhjfHwkztak45+kC/vSl4pHV+U0G+Rl22BAkfbZkUH9zuzd
yezFwClxMrYd7aGhZ1s7rO8Er+TNNirSXaNE1gkuluFcu8WTHnrQWP3YQAqw7fmRKmnn8rTuIus3
YFWE6MMYNJWF1JNnK/JsQ4iYVsuGlKOC76o7wVbvc5HJN2EgnbE9Z5Zc/svKZAB6MUmwNVD63cY/
XKsSyoskAgE15VDIfe+U1OhVACIP3KIajFfRqpO9RwotvyrIvsI0vZi3yhAuAOgrTlnNNrYYEuz4
q4DOBXlysLq44pw/wtXzprVPGxB4z2S+Ff7Ir1HpxTKO0Pvb4nnYf9JyUnCyQ5J6hp8/E5u2nASn
FhjKQhaIWqOqGHqD00aGj98mse4fW6Kvk+mIRAdmB2ftoMNn/pMDkBucYQ8T1JYJw6zKl2kaD8JC
xIKds7tYi4rtpnqTeqLgrrTpaTUjS2jjOdmgaUGSILqwCHbU3zD0BPJ3nd+UwmbUhrWuQTqpgjXM
dk3UQjOR4fksfys94AhvqYEBRvLMtsdJAFNyD08HdSv2+/G3+KHafuKo1eR+esuf5lupM8dsFOEr
EG6msg63Y2eVSBsywdPVU9hbZxKAqoDN/VNLVY4Hyu8u9gxmBsfr3pce0HbFd/oaemP12kdaov2v
Houp2NSZVcQMHhLjfqdidfWUMBLszwhvNJHFt0xAAHgRhPixzEkv9hTaBlRxKIbqPEvXqMqKj1/1
XF9iOhCrjLeT1AblaOf2lDuq7sn1GIk4DqYDA4XP+jbuC5In0uPN8lkY8L9zRCW9IYxkDALgfGqo
F6FWUHjiMqqQcGolbYp4UhqSy57BUVu6LsD25fs1XujHoL+0Hr76CUqjwzoOfTL9sh/wNuMcZrkx
9RJGDJ8hpxpAEgCWSeQ02n8dwpqWcYA8POdsNSOCJUe+50gRJaWI71Aj5Mdxb17VS2OKhenO7prw
A7rknDVk2c+E/X++QkJySXSU/pvYH063DpvRQ3fIvVfV3TRVBWurhBCTvtnS5KOPi7rfaMs6Xgrk
jwurtgeg8V0HYTZ4cwdkYamjAeofT4UVMPrJDc+Jfz6xs+tCRwNcryABDpTd5oyqh+FkfPPJtv2D
nudZzjjGPnOoGVpF8+++7X0afFj2SpSidsf9bs9KwV8ceH5/h69zJ1KPe6ykYRWT8uh5sVC/JQIw
KjcI3wmgGznGzVceT17tUdgI5iqAiHitz0OP3ljLIpCtIDmW8+5ZzFY/vvuUNXFTFk9m/hccGKU7
PB7S/j4dUz5TBD+//5e88gBcOeJ64KgomHl4pF7OdxFHR/zkgojUADRT38gxagPHk65fhRlpsnQb
iHmEadHCsBcnYcPrKBRKaBj2OyyidgfnJDyh5aoliqJcHN/vuZn9PojEED1d82VR+UmjQPCTWLOo
WZzeClJZlYcpPCc2UrAdAasfmRehv/wHKkXjGQHJoUtHLluFjjyBGXWFqKwSVua9volrNkmjy7ju
QsxWWJv9thOnIb9GFjyPbBWptMtnkmmvw8YQWhV3wWGmuUZ0ThO2JiT4/MqFk7sTp6gzDnSJH9P8
ws7L/Y/IhxWNx48QQoBe/ASLMqL3iKHUv/Few7E+Drlv7RSeqTOTMp686s7qt0Gqi2y1O5qeiVfl
q2H+rGUFVrOm3R6D3hAYisha08T2/hjPGsn/IZIgnNwHAVPxpSp5L2CM5ThJm9eF/0taPVookcyv
vzwnXDgz+i9i29/GrShE7GUr6Y7hMofTKQ0VsVMa2IS2+hy+kvkH+Jz+4znp9vJ7m2UwLJauXmvV
cNW24ZP9PALqZu71z8sV4Ihv33BfmMM5sPwrqfAXSuNzx/R9VGBzWAguZlEjTejTtJQwfa+C/RIu
T+mhlKCZQDozpPgJ/14YuRdTeu0krJKh0PdgMrzELvJdbr2wAB9De/gPVzQcHgMHffC9LlPP1xez
3L8w2QyuMDOxvxSzivrbTtYPZA8ftOirlP3ulN/isJ7lH/sVsn0Ei0mWfcsDXk/0ReyneuylQhXb
Kt3tZ96Q76ZBFiEDglpIMKwbxhQtTGVU0mKJd11PBhYkvKvWYLdYLZhc39D+1GLzvjdaBIwpJN/z
XrPKokpBgrn//iCMlnBELKyJ9+H3kt970HlWqDwiH9sD/G3/p1KiCYTLMuymnltjJ6Fz/0pPyGKD
yGqBeQSTEiv8xqgNVfOtKXsgDXha57R7uT6+CZwsXklGIKUHDBQlU8a3fxskz3BZskWozuMiDpJl
I4L7Gbv4beXlSNUsfV1xtN24jHsSS8lwv90+aKEDc91Tg+QyT5YJmTqdiGo/uJfwoNPaNhVsR+8B
9BWBjOEaxqudJ3/EFG9Jjn/G2Ui/hR6JMgrcTxx0MU3FjE3+IjTOPL5yYV0bNt3tNBh0NF3QgEnq
CbQcxyF5RVbXAArCdGwphXgFnXUXL7fUsVgppZxVS+nEQM0ZOmdhEBB5RiJONUz9nzRyagJvn+4S
QLbqVzbrNJa35R8W+lwBMdaa7StZDVJpBcZcYW0im9h44ocmeDMbkrfKw4D/Aw0/OYUHVBIamAjX
TFPL0hEp8hzYYqbwNki2XothHh+edjBBWxkG/86R4DZaEaq1Ph6uU36gkXJyhxHtRyyB0hzTUTCo
UStt88tRp3QtCLB0yxkDGcA1VMRKsGkt0BzVIxJrsivkJjN/mMflukCLdC3RI5ox6Mup7ciaqhVm
gFbtEjcVIKRiamZDPl4NINw1NhQivWktaUqk8c61/ILG7O5fOv7o3S9CquICo/+mZl0/y0KPRtqX
bOjkNjS1DKioMJt10A++Aalx+wt0jhow/UoP6gERQw5jOAYE6E2DVVnWRZASs0iRBheiEYJDOVNy
NUoMpY5Ow5PbKcnAyjfuqsfkLYTTQ9+Di8fNujF/VmLwtcG6k84UWg+3hJEwEo4g41R6pZgUHxNB
eyn5fNwnTiNarfhNhPsQjcdJ0YyQ44+T1cUTDCO1/9sclRcZLuSHm0/MB0KIaEg7vsympEv4+WKt
Y1dU+b45/+pOwj/MpHWBbb0t30CgzVjtTSqQjaAsZVwNaCnKFEEYTZ/gOQdDpwvi95y8auwiRgoj
tLfnvb/laUThlIIdft2kjcI6YzY+L+BA1Y01tck9SiXzVJv+8uxDIBH9uaMlWzGUNlqnwmQhSn+i
M2dQtyxVn+P4CJeh8rLp42qjWQIEyCaVfgzFO+DnnT3HSlP/Fic2FrdCnGXHHO/EuLaWPp51Di0T
kf7Y4xr0VWVUsewHbL4sxeiagYjrk1STVk7iDo7G2hfzX5GNRWJ12KZPozLYo6g4Fa0JATVRaOpe
QrfSoGh01j3DzW4xbBbmvCocYXNEly/yr+V7wpNWZHf5KMEsS+/Pe+7eT29UTUKuMGIu/T1jJWyZ
GhamyN+IfFKXauvGF4SWCQLdG42xJCainD70GR15ziU130TR/e4j4ZvRoxLrnAPP8RN4ObnqrwsC
s/LolQACr7PLPN7Tvwx0hwxpDhxlerOO/PS1mu62ZvKfiJkiQ9CNloxt87330eV/VGtPOcFdGUD/
yJrWXvBPqm+tcKQaTSAvgKU/mbnmsSj8i9f2qKmfv3POwH0tv7AtdD5uFH6w98W5I37+ujlyIEGI
JfZe4IhDwvDiOv5eSCx90Jiml8LCZ95j0oSzzVqSqieVmbXMbxc1buwNLYh6rOeTiL+xy37HDjEo
jBv6nw8gnawrRuycSAHFguo256661a2TjwZeNRfowHLu3jLmnNT90ZbqnYTwnLXOUWtnnorW7oha
/U4VPSm2CFpdumhQ6JZL+2h2xJOWZ/VLDGthNiM4snzLxq+n3ZPTZ/HAto2D3aaLBCg2JUde9c97
gMlxFFysgQ2dBuazo9d9sJiT8Rys/upDIM8zAmxe+pvF9p4qCw/UUR6Qu8I9MlKGd0/N9WNZ4v3s
As0ppr6tn6g3Axvevq4Sxw5YrUdHYrZ4JGNpRdaQc8QFvlr/Jlth5JtWoIjMSZLfPIm12Ypcazth
AdE/gV6pRV7tg6dbU0uCsd4mvtH3UZEwqCTciFvGxC1sMpzwuDRrdbKBob1goNjlZeucUXCDZFkG
54sUCsIpxnki3kimBGrRCltrD20DVAfA5Vil1qzRZI2/RrW916TssZT5AdtX+FSFcDA+aj4Roriv
RYxYQrKtcw5kgt2q0BMfAqItn6AH4WJBPfYk9ZGNb07eRSm8ZLgJ/JCRtoSvKnk+RMAiwkaXzrIa
woWQIUUKCJO7XCCTk8E0jR+AmtCUlZgIqO7NKI8zewusGnhKP0oH95f09k62bD/uMLOhUi6373S/
TXgfDYgtcG5vYIInQclJr4HmKp8oOLSbowH6BGjFBSPdpMMrevviP1Rikw5L1RJ+PlKdahs7uheo
aRFVTY5hxEWWWXNcf6WcXs1Ly+GP+eW2mBUG3yivoAm65TPesS3SO6Ummah8XLOstyTiAkR6crxr
A49K1G+L9arqn0IXBra60rvmmlAYy6LhwQTnQ6uEW6mgMpTfZ4ehht/zTuMvaT9uTx0QKsi6EQW/
SDrnmgsXED3XdFdaGceKdAA6odNq5g46u1x1FoiJvGKhGAl424i6RxklrurT9LGkZYK3XVedTVqU
5JfbR8plNfK8tBXEYW6eJjUar+GdJAnScSuFLw+Kb19yXi5O8QJg7zfnG8Cek0ry2paePj/WNEXB
RRtMmImLNWFxeDFRIl4VfcURhduZI6ye0wVnmuc4Vo4ZDEb8me6EcLSyMYA9I8DsO56PBCWZ079B
fUBljAPyUL3HVQDKfOQAXlgS41sVRXAN566iNnL0sYh4538Y5ahQEylfWLFo6LvD9unBPG+Y40SP
6zmq+GZJ9U6/zEkK08hbKzcDuWCo6R6feyJBjcRG8RUrkD49l0Z6odgmzQGnfJlM7XDLhXb0Z5NU
EP8of83zvkXgbSlZILN1TYj4cImgxhgntUR4HYvcwcZjCEj6KnXgwOKSI38zO539VSGfZHli1fvP
LYdeAD8Nn+c4mcy//Az7dJ+bAALhIEzcFXiLzJzbI5EAKIPBYL8vRV3I7PabtRMiw84cpWuGNOoC
Mq5FRSeNP8uhzCY7/J1IT/cvt8nrfBTFG73LQpwE4tC82eAwDPteo/FopMaLIa/9H6xIZZvmfQ2B
jV9J4gSyuzIPFks3DksuG2XjNvrUqtZMwzraqBUnS2hRYOXvwVhXkirV0kVFgPWnxqSpzcnr4Zxs
opiXDbGn0xCwQrZu98DLJWf6zm/4r6PkyNEwPpUBa3dUPxUfbHKzCta31vPnv1EolcPLSP50KWBI
r+EGnEJDD0q5c6BMFfBH5J7j1M68qNAtCE8qbH/LmMlGssW3YpjC1Bp4Fm88aB+6LYyqOFXXSIHG
Fs3TAzl09sxcSBag66R+iq92OjCuJ+Y+xjqhQM+c5Lrv+aZWiyeBZWDQbXVVUJDSevgASYfkQqPU
3bnv92wo6cgnoED2Ag3WuH/dKPd1K9IUnNghdxghVJucWcTZSnFWhwtE3W7ZtvRLOrM0a/leRkLv
JXkY2d6waGqCclIbb5YpPwVRN8WnWRUbXo866h3ccNPScpE79kwvwYaJ+tkK891kvwoiaFgSPXx3
L7ksaZd6US6H1YXF5VN1e9Oef4RKKQ0A6gbzEuFeaM/C5VqH2V4g2hCaNwO/JmE7VgbisiwOQyL/
g1ezXKgiqLghuEznzyfFvzaOtK65g2hdVutAsMjiKyJOqyBmviH58pTxxLNnSRUHxFVrnA+zwJFN
HIGOpRzZ4FgU2QEFpE4ZUON3ShYbMBd3C5eNMYpS2xfQBzm486GuruAKuOS1ErLiZ5kCNRum/0ZV
B+b6vai3kXJTvOLpJCEXdkcgz3qpmqavy5TbwDKBUHVo18PRlYX8RzboKvS3eqYaMHqh64EAITbG
GRkXdFC/LucP5NZrXwashvmcV3KVbQBEZP2jRXy6qMTm1hsZei2gyOYK2fQUcca8lvpprj7CW9l5
KpGlYWYIFh/HTt4HYq9cvd0ZvZ9DlfUlGihJYseK3jLbWC3Mv9CUxH4JurM+fBfkJ0fCzcd3V0iY
0u2JyZXfLVDms/v2KraXneCbW7ZH69b4pc+Vw2CwFEA3IM6ANvCn7hCZ1VHyLhRYLO6FI+42o4G2
Gwk7chQcfsjQItTbq2KGxP9RXKlNhslSpTxDXIZ8+py8yhm6PgFmhLix0R/cMLGEraZOap5L+Aw6
BWahI4IE0SHk6JwoY9j8NplxJOf3gJdzI7197KhxcBmQp0bWpxNb1SDUcwYzdzW+FVw6KB1d8+z/
LVuCFSLOVNiqOxxqqLdxAsnAhv2XbabpPPRS5MK60pd+luX8EWDJjS6n0sOJkFznZEmLqw2A02F/
oQgWyJqMILl9EeQsWUfnRHyZVBIpr6RFGeYYIhP3dBbkYzOtFZMDZlAji9PcGIAeOcP8HC1WHsE3
vFKDxECPJKKcMqd5c0uElvKThczw/oQVeGAIzZhIdPMuDB4L9piQFDTTmeuQTQi2eqyGXA7mP/3G
Rv4uXCGFWDjTcN18SbWA89L4MRTXYmsvhJTZh5sAjdC0I0lUdJSnyUwHJ1xsHLEvujIZ/p3ogYKh
XcKSp0RPoAHvi/OHO2U326aAcNk8Ibay1aDMjZYDkq7d9wK60rFH5fT0wIDeqieFKvl+O+5OE/D7
5E4KcaFon5aX/3n+6/MwUokjy+zjSZizMa8nhGQgXg+oMe5GhkmOh5vMmiHmDIQKerch2qSRjE02
AV/ipduNQ+GjTZm7rOO/OfVJGp/QD6Xr9CNnY/JzPcGLG57rTA7FPeOsRlQnwn4oPBUOYokjc8KG
PB3Mb1LBr0ItORYk7JPCvX/ulE8yKeJq1eTHbuZn4RmuWLfYCGlGPFhqq0IZ7T6TylMRWk/1WKfm
hQyp+Ubf3O1XRtnk71V4ojFaMJ/DYKMw+t4PdiNaBFmtGoJbPkQCL+ygG+rxxQfkki+nwyt4479S
+nMiYxU67l7jTarYCEUo5ufiNexl06bZUv4lgf7ze2PheMBTwtYZRIW3jTCvgJNdPGfw9eEaoDb3
MRCCgj+5GgSZ1aqMtjsTU3Xi6yBRUVm0X4NJL2naDqEclehkRRqSBtfi7mdrO37WqWD8rTNLGDdb
77UaBifXgBg1XX0tbHedufpnOCMbLHr2THb39hf0+hLnf7yQY7gd+CpUS0wUUW10C0WBnGvpCOpw
99R6A9LOUHIY6XtQx7XQVa5HQ82iOKZl4cvvXUAvOQx2rstpdXONUYJ0JWCnwmx9iQseDAhAYTUm
mfa/dNsDj1TyyY/xfCojRkdfcVG/x5NzatQjlrqR4qOvIX/tIXCFl42SnX00mcjCh6SyYxzF0QZs
LpiuQgVj/ap0SvzUBv2xNGQ4TB7IDmXfvOlz1I62/4FJZIhHKx9SShMaDcHCW+0cObcxt2O+Km9s
NZpSOOMFGBo5hCv9WmazyK8CNVJFjwdgJ2j+c+2VDiNr0vTDR0DssrG4eMWX5Sqi7adcnPXYpXbt
sbrw4OMihgBDUZZXjZjS7cUPdvSdX0frxqn2BdEF49CnWX+2S2RL4WE4HJ/LeNgs84ILhR3LB3SD
j/KEJf7CS/G9HgRKur0ElL66iE3n4jnhVtaGgekTYgaOBD2uexzeIOvXcxPkrFGRaUoHUukER/LS
AnRbFwhjL6rP6BtFf9wtT0ojDHXHItBiJd4KRNr2eJT47hYxZ0fyHiyYVnl9BcALArCnSEdUEuuY
/GUYZ4sMoiWfGSGxG6I/CazPnkeclR+b85ce6wAFujvjO2hMwrt6yj0ZYqVOWvq8bPma32WcLjAu
ehDp/9ufI7RSGdtJuMLv2nn167FpTv7lygpll1jmb7lcv3YlcEUky7kQyjZl4wZT6xO2UmJPHNSj
19wGtucpQOLR5L3jo2FyYpGsNjyhrsEMU93IvPrcsCFhowjPbfl1WKWS55WzY7LIy0cLgqTJpIlj
Heky2BTyqA1/gRaX3gMG5D/7Z1pzgBCjn5ta/bsOIkEoE+dF4JQ/3Tavp31X5WSxgR2kVsNLpxyx
GzNt8fSme9MVrJAjMdtl+OTvIf72MUouO2s2PU8MKRJrG0O1SMhfoVX8DHU3nnV3ynW2c4qDx6U8
tKkK3vYZEvPoeA+R+4tDrjOIENIv9bV1ovZVXGHvg1mhvjwOZaXkLliNgK6LZCsidFI+TZtoR3oM
1Qt7Sm6W+EmF+4K16A6qHBvQojm9qP/zI/TzQisL4ZtKYLCRCUpbEZs5j/lpJCOXX+xuJCn2e3ZK
RNvieMwYPi859UlpqtrGmTkv9m1GEXD89h73/U6etNVpc8/Rwht0FhFjgddyno2X3TXyuLE9PSXC
6Awflv8ZufTcBqJjnXTrv/mS8cPHF9bnLWgFYkJ+pb5LzLpnmi2cCTHMXp9fQ2r1ks5PkyC1TGsR
NiJo+9J5wMo2o8Y6PGjdqlqLVyHmqF+9T2ZZnVOYXbV0C+K6xDdVcgJnX/NBuI0oovtjqi8COMZr
tumqgRHg2N0pIEndNrH8bvlTU5Z0J7TR6sARV3o0Q9qaX+hEMD8YG5HkSCcbvWNafpUN8ebOjBVb
69QhfBM9h5qGXS33yZDAri/qehIklOgmwORR7XQZMcgqKySuNbQkTFQz1c2+dPxKquu56VzKECfn
mKqtpVEFalKpHonwoVcb1qfqtCJDxodvY+XLmhTrwfk2ueZ/eIhFr9fNYGfTCoifpUC216zlKMNT
kkAw0bl50DyoKWXqx7KHe6VtjdurdN/f/6CdqJ4FgA8vM1IHruNEwPRlExFlFueO/yKCDrRHd6sL
sQFKfLe+i320EdkN1oXcGaZ2O9zkRV4AcWe0hLSk2tb32LenuRgQRSpQQhj9Ixl3bTgXCsv+Bqyb
8NmjmKUaSvE7AzonuySK4Ie/5HlmdRun5zneyoJyE5epzc7Ng2IRXoy7frw+G9RgB9YqCMoH4eM9
1gtNqm0oj8+HpogylQh1B9VxtYEDQtv7+nZEZpmOQvv5z+ZU4APx1D1JYAccAH3tlH+QIj/o8X4I
jNDTy/1Z4Eo4pbqb+3JShNGZcoG7gWWDfgKNU/IYd2DIFgjWEluNzjaZumS948EGQ3Wp+HI1jxGD
L9QfEZWFcL3WxPF7oMGNIFBj25tbs3g62jnk+L449cMvlA06SpURGpwI7WX0A+omCHnFVc5Ilqrw
+iMYZMapi5CSKJDn8lOhQRWUPl1gWW4Sq0UODjPADv12KdB15h2snLO2KONugnrBAleUCriRA1lk
ZVGkHzlgNlejvv6Zu8Hgh0u8KhjGp8GEle0uyenGiE/Gp9g5mY6oNVclQEuE1wI/TEqJl9akpzbx
OMe6hZqWjPLNpUGRc81Fwvn81UfAWh8TN6Z0pWv/qMC/gexMexONR18qMHUXrfh5HqkZ5faW5oOW
HGUMOE699vD/y3Tu2sJE88k=
`protect end_protected
