��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjH(�D}�<y�R�S��a�h�����J�iY�m��D�H��v;��ݸ��,$���w��4�-���b	��������|�,+Nëz�k�
<��ǀf奭N��#�|�:��x|�>$_2���e�Mr2#;P�ۋj�3�<��b��kO�L@�n�)<�|e���e#�R�hm HuĘ�;���ƙ��[J%?���|m}�F�52z��N#�/��y���'�A�K�����c�?kb�+�h:ы�wO�IP���yY��q?w0fF�K�,�X\9�%P= ���sL�vV�US�a����gN�d��QM�����n�v��*��}����8����m�/#|U��z{��
I
�:k���m���WLDP�%����AEeb|Z%W{gFw���9Ev>�Lt49ʡ�$�����{uV.�U�EG���LY�������Z����)�#���ꪧ�\�!���ܜS@fD�����f�' M�v� �3����\|޽]��:9k`��Zt%��Q�z�}Ν0E�����dP8d���*VV��&�e���t>���[Ɲ0��E���_���|F��LT�[f���x���;lz�3S{<J�qi�ʓ��d�
$M��!Lp�fʮeָ51��lϮPzQ�w��jWh���]���:i�ރ�1�--PE�/N�X�fW��R$l�]��_�ߝ�&`@'��<��5��}=�{��	ka?����J2��*2��P�9u�T����(�$��QP�	����H��+i�?��ۂ\�Aԓ�ޔHw+H�N���! �1�)�GI���B�&ܤ
��V.5rD�X㟓��y�DX(1L�s=
�O��v�c{k�Jw�I����[ݻm$�iX٭_�7�ϊ.��L��0bf�۸�,�e5�)Y?�P����MhfH	���ԝ�+v�|�.��]�E;*�  ��adib Ԗ�j/����b���~x��:I>�l����Na{r�sf�&4������;P�N�o�%�a�͠�w��hb�l�!�e�˒U���?�ZE��8�O�f�ұ��s5�(XQ��hacB���>x�m�x���1��=�9}�Ӑ�M�����w����4�9��$�6����3F3y?^*��Kc���w&m%.�zۥϊ�:͚7��e�c���-7���s�L�i�+"�o�b����H'����Y���f��̤gޏ�Ti�D�*j��k�}�TV��|W�B�n{�\�ok�[�~4O#	�5������/�0�v]�N�*���{Y�s�N���AO���|��Cc��@j{zِ�M�B�_5�e�<Cxʾᦋ;�<�k���R�v;���s(������F�;~���:=��K,_=��ȯ$c�� ��
�=��&�H�^�t�%�����puZ֔��o����&)J�"MX��,6���u�d��������Ʒ�̂k]���NB�(��s���Xň��xQ�^D&�\�Y*��2��:�c�`��|}���J�p��rhh�頛�5���+�nf��R�s�w�
{�zh������0�>�����vz�h���3Xh^�ƚ@��a��jx�O��)�pG��"܇�}�,)CIh���*+�B�Lu�Q���F��Qv�{�;A
c�m��:�(�A�#�2�6,W�w�פ~�W���ZsZ����.�HY����!~����Ҍ���ܸ��,!"��P��i\���gm��`��#�	��rpe?�8Z��~�N8
m]0��u�������<�x4�(0�/F��࡟��!�b�$�,
�����.f ��AI�N��o!Z#l�Tà�Ԏ,��[ϋ�QZ�[jد�[�
"���
M�;_��I,mKJg�h@���j���g���&.>��_�CR�*��w��6��V�uX�yǼr�̼����!}.��D��[���zy������-�s����q�k�4>�,I�ςVG�k����)C�Ldm��+ʗ2"��
<�5b�I{�ln�$I��yG"� 5��Q��8D Ж�L�)�������ĳ.�C>�U�p�7�B��?5��2���{�;(7�R0ИrDS�>?�/����x^�"��׋�6��țZ?{N�F�eZx+kK�c�r�Tb���VM\Z����s�,Il�<x���&={��1-���+��[clہ:��m�t`c5�/`߁C �����(ey\���� [U�ԦU}�*W9�����E�`[bFL����,bp�u���\ZA�r�ߊ�1��	�j�=T���{{�兢��V\��t��(���6��j��(�y����gK��G���(��;@���)DahW����*�'�vz��S�w��R­N��SV?s�����Э���ϒjt�1�u������bb�z��K/;K n��j�~�𸈦(x�ٯ�����y�j��9�� �e�VDcۛ��E�$��"Ɏ����E��LY�bc_D��'�z�e�L\������T�9��6�����^