-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i/abaTA2yOs5a/cs48imOTLqUHAK2KZgELyFITh3Lrdt42vlKUApxBcDZoQ6+hWktVsfgSNIsa2p
GuB9N29cjfRYHyBzQnHzRJU6O1WJZgUjrchSUAvrJegTfEEu4Yj3kRgBF7DsqMYzSS5MwKPk0OvM
sfrrMtgFhxR/+c+Cn+Iw3hWp6DvgjYImUnPbHLy4HDvlBXrQj2Jq7YWC1/FU86J0jwNnsSkDhbJb
0KnFDPBE8WkwTt3958reebP/5/+/UggxmnUzeV38Czvdn0bpG3TPmIhXVuGm8+h0v15dKd9OEsJg
aJhqjUktKz/yjYMx0P3OZ9cKCT6yMo55tXHPzg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
AKN3dg0EKhsPw4m5NpqH9JmFhlrR7CrQ1PTPP3HdnktqP4EXlQWPtgUhcuqnnSQBNsG/RL++rPL2
OKrhWeAMp3ASOUTORpYe1+plw5sRdOdG+nIFfLLAbhZ+iUGMAgU8T56HLBi1sdg06Adn62Pf9sIo
ztjZJGowQj7f2diBuZXW+1ZVVCYDM5x5l2NTduyj8ujp7qo1eZGWj+F+TnyjRmchankTajwslLrx
oc04z1YKFJfgw/HnpYhUiXRozeAihJE0p+NvNFRTstnO8DPxyDL0RfrrTA0KSGuhZQyA0yu9o5L1
saWbgLBD0rzjouUaMqS9Zdu2vBP9SAD9clBklkkHl+iRiUoQHrHXGa4gQMnPDEH7dCXLmNk0f7WK
zdMXwvh/wK0DCzFa3SPxIpREE4V+qvo0RB/SkFdG4u22qnvomWfCzsT+HRwul10ZGO95Tzk0lar+
TWY+dcxCJPpUqZ7qA5b5ws5uJ57aOzC1myvUyCTFpNp2oN3HdR11LeUI0pLYbH7DNKF1y1g6zM4R
gjuXwx+9HuwtQmQTu+ZzmMP6ivYI33/DU5qjS7RCKjRDLEuMiOPoGrrVY6m11Q7JszU1SE4xkakI
RZwa+o60ZhEYp78YQcFyTfa/6kmt0QThZYUb57+P6TGDEcilRTeRzeQEijvTJmNun6UNpHn1NqVD
GzxqSU/tm1Z4DBnU7AJJ/Or+aacOyk5/WKIQ5ABnkFptoPMvWhXNpi4E4P+kLEXF+nGgLp5lYJrJ
pD6uF/FeZnX6HXJvEM7aCfNYzhtJjOVo4NBeGiGiKcVGGgkC0hxQToXEsupleu9Ms3flS/o6Nmfw
PHCIKKcklKgEK7IIuBKkzI1XChxkotu2COKcNLdvqeUkDs3diQKHerWs1mfO9wXTvOEIT4grjWdP
fcq7ZrsLma/Y3CBfTk7Jg+f0rGCBe0LDLK39CpfXkXNmgpXjyabtXBrPh/6DBujfwBN8h8yOYxjx
bniY9aWq3W0+sQge5BneD5G4CJCzPj0BvYeOCl25F9N5lf2zYUX+sy5O9w4yS3cFE2k3og5+nxS0
ihS5as2YmIbC4oqlzGWcKawkI//tEeGAqknFZput9C5JC9BbKBlX+9aHsMu56k1gsGiehekopRWE
S805oJmJyqkkhJJzB6Zk18WDIn/HsxQqG6fGyFYqbjIlLv1eqnSG/25IyyarcmQzy1tD4VbVcT5f
vwM8o7yQvPj5FOboNYAKabOGqmuJnEmllkpNKITNjhLha9GjI9vuroyZSsNNVcRQ4LLgr1vgbQIS
roXIzUN2zEEQ9rPZSAkUDwnIkbsOoi/Q1wCQKFfoWJ8xgog5RfKXp+JnPTbrACw4MHvEH6ljgZSr
RfhmH11PwW8W82K1uom34IWRJ585SWhbsVR3n22JX8Yat8RzYHY2j/6MllmtqlEzuHE1Cz00GfBi
aolkOPtkP7D4pfekNKtTNv/f11DsLDlaarYjUPurA5GsyTwAa1+QnGNLkjKU1kZgRLxpPhpOfFPu
ZT9mSgoSU4x4J8a+s0VAe9dq9dqDjRIONhdC0MQxzU8iIU7H7TWa15HClHl1z6wNw1StXjs3ngu2
jh7NK+9ELDv6jjrIQDYk7pzEWKFRHw8wGADRU0OCq1b3OqkglO4AlCe3VbA+tr2VWl9lUUtYWJTV
2sjzMxhcg0mFQmspyKoCuR16mTkoecE1C3V7EMtO2kSxTjZz0jci2/poyW84CSoi8pgk/WxP8QfE
8pDXDVjOIjvSFo8HTe8cbS57zle3rzLW/C9neUEGqrU6ofjNvn3QuGeXNO9F1SLWgyj0sLdeVz9+
E8J9HKtBiOOk7DKaS490BHt1oB6WSAy7/jeWrATGfrmCw4TlijRSICz1Bgjy+tKPfpNa2pxlgZDL
MBH2U5gI7aV3w7ZNY2GLfO3/8QiecNexsEWEXMVxUD6qUE1ouAXAe4uazWjgjOFKgbX4o/JVZ4g1
0pIdZSs5T66ObzyIw8F0NG6X4yvnRt3uO/+/c56VCY+oALkyaL4KoS0p2WPwMMN91TG3pdfhfB6e
/pvj8/nGTpkpMFe8M1tKVz0UrufFDHjPvEY849nxh2PxescY38xJjM33ile4n6aGshR1t15vNUCG
fTXWpWCOd2LMG10P2INtfMDRbcOZoAAwXWXNUHcAyDZVjAMnaYQMt4kFXWQJuTavBEybIBvzP3v8
LSACi/cCOU2IKhGmUv1O4NV4bIDopzcN5grXhlLpPqYpdv3u85aPTJZqLYehh6Ki8SSFrEVIWbD8
Es/uMy/M9Ni2Mm2LXFLJKrxHmNKwPUxxh/TVXSFVKC8kmB0ShdloUYJ1ZhYa2hahSeUCkMmbkmt/
SHJ4HhqiKUOSdjt8lP0avRJVGxki0bvWyz9LdcM4SZb/NFEtQjv5CJqz+dEd7ssVVYRJiTnFVe8V
KziNeAVDjj9GFzSatdZ59WWy2fJ5etIQMr4e6cpUhP6/UX6KTanKXEq+ZjQAvDWSeJ7k8kyKBGHM
CX2YdfK2p6D1adpZWUlBaMEROjFWYpR+pRJ8LXapabwPSjuwxZBKMGhUFAHTFNrPjpa6A3KXpjrT
QowE0D2QlhEj1kfl1zKn9GnUE/vVbD9606uDM7LlnWqhIHvVJr1s4bCZ+ibz+Y1ekTpUXz0xWG0e
Q0JHbejd+keMQkWxb879mkvcVpPpfs0CYgZk3Oc3239nC3h6y4ALbqd1GmPd2Hj2nIarO3x1BEry
GN65EMeYLYNw/GtHYxXVNKcxgZ7aCJJ087FrQrX437CTlBchZtg2vFn5MI9UTx0TaJ3bE+qt9bow
bnA4A+i2qF/2bUGABjrZzJoHyqpzhh0FLbS0yc3FjuzI+joOm+7LTysRqRplf3VNuqS0q6aSwxrw
GzbBP/alYmg1ZbWll9A/41FnqwefksBp3N0F3fSo9GTt1KWE48Kv4omMgg7kbiaKjHOZ5mhKsZNE
yS1ZzGgQNDIL6Nb3aZySveSrBmbeoYBPQT2uit8JuwB0pqIOtLdFN2h4dHjQakkDGbo5Li02M4gE
0OzeCYI/4jmtJsWXViYvFpZQ8s5qs29fVd+zTOSt70TPdUymb4EZbDHq7ucsaeFOHGsWinZ6cnjY
deIimEc2TljDR3b9rSnwpV6FCUa7Uvaln3kUQ6Wa8oDCCDXHQypMREjmvZh5Tzowxr/jkVobHLOd
AUVw8jfWEn6sA6qx7VZ9SN7/CYJo/JbQm01nMRFIAJsD/862vqTmCDVzBMPXVtlXOrqXjRSDNTzU
2LWO9ylC2WE7N33LnrABEbXXKJwBfecMIP09gDueEmyfDInnrFS5B4hcCJRicJW+5+f/CTEbhtH5
+nqgW8yx7n+maLPJe1GL/b5A58uwUvOSPthMGVV8i6izSxGP15rBmnx1KlTs0KdiWGnfFlPL5xxG
9HNMEgulPjuQgPmOrwky/OZQkod0IHiqkKUVE6+5Mq92RKGwI4HL7c54kdRi6QWcDrXvQnpitUtB
Q2+9CAGRSDu2JdAvTNUDgCneqPkQiser9aQLXnYsZp4DRyRT8IDrVzWk7r9sqIh7oIeywZc1gpIY
LHvQcl+nYduwyruFCgBC6ByKUCnFjqnPKyhHIG+6ul9c02Geo61mRntBatbiINlZCtRmZrhoiCVO
9H3tjSnPTkcGivUemX8Q/rZU7d+UK0Oj1KVbyOwainipiiWzLqOMkeXS0h9ZU3v1xPl0IPzqWnUl
w41F1y8oThh4Q9uJZ8HW95ZY1/Yu6HaxyzAmtl86TTF4uVvSiY4EoX2gIDlVMna0xNMjssqwvp0p
Di0csdnwyyKTK4zhIlPNVvU4UndZ1AAKkD8GTNLVeTkOkIdO5Bc68TIQ6y0t6oXxvdjd0lV2+4NC
eI9DocCZwQWFhmLpGHgWo/EvXOXMBzBesmoQ15NDOKi51Ie5dJFborOvTUYuxkLk/wGj/dRxK0Sv
BQUW40yajRN/enUJwdh194HzKev9oXJKgSS403Lkbyq/zbBWEexbh/fvufHRhLpYoWzpFqpW0F88
nz+sxzCWtpcVRqkoqlPk/0TpfKy7XBnyLoywf17UIlCxUZEDiaGWetpKsozDKetL7PlbKHNQCke2
RPlqQ7GNJuJGmdrs0gTGNRsUwq3sKTRlIar1wPXfxKHBs7AReLtojxPwb5ZDCyCb+iULzmp44ZCH
ttCBfKvvRJpyb2/nNSNuZ4sKXuIO7NM+9p0LnwA0aHk72bHgipSHxI2ItWzcFTH3wUFR7zsvZY1M
/TfZD8shwkXgD7AxbQqyvgUegtBv8rhCH/yx90SxncV/1phq5xkaNWvxpZ6JdNf84T4vhQFNucxz
DqHoaTHOxUTCZFqql/hKEwGXLHWka8/OICUk6CvUGTY+rOOqJCBEEdMb4nU05gbXnojEXReohapg
WyjwlWJ4NKRGeuMjRkqz4IX4r+fmyhjMhpbMndCR2OGGPQ5+hW/Y0fK/cI0ePW+O4F78q/awTL6L
ZfuGgbVSTNogXBHEjUPq8jDjcRlmWU/oXxNkQvfwzZntyt/1lxjqSuE7XMKrkubYUmVSMV5wnNvt
HA2osIHllU+S9VJgTP2VNwsWxRPnTS0HhA0vayz4PBHN0WMt4G3bAwdtAwg178FfMMTKUe49V6Iu
sAftbzwRcdS5WMIEKaYFPhZnM9dbjIPLi60tspo5iqx4YB2oGhr3+zaw8/+drHF+6SFg9Wuyrzwe
MhVmIeF5LMV8DfXq36hJCO1s7yte9eLQO6BzXIswg0FXcgU3C4ld8Hh4dZXBFDxXI+/Io4/NiEVO
eczik/nIHNfQbxsbHr6qOXADdrbGdbmJG0TDC9IoAWMdOd1kXHUMITrAVDMBvI8stldQhgCBqtev
7O0rus3PaU96U/VpeY/VWVA+F34Q9CAt6cHiQKN4mc41eRP3cqINEVa+O1o9gxdp0hJKbhjmVSkt
+m9eftEZZ7fS+u+kXq6PCf8CPUcOeHyP3gWxb5fFVTxId9qcsrEl6PktKhq7gUQUZttIC+fEYrIm
sF70yBiFYQGCKOTMItyBnhjJ8QDta0Bh2lYFfY7wQJDFlgA3F07/E/wd1SE61YBxfjlL29G1jjBK
jWFTFem18aJiZEyvRazt807OA/w+jg/oB3dAjsNnAfw9Ccl1OA5C+sVx896mbMBo8Yq/krb8R02i
HN1fEFlnvTvSF9ONPux3eUBmc7cRu213Bl563+uDGaDuhBcfkk/31YerN8lWgeAtgYnmOqTXORPS
uWF64QY7lhFNwWLWN//YA115solVh2bU2Xlv1ua5yKFET9xfzUTJ59XJScAOS7OJe2lB1y/GvaaP
50hqPTUw1bVuwwThdG8wY9RjUT9b2oGZlcsCdZSBVvUaay4YvimvT4R0Bo8DpRYdT1PPIZIXdoW0
dew4qHUGkr2PANfbw3GAk15esAgHMdhG/O8a9KVUXCiIfwDBX/Qyf7JKJH04CsKVFi32Diwqi7rs
aL7hLU2uHFCNPPIvuYhCWlv6hy2qvq0R3DBxKZSwyUAJOZI7VjrLhQ8+13BDXHKd5GraCilJtvy6
+Hr51T5yeFN7G4zoBhhTpEQTTghMRPVm2ElMqsbMnY4/Ocmjcpc849pDVQqwwuhij/st86uqy0Jl
5e24XfDw48hAhEJemE+KcaNkO42doEWCZxHA85E/DBH5nn4L2FphFT9fC04b16zZVPw9OkCYtPXV
1nt4mKFIpfyFVt6F/CSC79KK0XMcBhztCamgJQS/U26leCu8NKEmdA5OfNDqDBLr86Jpt8wPkCzK
hTU2Z5mc2bkcP8PHuvZjryo+E8UsUm6xvHo4CM87Om2c7ZSf6xuAVwS0ZdwIc/K3L70cxjXaJDe+
fUfVUe2rm+HpTUVZ7jQ59RMAKEthiiDqDIJE8qzunBszy0YytZqZpwFvcxw+DFM/EZScvkY/jjh7
ezA3AMVUL3HlIl2YANMBD4y9Q8WAiwYqjrr1W542Kaq3DBuVj1DuhTbKcV/0lV2QPT0FP9Idk8sB
iYHJdHUahP2pvA4AXRKpjqZXrM0KWe3rIy6mOQQ9jH473v1Yr5prI2zYXNIhKRhaG4dh/on6q/vb
k8wxV//EW6NWUihYm8t7hIReIsAJPrvVEP9L9M2Vt/3rnC6TPBy02KtJAJIBYV24zglN4Tm0PTZA
5xnGBqL7+UZjXKWRt6GWZyHoBsSyClm6pVosOhkZSx0dku8UHWCBVFVm9YLvBkCqDgRRBVcJX6gM
GtcGwqR97pyW7SEShUAD0QaqNnfLew6COV9lCiqO6Mgu+zcjYkd/xEGuqaR6XC3HAAH97X1zAgrJ
c5aHY204PxIwD3IVngGAkYu9Bci/dyPO4eYUyQLJTF1y4d72lCudeh2RWhE3rvpYoQn/C2+rdyvZ
/We+L6R7FpN6j3rA2H/n8qRp8DL8Yg8ysxfR3GN3Yp8rpmwLd9fKQadQRqi/CMM/Fn+uWZ4DdDmr
e7y8Atc30NB5sz6WPC12HO8BTZmtd5nusTpDSFrSaQMaMvKbewrUONhXMhzjdAjCfKz57LTFpvHj
5J76ctDu0k2KFNumbdT739EJzjpBjsyN20BMJdFeWouGoxu5/z6lOxc0E22Hgis1iYQivUr7e0CT
t32qi0hXyD/FOvAx4MazyFMqCX+uaiFPdVvkiLHgX9nVA0ZtOzpHkGSZwaEIISWpWy3o4/p7rlDG
avcDybSjTOOJ4wdj6tV0nGSHpypNHHmQzO5GtlkEcPa7hw+StL0HXrIgbKVzheRYxN7/lAiN7WC5
QaZsfR2A1ba0Mo5dCDXPmDZIcAXGaPrQvgGQjyAzFg+M/JxxniB/+YyMxRxGUQknTeUFpLW2fDhD
3fFisRsS0wdgDF2EaQl4oOB2wPRuo6rUdcFWEF9zrNpRFmcDsnIE+awxdfKiBUvePrXycwYrKLC9
4ESLSnOT1JOuF0IPlu5D29qpgEFfDRWCQ/nRS01rVgHOVKadtGArSaP2sGBAvrFCAWZXVXuh2/TJ
uzGMhWNYuX06ncEs45/u9fO3c5qZWXl8NtI1jsW6A+lFmTkvAkPTiH9jOpZcFxufwzE34u10dxvs
J7iAPBj1JYdovOnpAF69c36IjAtzqqD58Tahw4Gc1Pw75XtgdxPO4R3JuZCf+J5dif8BsWIXVcrB
0qJ0UKMtrylu0dNdzyNWvWqq2KbvXoJAhcQY09l/yeNKH4wB6ROwlOWyhCXR72QHt+iQSldQnGhF
JGf/FX4n4FmUM2k/plwBxC75aIhTB/PRTv0SjiljDxWV9sa+LQz18Xs1E05lA3ZfbFmNKNB2r/DE
9UtHAQb42h/1PELMovHm/vyqem/JetLjjVXHbpKDJ3+CrFuDFIoEtbec96k/Yq+KtCpiCoQBMWAF
JYLWxQL1TYVxbzdA7AamlZibUKerufkzhltilEFVrdL+/hedi5X5bfQfbafrI7bL/4YMkzzYWb2a
JzT2mp5iCgSeky5PHsvs+Ff8JzFLFOrPmKzPaq8rDr3xGrm34VUUzihTVTiqEdbOlEgOk8qh3a27
0U3v2J9PqfM5v1mQjDTMxVcItFlF3csJrrr9ULhxzTBO8E6Lq3yYSvZ/rumuEAbAnbtY5WbXffcw
0OWap3Kjot0LliSzjzJuhJI3waG8lNyLZ7fcC6NGolO3uxhdsjohqUrlKopbYQ4Xw2IQu8c6+E4G
eO1r4PYvJErNKQlT89r1YzO2pxRPnpJG2F0AyMyLzKWCc2/CYRhVl4O+YwuOHipKktuXASo3rR0s
zNmqrcQdZFzYOUx2kmtlqHFZGZOTmRukZ8FhppBdbIOa61POsO3XgL+/33/37X0qzxEv76wH95r9
5qrp6/+CapySOdPGhl6GZSAU5c1t8Qx2MpxKkQEUjE4ofSSRhpMGJD7TJyfafkZb/1nVW3gRNyID
JRkox7GxNU1YKcfWTfSMtkjXNz01O7T2/QWWas7ngyCUxqEnUrFenoQU01yA3kRQJ6kYrGLn5/qM
Jw1jPumLjxfwwMhNF8eKTy7CQllpby+VqGHu7f2sJj+9XwHqFMFLSsWChM9LNC79aRZ+06t2Afb6
q6tVzUw/r3ePdItIQW6DRChR6jAe5Yb7PXJ3PKoIsQgCBJQAMJPjaP1DaT4VEKiYssy6jjEEeXXB
KMiTMsz8cikMlFWDOvuuVbfDf0HkmJMH6+6iR5D/D3lfFNnDcMNvTNUtfmvPxLY53yZDGhK1u3Yq
MCLbEnc2r5PMp7nub39UNA2sM8ic0AIHkR1jTKC/SBbBHC0ih/9MV+tOG4L/P302UIq/GoXgxwvN
6n8OaOVgljszBoJDmHL87UZ4Ni0Q/L2fl71/8gIZRadysiAVGKOuGgAN+MPVDKyFxu5mZy72ZVSM
7iZI95wd0OVyD1Wq6QKMGs6aj47zVQ5MBnX9lvEG/ZIG5CTJzaVJ7dULtNLUrQ+e2Ll/ned5SwrR
Kf3f/7YkV2AH0cJb4DIDbgVcXCem7DdZEbneruYJinqKgkRmlKe1KwNdCOLDLmfy9vprfpz3GByo
zrHbfWijJ9yOkPxuqfev3eDUgDqd0IFUhSjSOvbC2mgGUbtwLmebQRW9mGVKBtIGrwQlC1veZdNE
QNus/BCQaKFpujLm+cCeTTxY7gMNOITnUxECiF2V5+7npCfNt8GGht4pFMBFhKfCUrOJXE396ugS
6+tomzngs2iv8ql+lEsbcU6ZyR2VAMmQtKIFrjZ75/IWKxHxFYucaQ7dUxXMWewxRsrfXNpe47a2
+M6q1CGkjduQCuvUwx1XUHt52BRd4x7q7kFW21WhhpHlA0f+VSlUhN+wMffeFuJgk2n+dPOuowAK
6H8OI6GiEu6VYo2JO6+KxqwrZ2xPNx/TsJNJt/jkGW8WoYxi1KKLt9qNMEmPkgvUtFXC9bqWHNjF
iSU46Ur7/iCee/lZS/KlDRuN0gtlrdrL6rEzsrEZCiPiXwjCOTIpggWQ4Bay4gvZM7wTm/oUl1z0
ObZZHC5O+UiMi5lzAHPfJ339WzzKNo5N+GfpER/ble8o2dAyGSM41pUCgchEFeldhyG2BZ1l2L/p
WktA+s0vE6Bbx2GUa7PwXj6nLG6RqcYqKWaKG80mBYvZJZVzNFaANUlisrJhmzDz+3YpeI19IuwS
YGaxz0NeT6pbpeF3K95yWz9hxe3zh527yUyPCvE/IbFMAJ4lMjqZA9Yp6dQ1hiAnhOaiYBg6Fqob
NCKAHipnmwQGuAN0DmsTraZKm9NqKUK1kOmq13pExMyWX/kSCuUpWmCAT+OcbjHeypfwJqGzXIWv
hxpe1oYSy2i+4I/uTSrUFtOCxJw6Tw8wvMOHYUzj5GfhCT1QV3iKDTxgILOpHupdjaBNlsYjpgeW
EmRVvFD0K31duI6hNl0Gvd++zrRSCUdQ4lScYbTXgaL6gMRfPw9PP0DlTg/WxF125g8TVcEQU0Yb
mhXPzIN3ebnrmUNCXKjKc1zQBcWhZo/NvCoY24mmSjuJeIxJQpTyJWhVL3hTj3aKTrRcut/IA+zf
qdnIflYSQ+VN60KLEDWREO2VQOsUj3DOYAPc5AX0Uw+DLQrkspYFB4EZg7M2jY5Uuxj24+9gusYQ
CHVaXavo3CocR3LSlfn7VAJ8K96myufhObCD8vDZX6tPP0U3ApsRsU4Y5qBjZVMpdCtQOAKcZEde
zBZXIh+DXMUkDwffvwdSNH+2AC8QN21N0MrFB1LtwFazyqmsW7VD1/Ydi3CZLICbkqZq1AGUNLwz
Vkxv1viLfobyVU89EMrv2MJH1+TAXlnWv5PQO05BEbi6+PvepKN3pXU8bs9/orLVAD6fCVxzdDb2
Z8mekJek9bH+kdzx3+Nlw1acuLzesY1XnQH0i2odAYnyeAywqevd84AJQgSGo69WcB3yir5qbHUo
BUwHIt2AoLWGIO/sXG1uZcxC86p7geXo2yO8Picq3zi9SzXZ5iE6ZOcSW14yZ0K4Su83UtqOEPIV
Oy5t9Mm+s9cIY2Wiv/I8DoTyc8RKlARBw7U981dqfNPoKEALXZHxnXufwQ8wtlO4ng72rWtPljRM
7mJEiAwVk1DPwRJszUiIyZxHMEKfsS+qrQPjjSZD0RnID7Sh/Fc25didMaYS9fCpRLXj2JU1a/Sq
hiR6/ntz2M0yUspwiqA7kON4pxuXzKzVwJdHOzxcgIuOUOeVjMDuk3sULtf8CWrJPCOC+JEbwaJc
hNy8iQdTGFbAkUcz4NUVyYS24J0aaWtqa6Rxdn68SunJNH0e4Prk+sXExaX/KSb4DUj/sy7koIn2
ZOwa9WsQ9cPtqzaYgiDIjhtsfdhwkyUe9KLm6zF5ViEO3mWt8GZddIlcRbW/Zr0nhqL2E36XYoIx
gN5ni4fPbmg92Fg3vmjlTsXBCoPlGHZqlkQwndc6XPWfclIcej+QXG4cmhK0CUgJCwuoy5Ln5v6n
0sl9EiHIp50jHMaLm2Dt7Ydb2iZhfYvKFJYY/sdk/ViTaBonsgXE9bTpTHIeSFVA0HPReGqo1gvk
f4p1PF50D5PaEstu9l3zbHKPu3C9J85RMLkXL5/N8R8lU97VG7TyTY4fhiEaVMI22ddb4b56ZoL9
IjSdKEFnQ+21pQOd/+tNNP6NzbXRnEjVqLPOsBaao1fffLlw8ApFBA+u9VHScGb0+QRWFBJM+rwR
lmnPgOiG2H512dkeEULJVcZO4bp5oX1derrRqihPoBvOSv04vexPBI+Ca8oqC4vJyxWbjK6tH5mk
0ZSvbefCowFUwiQl12gb2TnaqMKKrqu70zKn3QLzSgm8fI3V2lYGTqqsQpx4IFaBMWujW/PtLWBS
PG8OuGRRb80ALRjc/TvGaIgzsI4dmSkGPGs0nIjZ8icQfuSlEeyWtj4yw9896QnxXDde/EWSdxlg
KWACqz6XiUola+ct9tuBST7X8eZ2sw/+w8gI/3FuRuI3hFcriMLVVIsWM3kn5sbYDyKzeh7GB3JJ
QA8+Xg6L2qbR7tIyZZLT3OtKQjxx2NDU8mvT04tXWc1hXKkJiYZxJmtNWwMJve6TpKMX1zIEVX84
Hd9Pn+Zsa3Qq3FxUL3/6/DWQf+mji4GM6fcmgdC0OotJPFfpeWfHgaTiJECdJaJ466UV4Gfcw6ot
SgsxtpVzB62NZeQRCA89tv7HhmJP/5/oLkXnyZbSPALoi++hbX29pny1jNgr8lFJm8XVoEpmkwCV
8j4HrxwoPA5/GBBiN6/mCLwIlFWTO+tQKHlDYVSXtrQq8K1djkcPHxyPh6Jsb0Jwo7y5Z7cFp+PS
MlFhkOz6PByyB05PKeOkJx4qYr4AJrbcC+zy5Ko58yPHmvlpNkTD2/mTlQli4IMmIeUBD1vooJrk
+w1tn8pWiEN73yGktCL/tD6n8JWKNVsNeQaFATuA59sZ1Y5J9qH/03xP2NahtEnm9lhhaf4/yCd7
3j7UarGC3KC7zPpmEc/nN8X5e9fOY/ERSzatxIUzif0bFHgbvXWRSohR1yE3vOYNO7mQPfUTP95D
GOt46xp/3wP4B4CsKorQ+JFINUE8SojpVZhgmH+PtCHGyC/lXYP8CR/JBKTqbRzz2EUCrJWo1GKR
+RD01payDTQBy5TkDWlZyQiu1Q4OUaIUO9r4JjuexwsRzH/tdq0kgJHIdxR1IPmtkvz4N3UbuWvJ
p22n/GxrSwjzorJteGHNSroInC3I9PqMigpZ+JHtiWW99wzBIBw9VYCnUj6vPcg00yLy8mP3tjSm
Dsy4dfF9CQM0eRXwlGFhDunEGjCAqAA2nTBb5tJw94BriTDZEXHHZPOgskXc9Yh+lNlsUPyoEQ7j
5C97YKRfju6yH8Le+c6oTDSJMs+5vZ9Nv94yAEv/9FisI5Bm2YNQcsVaZt0E7E8lWqbqMZPYcMet
u1bgSySy46+rSpEw48sF4sSC2vd3Yd0P+TGcEb/5K85IhMruFw6iUapLKDfn0O8jxawRI6tx415J
TyxZMXgQrHRPKzW4xk1qcv5i1Kg8E0261cN5vNtkBdXPn3gJNHVdVqeRZmIa6QttZqjvv6ts1mtr
/qrpZgp+aH9J++m4cZa/LPco1Zf8D8SvpXIOQA4S+mv2H0ZpMnkhoOdnZ93Vcdnm8nu+r537rmG/
+53y42xanu/HLZ4YPUsRTU97Y9bT2yhdKP02r7SYt/2qD0fgBlR1GdmznOUDCr41apcUQSvIzGn/
6Ym6+7tTf0NHlizqr7Zz6ieOD+3pbDk8ob9ZEDppnJNxCDBAbUniqe4Mz+R2R2g2SlpnDjfY8VuW
EboxZRFTNxLjd4WCQ6+DlIkEFi3X91HW1zPVaMQfqL8yhm1UNIGKf4MD+38aWtsnIB3NuKSTBnX5
ijtCHuJPEMx3ZEjp97FCJQvLKrfM/mOfwhClRLuCeBczKIHdokz4Kmg3SM9UZteOE+qotdLsKYlg
cFO7njXH4roMiPswgraHCmGADF7n0Ql2q0I5AoyYfeu+n81BK1lnJ079z0x2S6ar1KCg5Yu3m4VO
h25DA1UT/71UV2Toy+o7H2hiCeiJ62Etr6ZEk3Oi94eg9yYgrv2d7HgteEoWM+7eNHKDUIK6P4KZ
XHa4/0A7IU77zLo97bS2c3ZJcESl0mTmzIgPlP8v8u2E91LmEGJpaIl8ed5XLNMy/+QsY+dFDRij
7v2VFi8tPbDwgBiesbdCp3ePFF+2a+F6Zy97tXlvUg95kQLd1QxeinALIstea5F2KNi+tY/IcuZb
4uS/bDgHEnKiwt2c4GsWtVZeqf1cjRQ6FiDF5rLc9spEV6HYqOdYu7cfZbiW2j1CfSwceEREonyz
qmot24vINUpTHaMA7lFeTzmwYHpi9LmG7yILDd+DilSdq+MwWnipRO8TWj6VC/3dakzSNuA3AwTO
nG24jNxDQWIsWjXhwxOG3liV4pPStfOZrdfzFg4Pj3KdF/8ciT32Wms9crUnAqGjSE6YNrA0P2xq
t5wwdSYExUrnOi7sCX3VL6gFqMEZ3oMieYKc3ooDQFsiDlHYF/LJ5hGhLlT/xg61rclwhi1Ss0bm
Y+HCOefbX/dGHSCJ17rLLVlK16j+0G5iVDs8PLJeGzfSCxI49Bj62+oapOhfcGKlotkAsGHGTIJC
S9oWEaYeHYQRE141czPKEb0Ox2XfJY0tuJ1UPoMK7y2KECFac8ehzjE1sDGENU47Iq8EvUIhv9/o
tW895cr6dtW/dCeMlq6Al2FHAuVkogI+hVQv7cIPl5lFFJcicxlhmoXiycRZ2/qZ+ellgo2riHX5
Kja9/hz1qqFzNr2GgAfrQomoCDC6k5fyr79EduxFOdEb4rqNZDqbViW/WnseKziIPA0/7fQ6VSge
5qXfAfOKxlh3lOmml4VISHE/tS/wifjPxVCx+MqJKxDd53A/VZdw3VAQ6AziR8Cu6s2PXInntUJ2
VDDOnIRKSNwSujGbYq7McpbLm6+zY979j/286VlBOsr1o5gdP8yIH6hHFCcuc7GxHROy9bMcfgX0
PXE+ANNKqFupglhiFGo+Q8sNofA5QFp4vCuEviTfztEqZck1IVLui+rfGmIC8PWM3kU4ePKuo64A
HKcIrqDeAguQ7jVmBLs+gXAQ2wXtz8GkKHgA7zN/jRmK6B1cAIfTdKPVytutQGf0fXulONbnnfOA
S0SkplAE4oExbZinMoEPsi/O55794XEFLzsMejEmJqckFT9FnAhOiPXw9yu/4hjQA9IQzhIzY+bb
SM1PUTWi9++MGGJQBJxOUq8kISmd727/KV3AjQp3Qs/UYw+Xetl33tnM3zahFPuah/K+B4EQ/cgD
MLIPnbPxTvJquyl33RmhwpsyYlyp6H85+6N6IiAA0zsX3D9JP/TfLWlqMTjUICrQVrQpzRM4UV+f
rFO7FVgv/zF8knoZNZKy+VCOLtoBptD2BScuUbEGCsmIoijShKhtIjZeT/yUrveHk/qNrXIu/L0D
C6FI93/WQMovHB1IyQHygRQPjNADGBJbdllCfM6lM3dpTm2n1j2fbre6eRbotBIwlPvL/tPw4Ag8
KHaVf9xxNVVeqeS30Ah7wi14WqbI6E5/zSc9eQVcom9MKkCARHADs70E3mPUQ8CtwGP+o6Xq9rao
g9pd8N5TB0r4h8jcDEKEgDlE/fIFVRcN5OYNgTC9zFHcMOHovQ9bTzazk5y5cUo=
`protect end_protected
