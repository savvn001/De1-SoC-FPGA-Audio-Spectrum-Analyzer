��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	;�׋�ŭ{ 4�1��D�����&^����5�U�5^0qM^խl�/B$�6�갚���c�����S�IK���R����紏�!�<�"��uj�_�8�˿���9h���OE�M��y�ɳ�F��ă[�H�sͭ�{Z�����U�[W�Q�&0)��	_��₂҆w&f~�ax�,:�M��=?_USM)�>J�PE�_rД�����"U��?y6o�;f k���S������S��x�e��-5�N̈\�T�mt}_��d&&��!�/<^̆�~	�
(ۏ��,�cW~�w����e08���š⚔�j�$�&Tx� ����9���X(����wT�<�z�����<�¬�{��_���ȍ-��D�����W�*F�+�k�FW#�_��O.�8(Fb]ǅ1j�K:��f��5\��Pը�p��2):i����ck!�SԵIo4�M�Y?!wձOC ^F����%2�+��_荺�y�B`=oz�pW�����:�'��-�&��5�ɠe�d��.��p�6��%.�2��Q~���
��2-K�G����5(��V�����re �T��>nd!
��k�'϶�c	LYZPn,rj�x�J"-	�FI0�� gQbc����GZE՝]�S�4v�6}=s9Y��0L7�K�ώ�Cr�޶w��
�5]�P8�_]����T u��k��-� �7��G슆�Q�<�-^�|�k9�����o/�����D1�V6��(ݪ2�b��'�&��\��ö�E�ok�zd���2�U���9� ��W��O�2
um,�1	�>A����c�US�.XK����$EblR��ؚ���	������j6�i=ѥ�i��lWK��<�o1��En��^�ͱU���ӪU� ʫr��oM)�6d������σ>pS��2dK�S��'o6��͝-�B���#�+9v{؃��X�l,��k=�![�L8�Y���Hdb��d�|x��>�n�X�Ҙ�1�XM�p]���O�L1���qV���ȗ��p}s9_�� �GZQ �`c�#���A�ZD�g0���)Xa��d��.�=������א�s�Yn`�+��
j�4%�c�+J? wؕ-�{y��"x}�;���:L�urŬH���M�i������.�O��Y�k@����/:�)��G��@������@q0���jt�;s�Cd��;߷�@G�/��!czϭ0� �Ou���N�j���ޙ�Gmm�Ux�Ǡ��foy�8	�t!�呵ꉝ�I��1E3��} <F����BB!.5Y�~��� ��}0Ï�s{[/ͫ�R�g�S"ʲ�E��U��RV����)C��# c�;Zi��fY�f���;Â1��Ke@V���Zo���G�\�"6��Fb8]4�S�|�N	<��~����\8�3	&�����m*#@���Jy[9��bW��������3z��(J;�2�r/Qs�6��f$�܌���w�N���f@���D;?���Ak"n���A�n��}��s*bC��
_�Ҕ���ʗ���<�Pz:�Yf�#�W���R#�!�F�>(�^aa���t?����Q,�v��9[�¢�?��?�<gkR��H�9��)B���TyS�e�V�3�^���l|"A����%|1iA�B}�e�T���L��
|>Qo~���͢������D��x�6�4�%��"�$�b5T���nWY��\"�+�1�SgC
r�f�Z2��X�Y����Z��َb/��d�A7�W0��t��ހqL/�5��^E�r������^CY�+
?�6��\����j�a���f�\UV�<�:�zG�)PI�������^i��ٲ|Qju֢��H����v��5lr<���`Ǭ9c,T����C�ɪB��j��j<�e�xz�6v���!�p����?.h����l�!qr��T��VV ���o�j�`���_�,8Z�%�ܺ��[]e��Єjp�*lY1�m�YT��A�;K���%[|����*B[�Y��Vh��x��Eq��Ư�e��(�Q [B[��O�(�d��vƢ16j�k������ ��4��75�{G�sF�S�e�[����S��4�D&�����a6,�n��g�r��	j��!7\�+NgOHgX%!���C�qV;��лT��szW��{���ҟǸ��'�B�ȌK��&R������Y�17�i0��%X��p����yi$�ȉb���΁�Fv�'�'\�Z;]��2�3���4��-��Y�����	�a�B)�Fc.�m���@'���w�@�IS�|F�O�;`�,Jvw��$>��E"R����P�{�nF|���mܐ�_�D��k���"�+c33ai�S��~��<I�.5'H���BFRl"B��bD���������s��<]>v��$�X	��������\��W�5�Q�:Q!�৮l�����ep�[9��.��>eՌ�u�}�_5�y�{eỏ1�*._�_.:'�[����V*EM�,�GM%�m֨X���#2zv����'}�qPe �q����b]%�{�8)�����C�3O��fy�S!2�<b�4�$t"�V#٫\7������#-�q�L�NI����"O*���,I�UB�:U'��=d��¬�.~z��������,"4$0��	3Q��g�m}���o�~4�<����]4�|	ٟ�6�q�Y���ǉ(�I���l7��'N���B���<�ȱ!/��S�����!��<��4���IY�}@m,�3�me�b��/מ<�8�kyKS�DD��P)���Ѩ$�����)SK����R��&�Ǻ����d����5~�?X������=>�s#��&tg�{bX�+���N��,����OF�Op���{t'�LzC�Q ��X�Yj�iUD�rn\�J5nޤ5�:n�����#܏�ΏNC�+	Q����9N�t�mj����~A|�E��ts�z}��Z:Ӑ=B�%dHI:	���xH\��qi%tp�˗���MHkrP�o�'2)٨NҜX�iY�Eɶ�+�%7�fG��1��췼/������u�������������c1%�s擓�@hM!��
+�z.���,J�h��2.�B"����[d�2�O��q3��i�0t]���t�h����$:�I�ՁU�M��jG0s�"�[��dB�)G������������w��u�g)D|{�M5B����Fv�AF�GaH]��or�~8no8�+��dR��!e���R��EA!����(�l
�@ r�zٸ	�8��*�N����]������e�	Zc��K�]�FMQ�r'4 x����ڀ{w���VY�G@��T���7� ��:7ɕ�6SuA��<�O�5�ё=�LY�bѯ2��Uơ����R,gA���`h�ȂX��?�$�I��xz/*?IǮ�ibeiU��/٧'���aB�D2z#�0��Q\�7i�����l����k�]��<��.֛�$Q���š��*��ط��T���4JR��>��~V����n4��y��-m&�8�h�� r�������޼ ���8��'f&?%�ڡc�E ù�v�P�R���/i )�3��=����(�����]�
w,�|�UObo�r��UP.F�W�6w�6�S��g�u�i_�%��ěD�g��	��M�?�����Y��L�ŕTV��Թ�Y��@������ $��s���1�d�H�c:�z`��i��,�g�����yU�_�����#O4��!��R�.��Gv���t��������LT��J~Έ�wp���EZ����לm��W���WD$'!�t:��z|��Xd�a<�I��x���G�"ք֓WGN�o��;@s0)M���2��}�ʒ�d躋]�8�oXS�V�|-Ȍ�u�t��S��J�eo�^�V\���P���Í���s�[��:�XK����WR��(a�g�p��L�`�o~���1p�7S(����zࠟeŶf��)�'{��ʨ�Ŧ#�h��ر1�R���%��2;��h�M>I���.��������[�*A������Z�ȣ*g$%�亇�b�>����۳1��:|�2�lo�aĴ1��>�n��l�\a@�F�#y�$o1ւ��=��n��B��T2���=9a[JB�ޯ4��w�D"z-�+���{
��V'�cO
�b�Tm�`ɇ�����A�'w�f\ܨ�um2�h�XD���h�DZ�Ϧ����!���57M�@�M�:�rr�t�#��m�#1���U������Ki�'d��LK 0���Q�])b>���j�q��J�S�n�Q��AiT����t@>��ܨUɮo�a��q�բQ��|Hm�LB+�%��~�3ݷq �A" �"�腄6�Ͱ`4��68���&	΍��S߻Qq�lS�3�p:��A�w��X_r+�G�82P�*�gq!q[%^FA�7ߟX��1��Ms�]��E���s�(�j;Y�.v���-���8ed�E�i���7ϕ�[3�Ah��7�o
;IC����9H7�m6�P�;(̭��m����!�U�򃄎/:��Q2�8�w�(apCm���0���u
p��m�K��K�\n��Xeh=�U� �7�KS����;�a���>O�N�8j^��׻Q�Ͽ��~^z���'������	�z�ۮ|J�1T���
OAv�!*
'�����{X3Z��%�TH1^�0T���*�D����[���d�`�a<4^�nK�(<E�_r�0� �
�l'�JA$y���Hd'O���;Sr��<�Ə���K�|���7��T|�q�	�6�>$�/e!6	8�-�Jl�F��������q��T�X��-y�b=����*6N5h�����na�b<�2>B#�R��C�$��c>x����u^�HOB_CNt����
d1����b�Z,>kJnnT?@�Vy���/�K޹�-1%������z�S����?`����L�[��������X��J�����j���GS�Z�q��!�>{�.�බ=M���S,@B!�G�^�V���D0�BGN^�ŽR/*�r^"�jK�B�I�[�'�oĊ�M+��6�z	%D����@�k��x5?��_ Ѵy����v_�.��9M5λJ��P��%?�H��"�(n�l^��$QAB#~0��x����� cO� $�$��7���-�	�宒�тc�%f���E�
VN�~qŬ����<W䶹S�h/{�͇\����Z����e��<H�6�Y'ڡ12/�C�*�]����e.��؏�b���7���F�Pۣ 
ؔ)D_����c-#��QP}/�˽p�v�	k-�m�VL��2��h��QX�&!N�(y�Чܳ@tި�-����l�?�������`9d!��� f���@#@�M5�HT/7ͤh�=T:g�i�����Ͼ�/ЍV���R>�naK,LV�����2Ӳ'C%@V'�y���߅f,�0�:ЈL�Ŗ|���c\��d�GW(�O'p���6}��j#[6b�9E��E�ٟ	]l��
��~{F���l<��w��5k?�P�t�Pr��#Cr��A�Yq��w�U(KYo4���1�uS}'L^~��qS����X1�Z�*	�h��
a���ń�^����\�����5�l���3�L��hL�j�W�C�.���j*�W;��酅�<�
�f݈�:�b5�a.C(����Z��o\�T�r�Tt����M����nZ�-0��k'8	#+��-�2����>ʞ�W��DTi��%����[>�k��-�m�n��jҾ�D�-T��X���İ�Om{�~
��]�Lʎm��Qg�v� )�`�թf�ۮF]k�2��P0/|�� `�y�I��xb��کQ�$�v�~Dү�}o\?�TOdE�<�R��=6�;��K��݀�qbha�G�3n�h@�J!G��qR e����t�<˻wvM�����\�AgN�)0�X�``�AF����R�eq��E���'��k�	�t���Ɲ�'Reϥ��ĖyEf䝣s��8T��lP"Ŏ�#�|�]�m2����R웹�^�)t��OǮ�7��A}��\*�s�$��0��';l[Y��s����)}0�olL������˛��ݳQ�龪�I,�-~��5�0���55щ��|E3��=�eL��)���&}��xR!X$��׃�!�!�2�	�9SʟTӭ ��<.׎�f�8�Q�=� �GH7�fhJg,��?_X�ѳd"$,	���M��$.�І��^>a�?����X��@�gC�5�j�H���}����T-�xtQeW�yͲ�T+�W�S���F��A��Eza[�Z;B��[�M��)����a���엝R��)��I�2	��mV?rV^>���0�6��%T>���Qi�~���޳(G�%p��G~}�P��ŪҠ���Ɖ����r���
��=O��E�f�Zv���
u�ڏ�����;�Y�W}�h�@q�l��
L~n�I܉�����mJ�����3����<�;�Xmt9�Ⱥ�({��w��<3�>Y�uf���Oh���n������=H��b��l�8VW=0�r��'z�RO����zTb�EuN�z���6��[�?�
���������5�-���xkocn\J'W��+�n漙J�4?-�ǿ��&N�-$a��x�k�u�����q������xih���'M����o������uL�Z.	9%�i�������~{.�d�C��;$�3�v��h���å�]eGB��u�'��B���	��d��U�����(�76ACխ4S﫬O�E<{�(�D8B�Ć���l`1���&ʍ�t�7��s;D�Қ:?��W�iLTj8w'SK�h��}i9^�����*�p�\�2�;J�_Q�G��
-sƘ�W��&�5@am���GwF�Kzao�~1��E���`  ~i�l���-�}m���\��ϖ�"/8�g�������5���C�ǖ����E��.Ŏ��U�WM7��~+Yi2Gn���i�0��X����<�����]Y��ʏ���2կ?V{d�-:��~��[`~�!0VCK��bX{�n!&�ѵ�^���S$���O[ &�t��k���n�χk.��4�k@`�'wt������=�"Ĕ���e}C�.�'��vmo$��M��r��k�
�U�}�QD����9X@��Q��1�;�w��L�Y�鿑t��j�B�~����`7:��F/�D.���8rY�c@I���a�,R+��
��O1�Z�f�����W��yP�Ro���7a#"J��˺E٥�5�����{�)dR�Ox�`�"�X� 7�7��a����U�3Ů���э>�i�T#����
^�U&�!<�1y9: K�d�lpy��)8�'�/��}d�؛?�+�S�K@���Z.ƭ�+�|�RS6�p�-�z�	�$M��S��oA�B��C��Y��3�߾zJ��Yv�u�cl� ��?�ݯ�2/V5|.!��5O�N��~�a�n\��>A32��Z~J=�BzJ\}�0P<�� Ͼ��������%�԰��J��֞V���}t>�r`���m�����e���u�~�t���{$�t��O�hxEȖx���3�W4.�Y8�; >oӉG���,��Mt��o��aގD��5���z��6�5�U���ؖ�=�>�e���	�1���^8O�SA_N��G����Lh�pq�!]<l���ɇ5F6U��gT0�W �,UtŇ	������Ҕ:�u}wX{����'γG�ڲ�& o:��o~rUY��W;���.FT}�\0q(�M�J���BA����T�^��1kb�I��[6\�*�~!{���+F�w��J=�'�e�|Pnp��!���1�A��Ԗ���N/�@�aVxRF�
�v�R\䓹��-AdT[/$�;Ǿ�賴܄��yl�2���`������?�X��-�7�#s� �o������ț����J���c*"�[�J`;ܿ�3������Z���'1#
��m{m�����Rs���eG���B�'�l��H�L�b����N��׺�LSnՐ�d��ES���P��E��޻��N��Ӥb-���k. n�j㜍�ȵ�n� �.�I�A(�ӴvAT�ZBd�r�}�/޶Iᮟ}�Q�6ãC{��Æ(κY�}=��k���]�q�e�i#Q��O����������!��\�(�b]p 6�e=	�cI38���>V6lI���(�3_�Yp�FBqwp#4���"X�J�(���}�Iy7�a��e��"��ɚ��[;E�C�ܭE��7�C�OU� 8������h�詓����Ѯ���]=�~^�RtO�43AO;�Zk>�ka�[��ѵi�+�`?vX�`��T�X�9�)�S�HL���r�-�nV��'��p^�4ͭ�,{�7��s=�sO$��.!,�w&�\lv���u��5��:)�;?��iz�������$�K!*X��0���� ƺ��;�\�n�g����W�I��ת�ɴ<4N�{���!�5~��
���(/�b�/,V�q�t'/�*�����N����.��/D��n'��>k�%�-��nc%~tq�9a��!�����6�k�a�"���4�ty��h�U���)H�Sl=��߅~9U0��?~G�:�̈́�rqp� et4�X7<wN� ���o(�����8@�|�r�E��P�	�,�U�X���H,�>��Y=��_����K����'a�����k�|{���~�	6�P�Gsf���X,c{������e�8�{�p��⺵�m�ܐ8��b=8��ם�����X�����H��A��)u����Y�Q�MI���Qq�7������YT6��B4#��o߽<?B,��s��D�`n�(���^�"W~1���݈��M�.ZG�Sf���oHÞ��<�M��x$�/�^�*�Q�s[�r�J#._q����t��D9�>��OF}�:1$��,�&�ਤy ��
 ����>l�7	�:�4�=������:\�tk`�f��@�`�!�Z����^�t⊢��l��W����ֱ��N��#�[���@���m-|V<xT���N⯶��� N�J�D�$_#\
"����3�\[F�	K�y�����|h	_���X�<_feuZ&��		sx�"5x�ѦX��F>%M۬h�*]:v��e47�FQ
	�"���b���G����F /�Ȁ:�����}Ȋ��"G�=#g���"�9.*�Hr��()���m�w��[~����:�B��:$�j�����X��@��m�e�k�lC񲀏	zE�ȇ��Jÿ��)�J�R�]��].F���{k�'�9����C�`=B���ɐ`Ns����AH`<�
��sM��l%�Sy�g�q��[X4+ka�,e����q��z�S�ԋu������3*l�Uң�*�y�U�Ar�L$HX�3��nK�����t�Td���@��yG��[A��$�%͜ӝ�z�� W��������Z�{2zC�Y�k��n�·�rT�N]Xx)� ��	�-UnJ�$⩵[��%P��Fs���a변�e�w����=�\K�����G�-yL�-� ��<�K M�;3�2 �Z��#Iq��}��z�~�F)����l_�+�K �!��0���_������"��W��v������5����\�����}��آ ;�pt!���8۬=?&c���7*�o/��7�XՇ���i���A��7��o�EZԂ�Zv�L(���ˎ���i~9�W�2�8&�ՆD�U(7j���M��Q$���
^��?&W���V_�r3tU��}E�f�ݥ����A�wÓ�1���FGh~�x��4={̛m�����&�v"��'���!4��eN���`���G#k�C��i��u�����8fx�1���~{L=�v���T>�����ޓc�����>��Ը���_�޾i�ܾ��4�q�X�f�VQÔ��p���{���&��O��5����L��x��w�_�C֟��3�f�l�G�d[���۬���r�C�zl�f�	`�[�T��d���-"1Έ�,Bo���������s�J��qu��=ȝ�����uqwXʹ�����ڥ2�1:b�.N���?�K+,�s_͌N�@��f��a�8���=�K	��X���C*����F��_s똑���s�Y]!��v�O�ք��w-2��T���FE0U"���'(*Cp@t�z�~nQs:�e�A�'���!Z3�|K􋫕��`*����-N�!�7���#Ro�䥌��h���.S��z��;o�㤹�����d���
	�p'�=l�1v3W���K��Ѳ,�ȶVP=���-|q0r���n���88R��P8 /�Ly#�����Jv�gi�߉v��en<�G���q�8�����6]�c�b�{ВM�����}�7�ȡ,��y.�s�z�����6B�-u1�o�I ԇֺ�}���xp�b=D�b#E<P`�i��? �q�c`n{��[���{I6*�Sc����c�Ьo�Q�{�'?��W�GZvQB1��K@�u���3��yh�����>%a���hVK�7�V�'�������ywkh$�J^��դ1ݓ�$N�[�\�+{�[�����L�#��6���^܉hJ�sڔ��9�g�������Ė��w5�Z��0��޴��Lҝ%�o�ݎ+���	�!ͷn�u�0�@`{��ݐ-"�?2���,]p�� �Z �s�����z+ U���h�)JQD�� |d�� ���`<��f[�7yR���y:Z��D�pWl��=E�={X�o� |���y]iz�:6�@�-���j�*].M��+����K�f