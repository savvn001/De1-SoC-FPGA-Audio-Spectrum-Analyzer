-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BEQiyhjNyuOut/JZiInM9BfQynz622mOE9AXJgAcjX/jYhy/Pif7aP8mR1jgfmatLcyH+yKIpJbA
D2TA/ZI/FeaJUQ9b6uhcO80HGrMdBgcD/TEsueqWa+jNx1zUy52YFpPiEYmjBI7Cf0+YwUdEwSPb
z9QAUyBe0mO7G0c2fqLqRRYtc4ouqKj+p4vvJbFK4f9VHKxV3cR6LQEMb4ZUCMH0MxEle6oxrLoR
BC8aeHaePTLopeKU8HuHfjSgk4wPHHza9xPX2X9+sO6n4ac9Z2iH8EET3fx7i7kjzkLMKhFlsTie
VD8rkgptYqKQc4Sz9K/f19NLY9/blZEcYSZfew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14528)
`protect data_block
kRNxc+W3UCwEXHPRPBxyet47TBhedqSOyyMF/u2N5q9LvvQrEXE6jJqcs1e/CkXEk5PLns1Kn3IC
M9KreLWPg9MDx7NsA1fHKY1jRuNtL5s2xROHsAE/NPr40ZwpJHu8YtnBIGWevTbPv1NRe5FDi/rl
COAcXlrzdixAdF49cQyivQwPDSKwfLThWY/vqenRlZR8OT87stMrA8gShso7oapQ9Aog+s4DHw+L
dXs+HHKbVGvFGRg7d8O9kGYAk3erihBxNJdZ9Inf7M/UsMeDFz4bgzsAr3MTSlcFAigpk7/eeF4q
6/XTRiDMbz5HPxDuynLh7fCkO06Dja7E4DafDEpGxp1ovYjOk0EUV1+78QljcLyuR9nGTkA61loj
r2k2hXZdAFMq4svzCz6lMG2d6brFItVOnv7mH2J3/3NIERBPHOFOqzFvsTzaCEMtyIFMSkHwQZox
oaywYpVZayqBKPgc/wcReuwjzj+eYvBzGEhvatM6Uu8BMXqUfW0Ck36XJRiRHKEseR8cftbqGaS/
FclzT17jKbiBzpnqNnKuEPW3JONr+lVUoa0Bc1VHb9sgj2MRZE1pUBNsIIOHhanXwyBtJCLv0wog
B8koggBzMK/oA8A9rh4OOXJUiMnvRmbH26qLdqBN3VjSoyJslAwhaSG1k/8KIU8lWBadoLuAWeZ+
uv+NhkzLijiMZshJWlnTsritZIX4H/6rNmviM5BsOKwGASQ+Trg5D/9iECs10eM6T9Sfr0Oz/61/
F4qH/m7ltTyILiGc70MGg3MFV4+iUbsHEuuSALJY47ounl1543DsqhIIH2bKAhP6qYH2rg8TwhwU
RU4eMGsJuIpXEUtYuM145AdCh+CwqAVFXHUctbMGMWhzOOLl8HHYvfOrHa9V/snCkZ9GBjOOyQGB
pk+bGghwUTQuk+ECwF8/FDQ8ijYuhZ769Q5uahyBibAi8KMnpBbvSnWjqm3mCk3S0uoK1Xq4M+Wu
zZMY7tdwa5eCAHKLcCarbu2UACvQ5gxJwwMgxkb7KJnCNqJLONpzbu2bUR+G4qaTdZXQ33qc5uVq
BmMwaa+USd/G/uaskcefsrOPTaes4EYrcjklZ/ClpyMQehimW9lB/n90ttGySKAzO3OLd6FVf9bX
7LIfrUHTJqPgUIycLUzywcjV233X/eBngvSFB4UjnZ+GsfUWjg9ykAB3jbBCyYnokapUh5pY+KM7
v3n9tRAKimF3R17/rZLWszdtOPN1Vb/Cm3Q9+Ft2ayvZS1pRdZePBk2uKuK0e3EFlAeFUc9IXPH1
9O8ytYDwRxYvBNqnYPNs2+0orWvflbGQ8K/uAX6PtYNAu+mAjXVryPFoNl82EqOn/SyZD2ABBGYB
Rc/LHOTrtws/MW8LQvLRwpy6JyxLx59QXuHOSkDDPsImomXqokzGjQkS+OgzBmENwg0NdZ/jhFjv
csf22+/1fUVkvxuw4CFC9XYvuOo44WQ6Rs0ExuhFczCiYkPK05sHJ1lRDqWmfZusfQoA6q8xG+bA
Yy3dg0QoWlP0n3tii9rdNPi7AqaM+uNF9WCQpPk9/CVITorJWo6QicA5Y9RgkhmdZld8i1qDnDnk
bvOEtM4FqheCcif8kpcenltSMVno/dM5AWMwGQ7UE5TL14ZpduIs0avJ4R/VHN431+vTO91PYVxa
qrs4o/PpH+JL71His8NRBoRRsycr5gT4dfdiuM9tfcm0Mb07QUY9E12Hgss7euRmZ2mlwLpzWYPp
6KH+sbUQR3f1xd81ZXKLNgMXqLr/Ef4rc35RC2FvIMhG64gDSUkIuyn6Iy5sslsG7pC2dJq+HRMK
pK4itdUSwL5uvOXx3+X44zBP2JDq7nCdO9h5cS7H8mAnoagxfJzfNu117o2fM5v3tBqIALrLw7pK
4rmLx+JDyBCCpLWn8WeLpnd7Roym9dGBs7uWo1yI2XXl1XMTj/blPKU0Qwjauuy18YWsp503BIPh
jNWmxZQLr9h34buF/qoZe2e+xJtmsY0E3sIDSqXHpP3OluQ+AcpSV+SN3dhAaUStvJJiRIaG4A8f
eZDh4Z4Vh1T7g5hhmpBl7SNLf7xtxFH31erw4lAtZII35tLBiPFjhHht7AJog7GghznJPjhr50V+
QWBT4UA7hSD5jUoWA6PGBxraODghiZJhCT/wJmxLe6LNu1bo2r3l7tVLfAPvewepLpG7NZvRhnMa
NQK48z2n+P0uRupY+QuFPsHSBTIOkpfqj4aJQslDxf0ymAL0FY5naDXf8xExtmHLzXEDauXjwn6w
fDznjsae1MGb/azbrn12vw0p1gVodb1lnT86OfFwtG2qOoa4yV19ZEkxCyGb9915O4+mj49uUK/6
Kaezk9SZJ6kQGFi3A/cFYR2Z3Bu4jAxRU5wf5cyNiyy8Gx6md2OyVXIK0qVrksIpu4zLXN5gNZSa
Vi2IxIOjkSwxuutNPHmFX/aiTqbQTSCyObqQyFn8JTivpvlDSOxbI2tjQcj6+E5E+jhtytAyg540
+U3J+x5OrUyZ2n87EmkdAMUgzAlDho+iKPbD7nFkP9KMSqc2jBdxwXBSQh0aC/0EJON51pZS9zaf
HjWjlj1OKOYKpRzdcv5l1r9nMxya/4VpRTJm4L14NsqSRNhji3XcDyKTwKW21KWgPG3QuoRA3Hk2
ATr1AUejR3vvD08cYTzn/x855dx8Ll3CJf/M71gmTZ86S4HD26u05Hmuab6H2POAUfoCa/gNI/B9
Bk+0DCq+sTAXGhVsDTwoTwBelLTM2btkD6R5K4uuR9AYyxO6nIgavOPiCTVY8ioJsAUridXvSyhn
tRJc/o0WwGEe84PrudXrFBiB2Q/yaLfvOntyFiKPmiB8GoXtWNGraqCbfNkSpmzoB9PnTCQaoW4f
94xV8nNcrVeU7sbCrFngy8/hOmNzVeXyN7hxBY0xtJL1Fu8UJsC77obQyAYvcYtMc/e1KaPinUbY
UYaNhyjTgaSb5DQSodG0bywKBzVNbxjU+KJ3GA8R5f4fb+GPhKKQSvGiV+nY34DHXXnhQhyS1mIk
UuDc/kVm0RpU59H6UBoH6wjEAfdLUy+wrxuh7mevQMOkgbycagIxNxkkzURmILgivuIIcgpK6oS9
YWpLBoT5lj9JBCoACp1dud3r7fmcgcNueQejWkbIgzQBj9HbCAqQheOdeKv86qYI4+wWTUxPBWGf
YMvpF+iiUo1q4OMP1x0ZvgOiUAxQ/d/UCJlE3YGLcfVDbNX9NKiKfE4XonSFmYuQ+6wrCSeKagqO
mvFhy20IHTYD9WfMBMLp/euijDBHhRK6FDrycj2qXswGnF3npQfns+zAZd2o42BimEzkbUwK1k/S
9jVPiMq0GeidpFVBCdvWgObjjVm4qqDJjOkvp4uGdTMK4p/Ua16StH360SaL1YU+Djal3ofJboi0
kXUph3DLqqy7C6Bo873vR+kDQxZhcjFkimrrPIn6EFbs2ReZQGJO88ODE6TK5FTq1rmBmE6SYobB
lpQATG2Je+ycVVg4rlYSSMmzIJAuIfYt5TwLIniYWr9ZYcR1Rlg/zIROzdkdk4D+X2rNrZjG7ZvG
cEk3kwedi4sw+IPNLiQ1kLjAZB910aJQNDWqt2wFfdq3ejfIflJZdrF7bSje+QB7IIm043XSduVs
ZmML7+1K4PiJXfcT4vy/S6TAsdQ6h6hbnrYwVKeoazr5d47mDZO8cXc2jK7PFs2E7azMDL0e2eR7
yIRRML8X3gWkt6wgqdQ2pSNohOge4OJd/z6TYSh3g72urIJcvtFPAZPJ35o2AWs5PSxHNbaR7dAd
FYStHrJmTiF79+PmrfjSarfBoIPVrr+FGnK1gxJb1Zl9Phw9fzQn/NNdmnj+h9igFztPDBOeNo+6
D5HF3Uy95lRtxtkhAEIJrJHezm1HLfKHRpX8sVgCMXtGVxiDNpulLkMFN0xcWkRf2Y8hDWJxRabd
GyOaDkfim/We+VFPoFgiLKaTJIxO86uKTbDNNpn9T6yirGhOLzmjPo9zOqLTNVUvqBhvWoLNTF0t
ygbv53qrXF1tIZD9lcohPM5wzvuZPB2Apum3mXvqz/yjdYW0pLAJJqGOfuf4nyige7ANUuD0NgMa
LQdLzQA7N7F+x/qukkEj7sb3ApcGXiygGPV5nCTB0C8/wyy1/o6AtLf2sN76I+LpS3hKIEzeGwOR
ZdUlnpXcTQBUw69GJbKe/mp6o77WeBQa+y0b9oGJFczsXfOreRJiPDzU8zzKaBuyoJr0K4r4/YCF
DZusN1d8mIX27fvDVzTHEHmQSG8RSECqZteXdmEEoLhmjdikURP0CTL42N5hn4lYHKLzYM2Q3//e
CKHRzKG37b4M5LD3xEFKHRsoFdxASc/lUGiThVyISiZ2ltA8Eb8Yyr2pBEOBe71gZH5V0zOqhKr0
f4z/vzIMEyeCfGkG537ttfJBWxlobN+UsswHBubS/yyJVaONEwVinDyj0W0Z5RKqdXLLuc6ivaRZ
tayc893z5y7Gcv1TXNhrwYzi5Gd4khECyPPAaNH450daQYBsnyUBfdbXwenDY394858nOydKFd4V
I+RB2xO9+Fy8WT2N++jSz2HYJcoUu285kuOmP02psq4q4JtyGNExBzsfBeosmvFY6RVoamCJEtsL
+y0q+7qQVD+vyxmtEWoiJmRAY0DxPvSrwmbMWjm0kMkuZYOW9TlnljUEGLLw/jLsHmdFve0P1mK3
wvIyHZT8gnKJ9qEEV/RC7BCytVWxQOaqO9qww1gZhgtYS58KmZGL2czwhOgctNDCwDpCSkNneime
zeZqeO7ibgr5w0gKs5085rFHzwsj/r9E6DvDLjsxnoSggbwdBORYVjVxm9vHGsjEzXHw76tUVkmx
/IjL9EnIUMo10I0uO2OpjVyx55FJh8K7Ex+PnOfYlyxxXozAKE1fIX0jgxfijCIHOOnj4LFP85bI
9h4RQysuSmNe7GlD2rrQxfZtdsbdhcNbxLHsUBzwY7iMX87oaVleObr8A/rz7RG1+/9OnCNU8DC6
6G+Jk5OLyXyltexPeZ4buQYqSlSd3sfb3ZIZU4FXxDmWgm2pChvT9X6TLVpPRrNvU6APuCRgdxzn
D8y6sMy8YbRlxzt9V8RAizvtFGRaKKmWfNDhEgFwFd45oMmZw4vQCG2dMXuo3+4jjiI4Xkm3FZM3
lxV8q5fI8/BvWKz64zyPh0DKFwHWuKXRNFmpsWPaUxnYGeUbIoHtN7F7BvOzuYXAeZtQ6DtojTTf
/rtzxfqjLKGmz0RB7ARoWrVN8fSZDy3KeSqoDaDQLiMHWRwraMARnZIIdyheGt3QU+7PY69zb99R
Z/OvJiT6fEAG4shtiC7FlRCiDU4odjH6LfpIbr3Yvr18m+gCCsdpxBC1/Kr455PMCSIUVOjOBlMQ
enn+NrXRBCK1K1jBrvP5pUdHjRXGwL+jCruNngKiFx6D1+t9tmB+PBWfQemQVRKUNK8lThFZ6eHy
MYnUHdzdLnB4fqJPr7UIthufRoPzY+4nJMVtDhz7cYDM6yA2pVwNz9nVYfuXso8dZpk8ZjwbKvpG
WKhj2V/fwP0PamXTipeh67LTuMLrKmS1b7wEasbloOnsG0a77y4yYwplB4y7xbauDCuW2ULPXkLH
H7BOle46iuqSuVSbn55my1B/ECYnpuBWpcj1qdQ2zYNkBhO7Qn46fUDsURCZl6yy9daRhA7v1qRr
oTRZOSlLKCHQa3e2zYy4TXJMJUFGNcrNMOWMpKOq82VWFHKjnewrd9R4cysv2jQ4iQgOOE0Pn7tv
PMRakQh8rJgLHnlweWK3T6dCdDWBS8er05US4GKGtk5oRb8tKquUZnoVjxHsqEQqdeiWmsnkBVdt
dMAVa1vEQwmTtfLiv0EQ7VReXCqwZIMslEeffUsQm7Xn1uQJ0ZY+D9wluO7wAiqlsj10BuXOXTNj
3oa0d4e6JI3a3bHEDXlKpQC0Wo0N+rMTkmHtI35GaAb3BKGjhdLXE52soCsF1grI2bKrVCugAia9
in3AlKIo/v1adcet6YZ30NvtjqZeI3uGZifunyln6mssDKPYai15Rn0dJBil97bfSLPyyPDGKeaU
L8AmhDtHu502g0ztPTn4l1I5PXGKcxC+MfIxIzq5YNqdaZvdSwthesbVq1/iDb9XynBXcg4nzaOa
cjuxYS1OwGDIx3CYgxZzYgEfmtXg2qB72Bvv+Id1//ooRW0Q31AzSipFiNq6Rh8BOhUaikgZqZDM
LobLvCDjVtjdMcFa1HFpaZJHimj6C2I+78M6X5dMnb7F2qjN/A6sbWhfj8j6FqZYykunWnBk5Nj7
FvpxlVA2adhP8WjYtyTnbm5lfXLxYlgv7FkOc24q7P3srF7k9qIZ3jOFGx5zBjDx3P6erGLDEttk
DMPw89DRjvn2M04wxBEKx2xrs3n1X1/5RH4VP0oLhy/HguSLyySLsTuEBVV5ynZCSj9s+XOk/j8t
T3b8ztU4QzoS4Ihvlx/Dmf3KuFLpM87y3TrfteDFIlq7U1xkF3XVpxJIcJ8NDsvILI6nKa9yQmgw
LhxEQuFN0McwZ+3KontUzGQHwlUQqFH1Esb+OI6d+2+f6mqnC2XFn3rx8wvJvRbHZmhuXzxWEzJ2
lLbHQVn3ui9lLZ9PO1lCzRgh43o5IP+lOA1hWS2usZOcuA4+uHIFETwTMFgOjyGr0Fxyr6Su3kq0
Er6ipPp/Qbt1eag2YpuvxZSgYZzO3h/5lWFV12w/37x4F6oUEuEP1gwGOwZQMwfyUZwB4mK7iixd
53MJtxDaO7ogw5D48zCdQU0Ew7W2TjSTqukWUOpyuKK0uLhmcCu6m6z2EwKWzCk4Dr2P0kmIHHUR
jp/KKZ8rewwTBq+hG6z75oyhRTxN0hW7N1jd9mjgtZDtQeOZAz1+I+nl+MkDztQfDOcxB5nhZLDL
hSJA5s/pQ+Xz2BAiBvm5K2q5yvPH1IU7Oo67NV2Sf0TlGX1teqUclPdLP8A/O24nE0yLQFJIFH6O
bivGdUEBXE6jfCgEPWa1nFu5Q+xCF/+zZGuEDHzm7Xsf6egipKnjyGU5sgsyMra3KFuuNn8wPUda
KGzddQemT9bybFaBV1SX7bPx/rRPLtalGhP+9VFqFvt1y4zJ/T4x3cJjQXYkq5lgPW0oTY2oSMBo
xsEXDoHv/QqX8IZCZVTbEnrRtOryJWflvBIK0SiEEeyyb64laq1kqkjuKXs87GqQ+2MVb4e1Ff/W
IlIM8GhQbAytNcIHOH8Y9B7H9kDOUVSVPotjw/fY06Pc69eqo1owkUKSMuPsNP6pimlPgcPtBPlx
Ko47iUEKa8/pB2pHssDAy4Yx7ZGBxO9kyH00FgV6XldI8m+0z8jdZPHqw92nV5dyXuLVeW2PmDzY
VlsWI55I1b3+XOA/tLcgsl5yZUxHlSulmsunnVZaQvZE/Dxs0JkBnHvdMkWGB9a+bFKJ7RY1rgUx
BxqRfcxaTr+XDgfCCVJdzakH5npl13LUE9/bBqSpaQEs2s+kjLuw8eNLbWgtx/dGqAhkqD+wrVCc
suz63kv58fznSQmTfLW3QD2CoiEmJlufkzRvzGRHx66iM22l3u6iOSfKJQEgxjP8K4gF8u417P11
PN0dz8PfC9GM0xZB+tSPwKtywKPekRHdb466lInEM06jlXNgiPHOjDsdozO0FvdRP0ZRHnTcZT1/
dET747DJme8zlo250ScxGOHLnE2WurXsueb2x8yvZIIN75JYSKJdf6wEbVSEG1eXU5I6n0bVYLw/
2mqUbNgbpZ8YqdW6kwX9ekFS3E581RhJTzcxzEdMFZdtOkeEvVT8zvFVQVgJG6+Pv9PncGP0b9D8
gO/9UonhjB9S6bUGlo/AnhGBdPfy4aK0t6cGToSlJrUxlPFTvwwGAcn6j3yKwUGloYC9SYpx+qZB
UtB2aBP+RN8MZu2EUfOyGTb9byqIMOCOOqeYon/RTBXi8g9Ug44z74/LA/z8Xq0jzDp85o3yUcSJ
OCrE8UdBUw1eE87Ivnrm8urtdefO9y3VSA/rYjuoCexyJEcv18VwXsuEHIA1BS1sB69iiE93zpNq
un26XpvU44UqiUpJmcmBmNutfERKvWTd4QBGpvrcc8/VqF+tC4TPEQTuQRsT8UaQSz5VbcI+uu3F
zT4cHSfQrMhzhHh0QdKTSbezuR6MO4RLxDUo5T58Ixfz/2a4Hwa55aGjtbUrVRl1XSaVSp6nm3My
Q5FR0QG8cTZF+AUtrHLungNNaqxV6BZNvlfV353L78zeCl9l6Xiv/Z/XdIgKFFSi1E7Ej+EMGPLX
I3ibFbpapDWAF3NE1qeDF9x7It01kqKM2QaCtrf1Be2pS4pHacNtPcMPS9Ffc2POgRRcNr3Qf70f
oj0Z4AEo5NUBfvegijloOwHjqSyiDvvp08QiT2N1ymYVnA7CUqf2BMH+qJ5wO7/yEUBqt67KNsY8
EEbUbcS0ksaYC+e6a428Z+Bt5iDJRVqMdNVH0hafmCajyLYVqyN+3YOrkt527lDBMslZNbvxDGjv
yTrpib/6pC35u/nKw5XrNFtFztMynkWZdg6o4anqrnQAnQwhbHJJ9JHRWhVtcAyv2t1CuUQgqPCV
V7w2RZIhdWvQjvwmEnL4MZQ8Lv+W3dsJOeREdpNUnyP6jIT8MPhjJdxDIRe6GxzljaU3ylMTm2Wf
XWJTKDgUgnb1Sns4VJNOoWvLroL3IXXLH6S0Z+7yLkIBGPQjNlP8//AxncxobE3NCj6tkSpnmS9a
xbbU5By2VxmYoL19Bi6HrklKvDsFe6fatfDMKFBvaD9QdgH8KfTPyi1V17JPw30sMLMze+jSralf
l0goiIsVFAg2NGPkHyTBXH8kULs6QVud5LX11yx2jOQ2bE3FcA3j0hTBqVDFlnmgQZL/LdtqfnuI
G6bh1/PgqtSYqtze3UoeAxChPoPCIqfPC2BnHslfawHcYRvYFHea3AUZjLhIPZyi+3VG5LEdOceu
5Waqz2W59ddKgBqJxjrPn8LXv8XwXKZ7GyzzVBNmGoxH1+IW/9TF2uege2M1BOP+sEQBC1Jbkm5u
uYeWsgVDBGJiHig09+zdQ7Ci8oDWlGbMHe2R8L/YknPutnbX9QbMWFYauXSUHRGMqeOJuvTpqNOR
9U3dIZGrEzhxttXho2M1tJd5bMKfp6WyGahzyR+/N3RxDn/cx8Fcl86W8FYSvGPG/sAz4faVORWx
WdUrqpO7qTQfnvGe6vWABK9z9E1f6+GRCqkN+ZbKnkB0rMi5I/fmSqRzNap3d3ctyNMXqDdjEYkw
jDED7OYr/CZWGL2g1NIyFYziihN8pM+5KibM0MMzRskVjxwTs91hDVPqTpC3jCxzius9vbInVQYU
lYy83d4k+wqoCAsUpsjzBNakPUbAE63s/bRPERImr+N+qUl95n5pJJg06UUB9Gd9LhW3oJKvOmSO
uONltpZpdHd3/cDbGxkbJgxYb2oaNu5Vexgak7hXM7OXsmHC/B2cM5jyYU6H+eGPhvY/YbbBRxZ8
QYC78nxxesgYJweJaHCTXv254aGpROcWaf9kKNuWyM6Z3uLWR/MfIbiXZLFzaYXJPrylir2a7f0i
p46ufEvvLEvxwkXQAf76he88duVvVq/aJHJvKrXDAO0lKmxDveGrjn9SoeJuucxn2m+fwZbkEUll
i/BGuxDM+KQeYKYwbHuyXTXyiKIl9woW2talSvo4ItRO9yHsaGeesrlmucPAo2yH+JFM5TMsoQ4F
VDMKGZrUyAwqwzRjSl3AjXvBxd84IO39DqrkpHQikJfvphibCngeWCQwr7Rp7wEHpxZp/RCxpRuJ
LbnvOg9zMHhaDzwAB7Jtv/fh0XPWlXoyeQ9P1aqHqr0YytX4Ox1od7a+eZNwJT9tBDTWSiSbxmvZ
sw+fPRJKEzYVUqqHG0vEB4Xlfx60s8TqAQAhPSHvSGxYM2J7edtoNzSUCu/Ap9yWmOqqA3tL39ku
0oRD9hQGQgtTiNB/15R4PytdK3YkFDM/BqP/Fb0dOAfxxsb+cUj0BEXr1jlyC3tOHzaEgBbjYTTD
yl/7s0gUoK4MNTyhWB2j4m2ybN+LvpjaRIwA0sMeKyxePf6+XJ+aJG25rX1FAbNBKcbYUCaO5YMx
HkZitB9O6K/s2pwgf7RFQRkDDkSEHs/UtnMBGZqcYLclTTxkg6BWtvmmTMzgF8JnhpLkHKo2hfra
/X9A/BD6thH0ivuYuSAkWLFaXDXtFY/aVtVJUklSBugDCO51orJ7pgjIxdkd8w2GO6hMk2Fhge33
dHPts2BADEdW98JiosBlGRgunIasEs7a80KoCwWY/JAW7vF8JsF/a5DvQafD+jpGtuJmJhTxeUuc
E1shnjx4lvcsv2bTB1oUsDSpWlbpVIuhzrOhQK+zwZ4ZBCWUkz6UMaxT72fmv8EMM536AVCZCxXf
SJfxrPmecT0rsgSrYZKYw5tCD2GLlvUvvopBAyeln3tPjk89kNQ+Rkv2VOyD1B99MJtmL7IHkq3H
Ncfx6hJNfxwJcUDqNgd9l/cYd0ucanMo/kncY2FeFS9WObR0p5x6AkNC5tCncgHrNr0TwbteGVtr
jokBS3mZsZdYmdoB1t4RTNHwNRT2jKjnfsWc3z+eubdTiQ1Ci/PWUdn15o6AdashpVhhzQhkRbRl
rKWQlqplOCDBh3svR7TSpgaixkBGQvpyVCGNw5/3gGXBe6heBBZ5yJybNeykqsRdOvU2KfJ8sIRN
S4GvznqWeXdpqYZi2vd4Qxaa3eqpir+cUdxd7gjPu3EAPFYKeeevtWyXDjYHxAAz9IbeEwCXf3MT
9zFDlP6rGTTKshn14uUxv2C7keYH6RXZRnAscEX0HQUpfL5B+Eg3IKGGga6XxiBNddXZwAOYylIM
ynAlHGsSb/f8Q7NXbZR9uRrvi1E0msQKl2DWcydneJfJUyI2Rcdzipo4fygufYhCorxjHD4CtNGr
kE/xICyMhYLqTAUfZaCvZeCzEBKL9UIcKadx61M4V+NsxaUfkyd5HSGaSd+CmlwR0gA73k6zQXM4
SEimNQh3+cSB+WanIwmnKu+7y6oSWXZPns+eNFIE3KmuVhk9TVHkwQI/BsL7Y9KcY54dxZN4rcbm
BPUSFPZXpBTYm4V/7lDqMt1eFJlt7KEiCvPOtCJqMJuWTZcnhu+/ICAVTtVViaVfQNDumowTIPBC
m9DVOhB0Cbb9+NIw1tyrD5JfiUwmorshHvfCpwJ0Nw+OCN3sd26XVyQ/I3jamQtgrNXcIDP5lX3I
cGKQj/8jXaB6GDiRBacanahqyGilIyV9wiPYgB8wjSvAAyH0KqztGPzuRRQhI05KRTLkDSlOgtIM
PaBXVRbLDN7eWI3aXCNbWv61iSq10UbTSJMFO0tUQROKci6ddqlqnYidkRXDnKnvqlP+CK5ETbM5
k2qYp1g18uwnnkAdrrgjf+kJslag6q4hWec255rBAHsCGho2uGKlgiX8/PEONYq56xUt+cUrmDR5
Q2+5gytSd9uiHCoOjLyl8vVlLhq3S/tj9IJml4ZvEkjRadULlCQWaF2KkzsHcIyLHbw3P9fGcsAY
wLwhBM4P+LL/46sngUDPrlM++qskITIuKbPeh2RuaBCMmmqCu/Ipta5Pn0KsEU5OE5YopAuPi6kH
YsRofNxleeDBBszMOiVt6lhmLv4TIw8606jtac+ZQCeL+5uClzSUDmq06RXML8n6hTRt6OHnaXzG
OZpYZW+FJ3Vooryr0Yve7luUjruedrlSwbsQcsNe069dXB9uME+XyDX/89rPD2fa6Yni3kpji26R
v7BgjZVZncMafiDzZCV/ZxT/oTxNQcGexFZRKHN5/G8onkaHLfyHsY1aUlpd4YZODZOUe0yvOPlW
z/uQLPS5lVg50MqEpb+KHpCF570g1Ez8VzFhtc9wTBarKeC9WQ/RUSMXmmk9k+z2vUC+ivs8Qt9i
9nVbeaQdp9SDIu8zjIl3CkOgFleQ3UZi1yWICiMNrmEEXaXIzR594lhk9q15zQjd1ijNUVLd4WKm
E/4XkV2kMkfl0rOfnxwvNKHMnAcV2cx0tpeCBKErlUyydz8adNh2UYm9WGgK/RLHLu0frrEZTCuf
ly4XhmQX+HSboIxkVrcGAfYkjjSDgg1bHIqr1vR7HguGCaX1EGKwlvchrSxA1z0RR6OsZjxZDtOi
DN14BgRvw4Ggm18fW/hIjVmo35jb9Wseoi4+SJvqCrj65qvdHUcgdRdZQfrUp+VS1a5XNeMrq8i+
D1dN6Os3VZmr+LGyXnLrlz8IGDEZJ5s5/OIUoPIKcXD9FTr+n0eqJFD0tHVV4lYgZYvyFO9R8Nma
RKkZHA5mwbBiMEpNSHh8m85/rbeoZSv/NWkgRibpc7lNdEkWn5xx6TetnaLbhjynSOt4T9Lb+7P1
oUanduiKHWHE7vZkWFwAy8Q88/Wm8+Vq/fh9QP4Iqy0Ev6o0ppRbObXMJAElbZHxfoDE/m65vnvQ
PZthBcDsBlkAQSLTrD6b+skCnptN3xQOvUdw9aSKmU3S9vESEmCbwrCsW+hrtOF/49Q/cl3eXuEO
OjQ5uEAwK6aT9esrXtnVSI9vW1THJTQh8+X+zzo9zUd2jHfR3B7ptIXsbgi8wDAhJEk9ZbSnBF6D
4XE3nauAaoDgQjzKgxabSbqj/TbaUvQ6lhyiBjQYJTGQQzZnbvVMeACPKBIa+UuvyT8CofJEgDAS
/9PQuahNTAnY5jWfywH/QI0dpmMWgXcd6ZQyHiBAOXzQOr7d9CSAgUCyk0ysQImPt9PHDjQ03ZSS
bjGJeiZLKV6po+w1S6ufMxNRQCFdcObCKTvCtsH0zXH5FvEs0+jBpkUWvHVT+lClmLj7kRhCh9o/
Q/6TSQcBc6GpUl4KnefUo0C+hAWeOvABUieC1Xc0lmrslUmIprU/aGpHPbk7Pir4kwhmJxDU7eLW
4KdEVi+UN4EXj7m2yf8IufPBJKk6f6/pynY5dy8E24ijb+HvZLukFu/EAvSdeRpHwIK61vl8wWmX
h8HhFqHqAHXm7s8JXqSWiyiwha81HJlL4+JG5LuGFHKOLYq/jCWjrV5J3RqOqJI5WIWfxndwzuZl
Of5Zv8Q1R9YvsAevnWfW5UN2u5Hv+vPstI26/+fGlrECZ6frKBthSc+/rgkxh/19W54ctjvGWcoN
CWyixTClLKIUd/GR6rdcuW/BjTUeAhCfVH1/jZD867U9c8mYKRKkimXuznn9A8H7jjl9y3a+8eeq
Rk0dWMpFclrBhTXuo7EZkhOrlKU8o8AWYUgqpEuTYCLU6JaACFrhqUye/etThud8HWtPfjm1bCLf
mhw/t7gHC02zJWxpSGSy0uGEOvU/bWtC/buLeDynn7keM5QHk7EXs8CJrxmxYHT6TAiSlblfeflo
IB98Y9PseHPl5+N9iOEW8xmbAJ5w7yDgTEqrnrPn6bvmrYfQh6EzwdrpvGpSzWjnUv8ckmrU1Xo7
+/jd1z/Mk3dThQB5H6D+Y0KVByeuBXwOcLrZovTtVUdWdpnk0M3TUtEYPuM/zn+1AsBMwa4SgkTk
e9yHonUa5ByN/cQV71js1iaAl9D2pIp74BoFsB7MKZB8BsVT5rorZwURcFeD/eaJ3J2t4TxQcuya
OOob+4H63nIUG/RWn5ZmcfrxkWkqo6U7+C5/Ruf8fubDQXokS23uhwXJjaYogLDekHjUuwdy0VZi
XMpwOy7/AvtzC8NJGWHcqhA7kF/PdcKZ/wNocpXVvCYXnwKsaSf4pMsv6hgiQXByu44etP47P5y9
X2BA3cLBl0+cg178W5jAdkeNgIOj4AVMpOOJbH+14v5u49rx3A/HxZ0JU9dADNRvbfH8lO6iIo9I
ny8h+fA22nOJ2kLlgFUEe0FzCquQ9OHzFGgJkMJPRYxJALqVTxI7/GLN47DSriUj+Z2U7ANDuMS8
3cq8GC2Y+R3/zqm1bqcwn//spa5qMr98K6MymvcTVHHcDFsi56uGsQ/mlBZpkfum+XjRuTW61tSN
MZdUN2UhylOBuLboJ6K0pUFl8euMPcOtrBpK0khmPCEvHo7AWPkxDGL9J8VyaUwgvHU7bUiABZsW
U0yvJYjNVYX9Dy/U5+JpUVAyyV5TxCeIyNNXimnY4slLJq66+/DgzXIPkUWDoUon7A06X37g3iP3
yU+HK8LKBWczM3vcx2m9/ejEn9rIyQ+v6yqaW/XXGTrAR5HzMzbB72xH3XVNmP1g/ELmeCKzvVYQ
voc5ueTY8+bBonlABHP18ycbDjLUtm0rkUuvw6fzU1R9yKkhUhBY6wanqBE8KmNkwlFHMnC4Vple
d6xgdAUI7KmsinFqg7zqurUMpuZbigpQOY971e5xrjY8Qb2WhvPsRkwq39h54WRZvQ5dxszKA3eN
V9+ZTrWXB6IgeBCGBnL/JLx1yY4ZVXe2ZpPt1hjB2H9/Uum4cKazcRb9KC0hd+FBSh1Kbu+65OEx
O1HQIfex9K8ASxsBeiHMmx8LvgigxEu+LNlm8mtfWXqNeP+oOjiuL9FojsLiTbsHcpMLOum4FD8q
7qCbWJkNRl6Vlqwno6MP3litYII85N5Kj4mwbt/bh4hwYMWlWPNjQGKIOOxA2vp0lpAertZ+RX8R
HHKSuTDLzIs53BovNKPnV7mVea8pMaWhGICHf2Is1iSd/v4DO2rKODZxOcjNCJz+UsUTp6KXn9/e
K1f4ayY2OfOz3pWfRt9F/J5rEV/Oonzp0iKihUDrHudGk3t0QzpfrIyPw9gGw+eccNmGNvhTPDEm
2t930pQUjEJ5Py04QTQXEk7hb30ZZFY2E120JXVyZFjj7B3DemxP0RqmizFSG0viHzcjlBsfDBpv
DwwGJzeVcBN645RldWRVUldNo1dKxiyMLzbiSknrWXGi+Cq8IMFKXx0nnMJPNRFh8cNrvw0KNn/o
RBKXQF8qaCbZcUlN0sXH36hbD0EZo2aL9eTmV10WN5y7RZ/AZKD8qp21owgKLv516xILHBrnm2z5
+gVmeFITBlBbCsKlboVqziv1bag6HpQI8fMZkTYgiVEo8GzcAWO0OhIisxdPi065rG98vLD2rAYK
WBbQ7lvK/GGHtH1zHHBEUAgC+U2S2lcU7ULJDgWLxeeAEw+77hs8E6Sol+J6NjK1rIsE+wWe3eCc
hK2UyaHFH/MwAIi9UBXnblkKp4dycxqrjGUORnvLIUdMSsZJ3Mkrog8sfFDVUpvwf1yiJyZPZCQg
rakjBhRY2LObdHRKJt4tFwtRVeWxBvhCaj4bqMan2sXkg3a7i9HD8TZbP5knOXdjQ1OMy1LwGOPC
74DkSQGyB33ws55QGtuWi4NcVzQgkIo8JMC5Sie82FcLfdrpGekOXx4AAWvASeS6GdLJBgIlSYgt
i7qk7navvoBNIWXLNLAjJs4O+Zzw1BtCcRyptzIPcKsxRDhqQScRYqYKoiXdiPph7CAQ3//+1tP4
ejOwtL4dfUgJKwmoRA2uP67kQTvADfz3a+b2acJ+1077l5VlsldAyKisbA6HjSgunXsIsxje3YTy
HoQhMSq5p2Pdr5oq05WeQcJZ51Gd69NZcBZVNXKUN4h4H96W6QIVWYhMyXNO+16ma3LwHJRpo1Kw
1k5FVQJ4aRgAUxBKhZzIZpv2J0A6IT/zXx5InU5BLAKxA1hY2ztlHLLSLBbMgFoCn2SbjEMnw1St
H8n7ba5Vwtgk9SguoS2+EY0wOihdkh9UWDdPIpPK/Rvpla4rjVUsV26cO1pYMQ0DkYYrMBaXYscc
a+V0rpzHq52r06vDiJlxRdQhUQowJVhy+95YtiB3zh2+dBdNxgEnyEnlKZLRLj5PK5OQCZrMNgrW
5GMEm/imSptbkA5Olfuplw78CXNykqAtow6DUqq3pxf97pLFGfY3uBAytxGMb7NvScxzuF17s+//
3P80i0P3kHaCQu1b0dZtb+xCcZg80QxNlRTLv8gfjHSbHLEaVYrfxakHVeS2PBmSBTMsiwvx3TNX
Qemo6pz2F75j6VUfLd5c+v3I7TZXJORtGFhHG+eKq1CQGZexPsDpM15kqYksHDTNOCeBU+r8P8yG
233PEzMaf0Har76XzFXNC09oCo77A2KwIB28m2hg9aNrMfNhVewwHgZJ6LzcfMOVvCY/4ApujiHK
XTwsArzI8F9Ec2O5tGUC8Y+DSzejvOVyAuDleeR1E7fgMVnIJoAbudIDyKZ2xaMMTERecIhAtVBd
PnDjW4lrM3oHazS39bqFMuXXH5XCHuko9dwUddKSZVTAjzAykXwOkjMY5F0wB7LlAI/fnHHfLhYV
8SraioehgHVcq41TvDBteqkaoPe8YQNVnJZCocRGUa6g57WWJDPq14KYIzZXnKfxv7wIukCrsXTr
VyvlnIiDROLKK3oSyfpu/uZqwCeLAg/FRCYtlW426wXVJWwWafQTR1ao660gNG9feLVKk1pg9UnO
nSH+ZDxvWedoZDuSe9RtCh+Z49mz7JcRO9vxaVXYqnF+AQtbY3jw5lsC7xeSzmngdSZFs0411Lz6
ec7tFCRUFOSqQsQxkugtMqUDVVmADwS91XqOJENDsdefj289XtKBu4hBTnSKqBy54PXNH3WG+pIi
lkoLvc+YA1y0XgZ66B2/mz9HnR/wl8NqEidnuwlrf1pI0zPvMKMqrWf8UgYF8lpMgIocJ0tksTMW
PYQdV/LqByGz72OIbdZmmaxtKRrWSAApFdok/R47GgRarWPhWl3xzQJ57UbGQ9zarV+pTE7e8wGv
/Hc4/oYoX96xH4xIcOVmokgsCSKasnGPxsdCvwrdO5JswniOSHwJw+KCZwSXIWG1zO1u7gx/sdNr
baZ6zIeNpQHh0tKr10C+ea7SsdioFcYFPzEsu/V2ELqX58chYahQEcGL/e2WMdYRBhtnKfWhvmjm
W9FUwm8ktrIPdH9PyXSLsMnoJjMjfq/b1L7oQ6lhRlrAZb0rR+kedCfvNM/Skk5QjmkPk9UA0/QS
tc2F7tLzV06vaFIyV1aSUxuKAWhBvbvTAXp5Uk4rQO45g9G17V2UWG0LNwd5y8NHBNv6xHRuuqjY
OAmuTBiJ7F2zDhoFeLM8O7JSriStTPlxEOskp8eQ9WKJOqGtrfEW30MOZMwtbU+ny8BS3q/1QmG3
ZqpbsrtInyCzeSkDK9PbILUUxTa//qSZREcBAC4/4OooMkFva7FG5YnRGWtd6Lv9CyJT8LcJ/D5p
XldQstP37ahpJ6RcZ0Wqbr/omE3mh8S+DY9EB1C7IeMyioSEtkzSMRDxDrj4DL1nv1mYhjqI3jXq
haP0+pf/RvmJIXMu86IZKAqmC5uhNgLp5h3KCHTUUyba7/mEjClLBt/P3JIraMZ0EoRZJtG+NPXj
ugOPq32E9Sn/Q3j/4/2qDiQ1mXQD9a8YPDftJ43kj2P3kvjC0Tgte+KxnFfYWwk5gIAh6jIP/iqk
X5xFGsfMUr81psvpY2lmMQC5LOU84DoOlWAmsN6HRpv7HjwPxFXWpKP0dPS5Z0NOg+VXvHtvvoMC
ly0OZwajxLJf9BoDwI/GtFfJWqE064d3NWOmkAVCHs9OAu+TDAOlwiAVC1tJ/7Vxl+hRjSaY3V66
QMUCGtH7x3KBRhNTioPHuDFWgjxgSYiC2bzXMXXE1veqibZTh/Bpz2rrQYU6O4WeyhlxS01xuyE1
QJ0XznWtS35fk/NxuaSWf5+NHthHWb6siWtLNbP0ut1sqtQtH0s4gbncf7XNrTiuRrI04TJfIGUx
734Vo9WR27PrxYZvZ/PvbWLqm6dmzuAUJF0S/I1gYhI7QenhQK1/kj7DX+jyGNoWKnShza1jWf9o
u3Y2oc3s4DpMQShPn101TZ+8TY+aUx69t8rZBbghRupSztGy0IisbkKIMamVgrkwtKG/hMZ6Og10
3Hsm0SDlscx7m42n9GFfXAJFJBNBO7ZWsUpzEOiTLXkgVwGW271mL+qJQMbjidawJZJeD49VqQAo
ub7A4D6dKBhN0Hqf8yMTfN/16tiLcdAsC9hK8scq50kaxrKviTkDvv35zR5a5WDwFtcOseEbZuTe
Rbrw3MMRCj5DupG5E7pQ5z0Xe/wFqVPwrxuOtSbkgSfQi7BYSLAuvV5tHr7M5baUi81rXIuUPdPs
+mw2z61z2U6CUs65RaDWJIm040/HkyuxfpuB+7aTCjMHlS4mxr0GeIbPloCUOQVv24GNBSKcFz3A
4bvfzcyTvbq199592kr7UNAhEndsFOIcTSctFw72xaIg4z0tpabpfZrHBHKYfmzm6BVC1iWTY0SY
waYUj6F7UcSqch7varo/98GUBJ779mOKiduGkZUvT//OlZVKL5CqQOghFjDjxKk4s4lKqtXmIwUG
mnurjD3PJNnmEPiND+x7FZqljiLHOcuKVh161Ot9cqYRclLIzKPgS2bXr/OQmKvQNAKynAGSr9tr
sjAZnrWf2yJCuiEeLsrM+9nEheDY3PfFqVsqw0igt4kXVnQRKMc8LutX+FJwh+b9NL+vgYhJSitI
S1idkwBdjrDwB5lPnhfDnNbeWn0s6vUuNWT3eCZdnhanbiLfQdEyPslYz5wQGpzeDmdH9ILc3ul6
5LLG1/qyOrQO3y7nE4OswnWWSzG3AR3BRlfoFlQtgTdEji6ATI01NKWTasx/PXkb7BWtgbcMQnW6
It+ZalhxF8WdmlxEcpy4xAy6wVpDauuEbmQxb8wTbcgZ2pqQGm2JcelYm1HPe9dQz6NVKn1p7BWn
hXulDZia0C4vNESLSNvOQWGX1KGYtF0y2F7sgoJHjPLH3IEPDcweziG0RdZYYM8K49E7aTTs7DiL
L4nAKp0RW4kWBsPAdzo9pqgCnMrc8KPoBvQbO1P1UTFI/kPeNV0bsQ2+DQbBhQLwvPVi/cbEUqUM
eUuk3vfQMOUyHe4OYEQVEiH9NMnuFZmcfe8l/wB1U29wb/ypBYontQWWE/dgTaoqK57GK4KtUJEV
nyHCWYKB6sltHaeQUnh5ZZWAAcVjhG7yuIdXbFmPRmw4q7IW60KR56clRNQSVTKp1ynXX/+iG4S1
SKuvW/7zX9kMMausGicxLvzRCkYiuilHE2EEyDU7qAJRxsT90FGwgaSeJigAkIt8BJ7kN9zfb7U4
owuAPfRFKB+YJZAM0pGX+H2Rxg33O3ws2V/QPMlnfgz+dXM+Xt2mhWLl9XlkzMytY0uJ3BeoICBM
lCQNsnYGJad1CLQ42nvwrwHmyurd0GTmCsHKz94pSE0h+SJsPH5oUtgwHo1v7OqxnZnIvk+F48yp
3Q6kPzLGsfsNyALaS491Eg052+TOChYCs3+loQiWqLjC7N3ZQa9u7jyaUv3o0YKxFGmnNMv5MfF8
YvNdW6zCmrQ5gV7igZOdBSkXrM62KXJqQlUc5hhFAlVv4uZw/S6Ab+BMAFj8HurHuB4=
`protect end_protected
