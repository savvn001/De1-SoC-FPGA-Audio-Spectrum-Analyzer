��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	����_��� �K!���w��}p,���x����嬄��m݇1�����Ww���������WR~^�ÿ����_m$<�)y{µ�	4B%��i�660��?g�Ac$s�k�tP�U�װƆ�t�;q'��˙^��<l���
�"���n��w����|UhzX)���YoW(��d�چ�֟�Һ�d�����@��v�-/�)�`�@�<a\X4�Gw\UC�������*�g�"�E��h�#�=Lu��-$XF�!������WmU�j{�������uM�2ߒL�/�D�����"_���G��Ȍ_ͮs7��w	V�x}��c�	Q��?�E�1�A��!~E�0���Ҳp��1���^������,$'�a�7Sk�@�L�J��(̟��
q�>���I�ݙ���(�j�**�|�����%k	�X��d5�R��ocmh�Mүp֕��6]O�hk�����ЕB�tӬ��¬�n�MX�*c�7���QrCK`	�@+o�tV�dբ.��,��Z�1��J�p��dh��I�̡i|��,�y����2uA����D�ϛ�0;�ׇ	r\)�l��=��C��>R\"4��S�NB%D<l���_��G�Dҥ�y��p*�;W�Я��>���cy��zBX,��<t9auۭlfeZo|@����2���fs���^gw�2�|!�o��&#0�pg�qf_�O�/�&,�o᭰6~�b�5ETķ?_Ãֽ{��,~��{Aq$)b�>�Y+[>�e�JP�81���&�8h�N�<��-���ԡIP��V�ڲ[���r|�2��1�l/D�+ǳ��J�l�Gp��6	H�u#�����H�僸��T�4��a��*��R��Q��Ziw��i���M���������8�� �`4�[�I_k
H5�C+u�e��P4��hK��D��AՉFi-S�"n���������ɉ���&�4�J��^_�%�#�}��{�{|������!��?o��NX��C~\�J(CWd�����W��-E��kv�nY���LY� ��30�ws�����_�X_�`��l��w��)xMK��@��0�N��_٣����OF�dn1<��{;�T�U�' ����jqY�p��q\N�AЦa�A�¡8��`��7m?"��S����~G/G����S�$Z��h_v��{�~�ԕ�;��t�F߲�CH��yj���`4�l��ц�K���_�}�M�~�.����>��r!¸���֮F0�u6O�x��寪�*1�:F�g��鲲i��3����$��#�?���r�"aV�";�V2."o��b���c:-F��TF���D�h6�<�����rТ�i1�E��j��N�Û#��j���i^��wJ����i��a+"J��w�:�̊��"����~�#��{�����·�!mi��I^��Ї7�!�p��v�8�����J7A���a��Ptli0��E:�	l�j�J�6ݥ��y��.S�~���z�Vd�ʾ�2'ϨҴ��7W�.��pᴁ�$�j���]l��o���n�o+�r��c�T�o~�=�o�l����仓�ӥ��vj�Dw�����o#��|��!Å���	�O��e�$�K2g3��9�1�H�,��ia|ư������ɿ�������g?5T
5���%������;�Z�NVs�`��-K�H���$ ���w]��,����e͂����Ѵ?0�� ه�B�s��v��p��=�/�����,p� 2����.��<u�m^w"r쮖�k��#�|��h����f��}��7%\�d�O�(UY�s,���i؛MLf�z)��\5��J��D�9�-/�e��ŭR��<<������-�1�Yt�rs5�:|�se�D�߉�
Z��D�����аH�[2O���.p�ݛ�}æ���s�G��'>��\�ܖ��9a����|��K�D�H����g�@�[�7���W�>Η���V��6�W�!�Zt�[��\в�%�� ��;��+�[�����`? <t� FYn��s�N��[q;���#U�.;�K��n����av�D��.�D�����9����RX|�Vqtq�MgQ���>�nKtR/*q�3�t����)���M���2:��x�T-�#�K|5�%����w��D�(�/3��&��1'��q8\�Ұ���J^�M����.���u�9-uE
����|�,�݋�h� e+D�y���F�p��.H���}�O	���2�=�
ʙ��}h���'=��[�e���քQ{����Bj�ϵ��PD��
�+3C�
,�iaj�+�xk�#ʞf��R��7�;�����f�7"��8����n���UL���Q/���/�����n��X�����C��Ti�8���F(�U�%W��S�5�\q:F�>[�:�߲�)�XT�bW0�W^��0��O5M�ܵǮEa@X��(��%��-�Cl ���k/�<U<�%��_+x�}�;��Ve����0�_ݫ�?0�L�D�H(��Z�_��Q��b2&.G���K�����q3�.cT@��{).D����C`�G|�;2}����
�TAx6K+�Y�1ظ8E���5��޲�Z�=�	~G+g����
Q	�0 ��H���噔������s���ZF�Rb�4P�t47�8<��7s�ޘ��5qq�h�7=��ſ��B��r̚kZ����O��Q=٤�<BɥG�z��:�#B�z�9'%<��H�v̲�=��u	jnב��ODx����2�3L�_�"�ǻT-�{�yՏ�l��nu�5/���q�^-1%�m�*+iR��Rm��|����K�oBf�x�di��qk;���b��1��0��˙�J5�|�}DϮ�x$���&.qO����/V�n��)��F��ׄ+T#1x���2�%?�N�-]�O�q6�S���R4��N�#�u��[��DT��+v"���/�k�xtZ��b��K��HGr�c��S{���B{IKs��=�]�ֶ����`g�7<F#���^$c�^ɰ�и�]6#T�����iV-��۳�.�/ov�vY��riV%�7�?;g�����8i�m��
ؕb9/񇯮��)���L���s�+��C2�um�N6��#�����H(�4:u�ה��^]���y:�1Lg!&Ÿ����Ș���jP�zp�t{w �#�"v;֦6U�DY���=ӛ,�Tx,_���ӹh�$�/e���N�S��%�G:��F��Xf�p_9���H�Ɗ��W,�ɡK�pk��2���0-��\�g��^��I��|Y��pU
ާ�qz�$���>�0��`��V8�)�f���ު�Ge��%R7�T>&h��r��gT�L2*�g��^5�,?]M�ʮA�ˎ_`�`������.B�@e�v�ĉ62����֏��B;Q�'%�V�N���	��4�7f��
T�f�@�&��g[��|6���'�s�Ur֬��)���֞
5;G��yy���K���M�.�������z���������%v��x5�IFQ�nڅ��Ĭ�16�L�<�ҟ�a�
R���VpҠO�yY��tF���8�c������;K
W�rp��v��D�3�o����E��\4nZ�sg|JX��+��'�_��K�l��7^R�O�R���w<L�S��#UP�	�w����M?�L�~�u����=��uO�x9D!r�}nʮ2�1��I�|��iq��[qex�}���;Q&��N�ӣ���G��f��Oc���@�Ӡ���~u��9j�v�Z%W��
&q�z�t����崡�2�sB S��g!2��xb�0l��X�|��\V�ۋ�z]�n���*n��e#ܛm_N�\�V��4M�C�~�B��v�g����A���y�==��<�����u�����N�Nt����}�;��!���l�f`�z��}���_m�n���Zi�[���]����BU�K���r�[�����iQ&��=ǐ��F������Xd����8�P^-���\{�:f-\з���!J��1�8S7S�XUd_Kd�Y we�C����:~�	z%V��)h�ԽxG;o�R�g���Δ��>�OpWN�h7��Bb�@��%om5�z��a��"dFk��Du���+&~gM�D��<�	�Dj��ꥸ�%}q��������[����VX͸�Htt|��y����C_1��(Z����p�h�wm��$^���K�,�lk��^�*��ڏ;�K�8Z^F�%�������
w��g{2����e��T[&v��%���q��ЯY� dDu1�5�苭���h�
�(qI��m�iMxN|WFJMJ׹_3@�+�UO�:�&�+��D*�2�/���H֝#�����6�I��Y��̿���jE�ǣ�'V%� �#m%9uٖ�5E��^��J��<�F����q�����n�Lv&&���j��0q_y���U3�0~ @�;�>��O �s��և��~^6�������j#�:��M2�)��X��Yfq���r�Ax�_!��]|��I�&f-l'�\E�p��A�{W���Q�Uj4�S�e�}��(�hك�6_w!az�k�"l��h�B~Ke��n5^�-휪«�`����(��L���,7*�Hy�a�S�i	��>��|���12�����C�B�C >0%�GFB&�2�ݘ�$?L[I�k<���=�����^q$L�]�C��(Ų$T�[y��W;�n�2�J�����q�\�����HĽ��>���2o�H�,���c�)�I^b >\�<���1�_��\��أ��t�)���7����Q��|�uJR�L2o�E������/����H� �ï�����;�L�c��%?~�@�8>���	&zL�upL�Ny}%��E;���1;�<3"��`I��6V$UB"�q�z� �y�yy�!Y*��ʬ�\(;%V���s��N