-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
je/Kck7imyISb9xHaTBdop/NENclW1MyhtcuTCvIGPodkC7bOaIFMrKdt0j6+ecup0YM/GeYwAkg
VusZVGDCpvmqLG2KhvT5uhWZRqBQEGzSOtE10z3rhRtdLYV6xhwLXeRGyJST22QrcQi48/55UUcY
bk4G6268bE39qsTivo0A2vP5NJUCRTsTXgrQQ2XWh4m6+3Lq/756Veh2apXvtNthOsFkb7v5WvjA
lFFuCsINCdKpt7YJxA/okilpO00OnbY3/6TgX6ASHCWxZANtUZpaQWf45U70Ck8s/S0yYZDJwd8O
xzPWAdiL98dTGJwvDKMRQZ8VVJQr6J//lE1IGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
NRP9qhoTUPqx4QsE7DEb1xG4/e+gOnG244fIMRS3eJsOBJV2/0jlXkR22AUlG+XWMeZLG8OPln1T
hTyXV+ld0TRYOXv5S3r7CRF9Wvw1DPGbBjA7WgNjfdr5vPo158tRlLu7UANBzuBzcI4XnfSh3MQO
wNN6aPQ43Q+nOvApjNFlw/UbAPln8lmU9rPIfQJC6Am+KlmXCTBel7USJXmiUW7v79Rkt1t3kTV9
oXgDz9mZD0vMF3PwbUkLGrEQUzXsdoKFNvHRKg4Obhtl5qvc0Ipxfp88f/HoCsnD/hp0fLZsJOVc
I0yM2voP7JBCEsAlJvH8hZasqd8kiOg1uaUL8x2fOcssEgs2YfeB5KAetd4roU5gh9LTeDFI6ftO
N+YAbMEPfSB72K/vWRa6KZRX5oG8uAsf/ESoXmDM/MoeQWan6DK0s5ErR6qDuYlNZN3xA2nS4NBe
C4oBJ386v85rEgOMmudYSOe7yqJ2uImyrLfA9ETaId8d2KJjepUPacuPlEiIP/rnQQiixRwYyG3c
83l1DRFw/RU09j65jgWT0H+6PeDzeYX0575fic3uTELninKgaDo8Qw0zmFLNI3J6IQb08irBBzX6
5PzHZAxvZlRYKmrxoo+LzDLLDFkdoK64LNbn2zt9B0Vz1f5sl0zVwR+ZptLH3TOq5xAM3ObKwgmL
1XO97pZKUreV05YKfbQTs+O3zdLJc7xX1HpyM7oNYtT2JQUWmwuAZ9PQ6DwVscUOr95hKTc2RHkm
fH08gBhsRl81JkJUAsuCNYbToBkQ92cnexXMCxvFt20VUAaWl86tTD6AxjMBWWRuMn+AxKgvKZwh
5a1lc3Z1/hWDUQ0vWJf0q/+OXiIkc0vTHGAiFCaeLPPFrjAVBYaV8bK4aFELJHwZvFfuCzGGpGdL
ReVdOiQFDU+ZBwnJHNZ52yzI1kRPzxbX/hNKoP/uyn9AgjP+AocbE4ocSSCarbfYGIBCnmIafkrO
zRHnpWmfECdFVPN9EnPiu1hcLP4iCAgYUuxko8RBhkkIqQNhBdtKhQXIiWSrRaMsf4Pa8cRrQMSo
z4RVQv3/oDnhJcsmqHKu0MJlqgICEJmUOFvXBSkiQq/qNqxD6xu7ornEkUooTE0WhmIISf1hW608
mSmCqrJLh5kxTQuVp9ifzB1rhBSj8l33Zcp0LmYH23ifPUstfEou6Cr8uQGIJH78CnwmsAzaHQN4
JyGFcAjMhK3/Rf8JhOvxZcVP0F9+XQoH7xZJDsJl8rPny2mK87DADvCT0gdUT/CuD6kp0Yi5y96b
/pSOivFHRyJeGgKCrn/6NuvtGfJ725OFl6K4cYKz862Yxh0TpwjqB0fg88Evkls5DHZh0Luwha6T
HudOXNHpFc8B+7CiCHkaWgz/VZiVmAu49lpH40/3DZrkvLXe2iVJevkbZd0wGf7/wlFnGrMHY6D5
CFOcv9vC3xtiQCnv85PQ2Ft7V5rCL4eaYXXu6Q3Vv5bRjwlcjmnlmh8o0wdvB3eEjsIU37e8cxBD
i0YqpN+bG764jNbBgBR/ZIrfOc7vg0v/6XaJon1s521j7pNFAj1O/03bvCQue/5zs8ou8uBMqhWE
nAEAKkRTn5xv4CYfo4e0sRDw9R4x34feDMLCgsVdvI2JsAabc7UO4akeA6bjXTSTmcfFnnHGq0Ne
q7iMFPA5gy5xosHAPA2XwnJtorzEni5jfs5Brv527DVZ6i0xFwLVVF+Hcur0A3+m30acoLUqiFF+
8khMvi8coXgkxIzgFiYFIjri5301WOVcfKCawkHmCQUt4qwztyefuA1WiG35IlEc8DMmpqzXpKHM
ETsnZIo63qTPIQlDsF9QU0XpC+OZ1MjcGQYyn8TygIO7+67rgt/XzPVDw2H8R5BmIAI6hZ9edjaE
v1Gkl227yBD1h5ZmFO5hX+eR+FhHwIzeT8AX0H1+o0vqZOPlmoIjK+9+4pc3V8+DoonO0qLD3VRr
giMCP6Gt7z4sktjHWe0tdZdjLCuBS1lzZlO1GO4q3Q9NKcyLUAzMRRgl634a1/NXsCNf5oEY3/2U
/6VrBmjDVUrHKieFGsmbmwng4WcXXm7ULmgyEorQx/Jh1m3MQsXZPUGlRPRmGswHBV5AJ5axDDTQ
WXByeSi5VshBoIy77blNjhV+Hj41l4jTAOoAhESjcnAzk+QMIOnACJOsWGvRNZHOoS354Tr2jqHN
P85/5llFNsSaJh+EhKiaa8Ya1AnZUDMeTUz8r0xoXmT4PXMYD/ABzfVwcwax505ssejODlvzmwSs
Od0Lj90Rr6Am+zxjfXZx7Avws7eipcBHl1nOnJ2hD16bQaO+uWmevoitM2443e+NLqutGpw8kY2j
yixIVNhXUvAU++fceifB16tnkSW+7h22j8Y16xMgDLer16aMo/Dg6M+KxxjYTv7AweuBXmcKqjdw
QFRThCgpusNaLqEuw7YvprVNhjmz4PBN5V3L9GTNJcvC23/TYICTyHXqvRqiYnRxeSYP7u9iOqHZ
JMBEbFQwpqIaFeP8jqrsI+TdWH5CEvD5/i8+Q+7rNVNBvcEqxJ5HDX+q2MvQGRpVHBkMyKintPtQ
bqawg77P1GIuBvbcQL+LVS/m1262Zbi9z7dekgjEg2qp0NDg4ZvikJOjMfawkp1QMTJWRC4oeWI7
WEPGCxQeeGS0EP10BxUmk9qYx+EoXMXOmPSv9cJWj2cCZG5PJhHfDcwptO6kdlS/kiWOhaNUxgf0
iq59RD7n1sUTwTvhVZO+IWyC0FfRcDXq/QjhsAc2Dt8F/F7HFVF2IUCQXn0RFnVQ+JE7nyv8kYvp
HOxDpXWD+CPJvE32VIDbiWrCcx9FjtqUDhR2dnRlyvjDAgl+LSGwQDNvn8PkpYD2A1KlXmy2oJoG
VSiDFU8MjiBDE13Djuv4bsNU/7GD27I4L9/uUVFK2D/n4GvWT7v9D44Bt8sqdr7IdJT8YFA1n3E3
Qt6vRnPrC5QrMtK247gyVob4DRPTXOs1QR8fgNdtDCOZRiCt8idiuju7gEdTSKkfJ21l+cnHNMMm
/nDTtUz9XV4HhGds4c7E3MmErAXN0N9jtg8PmKqRMCVGh2fcNMoLyvu/gLqQRsP3VSdEcqGxp4bB
hJ9ivwF814h9sMYgHfXV/qb2da6e1y8UKFLZIRdi0SbYnRU5ogZAaF7JYT2eAezF4uvKDl/pkHW2
nT5APQI6tjSgkLIvq8Zhbkxb8hD0LJjI9CTQBxXRzNyrvLnPk8eBcNgwDoLDuemZtXL5+elthX4w
rwuYu7fnIgdKrhcThy3hXUTnnDfcuopPC4jgB3LGrfZSqcnxPARGRpaPN31HUoP0wmo45U0S1jDg
yBrjc92CwdGl62msxXPWzEYcijWeNDcju+N/iRrQ63lx4F+XwKks2Vry1Q4yBfAcL5W4HieFzxPJ
CZeBhwqas9F8yajiljp+L7wfN45D6pzh4Kp3WCg5XLoyfA4snMNhPK6D1wMkoiP9dDRWVnJUsAqB
TmT6HoOkFDnZ0RA/rOMM5D44IOTFtyvIJe/YfrwOz24JaPtKhBk/eZ1mXg2PeYluYirL9jmMaRtP
fZuyQ8kn/js1zwjP0mhp3iZXNWyA3pxkwJi7qfKiB4t+eL1/0JUwq7lnqGBJi7FniPOy1exisEQ8
4GdikDejv5FAG8GLt/lP5tk0CJuEJN6w3JfKi4gm8Ep5T5XE7IdTFQXBrgU+1DM72zNpWY7w3o7Y
7yH0g5YkaWcqNguAOZ6bKYg6hO4R7sZdaXx9okHWZZ7FIjIIolFITS6qJDiK6e4VDxLqfgsD3+Uf
9yy80YTxkyGLpkGrvsyXDbTj5ZLuNwbhJuGSB2zKDb/bkKHEcUPPu8EOwQIyDSFpdWipkMPRcXK9
pc5LlZ9s4NdhcyIsx01SOlmg9zwEQnGhbMqRRW6s9R6ULDZkLWLYP40hygr7jnSEJbBCPdCa48cH
KR2dK/VmgdvpikpgIc3PsrwOfHvtzn16F9ZjJC/5ncs0cqttixGfyqQzIgr6/S6HGr2gyEvxXZax
RyTcSWUooYwGSCbKVbycl1Qvyu7MUTgBRylhtlKPiEiRKwBVnLOaVGdyuQ/yN6g8dzcBdxO+yLHg
EL2Sl6t4sWyWSceKSbfU6ow2m4cSOyMMlPY/j26JARTU4tUlnETpaXavogLLfkFrrnDtsqw6WZUb
v0hA0y8PF0xV5egu77V59Y0jhdOjguSsDcw7tai2NPoR6SSaQ/cYq+do1cBDMWCBatRUi+MtX3tq
WUrUMt272liS7V6x1cCl32wDBeypWiRNtlQ0RlXnQdaN/N1I12LE4k5iu1l4FQ+xazlW/7v8Gaub
93J1T22L0JAcAG3ndCsoWLc/TL6lTX+e+YsLit+AYPBKb7IoMaqKTbsrO6OpR9LBv4wnOIB34ciM
SbUiTr8vtHSA9fZTFxkRRJEe2kKbM4IFrP6NCi8CpDNuZkD36epHIRG6a3QI48R+FjgRbfSxp3h1
jw9Qla2tOqIx8Ch8afhoTc41WwvS4mW4TviSAnctwh+qHyc9Poz/ec8JtgM65W1+GSvh7KTAML6P
GMhpLGo3G5GgK41Mrp6aAy6DNDkE0yE6MeHhMUZ0hSb8vPX1vKAyLAdfWh1k1o8mOqIkItjgbp15
Q4K5R6EHtLQL5mWPZ0jeEhyKyAAlyV1wXoCFLt27hTM328M8r375wwz0aXXL/eOWC3P0oEWW4acu
tT0ApXziKvm0Yd2zIoXznaqHjUBv/jxDy85+rC1Orn0DWPujzJK9DPmv7K7j88QFf5yi7CT6kkXH
K5NOozF2xWOWUl3erP1Py4Xq2k/zbnEW3rl7Faodj8pREJ1+6nJjx8zuXeNohbRYnz4nlzEj+MfE
tNZ7RYp5Xj2r+FWJyT6gdTta/J+ijo2ZVyqJKfCts7Pfd4pq27XSnoPYe6bU6xq3GPyvp9Bb7ZyZ
1ndRIihnKJDIpWWvQCYx1wHfPnfWFN/nj/AEInEh9pqDeiDtyuCN+tHpl6WRjYv7wCxZIsRbLHSP
tn9PVw7xE9h4sopb0VVdLv5QAiR0xgX9kXft6VyLfqVGgn882sRh4XP1K1y9n9giq2rfu/m+5AxP
ekTWCOXulIVnnhch7FaBhkLdjvv15t1XDi0dWQx+RkZ/nc/5jrM01LwTk5oSfVRy8xEYQWUeaPXH
k3Y4a6aEU5tt+t/4TRCx347WnvbLvnvOGCdjDCJgwn2IZg9V7sYmexfwl8iHxeUjfa1bX3J0MmwS
V2PazVR4qb6tBDeZCnSIoRZCbBMKS1mlhWa/grTEc+CK9lek1hInDzSoVutsfQsu+Z7STIkOYO13
LGncs+ck/G7esvWwPKT9zaTxrrUIrLW+pIPfWG5Zf7mVO6nuM7hlLN+sYv5rydTMRBBRgGaamdUB
Oun8IVEs19u0ne720jEHvPkuB4Pg3i5EBXbAKHTB8WeHSV0aa4v2IDd6zZMPOelYD/oquwI/Ac4o
edFx9SUWKohp3ibRqxR8CMf4hskN6WGIqBglxqBjPU4BxcwUZpnLs5SfJojiSBwFs+KoxALE1q58
4UNdYBplaQLqerj8wk+EkT9+wiBLbANlpLV1n9/n1wn0GvDgQgMrsBKEAVh8dBJhGXNTVZyGyj70
MX0UG5Qkufix+fBVhfDRrQ5jLYWdZyS18fffz/6LIR1YRll03Y6l1pZtXkzAT4uQBfzkbdiuSxKG
0I5iHDn7OchgtcbCNVW7pbqKo1B3hyAp4qJJeOEJbtXk2VAAtQrdOzATCEt2/dAhlhEkVoYu8OqR
XErNQe1VFdmecYcL7wzviSNwZ/C8OQeqOBdDkmHInhpPb3zYYdAWtbt8Ua35sM69BcC6U5p4vMNW
7m3FhmeYpPgKHJ1a3QSYmx/EgzJI4PGa+wqYUL8uRWfZGZ87lfLqWMkT/XKC1KU5LKOkeuM1r5lL
K83JGxoFo/qs8xBze1gtk/EsocE2tbrXP2S6vd3/kffv6+uPE72TI1CRm4D5JoFqQGgxY0MWQoyz
6rRjmnysqpgivEt1weZY+JiFiJRPu/zXVvyt3LW0lSlAJOm/nT1xtd0CA1sudlbzJ1VOWiByWnFD
WpKvjXn6NNL2HeowvYh9y1BtESbyyyBDN4WdykLwgjmPHFeWVMo+VyzhEGVD6zvQpD4+tZxQz21z
4u13Gb8A6jur2aqBijF3tvbQxDItQ3n/O3mDpaYEthZt4Kap8K91VnmefAUh+aGS9VAfjwuQW3X5
Rl6LlGs74F/MexpeDNDP4spB0YGDXM5VTH1G70LL36eW+sZblBxmTmJtTrasiNPnFWwwyc6aWZVS
K4MNgzSieekEwW96kMjsaPtRvcPJ/r55N/LMOL7XsYw2QYFcVcmId1YmSP2DsjRRLAZm2Ducj8A/
OT3Tz+spjSsbuaN9jvTTmse4z+TgbxzJAqYJwI/sBdK6IgEeojf278pwvI03iMJxaUzMMk1BMDNs
us6ScF5q758Eqlv2KcggJsP9luPf+dEuYLdleNaDL3w1TG+itZQV6UFGFz1w4glM3l1fn/ylnFzo
XOsWK01f2lcN5mnbnyHXKIK6mAHA8iLATb9m34a0gB6q0ikPfmfpSL9gSQUJvCOm5rx/iOwtmUev
GHf2P3NxhOl+0OFMk3Af70d4nU9Yi3Er4z/fP46NRi4afCxvsaqzWtxhPF6qIt2sGI8CwitdZMdM
iLy9ZEcYHLkXVlzvoCm04qy9szU4WDomMhoKzCv1PaNieKypV2P9tHpv40mpMXsrzaX0hy++pFjf
VZPh2KLauMHawbHwvsRumYkbkPYkZLS2CQ3VbQbDYBR/zNl4NBpENmJj/ixAqt5Z5D2y/BbBrtgr
bAACklCm32KG6N2j//Q3cHattIJ3b2RTNiFRWVH0dL/3bp6VBJeUD0Ryp4JwfPiAEYh9HR0OnePY
HcRMMxj9xGoP7PzRaPoVV6OsCpkHPL2LG/6+op8mpn+lD0rclFykcWK5UDfF76BMJyclQHYWUAD5
VF3B4VtIooYqQfsYHG5xInzOVo3WkKwHNMYxX+LvX4PJ55RZrrfpgTkjqBFwaqe3dmcYe5eFiHZI
7SS+Iu50iB/O7djvgM0d21L1OwhkCOYQ7bs8DcmCLDarASbQzzz3zD4yR6aQ0+PVwAkFndWgQqrV
TQZfxSNa3DYMxqVRJjvuxqFVcEHFLKsgqZ1IRqaBHAb1GuTXKp7SaYu9nSMxr3ZGVWtUgVqXOax1
zgNWg2Z49cqvP2wDDU3xYAnrrNuLsikf2WiZ5BJdAf5BGsgoN4kdHt8KfFgrIa3qMoFd6fXh4nDy
Inv6Q9ZlT2vmm4EiCwmGPpqzpucJljo8AP1Hai2QMTV4zgIbNrMzoEcwiYKgu1sTKvuUkdtE0RNK
R/3IVfIft0T/Sdz6n+BXKBooiDRbvVR0j6EJPzbYHxSXPLgBsrKMLlaxAyLs7cNJYNlY2O6H3t/H
HP3+9IOXmyWeOEKuXN0Zd5/wUYxp3wsb/+UWGrkRlMj3A/VNQl4KoxcNgG39lUz+StI/G/u49jS3
1iW/EuSL/mdVlqYQKKjiOwN18b+ZAZIJLZVFDlnxpqt8o+VmSxv6u0rMa7pXXnqNa0r4MTpKgwxF
Rmj3uqAC1/F7ZLA6WACts53a2HPY9Hmvr6Nh0LcWUitM4wquvIemt6k10WumNcK0Urud9oif5bGW
EfHedSdP/xoxly2aLvdV6nIRzW2Ol+FOauBENZE7pXMU8tAlsshxCStSwDbP1RPrgcOr9wgA4VzV
Lj2zzgxXDy42tREYaIkZHFwKqsUALJ5oN+OPbgrHo774ObuNpfhonI0eP7iVbAyGp/pFOi6PC/xa
O8tXvr9IT5GHZe10RkHtVJHlvr8gx4fZbo12DGalFCCzaI3r5pUU6ZUzdFDOx9668i7jUZYnLUn3
TGEqehPTkqFFI/PnoyH5wb9yboscGTsfYipgsmpLd1uwbXA3LrF9bDjEqLYoJC7alaTw6X95hPKY
MfB/C37nG32D4SJxtUNVzx4DdJTHY/C4eNwuHCOWak4cPdjpHy73AN+8T/0CDyeYKwanpTSdI4do
bBMEhmUUd/17Uf2gvmHBRv4jrEL/O39NEwUtamdmaActr1pVT470lF+1wC3zdQWY9ujiQviKpCMB
gBcgpXf3279CraCFm1QFH2NeNl/BQVTAAjkUPid1Yt09D40XeK3mUrrs/zDxH/OWiHLA4wmf//wU
CXZx7fRoHLgWC0ronb7PEXiKjPIEssw0rvb/tbpeFN8bCg5BoM3x6FNtpSHsP4wS9nxXXm7dDYUj
JrcdP4gZFiL7/RQCF8WZBdw/pdxml4CZQSxBaFun4KR0LAoznEQXJfFTDwzn6xnc4SvQx6jl4eLv
7mI77URSPfKiBdCiuX1F/Ufn5flof+pYkFoqW6jfGRFTN49jJvukXcrVnffFsfKbrFzMz3ngydWt
1eirJe6STGSW7oaLSM0GWrANp5HoLoGEAlNkFG7NYJMU9f4aBAKqe94a/iWyRXKEVHq9DbDOiIVv
VEYGUAutCz/QkQL4Tigfgjphn5oWyHe1QJaEMHJMqRHrw5aLZTbnKurPlTTze83YaCaCZC2Jyfiq
4R+VLRps9+u5gnOS55S5E9pcsx9+WbM8X8lwdz+NhvHefBPOTfbt/TCg2T/BnOB380vhA3sb0NCk
fUV3tNV3FYriJQQrYrmpEIMevPQdrlROIEGJmnGH4aCQuvXCGLt9I6RKqH5aQhcaMVM50xInVHW+
NDidqm8YDYU0F6jRtA85r4u+h0DNP0ajk7pjc8zFXvKHx3ROY6CnQEeK3w3qOzLkED8CtbwSp1xk
YAfT4ClFy7WWtv2MDB8IDBIuWJCAPLRZjG7ZXTYe0hhjnnykSyxrbhyyGkOakAECP238pcu5Pb8M
Kc9e0u3hX+xYyPuABrI6FtTp2QeERKrwbSmkwGllhfrSkHs26HohAlFywU2qUa6MTQhvAlciIR1y
8geo8nHKc/zUON7ci/weTBu3AJ5qQmlkJJXTket0Ym1lNhCPq8vQ0c4J7qln2X4Kt3XHupH+E83W
2Zf+Iihn0KFYuySTusZdVMmx4pXWCZst032fvIsuJbUCD6Byevp1Rjvo6UEpC8equCTtWob3iYj9
38fbEst2q2j1pggaI4MHvveH2N2aikkwWkbDSGFFiUwo9GelWhyJrhuTLac8LEXNgKT8MXKtN6oi
wSmHCeCRkwAwnqpfIbJ+4IXcMkVap+mz8k7Wc+UJFVetwLqHKTYHtb+ySK4iUQNRnrW0TwErC3Vd
mfF78u8eWALB8l9FVYa58Tdn1+cEMMCiJCeYWZQAcCOY0Tz/XTSgdsvefMHPB7AG5USyd3A+AhaN
aBCBaA4HhyyEjZ2tNVIZvrZQ4g9yChHTn3X/k56R6gUx3INGHDFEN57F1GbGaWB02bFz2Mz1kQS9
9y49iWPYR3bJJRxhwf7xckRTqra1D/frHpguponTB5RvHpd43bKtcQ1Br0Sg09AeTQZ9DxlTIpKK
DLNzXZrDkArFqr9IkFg8gIOQAgCgBqMu3UEc2yemdrick4y5dkDhaDkyXmgFPPC4UEInN6tSnnXF
4vGbyOQDKBq9uW3YNhUs5aR6ObcPmvq/pBkDPyusDmsE5tEz1cw8ryXB6+DwHQxxCZLQKP1ZTrdI
adtUpdmDqcqxfHCZft8zAM7X3hbX6zvuKfb0wJr0oEoe6peA+6RWkpoYD40CEd4CsBoPtE/zhNip
1FhgWQaSbFXhZmT7IMix4Z7b0JijMnL7tbkNPuuwQzgV2FS8ZzTl4FFu4s+JslhfwwwB78stSJ0p
y7Jdeswct5HxaMmFKwwE4Nf/QlQ4zNYyUsTu+nIBYHmGRLx/64DP7xyryJ7wRIbnu8KE/n2b3XNg
38iHQxu2GWAInpfCAhfSg8/E4NO/AwKjphDGCJr2JFfKt7bmtCH+8JlgwQjb417N5nCMhh7FnQF8
CXxBQbgK70HrC5zxXWe+c/BBuQA21u4oO2oBwkA10y2PJ2SG+aNARishL+aUk9EYslqcdcmUkZhu
DARXkBdRFjSgUxcPeJKzx6JwotR6wp560oD0yEjpvrXT/ZKAA/pd+gJ8aYCqGmB6gmVA6VL/jmBU
1D+Vx6jBg+BPb8FJMk7m7e0/feyqsdskDtI7/PSlRMYjcZ5JMNZDrU3nHXmRa9fDBqCkLohN1dDm
Cf1Lk0+O7/MlJ0sdSPjgR5KI79SEmpqd/gn8twvdIof20unZ/TnumBN81HtDhq+cCwt7WFr6Xg7z
ZHPiaCjvvktz5IpYepF1Qgc47V+i4T7y1+np0jmYpMqfEzePTtsbV1+AyguFx4cuG9nSHGGWNXFG
QrQEy9MsKXsxVnLgNy6wSXraEdEUgJO41AMnOcdJ46nnHTuDq/Ltl0a7EykYJNXWvIOHiw75xrMu
a9engDhb42gL6fULOUJEEEVHEaRLhj43tTSjJYcN79wyAvhN+oJXHAo2xmEwpXtpc9EnwYRmTgxT
bndQ37kF3hQmf5aCmjs3LZOJQe7bHiihqT5wne69i3j8tIhtVDirB1S+ihA0Ruh8WmfjcWsauGRd
ZUsiw3wMP9gEJjF5pdZYd90AxeI38GTaHFDyMrX06vqZEyLqGoORsJTo2vLV/2HxCFNQoLzvOLQW
QrQ0bvr6t/oGejw/qcpMvCMIPRBcnLtP7epKP/lkDPufeyukVZq9Oume69HHQfFrkiq/w8A3bDE1
7ixjHtUKoNJzwOQe0WulW6rWy8U4u1HaEliZHFK2rO4lUw6CKE2BZNrUE3lCfjFfLtvozwbnoWfX
dNfTA1zvfq0XfEIbsZdF5JOkEBFK+mAgDMDVqexKRDj6cS2bu0JmpzrZqylT5zY0yxsf5eq4KK3a
KmeqH54hQ/A3JYv4YyZZCoVo4ALfeF2fn+yQhDDBiPoI6y7nPMfQsY1j7zBdSmkx8kVY8THlcz6j
05526eqAR2MqJTBCkl2Ow+1n7DvYREDa3KQU43r0RsrPZFySM20SdekU8ytyNzut7wDy8K+byjOJ
WgdmH/WSYlFMr6I6fqUpTAyh+j+PTq7EWAVBv7ZwcQCYIOrTq8lmyy55q1/9COWlU+fKDaNt1jOM
GVdi3eALdhdHFkHtJ89xUWtSYLwDvMqMDARs07o6OapY8sDthEvqozom4PJGp0GtOlhzKEp+gZqP
qitrE7QWTg25BJhrFDXm3bX+lmItAANDPyHIFbEXIks3758FLtk5PBeTKfBeZ1DmbPHXj/zbUep8
lcdJ9g/bEhiZ27XzGV/b8TXXNtaKTpXccEocj5v6v2V2kKOm6SrodG2UVtMrDPMGLp8T1H64oyl+
Vx1U9iYXrNfdZbADXpiSuRO+o/Lk7nPwynI4tiAZ7iOUh3TBL5r4wJyQpI2VGl9QPQTHIcBHeul8
npb5kaejXPIyHfiydQq9l5TTGP7yss02rET+BUk2PEFQOgtbEw01eYXWzM7ogeWhZSOflXWHU/cd
zDbTHT9BDZDNj495XrY13h9dhLroE1mi+JwLNZU3zJse1ZiRcu14JiDso+XuzNK8PNFv/l1hg3fH
v4eKUmI2oTHHg6GKfgzgY+M+n/JmCCQah/0zvWfq+dBnxjUNHgjhg7SLTPocEUygeQo/SIrRZ3qh
jzc9Eo/ixthAEdHMi1jvML6oAtuIz34rfZB8qMivVfcANQwRHN3mLjCiyv/N9gqO5iXSXJBWU1sj
cryCP0ZkWVWbCPzR5EwQr2+UIt/EHM4UzdLRNqK32j8OZzSIxr+ERt1UDsF8uE/viiJoGwUrpGvT
qZNNpy+f7CiCr7ou6xNBP1A6YHwgS/gdRRnsujWV+nVqns30xZBPvInRsmp40Ujm/7zR0alYkK/G
uG6t8Pm8lrgBLnP3VN/1duBEs3qVsHxhT8nY4W+ML2SfUuJ8x7rMvauryUdX2FvdIH17xyIQ3guX
H5ms448oW6i3fZl/x+zEFAah+D/cTE+bmCYzyskAn36vpaCAst6eHt2YbOXNGJmbdR4DYB7vsBcf
jAuC4ni+J8dos6eRQ4FY0jEjxZvLH/Rt5D6s3thDriO6oQxSR/rOtiiL78OcUOV1oiMpMOE5ccKz
rwP1iD6yioOrQmwrQJABqdhrXj2xYW5/pRpi6f7tyP/CE56OmGq/kzB7CG8H/AXez9nX9NEEV+bY
KM4A0PGDxEsPGJZHBQUuSC3ihyJY9AjCj1imfTQCsgXwnWJVJ7D2RBD+YUzbXVHXicdHzHxkgP9P
5/7o8aDeoeMx3DprP+63zT4jNczZVFTTQjyPHbZWeeG4r7gzuPQipXGv0Jk3/v9esjdDG+MMJ75D
TBk3H17lLzgYVvvBHfXeaLGSZqAKHKbj/FJuiQRwDKeLYq6JRv5m9BD4sAmfjohJj03F0uxVQmVQ
FMdCIvCLojiy9uV04Cqb4PxVgqkhJOGLxClNAnVjE9O76Q58zBsQWZICUbNmYJZDoAwYu8+9uQnt
bb8nFSWCNduDVRGde+j8P6brGBAJfx4ccqlLIFsMuQMPJJw2aamDhsXr8x/N1F1AO92F+185VDMj
SwsTewomlxF0JORp3drleSqz6LwPQM+GVe6HL02os1ZN0sQACAWtQxJxJ2n3yUV87b0Gv5M1naDT
IqlJA2J44/Jr74pJiUxrhtIjYUriuCIz+oyRT8Mc8J6dFOgZHvew/8SDKtk5u0/hZVt/HUoIVb+r
jb+NjhfxJkuxEnAUOI5SUv7Clb9d5zRJhpokBjCauiiVOHqhRHeO2NciVjkDUFu+7pADhLfrmqi5
rE2Lt7iCNi7SaSeo6VNAAXEehrvJIniBt8NLnqTDlsGs0JhYWL4GsUUKye8X8IR1D2PwiRRIv4Pd
VPy8Ziw2q8UqpwUqSy1vg2pj2pLMNLgTfnKHb+Yra7j2z4sE1OBbmUrFgpt0Mx0sBDPtOBm7AGAY
bhA3f/JIHkyRWwDg/S2q11vFzFZRbKu+uTi7fi3cqmL1B3ZQlr9Cb0c25AAIPl3/YTKgMDgmmYJ5
cLbhgibcrHEIp0vA6PZdRrshoRXYlZNacYJuqH+Lgy+yumF1TDKjQVS2/PpQTj31clq25/E15BhH
m0Lxf25P5mELFqTbg9ViYFTYS8pcxkf30re1PHz28XIRZj/S2Jjy6D/8ThwRpDQqwkzyRP9X5wy9
QF+7wBHEtUBikd/zIoxsKcszs6+Fy4rTVHIPojkcWAFU3w0MDMkI36Iz9zkNlKvV05xfbKKQInqS
elVwn4izxzb/gB8IHcv7PEur6x8S9AtfippfrBRCpF06TxCnEzipThPcJfWDSj5BB21495cjaRzb
t5jDjAdP/zjXgvmth9QRgXExggRq2S8n81qauJ6qor1zUxIFjjHNcVIGGlVLkB4MxE/kudkDa8bx
P6B0bX7ZiT4XMlF0i3A6xFtWatmv4TwH7YmPRKXPau606I2b0vRdKrmZ5nXjp4Vw0VSej8caS/4a
dPkDf8UA2NTI3YCOBlSCd0wimKrT4VQ3LvWtktB79US6qYWGVrXuPjo/Wfdo8OUNNlim67fstJUq
HVeUOWL+aBP8i8WpltR3jAPVmOJlz5odow+IbiY4tEokGVJwRUVemcECSiQhd9ssUkAc20mr8E2u
KLg+N7IniPG+9Kzb/5iZ7ihWX2AkwpkIiAIliT1bv3zUMEl1Q14X+WWFTQL4eJevzu8RiTEyGnL3
qier7Wubbp+XeAyVyVqbUKOWFMglWil7gPUhRUUTLv0r3z0U4Pa9nHSjsqD2a7F5yQys4pMXoeSC
nty+CvN+JJerf9b7NptPF9EpgNV1Cp9U4VEXG3Zx5iMffrdmOF+Z5Oh1WSq01R8L1TD39u3UauI8
H7ggchKZAAqBXUDU/g7PR7aHuvlmJzNHt0SnCFqf7raQgIth/1GD4/uzPqa1XGIkd8QMryQLjlEe
JHH/rZlypWuXBeY059ZRrzML/BCvFtGc8nzjCYDy1l4ls2PQWKiH2tnO2MB3naqSU5mCe486Jubo
l6DEcyHEPGdXCysvxsEXj2Cd325RQaCaWBEl4olyjwM7aNynQtlKRI0ifnBUMqSvPqaYQ8aCiJQz
XPRCBaRa/WV1aoZxdro3DdncGPS2vu4pk5KvJA9w9TztILXc+ukw6jzuKtGkvcf+WghTt8dgUXIp
VsdF9CtL2KaFNYP0alPEdgOoD30Eu9oH68DifmV7Pp/GEO9Z43E9ClTBysp3LXqj0qv14b8ftuFZ
fbLhkh4X0aL4KrHISiTAkDLBjX+6aMjhyuW/rmMmp5YAi/n9C98YRruHDN6jIwbgYSmjn16lSaJi
XnQJ1o+dTV0TNXeSCO9j5lvVQNj/QOb+P/AXdCZGaqKL74qbdpElGT43S+B290ARnLSy6qboVi7i
RTa7Tu/RKSZvcn/pU8VoakV4JblyqIwLrwesl+mpbYl2+hSOwwsGy5WkASIhc6oohtK/No0w6x4G
6lin0JMWq728f4c9EfC6ZKJEy7/qS1pFM8KEjK9R8tD4LHs4Od6WkeWyKcVTv58tUcBuaMUssKxs
V9o0HbDnqLK76+2Fg/pgryFkX9ReAN4YdvrKZ8xyQbA4Xj0fGiQVkK+Ntd98B7XeLi/GmH3Ziy9n
+e0VSR2BlQoYBj6ycVvG81IUTo5F2fEOaXsL+YVsD+KygPCZ1EPPPGIEiUSUHx3aD716zhmhZ65V
KTmkrCSOWca1hBn2Or7pEcz++VqcP2JmZYdPmHuR9HrScgaDWo972PzzLLcH3OdkIHPvvNo1I2SL
zXHBuXYHBHgfFkagK+0gIAWmQ7t32UYWy640ma9STWVdjQUGwrUEZHVQmdqlUYDfv1EBO2UnETCe
0p+g5oyvz62+0cQBBR0CUrgZ4DKju5P3XfditMlmHO8h5Lhv33n2HFWofUhVdTPqZp6xDcikc5Wc
Wd+S6tp533vvMtUMfIJaIMRTNVvEkSeltPNIjEsABuehKSwkf/wkeGbrSHbaUwn6s47vmwirN17H
wTNCILfzRTkdcNJXO1rb1nPZHp7xNVGJwKLI6GXNnhqGDXfmMxqKjs7VmB5IJjvfw/EaZI9OrdLC
fnwcjScAR3xknvo5uj9rA7/EhPxAWiJnypt/zDxrtbx9dFbYB+Q9zQ0XUSVtHQzf9/6p5r3Kld7M
lo8zuNv3ooGuqqk/4ocrqNEAyzEL9n1BqUGRbEAXa4EA5BuPfTe96s4v8JinOzLMKRgD6/8R5GIx
5vwPbaOiRJVrFCe7zaJ01WIyQ/LXj2AeinSqtQ7prU7HfcibaMJw3Ww7MZrdVP76z326O0PCfXou
hwQSlUsCBzah7jn9DhPHnEtLVKDhQ3px8m+gtwKlOHa2v4QvBoy3D73BGtBA5EK/g+v215l5qh8v
xVepku+gZEWSOu86GaUCmwEDyOIqHQPGarri1Ypxsw+1AL3tdC/yVVubcbp41qGQxj00ZumWlk7s
mJTAcEJSCxgr2EFiE+lNl1xUcpRL/reaoQ/dpOzAF/hdSz3vtc78hKqGTJbdwD/NCehnfLgEm/su
PzHo2LmJUH18v5vjazOFrBX4Sxk+pPtrzKPnEjUVxGaVbZw3HG6L2HtU3v3ggXUQW4p24z2ZkgnH
G5e8bhXU+Q/OfrFgx+fGYMZNjhpoKb6C/EWw2kSouika6L3kz3jN7Kcz0flhFfLmCEf/2nYKjQ0t
n07c+KnuqhMMee/ERBllJBVZbYODPgV0/FvTodcqPbgegYTzC39AX84HBtCDIV7C7+kJRGiFz6HA
JhpDzNTsy1mZSXAJZk3Of0iqJY9dl66mdjdY3Rpgx5pQprCfI/s86ldNgvoWpYpp6KavjC65twiA
akH0pVgLHWGS6E+He2VOX2cS4A36+BQP7BHLdyn2OhI7TrsNgX6g9Pp/Agq2ftCAcLGLJ+OoinMM
lB21LCgdWnCQ2/Fb1kOxI+Ma7topbSJrqStyEN15iGZW8516vrG6BDVS1ITJueOh71sItkRpu8kc
/KjzKX58gpM9iIFFFfIqMGbozNPTl5KG3rF/PeW5T3+1jAomQFnJj+kNhJNMlNeV3H7BpWCyW6Oo
Rk+YaUjlKpCf+77ff5CLP/Dasw2PPdHDEbIuv2vbFG+/VlPrMTRVeiwTt0OV+eCSl9J3hgvWBlQM
a5TeLM/JrZ1FDqnaciAp5VPSrawzeQPvdEBlMuQFLH4IIlfGtiPgWbsqWFFoA7x67F5Osg9ljtDE
3P6dim8+GcYGUBAo5shvqpwEfzUAIh0iEK92uOWSdKyp6W+uJPfcHy+CyNAjSf7uCLhR+rhY5Qrd
b8WAtXOc7DkzRlw5wOyuoCGf7lCX4ROTGlBnpP+amDk8tA/wL1jvz1f9qkPfL2PSIbEDTEr/Va6j
6gXtRQ8PBeNxugp/F7+98n8u+ora6JtE4YmP9sKItu/PWfdoIVGUYh+jShEF9NCCjrXBe1ZTZaLD
lSYUtOazZISbgqJ2dOSV5BcgHNdmkdogcafLiYU4/SNLQ1x02oT5AJSP4shkYcI84uNaUEKcp1Tf
P2jujzexCPCtDWKowJiaHJQ1T6BqDnWh5Jh6ZwRkIA==
`protect end_protected
