-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NvW5KaYwwJSS+NApYg8lxCQhV5TMvfQTSlPMxDVVlMUEKCwHWu8jWy0bObSWVvdp2cwTHl4/4qjd
6Nu8aF4N2HLooWstIVX05+wtaFuC1gxCE3+Ldh+4TfQog/wT9Qa7IvN7XPEDKdOi2yAjmAqF+Sgk
Nr1PmLAJf2DIfYZi56MX9iPu42wbusHJsgrMi0GkQFwYcJiPkWQ02A/Tfn2wIVblPz950neW++HI
EhxfT+i8P6NcvPEX5L4TRmdUXn3oIUk5bJaNP4voSE/4cmhRkOUO/RXo3xaO3aIYmgjRzgjDYMzw
EPy7BC7gdrUc5yG3VtXGMVRVhpbf95wIi7JGNQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2960)
`protect data_block
4vCza3nsps/koBb8RwoaqsY24cKmmE4IOtum5eTztSc3MSO+JBUBZbIqNhMXkNdNSWh1yzu0wPs1
t9cbTgzyDwdEVFEhSNP449nStIRXGJzUaeYhKwNitCWV+KyJKnqYVmTpdIUFsDqiWeghO7CXSb09
mHYsP3c4F9sNk2mdMN9tT6u1uie3+aV5jpb4tdsEpMMmQxV6SysbzoQB4mJafc4RTlMSSXcsf6FI
qM0406/LQakYeBOVh0e8qkXr3Ny6tMdBW23VflHuFoU1FbRgAOl+tU49y8KO7qkR1K8dgkgCQJX2
FpJhC01p1bjjwih5GO7HF7dirYvyUAwye5Wqe0tDx4ri9m1Pzs58xYVO4bLpE8W8L4dgPq+mzQg6
5XAkHGXP+JgQ9xNbAuvQ3GYE3912qgByNksCBwAOrPmHmLnPjopWdbw2IJaHC3Q520CKbDilB/7n
BbvfmD+/TtI8m6p3KZvg4q15yxMJtnVRnrGghWsDuh3vHvkmCxmSJja1VmYGO/vhfz/idUVbOBOu
pjXoKjZy71ephOyZUOWt1DUJbrbL0kJujdd4WAnE49lEfJf8kKFImNePe24pzVJmdJYqrrbJPJTf
UOXciidiIQfUAt9TKpI4Tfq41W4uQR+wluxW/G6c11k8N45KzQKKmTucAZL5z4G/PGxL6dG3U13b
vtB3NyPt6ylRZOtsby6n1fTs2F/eI30RIgBdihArA2f2mnbEXD0+AKA4N0GdU93bQ5VHNV4RIJkf
anfQgMA++esYfwmY72C9m4dEgfpvGpQFC6nuk1QUW4gvF1PqgfS/RZyoj/GBYexFPb+OGazQeorc
M1sP/jmCh05ty/yYoMgwa5GSvCudeXyBMFaTNxMHNvHh3zMhHsxCHa+kGgu8Aws1Pw8ke1+MbjSS
snZbRKcVSy2VeBkiemKgFH5JChCOBgfC9UgJuDGHrOfPbz5hqo0J7yfFf0+xWw397mGWI1OA1B53
C5WMzgEgvKdduNI5UGHU+wNOdy/WjXR5lqWarfIeH/HfZRCdn/1qOy+zWTj3IG4kzbIM1PlULiEu
979zRHxqky5xWt5AcNlfrH2LsS3ixWlBA/OrpcayS3984uRqVDTW0yF+imyQQx2MApAUSwEJ3yAW
VHpYTZMwJuDcDPAKK8CJvZQZM++0GoPSjbnK5MTrRCpMNoybovyDslWM1W3DQwiCA5gtQ4oN+xFi
ONj5tkPQCbJolG02xtskXUYLY/8b5TkMJ3cNopb7Z65E2yLsL7bUKs2Mwr6NVML971MpdsKMtAKO
VlGoYe7m9FQYGP9/uUHtTglQfRh0xq2h5dvFwFTN0YjBLUinki6/bJqHZpvJQRXxrDXzY0iVM330
lJd7FYzn50ZL/hAIeaQOlx+YXdtDKicdKFDeSYIqTUDW67z/9V3ql39SsSyui/e5LoV+oIOvjm+e
CHUzgXiUrhqEVfeLjjzXBpmOGFWVnj9pkY1NwJwK9F0p6hTfbPGT4kHSxIFaDidB61ckjpUCSIFm
cu/v8HDhUrTfSHidiZZ/itvEzrzbiyYML0O/kl67BhQpAgk2D6i9hAoO3faqRfPwjpcznW5VtgpD
1jsiwLjwijVvprUOB7RECkgCUto6bT04mmKF2ug+Va/epvLdUWw627VchpAiHdxI2irqwckuty6s
Yp8JOdB+f40yryXouoSJdodlktKS0/UarF0ANVMMfCwUKHh1kVtDudFe5QmXu8O+5RD3u53rmjlX
ornCAs0f/FfPGcxOM2u3G/2MKTFWYXYrCJQNzradIhd5epCG1yVNRzTizYxLcGtDkMiQbUn+44oO
3eveCv2gij1CNzLWJB4pUtRxyc/ja8Ywz3ZFIY3qULJ7XNKwnIBufmeP5RmPiLPrmmrWx8TxKYXz
E+PCxHy6fqNFe1lKVAzF0bs+22f7oCXVD0ASYYdRWgqDX96VkuBxrscc4px3GTHbJOO11/0dlBZ/
nBF2f+ep1gsFg8B+GqN4KZ5jAbRuIUrULGjH8BpR1nWisfwoRyCXegiPFc1VetZtOSE8ybCgk+Dx
rBcjnUTy1hZJ0phOP8DPEFeOrMj8J4gwiIL7+E5DTKD5R9SFr+b7YxLlNW7KeCwvmw/JBRvY8F/L
nEPkzVtuJZMY3T++gqnZW0TmdsKhf8aUT9i6/aucq1s33uiO56Z7r29Eq+ixSQOJ7w7Fi9sz0kKn
Pz0iBX0qyzhwqXo4cWD0WDn7TySsTJIgvcDqTnKYYOsiNBcIEdin2OBUM7tASCBlVs4nd/bhHzi7
YA+UCw3w4L5i055l/17UqMmNx+5CjzGuFLf/HO1q5ckKdKkwBzYasUo/4c3ziXwUbQ243fWkceJw
9sn3co882npLFVdU48LpVG3NZXGCiKtMMUYAPT+GyBc5DhlQ3Zg2V2Z7zyS8TpkVgektXaWNUAnc
o5dk7L/BMEsmTcv8lB7M8GdbYRKaZPUHSo7Wo1clmOzc8uh221iPokhszcJ1b2cHBSeFoZ2akJzj
jzfotCP9+S9E628az16UhxIDbcGXc3mcB1FL/5TJoGy9warg3weAUlQP5hgdPX8+sNejqaY4kdOw
nlFi/HW8WRAjyZL/8Q3ut5qLRWn3+Km/lXJSWeukvZlYccLdIlTZECZlnQmEPZ8HT8tV/TJsLdo3
r4I7VZ0N3HcQzkwIz79ws773UXpxgwNfq9c4Ka6/+ueTHwbKGHUfpDO521hhfgJi4ZnPZhRePJve
77KmlldMeg8gDUodLdB1TYSvDvCTHaFOYLYCmYFoGCAuIGPNA7ZIk3t9Ll8WvqTB+2L8tawWbnE2
bLVoS64U5Nkr6napG7SaJeKkUakTpZhxTdztpxBlGQFIzGjzlEpZGzCjg9SfoHMBiAU1yaGsxlOx
70qeeEQ5vpUTx2UtUssoRQUuTwYTkMXywoJy5HuaBzW7+kYG/APgc3bOTok62bQHPJ2ITitf0nzE
gH3ifToDR86n0uVGGpres+NFDiSmR6qh/i/x8dtH8V4QGzqC1QCq3GZwypRDtsqpXtg5PBLlk2kk
afxCS0YkRXJfNHug3gGH/w5KSh/gjf6p5XMQHYbmm3j2Uk6litZVJTtHyqOOrJFX6ELRFMlVQ2MU
O4iBPQ0rvf2/PdvCaDtAl+eg+VKeXVnHkX0LVmqa18HQlNnd8n9M3zcxL4ctnOTqL0MXnWP0KTq+
57uBPY2gEYVVNitXXEBakbpc5g3F2laNFJmqke3kmBv2BAqkqMNtcls3eoBf8JlEaSbnaEkLkU9R
yJX+zsvnxBazf5tORZ3yrVc5OkTM/gqXN2sWN2uyHL73BYPhLlfG8qaJwk/TmQD+sl/yjo8hFyYU
XA3KpLwrTIDhmyDB6hK4HNSD1hrLK1Vs4XKJhlL6dLwY2UM5N2C8eDkdycrNwliWfLyBk1A3rUip
kp+gGHIybYWCA+KnrFOtAdhHjyEZ/BPs5zSGHLTFT9E1CMsB5fDwfAkJMMsq6mGLg+OEfj52k5uk
GRmhf1wxqiS2Z9AeKkahxiTQCS6sF9LD2h1hoiIdh3zj0ehouoTK7ezqMlFTZyIYvWryULQXYzqj
C5wJm3Ho79QOCSbeP4eRzxHsSzc3pHS8AHEWF3h9CuxWuVBhNrc4q0lXM+QskXzYHyzZcimmmMMC
uyE3qKWxoBZR+KDsPnHA7bYyCQcMp/nd+GcHZBC1pQt8jKilqQcel/CUmK1ZPJE0TOQ3q0lU83jA
RmzpIzTegWE4vw/LAVtg7ISDA+wIHyJEtGPxLy7yzqIRdAVxsvu3UjU8U5BLKd8LRlngd50D9Ly8
0dahHSLsgsxM2fSmidLKtoLOxAlaNvQPK2tZtL4CaAnXiGu7lEH88srl7aTmk1+OkWo6iN1Ddgfp
kPpGuWypZwPc5GMo1bUuJmsyIn32MZH/9HO8KpMg48FZvKXPSeU/QiCFmDsTQvAZLpce+y0=
`protect end_protected
