-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LYYaFFYL3rCQ5363CGKznbc+SbdueByZM+uf0d7pRMz9XNQjZcC/hWDpQkSZsj4uGA1Xpm78trZQ
SxbCdTRselk8x2Yhr9ZO5lTQ16EOdtckI5KggRk1zkdtC60aWn7/JWRJsHn6NA10bGTS2yTmwB0z
VNk60t3ObxbkZ2sU0EUwMxIa/OHnvANd/phTBls4MmX36WwNqCUzzY1jcAYJFs/9oes6UijMcLkd
zVcrVicBTcQXQGstnimqlzU3seL3USDwDLL64x34M8MVo92UG2x0E/caJiM5Rn4rPVORyxBWRz20
IdAbL54BwRBN4qp6oCdxTxTE7BGuD3iPe4UHyw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
xvujyG3s3/HaHZtIVErScKmeeJHG8wCqPrC+/gyRjGE7/jalw5VoKmzAXdKHzAFZIqHFaTOxcU7e
T1BmNMUjk18hvajijqT4Ws63EPihYUAM6kGfB3CyoXT2TQKHKqpte+iu1bsuhDNXDHD7uEOXxqUg
U17lSFAYboDVNaGjHkiQ7g5fB6vDujD0+N5p0BdRKKz/IBh39w20WLOCluCRT6ko5LL+TtDtM440
tkMHnmIpA9y+FVXgoZlNLYI1M2RwRRJRozYixaErdr3JDv0PhnRriayzmxSY0XFmDEmzIEhwUq+g
9YBJP7953hJudYp6RmMa/ZB6AZsXoXBTnJlvCuprrHvSHyQTkhDQzehRsI6dJEe2qSc8+8WHdNQv
AeffwZSmie8Vq74in7D5ykEE7XfIQ9Thrbz7UcTVX6Do+fiiGzvXaYaQmoF4jT1onX7y2KwYmKB+
QkqHS0fkvP+YyA1Lxc9vXkuwdKhlre6gjQUWkHCuKmMvimQpKUIS0nTHUJd7189CAfgmhilJ9cxZ
BAQOI7ZcPY2WeVEkALN+Wm6cUXZmbjc8TrTkYH4dwD51P8+IJ/9tb8BfnFCyrXpeYRvPAN+JRDBW
zCFsaDn8V8Ruc5D/p7Fmy6H5FU4AjNOpBn/DSD41FtlrH5WaLKGXoOTMtsWHI+TOgLdszEHI20Oj
4GFLglFbatMuocSQ1YLH+ygurkOJAg3mkhqAHkxuS4zWd5b2ldKU82zgtJny/rd4t8Y6UgfH0QCk
2OxgCp3GIXhQv9KVZBtMHhq21xVQQWrYPGQUJnlZq1EE82lU8almqLOaz5Og0Yw+769fGgV7W9Gv
WQvTxKD6iQhrRus6K0+3VQGy+vMVGOitAlZi2ArfKisT1vs8BbRMY9DU0kzvM79TgrkLzgJ+eAlq
DFC9AqaywEIrekn2xCb5OfuBkG7T+TCJsMwwz2x9FcOKGnkZLV8ELava9cBGHWdcNF5uZMRuEKYh
4VFwWH8WXtkrFQuFLnJPBgJLDVgTmhiPNSDVxdT0V6O5J64EytSDkT8KRMX69O6IfTn0/PQbWp+/
aCBGlf591tY3kN5HIIPtNH7Cw1zZlzMo9hTqJYSMsmRQ9/ffPhOP6OYtpURU6KzrKfXHSFsUSPS/
xeqv3FL0ThnhMWo4T7A3JRKHxEqH0uSkzsh/W3EBrJtE6aN1HBMTAVFAs4/whfZyGQD+AYjSX0k5
aTwfLM+ytVsGPBAGCdlCb7knsUGmK9SjDTB55SxtX8+vQu/lqvhbIOWa0ov1OakFo5NNf1HM/AV0
lkaPxJQl2tvdiNIW9hGW7iPsI70p5Kye1yJ9HdCjhjpbEiCjNV7YtD9om73ZVKzQBv9zqbMzipqE
ULVy49HwjBLWAL6yUhik75o4lxeFFZPAnPCVx24dCaHCw8KuvFS6h80c4B0rcFavysGtClw9A8IA
CskXhHoKMezWVch+yAUkz0cjOdKmPFxU7FUgnh2p/wKRns4JSL4iMqVCmAoZ56iXTnEGM6Iqgin3
FesqUHPiQluWvJf5VGoDtyZ+D7Xh3K8Vi7OudWLaIRDcKdo61qkW0tro7STsuq1e1oENPYnncdzW
b/lu9dVgZE9IYFwEr9yRwQijBEfBIBuobtKuUg1YF32x1Szimq4HHkI3mcFrDf40FYIsJ3BmpVTp
XYAGeQrvOKl6qlGf/xGdocfHUQM6H4SBfnE2acQY9wczPjo5Lm/0+FWisKBZLf+JnhILz4NBmaEN
RobMHwfvaGQV9i9k/XzZkd5GunzoGwSm8CoMeXS5TBGXeeTwl1xIFka6elrzyLC/Pgx7iLhn7+HY
cMwyaSKE8JmY100UAvQc0yPMQBYnKgeThNfSko7AmXDQNt1e8N4DZRMhg2v2CIYk8sXdLLuVz1KN
Bfu2AtYC+oQAhQY4cajX00HQWB6rOB2x2LouibkMtDEPhDWoJyTDEJv/yeEemQoxH4LcjqznigWB
wIxIq/HCYog3Y9Bg10dk8Cl6iR2aobS7od2/UL8mIRAA3I0DYc0/OUpQ65/L5ow8nAH1cUALaqQF
VRFDLwB1st0peCvD4gdc19gdJn4KqK7Spobv+P4igywEz5e0aMhYvMjo6AEJ4mybnmDf2DWSkFlO
yjHjtCN+58j/4HpCtXm4QN3Sz2steNfFHQDXPjRxL4xhVATVQmYHjPmOQftjPaFBFTps4c3lxL5L
XCe/VpVXPIaqRaAx0tgszrjvNv/u1ssYBIx7SO23P7OoS8e3mFSQGXnwIjV6VmA4vPzjuHLxHTsb
SpPp2MI4En1jk60SoXaS6DSb/MLAmc3HlcxftCQ05qCbkfyaMt92j582WFu0b2NONc9yqPMelXtr
CPlbjrXrYFa9laUZuZqT1NqE1RQHH+fUv0Z53wYE37VTkTAWKMUpzektYh/jDEE8B+3Mtimuy5DS
LySWLTVt3GkvUWjj0trQ1tUEyCe+Sc7jO6KL+05pei2etlL84FDoJSN+hMwgWB1ODvKz7WRWCsrN
TaDbou2hz7uCJs3MomdsJz7DiLlc+0wInD6vTUfc0F7GVxA26lTcYOhbL7/UZBzAwRqjbzmaBWXb
bTjCDH0WaClwbNeoOosn2RjflgF3vyoNXJFvjywvenT+s4KzhI6e4HxiBmUiYQ0lfy0ZOJrvSDoc
0ny/GGxxdYYwGU68xwuLYp476MsqQqNgvivbCY2gy+74dFckSXh681zhB7spW3coxZ78lS5iMirA
CHOwE6lmjdXroAAOmt+S32BlnNJ5+OyO8KbRTfzpZMNGLUwqJfyde8qVNydckSmw8LIiklA/z58l
/TnVWq61KwiyzfPP16YhbUTW82Zdp8XVFQC7yVulJp16tMR3w7tQI5MqSmP8BrLgR9QSbwNnAMNM
G9c8UPpB1JSRzM2syxVImcgmEYkpX4mlZICoij1j0bw8GP2hAMndqodJVJjcz1WdOf8KNX/UZsJ6
xGT4YNknRAndvitCNwToyVzEQIkKFN/T+mVbyYawT3x3/XohPTEVZKlUKL7dELwfQDiLtZCjF8mk
4+WLHincM98YVmNenMYcoO4CWFvKT4QfqsjMafBvVzFouwr834ItYsDInVxAF4GBuvmcnlg3vy7K
POVXuH//M5AltRUZYfLoxv0tx3mhVXk+2azrSxgql2Jl/3aU94z3nM5XZJ6aveUkA8HO0ufH5YJT
eHHKy2pvCY4A01RjNyWfzp5RYkFmB4dVlFC7TVQybtaqB92yiwAMwfZ+/SshUC3l0SCiSBHWb2BZ
usxBcwNesUhTLUnjIMRNJJyTE6p1lxUOr29dPr9ldq4JIDRckkLduX5yshYYiICOyIlrQfTA+LCS
AuZE09KWPGu/0iIUn//WF5IrkK4EFaQEY0goGgStY6exKa7c0DJB6DjI3v/TGdahZnYN7bETB18J
j7yOm3rtBTz2FJvCrpIrIVdtH5+ytoRqHH01ABpu1duw6yDD8fi9EJtsRTYDWqIseEDHA+l5uFMx
wveDldjFZifp2mt2cVkD3+jq6qWXqrWD0lnEow2pXgKaid1SbEm2I+LK+ZwZgwfK/G1I/8AjBuX8
AYa+kY4AXQGcN1DNAZoaI1lEjNojvUuBMvfExCM3s9fU+oynVaXEn6+stmZGwnVPdMqoUI+806da
QcQCnaUv+6WmNAGiGNyxfyb66ymGX5tSyyroxZbnFh2z3P3dEHjOB6yJKOd6xRjZvncbhMcDNfwd
412BlfJEoW5/1yttf/WUTJ464ui+yEYjlWKyEaRKfULKlVSlf+xiVgX1VQSAaeXgRjL7NlIVEF/6
R4sTyCGuIb6b1WQjjCl+XLFALcsGGEMlGo6EKQYubQbd0MOxviqUSJJc3rReqT+GbaeU576q3q+W
OjqQOuJUfNEBXybP+QALBxK/ddsdmMw66Tjujr7KZ5SwmACAB9JcPpu8yLf9P/ITBvqHJ0PrDt21
MLQh2GoCI5zcC0zYNLj068QPgrZFWd0MZHg3oYxAmvmUippbDM2GuFKqc5YNWO4bDGnXW6Gq0KJz
aG7wqXTGBfD0dI24zSPsHQKFh4CeumDQavGrxx3lkBc/5n+8p6bpY0LXCL+Wg8dimvp+IajJH+wU
RrYF59KHILk8HSyFDOBgi2aVpzxMUWDu12JqEObvbtk1gZQUGtnoJKQL8T8q7MRlpA7htYmTP8ht
2v+adcUSALcaXYShBT2F+VwVihI1/SDMbv9vqYgGbykYqUXHpHKZVXffwDEo0vj9en7E2LYnI1Xr
h4x9psYCXC1T02NGo78VIDokaZIj2pHYNlccOjrzVgRxF0srHKi0ubQcArzjTU4RXQ6CRm3ZVtmX
L5T5lzBlyCitoBZAu8LtumnUyjJyZXC+pVEZYxLJR6vtPztm6G700ms0O/3FM00Xe/qYAzDr6WGA
DAmwnXrnQjtflt6E3srOjS8CGAWJD2tsl1lB4Ft3RostpxCryXL4tiaGyGaQ4DX/N253dlWC9eRy
fE7GU2nuBLMT1ZHjc+rA6IdK9Q5a/hFW7J58XuIHPLSGlzVmTYuS7Lfe264cWPVwQgyjkWFgH3Of
WzUal1Oj/a0iKnnevFMG8YP/pOkZdmpJwV+NRLvWwXJ8+0huqAqKFg25oW5b/RirPFHMKdfsVLwj
Uo5M4pYUmSEr6JKQaNLzVli9amOS296r1fDuo4X8wI4/ohL6N2DnlNsimggvQy28V/+L0eYYZKAf
CNolGH0QkRhluvJb+32W8mqS+tifxNsTvbOW3nU/N2cVggQIJcJ75y6Uy8DDQd6QHPr1ZTwRcw5J
Ka1U14KX3dI5ba3RxvCmse4hAcQKMn4GQA9JyA+UmmM/sJiwEKozWD3UODPliPd2cCjd4CtjzQml
6qbAEH9Ekb7QglcdTyYBhWn0MEmjgAl5eu5EfhdeyVGi245mfiJfxAfMHTP1OyWueQJcclyonqtQ
bfbuQks8wfZ96FNDDEEeITRIZ6IatTaAXHfbP07PJBwQbGRiSLoC/vBecYwAnVLz2RESObhTbMEL
OPfTNXftBX08HkCIok0vwx0PwzeT+LJjeZmlqAd5p6Z5FLcqLbumwimQx2GD6uaMF611WOuJpTJh
g1VvWZlsk6XR3YjqQVMEHtY4QP3gpzrVg2eNtkZ/Kt4haImA/IPfoPr1dMBZog4deHimEqpmIRZ3
zJ1cC/kdSgMHcxpDTuCUf0tb88/0LqM+gMWNNMwlmlcXPIuM0GwT9M/I14DmNTLexAmzBAAJUt4z
geWOrMXA4LZ87cM3bR8npsBLAZqXDjtHEE7h/WSwyokDBQCD+/4L9/oeEkleST6n++1qBV+Il8DR
vvs5M3w4HKQUSwxAUn41JB0AzVBMPBwUN+1SSndJHajpDg26DgO5EJuBr204kAWvkTakDzCR0t2G
m+fqVKeOrXaafAEQNo3Y4aym8URP/Xe0TFWoUI3Dtg8LQRRqTZ/NxG2f7o6d+YCtbNsCb+zVVROV
dtq+H0NE1i133Iw1nvBeexmnmGSp6O2jtKFm/4JEEWuqLgw7S9V8LY4KAIdcx7+mGTptp3JuNDHD
1OYfeLklXvXTq6vcgtBZgM94FkorARw3Cd7dY5yAP2Z+3VD52oOCYoF5AYDa7Jq6Oi1jjHcMV3XP
+eOT28YYzTLfWYgJPHyCNOTuYxnTfn2qm067jPiimu2+WdZi7j4M2urdO0/6So3kYR/Wgb7du6bO
BZBEhhrliORP3LP76ArEDmgUjOSdN8Hjnce+SGOY70lXxjP3T9BR41qr1h4Mtl6meaXPUp3+T1lg
aGv7BJXAQzxsvFY1c+JtWmONtCRq1g4uyqFND53qYeXdcnvXCibluaLFoy1Ho6dOy9enEDuQusI2
/sveRYdgt6G6JCg/GStkP8V5xifqzF2UcAhsFnbRR+CNnvH6vwqXpNS5tcyVst0nLpdisQ2BeskJ
fO9TmwSeM3kf4Sj4GvxNoOkzoUvMO4MIDmSMmtiS69wZn/FCTQgLzRWwum9WRaqrIXxcjvoHNxp7
BF98jf6wYAumEIqFCxawH1VVYf0x7NLoml7u5NeJ6gpsv8/gvsgUYEmDwEZGBhyCr+sk/N5oBHAj
ZjTXk/SBUSnl+rAwRP5E7ZQkxcEMb5JcgPWWhW/9R9dw7EYhfJAXRqqJ0tWOY5X6acsnVJ/q7FNw
pXNogQaXexYWGCBd6HfUp5pcMTVmNt7I/S0PRai2xnJmhGLKh4uSIJlF9SklghirYElS2X8oIgue
MO5sEHD6wAU3woYd0nrlKz0RNIsT8Kf4VU73GvYr+VhqC4u1UOTV4dsc0OJXV1BQluJxrZkBO/x9
HOzN43vs8UOQnyBK2BHDkIVHKTWhqC+rbDGq9y9JYJ9rOagAp5TkDf0qPWB9yqAN1Vp8Fs2X9aM3
fM1/5yaHG9JV3fBMykAgTtEjrC32ji22ZXMe8w2//VB0VnAMFaNCz0eZndsjEyIimtDW/4rwjLl9
r/vkGkwqw+x6nMmJrEm1ejS22Ikmsr98dEKU3xpiAqqNP2aaEmDcy+9VChOYOkLORk9EKIFAhPnV
FdNEoi7BikHy3Vw4Op77wncTzo2PPw2ioFBR0Ixxzz8JzEkbQ+BYqpAxtxWnM/s9NM1QdsninsSN
b6BJKfVaFbe/etKkqsUMHhPidNkTFBt6xmsSjcfFrs1eHEZsEViWwIyguJhRhLJShdD4hJ31Frsq
km9keFLiQidLIcJpi4DTLLaIBibH5l8t8oE4Zttq6SiVKc7yquUnosjqp/AUp/iJKbD75O1E1KtX
Kx3CYBRUQQgm0X01+BI3Fz7heP7zQ9tHcRggP1GQ96byjrS/bIhPBrOS36JFAyUs4WORAZNlKxmn
ajQZrKKR2ffJvLpFj7JiqfJcJIKPk+P56uYwb7wRb03JQ/KwjkglxKtNRYVCY9pFVrRhZjNrDNYE
63e90hOjQFUF15uSWfsdft88HUFirKGLwexO89aeZchAmmGD8N04CsIc3x4nsTY551dzrIwyuOX4
X9EfMiEt1A/AGNxt4E1e8LLL0mtns0Ck+j9vf6DZEDLZLduU50S9t5LuMMn28a0s/GdO8VKsGN5J
kyIdjDpJa8w3xbU/802LxgaJR8oJKUj9PwbHbYrh5bzH6ef86noyG4OYP8JywDbdEPgbmeb7hNXb
HOUvVZk39D6hon4Yw6FvMT82EV/IE9ac5XdvQl0pzAfg5CWTvNBuzKgMTXaQWGaLh1GUPrWQmvG5
qPaPC7R5n6wg7oYwx8buAL2TJzvAZUXu+Kse39ARoZplOiQNPdq+/1xC5YvhMLDao+J6oSoDFHRS
srtL7VWn346+4BnHCJggOjwbAr0pRMowNaaBOywEdmoxGjZE5Jsz/7uLZyXX8kDakLwvMKuKmCpj
Lp7bbOexHM9kkcbM3agBe8AO7vShlDUPh27mLgbmLV5TK8AbFfshx38lIa3FWF0omA1O6CAzP9Y6
mbrr3iNqvNuH90lNg7tNYR+XQB44kItyGuZfgT2ytiVUQzicDUtNziGA0Kg5SVoRYnhjy6y4Z5Xn
sazMsOCYmUWikIOEVa3EBtfImKB1sYeaLaX7A3eBvgfbjAG5C1xYLJ+HCK0jmZWoxcUXiIe8BX/G
PmLPjUBVfmC/4f+sSbv/4CzkaFHThURYoY9/0zBeF9drBcM85LweeR4hJmbg5gWt9woF+xdmGnZw
2wbkHc9C4Lg5mJ5uGWd8TcbhR+TnPIvs0F7J40kT0TlYJ5HLTHNf15PsSGEqDcpO01jdyGlXemqZ
un0hwxGj0UWEmt8v4TgakLgjiN47LXb3z5eNVj82G4Dg7IvrE3FUsgaoQvDj+mCjPSsXuk/q7lq2
8iXse8L2irdKJN7dv7peOus1E9Vo17JuBeR6DEJyHfGlJKSAzSlmF+m05gUKUp+RN0E+/WLuMoiV
khwXu7Yfm3i78vTHcRgpwdkvlWGAzWh41kpq2/EHpGoukx7RcYTX2P0ZoreyA5HVcHZjoZAX8RBd
civEcp1RG0G562IJd0SGXxzf3jnu46CL+76o/Zuft8wIy/l/cqQ5RQ7uhcA8eykSn4rzuB//6D+z
4N0ngWUitbkaZDtkQQNtKlv88AlE/p/w6OPs/2r1Wm9g/oabAOb8lx5Kc3EZWboomFTrllqRV555
sTUFU7/BHztzidlpQoRsp2GJCsqWjFFbguxWMLKwmU3+G1VM2ihXEuA6QkQUbzmjY6P8tCR6zxRf
76zYBWJ8kKhtzRm73xbXXs00fVwnr6n1ASFV777VDPdho3/Gg7s9JcDXG8LPS+y/xF/SB09IjhLw
RGIcbQvrdE9wpvPS+qQnT7nvTo+qWkIhsG12HtOPncF3HQDHKrbXm7CvAqSblBT6rtGGRM2tc/7N
gCOZ8qhHUHOjnXGxQ1m3aqgkA0diHDOZa6EH76j+ljDU3RGBiRWL/GjexF5wfMwY7UvU1C+nQzPW
BF0lhENtCtETz13DhhdlmVPzrCAL0ocNZ6Adx/ff3RdRy4x/b8x2wmWiUoMS6GCBsNYByFp0f6qI
6/oo2ZvGdQd589mjvTII1lMzhmnNZ5kcN63EhiFqRCGZ3lEzApUWkJ3j7gqC4j4LIsPwnPN6xjNP
UzyR1CXEWna3tWBCm3l9/oxoNNspsywwwXkUiJE9gDlZhdkzXm3bub2gU41/BHxZTebkCOmU0Fmj
AnyMiN2LId1gOv1ZF+jQ1ndm4qP5L9WgzTrHGF9kAmLMD93h+UlPw90vaRtHILNssOjGLM3RJAJv
0mX8n08guFdpxzDsOYwc6TRVV/EzK2WIZRMIpjQKm5WPU3qQnLr/8oyokycTaTgJ8UPeDG/V/CEU
7Kv8d/Xgn/QksPnALMYCrvXRXgPkArU+kxY1rqErLZuFUo06KgN7lm6VJM1rWHfAf8btsN++1S7C
xF/FqR8SY+vZrXx8qE5lrQbzGVLauec1VYqqO0FLF0KHZj0UsopL8LxotlaEaCp2dEROX+DUmDzQ
3chkOAQFOUwcnT+1oqw8Ehbd+buJi03cI0lI+runQZy+XwRi6hwuUqNkedUNtrCTeJ3kKJcr5+kn
8nFLaJ/rrb5xcKgpcneq6Z88H0gqkesa7Fdnf6rW6oie9oFMLYUseZ1QMTOlyOEctADo9uUXfJFh
HCET/ID0+tDOj9Qiox4U4wzNZr4clXjisf+BlcZzb1rS2YMAbjVbVmufRgwFgMR8d+mI3FY5UBOn
jkqbIYTR+cslbHcKlnDpR/NhY8dQsA5tfPqk0+l7bskaq5N9wieqO7i809xru6yihEJRdjnoX6zC
AgLrD5GWHNuenz7NzL8EVJL5mATfrj2TFNsJpEroa7EG6Y2a0jevCcXur0RIvCJJd02nzjyha48d
7xuRuewkoeBPIVq3dAjeaCVznVoAOC7aPJLZzOZyNUypN844kAPiYJT8gR/cKvgscH09oRjO9XCL
nvQiYu6nG0MO0P0QZm2SF8fOQPKm33XP1Q0BOE4ao2O41LJ9kGnePxWB5X+Ik+auyzK22ogpC71z
Dpd715zF1LHMyXvMDZaddVFeRfJZ9WfC4utPLuC8yeekeC/+lIs2xYwMVR+kOF+GVmgkjI+wEkxT
q2ZHPkezznFYNIyb2KmaSUmyJJ3ikvYaA8/8Hv25RWkickP5pXpppIi/3bIlWQj5QuYliW5IGnWP
UkUhsrUyxHLx0VnT8uvmJ3JukCeWGUIj/3F8q/q0tPvKkd2e/ozOSf4Vlq77qNyFUqVfjAdwzd0+
wxZJ/Esj3EBqKroQX4VOFVffJeOsRGfgZtRkRA4QxLfR3ENrcm6Ky0PiJeerR5AikC+B0KDn23Vn
xCoFq1fRs/N5GTGI3ug7oSqkiG95WxWcMo6T3n4ywMJvX3HWYNsscv+2pK5Hv/Uv8b6IL4T0Zjkd
ZNs2YFqwwotDXoE2nPbto3vTMXt3SF7QhpLelPWKNW8f6hKqOH6mpr2NTDpBCRtkHProIV79pXEg
0NhcpBQ0QZYvd8WouAHO2tGHDtFM8vTkhyXQkX9C4q2mKKI9w5ls3FMYHYqJKHeqvdztNrKU6vAI
UzujeY7SDj+Nc8whi9w2WaMJ7ZlvN+Zd7x7JdHiAuaE7oTDD0sq1OD3JFeT1FuJEXM1AC8k64lTJ
KQBPjFOJC6M3F4y/QIB851x3bCu/0jZnCS2AmoxhSvtopIvnAwjdAKfFVb8rFLbE06sOByMEZTBx
kfF5jAPoIySJB12tDxPC/sg8gwr2DwIUr80aoH0UyQmG3QuMewfruJiApOadpeqVbmdKp7+Fdjcj
qlHHU1Aw8zCTB+oBRsPvIna91zSkH/5JLM0DRqOCKZbrEXN/P8SKHn/iJV/jwoNLTq47mykcVAaK
boQSGXQcdV2Bte4avfU4ffbjGT/EF7qrpK/mHaMbimTHT7EzI7VlsZJmlD6OpeazI8AmhzP+tAqX
/G33bLK8orNuAMZnix7SH9gVWuBrhsIWIWFL051wWUSSyjQzf+KJcOLjfI1PmFOhDhMqSkxJd99S
nsah9rHIOy9eNGzIQOKlDspsGwnpHa+yAyegclwH67nSWrnRYh+Qke1cNfgrkP5OrilOKp/RnPMY
+rkkVhlAK+JHBhyMrLvZQUbV+BrN2+WibQr2C43paCvVTlkR8Q0zlEkxsyHhP94PndmyHKn6Flpr
J4YAg8Xwx6diNP+zsNt3aGMh4TuGuX7zJfik4n6pTqQG+1w2pZkCar1R+3YxAEJTYW0/sH+E1Oma
zQ/3pWexJS4CftkaXAn+1MNAN0h+OeUSTJoZr1eLg9+cnd6vDF7ABnFns5VCz8YWCB7/4eM4M1WF
L1leKjyecW7Y2wReAZlZporR/f/q8QnG6mKe2CfK+fPPYdHJYQOFmjyZlwAuJ3WbNosyYLKP6z1+
mIbpeCNVxGzHY7ySCmDVcrqtO3Xu4TdhNXYdcUPxSSeMD02pSZoXDLsIox/Hd6hwVXAsUT32nv3t
2UK+q7UhgYnTBe1K8jL3xJ+c4RrwmkCyzuThM7hXXBI6CwGTunF8XOmEBZKS7mB1eAz16hxds35s
aTZvOhdV6LREu6FrQwO6X64MOShTQ0STrU+TdFfHeFCMqDAuFK6nGri+XxpreJe7ABLOJqPNs6tx
fbVb69mad0euM6gFRAdCDqHgtontpD+ESAfzYa/3YQCpD8IblJavLCSnjG+k7h+Z0UJ4TCqYKpvH
UgXIwitAIa3/awNHxF0hCTG4W+rFA+tm5PEVjC/i4rUu0nbRl3a8jAgzkPF7U0j0K0c04qlHTqvv
lNUUijKuM4WOWZrSHGRnIk+xTKKxqY4Zd5lejcwYWug3dWc1gqqe652+852lilfMEF03e7M4pjIs
kmh4/doQfmMeTX+cEWD4sUrcrdwo+Lbx9x5QXEheXY92ubCF5LNpTL4aITAFIqzMJINtNkTAw7R3
u3SzmZnpRFaF4Xpf4A4vKbqF0m3FbNzxsOmYW3ledkjdEI6+f+bqG0WcG0axbpUdqfzWZ8K0zCjn
qxB94NIw/iwPFrV+YdTvA1fricv9BTET2iPoGFs7IwHhDk58Hs+GND04370PfyRRPjzN6fw2j+XF
AHXn4pRjnwp60vybJlbZLsqiovp/7aRRN3r/nWQa/2TdBHPe/2eM9dcNcV2R6/7oH/6+2yZfbwIX
jv4isXAyivPiqonR31QD81Vg8emp+E3l5GrNLkVp322MbuYegI+OfxxyENg9lMD8QBFomhNzR9O7
5eGZa/SmTNk+mn+ciYhmwyQrisjmz3/6UuhTi9Ym5A3AzSZduzsvRdX57GrdCldcmDtJsMe4LhvX
LHNYwKQj3HHRGhHnUoUJqSelvis2P0ACm8vkFmgpCI4g6jCFpsKBVxLuyVAf
`protect end_protected
