-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DYA7q9Jxs8m0V6/9GLEzU95rNByQiCZ/fGjNUjXYxLIJ+WYvDx3X3t6UdMMptw4o7SarAAsSrEpY
FCdHwnE8uZTMEev1ViH1P2Qj7frlz8YFBKLC0/QORGuA4zcjCZFVCf4qCqF7CUt09T9ZRALgaI3Q
W0nOl/CMz0o28S5+kj7BGyMyHZI/kpszhR519Acopu9M4PK7qMnAiytaemTv5FkrjBYsRq8LFlJ0
dLhFSalZ7IltnjRF3ET1gFqUtLlKzcRG1YKWFpVpE8DnodseIAM852zf+4/RDqL6dxpvnVBvrWOB
ielisLteYjd6qlbQ4hbyqhCdLUO10aZEvD6JcA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
gqV2GyRNcjMWmROf851jHbGek6GQYLWTkZ4blOtQfLaTltyLVf2v7snJDZccE382N+OUBP+vd2mU
CNvJfBKJyI4cvu+ZBllsFPsZxR6EpmWxD15uGmVwEg+iyJ8qatOboJz5BibxBgsdOLQSVX+J6Udo
eYf4e7FNQ43HzWR1OdOCzwYGMNgSWKZArWG2cv3XTR7kt+EZjVVx2BQZ5GCIRcDd+Rm+I5uDjAFi
Dyp8FfpZ8lDKESJu/sYlmPw9xZdp1cRCxMaboxVl7hLWfnpXkj7Ct36/9Unz7KvfgM3Rweo9EiVI
xnDI8sGGMIkXum2B4lW8p4CyVo4SQZJ1VS4gItuYAV3USycl3pTZBQ78uTDgDJLsDUDGJ5Os6r15
lInSYVtGYyTQdpbulNtKCtJ0Bc6/Df+GqUS0O8PZGu3aEqgN8gmr00kzQH+2Z6Z6sdM0IvOB7jWG
pga4S6XI4rjuMn+wF2CWx2QRJCm3yd21VH2WzGzmsKfxnYisSD9MWo3XOncLt8g0y27DZcPqzBRa
Vkn8Y74BBR1eDxpLQZ78oXE9TfvX4uVEZDnxrUukiB5SD5+AHPKQ6ziKoYhVJIeW3pBd2y/sCM/O
Lxp41IOeyeM9hYTboyFloHUOwpphGtMjuUmLtcwFmlX/FKvD/3Y4+9ZvNaFLemtI2zGC4WXMioXA
0mzH6ORcLc5R24DchrI7yQfK8WLHj1NNxCwdewx/N6qK3349pFjkVCEvz/HIMIJfyr7lD5frrST5
E85MsRu/N5qpg7+imXo0vY3uFKDW6uN1cvJMMkYHsJRw4aA6NgoHJdhmaKNwRZ0MF7iurhuLnDYr
8Q55q89sgy+6rDA868XXSOGJVtU6FRvO2OegstLxg9Er99ktsX51K2saVQefsrrIKRnAKAaaprb5
tPnb5j+81vGCH2RTGfXloGW+6L4lfeGcDkcZzn9yW9SEH8J6lQgK9jaSNsny7hh0P8+LDCIHtY6P
ROz7jE3EJO4GHijWEfvPgEFfQNiRTHEHoEE+3jdYyJ47Ih7ZmJilLgaLmxyeZoGh1Q7BUrpt9via
NZ+uvQSPn7gSYhVkSqXM1/oZjT5C76/xEMBSlzdiBkyn1nvAbds4foxnh5UlxDIveyAYMmakXrSt
z7KiFQqSOd7DzbC/oOYDPmTTYpiaGu95i7an3AL2Gn/bk/RiLb83WcLJGCZNinDYB24q5AJTkywT
VXL3t/nNEGseqijmCzwW6tpih3OriabgXeZx5QexQnAtjVVfg1yesWfH58GUaHRMY6rap3/OD0Fm
nnjFFoI6TeiWTlQ3uA8vVV0EaijsubXAUIy5cUvhhZIDIPO1R2mezWzUHYdeIbkWkj4TJmrhogkN
D3LLJzyoeeEw9honFVJ1HOe5MaMrK/N+78k/4NB+NOLttV5zQACRORZDwYUXBzmlGsJK0L8H8O6f
UXJ1tjIVBG6q7YfpStVWFBjTLFbUmB2TIOUpFA9tYpbvR3d7+RMmkUxEZiR8wn95SuZNwzBmO/Es
sYVhcQoTa2S2PD4JuBdQ1w6jFNI+oU8FpzhAF6xPKBa5OL1CUP/phSyyljqOJON3741jHfFYYvho
0uCc49wpOAnVwWaGYm8ad+KmlHwMElf1lxhmU6zuqldF7mmlvsk1cfuzZO9wyc22jpcyl2efsDB0
dB38mHViKNlSzohan7iIOq6iQc0Jo24xe+JJnCIqROknIqHGjjCBtpP9UYstMMe6nb/tGFP9kIfI
hAKt6X/gg6Zb+BV5uHEbLiroKtRhrskh2LiAY+PcPMTO3MMpdwS6OJWA1me7mVbxHtJGyULX5xs+
H3BXu6ip0/mOh09mrh/UJwWlEh5U65WHYmYB7oXN/p2OHrN3EPJAoLDP3nz/MhlbEncCDJ+YEnSW
kltGS5ANDhmoB8KpMEWoyFrIcG++imR+k3lX7QMXABIAeCmsrLCV0WNmiFgaO9ED7I0QBYwcxqDF
JMuLC2IVqfC2poaJ5i+34wQC2J2X1tWF6dG/uDUP3vGsnIpC3ZN3BBKZz3Vxa3JieEhCjjqshf9z
nxqn2FbKK0ctg3KHevSQi8bi/YJC0ZkY10keUtkYq2acvfwk/4iKp+JCZgXxkriZY4sMjtbWyHPU
g1DAB0Yzr15+Q3idddZlOAIwUouBW7n4dUsQnPJBnuq+6Io6f6g3zIzzyV34tKOhIHQbjkvpiEav
m9izLGvMwI8fpqq8KsOQn1yNCFBs/gd770m/qrxmlnj7KMXEzC8ixsvIUupbWsffzXJiCtcUWJhh
yym3Ne+Ezm8VNSvm5LeYpIKOohDLefMDwE2oruWmO9Q+hCxLNw+u9ee8h5xQKSo+p5sQqgkb2d2r
j0MFmAX81ZcXo8ZJZKLzCMgEjL1/wo5oPw1MNkB8GcK8KYx/6luSCRLbhc+GrRAB9hlb9JvK1ROs
ZlKKcVghQf46g9kycbXyUfxeYbKVhd9tprLAEw9CvxJ1F3Ik3X0vKgaS1feQIEW0yCGq5OtLSQRj
N5GIYnVQGoH6xuwND/2qCp7rZhyW0ZuAPm7bpJ2KYSg+DdHV+RWtpWszWXI6zFBlGSs+sKsvFX63
3fP275NRWaK0AvG/5rtGgUFcsuGmMUBzVQArCoMhZLY9/rTOo7iVB1uVatQGq2dPPGWP6pFkAxqx
WJsZBiPHRMPtnqSrFaTUJKNb4ZIwcx+2is6tQaYWfYlIWeNmODSzAf5HxHnM3kSvU6H68F+Qtf9z
k1LoTSCGjq0R+hfmkuIxSU76V+MB7wpmAmVf06c/RpcBGkmSubWKNyr3J8VFW0c/xKulTXzzBFK0
cl/eBEly6Gn5scTQaHEbJWQe3mXlO4vFGdd5hRANE4F8121zUDZ5i5L84NsYU8iCdY57UDyGRhVC
SJbyIhJe4+GEg8xDN+qyRH9KiVf5hZzm8F7WJN7wdhanYosWx0YSuUUNX2Jh4TCXN+8Mx7h9gXWG
jE8mW+VSwxqjaM3bC9BpqPqJoe0yLrJA6zFxmUls1YYJNnhyd1B1nmlyXr1ZomlnFqZ2evbtSenG
GjOKoomUYvoN6PPWAN9E/Gtx0ZKGvFFSDlchkHvt6x2GBXk6BArmfnAZbmGWZOlkGtcLdxQOJc6K
O8RjLMZW1tmtGhZ+lqSDiD0Uc9+JeY88HXd9DcIwF0d9YJ/lBNu8JLiTDVE27oWyEjccCU+Y+SbL
U/v63qlHneftl0ikf3cEBJlRU5oGMfRcEI9xijqWWeKJ29vZSLmZA5sfOCSfEMaUB9hMJnNLNsaq
u1bNgGiNGI67pE7mc903U7cZbxhPQSXC38UO5/1fFiRre+XD0I3KN4WDoWb9UBKxSTiHanRUJ1cg
gjzV3UAHZaauSv18Cqlz9WWtaqqKHzwGkXTyAnUmhHOtddp0nWupl0gXZljH7Gw9ASOsHzxEQFAY
0rUnh1W1I6RAelfUv+2GrKzHlYGCGNkF4FhSUishdJm1OeT8caIYnHXThNnmBqVtAp95dVAOEvMx
/LzNgOkePoLYbdoghWavcG3VyZ1Jiv4dvbgfhk6lHt5bfXuK2JqyYtfIu6CwW5lJoOIDmXG7hBg1
ZtZzKozVwbbc1rIrtAdvMPbHBXbKrHGVSL/jdMMm1WZ5J5evVi/oIcB64RZ5WqhSykjQDT4V3ctm
LceKB1pFY+3Y7B5nG7N3U2adeyFPZOeesQb5jBe/T3enicyaJCxH5/rhVuOmIqjhB2eyBnC4SmTF
jmrUIl7kzI4AAbzZU47Flhmy/c2tDglKneNrq4N/0NDy1qjTGt6/b6Hb8sXmLtYBSojgGoN5Pvx6
y4LP4dftEYUtk/BJZ/o/Fk70WUK4fFyPz070NxIQbsVHOQ2krZUzdPcmk2rypSCTx6Z7IfcbfK5B
hQW9PhB9it2/r8mJM2OM3AmIipShS3p6nhIqVWFN77Psst74H4CNhsEOW0nrzBz7cRATdJkIZb/4
ydX1oX3+qxAMq0m2Fk2JwdgWaaniqIOkYG7Rp4gciJOuD5XcKlHHtMfEeARXggtZuHoP1UOkGmn0
kSMkwgyTreGvpMmi+cxsRubfzbPLoWEPNiXaW4ohX09k4PqRRfLaSURc9KKg1jquIvwFQK1akFeV
9ae+wLRE8WtNfZvl7vj3jl6OZ9dO/GMgNYyI6OOtTPjxgzQxzh9a/wCCGQ9QzQeR86QDB8XhdTO3
+bFNuOxvo/Vn1huWn7H3WKWipmmKFEEBjhWUZCFdA5NTfNSsI2TUXrHQHAoImT/DIFrfCGNm+8Jo
8oaWnpqz5W6t//jYz6PHK8wDcjC7NRIUdTkzNi47iOSDsInBFt/u9DnG3QI0Ju/ZrWUSg9tFKv2f
3uaxa8MoCa4JYrOePNBceEBSwtonO7JMi5KQWm63nemVYiaVlmNYPMKjkVO7Wg2dwmK2Wx+Gkakn
gfGFLfOgso0ZDXfFjYoiRHxS/Qq1B1lWY1A6AtmKcfTaoIFy5d2gDHlR6TOubtFaDonDvH6Tpmzh
j0DYijrdAGlTI8HwONaGGiPHVb/Li1OfGNli6HeHS7XPNN2oGRWY1oMHbecoFxtQphIbpmKQhAkh
msZD6pLA96G+jtwkycYGom0KwlplouWA9OCeifHDof4BWSp0iIGcU7f2IfE4EoFw/q8f/SlBPAJw
iy4M5eaiRT1gI6HA3dxA0VKD/yiNScVdTNzuGd4u2YeB9ZpL453KxcZKJGh6vT6IqbYgVeCQr//B
NkAY7l2Zyj7VIWuBzJyQOhUjSp9FJoNmgoVAD3/VsMZfhFSnUNCxw19B7bdVMSj4H5U6drhseo5e
SjIXzY6AAKkJf3D2ywUeIold556xg1LLpUrUaiIeYPtkuaye9RRHX4BCXvbIHIQ9/1ayoqASFzSo
XjW9sTkG/e0lDpZhonaBrHdzHNfXK5Wg3YR+jzoHLgpKd9A2aZcv7nffOUccE3Of7pMKgzy8+70k
/6I80IzL9KVEva8OsSfoF8y6kPYBw5kt3MkoxAotu9+xbSaBheYIDLXjaVz1ZdM3wfeCN0IfoAnB
j7ZPArMTtNbjJOAVx5tYf1wQesD9jwvmgeVB976s12fhlypNj3WiSs2Jb7ncYtMdbamu7POG6DNk
tg1AA9bMI7kb9MB4tfzkIQDs+t4FOe9otSnH/c49UoWmulrrO8a9FWAy74rhIt2xkhZoUM+tBhbc
EQRjJhFgRamYCFG1Do8/90ExOv5pH/uc7JVETIQYK44G1d1Gno9DAwlF3kQXsgHCyKDtAzh5UkAj
vc04lvgkJRMrPZRqHyOrVonPv0nf5XwcjFIsqyNhJ3bi8/e+aPsV077WizK0IV6IidmSKNtyBeBO
Nr+diITqoV7YwxcfxOCy4E8nQy59UQPIwCIwkv9iae/cfeyqWw/B7rurTZ7/4Vy4QEn/gJKMooHh
Y41mlXbxy/8WxwUR1nWTFGPQUWw6nr2fJosVEXqB8Ga4vh5OhYaXsKsGHVtzgIkO/yKIJXGCx8s2
WlYyTpgyc98wO/0XMTvKUY6cbs18gSdEWaEDdVfjKUTkopdeHBzgj6rInpvjCCeXgIA2PjWULEoJ
1vtcJhRKyhcjAYzIJIrp8DeHgzG0+uqHdhztu4wP6VrIuukQ6FNbhyRpIpX2lg3vz4E3TFQlFiGw
D568iqnfcyW2vGJVcUPxmnbyhCE65drAOCeduTst1ajkzLswHWkgFRUrFHLrapDQxwXMQXYuXAho
piK/Ik00jXVl3h1ejvjOstL1YOkRSzZkuqljNAdx2ESVq3V3CXSVEVwU/yBMjKIGepdJjA4RJRNN
gi/j8CjsJU33q/WmaPs79TDReQTCHrTWlKeMG6pIaa64uJqn37TNcSO9zZouZSvsZ4iHURABgK+Q
0SaUs2lRmptQXxLcDEsfJ7erkRaRIzqyBBKBtwHPyFVS9ZOIuQrlpGfyWV2miU69ybFowA3Ui102
VV7JS5Y5tkzfVeCwousva1ALITwcnbMbvy02JLcldeaqrrhsA99r6Sqv1oxj4nmXYM+0LO3orpTs
kZ7TwPuXiIf0Wz7/IsTSLKafj/Z7/ujBMtZVWOrKnqIG/A1a5aJnn8djbsWUtyr4YZ/L1WhP8AEn
XPQja8iskUuhHU3kDvuciIUy8KYmxqqLY/eP5s1tztpqBd4ToWZ9bqjUhP8e51uKVE/UJPtOR248
rLgcS5u3jbzfBbaWu4Ffnb2lYoPzb8qe71EzPlEXyBbOqn38XRwm69oRHYalNHcuD4moA75CJzk9
4EMbaw4wvtwHWci6sBxWfxvUjDCK6dI1EwmhrK2JK59Iwd+mnjyRO/36yXICLY1r9BKPmz5MdcE4
oFEeTet1XpmnS8AcPl50Ob6lFjpGgV+Q6X3yCjZmdkX9lhy3EzDSeDYT+JY4UnWabgsuWm7Sme7e
BEJCgiNkyfMoAxKxvWJbG2JSErXfILpBqbvhftZBR+l2fXdJooBZ57Du5H8PcdzDINk9/xffgpB2
0Bo0NHHrtT08LjSD+47UWmhweDEIOzmIdmOqqwYcYQ75yOjXU1b4HZJv79Bbp3/2UCFal9QCb/Uv
P3HpDWcA1TDE5AZgH5ICH5dOBkSyqchaOxvtcv86fDi9ooTIo51G8Jx0gSwOxKtuIIoWSts3NFBD
3u6gqz/ZvNKoW0AoSI0iqFFS8XakxKNsf0NbVyC7I5ommWC8NjbF4u6tv/BbTdc43t3ERxo03iyk
+DRx6AimaDmkA38Q6CCeq441rQXtMwHEO+PlK3W5GySTI6NK/nhn/BiHbIc+s1fWkhLp10j9SGkm
AI9GZNi+EH1c2CNS9WK4v4Xn3TvS1ry2f3iThlDzN/3JjVa8WUx2sqlsdjuBR473cSIsNI2EuraJ
i7XXg9qRO/R6wvyVOKGHy8F/paXKaej4B3HcVY2hwwwsKclshmigEukq9n5wLVt1UaHFE7XUqZ/8
fgWMqx+sAAvf9rS/NKhdDZEiagt36w+UnCy3EdhViljLAZmotNJUbe68D9HG07tb3be46xQutPRx
Wj2z9MEs4ebSW/7VKzN5QYseXNmlr8PeXLl5dUBQCV6vUzo8qHCJP9NM7r9RvqnXSVzytSxkLk5O
6kBDFZe7mNzyd+Yc5bjuJvJx+jmLMjTIJCfkgdDH0MHmB5OYjQ3auZvNNF7B+2nkPi3cNAIHh0WT
pCewqyxsx4ulljPsKlu86Fku4oETwfxVpPMuiIKnnv5pBcgZ5Oor5qRrlKtmBDteafe5PxxFigRl
wzJ2hmmbrjXaPbCeeONDw00jjGddQ7s3SfiJC9tJwIceDL0stw5oWXYb/PxVHoEI2MNI1V2RN9e6
uXyjWX1qzjIX1+Gbv9NGo7BZiHyUKgQPc4rYPa7NobjDGeFixbuxKxJg6HDXdAf2eLFGSCqpaaaW
wTmyaUxTE5CucHaZYiCA6DI3BSSPUTMaoLhoW0w7WkjT/cZ+3cFcMZeZF8rwFz+xZmgna0C1b0xn
0xbHEsIEn2zlO+WGCKfmVr92LOHB/Qw4KdAtI6GB23J1FLnttw0INrrwtYMx3BFMaTLzzMEeC7Vr
qAg17+9ADC7MKJ8unUeEcQWULlJj+sELldGGkgufRqmvVBtKdHlz/tpn/RdkbiTgFQJ9pbMX4etI
wW9JjmVGcEjjn15DRnHGSeCEsYEiwB/2T4wxUxm0SBUaT4ZIqz+/5G+4rHDFbhsU5lnO55Jve65i
HIviR1fNo81QR3TV9PIVq3D6a8ur1Ydn638Nb6srLv2TbqDBZV5MBOs3c5QMu9bo20XySZod91da
sSwR4jpjAmCv3IEAZ0JaT1tjRqtcgazAGlKMxbAYTYFPaWmQ5gjzLxq+5BdEbk288BsSXaanpDK0
d5bNvkamcut54WJfhxPWDgFBk0nEWc+ZgcDpfufPA44AYIZYFSdsPiYGccPRFdC2ytqLJ3UqIy0J
D+3ktb/zbTomR71RUn58WuFjunYS2n7/3wRkmHLopqKrBJHLAVQ1R+grhgMMoMSWcCqXHXSGyT07
0HEXDAv1LAj3SsOdOf46XF0iDVY3MPy9I82E8c726NFiPiDVq18h2OIHqNoq5byQS0vBSbku9oZC
gofjwecvCJ95aH0m9LV34z4pHSzGpYO0u88ihdnum7zZtPf1ElMMbUa5CUIuqA1QzuSVdrTspPAj
LJN8Vh9TQx/KHgnTIZ3xnToK2SKv40E0wBJ9CAF+8pCdavSzicocudsNTmDgYb9bdHH5d+gi204f
x+I+WA+oMZfAhjcJSQoCxrzr0gTReE5tgi2CeH0n7YWXQYWQX4UN3GDrD+TW/zvwU/sGwwwzcoaq
+RxxjJc+xZ/e+ZqOulDN8ISR0KRqC2VsPfqu8U/VuvPgIgaimuKv/Yq86xMjBuPYChjmEDMnH91r
dQhVWX8uh8EWNejYg1T+LM2KSTmZgAyNy2qbnotkD66O1s1sJEHDarro/w5HKbdvo1ATZWLGyvev
c3Z/0u+CKFBp3/XvTwXDJELNUMT9vKGceAIsR5Sq2Y5Dp8xTQiBsmWyx6AFcXE0nP1gSPmAvizUu
O3V20QSCbFSa9kltFtQk5HMnQqrLyAbNjrv8SMsJ2NTY0THIlSYXS3ORzK5B/+Z4mtCeVsnPAwJt
gbtgC2z+bOQzStKE8huLTLlQyCxAKv+JyFu1BaVYeyeHCtwHQ3whPa9JB2wTfo9GeX6goezS+C/q
M0E5nDhzE0oLpN0j0/aTjJTeMIYbi3dENCGRtbJlARO8A9cux4tSllnz9wnDfHJMg5z+6nF/8+lm
bc6niRoWk5Cfz0S+fWyC7jQqP4JuaPQ1Z8GInNyujqCztrK4G2PEX90tt9R2dCJ68GU+gTXBFIfV
I45ihbqVB4KNBUz51I6V9848si/OAfeRWlFSJgVUt1kx3TESKhkBWllQuDXfqMinYFsHoh5ssRtK
knxlgbhXueN/Bbc4jKdxCYBsz/n5/oWIE5akJv2rHv/8BRenIE4dwYKP0iGjEJXfSKLxy+bnObF4
CaPXaOPXVhYrD7Uc8h99KCYAr8p2F7a+hePx/+chaVL4otVne9XVkLfxdULuWJo8YPeP7NepYj/q
iwbPtLgAZQ2+C9TV159JroJrAr8a4glUqyyxh9n86Fj86vn8sdiksvn10NwMRGU7fplyRBdvTWf/
WXHihkqeVSsP0NovkmiLN+7DR+5KnB2Ua2SyAd37Bys8cNi+Zl1u1dcZJFVGhECR1VP2blTxTRTp
tfkStr6+W3XznmAiSmKRKaZqKYaUAlJvMw6XclO11KKKTka4xLFuZzoGoAA4u20u/0o6tJTeZMy8
HjOAi7VriYL7L9w3GxniAk1FkwO6uTjS6hyW6J/lqxoCObE5RTHDEliSpyCRWoPKXCmML+GXPDG0
TD3bJqH0ln4dUwfHWybttE/uglPbZO4uJPRNiPvE8xSKTHHFT8cwyxcKcwhQq17YMCVrL0QvNMFm
PCNGKg3dIZx5wb8saHiUbriG9dlorY2O02tFdXfQwUHZW53Ivujw9z/LY9GfdUnDcGhfPeaRupqk
jTpTmXB/EV4Cehtt7PLls5kdgEB8NfBL+ImDhDW6EtgdPch4n9e2YudJbFFZ5NwKHHJQpUSSlaCh
0zrhfSkO1dh3HHyyOBJAS6nSLTi5LNpStPsJIW+rsTJTnozJvcXgOcAV5GiT293FtNcY4GaQwfZT
BXawqeLDwZRQ4SSHN6iQXH2RPAuRJpjrNQn8U7SEWpfXrfccO+VDoBVb9Sdkkh7cmimrDKOa2v4s
8Uync7d6pqzfpQ02XkKlOl6jTOXXZDID9LNFgwNdMCuOSWB5APvvz5L+qbXLK8CrV5GfhBvNFOgL
Pv04DR6r8QpMBRQsjouZV/1lGaGXVnq+YCZKaE53UwhmDoTjaYD3GUMFSEz/deXGJGrCto1q0opL
Js9nSvXn1WhnnwG7nwEV+xq3051+tgwofUYgVDHAVu9Dyuwb5egi/JwwVf8bYZTfFIgRGjfy0u5U
sunNb4fTKJjfRL+ghvdB1H5RLO0kk2BPayryS784+8uHpHQ8WGjp2LStoQ+UFViQQYAqPgoVap0w
a+BSICKkG8DzTdg//2tzUeMZTuvTIiRzYe1Vo9F2rPXVtv0TFHm5M7RSZRZTbvFjmfyIfsLUXjaX
j9msANOHmturIAxvzaDNQ2oX+eHllEPaP0xev2vqGpZ4jMCMLkT+4QKFowqtuLjjt8NPuNsVVuCn
OVAf2U6lbReqnhXOi6jVp27hFHr/HBucOpzsFyhzlpswXhg77Y0Bt2gC/zHI4ptKiGBvduXuwGqQ
ZYnpLxcc00SNfqq9+IB1fZ/3ifqN7d782j7RhWf3QV/wyxfD3aTI5zwxffk5nphSfmn4kA0GF29n
dvQDIQs4/q0xTre8f+temM2e29OHGtdDOyG6WgW/pm0q6mTdLhiX8Ld1cpjkb9rPJN1I9m5j4XvJ
ClGRj8EqwgF+b0jc8iUcPOxUj1ERAPmve7dk8kmT1ZN4tuT4eqhk51IFlcJDQbERK3Ns8aPZ8lBI
EFnz9Cg4sRioSkgrekPRmGYMrzwnnXqh/0mGotUs8UrDAuHkdAelR4X9ydCKyCgSWdlckNxYUbWd
bmUkczxexYYrBXX/9ij5LrrPaflC0rMF3SZjYPO6j5XbIIyy2gvS1XW+TJTf4miVNuXGi7Mz8d4b
xEd6mmFYcjEGfu30PnSrcJx+MCsfoMIMKRS5ynOi9bv+oHBLCQp9jxT+/TH6HQmd146GISlPSI8z
5GOpSfhqrmrixYL/oN6BV3Xo9t67EVhQIIqFn8mr3HPCuCA41XMbiAeXhf93c9J3odHT59S+wVaE
XD1x4n80qYQfFvIMUuywKbcyphi4ArBvfoqM8niMRkaXnUmz7E48w0qUoi69WgO0+7EJjtq5lCW1
15UScnttvl0e/ikOXmEN6jAbUMG5AYU8gRugFXAvd0/BIGcj6GAKecibeWC8ZexSY61WiRKNAwfq
bNKUs43ZSZnYvdQqv9LA96bK9u+6VZm2Zr2ooAcqk7NGMtNOGD58lI7vjKo2xfra3hAPVR5hZ23D
R35fPeqlXHMKcZFPWamh6048vh365mg0vSUiXFkg1azbGEWSGv9hnzEOYZsXsq6o7nusdZA31U4n
px4xWesqhb8dDUJ1pZSe0dG9s5qFLvNab25exIPY+BYhWZ1cE9w8YUw4N1GjkkytFhrocCmWGmee
RHc+t/XO0XzUE5KBXqbROWDz82Vkt4bTN5G8+QBlLW0oxAsOt25DrkqjMue03LX1zGmRGSJk8hrF
IxxHTRCaJnLda7rgxHJOn/sNPT0SK5s9bjMh68lMPX5xn/rtgPPLCSPWc1p3pTXQa11vrL01AtZG
99gH+s/JR2HBS9qWJyxqg/VUqfWVMsjGaLVN/Wy/b5YonCXHdxdMs2F4Pwgf5igq/eoMk3rnejss
PP6ZNLA2NkMBjblGyo8rpS9bVrFjRSj7GjjsWM+W0ZvLf+0mnlr2wCMTOdr+oePFRg0eqrdEz/dt
V/p1iBqwYIlAKK0IWtELCjAMS/LANG2+yzYQ277BqC1gbnLPzgS+GVcthXGkBo/5wML16rLFrNuP
42SzkVkkNwvhDvORS8ZHSJW3WJ2nJjBoF4eiQwV6eG2eRDOgiF6JJzsM1ggVugcEpcggDw5aMbtL
rUH6j5a0ZFSfyRNvBCUWkoA9DXDPld+VbqaB08RuW5dE5Jfc5RTjSR3kjPUaP5OJ6aLE0y4sw0BE
F1iA339mnuKxdTOXW13YWCCrXOLZo+60jgdiX7QOg2ttPewGXx0n77WnKHMRgmkqXLYxdU0qa7yA
VK2lMedh8BGQCbbfDaDQJWLl4tvU3pG9v4uwGbbrl9zk359MqoGAoRxsotvq8Mpxm4ry/QHEkEQc
Akc7BgY6qmNrsS/N6AX9dG2ehoMy/jphxf6+bh2JGcHAcIEMbmTtl7+Trgl6Xut8ZEdc4Ay07lh+
8vgzZvGWqff4g4U06UWeydqK4onnqBAaEqafrqur5RA/L3Kk+ZUq4Xn/GD5G6KO2GgtVkFuB6NKO
rmhkSKeA1qSVsXt2LZkxgisRY66ujOPL4QkPBGCnkCjl87B3P/q0y7ikRjMDPxNBB9kG+iRs/WWT
3mzlG2uGA+5iWszxyyzjkCeEtMY+8f+rDuEGGWNOHaO5xKC1PwAnhSMEmOR+FsJMyxME1d5VdTTK
HBM0pb41ChAxcXUoP/CB7ziebuxUMgMo3MUczpFuvp1YPXL5A1ts0+yGbH4AnBgMCVyOHWcwMXqx
b4jxifGi6oCsuCdsk+B9DmRyXJDvkJTto/0UG12bLR+XtA0PcZzIfCyUjhEdsSNv1Ogje/b6Mw43
pCE8o8TCHxCTROH4v0e88b+2F31yfPJd//JC7YwsC+g4sPKVMU/hsCHpmpYxd/2iPwxxsEuaE9u8
qvjC9+e0mQK4RhSQ+ea90ENmIUjhbRUFqWFz9atHfwj7rCCmc+2BZZSTfdf5EFlt5JoLURmHljDS
19sO08KynBvOD4rH+Fq8jZydH989AxGQNFIXBHDhNACavokHo+14MdEvStydgIVLkZfXFac71WNf
g5e1J3ismAbkzXAk56ilhfm2/2SladCHwlPngAkFsL3qQBfqmnRdXKSF2G39Cl1DIDIgPdaM8v0g
8/LyO5O7wr4KYVYu3WN3MwJIW7bJ2mK+3DmrKGTB+LpxV75V+n6bx+b3IJfwmtjLZBe6XLsrbohm
ktDiv6NHcSQpEDSrNP261CgWQGf3MVPO1X5SXWghNbXUUDu98puGmFYz7lo00JQYW7ArGwxYrKOe
3E/WKqOZrpwaMuVW5tx331iorB7zCMOqDNXa3N7nPEHWum1yBoDggHIfyclef9Is3rtutXIPI4a+
gb5QWOV8vHn0PyisSnbds15y2hrXsoXq54+ELoWYz+tuTgX4ig2pVV1aBJXyWmC1i/bUEhsShMx2
fRXg0M0oow9n06DoUnlw1teJkRC4+nztyH+UPcpggbN3+pEYXW/1mamg6ZiHahwVECAUz9LpO7Xo
AgXqL0mTam6jOO0bp5d5PeVOvKAMwzFhXio53GCUb1V6XiCk9l4wAz4h5nkasramURlxoiySHvf3
eRtB99trUYCFi2NUycJssJL5uw+NUUv96YifBJytJOy4JNXKCPA9G97by0xhGwa6HuC817EXIwL6
gEKA+tc7xox11iGT2NWJs1AclenhoQFIwXOZY5qJqVKnAL1OMFocVBuJhsc4lfo59wRQM5xMfE8l
GF1wgodcO0Yzw3C++YGnyiVJXfOB0MdshPcT05eDiS2pwd51p8xkuJMyGXavYlEERqPb5ch//nX1
ApAyG8SADaGmFeYy+5D50NSvvCN4kbJUPydfSmNmiN0HGcHX+2CVwfoy6HcMKv9V9qJFHViOeHzK
U9B18ucVbHWByeUv0UDJmFUjRg2p4UwSXnmIxa6iN2ZWiV1fxbDiccYAlEBtaSoAQ32INU+HRTru
PZpwWgmp1zb1otDoEiH3Yv0ViwZOLByaTlfBw1/MExrj11X22/FgTJKaq5ZyQW+ZkbqnjFe8CbJF
PXngYJN9ixxfPVPiF866omKJ1qWmpWFxy+t1xkLyc9YgyuMctC28nAkTmnUkK8giYl/+l5UhDC9t
Jm+UqWztEQn0i6C2hdKfXzr1Mlqho2FIkkUX7ZqENyEpuvve1MqzXe0CpIEH5+ErF0O8gZFingz7
TEKy0VvB23DQsyXswz08Sp6OJ72AIKPZmmMYQsSe1uvi/wASyHQ5hYDjgtq0ZHrI2Fk7R1T8irtX
7wUx3NQpP+jJ86fjLvF2jf3sS29b3m14VDZpYwjgdrtYN4OJWofsf9yzJNadMoMuYQleunQylfa5
AT/BlRGkBr0Akai5sRD5mId33wQ9zEvHrQv1x1MBLUjWnN3ggQ7mqlO1OzTyvxc7V7K/NQNpgVXP
t3b0f40A5/1uxpexkzgdxROr9htgswEaf9wqXIR8lryTQwDpUQgBSQonX4vMp3qNIjVMQx2/W6jt
EDsBPmFkOYL8+nCJTQulC5+wVWz0kA71duliIeswVuw2Cbbp5Q30diZsH5hH2G+PupnMOrIXPRho
BnpT+SagGvLChB4U50vdshtLQxMNtBW2gmehnq2CbolH1+i7yjMbk0FT0G6j8Vc4Hk3TFUhJ5kfW
G2qxsY2+9g1tOalAx2SkLZu20zT0jwMZE44sJFiJlWRNQ8pHSA10F0es2dHJzb2OUDcIjjH1nUM6
71FUUASvjVlAssNyDZlpgSQ9ie3zY5dhqZVNoIE694NgBUJxfsqPLv/YIOFW+xD/QyWE1pRgU7kq
i/Z5NQre2oetaKmGiDwFQ4Z3rRJzNjY7Bz4GwC55SWD8z2lbzd5EdLFRlkqraVCX64CUnLiAMuN7
Q54rf1sFSaEvJcOklj23RTtuqzJcw6G5JPiF+BaVdiinrhRsb/6Cd4RsPRnZHXjJY2muYYGG0sx0
spfdVd8rmtrocs/rmKeFQzP+2295lMMezJTpXUcwyEjzzcYvgUqPbwSLGdek+oj1r4nTSdjaMiXc
1+4LqDNNv2s2JbbwjsrjMwgY8Wqs/6Fc3Dv7/8JV6qdkG/bGONn+SwAhBIzHFUHww5wFIgpiD9YY
HjDmAftfg6JT73PZ23jkxyRE+qiLQHSzHA+R/PYYNyU3oDda4pJWXSpiyx7ZZ06Tpjow4emwBlnE
kFGS9oyrwiDeFaijYroReOIG8JhXN6upffrjH3p+guthpDt2PYZs1zARv+rEh/eHiEp89Rf+qcv3
ApQcu0jLvbjDG2KgYpBQl5E44w9QjNjtvzs54pMgrfeFrVit0z7aa2HpZcXHHUPuAmObJfx6wpt8
cd7zIo1d3bGmJfkxd9txL9TNvBLXgMcBv353LE5Stqk0xkqO88TEuGlWJoLw1Y7nlpeJ02qSlHPy
5BZYnXR8gSjbqGZWwVPYgLXyTvX4UXzIoh7v3Vihjd7GCRSupwYHK6qTY1P9gtvcjQ3u/+0oZ2T3
32RKzjCffcO8YiSiLNieZq6UdmtmNp1DxK+GORCB25oQNa0tFgaDOTEN4y0mWfkyUv4aCYmrdRIR
1ZzLMfzuk50v9QwjNEo+Y8zkLF8/+wOERbVp969LGs+2LOC7KCf8JWrudg7q5/y2feDArEmvxSwa
oJL1xqBgwEj6BmQBEleqQphUnNJqVgWAuv7YqkqjDr4/9cXem2Pi8JLfPGFKXxS9uvOPCeDjVAHc
VSKfBuCD5YhDYh9qaG1BqYGARZf1+QSg19CD6cBaBcjqJdVNKcrI79r3lCqxMZWfmGHZaC0+Rnyw
3k9OkLyvCuawk+hX5WasW//mQzxVCLK5/XStsIMsWoZnOVsHNUrp1CN1SXvBsH/XkzFfQcMwKFZr
9U+f+UTiDXpFAwAVPXpP36V7lkEnqWzHMJcFOVXwEZFxUu0aEYGxRBBjaf7E1mHih2vAeUST3zlI
i/ja6+yM6pWrl9/Ymbk65/IMiXrccmFBwu3x5AeaIbKc3MW6S3CcMnBJnE/ug4sQ+6RClsBL74qO
H6ZpQtT7MKRgqcDeOwjswWSUrjkmgFoYVBzcp1SkygxE1Gorf2r9x0n5E7y+/SLi+ikgXFCS/JzL
ruLSU47mygcGVjoPVK+zZaFqAVPt4UzZ8iWJw99RzxtMw4CRo1znr3PGCJ1e70rjCZEAojZyZSBY
/9udo8EORPpB6YPnB+QaBy1qROlDXZb3byJE8aa+lYYq3QqV4rVolnOINv2uEHGdJWFE7Y60aHnn
HtTR46up02TPXD6s+Y+g5UxCCoCMqnanGxdKT7e2XUI6DsR7ZkZJGdFrFHGlAAXn0+frmksEvM2o
FPL/MGLcoK6hAJDlGGNmZ+PJ6gzHgjJR7I51Kpd4FshNimsW9zEzrsmAzgCJ2PVbH/VJecb0Dlbc
d5cE7Nn7QMx/ms4xedHpk3Uspb3GtV8CcoiR02H4sg1iMws96zsdVnbRNVKAFvvoQwGq7Dtf/1nh
VkUOotG+LPXxsNXtqIIj0AIQnukkJmOjSjjorFMqcxv6L0j21+ZqbHrAcMJDWKc0h+kDNag8hWDv
7Cp6nX/m2XPxzrr5RY0+X4VmkEMBMvPbFm2cA1QaP1TxkdnaOwZnRoWA/IfzPDhmhrIEAc9vxopi
jwtbSbOtZVWLTkWE2tvtqohcLIhVXQFDz914/4Y6bcwsIkbU5smoGIEs1YDZVa1sLa/8FVVPiGNb
OCqsJvfZnCSNSuvsSy9RxtYlZ1Vl85CliVK3DRnq7MI4yIFEZchau4dUwcwbrPzlmZBcjwepCeSo
4A2H0/6WkVvIrnmWqbvL7r6Wb5Qed3OknZ4hA0rxOmu+EalHCA5E+bC7IYAdMXfUJpmpB3lwHEAp
YkpVmhN5zh8EwuIlc/QRN5TDQKb59jAz3hvk9QcSVVOucTKzmN+ONPqqUsFPXrmuCMQbnMquJekB
fmJhoR8miYUl87hA2uWpU4t1JXeNiOVDdEtONmV8tpB5VP0Rx9paOaN6BYZYWu05I2ufHvZ1UmsW
tUUmc0jjknWiMGmVdNqeCcHwdmG2QeIsEKiKjhkHWyQxyE879NCLSjeki+qvwnY+vyLMExqovHE8
5U+1IJ3jamUa40HM4oMiSx1o7X/oE9LZDzHpCLjKgfmCDwoa1OwP3i0UB0kaeJzMVcyboHpy4plO
uYK4YvRRNUsvsF6x46ZzKIhiu3FEz4uJJ4mX380SF5Da+wehu2hnhoxpS5I4PRp29Lt0uV0Svpc3
IiT0Fdw//UUvIXcNfMYUNL72qaaQnkbUN0GC23YMtsFyTz+JUncv/fFSfn30PaAeW516qa4GxE1m
zjpmWNBiAzwvaIDcFu00R+x1PCla12LSJh7Qluje7eF3E3plQFs2RJcCDrDB1rD3XDRB99t3P2Rg
V5Pjry3R6e+erEeBU0LfmPIBkTbrnyO47OZRTZPLcZ81v3C5fWuaPCVHXkRtEAUZ8ThJIRpav+4m
QiXxMQSrqIxXGXTz67RqK0476DPGntHBPahY1PmGH0AO1zlk34092NqtJCL1/50sEaK9pzIPIJqM
kRfSrjU4mIk8ypDk68zJs/5DwVLln9zJNGoYORUO/rQtiZ+qmOCEHcAx8LBkfleCFTm2t3AdEC02
mQbJhpb+gSIpbX0/IRi+pAZyrCLRN/fBJ2TLK8see3oK7STMeDBQAcr5PNIe35n+U6au/heUottt
mgPe6daFdrqNteDZiM1EdyUkl6wMV73MRUN+Hvc8Obco9bYR8+uKagLU8IahLrYUOjZyEjzo2H+U
iiRYIH0ezR3pTrJXt8kgyFKzCeG5+7/TXYvcHBDVhrf3CzOTO8Z50kz6IMZ7vlQsW7NbfDjMPFe/
JDmhGr04Lq8MXdrSjIL0tCz/AULG7jKyoBvYFGzC/jVCCZtf4a4nqXo0unfsi5ZgniForiI9f6Y0
KWQfZA/0fRs0qVOtRhO1vtf4jys8G8jfIG/h6kCpaFSYhuEEUXQUt9AF+RAhUaY+7J5RkZfxTK6c
iM9ugdVE5qAczTUL2ORcMzjjzebzbxvs2wz1M0RlrrkJG6Z4cACfne47aeh9MoDgfqYqFNRTeRUZ
qZXK9nT/ZLYGThfDhOLUBu211ZuZDWENEwo6iiNmpZ/Pw+UJxBOoGX5Pt/zeV7Ux0t6fEvQXJgq6
023mbJNbphix1yKfPFMEIrlKeeb/BRpn/ipqQdrshy+dutYDP7cn+vpI5sHWzhiNmddOBjzPA2WQ
UJWvvagJPyBhkbMIQoliC/mSYcXcfl83XcSQA/xGQ1IFH+tH1xHLwTRGWlYgoVkaX9nlwXFkKt4A
d2MTSJW7xj0UUgU5qUCsXjFPHo5xk2CrlNiAiygMF663hNtBhSI93jB9Fbl/C0ZZfsqD64MU8u25
ubggAqi4fshwLbZ+eL8gmqzYqqPOdQZLhCZtArBdQDf8Ivv0OFWRxfeVmUBGnyi32RiZseHy+LAj
yib96qU5SUVUdaUZe5dzzPK+yxvUQoHD55Z53OwHxv7O41aQkQ2ieNi6JNHb6L125djEl16jEYYu
KqDfxRSQ6pmM1Xmie+A+x0d/VEF+RbpOeJmxm5t1+NG0DnsIWdwSEQjboorOZOIrjyhtcvRlX75H
WgiXfjVDwrz04W3n1pB1mHLypfNOQVpmQADedwLEP+sSrL7sJgtOakyznCm4aJouqg3fgCkfHKC2
8fgbXknuJN7pMqNolF1889OlJzBbTZ/vQnkgbVixYmScP9vjpS+1wQvGKqdllLEf59UZRY9S499a
7CvodAefY1zfoz+gRNqFuVWpMT4DUDIq4vnMtpEklDYneQwH17MtiiGEHkAJiYyYzsUAAng6XASj
Zo2Q66Pw/vdKXhHRyRx37nP9uW2muVdsiHiimOZWkNEzJWTtywiTGqtl+L1MSfQjL+bxstp3wLDo
EkrCRL7jbvtYfA3TpYcQc6n/1/WnNuZSxhhRSCxGqi9Dw2oHOhQpLAgIs2KfW1qruWmJ0AWXNwUc
m64QtZj+eWoF//aB6qnEBBsSXVT3DRasTS1pY8oMMXWgWgHUAevAouisbr8N3Lbd6EgbHhfSb4UG
IVYNP85CQN6/tU/akjlASVG8/CsYAl5ZEXrjH8MAFz7MAphmaAu9Gf70WBCy9PLFHGpOOH1cad2O
4bwQeFNGbAx7QUaLLzM/n4Ef2gNTNCsjppoCBLtdNq8caX9E9R42u+eaFD5+wZGpWdpYp5PGa098
rgwDmMiroFBAeY/J/+L93vmcrl/44O8fxYYLoGnn3+q1eaeVAGma3NYgmBvOGcfeAHWMHcP/CojV
I2FN2RpJra72mG+lYko/pAXLI7wH07k8HaUDusM/bzmT0gGAeuX+rI3+eoT3yHjSa6J4CxZFgTwP
/bMZK2L/iI3XqoLFwjZoUj/r+BKbmkJMnfOwbj0mPT/1QQihoo3c7Ch8krNW0jnCAM9ySYFk2Rwn
wLxq+T4GQj6DReHj/9HfQjdJTaAtd57TI2SCirFARF57QBeu/49fI2QCPfLvgHQbohjZjS8+0zqM
xTrJPtOWFv6TnpSSlH+7AW1v+APqJNeFbZ5ZQ5pioarue2W2GJJvF2SkpmOMPoxL5FAg6MFYbjTW
2ibD36utC4niB08q8PspnEKT8gpiHicXwUDW1UctsiydDPRgTGF5nuZRLvkoaunoVTMMByFPs8aU
aVKxExbvdmTUzzJQ99o+j+cqYpkcnl+LCUUvub7e6Yf37tBTaGQfCHibsoyD2jfS1Lv3aQzz1vXZ
azQsS1RbrLDxFy2Zdag2TyWpLeJl9e5St7Rxp9NkArhxGSQFOqbviYHoSTKpEPPtYaR6dKI176lt
//dmpaUJvTCyGAflqGevc4DBKAHF2m31MWzox7nyeZViWAwYSfr678kkajkunRASNblrSesZvvEv
ueHE9DOk4rydn7L4tQnHWXHSrYpBmK0C5LeLH3OcsCkKZDJbgq697YPaKf7W99T+cOuUs+Le+yM3
UZY31uziePHs5w8tGa3bXQx1gaduzlsDdulwhbNw/XyGHFxv9cgaTGCJmhvr5OAPVYdsLsilULoi
B96nVLyBjXXFnZ1BVzyo3uw8zOPbmo7IM1qXhprLgR4gDGGzo8J81nR+b6daFLhesIYfZ+5CfoCJ
03cmutqlyMnRNvjE4+duLD4ceVdSiCBcnbfi84aspNlYgMEKtd4MhWA48Iqo1AZTTxNOYZDhA3J4
1d9OKU4fX+eGnCuxnGpgxVKcuuUVSSmGhBxufdETH8r2xl2uqKrcuWPSqtouUL1aRRRwIOFjFExZ
TkHBrqidax1b4lgqskURUKJRAuQpkaPx9ikZGUNjHmRSz4x5Z1zS9/C5seITNJXjAs+KADOGOyFb
pFo/Jod04c78oaY1PDEzfN5l6EyN7miiK5S7F0e+1WXh8N8liVnYG1e6voz+Ipx5S5z6YQEafCMP
69lIBF37wWTKdXEylzYnyhUkykcIKSfuj/EN/zq7z+v2homkjZzN6RCA3ax0YlPvJ+NyLOkHhgiu
d/MNd7wZ5uINsSHnSVS4K1ffxfxzA3mfFJa8HKliwXaDsMsxgHa1DdkmweMs9Sq52bfyFNcrrrZ5
V+DmDACFBiCicDQHpTTETaeRv1bYwXbkWkBA5Qi+qmfNAmHq4qWZ9vvNi3P3qRRQ5YSAXzeKHSR4
ctLoJjmgu3baDfb9pjitHNiIDDEeVde2XwU7oCotJ0i9Cw0hNHEYGCyAeFYZzksLGxzqN6Q7GDoB
N9FLKXky9h1F0k+Al5Hcau3LvfRl7lblAnD/r50WDc4eGXrLEzWxdoDwU3I4BeahiTlpiW7P6M8+
YFX7uk72g8uTBaCjhrQ0VgUC8aE0dJ5UlZnaM/6dKAIW24/WHjLtdltsHee96uXl+JZ+64qryPxo
w+3TT2eQN5zbL2MiQabo7C/oXv+iR1btfA+hdxcorQO1RaZ2aM6dVlRL20kFo/WPYEjBiVeklcLd
HIJMDZPh8rB8e6qPMKaMrnJU7geRmYOomFQw+o0M34LhsUnDGVgvrhrxnov2TNPOJmEyXJsUQets
F4kWPE603VwzEgSiqPmEE9UzFhdC/6EkcWYNQ3VOuEudiVXhaKbsq4wobSNNedJFuk7zoOT+23oo
6kUYF9zpFhLT/IZeyO60Gv5Jzv6qWQ0J8+tsrL4lysKWuRELnMijD1e3rTWzE8fm72rkE/WdLlvj
UC3s3hQ8CjrIDLA6nxoAHZNdK6qNw/IlrurVfrMdp+a6d8VlWsxv07fiPrMDf2ylT1O1+/X0shwY
TVZwMmznD4n3juFXN6cjmYjaFHTw0rKRRAEisHran/Q/DaV3RlYM4uRLujQfwm/NtpzIngHDYHBa
E9qn+KMrSGxxCiFtEAXj7+PR7g+qXoUcNKQgyQbvCodDCX/xbh/ZuAuyUgOvUaY2ecbK80Po5/vs
b0ugKvtimCFk6vKkB1npk4b5fqDzb7saFiP1p6eH1I2DrHKjIn96FBMDqSWa/D0cyg95KKqqJhuR
RcXk7UGtmLpaQoNJOO3BzDX84/ZKEARPoGY4k5qvJn4Q7rVLIfmMDQwJYa59Vqu28gw7oth8N6Xn
0Pw2ld0K2LRYkPnBzI5163z2cBChBAL8Mf1d7afLL3rDxtUaPtt6Yslhju2ts6Nim8yeKExcod35
W0XyfMrHQ/1TdrpUvSIWMhBCC1+d6wyV+AP1JX5wWSzRRj40i1DzfZwz3gz3Oy5RKcEqyTW0RUN8
MtjIS/KPRYgV3gZgYzWl3CGa9eyaMAU8JCHSC9wrnoewdbi/BKU1xNj1ObpL/yc6bDYCWeVvzEsy
WW6vw3tw5ecpMaNFUs0sBDGNnEZXnpe2bM5JFqZj8PoELfeH76q/0jpF2bnTdYQSVvynXg/X1gHL
CDBsPlcgZM1TAYbi4CBcQpOBKksO17k9hqG1CEuQ45vbgdzA60W0cIzXwOvnVFEvsHgJeNYmBRLQ
k+WvF/NNuY1zG2EEQWwxePMHU2Fq9yrEe1vxKM7gZHp7RgcFMmdgZvOEg9g5rADqp/87xKBKbUev
VdGabaBuxLf5zOmK4DrCBljIcgtTGcl48bRR1Xr4YEy1brESo2lCS7riwE8ZBtYBOWA/ANtO4PNp
ByN75WrBkslksmGFtwpDBDjDgWz9Ls2gSHr+2KMPOH0EF+LfnZotwQ1GEXKapI8uJ8Cw3ymBBJxT
sndDNG8WxDkMk5FH7J/YyzXSIHzQqYosFE59/EKC+iOGBQd49SC4seFwOUbhsEBoQUwxDEbXJv4O
OIn9g6aHM8U9lVkr7QS42fM144yj9tivGw4IAUXBOTAICe5Jr4oyMJRsygrJGNf0C7qdz/In2gbk
OPQ1ZmgY4dUdRmEsTh19I6cgp9vGpYkFAjqNSxmktm2QlIZkgxigas1ynw2IThmdguEF10SSjGeP
59gsBScx8/YcLWHoN0Tr2zEKEJA2R1x6DGDkpeGLBGKX53LE3T51n/E3Vt+wRk6OCntW59d2/CA4
KOwbTYG2w5kIa2KPl5jXzwxq+EjXUqKchqymuOOTRj9wbl//l7nE+QqntcuILGbI3D4NXAQcuusl
U0AF5dMSnfPX2Rgg1LMVe7sN4SdJJKvIwJiWku7CupMYE/fIx6DNTHO45tUvIRoCVhDIkC9aIw+o
KS5RHn0P80V0FzxtxsxQi3bEolgKYo42Sqgh1AU7omVO/GEIDuEJaMWZFPuLvDugR1CGiqaPJPOk
EZaK144CkKL+nJzaqzfZp5Ikmw3H3tFacKiijwLI7GxUJx9UOIIc2nNrvkac9j8Kd1+kQd/2UyCn
SzOEvBnYy/9ZHqvJWCPz+uHXe+xEvhxEXlv88E3L+gcN/BwxcyJfQa2g+C1agmbPDvKN2oeWDnZO
MeS/0xUniLEeqb9gd5jbOeugLTLWm5kOZgiTd7PUYJInyjCrfKe4+bJJtl2x1ugw0O3ey7dVmi5H
iptF6pe8o1MTeHubXDO/b4BrKAUCNhL7mRJC6+z4cH4mcUiCk13j7pCNX2JzQ3YvuyStZlIbRT2T
YleNv78UYlQZwbtIhv4WZyjjKuMGrsvJMHbdWRxgUgpUh2OasGi0vGv4dNxEwiV292hLNogQbmgH
3mzMdVMgTJKHze0RZgTtkBR1XZCOLM7HOWfoM1dLkpvSXkJMRkFLuUv7M2HxZNVnRUvQqQwpbONW
f2TlRACcrZQUdQZ1x31T8bHHaVfH6/UmnemJwrRELixBkgU2rEiDfZIApttjWc/lzMeHgOR93jws
ASYr96Xx0vDGk9f/EPNnz7huIAwfMPz2oyau7T0eMSCKon53mO6rvvB1iHHkC4ykscIcWJeWWsLk
iClTRRdZjX9nZAJ3lqKgHNrh+JEx8p67UW8IYv1ThlvRZxmGgThwJuID6hEmHrkUXD76aA7iXyCF
R0w/BO6pWYTT5uNqzjtDG7FjM9ecqTafcgT8ptVKbfZYJ83Wi2sfJZkveBCajjxDsnA7+O0I4/xv
ZXgG6P+KJr3pzibQ7X3uD2RzaR1Rc1GHHadD0DTaLLLyazCoXF23PsnM3FYBYdOZm66e5PLZBuLm
8ytqCHUsp/K5S/IkavXpiUQhvSSMkysVMQ+AotUZAk0vDgqVD7Lt7032RrmFZK7tKttIW96hOWeJ
1J+5Lq56FeoOcee82LrLquFZJgdnqGmjw51XAkRAZlgSXWYndJG1IDbl3eW4Gqc2KWORyb9oJ7LF
IUqNDWXaPYqeqLj48YztQGVvMLnhGrT3AgKT/3WcJdNXMC1WlelfryRVafCwTVq6rZZjjE+cV52r
GH6XSTPtktcN0b1TGRkORXT6tmGL69KxVYjqYfYRuDAIF3TlCdgoOuREez0eGKE1CY+7sG5RP603
ibOquGBeSlsdNiJ+SVlU43jRMsNaRPB7uOLpb/NeO3nvgl64MA65ff8v5vID5Fw2k92ZGtA34K5U
EbsPyY1anHHLotXjoa28CAOpREwAO6D27cKKtaAnuwq/6AbbPIiuPxK+6udAU1Z4YkHha7AYl1mC
ZDPpbb0m28vt731xUY/ijAF3N+dqhxG6/ydjg21tw+Ziw6m3E9kKFXYxWqwiLc+DBWSe7PT+N7UA
sqJiKyojjS7hBtmMsC7pxafsfhFaSl5zHcdtQGaOj3ZPU+HH0PU/RfErUCfVE/KzpcRWHJ8Sz7AA
dpfKDqbhesyVXdLkNMHIamT7DNsUzW4CA3lBmZ/TAuxo8PdMIZCNJdkL2gWvUeFbedHk42WbJxQi
smOwh3R8KlNh+2pUur7YcEbncx4Br4AXUhW9fGGfWdkTjgsRwBL+OCONx4HGWTTXon6dpNeGNVi9
dycZVO0Ky7EZThqm1KTiO1Pf7lyg6T2krcKsEcX0wmJzfxs+1/fG6Qm4Mitw/nEWTReD4j3fmPX2
U6m4D/RtD0AfPVE6j8rlCfzSMszfs+cQZX7Ba9H+ZRPVFiDoOlx3bVgqTTaLltXpFGoyiIt1+GON
MgBEzK/tQJKADrGliSQurqtidJoXcQsCkUGYpBShUQcvQCEg6oEnVY5cU5F4Hwwy5oXuys03P9FF
fv7y5dz0Bj5ObXsNG5H8wVoiHTLu4lrQutOTvM3kfPoA1OfxJITRciQyssbYVVDi8fY6+4L2Efjg
+zjwcCkEjmYGaUG7Wmlg6j568jTYpParXYjBA8bG/sORbx8sLiKCKjmwt+JMF6kn+8oLbm2TyI7Q
6MRBoTGlgnbE1A09A0vyfDVZoByRYEwDdtoQZB/RSDcaimJZM4D+hJW7Ca/7aAGIVE+sO9GivAtm
Cjha4X9gWb18H9nLYXOPml1NPWIBCzxF3XBCRpaC3MfV+h2ZwlKiVvc/djyt3MjUqckMz3AZTLX6
UEfjgkTfFJBQgzT+fipgygYK1dPkuOHs1htwAvmMuj7bcKzE93JwVyZSAZIVDhnTS9Eh4RIhJaIa
x4+Jov9+KZJpHBiBuQfR0OmJ0Q4T2vPf0zyK8rjnhhMHDijxrJUZKcUgYRgWi5NG5wehU+q+OJ20
mtcuUhGguQCKHRinWWsaWNyeq2GGQWUtZOdsnbV3QGmPY6xrDDBpFOAOKj2npI4PvdjrPlt5CBVJ
XHX/iLg/AfxSVUowmOy/eE1qRR32QbPldne4lAO7niHonQ0Q1PQeHZuvWrZhfPpV95qkAuZ2B0eP
gPFDXYGeQ5eQ9baJlImOuxHR06aypmqIfrqSRnp17B3DEYtix7peyRDEdBJW/atVpag0g1PVdbUJ
5za3fbjag3a+3ev30zJa3KDzU7dEJfBrTEvru+DeNlAxhB/0E+eslAOIFod4i9wKM3dY4X288bM0
qgztFUp0CILAliXj7TBuWr/5B/YIrYyDx9+Xoi1OgWTvx3i5X+I0xg9vLpd47hA0fMcG3ffk1IVT
OtKuuL73GdD1l/WluH4Qq4rIaiD/kbCTwGEd2y5cyxOBvjKmJm/mVh/VEbmU75knBMx9EfNLzq8p
g8diCtEhU5Ulf8PVeQfNNVgPJka/H1f7suKA5wEpmKSd9aR5R4zx0uzXgkwpbAy7FisSfVwhHjHM
tksfqFgUc0W1NQSij0/bJqKvgU76bWhPH7xQvgCSXUDgEbLcyzC+USUbKAk8NsvO2lLvHSKcB88D
fwQKXift1UNndqw87IpgFuO3aC5zeDO3ObZXyK2LSokeJ2E8Eor+DJz+ufyAyqqd+rmAaKDzVSMf
7iTy98unT5/KuCSaliEkZtQeVOZJPE/Zg5P8vBnWq4nyHazKgNhQtj1a4sk1XKp331VaOFpXQaZ3
WgFzDNmXLZXunYLSuKEHvxUgTK2J32iJfIQ021il8ZX7LL325MPxd2rk/mrl9p+o9CWCvCRa79rP
vHQ2oYjiUoLVHj62KbakMV1A9Skf3QTi/yKvWU/MeHccFLdFuktIwlUvDhtyMMKPL0c6OjnSQhE/
ze4QfaWN6DPuKTNK3/yRzWeVGZ9sxLFu5S26gV1mYSvNg7TYPgVUNsL5yZWUMJEAzb2KykSZf7Z9
FyVJbIPIbxXXh68dvE5Q1ya+gkw7Z76dyCVUa5IbxnggbkTuGzAxaRdA9usvc/YjMRpsOI9aOnwH
/QCPkvKBhadIiFIu5r+/nUV60CwZ1RJwJ4BagREz6lWJ4E+wiuxddEjDQn73Osww/Yi07xyaQnVE
SKzOjNWee3JwLeaEcZSXr8IEWJm6udgVatelanlWfmxnxSj4XjLe3Q1uwMcuKYf3FnRQ3pLqfGer
9Stcv1osxwgWiQxdkQfSo1884UmkU5IpS1iraeGCKotT2v+TaySh8Le+EdVo9npOygdcWyVh1+0v
7XvQKjej11AW6pWSelrD5zIkBnDTehgxXa0X9IkCqqyM7DnVdfcWqlq0sLm9otGGQ3fAaquUpEnS
9P74Uv6I41DrvyOlPMxZmQmgJ5wgvdxE0OoMiqa9goFPc6NM9lXX9LofQfOaqw5eBjG/GKkynlwb
LdsLCrn8EkgPwPguu5uw2JJoZeHflhCd0U+ny7js+aHOFL99V/iOPqRagrQyxcwDpfls3xp5L/ty
lq2poxMuujkVzJeYtyqp9+gB/sdN+AuAezEfZYJHk7SIjsde2SbJ0JyY/fOoVwqOYHShyIpWDQJX
AMCKQwwyer0ksCaGcPsUFrGdwEgUWvhPaDsG2lbvfKLEwL18dWgHSgPe6BhQCpAFaeOZsIQuFIrr
1CX2ktwdhLss0GMpa67STTh1rzi56uzxXLtg5ymK/W2BVzlH55+Vk1LpXQ5BmAy7lq8Z8qnSPbpG
f0K+Jeo05Bv3pwZA+qFiAXfHpJbcKPAwXWpxOIpD9191r+LGbo85NuU3zMZexFWRNzQnJSi4IVjT
KdManfNIOXL5ftE46k31T/MUNl6KoXhqc74ZFBBjzNfEjgkIe4CWrtDX/VQ0bXbvtUZBO7HHNO0P
sJ7jDMaNLWDSDOfWMPU598hdYCTgBCx+MJaai5Tz+a+ZVZGVf8qBVvMM8XtBekgdI0a8Mv4EYzKu
BL5YbCk2P89YEdY5tQmiZZZ8lTm1vS8mquuxOw5V+tYtIcHuagzV7fqjOR2ApfjAq4XL1AQe23CG
jtHLssZo5V1/1BKhYD/ipdQ2cFMblMWB1Z9/SWaig4v9XEPJ6TQVa72q7v8/F5h4cY2v3UgXxEp3
QtQGJgP7swO7yfhGhFTrNuTmR0WYSTIenA2BiJCpIS8exDCeov5/k5xups/M7/UEaiqqx/CbAw53
JhyNt1YKZrLuisCLoN9+t0ITf68NSlFiiYjHoWQtGvX6V1TqwilsYvKi+UL0+JFY8yspitCBHKf2
9Fzk61NV3MrXNJw8KLWMfCmE5xIpTv4h04aa+vgiRrWIbj/QmrvDmUq7vtgiVNro5slOWpDxWzOu
v5o3/xCEoa6vODGGCKXCvpWdZG4Vk5LoklCWyPxO2fhJcSEx4D04URqq7VQQRi5KJz3TldnR1Xk4
0RjpBt7nqBTGKV/kOqS21U1XOTNENG40IXe+Nuf6mN34lRCoqcSki8fSVT7vC+LuSYmvRWZMKeHK
4akF7Rb8HghvzOPof9m0poCwxiwoZVqXNnoK0pFBH7IkNR+3abtb5hbC9a2Y0QtOABUuvs4+BcO8
z9GbMMCO3n4/vETZDUCy3dqZ5Qs782pL8mzB5ETphcbVKS7DyVlJ7AIcu03uxhQZwgr/Bf2IXhVO
T6i0CmY/s4gTUPPliMwpOIRbzl060eFWfC4vITYXajpjMKv3Sp5YwK/cua51UlBfRcB59LsXop3U
GeXe6jmbpsjiuNYOIObuVjJqIAi1VGX7D2nZ39yjVhJp1f4aBnrmWtqCibwMqtSyhsXjQQD6XrC0
ITtRF66/VK0ts/TklA5Dgedady0DWKtrNKJY1lQeRGex/b8NFMOULznc5mGG1f/xl0qolmndw249
fzHpkRp0n8Kc+gWUGYLTC0bBGqyLRcMsMz+VCINq702q0RqQ7KdtlwvXsvqP6eQyNfa31vhCMvaW
ri6lubCXEtGDjvrEpgjY9rxVdqYKv/Rez4Xfw3GbGOy3LghZ5y2ZGdsfdrpnW921qnLfYlw344K5
urnfjqQ3oP2M/5KXO2haiGHLz8fVVZrExQagd4i8+RTHdeIjvJhIJoNlrqBZ8BMY+t/LU747HUEn
/KFoiNDSjrpjLnMfwv17luqwQyDftHtaBT/07HJU8fTCCWiIyHQj6uMieyX9CQkOc5HhuQfWeFQP
TNC2xk7RS6Q1OaDQDGXtOUoFCql1RTNV09ICt9vZfPQgnXCpfBj+fVh3GYzaJFAtD76BczjVpEbn
nhrJM+Eaw8l3RWx1LdZ/gNXRgp5FxZCovR9CJJ1JxmgbcaYjVZb7zaAyVqS9qtFOtVW/4nX9OgkN
BuY6vrFJGfAhMocEBZy/DZzsYRNZFYkJPZ7nSfFr7nhaltbKDQMAaehvaX+QdJgITr/eGkUX0m4G
K8qVaESBhWAIdvj14gwh9oUu4GVtuLYdQccytKd4yfRxYhI+3ColsVUDLKGN84gJTrfVTvaY/wi4
CNvBmTFR4/CqajlO1KFMMvk6mfS0pv/OFae4TJVId/qBypqoeC4a2dLpRmQ86+iiLvalY+vzoaIn
OxXq8ggV8RqUfVSbA5C2AOJ80aq+gJ5elUwzwFAXjPm8IwbcQCq/+wI43dITz3FTi0NGGlQKwZp4
MIPn0YZk+HVDy65xyqtzTKvQnxdUtAYn/4SBZ2P19sTM0NmBNKZu12v29m0llxTvbNOnk0vrVAHm
zle8MlXX24t5wmW4hHZP630zyn1vSApbfKwI53Y9yFOr8AcOX/Dw5uhZxGeSOMXKXZIDbbd+gDOy
2JjBzOXxdyvuP/aVwySgl3O2evBd0ADup6AFwkysZBejGmYhZvR/CFYa5V9K9EwtOuB38QH2R9Gi
ANbN+FzrfzN0DqmwkpZOdRZI/JDUerikmFzkklWUcDIeMIJfVhXxE9rqXT8Jfdb518huXB0kUKn9
thxDehhto17A6emePa8Lk/pOzq1kF2loNJh6FvepQdBtaZmmcoBtYdGT2nfA/Ohi8F1NhT/8SKGf
/20hTmDBDXEKAdPuY3yMm23LcfNNwUdh1U/1Z10Ty+t69LXVWXUGElHuwm12N9BX81shSzPEWhHm
2sW5axQbqq0C85L/HG3DtO9dDY8waAd8FYmKSiQ8RP9ruL/bNRD0B0K205KvRY2CzPdy0BMmAJSi
9gDhmL7An8Pcl1k91czpnSDP4NpidLFG6ios9rfpMnItzod1rx+2u0Rvj36AhWi9YXKtM8Zb8Bvk
G3vNl2tk69xaf+9aiRKSMbA+FYGPXxssOiuRSDZmd4E+Ov5lhgdHHByEVlKyXdwUdTyHU+JT717p
osS/7VwLYIkrM1sv5SfyuD+fqb30oUCtce8QEefdXObWwvGzdaN3C4ZSgxaVywnUmdnEWxmp2bbR
RUcO9TEjTUExorgCam5OIbrf78VMyN2u3qXo9VIN624PzxbVRoqKW+wCqcGO0J+7WR+7cLJ50V+H
bPVYBCZwuc9skpv11ND77lpw3G5f3ncldAkvx2ODSRaHPiZ9U4YnQJQQ4wv7BcBaCPW+jQo1lZjP
X4nwnfK+uTg/3nx3DbYS8+fI99O8eKkFzuuBJuJzEAuJonWH+8deLjbxTt9QT1G3YsSenqrjHXD3
XZUEib2+/Ih2ngzrkrTxS0J+u3jiWG4ssPo7cAm9oS8MDs5ytziJBRkPewXt7QMfzrxx+OXSH0XH
/8bXGnycgHh9ovb7tAH0MrEyYl56zsqV7tM/LSNAysVAf4JZWjESLqCagkA+TtRSaS+NHHpRPIG+
h42W3ZUFFzp1eHmOnfK/GjfNRhQn5DehxjifXNKRKqsk6ccIPIo7MB3RZNJKvvsdAH3JkUDQcGdv
xqsDjJleC2RDFia/K8Kq5+9uOxQxynzqqX1pJdl+/9PyMNIC+tuOhvbPEWr+0uYrHT0YzyPCko77
5r0RSEf/KUyBWDI7yH8US/AwQNAPe+mCive8LzgRpuOY2TlhStgWOYMsk60P8mYg8o8VQVOcE/aa
Uv65JevxBkjTU6PybuI1vq6B9JZrX1scPrfObeT8a5oIFTH7Az/WEkfwUwDRJUMtnutC/C8PjbSg
FhJxRfuagCekkRHQ7jffrGQu7kHfqjhfWY4Ym4DJ23WnCQgCyRQFT2ZK0Z422krr8TjIvPMoETQU
SmCNgdPOFqPVsC/3kkIRaq3lQ8NgHEWamtrTdqpvfu8pOh6Q3Bua81INJ8z0WlMr1ralDJ9+Z24n
5gihEmQtI3T9N7dsKLGb9o7+BPuA8jQoF/SLNwDpFb9WYeNkpzwvM1Odwp9ukH5+ar4sYSE48dIv
TpIyC0x5cPqdnVK3qpwXFObkQOO546laOa71UHPiyNhccammopaOtpXq8mc5NrYMhxLC94LycerD
anRJFKjSo1bwY0vL5DuLA9Cngg41csdpPw/JyMDIVVjGzI6IRIGt+N/GmERPEnzZg1zjiq79TL1E
iJV7gR12n43a8jQzq/vanXyyu5d4QqUVXhdgnuWXdmSSxbIYqgM149LKZxQf719RexR3ZigKJMBd
jphfOUd7yEW00Azo4royyHmoFs8/XKJnQ6cdA9nnC7pae0GG5sr9lJlQH5pkjPCpSn+bhfvyS44E
d8S8NPGEAKr5o62a2CSy6+204Y0qlkJ8igJlS/yssP1J+JY87fQSDh1gA264zqaZ+WvIb9oIOdKG
sKKqnDOwiE7CHPHD2B9wN7GMMOHInGfeF4FbKBgLecI2u2ZQfce3luRet0eJEVT76vTeU05X4/6c
l/bGHc3jIjZqy2DHWOiL0qXMQOVhTu6CoLpgJP7jyTgCilvaF/xKXWVnRpdlU8znnFzxmOwwgwlO
r6UlrwSui52yJHCaCGgSrQ7JpTGyEqexsuVA0OsVuUR9ATQTkA8SHM1m/KLZUTpItGdFPY6dyZSw
ynGXlJxSjs4bDU6JJ/Tn3U9NEqkn8mIMuUjb38/spOA9EM2SqiSgd+Lsd9aZtRuhhOieY+xl6UI7
Jt4zTE63exhCkRiVGppZc1IxZ7ihFKBQSYCz6dq2iSxuTsW6/yQz6RMngxHReITEn6tyrIj18UMJ
svJ7s7qT9AsplIsNcQuBUSCzfnL7WUQ+z+3pZkkB7uh5IRY45o8AzN0I5i6YYRRqmfkVSZeQ+7TO
Y+KmZDuajGFs6lHRaGIy333/aEh98TJjU45Sp7cWhEkpKVvCNwCCBu1eCdcKgd8y9uQ+zO6Mw/gB
mt/qSL1bWOc5QSlMV6YhVHSRy9Cr6uf1anVKaEFmAafgylV8U77L4D8EmU9p7TDzZu2ivyixYIkA
vpHQe3S5jR8HuBrcBBK1hZv3V5zzpHne1BhXLh7hL7oqAjiWnindbuC73wBa5Z+hjkWK9KBQNWDN
ifvm0614gOmeSCvaFX+LLroi5K95c3tiM7kJvKTj4+NtYSdwRjkTB4P2IyiDq1r6S4+PItgKnPkC
k59+KT9Or5Mefw9k1lOzdlbvnqLC3XfctN/C6arc8YW8vL32G7uYoM+FuoYJg3VzUM6zNlBYY0W9
bqNjiAJ33W3778KtIEeLYgu/6N/oVOJAUlpIlZN/7M44Didln1B0NosXYHR9fAkZg7qdEnyoW/l9
DSY0+NAheOBX1Awi00zlGWJLm3JuG/dOKWtIuiwUgT4KHoxz6U2IwWK+gfFHI0dB//eMer69q9bF
7R4EB0OgGFDKAvzCXFuI+Sx0+mA7ts3IwMtacnExvro//3RnMErsmF6BrMlypTLXQ5LkXs4L4pIa
yprp0oauV6PxW+SQ7d75Yw6QPfWJrEcH1nn2NuJ9DeN5r5M/f91/+/TAtx7Ielbmtj3asAJ3mpLC
2yLtvTb2KmFhOShQlI2bjfyxJ0NA6ivIPxRJiq4+mTUo2MPkr0G46htJsRq/bVbyE8eqIOn1IVWO
Hu8fsqfNuAtp0ziC63w2m5Pj/trpS9UByCdXlxRcLAO9Mr6mRNEhquiY1Uso38r+5TVqXHZ+caJc
2cJR6JFbvnMwp/Kf69TRulmCBSPB3WLtY+BypRYSAPZj0kvFzSdVWV09rnkJLYQwaAMujOfI97ar
x6VdIqu8A2sE/U/cMGNPZFNVhAjihVmZ404v8FxtFcoZgWyfBuJyJiCzFN2oH6vwcXXCvaMqN56m
OdqQHeWH4zb6gredfxhWGvNdaSUvHsz2SKlpdtOs7x00EaXaL4NvM7CqYWjWAPPD1En0JhAno7JU
PgTYaSCLGYuFOjsFE+cjxr7IN4f0xWhe/eAi3vLDd84wHNGwzklM6qZs1TjqZ2EiSzIQIXXirh/Q
B+SfrqlRTJGdx/kkzZYHnoR+NLuKcC1N72zVRCJPSVRKSUzuPkQ1dFlTC7wNeXBG7MnjoYHQzZEb
FYu62AnGCoeYUjivZZvx/m7Tm8MF3a6FGUAwIdDv4daETufq5/A0OXz691SRFV807ZIrzae9993r
hKUtcpDUVSSllUTXT1K8dcknZ1GfnYpC22+kxR1Dws0IFzlNMGeyVBMv0NjOO44M+ALhfRFluRde
Z6Uguu6yw4yXb0eU7I86tMQ4b3Rpc8ZqE78w4fpkWpIVbbS3LxGI/vMQ7ytynH8o8DGt8xc1vv7X
ENSZJ/0HpoiP5Svuu4Fym4hWWpWbrMphduRERiTrLEEcX2bXxK9p3rK3r/cA86UnqxXv1Yz51nvV
bry4LJCgfS1KXLir3LqJ/L+D6kFUzutpbtYd352dgCdRRVGF2HiRc/IfvYEMDucBsUTHx/RBossE
WnjSryluM+B1K87YdXeo1eornCnk8i86aEWnpwJ84aXo1u6Uv52j71qYTNpFRQrSpgRcibQnvFu2
sLuIG8bRXQAOZ4q1v78gvCx+i8/cF8/8NqWl0hYUOD7a+qnwZ94rh/UommZAH4f1I4p/vWCdp7/R
Uccbkwz4b3mPPoAvcevdmE5PpHeH+aQKWbnS+4qtFP5ZYptiZiXV/3SrE2jjp4qTFArvmfm44BFr
FhdzhN+UTXAeTozReoQjnkgHCQwK+XxpJN2x3lkQ+x/0FZ48q8WFJlSSJjpeSABQHuBONKvg5tRO
aN37qQ/rxFseA9teYoZ1nvQJLVlOrxXBFXEDWE/Q5JGzD1y09NDli/nAJSRlY6igEWNq04UB/KBe
pyxKWG4c8x5VtYoySbGUL56oD/LuB1ZINwK0BeqPzYZ/5qm1+mvt2EMRKGMF3tS2KTb+ccUfnHKE
QPi9SNff8MkIw0OVRwGINRm5VAXOgAfC7W8eHCyXO1s/GwHoL/wtShyo7QrDtj1aElJOaf4/6YMK
k6G4zVN/HPnckogQS0LFYG8V4COl6kDxXUaFF57ycFZiKHnQpTPhjCDBX7Anf4Yt+/xh1JGoqvPD
XXlbJBctus2Lz3btCcqPJ7VZHHLxeqZDNTVuHg+wbrnv+FVLN1ECZQ8mUxJQLaLXsWZyc2K5Zz9e
q9jSrChBCfnqZwyU0CNfPptXNYynHCwctGaF92NeHom0hz42sb/ME27KPZix7e3qBLGILprNFqV5
tFAZnzglhQzaz71Wkbj8b/pFwT04DLZZPAQHQMR3YEWjVbY/vseWTQYXU5+uR/JpxDbtmU9nL0LO
ijKeR8fQzL3KT9XekY2CzZJ+TBcnkcAAg2UGnbH2UY1aDqV4mpI+o/Wg2bucnnfps9yFBQZhJW/Z
Jjnky57KLeaUTVHCYH90xJ4sSQxgWMcTFFAc+tuuJ0VitCWzxNQTrFzO5q9AiQ7iNOyuv+xS2UaS
t8hXpqgd1WwgCWekJIOR/pRPTAZWqiBzLaoVL3aQdHVLO3W13dzfm6dJP+j+yUem9FTr2Ls+QoMK
0cbLWn4e8jA9Jx/r1mozFYoVHvPV2URcC66Tu67PljSqLkVMoc2IebaDOKwoM8AyRurUPduHN43B
ZDozPgwfTYOPpCQcqR2UC5xyM+igeIRlsdtDwohclcWSfsh1iwNpaqyaNxZDdmv20bxck5Z821MO
PqCJzSvOBsYypinh51ERC513yd668wDO7AE3DkfAhBz72KnkFxGY0X4CQFCIMQPPnyuzPu3evOgR
Pvz6AIJS+2viyGgv9FBFEZfmY0X2a/P5BYBk0xFywFvYf8ozV8OZ7zTH4Ah89LzF+tDIWYrHwt5M
YDp9oq63OeASVQqe6g1cLBrLziLwRKm1Rx3A3voXX9z39XPtO57TbEhjRr/AD8H9fGB3G5rKPIgP
qu2YomN/5jVv48wDd9NMAuGJxAQFiCeG+qSzxtUzS06HRNLmcm2O2bMW4/vjigdXxoHu8/2q2tf8
16PvtmiOKeJqT+9XStu+dmeXFIQtWscGiTNcGTBplOcgxgRR8PLntw5P1UDhk2865j1njetkB+l6
YWmnlfRXYZlFj/31VEZ5uiBzhs2n6FQVVzXFdbMNBk5pHK1tridj4RCnVb24I92Yx2pkON/NmV7I
HBilaLhcZn9pj/Dxb7Nq7NLmvtgdtfYoEmSqOGx1cdxWghsjMlutqjqBINRsQANGiDjsP6zt/G1K
uy0IlrCc5pgFlUEVs4EfPqyBMHGE32v6D4/kbDTfJtuTOcmhAaCdt/KpMiHdYS1uv8VMY7XffyMx
gN3T3eRiT1Q5MEYm5wgF6iPGpiMJ3oVp/uFrR67yCEOBlOf/2PcdkpAoxWhJcpEeY2zqSYiH3h4n
8DJNy128ICXvz40TuTBHOowpisTdxB3hCDOQvPHVpyOvIFHhG9K95vlEREp/gCIqB2gZRFjx33RY
osSoqjYnKhwj5i/kI6+/uSxoL96wErBKKjsN41Mc4UWs7InAMZKKSaXH+0cj8Y9hstc0p60a3zpq
uVpYLrhz1GqSfS9zPLZAVp/sJjkWxJl6lPe1I+j2lJ+VBA3wTLMrZ+4yrwUdazoMsK5kunogOGbF
Tif1MIPp6PsqkBjcwRttZEGzfP4geJFLM7KdLYskCXNT4b7P31ClFsRpJU27M6j088tvW7YPdD3A
uAYdv+imAE1AQJPg14iIVCTZUeanfDwq+S7kvrh3dEJAXMZcYxbKWezGBNSa4/wLeZqhuzBs+lag
l96xOmZ33UNCtZm493n5JHhSuj8UFGy1/MBe8EG6F9HvV36iV1KXTNYTi7S2lg1WdcamjeBT/p9O
+aGCF6/vpDCg9yMXyz78ihs2/jDGT/lZztn9iYZK41tFe3khvwG+zrY/BEsFAG0NrhgKJSoMbkHS
j5r3lbr5nXM4vPinqM+nwQD1V/6OC1AvpmgQuQgYnDrDokQMKOuLAF9Hl67S+UIuC42YwSz1FlHo
iOUOvD+6IqHxfw6SkE6L+0SrtfBZfPKT4KL773AND7eFKmXP77rvt/icVtkviOQiDeXSbMP5SlVw
fUnMw0wFTFIeyDEr19ScffgIjXfUHRIiMoNuD0uJXBWSVY3ctVVapjQ/Qk9EQOXGq6a6KtmCLlnc
g+HailZw5pXcqAtlOYYIuhETo6/wGnLdmU0aydh8wz9D7kn+gTRF5L7jQgwCbxXSj4BS/MGSciJH
4B9haLgY+Ipopp5gTH/RRnuEq/vw65L2U791Wn68TKwq5DF+nch3GZlbczrb2hM2dnUMo0QJuSdL
mH5KJ3/sLfJJqH0dPnpspYOXXmpkIsO3zzuUixKcxdgJGwavLoFUe2RCVNss0k5Gk400tbZ+zzr7
MZShyrlnYE7/O3KbnXkgZPO2PEN5vPhr67u1a1iQNa3ZGHIQGdhaKCS9BIHi7JlzFnuw1S4FTHq0
XeTlF49MOip6ijF+7zBrDPESHSELpkJtweH5fDdgon88BUEJOOR2SZsNR8DvyS5nEwexePxl23zE
doW+dn6Nxe7uM0OBqRl4rLV2PpC9MqxeCnXRVTMsqhJMS+GoOo7QXUoNEPZYGNVmfjeDvTMv4HL3
pKXDmhzsgXXOkZYmwb7gk9/TR0QD/o+NhHe/PIj3Vmf6IzK9h3gVkAGQqqccjyh3KO/RAn5acGrf
UIIyjAPhSTo34b94OOlvKiJ9kDbGtnd616tTuQVXshWpHQ3F2Vm3ng9+ceJVfWor2HvIp1FgSzEN
Yk2uSMu5cCko2OnLaxS8+Iy2qKB3NF7+8Y0CzhYH3dTEqrAjnrBdb+lePHPua8Wc35pQOwHH2B+O
uIvAGTWrk347sfb513DJlYEYervrjrrhNlbiTHZ+sHaPpWiO/MNooOmr6RISdS7OI9Z8bMUu0AlK
9jPUG//sKtXQ0vPZfaSp9ti0+3Sa17uGSK2FuQia06oZTE6J2/+eKgUcrqcTxvVmwBURtvdx9oXx
mcNsyfxNeBx7JrMBVNB68iq/47NgPZwcoI2Kr8k8WEaOW6+6PQd54h6//JHmPSP9xbl6+sPKv/LF
9Fke4r+BmLpTrOKHABaJEX2/7qfJlm646o+EHDfalG00czRrKuGwg6g9qP9C09Kx3P0SWBtIgE49
efQtkHCRduHMEg6YIIX7hDs3MlkoWUA4pXAr/ZjzCxpUiA1zjwrb0WwexpbfCanE4PXfBNmhgogR
9Pm5LvMg0KEb7FaKomQwbpMziOH6G1uADRFL9KkqkwT1T7B21ub5aPi8eYDXweTbPi1WaKju/4dY
Xx2jCvNh0v9wEj9KCqQ/yIN8b0O7n6FROZHPuPrONMa71Io/4HgqB6B6rN3qnC/QNMQbil6Dg2FU
2B4ciUI8iekmRWlipI7peZ6rQVwK+PHc7NeaGleF+GiIcLZo4MSqPURwBKpHtnKcIdfkJLDh+Oav
cQJJ+cdBqGJJRWWqXXV2xOdiQt+qEWkHmB/kyYtDX3Qcn+OcqiegYmfcNubXsyEp6CEUbh3U0dNN
2bexMvA+RQyD7jtXyhpbEw4sJdCRyTvNJ+p870nIkJLsjLStlOAfMBGrM+Tl1wpHeCOAYyGrZolN
GDUfKgNo7DQbkKcapo33cGlgFvSw4PQD8JXK8hz3cjWgkTHbXpgEy4ool5uiVgGYvmfy6zlKAkDH
fpYRMZC4we5QDm3BoCkeHkF/km90lWXlfUcsUKjLkjh6sa3VngWW9+kk+NFMqm6GMGXrHa/Dspf9
uo9tV+hlWgUfIJben07PbzwyDxSRa6dtdj2BlClb5c67j7AtV3vNSjWYCYmqKfcdEZc0CcTA2CLa
f2hzcTUo3YTgb0pHMy5fxesqfoP0T0Zykan3DfNIZqOM/XYwim/ydB1sRtsP//wZPtl7FxJOx+ti
P7SCo0knZbTy1/SddLWp96zsdcrZR0klS1RUWTAPOxYqdKrT+1swM/k7+tVUCzfhV2I1AucsFhfM
yUNTiiJWcFmfOkIqhUuO9pYOwrbvRmSKo5ZI0yH+xniF6jsa5YKjFQ3pZtUsNl4ZIYb4WzJwbo6a
oW74ASXAWH4nGUfPIN0ARzP/RQw05MAtIaMPaWLLu7bbQ5AdnvGDLDbx72SdvH9feGJc6K1MuJJI
u/UyHnDrUxzQo3k9ejsyUEpTuDHZXk0YQV97MwH6m4n0fwPuDkKTFyZkLX0jViJBs+K96Afdp8rr
wVBJs/au3ThG7W1D3cmQJxy9o2Do8r7tGbkE64+qxEHYJsayUPGBOEyZVllOOfRU9gldaSvIUiz1
h3yK9fiRHzMlNOhimlT7cGeLfe9TH+ixy+kuDF5uvSe8QVV67hrogSq1Jx4RrUzTUxvWkUadvv4k
EhPds/1hrY9YdkdaHixiDwmMhQI3oZY71zBfyvf02Y11hwgxrW7DJGum+x3CeWB/Vc6qPu/nb/0q
tJIWw5C8B1JsaCPv2cLESaON+oZkLi0I9YdJF0oNpGS6Aq354prj5ZA8W5pzYdphFBG703c7UJ0X
QUMuEpOW0JPIg0usKkhH05yfMND9Mc7+ya7fgqwcZw24EH4rkJg72Kvto6/xq7Y5I1ugu3r4p4cM
mVeGLVLo2BQ1GmtNxsCeXmukTWI6aHvduClon8Tu0sNcxA7R5wbZ7ZxNC8QWn4IuPz5If3as65QH
nUeG2rvc1OpuRCgkCV8dLAzMgLiy603Nlv8hfMwFcL1a/jcgd9B1f7t8icHCN4hAZzIV8MILcnKH
gQGlIEJZiCd+i4hB2odGxg2WXSmdC5z6nxcadRVL3NAC9FhmPcbImoksDmCtWm1r9louTgmrWOGk
uqjUg8y6+nKJolpQUFI8iE40X2sLdjJu1uYA63tfMwX2wbzvVT5O+zenq07t8CorVlU6wNEqjbqY
T/FagAn0ikCGrOkxBdRmbtrBMhfUKLPnxjWXKcJpCXbXjM6f5am17KUCl7kOZRGw/I+NGs1lUQ9H
57pWOeV9bNAhb5xkM5W0Zfl4aZeUV4HIWp3suFkDsAjX9wyDZpDQwADZgsZCXzoCJTvuh7bEHMM6
uEWPaL3t6h7idhiM0Pr9ZUJERUkm/+bkR05o4jMOlSsGVeH9L/qzb7KKQzP5bNw9xW87NwvuvxKb
apgTpGyaKVRZLCBE0gpI55nI1qQfgsj3peCGKBb0PR/2wyU30chbKsSTE7VBcKnIVSN3aBy5HahA
6rwhxwG0bqtpLq/RpxUcp3Pc9p4LdS63/B5CDXrSIG5BRNuafpwb5lRB9DtUbeHY/tJOnH82kVri
HhFMurjIXC1HWlQBBj56hdURQn/u/RyFguH0kmMtXTs6G+ZVsqrHoaKmTlj1xqRtBSli5DitUU5Y
UynL7qzojsy8IthfpomVMlWOHtpnGCWl0wWcy3n6loIZ4hqP2lVPbgfVM7b2EVrk+9lhceUJtrLw
nEyhyiR+/FbLzqKdz/v33OiRhtCxg+WaqjOfgrM19zpECE3HpCR2f9U9hqkCT0vXgphDDgs/vEFn
j2sPMY7oDNMeBvl2rjwIpCLOsKwZUnAVYyATsWVMI0MwvrCD3MhnjuNYRjdr0aRGToYPEchsdffU
d+pncDOIdUIWfojQUH7g5GakdrUgvsO7cSjjy6X/D0v8OiVwQWAfmQ2Ccbq0Hz+rD1Srlob86dhh
btEM3qB0Gz7h77NZT8sS3pJ8ommwwDsK/AVrg4zV+8nDm4MwJpzNtQHhvqxFKoeYkGsya8AVthey
lWf0rOsk5WLxeKZUgxyorIIejPr1FeYzX+rqkrM6iqQpV6FNm47GG0psXBVveQ8rogVb8D6na1Jo
U58znZ8B7vUOgdNzfYFgLP5v+SXvxedHMPw4GpQST6k1ZLyLiYOtWpNb0y09dBU9J8z3t2vXWBsn
0X1+ZESUR4oimoBywOuBPlE5ljfE3e+31xMbTSEsuTQ+SFAsIHQZBvoqC8jOhdK+zAspDABNa/8Z
R2bJF7UfIIFhDwXYdbF+dIBxOAP6j7usKuDPIW8pkGx/kdkNhhO/xAej/to+EBUISo1YT9YK1jox
Hhz2b5gsDIdv8wHgOoxIlQqlJIb0dHRk9GnGXv6qqBoJL7n+oCqCGs8vwz2hJt1qo5oBqNjuU9bc
qOhK6FXmvkQiy4ZD13dhL0p53gWL28R3guF5TkLP2mohoA1dSwE66e97fV+SQ3WvX2qCvAbJX/xC
fb06bnKb5DKA2OmGSQ8vRN8SqK/UHCIg/8mQ2XURj7pVyOXKe+ix7A0Dr9RHcwBF1atUFZoXnZ7O
FL/k5IR4L2HsDAw6fWJdjO2gHg8qJxiLEKiDHlPHLr19bNkw3aGA3b2qBp+ISIWLBN86dxt2xcI9
mopPQNORa7HYXAc+X3wJVID+d2IcHLWx0DlYU7Nks9+mcV1Gonqst0Ib07bkt/i7zSoPp0MtlwVt
rAk0BSxidYFDxAJ7dIFBFs7BuvkDoyIlq+bdLMnhO/LiOpFYonhcffjZQ6ZsAKy531C7c8O4Is/t
0wdLRZa8ft+19JhJ6RB9pQAcEnF5hyPOsYOBwCF5wyeSUzKcV4b62b3QFjgcxXdbM1VdqQjK6fNh
pl7r+/WkGfPPAcl3INg+D2w5jVUwLLcpU29RBPJknbAOvySnDk3gOUpY5gLPHIsNEqSnEuiCXE77
pJe4BlPG7G8CrFtDEjV3rkGPElg6os2HwCSs43i4QNEwZSnwse5Im3DVHKpolUtLnn8ldaEMMY0/
T0whbbrPmKJWSyC4Diwz5EHu8X1fQeEJw2jeOPUevVrTg4gQ76uKOZzGf7+HE0Ceth3bw1OCXqyZ
vm9N0ruEJ/vw5ocUOzPbQvRkWxCvRRWv3EZ501lk1K/47olBAMs6nPztTORELc6fX+r8/JX1rqzr
gXys8y7x0reTtTZgUT4Hzza3NDQ+TojkwL1MELgGYBw/R15FkIBiK6VGR4GlH87hGk7Bv7s0kwkw
9VjwIxAUEEEIMCR5Hy8lmgm57jIoEDPCyeCqxY4xxjRGUCHz/Hig0HyizAvJdssUVRHhy6ZCNY47
rnbVvgnhZbEVaUk+7fLCZtFzw4o5HNbJsIKj2xqmbDZSXFxImyo9XtLuY5rcumbdTGPSeJY8xPw8
2/I9nC3xrm+a2Ve2vRVoxx9Q1yPayNCr5DpCrJgxplmCjHo1QT0Lc6szM+XcqnQlruiHykBCN0O4
2tJVmqSHo4LhbEDLh+FI6E2R9aqgfxNsHfgR5sNxUgj/WeGSyjV70q4kIq6Egoufz/hpAGECMVah
y8TVVf7w88s+KlZvyJcd3wJIWrSPKmPJsfaqG21eNUMDsVvc/aa20EwQjSOHVUBfQt0rb65E+dhG
klPQFnxNCOcztQpACPDO/12O+GUR5I+ZNK5RLuY6b8hhPGej3S2txao+H9FaAXC5XUXhag0wzCx1
Pxczmwpi0flQNEBqyswaOd/N1jpqlK1lar555ynko3lLrpCELv8MV6QUId9Rr7SBiYmmy0B25SFP
n5158ejDgELNk9DDuxpZbtPWCCvNNLBXrIA2GPKfkx28omSlU+GexJisGvoIDQvRNLK9zAtIdZFO
nsYKSqwstaLAEmCwYUhYWfxrvQEUEIk7KG1fRnuF0eeFaedOtrBeqbJ9jSJOgM8CeT1f2riSyPog
QxH72a+XEfW2Iv8jD92whDI6oq84W9W3/3/x47vNusyuFpiAMzaWJv84893JeTNfi7yeKpsi58AB
bsrvLAi98v/1mgBmnvwoq2aGFx7Air5saNrxwxIUV0oSL43IKYs2SMu/wdKjn6AV735tJ/FmNVOh
jBR3xhEpBVA6XXl8uaOwTXYrBppGKZotTCsRrzD6AIMGHaf3A+40tNp8QZ60OHSfZhkggob+4U69
BrMhW0Gouky5iXKVfmLVRglGLy9DUxn1BDZx2SCeZnbsUuTYb72Gqwf9C46Bvke50uUds4Yf8pQR
fSmzJVljd0A+XEw1OHVGn5PUDZcA4Tn2hsJjlSLVQooYysOzt9AgJJ7lZfXmkMp/lDCkF2b48ZKC
2LGoxhFtmESROa2rJHuWaLDOOB7cvGrLtnr4MQbifyDHcwQNGxVt/9MHoAAiheq3SVcE+SVFb1W2
deZ7uqVmJ7bbiNh4QmdhWH6CqStMmU9fUvidIUn3lPxVj4gjPZtDJJUVQn0MbJzyJplCvtipGLPZ
FsmWEAWmkcOINNX4XOc2BZNhZnqkD8y1UcMsQ+h6gGYll0+geI6ZYcUla6x7gKhybmDSFUS7cU1A
morXp1QRYocOsG9T9UpKu9TGT3GiWd7biwDciNNacOCYua/XK9i2gqbmPW6v0qH4jAg50w3KpqSI
EkzZysYVUXbUtRAN0q3vQI/f+G3xVJrvaTeEJD0vf2REDQEGTUscaZzV5E4JwcJJLQXlEmrW+ADp
7SnHgoxeJfAlgS6LR0dYWuGIlTeBzSZJuU7ofurxciEgzrFt4wvwpr4LHFtc0yTOigCzFMKJ9Rv0
Y8DujStJG4F0iZaSB4wqBuE7B8dh7dWINwdYFRvtqDRmCTKQev7ocrCW+nS/JtRjaMfMjFQYPR0M
Sze0En+Wq9DJJwt9eUd4abvyBoJRNdvIbCpTAUnwqJCUQs6cPivDLgDjYCZu/PWy5UNsxwdE4Uqk
mFxS3UjEGeCo+bfZz4mLx37d/3ii25yU5wM+AXQ0XIUlQzdLO7Cae1gXu0AQKiN3rMUaK2lvhw9k
wVFGeULHm/oojQ4wwsqrRrmWmcTrzpEDBjhRtzKQoXigQQDEWyGFuy85gjPwPpO5J+uUgYc6mmbx
VfUaWC+MXlsx2DB5fvhZ1nCn1GWVE7iyNOaJ4g/SNWwpqiVbDLL2Ml5DwDZrY9CV5NEawXI7Zhse
Ed1/dUYv6pQHiFdfPBAkk+ZcyKuze9Tw6nY/gV7FbdFBDwta/+WOW3RQezMPB/4f/eXAYiTLEFLj
2L9HYsAJ7B22bxtYrAtIqOQvJ6OOX9lnevh2WZyHW8r6m6va6AIrqL9LRzShdZHnUMo259z3tbQ/
3GOFwTifBd0R+cVFWJBO20UCe1qUapD2sxDjYZdm+y9gqjJ5ZX2ywe+wgPDJPSuEgVLC/pseubN/
VTBfKk6hfM959p6KNV8EZ7MdTOwwUjFPRFmQI5UjFZorGy+/ELdc55Dx2DPJMCcHzTjsa6+68/ua
WcVi5ScNxMMCWmiYLrqLx8Hbl+RJh35HZdpx202dZF81C7uaMGsMLFGCjy+MeuezU/qnlMAEYqpH
wqVsvuZ8xkPmDQIS6wZ6FwZmlLdL6X/YnmK4e0MvZDu0CqGI5a6e2UlXplm1A1jNnh2OvIVZalwk
YWIBTcNQsd5LjNcHex/y8AjCJAjZUwL+4DoD88R4EK0DD3J88QEfJCJhSaIw04/FxneNH5l842zm
XopVUaiE5284niCX6lUr1j2SRICCjpy4gcHU53UMMooVUVMl8zX1bl5fwHDJ1L83zPJTj3eatPEK
0BbARxXnHMv4LWEjF00krfnV8j25Gq5jRPAzG2Bp0rrCiOU+WCnGzhLaGMaJyvaUPJzsKPljOSNV
8DFhRyw0OqEM1JmMiQk75ARO1Kx4yFBluUd8uyS4fFdSfcrRaN+Kc8d3Yp+HksgtChOwlW/yjjza
fEF/pQZO4pLDo/aQdSI8vYnwEBvg/tzsvGShoA2gUHzYRF1FfZszjknmLpQwpNEtmw2grXHV6hyR
SzVRINJ4BPazrNhy74q3Fev94R/9UG7Ktc2gB3VDSyPw8UDQy+CbS7/knCjpA3IcEZNE6myIZ3z+
TbeN0Dzafl3iScIpEeAExu5vjU14WaWgU6w4lRm809W6Znwm9CV8N8GHGAijNnPj6oYkagijxRa6
ejmo+9lWE/ty5nSdYT+2JF/LI2H06wpnsylTQSTTPbktpbWE3/uMkt5xX4sv59e3l/c5QtQQeWdV
/bRJTNirL6vVfX0ygcI42fm5VGzipgEOR4q5wGMGM7zLN6Sez1ZrJqXWKXyJpRK1MayxoFNfj8gy
oWS5saQag2B/Gmuzu31ZqfZ1YSunmHgTmrtxBrdKNS0/P/HSR0/SwGhgm08W4ZC1l3/giskN9kks
FqxWu76I7ebyb6vktE2WC++IL4s1tyw10HD2wfWDC27AUjqnVDJi0GhTOaw7vXB9NfBDKeugcwbS
Y2hKgl6vkMbt7AO/WcXWIQIOKuUfc/swES1bS7D8Ezm4CGgipsOYTS2K88Yj7RZan83P9NMHRXXP
Zq+4dwtyVCOI/EJOlViquPaNJI3gO9czuPscemuX2yLXQV/thw2WFu2UZMPin1cr6ns/WZmvALNh
cYPXNQiAp0CVk1WzISAVmXYFLKMVDQG/bBXNEeYCsQyKdlUaEqMgpmfg98saHWIdL7lc6CXRbhBa
w/hH91oGYxsfEICN7KLnYyyMHshRDw/Ufg1GuyVHucIMux8cSzE49DL7AUbWR29p4R5Cz8f7CY8a
fmta/HAe+aROrxUPO6EeuMV3Moqu5Z+UDP4N7SrPo7HTzKY/UF+qNFA2Z4Q9TlVE44x3GnHKwrFc
2GHKCu7gBi9HAPBZgI1ECa92Q0PyuRzIhYIGoat+Q65Eqgbyi9etBlpnp/vfq0BUXw1XmPhzbl7n
egWnQD530YMI7Ua5AL87LROirV0Q3b///U1udnxjH/I3Ei0P2WdtqiC0DBGMLNG+nw94pPqkJ+hZ
qLxPgBjfuo3zUx4nDOtSb/N6hijVrK7a3OTT1Nn6DG6g4hMMNxKBNIT3d3rCVrXoqzqmMlJIVBYQ
TrL/pcqo73ESI9oSXwdYXX7gA9GatVl0lXBftP8uQTHDcaU5ZYgqGS4ET6+NsXxkasD3vJg/yT4Y
i5/OT1xwEDSdRUrElZiV+S/50Kq7Ht3c4RaQcUvTYhstFNO1f53IRdiFXDH8BKDbjO9TDob0tN62
KNBByUvQDGIWZzVQ9ib8yVjCRrC/SPY7zzxVRlgeyoUSKiYiWrqsG86l6HGPT/B+jF90NdAbGEox
Bz6OLqrSixzNbiYQbzIp+mYRDZ8GapsRJvpSJ/TmC3+sjTgIsMXPVKOEsrnOoh+/xWGcB/b4eXsB
uQoV4a943COwhYMWHeZ9Mjz4LzjpGov96XcTnbfCz/Tvm2jFmZvER0LubY/fJzJqEi9Y0fIgRvYT
CHsMUgq9pdi/lLdWsOneA0wPQWP+/ZhvFbgvuIiqXOEuobHALWJ054bx5oiBlyBVDZESn1xIfmXJ
YLKHtx/OjKT8jlz+YxXGZhksSNuKq5ctcEtILDaqoEwft17yqJtcp9dLW7BjlTdcyHw1H5k/ts3e
rFCGMgNQrG0RjeJANcs4hqUGEx2S8tdsMzEG2L3el9eAkyZj379xDJPfr6UBNp/LdHZaumL9nYA9
/7tFhZwU4OSrtdbutS/ONGTbPdf1wiTh370REaop3ryZhxcczVeupPvVnqA62iVXIlCFsuBp3kQ/
l2dGIw5JdURd52k5czGAXcduaDCcedxOHGINIOqvWLsvybLsycoduWu/ayrE0B+5geTzEG24pSBx
7KVoqVKzdsQ6k45Q4QQreX9sjnldgJwNGcuLmWKyvmE3yTZOHHUDS74WuQuby6grbryiK3YwQQ3U
8Kf2wSpTHoYr85q3qzvrPP6FxVGcpGUk+RyWV6JVD+6DtP+lzgs4wqGF7m6oM4UVNUo9s9POiTMv
h+hbsoSVZ4lq3oj3+CowIZjirdzCE3aJ7QInRvMKGKOZyk7PfTCEye5FVFU90TmO/DcsxtAnwCid
sMJDGsuvF/Rp+YM8OUfZMs7O/LfqdpadeGmY6chlvghXssaNAKa1IcPM1ozS5lWKsHFy0vUmQJlv
PngzoE1X1E2SxWWj0iMF6KlzEfCkRVdgfQQT0xcYxJswiAFGhegGeWRq4T3oBpnNlpjBeAhsUDEU
7+ibIBzMM/+2aJF2nDU/PSR4I6Q5F2ElLGJ9PWww3HnFSUGnDYOuZMR7/lrMwRAnevLyEHRumALM
CUqZTWboOkFZVylEhAk1iSlURxbOqDEfx1wxa2QmX+l0rEX9oglRfCdFh+2T3W2jIx7wtyrXQ+Y+
bdoFKsY/97BmNO4YKwM7JoAWNEcEJeK6yCPpyA1SwwwAU3oyckxtSWe7QQx6J+/zNXVJ1eIX3vcG
cNu5BOQrReO77vaJ3VC6NEqQfcwCvXOIpVOlLVASnu6XMCQQpVNpKl4Bb0EwtwjjSU3dg2vKsmo0
AMorUlkGYQyLAUEavaf5SLQBhJ3AoFE/G6iI+HPJ4Q3QObNd7TRSaYc7uOWoBePUJ5RBuhceCUa1
pHQc97y/9EyoEUnjJ/qRu14HjsxOU1mNaSrARGS2z4Bi836QQsW3oVfuSUP51Ydigg/xJHNHNUqu
NOMgSI8r80atQtx01zbqv0TA3aweKVHX1qlBzTmme+9OjX9IbYzmKGcaj69uKQCw4O8CPha7pUnY
AFYZbbCIVSY9DAhpEaxNHEhhk9rSTnYZAXjHtKSjQSJcitT53xFv6oozpJ+2DL12O2xDz0Cu5h/H
rw4FFwWOw+V/Cbsb7N+mTqkBJ3B34wfmqeNiJAcd0MArR/ePTOefpPlRY9afoNawPdA1e+jYWDNv
TgFQ60YeCR2S38xsm8T51BUVAKOjlOE5y9+PtzddwuJ2BK7J0yWiJDZyFyVWkZb67PozmFXXQulw
1zB2WTGQMUqZSPNniw5Fwt9WjT8gBVkwA+5hpC+jfYpV/kiJ6N56Amop1ZLg7Od1AVU6Ce8DGPED
VPuLj8mIEV3+5eKonPbi1Z3wLTRg/Qc0FV7nTWX5i5bJcWmOXCEYmbWicjeRsKgDndB6NsVtISzX
vkeDd72jIvQiJKzsZOdiJMNXpWyv7hTM6JAmiOQMumFQVSWscId9nJXv+IyFOjOis4ASnv2cCNUP
pt6voBrCbjHrSfYhxAI5yt5FzdzX07gweUm5jJYz2bln4I5ZayZQ/VyfSuKiSneOTZnwACY9n4tJ
i+fZkUcPT2GvdH0vcUioyHgXmJpaOaPix9AHi7HWxEQFNrSZzWJLH6SQRS+ZSs5Xs7vKuFVxOBik
DG8GsIRwc+f6Ua/qfASVMW76gcxrwbNsIjoBioSgJn/NhC12ygY2QjWPPpfuJvfShgTLoFS9jPOd
Kp6YhRgu4JSMYPiJN1NwoaW22aHVZQa9cTR3ASkD8sY4k8kofoqwjIrwjzUayAs9bX+5jlzLUj/6
Ez0eoN//61b+k/d8ofMTBrw1Ppnanxbf61UmuUr+VVRlTdtOWsoYkNn85GnS+/ZEH8sB05DDEjLT
5AgHKRsj3WEpdyhr+Nor64ZAdn1ZWzR4UqtQNKM14yoG/2MfF/u4BS0xcRTMISwGd8ymGHVZWqw6
kDiQX0b4/+vGy8ynWqW4Ua9splOF7Go89ZIvjKIRHTvveZOkuPwXJdhQNUvNJ1zukZ005jcEMSLA
xasyhCUOZpiKak8QS7OANud2lZYFw11mRDAnJNFrEUZqipqmOKWktaydga67lgARvo0Yoc8vWPgr
TXkgVhhqjT7ss4I3j11pHoQ+4NtD75DsO8dl4ZBiEg4eAKzccCFOm6EtYpk7YLTTcGksnTld2Dr2
ij1Bp1W3gzwqQAOBaub8xgmORYgi3YtsCpuTS8mG4HHZyMw9o1MSYP4+YWwTVpeBnI9Zx/WPYN3I
xChK+Mdx3xDtUi3bVeCt6cnt2stgS3Ys3IhlLZ0sbVhDXKN1ZSG4UWck5WhvZPpIsSe63iboqjVi
ZWTCn32fgmdcpfGCGENqTSnfOkqVG4HkPYMjD21FwFbeEw2K6j0rUstp9YQlf3NYeZTVG949uTK0
nhktlvPjmVYlWJ+UfoChQBcZebV4VEK4QTQtC8WJuVN7fdhEpTgmalQfoABzK2+oFMdUNU0PFLJ4
WVA3C3YTnLuIUji4F7w9ytN1vXhHFzRfEMgykyL8r5CAHQPZ2o0HKGZBCUkGYRKN+DsPhRoVpc/5
TbW83U0iWYHf//56IAtoxlJrApGMthKXHc0L812l1Lp+wiz1fG1TG7At9CNMNai5lKUDkEzcmFoA
OYlLslZ89JWg/UG/OrScQZ3sFI4Wk8Z4njX1eHwoBQUL6oEg77tXEjYyPHSIMx/KRGfjBFu1AZ9Y
uPDj3XYWl/SzGHEOMkDWE+42T5pt331HpHv2/vKygDj1fiKdjtXjRs7fGYYL1f6OeTuQHP7ms/0w
cpVc60ZMuZmvRJ5lEPKevNkSmKCXFH6Bt+lPwgCz7InPabL0w9l3uxwcRrWXv4TyJZoFbBzX7TBu
CcbRrO+fWbBkZptWl+A3Z3DpYZydLdt4s+9TjMe5O6C0Baght/pfDFUAxligyQlxshxxzjDrAJSw
YgKUTTFVg/eu9jWr6tIi6jeGC5T5dvfDX9Avh4WVTxXOYSmm5WehNQ8byGPH6XqO0QUCw3xnymtz
/NgG22mOXwqRcrtDOC/00Vcz3vLNv+WxlwT7e9WUsYoPiwRU3Y3oJrn4ffGkuqOX7x02c9CHZuxk
bLLdi8aXCjVR6xw0axClDpH/eG+zA4aQjbyaGEaUWMRCYUj8CRTx/kYpNPxY4QkMZdBvm1Y/pQLI
u0tnKQk4/BfbGpYpEBYDsU+Mzkc9Q1k6Vin+j6WhyXONpVRHCiC0lfpozFEX9oRt83eABw/slnAW
BO++jYff58vNeNueCUbYjqjTAj8ZuOaeQoF0SgzNyHsh5lJrc/NpDfmkFXb8o1ISreXiw99MJPBD
MihfD4a/vjaVN9BXbK/4jVtjbyuT9g1ELGF+HQ8ZINPReEDY71lFMq7sOHFl/MdI+f+Bx6h4vrpW
HxORylTqygLjasS4gLApwf7ROhoiV5tZLbgiPl86Sf6CBskpFzOiNwfMyXIuWMj9LWTdr6ZKHhNH
lFSqWRf+layjArskiXzN7sz0THPh6hgPcfXy1Bo1Ym8g+mz7ICBCS0yXNujeO6/tn77YExjG8TuS
Lpp5lVddckZasc8yLkJ/5L9m8Zrq058l3W/36i+GLuoDL40JDWDXpKFhSjOxk+yyhkKX0lnL6U9e
kMe4Cgh51TG5GnJpSbKJ6x4Y+JKNnRh2hdHmGSkY1yGOjOwPXx3dQBImaUE44pafjhEbon25lCRJ
nkP+NfYj/IGrDH/1sQ8ii+p319G9HV3dIzg5jomVagcjrk89X/X/inCeY8WCieWRurLN4ODm15h6
dl6IK61n97WHOoUhDJiq5wfCPg4p84GvX9KhuXGy4uODfUBj4Epje+PkvtAkJHr9JiLiEiKmB7Yo
gMZ4mjF50SWLzw+R7yZpEdtz3vtws+RfqFEt18OsGeJbt6GxJy2COdeSyH0aRJ9Fh8WaCf6GDcVJ
rxGKDlMANnq83AU40XBY7jURWfG6t/I9qcuUGo5UtUSM1O4TeM1GQY9nNlK0GQHiIlusxs7HscxZ
MhzwCQPgtj374VRQ2Aa21eQJXFEaUCAEcf5mg8fekCudqWH8nWHN6f28QRxcHRroPVCpgX0Lx0tU
v/K2H9apTyYlvs3iMDzCdohWHrpNVFLpdHfG/D66cWXAMKPAwZdEAys9wBw1fk2gLm20JhU678ow
48D3MAYJ7hxboXOFLxOYPYNQ/GQLYIwHQwvCIIsyp9eg9ZT+n22EtaY0YQjdbEKyXgXBU/ttOW1w
6+jqoGph+Rpcgk7PKs3lYkcr7ZT27vTIDLg8SiJHsP5Gty4lr4RipqfLZIEIVr5/EpiLZnWI9LSr
zldMmWcLcwyW/YJOENctMiA3+QVf2v5r+hLwovZNcRsMBPkSubiP5JiZX5gYHhoDHhzK46uUjDR4
DB4aIxNTR8hILIB36S+MTxyBF0Cc6pQuK9uvo8bXIjc3c1p4tuUgneDojdSqJuMV+AeN5EM+iGXQ
6dG5c4l2sW5TOUOrDbIBOupERS1tvwUJBJE4WEN+r5B/lK/CmpfS8p51xhvw0G/JAHJ0jb01nOui
eP687vjdMtK0vniXa80Z/TNKs1DST/5jbqz/vKoEopfSd0vq+RYz1a70QmWTRSIFO+Bx6Sp9qmn1
RRVy1Kksh+u223ORVEPXNzCza5eAzV48IqmazokMw3vTp7gcw2kgvgQrJPGfv6qiL68kRyloa+ZD
USUaaU+cfmur6tnNDwNt8qp5Nc6kBXSBTOSVLrd/M1p5stmw68prCpsRDcUPP9xdDIxQsXyhagVq
UBEGo8xsNOJXJKf3Vwcg25qRqfQdq/meNA3b3sP443p/G/fqdjHlT/sbPpr8SqubDQ/fJKOAiPWg
AnFUObeCKBWWdupZw7sGqy6db4drizSJlKFIhduw2iWqPQvZpHutaw0jB5zgkzETD9ireiIlVKXs
/aX+XnjacvnS1ZGFP1DMNZXafxoV3vFZrGm4CvBUoTRgKOhohvdM5e/mZEUAjjhZFltjG0XFTWEB
i/wdyYK0bh+tfGE+VZQnl3gpxmV5fviifGFPX/J/8lgxMoyQxeD8BZwdbrfwbGqOdZpte31d0Xe9
xalkLvk9jQy3B6uE55B1fWikCgz+jy8EZAmJBuvL8K8HJY3I0rlffaGQjrPpcnfNS86OGfUj7oEz
SQz2dGrR9BISrfGvrbwUtYaJHUJED343/MC59ZEisYRPFhvTRuw8sOhAUyfdJtznbsJR+aOUQA9a
SRlZC/7bVx4gdbUrCfKgyhap4l5C0+vndbHMAkfOVAa9RdklU5Ft2ISrRVjJGu7F9M1b5OcSc2Py
1lRSfbCsqMbOzfXDFBbsOADNQGHrMmK6Ic32uBq259oSC8MD8KA3s8zt6hK1qGL4xavsQtPmo7sE
F2BgoIJqIT008bCYAlt1XUI2VOUoEkmOCPCY/QdTiAvRJ7NFjp88tJQxdaGOZPyqQUN8WisaWhtr
3NESyrxN0p8P4JRXSlfrm7zZEivkiLI6zXLnBl/gv3yG9BCr54lV0H5OEIYJlJgvZ088zPZDweRA
jHxBIstOtnZHTCRi511yS1VyI0vDu6fDqO68BdSo7LC7JOsZmDMr7AoTrpxV4tl9l7mGt4gskskQ
yLklmynoT9fHVLS18FD0u2qsvzBNVfyCV2+rnrBeV7R4efzhNut9WhmYop40E95qnsRy/gfc7sl7
TctgDTSJfPgOx/MR3gaiOsoz+hoMOXppkC/7xPDKHc3bWIRAoVtFrzb8vaTtiKlHllmH4yU9EA5X
ArlGB1OWAz0095C+jhFIt3Vi0Q/sjOpsAD6yH5ay58b35MiKSDHQw6RYonBAuGtZaJQq4RUY3az3
minzTFzrv+yknhYjihk33AYSkLaCvHVfs3s53YiTF3qOhye5ORaXiLWuODul5UjhjeYVw2pBZIiE
a81yYb4gJRn8h4UC0JzCBK9ky/OKq6GNuDyifwrhQRTY/ViP8Qpv3bhVIJzW8vTHZGnv3OuGyMMT
JXa0vb64HGLVfV4HHHH7L6elqk6cB71MZMuPvFVxlgGcIY2MYp6zz1L8I0Oe0nmtWR+O/EWEZNOB
039ajf34OGFh4G13EFo/uczjz8lrlQcqJZCmpefbboUzwoBTKNu3xI/s8VOsV0Ew6O+jSVCNu4RS
OkuaVQreqpI5uEVxaxpubK9dIEiOBwYkegHj4lh3+tzhBgOIrQo3Rqkodo/FVHTUt7oSZ2mxyoXg
uu6kQ5Q/GbG6fVu/5VSZeQWvIGjJmfNS/hf7Q6hVED4t3mwd2SJGQrJ6Hl8fnMkKJny2rhjpNC8X
3aLKNzIikrPLSDSve4E4QBlpP5hvuvCekbHfRFkX4HJGPEk3FqlkMCmVa4IEVz0JLQMi+5osfBWr
ZEi5YJO1xi/hxDCJplffpMXBvFiG5LB8+aUb69xEU5STAfId5ZBQzdk3eNiytIyZVdYKJh/UB/TW
s53EHl2p3LBnhSS8H1gpbT+FfvLZDd6MJxiHadvg6ud72NsCz5pFCunjONmSllmqAn6KZCCTzlnL
Bkq92HitP+PD4rAaPo6tacdE7H+3ZXfYP+pnhvt6zOpiY02oUDuXGpHwk1OcLPFRk6lXE0SvUWUT
+wHnv2cC+CmkOLGR15X93/z30ku9D1kKqEg66tQqHOLlM9mfGqr5wZMAv3Ke2uqKGA3RHmciPjIT
idKRhDZErMBtNyZg8ppcXxd3A56QlOzQ0KlLXShKC2Lqt1R8ViHPOw64y5Vu8mQgYISrxJiLpRb/
1W56i56eigQMDxutdZzaZJCgcYw68yW6XnRZ5RA6c2nf5fxi56EK97v8XXWxdIzDNvstrAThWyWq
kRcPHmLjikdNFRYlE2yZ3qjEkyI4lG18/rggcR6LUu1Kp6eWIzKmxcyTS6WLCwXMGDjdFu7P+za/
6+cAcjLvda0Nk0mcarKsP72W+lZWNJiUod5x0JwrCwyNRioQUi4nMwZwCMPOimqFhp6bwqAEZ2xV
yTEygRMKDWCMjoEw8LPxbjkn1QchnERqmSCe2y+MWAMz+1RFZ3MEDKG9WiO+XSb9kGvsoQnOol4c
PJzAyNGtahWz0sWE1R/LEnCikOMToptiiZQO7ysQK5FsY/SZmUx8wo7iSyKSYXgz4OvMF0YtX1E0
ndwLi16/diflIIUl6z5StR31p0ikxyHLzX1C5kuxMHgIu5TXWwq+T1AHiMh84xlxdPvl+1678GYC
0Mp9/ZYAN0KDCd3PoChXcl8/HPoyWmmR6oeBAzjRmR930MTLC4gu1iu8t0qk6v4gGWNQKWhjhsau
qXIIJOHsVthrFMBwshRtGz5nTVk3b1wOwE1fpgiG/W7UX/ZkkJkYGjdHGHW3oFSrfJkQFln7AYeY
NXFu+57xZcAyxdkCFkxMUq5Jbt87nWJmPglEitII6nhUgRH24CYi1yJ+G9uQlu5GnHa6pIqPdDpK
LibDB28O5HKDQn68s5/cvkQdoQqqaQcGcPo/cGSPLi38b//wGgmtFy6KQb+PdzUa6EyQYtdSRtYV
LLpt9Hb1QYnZ+Iy5x0asgXjKT1F/+FE/gBLbJOTsC9pX387UZMjHlQ8P884XlF34nvNjkwUHTtzF
6zbztdwfB8QtzLE7Y8UMKr6ESIGX7DqInsqwNlung9IcBMGxyWsIADgDmgkY1f4gYLIvfbdCjCT7
Ixyg+Q/PtGuEKTnJ2D1D+hWMTWjEH2tdm+GAuz7KHwvIxH75FgzC/wYB8r1JM7maorvXflm0N5kh
7gCQ7kKC6wm87XoMAVuJmYQGCjo+yhzUDeSsEvzdJrqU9EHi0SJuc/Pw0jH1qJAnwZuUhjlqLadn
vW7JFsPXtkz982WSwn/Wn017AhVHbZjvUd9OFtJT4zqDgp1T+2ZUcpPpTKrf6wznEk3wuBPHXn0k
VGJrmse5aZ4gLU6vyCiPgnUxhp4UphhZ2vhe0wYSgBds2U/fBh/Vz/J1SkaInAZzqjl9hJG1TWFx
7sucXKCO9IHsdp2zUut7CPwfDPVfa3xXruAh0uMLaCNO1uDDf5TsxGjdJm/qem/kZO2BTa7of15A
bASpamlOMDh+DWW0xvZ5sOFCq2GJlZpCe/4PRusgPlGsiVJ3wydSatDOlKo8sMNNWG75a8CNZagM
SgKE18hVQUgifANxFDior0+UBqrxSb11R9Csv0jSOI0z0Auo8NR3Sa2ZEJXWNx5acxrKy+YN72IX
Ez+9u1V2IwUrrjA5EQps/PujUf1TBX/XjFKlkYLw6HQIO/FxiCoP67R9ollrfvhE6R0IrtgIa6y5
3vJApPRFf7+ffQqswu2opci+OLb0/BbhRAS14sM7ev/cE0bdEoTY3NCh8A7eUcwiyvw7PyTUWvns
+2++2UjJw1v8laZgQrMoj1KFlVFDkrH6VNMcxZExsEn/8TIjG0kPJkGmo3hv6LadLd6iQxF8Oa+2
4gBErWyGndG+I4BWFQf6TqGI82v1fE2lC/gfjj1Dxk5zxAvYS5AYdZgp7nmkAVa/tq6kp+Guokkc
LCl6AM17E3w9WmV59I9Z0IH/okhdFqq6awkF71sndia1eCB5ANHWrEWglthiLcxxCT3QG5uIxC/W
0XvkNTEiEqRbzAwyoW+XTNY0cWTUDuKIc0/0pBnxKxC92F90HNh8B033QpDNP/wJkr6N9cTOnN13
3lELprILkaj+WDlrJRMHiFD19YbvrcG2zQ0G9MPDuht88Qajbs1ues6zL/Eo4tHs/9Km2BfAOJWV
y6CiF+DurSEKYljn8l8YeHd8nXmQTUBw+RnG1mW3+d/SN7Rde2kHXjuYPRCli1Dlb+MvuBTZ63qY
odaNEV9MaTGYcaNTsbV+5ULRen5lE4thUbIK0I3xA6fL6l8GstZKcwP9F6Ash8LYyW4x916EreQv
cMyd/bU4n6lE4z6ExeM52LpRufa38OyoYS5Oep/tAzDnlfot11YQGlUxVmWFKMDDnxrbidpWPSjn
3RbEeeVRBCoZjyTzSaWY5vjLlRpwL9N/3ZjORVcb40+nOaRSqE1ybaELJMTy8KWQ2DEmZ7g8Ccu+
upqi1+UXVkm7HGAj3ONF9BWtbqQZkiAFjKKUk/B5znIbeX9ZovirUdBO2cXrnbY5+Glh1LDHx1VU
3KzOZLqm9VQw4VdkHQbALk/7KDtt/l40bq/djsHSD2Gib0fLrrpK18iLuVCXmVAT8ZNtwbi5bDfS
9+bLSCHhrnuZvDbNXO/P53fJXXiWymDKmwlTvly4TKE+F8GOE2urpeENGIvMVGv/JfF+idQsonmt
dCmlcEsvnhp4AKkLDNUAHP5skcujpg/GHgu2pSs8DMH1L6P70Dp12f4fZWZQthepiL7otbfKVTAY
gr7sEShvX9gdfJO/Mx9hALLp8B2z4E49o//YWu4wccwCzxVTswH5W4xNMvChqhehbkT8T1X8WrgB
pqu5g+pRdC+ZPB1lAoNaCNxC2o4zgy63ych5QdnwJxnnViequqH/C22uJBLrohYs6nLOYSKw22zS
xiRmb6l+Uto6SPebpgpd7gGONLLDAvJHZNpI4eB5svJRuM3GU4iPd5BSOA3TJjXE1ZMflGsCH3I2
JKHv9XQ3yvvTQFGKlxLfzwp+4oEYl46iEUGuQHfTrYMdUsh2f+PTifLIEQMj6ewBD3/GIQ1BLKAK
qta6DcOoYsxMewLBDo5eOV8MSZ/Mf8UiC3McGCoOVqTtZwajAF1p3hHOKu1ExnoY7aLXTCrt+9mz
9MAH1d9+NRRdnx6EkcBR1kJojotBxAqbGbNLgya9ZyfvHT64oAqds68wrOxGpjf1R2s1GB2TAEup
HBQE8d2E99GYQX/jEQq4nRxEbV0HC9QYzXMC7RnmyBKqQHLEKcmkYNNhC+p5fWCm8M43mevmQ3h5
Y5YSBq+9piCNtT215LEFoqtBGLNaP7LPyIwaJQ4uprA8lqJejLK2PyNmrlbtvo6+DCeJnbREUwqg
McvmwgVpRqQ5TagSn1wkDGselphrzH3dAnVzbGU6UsYTzNQ8syExK2YHkH/lE7Mq/9b3/0FsYXKy
1kk3ncskRwyc3bHiU6CDeLNFNGZU2BwbwqKK1MfnAOCCBHZaHc4hx49ZpQlmXVCQojQZo8QeFbbs
CyHPlJrPSCz/SFHRXqd/CiLKfIdIbY0Lr0OYR+yVCb2QEPnmYlLcSBcJkqYiAIW822llYAmbX7ra
JTESAAuNIEXwsf9hZlH7+rgdQ4IkbOn9HoAKjEuwtUUc8QDjj9temmndFW43W0nBHv/1UPMcw/LK
1l2fyrO59UtiOsRyiviz9LF/Eyln7X3UbuEF78eeow+ydKkrqo/rojbbEKoTiraBa68D76gcAtVh
ATVuVnKbF1o7eE3eRi96xdTZP7+J1sXt8FRH2vWdigVCq0cTeydiOnWDzO0+2YwyTYNuPJwON4Qm
a7Yg/LJvkeu7Ll4FW2UUUOHdiqJQXnNXv87kzvkZP6DWcmR1jqfyo9OzwPsdQKpu5VVGn2kXWJfW
+u9SK8jGPuHN78Y2DPhtxL49WdawcmbsKpr3Dr2OukguIQaN+/n5q4kmEXkGLUGqOp5mDCtyHLPE
rszOgX0KNLqfhsv4FzIe/3kEnk8b1XK7UQGgrXlugrLWDUuILyB+li9Sw6wvjY17z3TUnYEa25cB
pVzp4d/mDdfFpVA9UJrpnZw0kNbnCPO8wTDNNlvq8I4cDmlv0Mx1jE/ilgZNmFlaoE6IwxNeruHl
AtWsZID7oG30HT6yUPfD7PSayb8dyrmoRBtm/8saP3zAsRzARosDJAVJKiBzVbcntzQsfrk7ZtiT
yM4NKHjGnBLuqEkn+/QSSG+D03hIeQxFqyPAy7UO/i0zbjb3UZTldDB8TwtypR+ZjeOHW52vwGId
1t/BnTZnCKTAaUEHYKIfFFBNmcIEEYmp5FDVpB307Uq9gZTE3eEoSGmWMBg/q11YooeP1hRM6zkg
u7VW5TvIPpnJSyo9mUjdYP4cZg+3BdQwy7waBk7ncMOe6XUA4k0ExyR8guQu6ZUJQtwEw7bEbdKl
HSm5Dy2xL6IG/++JE7b4cTOXZH3IVRlpZuCz/DaHielf/lYKHLmXAeackJD+dij4DvTWl9yT28hD
GchFsulEYwD+mhuUaCvqW/92elZW6GDimAo4r2L13EIFp7XrKPy7s6BSpqt42FpLU1eb9MPin9w5
mZmG/RWNSKxqPNSRbOTrssSO+JeXmRicJXjmCeW+0iHE49/qGhaHEY1ecP7NxLwT2uFN5TZKCdFv
9tzBHxwZZSoIqVqpN3jCPUFdkcEtxFoM7w5+jjd9qSsIbqnQcQ+8IUeSfrOEoBA9to6TD+PvNZRB
IBAiPizKGDwQbft/iZ0mTC01qMzfwI+rxNzGoQgBnP9LNVKYu0JUfmAJS4prQr+MRh2aZ7vnvs4p
Jeaoehtlq1aM2K1TXxPDi6JXd7QO0iAn1C6KMsWUpdXejKTGex+75/iKuyOaJJdWQP3j2fOMxqz/
Qd5JZ0ub6wJbirvmWbpKVkcArgoMC71b1RvbxlrjAB9/QZdxoXiCPcAmcodg/plx/SxFj9XjorBE
1u1zr6Jdioyi8CQIQ/x+6sgN1LkoUWYCMHA+Qc0lUFJbUKGnc6lPd77ZAmiSXUw30k+KkdxQ368F
DjsgwHpBR9U0aWNQYy6fmKTwhfaOCQTQjiS9ImRBFTBAGLWmxKj7FVYtPkWxLUhKB+6jUhyiFy/l
y0slIwosrU0h0arZv4aRxF125xfMOHM3517cQdghMZCozcf6dwn54LjJlD1Mx2Zex7FHKU1cE2DU
MvqDVr6Ec5XOO/9KEewTQlENv+fpKenC9ZNqiqrCTL09dK0ctUBofhkGpY7rB2MkwQOaEnqdhvq/
638bKRdYnBPuWbpzvg5zTgZLCuS76Na7DHQsItG5HJlSE4WAouA4D9lszjbSlcNMhN96JFq2HYj1
qD3smlBDaq8AsKcOQSHQtsMB95uSCIGUfv+PE4UZVBoaS2fwCZhGonPEXX4KtiMj6tWbf0a8dTC+
iImu0lpZLNIu9Rjx58cIj1/DELVwdXjmqivo/JQHiX7bzz48fkxbE2+vLWPz7oai3eSYtQdQU2S6
tNtQ6/GrBRaaytYaWZJcooXrEl/SBKjgagTibuWm/Pk/Hk9lVMVbELtg1zEDB71Tyk/OE5KuBvyy
ub97o1+EGQSQcxbU0gAj5R7cKzcNzrIZPcL6KoXdjy9VdX07rtwSZjesHjVqiZm9qe1UvieQ/ru+
gaVAxLvLcAcGvbhNshmI1lluPeI/8q+PX/rbE4ptEJN1q2YkxqFuRbVDAXd6l04qDe59kI+omifP
gWCbsbc7PKrGCE6YtwIzKqwK89wy4YTFONN9cBq88I7DkJ4PoA/vhOUabuVYXI8nWt6RwLMPkQnd
t/B/PpwOyoiQ/CllQwy79W7xCDUrHOZiuU8zQNn8HMa5zw1MzTG2cEJmbnayHkpSDFbgDQs6YD9y
HXve/R97DRckYO48bR9vBLGw/cf+dD/gWWflneVA39qJLA4QuC/IrzQn5C2LQiyB7E8asSbSPiJk
yQF9nN2RmQMxvgoyD4AXN/8lF5KYywCq8pTXzZe7H7yMIzBtE+P9gJK5JNvm4jTzuhFM6qyjNdk6
jJ2riNoL7Eup+fiC6u5sASEeSIs23Fkdlef7MmVCBkZeFbx5f+wVHNNUXqt/bx7M3FrIOPo/iD8q
gFHsF6TevD1a6Bg9fsOeCcLi5HkEhJOsAiSVnhs9R7kvT07AoTH2B7rsMdS0bNQUeq0tvvpwiKeC
MuVb2Q1VFJtVsRU3gkCVCNeC0DDgrFpspn7A+UTLpBnLrUnvOe9To6SEMoJoDMxbwRVfpyBN6NxJ
xlvZRkcX1nhoQuurh7y0n7Me8XYAUh3Md+lgYQIC3AFI23IXOvb93LJvhwIk6/B47CrUVm7cntoJ
T77nVRTiMbxc966mRTrlxFaFK7tds4eD+qY2zgFM5VftfYuRnzw/YRJQipNf5w6BE1jgwyORFVaj
gKOMT6E5NHsAFDS+v9mYis/eH0Kv0Tc167B8BEojG3g7Q5sWAqzt7AmpUDAUhww1Zds/IiBUfab3
MC5PWG1xglQ8pxNvEy4PyrBVG8u6/Fte07uqmBpITpwIOy+Jqz/DtA2TcgDKupEcoQACv0fLaEx1
uaEvZiBtbmxULntM+dDK+VCLgfOa1cL0Y0KCdKXs6b0SCNiXvWHZitgJrbJB23NcRa2ijeGc7J0z
doQxBxirCNga3O2SNxjuPj9iVmlePR2T61xPlb6Ix7nSAUPHuRb4JF78TE8X3Y161MLLmUY3Zlgp
tYAfzX/XhWkA2a7JppHvv+tkLCvjwcTrhknDCFakmO/08ktCmk7iVIDLzBJqv+hIuosqByJE386K
Ngt2Vz4JutmhXfujQYUTnx+zpvUXZ5Gzu3euY9RSYRw4k8d3/Pv4y51XsDsT2qzujZhSrlB5WAbO
OUa/WVhvGvuo6nuZ3HSmqYHiT5LdrxK/G8vmL0kjzEVk1XOpYJOPmTSLsj4zfofd41914jC8MO1Q
9hn3F8v+aLZe3a+Ir5w2oRu3zS6LopcQNqpOpJsbKJ+TjZ54WU1YkXUNgNrhQjQepMLVrBzIjRYM
63/sUBFyAy/NjxQCkP4eigU/Cd9/VfeEB4jQoeu7fdDqNET0jp869gILQUkhYbV/Ib8cVioBHKSo
DSppN2uJsY8gQnzypz2YTHi10g2LiKRVu6+QUze/fFVIr2SULsj3E46KGrNU7x06vq6fQNdXz6Q3
Nza8qR6BOLh28iqU1Rdy+4MtCIcpIqqpSRQ47V/Cd3CzKGe0J84d2lEl5RsI78b/N2UbUm4Xsq9A
+zPqeQPrroD5OMzhOIgUHu1j475fGZBpWkqGSHqki8MUZGIvpgqlfCB+o19EcJIcNmb9Ulok+5oo
t+bLEpF5aYwEx4BEg9TGfHupeIK4uoTE8eNm4oihUmbJnc43Gu4jGpveuq/GSgWOaMByJkc79EMQ
Z1qXHr6/KeNkDOBmRnb8lTTDl4U+9s9X8X3gw+AwTjdG6VDlqIHVAEOzCqLDSTo+yeghND53PYu1
aePA5Ra9ghq0+p1iUKMRDVzUMLhxV33csRCVP0c+3N5nnfBzOam6Ihhfi+YRBnG+G5CbI7yErGTA
qY9wE8xjbFGTneaxrLzlbslJyqWkqOsTioM+BYV4CiVHevXm9/fwJfklvpHzei8txcKXdhy949R0
Uz4GCe6LMkPfVMJhI1haf3UuTR2viI6eDMOv3zZtpeo/L7OfnRMX0RYqtBr0ovaJhqfmpTN2Ao14
WvES4c92kXTcXZp5ZfX7ap2TL4YyoZylWsnkXdA9/e84CGY0pRcmP0nRHuQ5txW2SUhoWq8hA232
22HunwZPMYhsKPQKKLvfzXzulE6yZC2q+fuWutVNo+55xtwak9jNZ6vwtPONqpP8dGh8j2ZGXeJ/
XcUzQXh1RDMeUG2mujFVkFmaTT+WF89xXIP4nTxfAOKM/TtK6lTkDY8HPZAi3uqZcFNRwIGUe6+t
Lpj6gOJhJWhwEwsjZyV+9NE5QfPKan2eLQHaxX4KYkYKNRkBBjO345u0wC2YU/pZxrSJ9x9USQ3N
KzsCyU/atejqpDyYz6dH3X5RHg/TcOgSug4fAZs0jlOcxKa4QJ3hmOhhuafCX3Ln5ZM4xMWaYJL8
UKYhPmUiyEGpFn6p5Tkdvaybw2JOmyR4c4dNACjlguUInXxuBUw6dJBbPgB+iEvX8D/u+ov50UQq
O+444RC5vNNSM+AtZ5d48aRn3V0QSqDmVUIUcmoXte6dLzsQ4XwrQNWeMK+3QP28sb5aVglHnzvf
dgOoPMPI/RCN8Gk1DKuW6k5hpADA2zWTxR51snzqBYUTofTu6Kpff5VrGPOBLo3XtWGge1+mZswl
V+9H9SSfjqPITEA+CEAqCVThUsvRJZCBBbiC/h10FgheVyAm3w9Gbe9qQVgqEXdNopzP4r0c7UYO
JiHLWNaFXE5wsajskPpIRPi4UT3aF5iWWLLiknynPBR9Qp/ch2Un+lCSmplAoICwEihfyinzSVjN
NEsLjjzfDVqa5AWzHbHOaTDL9caaXJmFMLTUkQCoP1PuMI9IxwYnDj5uKdi8A0pjGGCMh1FsOY5d
qBDfOBjX7PGmYr+YRE+0HyYEGBRg/SVmRzaIA2p/089h/HIYh5p76KVZSkZfFYkdH07L67sCcypK
8fxGIFC0DLC+jjcVRjd4kG9GVz+cQwoYHalxL2eTdQlUy+W8eSxeG7x7Y+WgIlQnlq0lzm8rPbJv
a67AOIJRfVMH9fyYhCinVst07umUH1oDFbueizqCs6hlhyBYRYYrlqpELBte0khelFQDPFa5lnNC
yPfsuK/iY+QknNHCxCdrnFeXxfTu9s8wfKKehYWv15Jdw0AtOF2dDujEaz+YQ2++/VmNkZdMBjgX
03nlgNR4Xk0yQh83qsNywKzhjSSKZ89rg65qAsdQpkEZZnzKpYVNfKGegO3n6dfTC733DaX5mDTP
WpD1jW3YPJg9E0gZ+kCb+ZYem2yBQrBlP55lV6Uy6THTx3XQs3ba20vOzuSM+263mSDJ7w6mQyKQ
0DtJ+fprGSHtD+qCkQvCTImM3o5n7O2fbFlca+5sJDGXYyIKpcqa5encyxxHSgDtUhOQnYrRhHnB
/iG98QDfpnPIRbZBwx02LOEBK3MbanDQjNOMmJkmy+meDwOrUWMRpdXtipmceEUyDdjwCGVYbG8K
ohpUecUODvTu+2f2MRX5HDOtd/u4BXvJ6HXtdfFfqHnebnTY3AD7jBK5tiUAibAeKjpaUeTWSDem
/6DaBpjKjbC+/SbTC+3R9d9KiyFnMauO6MjWytuI0Sr00W54nSvxTc8BOsnDOQQ828DiMU7cqkAU
xbTqbE0ObzdSxkw5bi+X80eCQgQDdYOQHyR2U2PDJ7xQHHmwnbOcEURgfckcTQnDL198gPBg7W3l
X20BDBxjXCwYd0kNu/uOACVjXD/PLKhIajj0teZqihQkXmNizznN4efsa1h91PDfbMBCz+zhqnza
roTPj3HEuGRgnt//52t23MDqYB9oRKxLPp7sgo1NgxOXbe0V4LvzcqwcbHQ3MKnl4pIQRsnKIcsW
76shGZv0ZAdIEs+jHMZvtYs3nUJErtGhu0E8N4S8lUT7IphMqNaFoDY/8+40+ihVz43hzlTslD+x
w3qiWsl4SSBXSnR8r0jnauOm1xnGqg3NUggsc3sMZJxeyAnTLJ/jkAdcAHNJuEgiy1B2w5r9VaQ6
HE0IlDUjPzmkVsb/TZtwgxULXtryvpuIRHw2ZT6gWOVR8PlM5nXmNpgOUqbYc8vh34PwzWf28lHO
jxFjYkYtLSoNi5ZVBBZU8Dh9ziOvKDvuDQeQmKVDq1wTIayZImYzY2hU6jlH2z/LyEwg5TiBF0Sq
KG39gWDfC8GN9L45VcvGV4pAoQ3ce35+XTQuhM5szHtKHuCUCozYT7IsNPPz9NfyrG4P2zyNsv78
pBgEcb5jqs10AWIA8wIXt1o1RigDG5emnWndrn9THJ5XzjlpL77d89fxj6PBsy+3IWbmMspbRejp
swY49JIGxHKBuf2I/dS0v0AHJUKRD9lCCaPFXLHorlARdyjk7RQ9/mmUH6oac62lZKcJIUqj1haj
VacAjOe7A2w+cEsJmHDJEaThs66Iei2ZJwSwXA6KcizxgwAaidVDsA9kf28zEH552r1jaR24rzXU
CgeG6i9tMmzDGph5sBBbUl4/t0puvDWQmD3KszkDP3gdvRfhwg7RPqnvT46TdGmoTIr4O8mMVlnf
7yxiQLwhXV3sw9LjFT51zUK+TDbPbsIL9hsNfcnbGNRCAb2EGrS9P/GX1JJvt+nZ4m8f3DDurFjQ
FrNd0WvB11Oli3QqAm5Ne6mWsCiSk4LFwFwW0XCe5+BOc4sgdvBnD9tSHS34AcTrVnFYlzCOgYGd
Rmi5zZU2+60baU/AG+3/Hlsgr93wA8GThCfNWe/XaGAN2HnNM6/NpjzZN+4OWmsy2inHetcyOJ15
yRR1Rc3fpFj/dO4i4lnsI2fU5d8EviLDmvP00oRRh3GOZ1TKsfkuIAa50U8YudfdX+iVeLcMA6qd
a27AV4SRoUyDFK2GyxYd/urwybRCbQaoTTVB9o8C8Ib0ui0FOj0AtRJJ9+1w1JaZJ0bknWB71Nqq
pIZCKXZWo5+fKnErWhMhR3exIi5v036wMAfrY5kkTP1hdbqwXnqPxWHZpB3vAKUFsPQ8UjX5Xr8F
pEmNyzeV5a2psKVOUvZ1gjHsLp7SnnwW2n6V8f/5rywlyWsg6ZajPHw78sph+HfHJTsUOqqpGU1W
RqhB0Mmq+ikjbsbRQY7wQ5zkggS84qlBkXASP5M1n8AP63F1fPhV5hJD1r+PcitZHM8pQJnTeipt
Qyv+H/vt+YpIKUC4jZvAqoXNknyxNPBQRkfutSUdfzfk6K8VM8TvIaFaIN5Y/ZX8gyytIq/AMA1K
sggxjbMA2mrkG+x++B7TwH4hC7SlnARNHWZEvwfKMwpZWZZPC01zqavXVymV0d6MoUlUVppL563n
Q7quge0oHpzHoPD5USsCT2qdCeo7oEHtYEo6EkGXGahaTbKtRQ3yxLLvfKUx6qgDj10MtED+FjoS
78AVSoFisYnYb9cDEoSlVw1pnLK+34KynsYz4k9BkMx+WYIskosoYVZUcu1ZvoAbbdhpa+XcbDe+
7CdjAARePfu0fXEXW3LBUEgyIsptSBu+yH9f2UJG/igTyouMI86rJ+L8K6AWbsniwFeEJ7vvqoAa
dr8d08nqIA8RtnTt1n3uNxYV/696PtSOxMveHVY4qitweHLJDgWznFNg+bh6xGsZKjCsbaQDET2A
8VRQPsoBx0v1wGxvAZXouQXBI9eoAVm2G0Kd/s7QmVHW4NzM3IhRSUpGqdOtbZyNGzqxrsB9+h2j
gZCwEbuN9TuJUhgp9A2iv8lIXH0VSsqhZqfuA+qjWxSFqvhFkCmsiEiQWY8f2lGOo6G0MlKWzMOC
nh3GYKaMHvPNjYzIYNabPPjDtMTpYnPCeVPU6rQYIFCLwU0ElKMmSU24x/RApegG85cZVnxrj1TZ
wSQ11FagyiAWee3MGMsWq4Mp2qldGyLXN5g/ds/q2OROu55AEosXmXw6L2BnHhEX8ciSn0QLZLH1
vE36PyrrYLBLJ4wsh7lF5aI1nOAgXWqGBFsQFM9n4dr27zOK5wUnW4HRML2B/Idri3Q+ofOJ8z5v
3GbEGpii7pd0Oy+tj4hqbE0K71xSUBwcfyz5kqbtAPqZstJdckJj3N1m7TX3R6uBG9eFR4uxodzY
yG3TViXVsH5qb/k2aI3qs5d0CbTh5Fw7LkqKDLjAcndEGq81601I53FlA9KW4MBdnPb4zEvivQo5
vqAaaiU7VrSthB/fmkM+K4DZbBhkKZnISKc5qgUN2EWpW/PsqmfBrCeNpZe5NOrm91p3qlGNJ1bS
F77m25SpFaygFpLi22qNJKct/dYlAS9KgJyzfbgdntVRYbEh0ZYtnoL6cVnl8aKAGjEy5F7U27ds
L6RgTWRkfXxQSvFQwOx6MmMNAmsvDz0BclShQlfecqHHMdKZxHoBmM9Ql/KzEwagSlElfg/v5T0N
UowRoAISB4A6W3JBu3Bw7HK5yD/gPTDciqGSrxQOiCOqNB+upNaocbm9Z60ZoYFXv2OkyVmJfY+G
YQLnDNSC3ULm9l7+kvzmGWsmKxvVSGCZwybOmYzdygZS6yt/7IUClbWoR5SP20+jYpUzfEWk
`protect end_protected
