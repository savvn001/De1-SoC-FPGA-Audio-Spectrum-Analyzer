-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e8sQgRQa8SHWI02+rDOUlZUr+BVM3ij0s0g18klPu1VwxINaiBeM1WhftHjYQzc76YNZ2nvoJ0XC
vZbzeBT4g6OWMNlTTQ43vmllIoB6prMMXRxagsjpflfvskGP/gy3MeFDQIsiuV0hFT9XyoWejmQR
iyZYIcVzSAVp1wcOVkKX/A2Rf4ZtFxiaQUg6NBZ7JkW9HcB6UcmI/IjAihfPyX7Eo24vH615uWcJ
pTzgg20VYuYgOBcHa/gfn+FUzm/JiXeQgyvG0sV2NZJsIDtOaHH7EuroMq5SvxQBoYQqqcUtnXcF
0Dyi6mCFNjU6R5hj8GxSAOniJboEPD+fnqNdsA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124960)
`protect data_block
XVpRCWTko0HVv1/NK+V1cfywv2Nmxu4EhFoMXCE5CnOQXtMUqb+9Xuy1Ged39tiGpyRY5PRGJR1y
qL5cjMLqH6XZ/DMm+UKQjPDQgqQywEXjv+rcIKaWbpNmqJaOKo4TKhcNPAw3VYCZ1KiDHQm2fMSh
1kYiDKAT8ZesfOhH/a2hlSZorvXJysYBQmXCnuu9aZtpsBY5Unyy1VPUFfk1tTdodBBgKm0iD+Jb
L2FI6ym8RKlAPjjzmReo7k+TCvYkh5WZmgQgUsRLbhoUDjrZq01r/12pFQdUxvPiDpE/LXs+BRvj
LT2OmWTsjGiwA/qM0EZ/s2yO9ymWk+HMAae0CJ+4RZNfZWwZnIJqfhxDT2vbrxh3u1S5h8YBJ3Rh
CAw4KfqigCgQahcMjI+/XYtktaKUBqrxbgTI6ljupCmtpLON3Agy7rK1brVkMiaOUcZj2tGCmZsy
c8PAgx7pyv084KCzxz978VAmZO2NwkDEBSo0DMQf2cYHqHkmsEAbEDRg9H7ISpTQ8BU4Zbpn/0pz
bFvW4Leqbm1uESJtOUaOy8EqpPqeDnGrcEoJUk6wSSzn1bsgX8IPdDRh+5pdZxGWAY/axe6w05oL
Fhwgbo9syfErlo4xzlRbIAM2X460l37KNXQSUr4ldTsMeCaL9/WfAhJlJZ/BZ2YYwzNYzLQRk23n
rMNxsk7Q8Wbr0bNZbGnJFJZG3d1yLyNiwsMOZrYuQEBK0yeL+qxMvpSg+lKhQTgICECU0WW3MT5U
/DmPqKzE8lPLNxe083P4r/4mFosR1bt/E6ApT7P3kAUMpK5lMJmSjrwJwAhtMPwSRwLQFLlqxjRt
ewIP1hN1d/Vt50E0HEQGM4MGSnJhHG0eUMfs+O7YpBuDk1SA2RhZoG4u5xGWMQPgSeLbNIyzZ1UB
MsPvFipBe26cXRNF+4yqNyg8GRdQE/LcD4SrHRzWchutl6wlX1pU6gPUbKLTWb1J6K01Ql20oeXj
Z6QxIF+8Lmi9aehqUtm5BSV2drZONzZ34hx4AOjjv1gMgkSFI4oc90iBdQAFXe5aI3WbgPlBdbMU
iQyB8bzQ0vmyC3hwau7JCwzq9/Bh7Ym61OfjPjJAaN0+7qYNboCsEBcZZU5/itcda7zy9bfUAc3G
bU9hPZmzvfYP0XSyjZwez/SxRXdOop5zVyLWdE/3XWJQ3bFUSl2A8G3fH8uyV/gHVjFWZLN75xi4
1uoEoqBQzUhblZrybJXWlSjFaG/Naeydwot58aQNaQWtGKs62a/rJ9KnClX9ZnBgWZPZDmY86S8P
QY3rmB+eFAntOnSfrnuUCgHZYKsTMAvb7hHlDSaLyTcF1DSse9C1e6k9l1Q0/Hn+ZA4WnmOEIAho
CsZpK4YBReUNA9R4bIQBzdFYAu6W9UeXUbQXMjeelBZVzBjnLLR629ZRrOUPwZHotkQc7PgGIVCo
/BOGxhiqS6L/YcpZqJOr/MHNvrz9uxlDLQocLo8wvgoBRn9+bUi+ES53TvFT0a7rW1umRz/I9agI
IfP82wMktxw72bHjzW/8W8Y9JMr6Tga/AhCsxX5NI60KMg9MDaGE2XosDrs97KoFsGI+bqHCbCnk
sbRRKd0LOt6GnRjS4ZDfguSJuJn7eXioxUSI2MlEmsj44viGTlMNs7W5ShFxKzGzSgsaw4F+/ZK/
Wj97qWOhncpqHnUGNEe6g8gQyoq6l6uYTURga+GH6/tjvQI4yZ8VYYIFhx+aoGdCewKdcI2o/zUP
HbAleZxq6+hcPaVJYGC9nz6qyKgjSK6sV97VplghDVo5DZxoVWd4dNyrG+w21d+P5NyI8k218GMm
p89KPJ2ZYATRwMMRhjkmPZ0JIxRw/qDkbe7YLLuXAQl2Wzl7GKeNLjsywUKsXrCVlWxH1u3It4yF
0afQo8MeHdn5mi1nEwCXgWf5dNxQgPdX9TOhpdzqGA6so6ZmYY5TYJ5z7wx80Cc4Koo9ODghmOVr
fkTJYUjqxbfFhbJfZEbThoJXv5SD+lO1lyCyD/BI6lQzrdneRX3gLpDDmLUsuf3CDSLGHgCgDeHC
1mLxo+qAfSpQdp2oloCuZ/UwbBXOxpuRqam8k8CatuOnMcHpnVLlfeg6s7Przfisd5DeiFPNHepH
LXTwgEtks95s+v9gA/Y2FEFUPGGVbACKQHKGXETFkvGS6lW8yNW3O4nAu68y2yDKmOau/Y74c2cj
t/DgMK7Zd89xgV3S6HHvXy6miN4XY+6dUVgHebMbrhbIDqHB2a1m+8kJ8Y2+1ItaY5y1FPAY/nDA
kJeN35QN77y3omCSQTKA1YLwav00Oe4V/KVsvDMgIsLE2B9bqDisnrnYGWCfJXl8V5mv3iwFF6t/
2v/vASINvRatnsOyyQIJYe4cCtd6DTr+InfttpqiSkK9FI3iI3KW5mHuBzSgMLOYN89zIPdgjVe7
hDbJFQzRJsBarTpqhL4vpxfqUQMeTTVWDfGfVic7dsQ859yhRRYHFsCPiW7rz87qXtkGULCOPlQN
tuCC86xNuTX6yirjeQrYaX1aTbm/DPPW4QbQwEjklEfgAn64dn5MavF0875fdPF+1b67AwodHXiq
4W+69IZ+D43Y4ug3JOf1RJv4qHbncf5568y7NuuXj5oAlmsrOVIogRGjeZgBZivLQ81ZeqIaW4yB
RAM6nhINYCpXW6reCJW0rxj83Cg8s89yERS9Ydy+N6bt74t6i4Xkc0ppo5/5HLRzli8X/GCIAaXp
vSxj55aIF0fDh+egmkCZ/4hx/lswpZNptKAVFVHQFM4NXy3CJef0I6P71X6wXrzx7ubjyLmtubGq
Hd4RDd6GoNFeIkrP+YUksR2u5CnNoKHa25mPPF5dpju+qgY4si1+v9YLrlx7ssWMk0QIN0OVG3Zh
/HQrx3tAqt0QIgeWpeyhjw/7E+kGlwTbxJPMb91eEHPj1SnC2vofJlqo7ZOPXQSYXCMS8xMAKkgQ
1OsAEun6AVytaW4usOgUWqDeuWFXWyLawPQglZ6+hHPcQ3Pc7SQgaox10aubNbt7h/T+/mpwfRp9
vr9RnqV7VTtL3WWotkky0q8GzzbZCymhCPl/0ZKSu9QS9Ve2dfWN0MKaXcyAzOXimAgp70aC3LMx
1IiZGWaYDYppNnkbjTAPUNMR4VHIpT37lMwgXMS/lc4LlebtWphzsigbE6R2S+UG5JIVlXMLIQBX
GgFF/eMqCiH4irT3BmBsHekCNOw12yjXVdjDCvRIfYS2qVB+gWuS6FSWjmDaBVlN+IxGqZvEOouI
HIXdSsH5gywomZ/LDfG770ubrS5FZfPsoq3tNiav6hew2yaEZ2P5tOhiCeypgOiIkrVfmyAYyNPf
btIR/Q0HvIUjWRhZjCB1c1m3/mdWGsQB4Q/G2BnPseI79x/54MQYtyu67PiiM3J6ITU+MQrY+1Nk
hcT56n/6ORstKJpgN6/gY7+sXi8vYYSQbQJ4fJqR8nS1CXX+ea/PCNE/i7vwzyoYkJncULP9JlKj
ppNFoKKH2eH7kC4LmFPM/wyL09cmaHgubiR5aSplybmgO5zkveGUY0F3K+/2gyb5pDzVt8qMoTAV
bn0QiNPYRhvUlg2kDtRCJgMoRg2h5IBerocFlfONkFiHz2j41RhDbxupxYgJHsZzFUXmW0KIbJlR
Gkv2532pJql/ptqjbrqaZXHH7TegnAYJj6rHBbHW/OTfvLKkJolHk7igbgnFVaj29aVEj7w/BhdI
oXvJLznNyMM5micgYunJGwnFrZw8wRY8SbTw6sM3xZlBk9r3FFfnQo20c1VgtTCUFpbYu8pkXv/4
FxvZl2avj1SyZ0RsbzHr11VLeS5Mgm54vwqs8dsYE+fBArJX7CkWOsenv8hg+HD1vT+czfoClclS
n6MLp/LmadvV9H51SYSP4123vf2prTZGbW2pJnkWijhJG38kUkheehLNl/A7Rko8F5ppszdXPdVp
ZIyJLtZpK/6uhHpdGbw9+hy5g28dNpnJRvXKDaFiSXqjJ9dwK7nlzyZQOYKQmK5w/KE/ylAVaLPl
9hgL/uUvOpDDFVSSg2eFy1lPIghIGDgOoSReFSbpZVvbIoTYyHvWtIpNuBikXH+e4YHy/PKSijr4
+oy6N6KLxsy28w+VeP0gxJvxOMz3VtaNQ8HjGGMhc5Eb0DAKn9CH27mZjmkKbqOQyydZ5scv+UxK
Ya2pbVL4jSSy2iqSABuJEXx3/rkUH/4z5lQT9R/m0J2lmyJD0IH13rMi2FONfeLFcYsf44ePE52V
mbR7E3DmnZtOA+m4Qxm1x08hQZ06EgHZGg5w23PKNQSct6zFvSzbym0XfP0c7Jyn4oDCTqtNhnE5
PR3QeZhw5tYW3iE8Gz7WbBGddZaQlf/YeqYsUw6N+9qaABhJjEdyYiM9Aztv6NJJ70W+HqMra9vY
aJzm7jMbSNqL2rrl1lZXhpzVvoCp1gSJcoza5rdxCa/6trz2uayeMhzVsWn1n18/CYYubaViDAJa
or+NeOjckUqGj0DSKVV3ncv3vz8VoXyS+prMU6JEn3AedRDBecyDfyt9di5OI2XEs1NUUBnZ/ayM
+2+a+nfdySs9uwoEXiBMpZ2poMivhsqPf4kVdcLwUR2pp2xC0nb+8nIOmSdX0idn60VxLDmexOri
9HXrr5/ERXiCswZVRdEQ9GFUItNL26NI796laEnyn3zj+Oy9w8ETqpT343AxEzI5IR0DTiNaU9Hp
SxcD2OKPWCMd0aKttahF0T0ujvjQLRNznlm/jEuA0RPv63YIsqklZnQZmv7qg7OGwQk9J8RGlqgj
0FePlSCciA+/bA2huvI5NX/I5pzo3ZNDmUfN7Y3UHoj3Ol/5NBoLmzLCwEswxTWDpKa1HEJEHkq+
o00wHaGbcXoV2TZnVIrMnx5SZ8tNZKnnKY1z6btBtMXB5fOk6ydzwA5qWvw26/GQulie7PfIPU9N
03oEq2Am+7GcYUGi7lJ5ASVfyt1lex90ZEvM/droN1PkcBScIrqj36DU6AJbhfWdHMUA3a88Mwmr
dGTBx3E2VrlNJHh1cGiFHNSstFEg3ULoN4EOCqm2330XJKdgkERhsSuIzcKt4RnjuHAmBNDyXlB9
FRMD812HVXlwjIs0Z3yZN6vGV8/X9RkHP9H9hc6PkAtMpGWbmw1PuSJaCEaoET6YZNxAQVST9EyF
25Fq9UuqNhXGvRRr4kvqoduDUE8HEBnqNCaWm383NqRcqfN0qfLMQf97HDmk3BzEG5Q9dnY1VSzM
+QxDV/jhVIjxykiXi0SVBCSDt1Q+KI2qFQdOMoErixcPmkoGdWEgrmVVpMj2xqdlpTmNhba++WhX
1SFxOrWLyS+IFgpJoyRVOFKI079xJhSeapEO0z78g6yevYr9D3iL7e4+WvwIXlV0I96esH9f8von
b1WixIDexOozrJBlADpw5IG5twBihQAQqH1l9ZA8Ta3R2MURxEA74Nb1CvPqGYLfVSDmOOS4ls9P
P5go9af4RLf7jmeeWVOIMW16hbJ7J7x7J/WmBv3E6rMjvP7XrB7+aob7b80zHPcxOJs+i0iypgWv
r4BGdSmhoDMyWKVx/OjeNuCBdybvztKk2BiFYmjKIDh3YCZem+TiS5u7c02fp7l4UxyK7WgMmTcn
y9nSN3cyaR1HPCyYIPOKimTtyLGbjdxIzUVARwlUvm/iHUnfXwmuAyd8KxP5y+BYiMdJRGGuieLz
tk0iUVkHhYr3ik1djL5VY+tm/AM3eXD7RrVd029O7dJXW5NwB37MizUTfA9yXFOh5ctNlcjpk10K
LO1ibhfCX/rSjVQMI+ViDHYhjwVQTFMDmmxz07oC9YTxznUBaYXRfoZla7KUl4Ab4twsIn2uGTuq
6TrjBtC+cKVLDxiSoGQic6YuAzXrFl23YEGeqcI0i/gX2SRExHupb24uHeym1MqwA74cfE/cLhki
yIrUY89cy984MEATOjvSSCk7D0Is2X3G4wBXYU1O5hjtxOpq3ZfCv9S9jozFyEHqL3WGRqaombmD
u6vbC1XuSFXbbQ4S2k8CbCVImrhtEDUpoaynx/B8IzYqDSTNe6tWixKYaeZvwLFvVDYUBV5WrNJ2
dm8DR+4vQ411/AbOIQFThJWTXe2BflWin72FE4+weYEmqdyib4uMu7E8NvPrOflc+Hp5NG8JbRZR
z7cYdcllJJ1TmtpaGS1BbnI9+LjhRst57/aFHZoOomfGT624ESNRFY0mKYJGvfLaEGG1mRghyO10
yoC99ZQUOxLFSV6NDgjaXzklBmPc9vXhb0it0z/ngl2NyC4K8T5kqDdylEjtZ1+J7Rjf8MVvzvDV
oU0odZudEtUYwU954nZCGoxD0vZvSrkFo6ePFfWNWLwg0D+ql0/VpGGCuiHcbUp4C+2Okc5gYSm+
15nAwzLAjVLX1yj++7esk63nX5rP4kDIYZAscPBz7ZWO9MP4hrRGrvrnYvN+0mAXwhTK3kw48q1X
g0p19qJ0QcG5z66b53vEfP4WnPmtmP09Krw/vJW5CLulVRbnoZLIStA91U4MkrtxvLpt+Ts7C6YG
fsHqjBXoGx4KpH4kKbQGjCMJDSX+9x910ovC6N9rtp0g/hHbCjOyW7kNmXjSDYn6ehWFw0yIj1Cz
++jXTzWqNsCHndP32nzNNH2h5z9cLMPMZK4KwInPgw2pWJcfggRlMrLMA9VujPuBCrI6LkYTJTNs
89BoFsf45qmYdf4P9BY9NSFqnkiOTki6tQUFHp4+pFK56ISRP8GRZOWrhxo60AeII7Z3xXWxGrjh
dLmSPhX8Yh+CNB2aXZ2NTb76SkubmVQPvYjFbnGoqpfUEbB0qNmUFJdd08icN9a+dpMizPTN+PLG
QMA5rLuSMXMkhfILwe5GqWTBsqm34lEwPaDI6n3Bao3TbkWKxa5mZ0hZ0TCHJHs2ikhG2w0Dc281
GklGSoHU/mE3e39VviSEhucdT3YVYDDHAoBHbiaikgNWHDH8f8wDSd7xn9Kl7V545xg1bJS49GGE
HKgAE+T414NerBtfBdZiEn39CKuR2XVh4UfkhF4DI8i/voYyWxTEicG5H/Pf/f5Id5PXhH7Nn/JI
HhGVhHEtwu+gk94erWVmvGlCzwrHnPgAnlI2l8Hz+Z/Mtz9aG3/7wyGCVqD9JltoSz4n1YgaG57h
aSJhw5vsI5tk07/zXaar5M1ssgnjYDkEUbI7Am1DIySyv8XFAqAqUztf+H/qDFknzZMNLOr57TCK
aLp2ia1hglAtJQkB7UUe+q5FnHUwmHGQSXpFHVwFnnL5qAXyvuSIhqDvP/q80JxC0AXSfSy7al5B
RgFT+OBmMUfxr/T9LfeJC7m6haneecTi68a1x5Dc2W9nYyDQck/uqPP2SKHP1326EAT0foXis2ku
G6IAyuVe1MudRxCdD9PrLOlM9F+JGssTIM6ZKSoOiU6XdjMj9TTOM8yIqy72847JbYjAqF5LR7Ht
fO6f4ej75PLsLPKRwjubI+lCxTf8u1fZoFTWYBMaRrtag+SNwGOHHwvPa5px7Lsfo2dRLJaxCiHF
v/4Be7rNOj31ywKSdrhXLEpPWuToA1vRNJdmb4mFF5N3mVvp+CwzophoFBlTGmyFaPhREHztXNII
UIdBzEb/rMtjSxxCu6jf4Ibh+e+T/Eys1vzXSuad0jvuXQEPwORF5EB3cAXl7AnyiQpMxjouHPzG
VtoE4HXYS4cNU03K4v/s1z5BriQqNAJ4UoXYCNVR4rW725vpcH4wWikHXkoxZgMdUHA2Kvn37iIK
5oKtlr1KFNT6OqgyYF3wpJZEdweruoctkjyIprwKjYtsddWExHDyb1j9W93fACsee0OqU5Kx2Sn4
+RGYYujVYh8FLRSa1EF/uUE5vsu4OluAnRnuXnCqRU901zGHvXPoNA2UvR6HFup1YvGpA0Hi+mJy
N0puZ3sNVlqrLGHacjfkKIWirDoCm2AXfFh3WeFFGr3C5R7Wdxob1Nh1dXZmwm34vGob10HbiOWl
BTytJYfwX20brkfwolnt+JVq7Z4d0ec2/33exRngHasB0jeFDXQEJnpPJda/0+fwig5bzcSHafxr
nZ2KbRgPcJeRXEt4L/OVW1sOyMtPZzIUUsOVKV1dQ4VD+7l57vzRk6Uvkm3OtiDsUNeI9XzrZrm4
VU6G3F80wY9w6cSGDR1m90kwzBr5gZGjS9WuChAJgavNRe4TQ54jF5ZLm1NW7DS7drPJlVvIeaiR
zQpG96NASbQnn2jZRhdtEo3soj24vxPGwv8JaQ+OxHH2CyNCfNS25TE9O5wW0lyHN6s/f+En0WT2
Y4xGs6sHC+PW+tnSO+k8cRkfIVHnRrT2gG3Bemn6ERveZj90k3v12/bsPSnneQAvYy7WP6SpIw+P
RaACqo24y63XQqG4qtssBOZScs8MQ/ged77VylbFm6gx55ctkb7E+skOYHQA5+Z3u2d7FbhNav5h
j6H0DlcNrv0afXXPx2CIdYPVKksBMhi6nqS6DoEHrqI4jTdhnO/+ZKkVeIHILDcF3yZCSQMaDQD8
g6jV5V+oUd4au7F3G3A8aVlCJyoktMRTVCP8gDalQg0JD+Oj4rQwsAozmrjvj11a27QzetxyrQF2
PP/W9czJUqXTedpjZrSxNXEK6Asrow5zwT+5TMewbdzKiLzSerANxNQ0u5G79jyjTlEtCUbigVKE
YKhTiWuWYqelFbEDtKTc/EywFF/YZzuY6ij+oW2UYODEJithEiJkWc4QsC7qaa5nX89LBShh9EgJ
OSUupAc3hUzR5bG0CV0QuHbmo1P0aH+6ELDhDIPpCMqENhf0LFKcCjI6oxCiXlkWo7V82/JsipDS
U6G2Bn3A7sdJobDVi5ht1pL7Kr/57ruJjbUAKZ+NKMiSnwQNQ6F2jg81dQpDms/xj0v0Ol/RUmza
x3rdjS2xTJ1pQPR4a2LVmIYQbPZ3D888f+5adDbvIa6BqWKXDxN16QJ6Xo+M3FOgzIDKQGLouFsP
OFrQUvrDU9AD91r45ccR9Bm7i1wGqk7/C+1pZH4Xk5JWu0rnV/bD1cZPALcA9QUq2DekMZgEAoTj
Jt+KLUVHOfRZpQDCb0FjwpMik1TgaklYATE++8nu383t8uVegJHDtnJCUcim3EogR485x4Bm6uxj
x6wxWSD081j4ECxS0H1pSgoLNm2pQmA+JMuzHKTQRs5RRvKMm20KBPfRMjF5rVFHgY55EN1VsltH
7ztcjHW+gKWG7+AE40iPVYUUYSfmB+r9qvV/oftcYTznRFbAspo4h6Btu5I6G/C6UsqgPfTzyDdk
cewZhaFqQDnfHfwUsXk0kTMKUPKXaXLZP6oLBPUZzRl8fUrlvpE5Kalej6DbbtPMEbCDpun6Qwot
WJF8dKgjYEM/LvmsHrVbuyyTKE0Mgo2hAyogbS1wb7KsjlXUzqHDzhgPatHzUsxve5Pe2J2+k9Co
bExn2H44kr2FVcmHupzCsz/SwOgcDYncezHdbj57bCGieFq2mPyZCE8N121ZEt5q5DBgNpPnpQfa
ai7T5w09Y3TAZNJTQESkWuLqxooOKNTVQxavekKJUtm58/8mY463FofVXOMnW0C+ioKr1RHq3M5r
B2SIvvDh8JfsMvUQSf3J57GacobAUARqrTZo0wQUgngzxym61hLUySlqOtmdRFFBduhQK7N3nKkt
+CUg4jmkBoATUXokMwS6PzHCmCCm3uvR3eugJ4b6QurYhqO5vybHdxl8JKURHyRUDxCqMwNsEhRl
DsAInPeSoIi28u7IgKNtIv692bLZ6IW/zPlqBL46FVcZLl3EZ9YNOQPIvCgjJBfb+q8RuZsgb0lB
yF2jKNlpQUdalB93/WT2m1oHLWlUP8m7Gf57HFtYbZku3EiI8cTxqVQ7kHi0oxNCG2p8EZRir618
jdf12c/+K1rBf9R2IuahZg3GEoQnHmnLshJSr0hWMmPhXEbKAetlLdO1jiKdfsbuRXipOr8dqgVZ
M9uje0gqUCTadxY9/VHV4zoALDTmhMQy07gXUaO7q42hp6sq8pcsbkM5nwEKbNEZrlb6sLExZMxM
tOiJ4wzYALk0y/Mh+KdLkNhXfdVq/jm3WoZRwAk7gEVvp6ceflYOCSyZi2wA0DDWbtcUy+NALHR2
p/gMfL4nK7JkOOKNARqHxpraxeweTCDywDVIftIPJ7FCAvJOMGdBzxDioDOJ6En3o8MW5xX0xxYS
iu4/vwAZXx4inZuknGU04JGZuDRbx3hKFOOHGBA7LJdAVMZgIEACwO1jbh+5u7dkya5Vw3tZ9Usg
UBajG5XQXBBhbizhR+e8rEXoAvWDs8vyGogpJRF+DDcRjUCv1WC0K0ii7OjkfbnyDUKxnv9KMprk
maT9p3ur7dqR5vO5gaYJ6EylEmdT0a58YgOuTumN58F6cDUpQvyVXMiyylkBBzxgFnZptH/4Wd2g
UV/EpV19d2wMgfRv/XQRzgIWYXAS8OrU5IMlk0N+1iNOW2csNLI7n0rGN0mpm3m96CIB2QGvFyGO
JaYsfnoWgpc2R2sILX2GB8RKbAcIFJWcHMLt9TMa78aRvXNzzG1sDAw80I0fsstK8CKnC5PYEVul
RoAbo6o5C9v8p+tpAWctbThnRjY5CPwqrGxmDjmfg5u/gP2NFONIUmHbvtl1RoW04oGkfFc5dX+k
bgr7KYNzJyrSsa7e6SBZogOL9RWdkvbb3cUyU25DHWnXHEGizqxVqEm9TZtV+kYA42bqMpjTMcIj
GxcPZ+yPQBezUfMNPDjmT9s2xV48OMYt5GVyO08VZxy3GYuv8fzlszZ0IiLk1Csoz27zop0YLwNL
JwSQfM28BxYAroLgncKj1gm0qheR5vXIaFTWgKqKbJlZfXStvXMlzv2PROaUOuU7zxQ8olvM4/fM
HpvlsUHwPZebIV9lDNeXSNUyD6Pr5+JbQ5ObOyZkkoAS+cWKUVSNz0kgY8SqQBcZGL4WAEQzyCno
6yBZP/WMLLOYYPYSFUCw4OxYpxE24oVBtP35NmEj5Eq6RrUsAyUHnscT4zfr7J/5JLVthRIIl842
Ct62GuPw92m60eU755eo3Mie6ux6AunsOPjFpoqJyhjR8MRuwJjIY1vvRUf9Co2Bk3ZLhbCkhqtI
6HVctW+Td5PXN7aduLBQp+NVSfxpMTf6Sk5R/7AcngLXL1GpYe70V+VF5a4SmtR0mFfrp9xPpoaq
vR+Ec2dNfFiiaSCClP18715Cc8mWDFtLOHX+SdDiVkHF6U1n2JbmQvS4r/r5u6bGWF04y0MDndCg
2w5WCxybYepH23qKwzvH9Q9JOgwVW4LyjTFDYMpZEAbfEBgUYyvU6pdZfJS2FkznEcUaZWfGDioi
J+5ofwpfnc5m5tG1nBEzfIaIvFMf/eu8gglWIqDCi0Axtt+HBFvkdm388mu+ZbFfeaNl5AsyEw6I
m9xy62gC66KFQ5YK4qnuAXPPQXBCjgmbxr5fnDKgK0FQ2GUQfhwqtsb2vtAQZcqX+pyN4nmlrrSj
uqJYA1ZO/Knm2h4927w6pjEwxvwOIK6KzmFFbss3A+ExQ5Hg9J1HmzbWMxoVDvqRh7AeidfRqaGu
4Q01txqeRzeD2qJHGFn5MKDhF4wZmRyD4dY9P9twFQw6eSUjm6G93qri/RANII9fAjYNOVIWBUVS
y3bM87verli3PTn/tAHWyncZz67nyuLBCl0csEsab1ixcbxHGUwnPG1hgJABYaH5diOR38vZfeEA
usUNEciwaJ+B1/yBz/iWIpg5t1Kiqs7UE0gBw/g+dYQTy7WrNsZcmrLSyf3493SXsRW8UAHRj7b+
IkCkaSZB2MVpfe6g4AwPmnWtA5fmbFhO1lA2UAl75apPVbJKV2WWX05cIJCJp2dysMo3wLURU/9m
Wy4ZexENHzDweJJAuo82ZEK6n75QNXHN5HLgKhR9ZFjTz2MVsHgznjMjc0b6V1Q/phPIUDc9JH3q
dX6ZPoJ2jao3kE6MtEZsunwzMqo2tj8e1FWUyOfYI5Mi9QClsvNdJikC2GctHyzx07+anv27wRi8
cMe1WRi/94jjXUTBG3UKH/I9INkZT9DruHksToL+G1coaanzx/TvNF1iqTkfaXNMePm7NScoh0WZ
gTcptS0D9hz20HTmbB/v3jtsX624TLWCZbjwOvpeAZWKOOT7GG6aWE2wtWCWYyhy4+BuUuQ2dNvv
AmXIAt33/wYQ9iDMDEgbOBY4LhADP77IE0Gt0dFpGPPm43yzGWnYeDLst3WgffbB7ikQUEx3x0Tj
1MGkBm7F/UFTrU9OanzyKd1axFR3s0+II6keDD83r9f7aj6LJElW+5nP+LcQjxVHFGEIf7RrDk25
t6fnSiaMtwAdz3Va0poi3SxyUEqtLjQBYIb7UQJzovTk5ZXA4GNUw8Pc+zPnOM9MGabDSFj8OnYX
0oJdoVCU5PGeHePfgcYdrDxWsFxQkIa6Giut8pZOGeb7wW4e/uuS+SQulv3ovUNYv9etoloW/xne
d8dkG+BsX0XjV1sZcXJ+lfKwL2qxli4V/XepgIubDsUybGw4yYtd6HwbHM2g/Nm/R6npUxb0SmYi
caH86wPj+tBTrVvRhgCh94gYaZj2h3dGtt2vgiTzjp8i4lYw6v4oiMotndPWDTthDvgd2Hkb0noU
mNwu9/kjxzv9nbpfiW2ML2A+4xEHLJFCtlVR5GokUKai7bJPBb4KGXm3xc4Trf6o4fpo9h48aVbG
ZOTHcCC9RxCBxxp5nXJu4PDvwNKs7/cGwRx7HklnQbQrDKRqfyHf3xfyhPGRsMhxofKYK44OTZ94
Q1N2sGtOE0JMSvlt0CYefc+6sLorR8h0G9GwbPpyUHOM8RYAOeC353dXgzrgjQrENaEPXCaDFz2l
QB9+ZbGyWnvS9VMW006efUIZ8yLoW5b7jjBoNhZgaX/m8pF5ym9rNr3JkQ7NAHV8DbMIhRdErJDn
HHL3SfQVxH72f0R50Ig3oP0/vbJo4R6w97LehCn9BEO276cg9a/aTErDHb/b3LgQl+NAGVQRmMbA
7cf2l7FWMUEQgHR8P5EjH5dWgscwDBXSHdgGbxIPZVTgs0k01hYxN1BOysbLs9PRM3YWs7T+jvN4
vR8u9820O6QPK3eAa8ruDKk/IpUhKdfBm9qiQtg0AX+ag7W/fv7XiNytzgY3enqVMi0B4tzjTqmr
SSuQuoMyk5MxXmhKzPdIPZn04mYV/SLyqUtiCQbROdjO0T5FInA+Piq6JmwrinoZTbpDEicQserc
avhK++7yNikU117TtFJdDUWXxhuY1fveMsOgJCEICdMVeR3bGSGilE/LswtpKXkhLQeOXJXHBxb8
n9qnNJoqoSXvmSIwti5kfelg8VIB9I/6ENs8hVTYA/UsocBCZ8T7IDo2zbx0rz7uve5Vg7JYbEjf
0gnlKVZMOD9W/w6ayYdzfIMCWTiqhfDz6jDE5v4yyskAnjwdn5XDYzGefHKlQHFUnzTT/dEyo8hU
cVQ2OuUaRTooN4dqu7SXxU3czQb99/XAOet3sPWEDD8CzRxsegKcyi6nvCluXg6TZ3YpoJGgOn1Z
pb5X+0YlawBez92Iw+MQYb9IaCvHrXzn3I1tFBAOiJYutnQFJnJNPLkTU/OggT3wM9TMK4013fL0
XP5XCP8vYSOcRYGeEpESBvbve0Y/9/O7WFEqfouZ9TDorhqt9umoo8mz2cTAD+FEel1kQe3XSFhd
fe03mGP3nHV5ChF1Kk6uGJnxYrhRyP98pS2hhyMSy61Ibf6hxwNBqaU1duhGy/7KeWJrxfCzQS4u
AS81DN6XoTCXuyQC+QcEToPWVpMQ/3gU5aMv16sMw9RtoRX2TcrK9d78rnjkYLMMDwcpR3Itd+5P
ziDZshZOUG4sMfIY23yViV/ZSYAvAy5GjyDoIFEzqormRWnAKiEruvLIM+l4RqQiaxEKgg5B/oO7
TKLPANqBtoxLNuwpDLFCNQuK+/7X58aH2IM4noAQyL9leARRwXE5SUJwWUEiiavj9Msq8uhBCzwH
JOg6EZ2r7eLjlXgB/T0JrLHWhoAOCcNcs8KXoxAUh24sTemk00UWmZ+PCS43WVwiT8ohEsdNLhc0
DR4fnMSjqpDgVTZ5ylx+Z9T5V5FQt/xFqnZjs0WmgWsS36MErcObfWOSCr+L9An1CwCowLt2V8nQ
AMiTPYiq2mOOjdX2WQ0ecbp02G262I4MqC4Y358ac69l3S55n2JCeeFjlQ0hehb7Op4uqJAgwf3D
28JEzJoNaBCXYiEKBZgasyLFOXYKILil7DEMvWFXb5ZAyMVQkasxWuSDmoL+rJouPbbmX/8EblWW
vJdmBP2UCN2nXtbKGMubwXy17POeKOts4GAOGeRUeKTeqiFk/z99HpZ/AVG8tZglxcsCC8BljvGp
T2in+aAwF853fEwSFroarn4FDrW0N6xy24K3zVDpj6B06co3SxlatHJqlqwBfLYhs2D2ZX2CIz9+
p7OMAExtQOTw7pvICLbXibLoHBYUeR6yExHCEU7Ifm/OxtKi3fDQFXD0v3MM5nQ0YpEAsDn7Bmhv
rgLFFsq51WLubNMr16jPo7ZxdqqK79I2Y7X6ZqZ/8CcKkLDP49ECxkaPL6fHe1yaXiGrvkM5xNXE
bYz2pTu43WUTy7E3MpyY3B/4KTgLwFjA5Vxjqk6vkk2hk4YijifA3sJxU0ouiJKZGHssPsawfePS
kpLIJzF64eh7+F7hTN0u1BQRCDjyHjbYOFZUhUW/dAChjpBLybH4uImD9IlgmSHiXgZPb7MsGMJu
1Qh6pOhexnWC4pOIFn5NCXJzFr7h0OMXtQv1H1oxZmRV29SmrOzX0jrgWF2/iGOoWgoDSFeot+0A
6/OOuoptJZXKAKIxY8micWHLtkP9TTrMWHeYBBNf7HZIp7AbcMrNI5ev79SLsnMPr0Rhhx+3ON7X
Ztsy7yIfeo1fhQNoUH8zzuoaxihUUx66tnhNu+ZEJQr6UNYa2fbqcglBc+5GKK4E/qpthYJhQ3di
MKzii/POqcCs3Zawc9ESqXJ9/+KB5z20BeKfElzdJEyez34XcgLGaL6CbxxqWhuv42ooLNCrRxex
jEokI/9wdxmGbXe+X+DSD/21t2eTm4bCkS7p7IVjKkL3ZogmIYrdTpqMYo1RjXzBOvbL2CqsOdAm
286NylEVEehL5VA3AO1PERPo1PW4HeMmAfNPDmDLh+sxJwgOj+TyjIgLMRQSa5SNFO0JuV1YpzRq
+7wDu9L4GK6CL52+rpGeDZG3QayWOGbs6Xe/zAQ8LKqO21ZGuf0OYtG1rwGAeodqWFNHOJhueFUC
z8EbsivO46AtadfBmvTpuyCTsLpt/IwKh7EmRK/iP8XAzVc4fIznH2EmfpBx7Qp8WBAujwBAUzqj
n4cT1K58L4z4ocsQuZ1Xqq5ND7fY+mfG9/fawcNMe+ZZAYaE2sOMbqQwiBI5QJDleneGZf9f4d9Z
u/Csm9GJYWvUdcVFEi5gO92/Y5IgUW1P7a4SOapc6wY2kLo+qE8iIe7Vw1IGvLOYZXsQW4EhIQCC
mpWJkwE55Rd1MPG2lhz4aCCNsP1rEAAX76JOZZpMO5QpBFwz6JEoAebXDx6BO5dnRistgA1jwHDO
YVa2LL0JduK8xq/SsQlmyJEjhHHrkPbhQnu2I4xOIpOw4HYrwO4ouswN+qsDFrxIIdx341TXGKnt
67H7STSlams383gzGjGtEX3i1bgmt9g0gzjgPeq+OJ3AwMS+K4bScUXuGZXhlCDuNTkV62StO384
uVDZY/irLvtcvT3eBgIcC9Vrk9rTkhUxGtRJ3A/iy5xjPOpwZx2PKDc28oKMnD8K97PkTNporOui
iZujfB71OPbzfoU+/BcrOYsAQ3KY20j3lVluF+JgqxcjRHMIioBdPJ8szcpSlHH5DrfgG1t7Ak1R
SS1Qg4rEbLDTA63fWbg6pKl1oeXCKpWkHbvzByBB729FcqRB45iqYvDMYdxx5AsZC7uN6ZP52hw6
aok+L9vYN71gT5JL94tchVhsQYBPQsKv0nUru6rOdFtBheoFI8MvmiEjfMpcI/5LS9jZyXSyKdK2
wfHbKwRtDy0X1GzfF9iXBE7jKK/SAEWk/ChYcQPeNvixrY7IbudtZZykqghEYB4kY3WgihR0mUWi
Mroi2bRyxw4QIpE/9+Gcn5M/6fU55F5zAqCfG5BDYgulSA/D7Zt0cTwbi6Es4mPxlFNoySs7XSdK
EMN6RAIE7KcoYr2r3iY+pER5zJdkl0CbA7lxaGjOC4GVopOupd+0uBtABNnN5w8c7NSbBPOFKAQT
eGxNyPRMWx9n/kr8PBszaY0xZTu/wTeFJyxUl1Meb7kBqbDWUd31B/DXPHU6UizUKYLfysCZvXQv
gI3DtN/RxfGAZi1qIk1KVGQH2nNVlLjPGX/WOKk7I7TgeC6zAOwVMj1kQOBqjBsIG9fmWMpzcbWa
cm/47OcJaOGrEtOL96tfg0hahvIYun98AgZPae/ADtT6d/5nKmwPYLmqVK0xX+EIBD23mhY2hcAa
emGgOxLlpvKj6AtJyyQMZJGkev/08CV7KnpAgWlCCY4s7hKWrLuiyuHVYH+E4eGNDbERqAjAE0Dc
pKLjpElkmacrpd6i/jd00K52E4gEfLDcoUCtMl6eO5WXvC3WY3JnaD2osX1xQkIfj3FfkicbodM0
gXmfVeR0RQ1Ct2qOdMhdq/Jrkm/LjYTkxSwoi112M8lLtHB+XWhZre6csZZCdhKcSuqm//AjQBMd
0xkBhaygK5m32Dcb08PVxYwAacHJWrwn1Akbvr4DobAAPGR+TVD/U3UkOhHTXOllnDd5IY8EGuOI
vwzpJYTejCGRt0RJAfRPdgHM9LuQMbLla5TX+/SS9nf9i3fOLmuI2RnSx264LT9/tnsjTq/zPSmW
4yBgihvJmSRZU4DIW6XA5WT2peCT8jcnXYhgPToFHE9uiaPdMkzhx+jmes/Y/Em2d/ivhKb/3Gq6
MocOS5JzqLb/Hb+9nzxgXXHeTxXaoD9w0xEQrglgXf7hxpyR70s2XZZFNUDnrS4rKjJq/PLrJzlt
m43fOUs2gNfbhuDGf0SSz4/cRtsEGVqtOyPGOtfJoHOB9KpnxS9mC3el+x3sJWNE6Xxbw5uZ08G6
w10YlBgISrYzurhP6JV0Wmfx1ausZvqkkkL/nSA3UA9KGp2p84p76O47E3F9Er9S7he9v1gw8kU+
6i5XvKlVMXYr00GaFDMFh+CrCpt+BZnHd7Wrldf3mAuukAC11QB4/sdQoFTlHjXuPl65kocx3e8L
Mhdm/U8vAWTmSpDaPFAlKoVPYXRAevz12QVl0OCyq/Jgl/r+rsuHx+Fez8D5IW3IKfCOClkP05NE
CAHEq8umKI47yuqIEgkjRk0MaioLntafAbwt8VFRXg0da489ouHRYWR2NIj1QYICK1AFoI1QuD+v
4aDAE4QncJRFjmjn0EYFR0dcaHoUu626WJeC7nInxKtNV3MH6qQasow/W9NkQl8TraezWS+xBsve
5XHir7VCdcFyRbPMwpMRbhMvtY/oDLLPV+/h186bGJdIPb/QdrnsvR5VSvTuUQ1E8/1sHxJF7/q/
oy/G0+PbVcCC0500ozPxztbUgsxlFGsogIo3FztPCbXUZOVDDjgnTYIwWIHOIbwurogljjZdtgWy
no4rLgqx9LMfOX+PgOoh3dr7RER50IA63tqJF+U5Hbk1G4WWfiAb3jxnW19Ij1s8mfS5ea/0jfM/
20vugSn5jgx/rkWkAzRq2wEZCnXh2aEJntq3eUKCXr0RbVMekyYrb9NkvMj7XEygKB6th9DZLRBw
N2fuTrx7Nd3t646KDQgQPUNCUz4uNAr1I+tga2KcsMEJCDtpX0YtLwgBKFb9ypPQsSr8MKWuN7qz
o3NJrNiatiO9zqrlzExrrsrAMLvEkmwjMzvMjEc3gJk5JRBRSDfvSXdsWNuSamQYA4Xox4aNY7eI
w3FdMMk3J8FGg9tvOOg0flaZHK7eMZ+nG8B3SxAWeg+jfxv7ivLEToxmp1r+UtYVTBc9bS8oo5Ay
81IPo5xqGfaiOVXwIKjZQ99PsLbZNpKQcY7oWCItHjwUZconekqVCHTTmRX5Lkc2/wlKtRGCxhGN
peiZwkJUygmASoXVBUUGTUyBapxUA8fOftR0oMm1/0WU04MeFN72IIUoP3hpemzPgfZAjqeIVzjg
JiU57Kp8EHnOFm4KXxrzqxKrpWrUixHVYe+6gY5tE12bq+I+CfDiS02vE8pY49CkHtCPqIFnWejo
I+dsCY9fk/x5TdckAlDwasRoCV/bA/WI9F4xON+z5IVBDr3BO5Q46TmMLOPj4vluh5IoTT89166T
shvaJX3AncFUVxisBY7s7LZ3jeBSrebAjZKVf2W59fTH+TfBZVtseV9xTIWySH2NqFzxss0YJ2lv
a7UmEb4noDMzALF7YkybJeglcgVsirBjYSl+sI0lZK3UNQmI2rkslqqZT5USpWp7vgZPK6AhE85h
Bxhmew88GRVVEXUgAThqREs3CArkpktdBg+nY1CeP/NstMl157GeBL7BrIUSGlW7qYLeKLkKGBJi
KAVLQaQU99eV+VSHBa4JVjyWLIo4Pg9dFfm3XQ5yDu9RJxOLJ9YJzatIOn0C2lx14kRlVhO5JewT
A0KgMHbKh4WGH0UTmelcqYsIzT7+6xcTPRKUKs9T8hWIN712NObkf+deqUFAkKpOb+pmvFO3b5XG
9kn9UH83YIF5Ztz+oZPT+PbhDxF0ZTKElxddc2jIR1z7vUpaJdu1L2OFjMeGPSQte5qwz3maStZl
SgFuy8kvRoZJYwdUzGWJOWcmT7ZY+8zMPiVBw6ojx0OTCVQ1BLktAsCVpC0A4tEdtLtPXSXa/oEs
vL/+tcg6ty99EwHHbpV0GkRMAf1XGGHC+1s4X8dSBv1nYB5FFSvIornh8bnYp3rLUXgjlv6XtQZz
84/M+y7TMfiNF5UUSxu5uqcnLHjcS0YLJox+h4T7e+vcBkVl0nv3hTSNNW5VFpVjxFiPwXxbhG/B
JIdGlTpxMLDTlEQEDsDPtb0hq+oYJsUcDIOVkfbjRh914cSimInpCHIhysbXQrJrGes2hURG4aoC
jf77YO62yuoZUu1viT1hYw85ycGeWXyxdApzcl4rliQShADVYwfPViFdMbT59EHr6PQ3VFodfi2J
vSIAANn59G8asfnlGke2eqUUIrI5t/h/i9wzqxHePv5Iti8FJs9qvOgSL/9CHYHOxhXJgZYi6Z8k
PsFclgbxFAmIpdo2+VhbuLQWqj7QH6DOOXAeT5f3hfKvAgNqeZfUfIkljuC2CyBQ2uqS9QWXq2hz
JY1aXcXUzj2Al6zVCFGr8BSKbux/BzhWnMWIuQ6SNd0oQaliYpA2vZv6oDsfUKMKhqcdVQhkwjtq
KIxC0IJxcpSG54e42Cf/0bQQPpj6z4bP7/QTMtjk148r2DPNl5oIBXpDLHtXtstOc96zQndjjAim
BjzEVlwaE5fX1tiYpbC58n8VtTORonmI43i1JYJQ9+Gp2sZ52eI2VEXwf+XEvAshQdT6lCvH7VXg
oI5r3pQjkj0cB8HFnNaPysyjHfh8ZEGrfwerR4f/yym/2FXQ9/lfTocwQqzIqJXQdmgsdVfJjrDN
HtvXpwRQXvPFbQX/O+U+WvXgOVKfdBI40dAKAg0N8WXeZGAPMqzshDRgBIIJ5EqXwSAvKuk9eJBF
GmuqGKpeFxukN5xe0Cl0AB9Qx5W9wrIF1bMaXb1hZ0V0fhC1FJZtmSBv2+6W8U+K1HytZ+M7CUJW
tdWokapHNVQd/sMGhTbkjPxjYepe7Bp8i3mzABiO8I5sgS84PagXX2uZUQwl3UsR/oYZU/mnqaQC
uC/pPvLuTHVjaKrjHfFN6+FGcuDAsGLUt4nVdAINh0azOJrf/aAiw9Xe7UtQ+N42nnM14ff7xn8+
5fFAdzdT8NAlgb6XdAxHnq5V34wN4nwuzXRJNkDl/+QsVJ6M/kDFHqqYXiX8W2RtmyNzlmK3lUQn
4CRF4yyPJWY2S9jviU4TrUB5BZCHmX2zUhaWDlAp13+BwmRJ158udPuBEgl8bkZpG5f1vgfTrbxp
jEsBMFFhYa8YpUz58tsXgoWqHpXS3MAdTMAbvSV0q5d3D4ouZEhXBHIhvwjRi6aTNpeD9saCxXaG
h5G2oms9Y51O98WgUm07PC/+J7OyYBvnHFmva++dIxeIdklCq6surFeq7L8f7VON2sgvMskqk3+b
0BLDlcRBPMCzoo3kKDdGljs737o2cA8ETmIuEUuDfyPhCA7zQjwDQFCRiqL9PVZ7VB4UK0Bhaimd
Oxg11rPUYt3basciO7f0xyJ/+81Ic7792aCO+6oyFTo98QQyZQUFpqdGzER8RWyw56B2Ip5Us4mq
QNsrv1wJVLpgHrY3TeBoW3twdTZpsjbFOdNJUgxzaFwC2Yvt4FzCTYwE13XW6kTmIeRR4HXTwnX2
tKNPzbyX0SHuwMi7H/mXafQNSsrrkzOumdTzCM92Oc2qdUZpphXHx7uKYV889H+dN/KlDC6TXJH5
HrPkIak9rpeWt5kQmAaaURtGj72jUCv9+k8NO7Kq6er5ZJxr8Jz1ZPp23cTIf1+LluRKOlwzc/IJ
+b0cFs1lbv29PSX/YxO9uS96LrJQtsUI40Q75IytvgJ+7vrHM9dWXnZcPUHcLNB4EpSyiX4G4vPR
Q8VZCD9SM+p/zNjccocDGLMu9MCzZjFfsXcs2AcVYpEtR91px8MgeXYt6YuKUecR9rdgrTOsO8L1
4GRmD8rXtisgg2sELdI5InwK9cNyTvjALpoaZyN4+GMg7Sw+iS7CwC0z/NmHpaG3yaao5o6HHZZn
1S0epjTQ4ozd9UAIAoy5/hHjVTSp49bNyFXK3pAsurqgyn9sBrXkzYaPD5KcTbzXjksxXq4qissX
6FWJHXrZaaUFsVHLL0JTeG1+b4Qbr3xzkw9AL6tleviEJ3FfPBiizzwHieRj1Pb99s/e4TyE1ISe
6w6ZSdJsEccB3k30xpMQlQbh3+1RvyCIaQyZv+icHHvbJfGv3DxfEX6dlFK4HAyg8pawSUvNinFl
NxqiafcYNho6ooW8WLZ51ZbDG8aCOI6I6oscg5KqDj+aLeKchF7oEPuq47E1OmGkJTJ/RaBpX2qi
Fp7PFlSVq6XHFoE6H55PZ4okvMf0uM5pBp8yQOrtzM5X+mT6ZPxXmjgEf/29yUj/57jByoy5YltW
vNMXpsJ03Ae7x0FmrtqBo/QjvcaddrpoW18ahux0OT17EyPJL/lg135KqmpFmE9UxoLpceMOz09p
S42OEHaNKq2frTXOyH/t7iL4gGchVb+DkuJOMzfqSoHhc5I90v/XXUp67070CCNkm6zy5CJv2Hgq
FVzVMLzYOPKC0tQAD8iTb+YgYC8Pm1CB5hzw0bvmuklvBU6Zj/Pb27wRzLtOeb5rUZ1fn+YIjxtT
E4RQK+P+ef/dQaoffH2Y3d1rU5cjBWjbiCVAafzPpsq2Vmin3Q3qLXWHfFKSEXWU0uwk1DTdQ6v0
0T/piIwFt9JybDoBBR5nKl2QUj5oJIyGK+Gbuk4MGzrAcelF0BCuK3GzQmfs03oDcYzm1K0UA5Hr
YliWb7BQe16+RCmwET+mIuOuhvBlO0iorFrG8Vi5dkE3m9edLnyTrwjxW/h7hQK7TJC5bWOdGZX5
U8+gSNwlgMJL0w8d7VZBd0a0OlgVsJ3BDQtZ4eEIEjb34HwVsssVonsAOexhMMD6vJl6VfPjCyYu
hBp6nvGm96n0cbR93uy8DVnJAov1ZmphoDwWT6nMbkzJyqZ1q2q2zONeK63orMBfFZYK5kGPchYu
lPG/LLrVnJIaMkaRAOQnEZK+MMKPoYd+5nP6JYcisPAtUUheNU6d6rYjcqvjSZSVkx2nhotI/Di3
ewKBye5DgmZ/nt9EaU/H2D/8O7StxXTZpJ6tcM9Cc6PGc8euaGt3tGjWR42aMSP3OOahwLu8kBLT
yvK466V87VlzNPwUTE9HrKF7Q5anKkJLIDpirf3HTgWNq3m8/Fy3fqYstkhR2Ekxm4s/le+o+Fy3
KKxyNgklMWm8IBbjJ3qufvT7j2h44x+JW0u9lLIJ6zezfA1ik1In+Mbsv85L2sOgOGM93+jc6fow
zMjO/+H4fz161wwWNMgwCa7a0wusZJVu60zvQ5eHeIPds8qgSRD0z0XnBAQppuU/srdH6uT/rQth
ujpNThLb7XhHOfaKd2ZwXDCyoygBQQ09AWYbr3AFDWImXiS/1DPxg0W9oIlUlR1KQ5DpdnpOvsZW
A9J1Af1UXdCeVO9lYcJWJ3Glhi4X6uJE0XgZB/JWFJ7bME8SM4IKhZ46Lk9R+9zgSMZg8bnRcfDs
dQmv5CDvkVL7WKXEU/gZixNp+5ihIXcE8/Gzxgj3E1NIILEWwcVrCMCxi89p85iQMzVKneOF8oAH
6K1xZ6e2Y7MPlkZz4unXJNWVDwe2WzfkiLk4ThZNjiHMk9xSe/kNYSNOS6k8sJ74isrmGyPdn5lJ
4h+fsofD9sasWUpQ0v/24Qf7T7W9jmb5eVYW/EVHS3ht6/SE5sf237coh5tD78pxOjFeN8zV7oqN
uluQxWc52fyKg0TfQRm+J6xhRq+ojbVaQtdsNJQQPB1R6yIeQO6Ci7dC9RLEgTlgGmqqGL3g3A5r
VwjAMRTxrWNhrTYda6jCOYsmRznbvFFoYWCHRAG7jnj5GL0X9v463BZ8siMEzyIieNzilAsZWXSV
UItKWp9FWYkiJAnMDcqWt6K6uqsnhzAEcWlrRjMaT4XPTzz3KezP1E+dnF0oZAZUa6tS26HgKPX0
5Ao1NLgIiRZ85KCCEP9mHzk12LabQMYZWIwSmUZVZLNQiNwJGSw8r8SCRXinHjXczduLt5OjP/cM
ZTNhL+3H/ImRtObCQ4tqYqiQ33h5/HofyJDpuP2uSv6ooIO2g6VhfXUrQbJfBOImYiAzYR7uLuZR
zhe5YRSFQZhAsqpdOpwBC3nxuKLvvkEyvh4wEpLf2EkNjLJvjk3Sis6oHbdQ1RGwWuYutgh+DeY7
pPpOpsdKNl3qOp9eZO+rouG6WHZ0cd9G3hHCgd9LTLWq6d/BV5UZS1YcgXhAKvVBKgb6des4hgVm
RoMEOjb+8EkEIcoktHzbZynyFIo3iYBDgz9MjM/sPNy6BUPN7H8kGWxVagKLRUIsqnsOUP8l+gAt
ySUzcn9QS4eOr6hykUBNAiiKlzcI5CJi1sPvZVufQtE6NSW99QV1Q9CJU54WbRKifr75Xh3Lodmb
otEmL2QKPuEpZQqxywVIk7Z3RI8hzK7iwrjxZk1D/GXdGeS/ZoULogZoa1GEhrqDYYCNvR+QzMV3
lnWyB9wvD9N1zOvn2D1vvGnauagmc6n0okEtUf+49io4/SEO/P9fccjqkEB0/S7eqwe5MGO2GHc1
OTj89nrLleRkqGSKkgOmqWh9VJDwPQ7gaWXaFnH4iupxKbTNrBKRg6IT75AYuyj/Who0CrUdVb+E
gExlZgbI9noUcoQGMQ3uZF42PE5ddZpVGbR6pqZrNF/ss4+KfPgHZUGZ1srAqqZ8BrjF3mMiYfKS
JQkadSRd015PR0PKYuHAyDjibH5Pc3GS13+vwGb3hhlg3s2Euqzz1yb8BQLxOqI/YLQ/pfokJ69T
KWh8yIgOLAd5dk1rMmy4cNq+9Dhfvmjbj724heNhNLOzak0nVEcTPeIu2tSUQNjxR7J7hFoDttJd
NqrgRNvDXP5sokJMD6tS/eFpgzyBfqb4u9EwOn4ZXAdURdL77sypyU0ubgM6r27HwLzNe0XN0yH7
d9CrTvKZGgWnD+A++xmrCW6Hqns4sFjSP0R0LlYKMzELGJrPpJkLrOaL5PIGaJjo1gwqOMAWL0al
dWMpiabjqyHiiAZxIB+V2aEoR24Jj3S9VbkfVpl0m0ufjtcjMcrohysSzaXf/EHHnfoyoQlPevTo
Bjcooy3SVsp7om+GtphdjQTz48hT1r84tD0+RpcRoqMNK1x5ZUGXCyIlJZjhXigCYPgYLZQv2V41
nocTeO07D0XCJKVmAo+DXVfw9E4AAxEk1N9Ej19jX3HQEF3URbsbgwJvp4oS3zd/Vxsofs5sTXYB
RHnHhJU8NpxNWqzqX0LBpUugGbKCl/OEtyYBB+2ZFRkGXHk2w9qwmk706TVJGzgFt1bCQSzPtzpE
0vio0n7UrbabAdToP+y90tb20LZh/GTHQXO+HrQypiUT68cgsHiVOAjipYmbnb/3Y9SlLQahw/8/
HGbn80ySLNYzGxDksvQ2qvitK7NloPmsxrJ9AkxlpvFSD0azIAmu3d9zyUlcXmoYtfOtPAuW+Vs+
3Sm5zGvYWnf/tPPO2AiEDCciPqvTcx7sgTtCKksnSYfYclT0CKPgwdPGlDHG/0Bu9ZK5XxCJ7ER1
XTRFuVnGi+KQS5yN1jQrTQ9pFD469H1GndD8dGeFO0/t5cA2KJr+mtVu9iG+MYlpM4XeGKoW5jBn
BnfMmuLd77On23kxGwpohRYWnGX6xaiASq3F3ZegjKQADvlR7l5mhxp6wLjN+U3qD55ulhLq+uHl
U49yJJT3675DLcGP+yZax9MqbS+QX4zuFOwXJLp06lhWKwNXX+0sbMAzCpoE3YthWFU1+DYW0r56
7ebPmtVSY3UHf3mG3OF27DXJS8PE6wg97oFnv3hVay8BsFhwIsDt/usrF7EIHwkgef/o9rEdWiNg
wyJzeHsaOYuOblUHKfNNID919pmNyM10MuMlr2s6B/H5EafIpx0/ZpFgOzo4Q/OqTozG5Pdhzje+
0vr0Pgx9GQSx+cqvRIhIhBB3AiB/KzSCzQ5MmrRPT8ax8MEVJ1SEiEy2NaICOnNcoKvHWleuxdnb
erOKZOGjAh2LuZhFk6hYNQpBYv6mCVVHtABPULrvc77QJ5K3DNTqFptQRIFsiXxxnWxekzWnAuJL
3ycnLlqwAEfzfON3zwgxnEbfnWpIxtP1r3gCvjjeX41Gaum+caEOx8Jmjul/JXIQXSCSYo2E8cet
lGFrWrx1YBNm6ydDhA2fk2Zf2MimbBcSiJ9Eq45GHqi8uTpvqzu4fvlZJtOnGD7RRIP453tteSZ3
IQxXUW2bIfn/SRiwkpuksCjxNlptC86wKNdSXvxMnS4UD+hkyAYfMj5iFWH0fXfEh5rGDPbirjOS
z2SLXJ/1oG7kahDQ0xgbZJ/cauKMOeR4FGJBkezF24GQuv5XbS1zxmnl9bsCrWFutMvXnpKw8Jfc
7N+BOXMUliT4px7EZ3LBaCKCcg9pCF+AhFe5i1/UGAf7hC9NF1M6ouiEqqqOQyyxaPYQrcb1ua2L
Wsm8MUDMT8yuuYRIdYbnTcki3rh+eKQqfZpV7dMZE8BlctPBs/NstKuEWyhfSTD50nL8s6Ffg2+A
PbQqADgHcU8Awtp7Uh96tFKWb2lLmJdzPYiJshlG98tIaH1bZRfZcBi2tE4GM32KzYsjM21hhdUh
kOQlzgKqEt0lpOuJGBWqOA5y537iJUMBjdZbSNgVWUYrQQfd/OJ/r0VsvZAsAytIl4ZgHB3JHnSo
LilKrRTlipDzF2GjAcFZA75LIY3SxkUDBY1yGMzc5FdJgqDEJ3oHK01YNantwEc4mW4Hf8Oe9OdC
+Pf26K/gfEtYU//Sb1Z0vloi9tsFlulC+EmvXB7oHMRoMTdK2Mmg8KJ7qhEtKdaRowyCV0OKQHtC
Q2x6LCqTUwdsqvRFNt9JHhWJGhY7l//DJK284//kBwSs7wvM13dzPpnpWzJ2kt9yWUhvQ+P1Y23M
NTWzThMafBnlX88UdT0GRbTGU0UVHMopGj/kMIkmOjIIF7YBl1ezIxGgo8dZcGGqSs8+JgUSPW0u
dx4cyKhd7JNQVHK3rijLj7cySX8dbk9db00HR78HDwr4IV0yVREvpphq5ywCHrB2UJ0X+CXK6UbZ
5Njc1thQ1ZV6nsGtMShxmVCN+IJ3HshLCyyTvOilppYccPwp0V2dvafEcZXgHriVwSpx2lNosdm/
6600JeZPR1s6uNuRJKqPBD5VffvO6g5CwLYtDiUiOTKwGNvAiLJO4WhujeGdltC9wQGbnohswUhi
oMhme8qtA38si14xIJBsKAB16iX7lKvdPpmJCPpdytI21LXjgVAv4cOM6UafrAhOtyEsjLeBvBRe
R2nZNFVXCrv7SCeyOqgtWYIMNQMfWgBRwiVjF9kfoWrdKOYH+A/k8RoVMyi2uf0vV/Nm9seNL2Pw
ZjBhVVmOZN05BwIj1lx0Vs2WqtGY8jqiX+utNJGlcta4Ia3b8oZtHiJ5E1lez13KkeLYt83c2CrQ
rB+QZVizNQSgWdSEWC02A6MXYw1dfniK5+jCFlU0/mtWjgDKQGuVpariRiAiHrpSZP+aVb73d8Q9
Z3v9P2Xu3mJDPyFnrByGcpyHNQ26PUXv23wvDFD9jtpOPFk99lT5FsuSpjezMdyNqFN3ht81ywIP
HXuMD/2RNyLkxr1DpHh8iswSeCq7NIisrKjqu8AHwL9zsVskMci8K7FpBxlrHqsAor6R27zkRkIj
OFSt6eQJPnxAWiTrt725Rg80AxP0AEtacWei3ycvXvrPEoT3OEVd+aaGQtE6nCpXye6eq3/OaZV/
UfXLwU5bZvMOv3MTz3K2d+ZxzSDRDrwhyBeNd/EN07Kh1xYC9TE/CXuIndraVxavl+EvbGHUkrwo
jFYAzahCoifLo2qF1WGAVbrNtJFNM3rm0mF2dUBzoHkw2jUNPvhnndw8oBBNxGR3mbGzGcZ89Dk5
YbPqp/buj3/DSUrIUPyPqoVdFH0G6caXQ6BpQfQR0wK2jDd00bgZ/9pCl26PdGUikoqp2n2i/OaF
J437H4BApGnJMsYlYI7HHxnS9bRmV4KOZUZcqKJH2k4/cnff5BGXjJ9PTnP1DWZ2XAOc73q+xqRr
PI+9Og7RTaKrEXJVkXYTCccCrOggbS4aKAWhjIlY33xm3pK8AlQ2E0K24Yy+9eIcv85gflFw3pms
biKDHZaXnNw5dPbd10l+15bFkXDyKICdTq/3f7oYMf85oJTb5AXvH3U2d4rWvsFsif26Ume+QQHH
5qOAx+oraByWsTwJnyWU/zj+nUtJAIRv+wP1aMHPli0Ea/YCCLwxwuWsntVFgiK5rKaNmN3IpKFb
1IGxxg6pyFU73bDqTa55jD76AetLbIPjQFZ1fER0FAjxSEE7q0osO/oGa3AqP5xBnoQZEGNvsfR1
8/fyILyg4x9t8oIHVDzPmC55vuZGUsJ+3gdyVmOeuyLrToXImmSIdALGLd4Pse7vDmmY4d7yb97W
DmMxcRTFAexLaITVFdSFQmt3H5zPFyrELQZ5yB46s2TdUQ/bV55RZUQWYUPgZ5zvV+fHsqa+brnX
ka/GUfF5AaY/7cbiPSvv9f3rP9a2jYmqqGh/1zMploi3o75ZXnlvV4CEnOi7hSA+oEn2XJJk3zF9
bi00yiLoa37/w5co/YMcELr1kUH6kjlxHMfmznCuscoOaAMltC0eVKXWdydZxg/KB5q/zrFDIfQd
1KpN0T5xozEqierm+xIJrz1EKkuwOhhe9TdWU7s7+sXQWLetwVZp53Dp6d9pxv2XUT+sYcXCIDMP
XAFz7Bg2NqHGYWKbuB0oYyhnf8kjqpLVSUw4/oyB653c3NB5UtOGXCfMYzjZfhG+w/BjSIsRHD1+
L4L4jSYurDFxDIgODlp/KHy/wnoXpDirEm0qLBHGgouH0ClHbXwzWR+JjSoMBUXCY/gvk/OgTDo0
j7cdjL+TauIVTdDbUFDZfgr9vRYv3AFdNQApV5X/Cw7+X8YWcfcC4R7LrLh5daoKFBLkV12ppDuM
k8Zpe1gPo7Cg+gVutFpMaG+BEwHhvgcpA5c+Kxo+5dTnKObAezEqPbwQCYM2Hs/aBC6a5U11Iurq
FHe1x0waEBhGJ0qNsMT1e5958w4Pu2z5Bwfhla2xL1Um4KYb3nsvCUwm4Hfl6euJr2j0Dz9w0LMM
JI9XrJo8pyHJ9mo51R4BlvvNmrg1W0HFgZ11H8KewotrFme7jWigwVbP/un/aFU2N2UnJf7RqSZC
XPt2yDGQ6F8yWIL79StdiRaEeszs3AQoS/OurDUEzOhuabOpW9g2E94Su7PQ01+C1DkMe6ZAquGE
AEH/ztKkBgiX9uAz6iTaMTx34HiNIj2HeXlJMB/mfxE98hEVTT1gD+Z5fu04a2KqnW+urxsTLD5p
eUUm86nq5MqjhDo7dICCWX/bQaG258RxgAOiTqf/tq71W4T05iOukoubLOMwoFRE1rmsbrqgfWJD
K1g17PXndaeED3g4Vll/34UNsd33vxfTFV67j8C044D5rsqDYA+LyW1q36QbUK1Fj0/RmgI0wXLr
SMeRCtskqtsH6Z7C8iHNiEr+iJai/21492UCax6MS6zIBOJsCqeJnxBo7X7rUSW3k8I3iehX5mAj
h+HKYREusuujM6NxIu5xb7wG2GoWS+tQaPGgzvL5OiMWQcfuW/n5rsnKoNruwSqCx3NWHdEyFTdT
Jrrph7wW8wV6mOnsr3QkUcF+RSiZS5xlUsxSvcbfSIhvBlAmW2FUz2crygaeiZJl1rnA3b0tfRwh
NzA0vgO7qTWxhEBkKUiDxEB6abPER4rM6O7s7x4l5v92j382HXra6Lp8OkPHbiSBd/bE/Mr2N/f6
bF58MCBG51Fs+OKmIlcbCwYo0eLlsiyAP3nZuK7NQK8ePCU51GD7cMCa6I4MISdSze9k1HfNK9IE
rCQgzC38KHgnLR1y+v+S7FN9G+Y3tOv3Y6jGxid4VTlhtTRlLh7FAo6UjW0JHUtVv6GgcwATdRLd
wzbeg6/iKhOepoWBuhs/RQsRksIKfEMUFGdJ0SCNCEDvFd/ZpeuLQ75OrlF4s44wFKrubYC9YkOb
3W93Rcgk5y4QOxQk+S3TuyjBSgQ4XKUme/3n5hWSXTFXTMP50beOEG3an/aMM16KYytcF5dd7hWF
1qIAJrJZDBy7dEDYfENod/JpnLix1/5drUd963cKWmHaITX9/8cUgVWj0Pl+YUiKHL+294vX9B/R
6FpXZ/joO9paGaTU05NINEvzqhQZwfPG7QUYL8+7+lSJ/NUpZ6MCXY2M7j2LUyEO0Ic+39zY+coe
XY9xhvWSpK0/Az0MRLgE4eDCBFwMgLS+XUWLgC8COqF+EmS0M4GFbA/nIHV5cpCdSYCd/psGA8n/
GKVyhLnYZPslZrvqvHYW32gUXYaWYrZJuZvTfK6ai26A7nk1HAPIGq2P67/eFmdUzkAvPMtxxb4h
/xEiN2lw+2OmI/8D7bQ/61vkl3FvCYlmHLcQpMfrytyfAoEbMWY/3kL6xbugPX04QdNTe3HGi2a4
LrKSf8lE7tZ+FV3MgOs7xMZjJVuPp5AQtbOtia0aWSUyk3++66wQjkOyvqs5xUl5W3xwxNcpkwiM
bVTbu/ma8rQQ5ODTcfZEsWvbAZm8FMsw6uN154bPHmQPvZt1G/eFEP6H0VUxD+g+p7BKlYhNrbZr
BAKdFHJF5t9lY7nAqL5xF6mbyC4iQAnzT+/BrSv+Rluh8ltwrHDFD2mwO1117IyjFON6S+1jqYGg
p+zNAsLLWGJq60fMOZNiD3zEKD96xRxS/C0tOnsMk3c4htZik/N4r0srecSGb9TUJRLy5LYZmtAp
HsFXVjmhQrn6fypmqPE5VMWxHRziPGaDFYVxyPIUzDx506FegUNcB4jX7vtrnyrGxzMRRNhBUzOb
12YvyJupbmKFiQ+NalDylIEJtdxRmz9+cruZughTt1howaB+7+S5IvMqAxiT5odDLeu31U30myuu
Uu4rE4hX81JFswnjfGHxuoZbjfQagJD9gUB5NQHEMvTL73NQwU+80muQjTA4pWro9o/bW+l3Wc/a
f9Ej9jCX3JTFWqpbAamrGsurVAIs49TXvxW9W3JRMFQ4Ai+rO491GSiTR50x1/YFC+cq0ec1r5y1
K+S/MCbKFJWM1YjWYKxAhxJ5fkvlVfZCUuSSSEYc92dpKb1kZDOG0hxc8TQ3bap/4IRsXWbhCbCe
13lCX0XrYvjesEI7SKpaHDGFWAoezzOVz4gnXaj871ysqoPielj6sVIs/1Ruj4onLgd6VYxpT8nK
gG48djauPyPlVbuAzQG1/K6K+H3URqjBPp532I9oldGpXcZU9/nOS9VByOGjL2jUjpWnALbOMhUx
0udr/pdzo0Z+zfd1MsFCFRe6OOV/NUG3cQLTen103lm9WCJ+784ULV301MHwZUXgvYAUu4ON5lx7
RM7RUt55zslo+tXK2ksZh9Sk3NbYcjmSnBsVSWyjhpkNhL0PxR8Tqk31qSikUcLoCQY3vdW4cKVb
scKehxLCswbgob3RWnkT3BGm4UpVvmdx5geizUqtK6oZyds4urEhIBsnbLTRA3McTd0ag51fF5En
O8z+oPqyzW2O8gRJnx8jtYjFgK6fc1W8Zw98a1+8vvUgL1qODsXwgeqfn746VXhIZA4gHQ3gfeTN
zqSASrEn7t2VXCCNC7sQBu0y1IwSyjF0U7Skta77Pwx+DjEEOD04cSVBCvuM+BosG2TfiZr40ksD
ClXT7UYvAdQfVg3MVjQ8Q4OhrWDBBB9npffWLNwpQlus6fne2ukhjUkrcFRMj0sNMhJu07iZ3P+D
jgLXuvyBnkeK2ffFj4DKZeY177m8DpqdOL/7qPLDrgLMYkQ0XYOnTbTuXmkUbESqp6Ka062qpDQD
00V7wobVB0mWVGel/cSuOlYGcC4XzqZ25qTiQlzyLLUoaWlaebvnOQbBgof3fZvsPODUyKBH/pBY
9GvjK1ucVUZaGcO0pkgFBo2Dooibg8jL6y+Wj1R+wGpLQp84GVabwIRCUgh3bCcW4iSyaA07lhMU
aMzBCw/zrV+ahQV+z1zBHpDc6CL4CDm3DyivmEF33wF3tj0iL+YxRibhQQ5hZU87DwLkHj4olGMg
uSBoTKJ7BRut85ZRbeX5NFUenvQWlhBw1Co0czra8f0I7iX16cCTCfeo8WyZO6ESJr/1lab6q7zh
lNQ4mDUNt4vDUErr3pWiiSNYQcIb5BoP80PcLLCw0CzpHKxpfq8+kUTD87GtLR2CGz1enCd3kwXs
YZvHcBeYbIg3JAzli6d4ymgMDmXbNCUqZqpRItoc8/PAZUNCzXgLZQ+D5a9cPliLExvSLB1Fwctd
jkyOjPfRcuCmIZQtVXnNkDluvMs6E+sKfGub6B90ItN5BbzT4KL+6z2tKJSkgmcikXSkBPcCQp1x
Gjpx+RC4pf5LkAAWM2T+5AD1TahYMuJc3QBI/t8t3u3OQf5YvVllOLgSIegcK0Xqt/sU6X1hci0n
N2K3FVhm9Efvme7AeHhGDMn65ruGPJDS0T9i8fsdDCl7mzo0kbPrQCbLufwsmhBp/7iGbOCPrkU5
6SF8KnVE86l1rhYoHAeEHuYci/YzXNq7RYSLIrR8Oh25Y+o7rPHkrwkdyqty11QhqNUQx9WSfCmF
r2Tbd7cwEksF+2JAgqlOpM46VL9eJVic0aMV7Ap3oaTzVQO8Ci3qY0322z9B23NkjFCRSX66Ws3W
ptduTtMabZjn2rR5uN6HvMgNdrWH6wGS172Yp9rJFqjTYDjvlsr4JVDIKWFwRh0OvVrGgK5xdLwx
j0Dt19YP3YRdRmsBrM0W5pnFb/XeJlkYfpTS/1DPvUZQZRXFE18ladO5fOloRWS50Jr5b1mefAer
GGBBdKEudHVhMoZ67hqcAUgSsqXyWebgdVrokv1D52uTFQVEUSDI2CQlH8JlyOzyzhqKhghiYVhW
SQsloREcRzb6qAb8W+0HuUS7/NJJPtZ1R71NZ5xM7Np2Oo7xHqpKHHWg4KmQTcZxACYlW29ZsKVu
Otmr551DHnKuT++eQ0SAH99OxjKBTUi1/SMY9diw3igFK06SlE4xzx/QSyAQMNWZhAsF85mCt3xt
SL3PIFczNa1L/+9HqA9JhloUue8SPJvjucw/aAU626VT8xYl4OYldXjwlqqsDhU5Chekw6zK29Xo
n4A+ui9LV62jwqw01hLJwIBdwBMgsXc/FETm2EeoDN2ma2amv77Pmj7fIyIyHHvHgbC/M4gTsXT8
I4PKlsTE2VKtbrPwaly9RE2JSpjWW57gaWOI+lY8pxdmAMgCjz3h753IUEk3f/FHofAZgKuewSXh
itLYSYBXl6EP5RnoUoFIe85s0XMubSiufVH0GQ69FT8V4uyBDEyHqu7cihh95MxYIxFIUlS4oZH7
T7hiT4NG399U6A7dHc4PqX35PCMglnK5f32jBH6F0h0RUcIxJCD4gpa7uKeL4nxB/+JqsKa6ZRvT
rW7gEy/+ggEv48jhNBQAaERAwe48n2sdty4RVep19QSq5DYTi+pla6WXBQ+r4xTedvZpMKur773e
aeILDeebZmQyXrXpsiZgiaEH6vtVFI85JCqpoU5UtCfqerkAVfNVCYrvuJnFSXOkxkPm1Z6aIJOI
ociG4G4MPdZLHeveXKu5Doa3VS5I8nwKiQ0MpILiXxZFvu+OSY8DCeUDzUXCLcpEQBcqdElp3eGT
4zXba5zjvMQLspOx3iwmi08uU8De0JkSKf54/+VksO60QCIFujjyIoyRSVexIQzpv085jbnKkb2D
MUAhr2lr4VcaA1Yb7wyJxo4RoTw83e3xRTussoj7wboZ6yu1KmsFVCp+gPbvJ4CwztffFD6apuky
Qc83QxanD77WTmcV5HhofxrnYqmRTBSeFT+t3bfrAVM+oa+ACiBoIGOWM+REIbf/gS2Fo2F5m1LS
9rxbBtXBKnlYdlJvpxWnjeZpE2NSc0D3oPmw8xMUE9slOAVaZU6RZf/uMpGRjWfpzeB7ZcowNI8H
SiEvI8sfRIwvpSVni9l43/a2wYbMAdzQ/Pv9Fkxf6g+h0bfiBTVzaD1Rj7kBW5BFGPMXq+MQlXoT
GfPjtkLvQCOpOtnkZQ7w3yBRi9lKhIRa6tJEUbm0pkB+QlByQJ8EqgY8dMA8pxPsgIbcVo8xzLJb
mSJ+OfWbPcDR5eJis6s+OP6xx81C3FylfP8Dr/YsWy4JINBy1BNwMlLjA8kE10zGS55A3Rqxba/v
0KDpgNEcr1mF8+Hlhx9fV1hRwX+JJNkSrGbKfUA9ZtIQv1niYHjzRTee78qi5G18yjsBmkb72Eyy
o51Uayxe8cb0d0SGw54kSRriI267On0/pgrzONyW6bgb5Srff4K+j9mLfoeO13v/919Bh9I9zle/
Ud0h11YH3yzVNeZ6X/o5PweerEw8kjDGfhuTUjQGNpOF62/kP0ZTzLcShsg68m7E+8S8nbTJBsAl
blk1SOLduJMZue9Rf27OBkjW45r6+jh9wbzW1GNpk54vodyhBxh1UMvat/WqLhp532lPtDzfjEko
TQi//FerfcR+U4SauZDPLJtQJpGKjIpqvCSS8wtOiYlk0c8IaWEzJVHytiAPj/xOIXozer5e5pXQ
0vLfweU/5hjY1+sZ1un3alwxOAfadwml7FXXgPuwcoz8altbUq6ye1zmbQVAD2IoZS1xRDQe86Iv
yUmgYqlBpIR+Ay56dnC0PzBmLIYtKy4jd+x4aYAHl/ur8Jft7DohveatT/6t02CNxETj4gH3EBL/
ZUT5yeM7WkLTMO2C8XAZccIAFZTbzOMi654gpk0Hlr57bX4TF7Gi+WqKEJqHX8+e2UvDYi3gPF5q
/bEGARatNNVhTqGG+tPRgJ8H899TKiyei7m68QK60g2zHS951zXXLP0GjOE/+QbOr8T3jbGfxvt8
LSvkO0E8Ip2wMWFv+bvv5x3Z+qXodkHj6uGLH8ZbkqCdcp+Coyx6qywJhandGyYJSeZy93GLKxDx
BZcvtC5ztHPEiX/Pt3zoG7nL9CwRhbaa6QiGbE+2xMRjTlOGfSarEmxkQRKkp0eB1JgBn8b1GdP6
u97hLY2rl1YQmcL6j7680737LQqdVKJQwCiMIIbCBy8t+nmB/WOd4e9ETVw8llVzgyuebQWGZ4Og
2Y4ESuQP4CMiP0F+vOECwHi+f1yxjS5f1mcWjQeaDzS5KfNnWCxUTWTLX0OI3HRRS9onkahD0cRP
sbgVHf0uixhXXUo+J4QhFd8qx/jIkWWc7aym3GC743JYxE7zVK3161esnfbw30EYqIhrn+gk/s0c
Yorbq96GxmcSwkMaCprhcqb9pjKvUd/gFNfOAYXtQacuJLnIshXEhDnb9BZn9g4NMkS/0omeYAe0
wPSdKBKOZYLW/eEPGfs0gZOvcpl8JFy4ji78zPaIr0x9ect/cHXmcMg1tMBujY8ae3gnxya28zkh
SMUbs6oFEYSFOc2IYTwEucYPpgrTSte+bih6w4IA227fRssb4GIn5onBquXW+J8MfRws1op2ApNE
22K4qgRglD2FZapjoL+3b7mK3N351h10O0Kt2DIPWMD/S6Eb09vsxFCfVq9RQ1PXUsdwY32NekAa
aEJCMPPEv4awndzCaQYAjwjO2q2taht3OKOJQv9pD6lIBOYJ76mUg0pu6veQrzNnoxk+KyqOSliF
z1CZyHx6pxmUUbwVi9IhgBM94cEYH85g1q7i2OOxmrCGdnilH/2o+pP3UYyzvLlHXosYSjUXrF9g
aWfIDEzXam4AeyDOKRnJiCt1SNTSDTxClW9hBD028qkMOjPnq7GjgwdSA9/j8ZAldCLmYXdvDKHZ
1N0pNYAVSIlSXG5Pea/lH9FggahvRbmGoY4Tr3wDmxzsvohfTDU0jgxdJs0mp6VoEMaXid2whOPz
NUNDcEEvVaPYKQxd0gDDI4VeeGW431i3hyZBHXWgkj+zUIq2xMOpqNbBeyxuEXp5HJrLbL9OUBGP
REOryXasc7+gIdmGtvvspGvOMdlijAeZjnyLHkkmfgwCY5R4iNwHuPflklKTFNVIXBIRSswqnw3B
rgSY89vIuzcbyZhnWd6jx/v2NgUROr6gxSLpfgYjRWfEtyGhZVp+YcuphvpKXcRBDx+EoKobJjZy
6FfYa73G8GNH3vbBoVhANi3cKRg+7YB99DSUSTLDbXYAP5zNccEjJaLsPZKYhciTtbavWNDiHeHd
PMN4+IAIzDnoaRTWbpD+ZPaqKPknX8qa2t35d+Vk81BskyMh5ONqx5SYJFWPDfcuOej6fpIVaRxI
43i0aEzMLhpc8Hsj7hGKhd1ekx2P5aKPN+cV0443zWt1ge/+XqLs1hRXN2XShNKvb2fokZsXp+H9
CIMfihiXDiV0BQPlXyemvRxJl9TeMiRApx4O79Q8lxMr5lV7ya8En3mH7i51sdgkrVaC8A5UKqKp
kvWPQgPxTN7nx6QvfOvCf1xGqYhU9wkmPtJllQ/FH8gYfT6SQVz6wkRV2KvV0LPwQYMxtFaHTic2
AqRhoHPz8DitrxgrX0p9nBgEGPuqjYsrO0yTmTfk4HI7lJ/pe9yuzz+5F4m5x86sfEGlHUgGb6KG
ilmnBhxOhpyQxHQxg9l4W132bROrER1g9ZjEdhzVpIvoTbqvpDSfHcH/RDQdy446ata2xQsu/kJI
pIc19dCY0IN7TC1z9egYGscbjHXFH+bst3+CLkgJ6eUT23XNdVfn1bkHWiosokkiXG+Zn+sZBchK
RL3u0RWoJMFejq2DNq4HWxLp0rXQ2Cz8terk5H3SrdvyHBxs5Tw8qw28fCB/A6w0kDOMDOHDoBJ2
G+ntJttVSrX6BS2t8WJEPWXOkH8yK/dimbjO2upCS9AxKi3HeWKU3pSB/Clj+/7l+2LPD1vvdy7S
+rsongQiUtN7HOvd7qDTZg+sERiIsiA0k985IGnRIbH5hKLNKL2x/MTSh58yUIP6DNhndgCO8djE
3aPeGGHZrtjk+Uqy1OCVY/Q7dYDJpVmhnLwxaThPuKIIZWDuiH0cJqOPtexMEXKo6L2Qw1Oxc4Vf
fdJ3hx9iEq8W38wnxLWuhwQrAIMhyUTuMUof+Qkz9wWuBZTooXQ1V4yS13vmV+x5RrBoudrxEDg7
1HQ+tym/ERLLhGnczlybWT7rpNT60gl2IwMP5E2ZHb/5ndBeRj9VVuKE6Zd0FClMPpBPv9zFBV3c
ZiQYgEnliu2GJyrhxYlh4gy87s/vqdm5ymsFseao1A3e5RpdKtVxAEA9qQSdozhTqwBjASrvs0+k
ldmerxwlOtH606dIOoP0cRabxn76kp/jX6Qy1C3oO7dYmtH6DMCGFjwFQkEDEILlHBkVHvH+YURe
JYTCf7pzItkUQiNaprBy/Y5NvkahO04QLsNGTLUg8bSxjslNkQMxf4b/Ayqxpi4rqBJwxDAkOW2C
W/XvP0IG7J6d8c7BYJDtxVAkmFSMNr475vPGsyeOnaCnDkCfYcXTvnJpluJ0HkZ+y83+84jjkJJG
Fcmd1Qr7t5hXd+R1Hapz3UKvCS1tFTbGHRy+c1P7c1FQgRUJlV4/r/swZ+qhZi3pMwPGOCOcPBBl
PUmdvGKsUtGRgO4a9lwEwhjzci9gKMIw2oVb7ORqIYjUUHeE+7xxe0+aoJamfpwrAq2wD77xDrSh
Nq+6qbaWKUgeJIQKXfD7uyAf0bMMRpGxdfCLX84sbK2BlWB3NkAqOJUX4leDdLsaYLH7oaGWq8m2
m//Bb6yYF7R0IdWektH5X1wGHN0R7xXmi5WjYNMXT8mfi+DuHYAKhuE91/qDgK8dcKpH6SiZ6M3c
Cg7vIwZEWY+12+4j/U5IGdUmZeUecdFcbDcFvKIQ+dLe8Ylljbo1vpiG1StC6XZVIll2X557d4/Y
LZiw3am6BvcfAwy7Nfb7UBqVMTB1dp6yfB+mQzhGBT4C9VPUpZgf0BirW0Bm8z9bBnfCb3V+CEmb
0VdMebZ1NR1mb/nhaYwWNarsEe9rSvvznAmI7mBxQUk8Y2s7SvkIK/b61SxofkB9ScO5Ro7RF77F
1ZbcpnilKrhqN4p+aosMt+UDHfvSdkIT84IGZQ8/JYggxazNjmLygEXtN9ZLraBK9hn92P5TsUiq
A5wXygC8pWoWbqOCGA9ollrtNEVLq2HYwdrFQXF90pAQN3eZsos0MF6U9zNCVK0XYAHr0Jke8J5u
dly+NCfmr/ogvTjaT9NgG2ujFKdhT8WWMLDsjPvCyVDQnh2cGlz5ueQwEU3nQ+wmuxltVSIrJpPq
bCepkP9ICpwTrKb9330eApyvAFERd7XJgF1ri5mWHaLwk1c4cQ2u8Yp5DEM5FL5b5MPDfswd/QeI
toiBKSpWMSVPT3myEA42Yv4vmJOFs8lWFGUV89EHoT84BqLb0uLQUYwY6kuAPHcFn1P8ApNzXpWN
VsOwnkkLayh4PCnlH6l3BAQhdOxLui7quoYka//bTjnmXhCv59E8Zc+wLtb+VdSN7ey1WrWUKetx
7rmuzL6uBzEmUcTHNijVUenpF/ll73hvBMXuinALa+wld3eNw5YDFmRHMDfzOkOjKsEofoswvXip
Sr2j6mTsv5abAkD4kZut0ZGyrigi5ABVuv7AQrb2uj8XXhxe5sGYpvlLJVXmr1eiECzGIuYjrY6a
cX0/HnysmqCLwDzKXmwkkPId20hTcy3iRtY7MRr8SjRPKspX6xZU5CvyQ06RFYTqCnLURngmeu4c
yO5pg6IbCVPWXWsljlfE6rJ5u7u57dA//EyEdXkcn7qBnPjew8hyIpqFTJxaO37t8I5gRCS+mje9
h+XeEgqQJz7IoLu88h8cLgArXcoXOvQ48ItTxxI2dtBqtb2XxLofdj8u3cMqZiThIxwEBYR8PW59
Mt0e1DaK2KNpcqSU9Oy6Wo3mokBqm7aR8TlLTYDS4zfy98nfII538nrwIxEj8Q6y+aF8rUm6+fpH
PeG8Zh0LKmnLaAMrr5boYeupcox2DnvGpBaZLpQ1/F4KFnPUvxNAiVcgFTNcrCsO5fEjfSsWSkbW
j+EJgbOeDWPxdGWk5HpcaZ8u4p5WsPaYbfvV4hSppZEWW1VUtdTHnzcOOaBvIxyRhsmyqoDiFq8c
EWDN6s13SwPX7LsMh3XRH7g/BVPiQOP1rw8vgojfR/Y6MqKhd2iibUExFxx258/Fk20VFzors2za
L/2jKboBrrToXDY0IaT6jSQeR/nSTeXS9bvTPN+kP26RwTi9O/2bDbhMOTPWgkIN8JtMuTtI6bcZ
f5z9lLjWMP1CMJe5yURi3KggOqUeaxJTnQrGdkyTvBAlLfW145ZDKvw5g2lyO76pkHtEU8I1kAlZ
K+CqD1FK2ak7kEFeAhjMrnpBZsaHLRY5JjoZvhd2284/Uc037cviuylrF+34ZqPXpyE2GGfDkkjt
0e1z/OzosS0FuCJj2AAkfzmTbUIBlNauEs3zx4qHCLAtK5aeKrxHGbId/kzmdnwciydjVp2Kmn4Q
OM/tQStxxR36XqYTBfnQVC/whiGL2g/nY91w1dDjeKN1U/o58yghl2SQQZWXy5ACApQhWmCrEcZ7
o5hzS0DXr1C2imog9fRZs67FJSt0YJER0rLX4pGntbtpBEMOj3/YJxRO+BZtrJM6It8DLN7EItth
Ose+3Sw11oR928Ym+sQQ3OgKg+CBT1tgNH7xSPZoGQjCezadX5UoE/Uien//qXrGwoFztd6/se2n
QgKW6gJiGYTdWMO3gMhpnSf3ynZ/Bzc+gHkdtRmXMZqx3uYRINJwJTeUsEbrqxrXUL9UgvCNwtJv
VsWDwphOBcdqSCMDJHQQM2K0ldyz4rdqJrxlil5hNJ+Qpyu7AsfFtdfHwmkog/AiM8zjZU1q97JH
zHHRFHP+/lNal/HIVsIEOFoh13vUdtP5wZE2Dve56r5lyR5Kkd2ozuxahS+ozaiFZD96O6GR+Hc2
CF3Nhl8NjdtsnzRdCdkC/JUBtxq0Unq/yTjgP4mz3tfuQWrVXg858MVms8C8pf4JFs84mgIB4WKK
wfVq/DaFnkmspIQLphT7DGtHWRoDNYkS1k/5RxY/zl4tdRJcaJ0lrZGeAH1aIqRgHHoPZbXNKaO8
L7ZbzxTUbNCqAcATpZqLnA+vuPJBWN0VsoUQCzrzk00HJpx1I3Q+VMPI47bt73561FFs2i7qpMWu
Zu3lFeh19VRlz9QvRI4ptcGcD2txx8lm14MArDd+awJaHDuAOqvcXANFtvAs/ljJ+Wu1GhdjEZdt
53B5+0zaNox8tew7AogXQFiPuA9hO1azNTnKFb7xY1l9IV9GcFX3oRQCQRXm2w916Knmj7/Bo7X+
kycInMFxI05gbJJVaGCuI/4QDFZ+3+wKdu82C3lwrUjlAIMshMG2hQc9CiiV+PbcyxeCotZYHmwe
IExzm+SXAsd3ug1Dv+WtSEV5KTGlVAvB1C/fY8PKIpvdIltxme7d3HaGr193Bpj3JXIFlpeJzK+R
kO8e50C7lpqQfW9VQNbeCPsfAID71UhwqEeW4K2OUh7at3IFVZk+9cxI2zsjNfskDvvtrkH3sFGA
kv9fSKaE9VzfZFpilPeAEeNUKvk8csV246V6yE3LrZwoq1o5/UfGSzzTd+9spwUOR9gQX96BENFH
rBzwr/Qekxhv0096cFhVlIczKX02wU2tdgKR0KrI2AM70T1bbb7wB2PmGgHn5gKrGRJmiTKyOpNP
phHDGmROmqtOlZLcJMRGSC5fYFFJHz15Lpr8iGWOy7kq5xoI2Qfza0mEFvjfPIzJgRa5sMU/VTn2
udbwb0dU24UDV2HEAj/nmnLmpw3qhpvVNKhAa07IOqIpXo3Go6X++dlgwhdRCo63WeaQlT4yMA03
gg74kbg0Fqu9jrz909yHNFdCAphDDh6LiaqOFgo5IhnfZSnB1dO7Q5Td828mUHNOz5M0EXBuTFFe
5rJZzQ1G5WbV5rPPrf61bD6x37JN0W/dGa6djixfTuR7+0TbWRydh3aRJIqWYQRfYVnf4ebRBCEY
BGyXvgiUQAbScKuqT3MxEx5NQSGX7hZfgHJzFaPOVW0GPoRhDjknq1VrwY0FhmwDXGz6zbETFeyk
Pw7u2LWjVaek7hNAa5mI6QoS0zsAmaMb5D9BQPHBAiNuKEgFmh7vNEhMj0YpGIuTTI6sqQj75Gzl
0l8uL0I7Y+r1TpvpnkREZDj/JqglqAq+l4pfmPk/0bQznoBa6Q0KKRZfJCFJ1yibKgrdVrJ3tA8i
lZcCMBr1PQDEkdfwMeURLc7yJSx7wZRdzbW4tsyCJ5bJSWgZVQQ8r4dhZAb41M6/SI+1eZ57qhzH
eN7+uRItQ4RBeIoGROi3iNJmc4nCqD6jKLN/2CaSmVOJI6G5GyvGOI3SR/3T3KkKRyCVgmu0aMnv
bPsEeHHXzNTEarg3crUKzJAiNvf4hUppmjh7vraYgqehRQCY4Vsa41yt7PuywLphYuUFdcksbIOi
dp1MtZIqwnVYIqLSHwfmrQqIA/8JP50xqszzEEJg/wofRuWg/wq2mPQl8EfMKzKrJlqJkvSbx1vf
XfbQ2QjQBHwanjXoMRnRyPgsFuTiZG24gfiIxNIq4fqZ+S9eT1neSp2WubGt6lVpWGI17flRH0sw
STktY8WyJ2HB0iiX56Hd2Hlfdir///Z/rOf9tpTVwQeqzfvsZ6iLZrEGkQzeABY8SO88gH7JfBQK
CULQtP0jK2E/yv2Umom2qtiboK9/NVbOudf/mfkaFXO817gSC4q5OoYyCzX4lJE97RFfpZ2+Vuop
Dc0kN9sLYmnYGFSjEqyvaM8bZlhKjg32tjwk0HNrfBnqBZokp+EuwdKc1xbdvTYS0DxdtxdCceey
Hvlt6pF5OVGHQDE8zeoPHTwguaBW1wh1xLfxbYi93k0cW4B/Zxuk19Vf4/bQA3QTZQFhU/LkRpLm
8b4qc2vwKfvvtlova94qcqSbj7h2WGV7GXH2QGElo8Y0ysXRCoBMZjhoO9sZbLShKaNCnCpj+OC7
756sEOFIz9cGO3cyuoydLX5clzBZa9aoyS7QXZl57QV6lrOZ3xYA0UxmhRlBAFG1f9vjLygkNNtF
qglxA1GzK0Pk6Up4b2i65zNdRaoKxt7GRt1YLgsqzYTBVHhyz993zXNrJpuah6fQscUhdBiuG99a
tqEfKhT219OT6CSM54cD5Cjvmnei4faGcLoSJDOAzlzha4Crb6RG+MtBSN/BzS9O1CmKoE2kER0C
8EGh7phhZs/R0WpuSS0EZVfoH7IPYaRpjTV2OC9LQ9APBiTfL+DHYPJnAdHV4R/Qt0bEF8wSGyw+
b0i/9q4B+fx1IdmBiQIyBx+lcXcpGJYtNZwzb8+KHS0YDbZyh55nb+AoSge4n2GLhgSpSf+tPUUQ
O8+qkjS0LIOJl/l/m9FywuwL0yq9cAeM0orRq1Y/dLibgSWxaaCFcu9Lb/JcVDArfZ4BF32JmrUQ
bU39+43KpN9kTJgpJGhhLH0hjdK/ENIEEIp+Ai4GTIOdKtIW9GEuBk50ZP9fOFDv0zABEN8K3uoM
84CO4VfjWaYP07OdRMarGarUkFX1J72c76La7Y/PuX1FANmrLOJkEZ/J3bf1g4AZkhp9sq9kvcy4
bMnS3//TBFls8KuxPHqdu0cYACWMoaLUw0DnIGuNx6DlWC6EuB+rn55MGRg9IbZinYrrMB78eznw
UcqYUHaed9GBeBqrP8cTP2GdrIBdUpjlH12yrVzmT8XUuMfNcPapEFNU98fJPZZ5TkVfup5BVodL
Q7NJCpFv7vA62oRLwKfe4yDqtAk9n1sFtFzvwG4Wt8E1hc4xix2BSZJhbAThipQChL5woA1n9II+
/HAI7L6+bO8P9ONXmQxuGuRzUELa7xh/LDIAdwub3OsIOvHd5p08+FWNBAC7KsYDGap0lowU5sf0
cIo0ShmhFD2cA2xNpRCmN5ncq7tYpGiqDSFyXFT+ux+rbzi6oPd1mnTgf/Wrkaya6KfyL3Z0WsZQ
a5KrQTB9VEB95/1JKcZpP6u0ksLjWQ3DC8ujUfGlmxNYgVdHurnbf7/WhFJNjnmNhD2VrtGcYXDE
/iEepLLeGhnbz5bpysI4g4KFPgQqZMc5Yjw+qdTB4ydqY560R/uyoZqx2ZTnbWZaCP4/DYsSS4Yb
QHK09jcJMgEugbnHcdnRvDF/Mw+0nkiCAU4sxLMzlTCVhqw3jCjo63pfOkJ9KSYvXfO0JG+quPae
iCt6MNgnWwAUNsKnBxn6S0GtsYkb+OkMXMcL2UByNI/YInx8f/fsvDVAQokbpcL2K6av2GpbxR/Q
cuYeVD5HPd51YcNVc5LTOsUv7+O7bBdMMLPrx96r5AFS1m1oqHjKHeZhrDgKB4XKITkRRI/6WT6j
Hz8lzWVQCOnZZWhB1kjPfsFGPO0Pj104gglkw07oRr+lBXeL1jh6+ieUONMXmy4ihCqtHCwoj7VF
9o43ehSV1oGZjjZ1HDL1Aa1QcJysaXMKwh1j5s1gKTV4eEIpqtL+DTeSdbPArdDg1AJpQMYMhpD2
8cDdups8k7rQmcO/G5cNq6TqK4BXFO5YJbR3N5CqKIGg2+6ne26j4dm9/wiTwA7FQ3cF8j/Hmre4
A9dqaIAxNd9GAbD4hCGJh3xto/xaquIJvl224V5PBMixgI5le6oKO4fNYLqsgBB8Fx8fdfxVK5Om
dIdEom8YllhRBSFk7fn8x+CaFDlXtenW/ytRlt10dPmYn1C+Jwskql5/8yZQxpxMfv6E1P76PRD0
7fMqXkqCQApWixWpiwk19DCASPU+e+EFIBZsLFn/Jg4LCUcrtUYoGsiSTgjETpdCvJ0lSXJMm4Sc
FGnNDH9qdqn0nI36CUVurpklBJok8CD2vdswQHtG+B7jVzOvl9L+qjJzBu4XkZT5yRN/EtBGJ1P8
WVxKrVfDhLsZ5EMHMnfuV6v9oDnhsLjHHQ3gl1xSV/Q/Y5Mzf3XTWpjLWLSGn65xposjWVafPVo1
kkespA74a4sJDDpd6ZaNXG3CsCuBmpdL3+koFHJByzyTl0dOgWmL8FkLcUGrF4i0lv2hJgEUpLfX
nQxVGZCmAIzi9hsaDm/umfacfN9pd+r4qpsjD2rCNDhlFT37883Qiw3nSADiPVwuJkUrO+ms136S
Ve1wUdha6HnufS7Q9LQBYquF/GVjZWV3OdBwyjKvXqNBSn9/0CI403CaPX/6Ol1iVZRFFFc8oG9c
QDP/BXvW5GucHx/MVpDW1Il2pZV4W1EATLjG3wKsYxbwwLpy3YI1yvZssSdm2Yh+YvRShGbTzZRE
vVFBekPrf/bCycRR+PkbJpXSzoJssMBWArYZiEfPOHxEL1gjFYedySBDrqzJI2y39S8fL2tvTgjS
QHz2g3K0sN8Tzuze8xNb44y80MIdWfrIcoqo9dp8aHFzsA2sk/RxWhQWlKfuL4hf6GQ+Nm2XT/ul
PWLcDNKc7guZ83OTValvEk3Co7mWZ0BOged3lPsxsDMcpFQPx2KEIuBIzSJG2fD7f0Ny/PvkOE4J
aJL+cchLchBC8auSTTDGUOgsFI7hXh03dWcQVR7A8nfu8ZZg/ra9HL4LsXnK3qB4TbnwQauzoptZ
HAZh2ltarcxuChf/mfj8G8R1BGqJ5Ehk4wLE0AH8AKE7NK5fstS0V/JrmZSRVpGUOzI2moJz9eyF
FXpj4jZ3if1JLQbiUe1/kmxJVBX7e78QJI7fVUZUa6dP128H/LboshSOx1GnlVZw05p2AoPVTQQb
t+cfvui3HTU/7vscgE/rh6Ga2Qz7UG3UwTPc6lXFEF3u7uD2cjoLaWG7Eo71PQ84WK8QWkqT1hW3
Dd49ly8WMMk2DWOTX5yicRz7riU0ykWYoRyWS8MyGtPop1TU8oR8O+1775csaeOwmvidFhUkVz6S
llS6XpVwTD8lfzCFMRNzS2WkkVqaH8g+JTmJje1RHd15qdYMOvzlviziuTNxROANx1voX8UMY8pk
Li8h4QO2dopp3a8KQRPvBb8iHIq8LuEJy1I1uYka+t42d4ZYpFa1cRT/+CcFQS4BjL1OtnzEgZF7
uGhrZisL0QT7/a+VZRiJwR92RIJD2kdmwRY6n7Kr1zYY2UUTA16yEBiYkCoK4v08nIQq+xq6SfIc
EepAw0GMH1rCaL7fWxmQCWqFoX7SVbT9dvLIMKXFPlEgNkHCZBizxTVurpBG4bf1H2wArgu7rW0T
VyJ/+KvQPm/N44U9rkFujY/VEqpCN3+Pt66M4pPQrHxjrl+2oz4SDZSWSd/psrm+AwQPHUhz0QXi
8h8flZpSXXYPZ8FvAbd+0D3Q+BaLdGN5fqyYFeRiNpda4tjz7SAs2ulQM5FwilPz5nJagqK4jPUG
f2sLenX1OYyIgdRfcP6L+oLs/8kc1oClrbMZOAYrx6Nr1PN80/ACwPjux/VgJv35X3c0fo1FN+fq
oRGrpfG0CXA2plejgkcpPnFj/gZKTyqhg2VLXiTWGleA6d/+N+kyrwZLw0+KlXo1eyHBYdqd7lCr
m/DAzz7Nl3x9NaOUEMSywN+eW281ijSTTQBVbkkzQ5HC0KpSLP15jSFZPzkNzJeTZVqqINfuWpY+
neDZOP6IoRWaG9uk6CiTG0zwOKoMu5o2QVZqnyNScZMaU/9EEwRMImBOxkbaK390+G29qHVe64B/
M7OA2XKeJ3d2UF8jA9KkG414QVpvh9P1cz6hnzErXZzueTJ3kbNBDnMVLN3MUGf6KfTFy31lGIta
WoRa1aeWYOp3pAXrAWxqWEWAkuF8fFDuB+ovVGlCbFDmtWuuWlzM3Ky+H08ZxoNuLeLzfq7cbbXs
xydnbBAbezutc96nVLKSDjSM9bDsk5UaHYh6xrFdP05HIQjqQrPG8jArRuOxrIJsrkYqYe9CrfTs
2BfVRTD1RLeO7yRKzU3Q7I5VgBrVj5BD2Gd8u/tC62UFqX41AWrUjc8YWYXgOY/n0gVTQZG9PABA
M56Ai+uEEVAn9YLHY8XiZJE2qEUq+CtAQaXwh2f090uB7xGNyjLUS5V9NI/5L1smqvq+MLVlZA5G
WIW0oCv8vkRno9NxTLi4+RVfHdisamaxLxBPJhuICBDhJluCyi4HWwZ1A/AmazPT9DDytOiLDhxA
AABS6RZPThL7WAZa6npkoNz9fFmh1g+Lfq7DrIpb76dpXottarSY/ed3z/c1y+kZGsmvfkem8HsT
1NWOy89BdddXQVqxaVElXEIYsoCIM+3VzF2g2eNDsXP8W0B6yLyFQbQcxKaXMebpBd605qL/qGUy
i/XhDYJOy0AXtgFWzfa6xLoUA5Qvj/mg8lII2ELiyySwtqywfSibaBqj5poDf/mPvwvEhKDDgY5i
KfH/HeGYLYW1SaBjs5iPGgyV41S/fw0trbAkyDavxFjwtDjHR2LEkP4/em9W5uUfp7YB3Ir88IGT
nG+4txOjkJfqH6pOHLx/WIjkPca/mm9Qvu+0ar/SNb9l9rvZUPohTdLhKAsRhefz72lIIFc+xGYx
BQPqZetcsOzg4BqqX8HfLV6Z0qpkdrEzUMzXK4/jKhedANt+vxipuwSI+jJvj/VnqsNeFB8i+ln/
yTORE1mtliEJBej1Gp6Qj1pIRatAhxLO7fG939TVL2MQKJsRoeAiSnW0XqWYu1c89EG0yM8Oi8El
pfVHK8oi/VIj41KJEOBmUO1OR/kerpsYVCFHdSTzoXOa9MSVleUMWAQ1ZcIXKQWTDm4sKi9rT29a
x13pxtXoeexf0YXktkp9U9VKBkNe7TAdzyzr4w4pSsCNDA6XTmtTydStFDw0sZVR2cyIYyMk0BMB
Of8chyEpzWZ3b0cDS68rmEhABwf+TFvMpyWBv0fhxuWIPEP2TIPCws53kBnxWCFx4bkjEvtkBerj
YyXUvKSXgfXBVI4eZuS18xH4CFy8E6g9WXZJwjkLvhNYeb+PIJ1+ndchqfAJzhJTOE2D5ZF03dk6
qlp9i139i3Dxn0Wr+10iHerzE4hoSpYB7N1ep2yQ+YXOTF0YwLQGa1DbxBHy3QwIEH4KHat6NOfp
eplBlikJl+l8+/sVmPTrLI2DCjuEX7vWHDfw5QP+WNl60uKUwyH5C0EGFuNmDHD1vEXpFVHIJKw7
U8gqBNA/Leh1erKE9Zmg0RC5egM+nlI5F3rzTnNCpaHkXHFhkM+HKvXm8XgzSbEU4SF/arGvGg26
Uzm42rMTWqdUYSIXmhD1wXoMQgejY6K8sS0Z3rNRF5pZ6wr8eLLQNBPwHHEY0nj9Q2Ov+WBEqyA/
7vdayECm2g5RaxmnCbJfAdht2HHo+JpYTKy8FtNt3GttsXK8goRZHE4sZzIWNZxubhOIsqrJWI/1
kV9v79OknqmjvHbllWMtZlj6sdGB8PPuaAzrCBoLTNNfwZ7f3E7GzyVqt69WfwhQMWSqXbtpCdKU
T6CUgD2/ishdsLO68l+xeZj+5qJSFujiQMHgmxiwhIrJ16LbFtMmcGb+ry3l27o4G9a0V+i99LyT
v1PuG/PPdvu18CygMPSquvgkEQxn0d4AEaJ35cVKhz9cAzDFdWFGvFpsjjZzkzPjRorg3o4RZkfC
rTWd7gYxDoVjIDQMqtFwdpdq24JMR+pUUI24ghYwDNAs+DB6y06lFjWyHIa0Vo05/5PIZzqXjlhU
z5K0mhKaAEm77TcEDCqEVtoVatJ3bUs0xGD6pNApK94kI+Wvz/mVxKCCqSfQ9Y2OC0C+q+4QNx1K
R7Gvdl0AAIA3wAu5HZ7F5b6892bIB5RMkhwqIyKHa9RPEw43GbSNoxqjwYaokFek4T9Gr3YnxJZJ
onYjakT8s1V1MrMYf72i8fPPTgvU6rHGRm9my0cbfNAZUE3Hqq6dfv6GEplnKCj5SFk7YeeUcbUC
StJQN+hD2jcwekly3dJIjsoCqFTqXegow0kU+E5nD7f0vyAetMcmNwumS+eCk81xnLwgeyVpI9MN
J+FBQl9ttrBkiUs5CkfPNH+gWaGiwZYteroSx6xWbEerWoHbYkb9JIJtCK9M2dtz4EzF4KvBskBT
IHdAQbpw8NIAK5ZaVmywEVWuJJpKuzALhVgLEM8cghu0Fc1Ou3PAUe1Bd1UopdNwCJiFyuiEtYhV
FB1E56d5Jrs90RCVp1N9ZBjA4Q7dE/JdywqWtm829LHeIUTjWR7BWkICgEB8Le0vEIYIEA8SDi6+
sB+t1vJWneLdsq8eJlWlrxLOIcRo0OkyOMrfkb1L5M/YSaVIBaH7Uh0oIH1XdjryNSSohoFs4rJL
66hg6JgNwmM1VK1N6hz4iFLxD7/W2WP7leKiGCa5lZoh94aSyLzI992AwdRs2Stc+ChtvRFwLiwv
1FrlXCVgpaoSE9gKef2N+nv5RkTJDOz46I/mf3mbuxDIN+jIa7wzgNV0GnzbLEheoSEUaNkt1it0
tMkegi7ODzR6NX5Vxnoer0JOrzDdd/G9ptydbEZDJ/RvtIMLI/GjlSKhRuw4b5JydC0WuHHS3nS4
fC8xiDUe8AvZ6y4rPc0ITS0aeEbliaEXi/0Nl/0BI7xS9ijjcN/puy2UbuTwiLBP4LdhM9p7MZHN
BGY6cV9P7t9JoJ5vJ5kVWno5Y1dTvOELPULJDAaNojvHESKoOCLOn0WeFsqLSJPGFyw74iNXnuUV
0YBDNGRrZsO2HxIepsZuOe9ND9h6xqvQmHkgwvYRN1Rxgd+H1upOfScLWnXE7VK3BAfdwET02gPu
sFO9yqJzOtitaPyaNQ4RLG1mW24wRp+k/sbllGByTcEg2q5QDYuS0AvVZBpFshG8U0P///Ze6isI
4GOm53mmpLR3SqVezSwKcx8S4OJP3nxmGYbmCXBm/5IpFYvkfbuXVWVhQ+meO/g0XK2UQ9Kn786V
uOU6QaOJ4kDvyXrPXvwtlX6wl7INl4vhi7bwBVZ5BpUCQxeaoy8+zRZiY4sMI8JWFU270wJEFsly
jfwVouV88yi4mNIbvaLAIhWOjP5bz+zJhCn1WEtHv9P8STIs8IYlCmuabCS56//gWlnk8qQSCiXD
iwHjm936ZXjSMLXu/A3/EBmMBY7NGm4GLurlfcdgbls2hbPEymfVkmhD4ZnZwAMjAz4RHc38yVfs
ZhB8+DYrZTtEKBOEPsU9RBckqN6zci1vZI7gUKFHpuqKDSG9syPojt82fM3LrZaO//Q04lpQbBfP
XR7eoYKP2WNv7U5RQcTG5jpg7P8sohfTe2hiZKTeuqUl5rLtcV+A8uhecVw68LI9feO/ALlDC1pz
BGS+eobu63GUivvx78Qw/3xbNtanEK+2kYQggL6Bh4qLBB3m0SfhpX+1QVmBlIxg2jtSWif1y0w7
X/17c0MlbQfb6Sl9Zjb+FxfwSZNEkY2BO19teE2byNcQpZ55njwcp7jb27Ko1tFrAgehqftKSJwo
wgO9Fm4W1fOd6rafd0KvVeROUJi+aaEijCnNUNY9MGZXTu+u0rIZk8jQY5gekYyRq86uJ1JOhSsK
u3e2bE9jvK5Q8k/TzgwTRnSNlk51MdWohaSK1BaN8RtJ4MdGmsVnjzvuR0w991o5Bl+0yDfl5VsN
uYHWTTUwxaUk2+htgnA8WOG6ueUtqObocNf3j48ofEUNjWS6QqrE0mtW9flg7hr/m9zI2lRK5iVB
m35xIk3cVuDA+bJ050e5/mwSPfq+ZWwHAtJdpCbWi2OvT1cJSYEKJ+lX/7536I6VGbamhaAgvbZ7
dj/R+dK2lSrSMJxyYGiV6zizULdkn9Hl1vN7s55wWeY5HJ4tzxjVHce2eMU8KI8gUyzQztgGT5BQ
utrlwjUtXNF6KdgFkHtKKkva/OY3z4XFS2PM6KERE4n7D/URu7paRBXcQcDaOe60VgWNHuiyCsq0
lurpb/tvHUJdKqUEtOT3Tf0+C9bU1i7vMeNpf2Po5S7YvfQbszz2mfAYMaleVVIZ/xbvMj9E79rs
WzLLili5wjM1AKU+Vg8Ceg6VIJYpdeIWkih0XtkFwaPMuvuNYPetpFPAJv1GTAsXfRuRoSiJ1ycm
7Tr1RRZahyS/UIaHuNaQ/HCsC8KDpNOWI6X05tvAAG80EsEFRbmYYti+w/gk0sipC4nKLWjZ9eaH
ypb43WsOHTNaB8t38fFZNeUS428jqZTGOs7kYXU4WKgOGcDF0PD63jyk1o3m3BRa2hmj9io7eJo3
uHGtikr/OjWeYHTUowcirheqEy02JOgI36Sdry3qhT+6QftcqNtLZm8hYM1aXCSXUy+IR23RJJe3
Efn6UxJ3jzknnLQso58JD4OoCCL8otLOSLH5S0IBtqxCWhXQ7wtEL3/x9KVOS+oO/pVnCfeFz9wQ
JmSjzwhIranISbvQiO93GR+qLBiphp+2TZ4u777PjGZes8k9Yts0NuiKVld68/9JWt2MqzL6dm6E
wN9cGeayZKM0rreTqvpP8Gty0tKwikH4hOIBjPHhbisQ5WROv4f4EOWQrW0oqdj+M2Oh4Y+JL3SO
+gnLKSavt+XYdyi8XwNw/SpbT0JdZ+zbr1+APs9S/RK4n85J92dRNouOyqO4q/sXnbsRwgrmRIFO
LCh7L7gogMgv88Ekpj2Z3gVHpfuhnCoIsZn7IbejPwQlJ6No35L3D+57m9lBOlU/5NJoDdQoT12I
8BnNSulOeOJUw+Up0RlVO3dhZTUWTooIWNr8BcCHxvkJ9lk2Y7+2pYSDzejI1ePgZcoZ82274JNL
N4AqwyBwa4ZPfQHHS/LplUhA0CRVfu0hXDQninb9RC0tmgdsbGlsNQeZHd7rrekMUvOhZodbI/3J
rfePpfnHyZOQ7p8sGpDVLTxgTiZbrmzhOr1bUxyM1AC6QF4HL77AK2wAc3B9wGjPDMlfalb6PUuA
Ah5jpx1zdQk5Pb/3a6t016UcfyOPh2sAaMFNZysfLrkzhXLJNCibI1lM/bDkvIIWiuQQtY+cqGHN
ljBkgDmEaPCY8dfkhKpcO+OWT3a5fn7SQbcNutWdhI7KEM6bhllmFC4H9tx+cFY44y+0uXdCUN+K
bF/EIZifGfOYDzhSs9n9kGRv+8o3qjgtaZZZBZKaDfoj9AxaVAtpQXz/KuemdUSkd6cjroDhZVzJ
ZWMrxFUd7s45tDq52pCxUqszb/KFmWknBHM31+eEvRK+OKP2Kdc8/4t4WrTiQP9cbi8HdkQOIh4p
JiSs3GUjROmPQjaRtmjKjf4jqCg6T9mk4I9Fsv+GFFp07hz5Y26A2w3Si7vlCFIqRB64xwwkqQXl
7XNtqGromxxVAlM8I63xXz6IzOvc1mgxxQKS4k7zFiduvzvxEyotDUU0tdkm3sm+w7bLTXi+5Obc
TECdWb3ySeDE8psYM7Dcoaj+VJWF2e6KTvoWwZsiUxRnF8EMzQNc4oPjffS8mc4n+g53P2l0HwV1
syKoYg6l++uguW2HAjGq71CMbVhTwO8o3TIW9g5XBz0z9jvQI6HQGKxydsTg+oXE5p3crXvOy2Z8
Vgm8sKONIfg+0FRqsKq7byCvMe9fu+XqD2M4Gh7ri2XB3s7OYwpquije8V4w+oRyVYUSLosPW9gn
bg+rQbHaP1vkOw6nm4D95Wo1WP8GOdmX8VIreMV6D0RhRQQylS+fXMOsWttxcNUu6o6LZs8dF4NR
71SIwQmKzn2zWX1R2pUOkiX2X3nZnxJkOlHff6KjzT1SDsCadCfzTGS60URJMfsUhJGwP0OxNotT
sIepwSa5VGrpq0+CCl1eGLPpu0M/dMlX4NKDW+B4O0cxj6Q2dLZVB9xEXxZoeCymdA86t19rNm8s
zA3KwwxHyK9zneLjdqqujKCf1tQdO6mvjO/+TsRZXpU74QWZP00Z6yvjXmFOLYmRMEygnO0jJX3H
kSJ+kNLQHuAvoJT10a8Eycr5BH4mQO8S+0+OBKJfGYaH2jedlGU/CTwO2UQMkkBnYeEPcpFZZUfK
+uGueUS8WWY0vnBIZYvB++JldxeRBT7EW2Yk51Bug+khVfNluJ31odppoPsokgwNUoVwfkLF+5KV
kSp9P1y+DETUeyFo/b+/MjC15mOxYpminNHq6Z1QwZGAZevGEF/iJHDJVhiJRNjyEGJ/2icdtSns
vD3F1rV859tKDVrjkRl7Iwt4pHSvgVMNVAh/Qkmiutu/D4o/soSNHq1HBKQ25AtKppYq/zz7JNcc
DXoFN4ITgk9G62Cud31K5Y6VFAVFQekDUi8b/08B4ZyLTBFm711sPR6LSn0dYYMXj/V5Nx4elDd2
BVymPGEd64lClbDBYvZU5ks4v82c4TTMWIW5mfnIxvtGjtrBmmjD0tqJDidvF8iy3U1b2gW0RW1N
q7wU0SH1XSEBiSHoC8o1isUFdyHKKweQg3HRBoBqS6vUEDwkT8OGjDpvd2f3EU0E1oc7e1s8H6Xe
QQf996Ux4j2RHcQO7Lxm5UhVtngkFRXiuSkYZlNiPlzjH7bI5RvyRs6D3wF9uxENCQkI99aGrhoD
kEDv170L3AR9C6/KPiYuXo2p5MnKbFrla1co2YkVKjTTT2I4wIpiuS7I9sGnw1Cj5ukKHpo29+3e
qtlkE4WWe7032sA92XhFwwcK1PdYvL5GWTgvhQFzZOs48W22a3vAzEBGn0GFvAwo9wYqQQv5v4/9
7YnoutwY/Gfh/i6rrZpbsOgyS4I81wQALiGIBH1S5MCefyMPqZJmBPPkO5E3+7pdcCx/nbTVxT5B
FLd+7ta9QTxH8nJpMoU/l5Ew723SC9c1LeIkC6E4+wANXjp2Je2FjnzM9LvoYAmfi1py1uGc/6xL
MmaoEqs79s0URLjoIhPVNYSlZa4hB3alQ5PMfYbRlQ47U/ffHqTyNhklyR4FTOP7xOWTx9EBpF0L
hFblEgkQQAIPgSfh0ZD57AYxd5HyvyFb/S5rDO0IxP5J0xm0zqXHOh9NbZNB0tl7p21QhiOukZg4
w/JJA4fAtajiJN/SKWKutzY4tsX2nBzWTRbZbWiq95jdIqSLjbOyM85IlcASVWJ3ftThTh3E9LV2
fig/BxlHkMh6ZTAfoT3gVwqec6ff8M0UlI7rUSGEPXlCI3DP3z01yJNdsjuwyMgL/yobEQkSRIcC
YiFLngOUEpC0FR5M9J16aY8rrmUNTOtyqI/RRBkNH5LB6U6Uvw9FDcgaRHOXzWhJ9xL9UlozSFAt
YsyuekrayDA1gF010Uk1tZoj1tl6PtsgDsYneMbSFg/zpzRDm964dYJtlSAlqyOugCzdq1Y/ODe+
yLD8iz5cnLO5R2NPBqFbFAV8sv8gFn+cJeHECrW/ypmtZGar3a9O5/4Qm4AzyUrpxlnjrw0a8w0p
LhuLd/CASZDWzUftF1hMd628DQM/oQ2jhRYgAT5XmRe0kXaHpIP+zYUJiBNcEcCD2KuaKmcMEx+i
vdOEH7+rvbc3/F2LuyrqiXEbGJa0DnYvQjOGdE3AW3p/j27v3BO3Iu7HiFWhn44BE2ZQqsqzjzzi
qsgp4CQc9+ZL40OFkVewh7scjIdWkaUS1H/gggQHLZ4TwOQfMvB2XJ0AksQPpX5IjCP7UAFp6lx4
BqNoO3DXx9G/zdVZRqSjTbMhq828hqsLJr6f3VN5fEdbLAO4rnXnCxpwSYWWqCY0Aa6K1V5Rk7/M
+EzDyyQdi7X4WXpC3FNh9Y87+uIJMpb2fhFjbDWoRQ95sOhtVZEWhulkL9tCKboxcDgJ0aWWeQpv
oxXVBLcIerhba4HoKRFGCgjN0E8nd37VrfwPPm5sNcVNUIxljGvawxc3KJ3Cq8ZDVVNCkWpk55ze
gjD5QUxA/nxmOv9nv5gTeKo3JAqzf3bteOsaSXmhq/JH2xmcd88n+R1IH8E+R6kHtOBxSEK8ReI4
w9SddUEPR96YzTY2kfl3YBzLAVsW1P6eS09MtLv5+holqmFXf70r9i47niCKSghkoTdT5CjHWSmf
Vj3IVyHN5haH/HIkMnOrb03Dg36U2N1id9KEIIr1193FdPYb4y5nsbAqHzz3ZEoAjmKlXiNRaDiE
WYnvDRQ0dgTV/ey5bDnM9BpPozka6cHlJl6LjckJUpMmUYw2gRV8uNwBzZPZgCqqk/TTHKuf6Dba
lI0ZP8EKaROPn9zPbsXd+XOFGTJqjtjrwBSL3QFwHOJyO1zT1+WiSqyjdKuEEVu12YFYHAxtBupL
L5iX37agu2AF7NhRHl7pRzZPzhkUakJSNXN/rfNCGHpmhl7AvEQhLW7qFfELZfGwPeYhzNsuXz3o
/1r5bQK9capcOZHOoAwXPWPqpCKVT6LTKCD+hipU0SGvxdRy8qoIlvL9HC4SSexVil7j4r2QETBv
1ViTdjgc+FlAnr87U0C0oe2W3/RKXjDTlxFJIEtQ4SPwIC+yypVqVTe0BGy2LBb5VIXfQI8TkeqK
7DLaI3o1SxsMEYw95bsXwUFngfdooDAb3bgiVFXuUry2oLii9LQ2jvYc1tfNUixfcb4BssFoatrJ
8EsvHNPbyiF8Qoiawty3hu0t++pLuTNygG9SzBUa9ThUavV5Jv53j2rlP10wIwpGdhIJaYeso/nL
QEyvcMk0B+E5sUny3tdL1z3i64fhuBvZdwlRYsR69AsQjHv9JCr6Ozixc7kAeZDYoWUtjHq4jEVT
q7UAO6B4Ghd9qd9Q60PL8aCEyxV3AxRp8jDm9s4KUtFGNQFdA78bt/Zssnl9EYDqkIGggSxYhDn4
+9g36wuwPCjTWxuMylTTP++oHJ99HwMQGlMWVuLJx9bkwY8ta1VU7urFkvX1CSUx9Oa5s0L+oI5Q
L/Rwn4xF34UvafQoyiSW4RNek2FLV1HkMbPBcTDFxhX9Iw9TbilVqf+9LOnQYZSJOyCl3JD0S/kS
kkH+qHXIGTFatfoE5FzpcRExwsJso/FhyzRncvVup+G8wollrBbK74nJvZQTvSKQ1jF3bgeMdHJY
cEvvUoKj4zEI/643U4JFmXdtSK121OFXZVWAZ3XGgE6qIJg8RngngbtqahPeWWGL5WqUja4HkGXX
aR+nTO3GMPfY1h7J/Lg4JWeDXrJKFe95T9CdBbVbT/RuYhJ2NEnrzaQPypwax00HOh7M7612fOGZ
2ceuSh+npvsWvTHlRaOUEz4j5k4ddX0bDwDyLKNk51TmqPf4kkH3tV+RIqbPXRq2xdUiqQG0gdTq
yykhgDscjElWKbKOShE8pApKbjkFfWxC1mnt828UeRZak7F/wJ+YD7Gnn4Ie4Dtogl07L0x1XSyo
kJI49zYdh2mM9SjpPYvC9OGpbteF2NGPeXMMJIhppczX7LE2vZu2At/OGooiBuoT+1M8HK8/SjFG
wtW2W65NiwN3t7lz/isMqsJP6nKLBisFBfP/WZamqoLyyFzpLKiAYU8X1v8IZS5QZwughyFCDj1I
6isL2fvihiNYuoTVG8xoHzkAx/g8Yw2eNeEMTGTlATJ7t/ok4S+L1cro7/ZtR5jGnGJYiPT/gkwy
OMWyHh0hgVhWd31JaIrNn3PGkyhW8SUmoJAUQ9IJIaSjf2MvqEEXOBSvgznBA+Cq4Wl0oMP+qaQd
BIrRa2+bT344Fd8NGx4Ihihe3ULLSHbEcSAFSTzC+ztOLp1eUnZABQWsHhfOk7fK6PDW5khDxQpx
mN/BGX0bVrdIzPiiyc7/QTZ933/K0ZDsX8+PTdpKcGjoCA8gP6yQTw3ihg1sScsx9G2CTSc/WT7l
1nJglWOuQVeWiKjV3hLpSbjNi1YzhnHcgpI7smrdlsP3fIR8uiJt0gj0ThgPVxh8Ux/3wJwZ6UOh
1h8f+KmbXb2QOLTDuJBeKxhntcBxNBAxzGhIc1RgcdPFha7lbwQDVi9h+d4TfjQk67KrCHLDjnKX
X9LDBdQxJiFM9QyaT5eyie8O6ErS1tb8USI4ZEvHk85Q517Or619uoHcNEoucNHYTLH42n5NfDJt
auocxUZhOUWBnj+FPgSBU/pVq1BvzllRh/K1oXse05IV1II1hQK1JbzEkWHCPvC/kcamdf3X+eDo
cGtATVBMAaalHhXHYvmuDkJJQwCPd1A5lX/GeoadHm7USE9lRHBlfDYNoxPG0K3Xs1Hr7VzEZmkV
t+2ryfnciHqKMjgMmp5TXqAa4eNCD6Xppr+8dAl0fdBx2uvWHYVc7/WXnf8By5nQzvzFFBCmHgmW
As5211oGiEUOPLQSw0dhtoK27ve0TgoNFA+z5N7JlxXIexE/a9k+rL9K9H05Qp7COMdS8+I3kP2d
x9oGb7BaeTnw03NA4G0N/7kjV9N6MrWubZ60arGRcbQmxgSSuK5kxntHXNbYObVNacF5EDXF0trI
lLTj8XGoHgEi9HgCnjdMJVbLlsEYXPNj6LBwfr1pmBDcA09W6pUAVSYA+yD+yfLBvdaFBB1Fe4nd
xjHchLFsZzGDtvBxQj/sdn0U/Air/PCsmfAE2TQE69IIqRalOCQy9mkJ46tLpz3ZS4RFk4FOBv/h
cipWvmrD18NkGweqsbHf2YFFocY8DZ6abVEyey8YrtD674HtWD2ujd3nw8MnJs0/LuLY8R2VPLfb
ymuIYT2qgX871omytlH3Vjnm/OlYWN59Fy1b3i0qQujJ7U5BMx1aFIvnaMxVHV1LOfdmXWmQZp53
vxybisTzA4IzNKQ8UwXYCZRZ6zyY7O9PlKN8THVRWgUXyAfZOismHqxbm1oygP0mDAi8fFMxEW1y
gXaXRebuW4tC5STInQFSM5ky2fHebZhd9nIHOjSdLKWwxsraLuDEGMJyuh348mQbirn0FhejVGh/
f4Ga+0WKcvWVjCLDgHpfnUmwRnrN16S2mRW3YBGQZtMFSO7qK5Wbd3yTrV8OBPSJz8Bp3wwVVvD2
kdCJkKmq4G+Aha1GPLebI6kE5wmn8sMlyNi3MTNZFdu57KJcgYbfWfSNBWcTHvs0luGhsKPGxeHV
45Zd1cP38pALOit1vTB6RTQrywaSqzcALZxAq3emL/4gDmYqIZf+E/osD6cTaH+LFBaZrLBVKiL1
Luf/JI3tthYtSCcfNcyP71sWcoeXfCYgNPuKdf2MTPwLXw5Gn6+TqWLEO0sTmsoRc1vdSG+37TtC
sQgqdW+mHDWavijI7lW4VMgGBZQgyouy3lLF4uC7F1r+p94JXAwVcdwMYqrHgMwWPIbZi6D69RWh
i3m/s7kW/SydaDKKShP0x6zmCZf49yPAoNJgG+mDTO/fOl5feVo7Cu1uG/601SWamXCL+IchF0nY
upr4aKWwPyJTS764AflzyUnvF8ZHGjHRVwcctshjazdDrZfleqqGWXz9o8mpukXDPL2Jeg83Uaiy
wYGq8Gh71L2itS/+irGqwS7SHzpxRRwVxZ2C2A2/y/ijj4HCgmmIguspO6tvG1tdz1ccsKxWbiD+
NOqZvWsfcez6bZ+oajAXZBnDUD3XbvXZ52ik7j4FQpN1f49ncMFJ6GRUpzRbDTThTe9oM3BQpXBb
oQ2MvIH4UJD9Uuns+zQ2rqIGkbRHzhV1aZeEjfwHAZBvrGdd+fmjTWdWawDYLGUNc/HOK2XfGuyp
kuDxD1esZmHaZjVxFyqeZxVd5NjgR3EWgGsTwYH+gcDsRdNLVKSHyMSu6GpaMYAQfqhHP6OLa85q
q2RA7ANTCepCevvG/VA0vGThGkXJ1j1jgMASySX15tIVbEL1fi6DzsbQ84KbLNJ7P0zpsuiG3MIL
/fjFV0YMPYu0BeeeeHu92vYG6PjX1IIRO0tShXa+zUBbf719HZNEQiiXq1l9DYM1H93q+P4XTf88
RX3CduQqRozSiwmkYquto4Ry5HVI7MRu1FY05m2RQMudtTh7kKNAIjL/oQsmH5onOoT5rHWFJ3Zu
NEo0yUBB2JrQ0GuY8LQyh5IBIPFMBKu+mp/1BF1SaRndU28mAGL7e/KMP1xvH3TcHVI919Hb0v9N
LcnX4yircGXePZ+3SwoUL1SAIVYK4wB+WJ1b2pOMcHcz4kQxCxjqyRerX0TqfzW5mGrMh0OXm3fT
Vv+Qf4wk5F/uRYrRHRAmuOSOhmXvwjxdoZJ+PTYuNAMFQh3Q3XKvnJ1HDEdut8KHBnv9M/6Yr5IA
dsKRHUF0lMYgCHBOMXRHiK8ZxgnYsuhkc9cG4FhKERzEKJ+y5idc5p5rus3Y2gk5fmgfRh/jVmQA
Z0t4AWWLknrcnq7AYAgrj92kTRTbqLebTzkc5jjxM7rXZIhNfEvJMYgEcx2eV/BUKGPTk7++KLJO
9VH2WB56IY8x882WfzzX97NgpF2yd1jKykssmxqgoXSIdLqP9JOMlJV4sYMp2oR7vMRzCrO5VS1Q
wsGsB4KFqx/LCzfiFyz2v5fe+NiZAnYqEaH9bAREQ2vYkez+ap0f458zRgA3kL1Xr0XeFkI6HCpm
bndK4qTPNWrd3uLJA/kIj20dhfCp5d71eVkx7BOVgYp7I29f5mbE0HtNxhRyoh2lryNjQrtYyTIO
KD06o1fo3X2fkwswk+aJLXT54Y3D7+ZBCd6mJyArdBEsV1Tnnc1meMupNuAgp/9SSxn0eZ+tzvGO
tGcpdVsBnPOTD39qgHg+pC2nPF+A0/jGO3lceuGd9TWiSdE4GqG2oe07OZtYDasUW4/B2rFsnh9q
8ULfUICFO8tLfL+4Ido66vkq2j6ZbWung8+HA/AuDTlVOeflEV64pfJ8nua8yuQlJaZ9vf9I9iso
lxJPh6Cmf8UIvdE+8R5Uf0BUoYWyAyW40tkwzDUX7aSUT0GHOSTgyg12sFqe+Tfwml/2qiOUnCyp
1x5eiVzvjgEFsJgG72h/rj4Ck7PdVvbQ1Y8+1juT80+ar3682DJBRfrhqJcB9L55s0L4uf0Y7xgk
XMQ3RrDEjd34PQLM41RqaBiSqTI7Vwb0wW0iBdW9NChwHHFbs5B7VN03tSJvK+dUByBSSJwP7Qy7
Ebf5C8vrEe256D03QxRyXNBJ6HwkwAsitUBTI9/bkm4wIw+H8rqPZltQlhqPiTEOdsQrlpQ/L9Qo
cEWTuz7peopN/bGUk6HLsbfNk0E6cmoB+0UE+Q4AprlLOa63QhMVIGh33Mnu/txm4DAkHDwtDMyL
RBJ3gWYqARPCWrdsEhtSctepRcgSm7Vst47EqEG8us4O63lEvk93WZNrR7nFI9uiCB6tBmC0ZDMz
GFI+OstAZBHL0tDbz1E00D484GO7ZsBUY1+FMdkXdOkH/cVadaGsr/Q1Qmb8h/09Ww+HfrtUnpMq
euhIbYvHLGlCET9EdgGkGgktmx/Vqj3PATACaO7JfH6tbbg5zVBq/pN9mws3QKtqCdB6+JBEIstB
WaFFUiduwxSah9ADMEmGV5ndA7htf2XNwc1zOMPPZ+XzXp+SnAT5byu6refpeNf5DHR48guvvG/E
oxwuzGnm16ThPpj4MPer4HoDdm6sWM1mxoteS5gR+YrwVaP2Mr0zDUjONOIHKeiv0yx/XWv+tSHs
gH0KshTJbIkMm6eMiStLcJ6TjvtWtzT1QUJq/3QdWkDqZ9Xk+pFhkZNCe68uCNjwMEMpFqY8xBK+
emuTe4e+rs92x/7BHbQfG/7vTG0Ad0w9CYphRBpEWHXu8SyYKj3OZKvg2tfbUdfCL/ky/xJ6kZIv
B8KGOksbBkOyWOnLdT4PQvxJGwbBpDFCQVWpmxy/ydOz3rIVLbSS+JJBpdugU5NhQI58EniXvrr7
7Z/Lo5LtWp4HOcvDuxJuyr7yZ7As7IluBA9wmevHWbqJ3p9Je66dN/53FujbE+tKmVzeGTawjksj
BnXiVLP45Wzc72gLA/qkidnENM4/QrpiBeUclqaHUI/rv3hVIsRJyhSxTZqOouVaQ3mGRFZqulkF
QS0f9PDo4kN5+VQ04qc0JSXHZ8KDlV2kobfo7gax+tlG4SG9nI2b4947/8Li5gzrZis0rIzPWdSZ
HwJ2NM8Z0arkpFhlAKAKKMMwq3QLg/LhKFY5KFbcKfu8JliRoFKQtcIIUZykjxbsigFMFn4DKLpw
MzVWQIIlYWQfEB/7lGnXi5TnMC1JUDw5U1mJwObdSB806SLWsUwkk4AM/lZ7cy274+6lzP56Xfxq
5kP/vJNyb+JBuelKEgNQGNcVkmwTW8ijjy28OrpB4QU/2Bqz99bckyuJXHoLcOfDSQHqgSyWUin/
rJ6LGoLbiCfAtLCr6YpOwWP7PWRhVGGRCm0xk+e033Ixf13L9qv37w17JLrg23rqAkP2/u0NMsKU
vUtetSrJ5hEEFpNld2/zoJZxgTR60DkYLoftG5ewYQdjG6I1zng+Sh+ph0z5MGu5oL+YXOZhxwLf
KgVTwIdsIvAo41laiIceENQAo7rf3JyoLlJJWYB3vJaJS+S+54Dv3RyzHQwxWnSiflhxnHZrG2cb
yv6hTAZf27C2IRHNlmxKb2AI4Lu5zmu55XM3zRsMdX5G/131t24ycHSKvvvOvO/cZw8f733/GT9m
Uo/rZQJ7dPMpRpBK4RUlZeH4vT78Q+vBldFiBuOWBwNvpjrKq+RrKRxJ7T3ewrcUpb7xM/g6KLtW
HE0/4tC0RKCkttDCLSvgGr+PeKQxruRTfevIjv3LDKYsJ+/6WjK0RyIUJgIACZctRfxw8DKt0lya
R2C4EOzybBCyHOKIb2a5NbqDBPq6T8xIz0xjK3h4iU0jbWKGTXFqPvGt1A52LLf0Run/H08AGDco
YKmlGTFk8Fk/9qDI7QxdauA88PHscGoYYV8C/PrNBcN9YSsns8q5niKXUUX0/HBWj+1Lb/1NU1Hx
1Nll/F6PZAvf0jC6x7s9g8hdjMNOfHus775OUjGYWMFCFzn5tHAHLjzahcgPTfRq0jYNTPuosRdj
QAASl8J1Lhm8UseGrRuIoUIDPvPhwK2UGJ+wCh9MzQUC67i29244HO5xKdREwtjKvYp20GDks69J
+v2P9OdsG7WoWX8L7dPxni/6df+oXPskCYdGct+b+No6YBA44+Las1nD1J9C43xVVKwSri4FTzmM
qPbmjov4pwjZ5pGKil3mDDhlDQUVcII1SH862YRh8wCR3KRFnBtUnsOG2E8VwJIevFaB1mO2zbNT
NSp1glbNoD7eCRa06PFm02lXPWOqeUA8Gessm0FSHpz1nxUBRMM6h9GVLKWCytvGvZHoziCFm8Hx
DrvwaF1Y76bAismocTdJVxdnjsEXyiycu9mXFz9gj3xv/n5UuLqTDwy1axCKKYp5p0VFYc6pie4n
RAux8U1gDh2WJfFWggOaoey2I3FTZHT+g4R6mrEj6veFGTjGupZH6wB1/A/BVaMse+vYGggArDNX
iwheknBOeF1Drm8zjwk77+Vfr1F0ClQgYZPm/FToE8eD0iSNjP3814fOIcGjZoKRcEO3lCFi6Xpz
/zl0ODSrQ643MU3/3CVRxZl6K1J6bfd5gIUiziuVWvlr0XOeBDGxeNLj5qHgqJe7myKYyNbPnM2G
XdOuxCVmV1nT0KDbwFOdDGgGNKymG/7I8taHWAvhwzSDDSV9Yff829RSBpSnpjD7yKDSEFEvfmqY
2c+siKNpUDgK9felPBpTtYBMaCD570ymbxJ3hzFpDoX7YVLM+S2mH+w37CXkjqjgZqYtNorJcgKp
Q9OI0dujsuCjzVVZ7lOhPKvPHP8UdmSyxsR9h6beXbJ4qH7ksjtQ63kdp1BKNx9TY/5N7IDKExTw
1OZxOcUvpQCBv9Lus+OJ5LbyNvpqRw5nO5xxaKplcFJIi2gjbltOwTju4leFm9Dgr7PuGVUZ26JN
S8rkpNASN4UuEwfGKYTQ79c9cV1bCND34QhqTdYYbe3l4Lri2q5dIsyTm/1WBVxhrEyQYNZcbdtw
/yTIJkj9d40a8ikRJr67ouKJx3+EAdZPlP89bL0GKEIbh6qW5NWWFmB0MV7ACUuUXg2h+osExCET
TnQkQYwxWW9SfZlDmLak7FYxRI9DTKxwuUEoYJ4uvltKPyyqsRI6TEY9O/Av6xVea196BZv2vwVW
9eDON8vKwbgsPUVJPSPXb4yLffz7k1cil8UnuPh9+x//8XXc5e4fOKUiCcCfjHOIqhxaTpyEs9OE
5ld/XdTMQY43DkJkXBe+TPFxt31uPCu09L4g70EXZcydwhzf+NK/KyKu6hFa3zNPgqB2RXjsCjxj
imtMdR8IM11TAtAUxsoWxD5HCLI/E9GDULwWBNOlOoP0H4TFRiUFplG5LVjii0GKreTZpOzXMRTl
F5Gv1lZ4ayM73FB0h/is/KjQQDVmU7KfMunnklOw+lF4YY7ZNA/83tq4V5d21aM65WEiewn2uAF5
+macNcdNXgssbLLfIccB2JSO/jrBMa6xvLRLuarAiut8Srr6E9R+HGmMoHzAM1kt+PirSo+mpVxB
b4W9r2A5/1oCqt5J0MgT1BhiQtNDc9Jh5odjytDaOv/M/+13lOrZOXLnt/tgoa9L8U8zd7L3KBiW
w7L97Xfvfr/vI7X0H7aK4aJn6DDhbW54CzOBBBcqqHRPMTX655JaxE2EufCLcmyOwoKgnns17rGV
VmMlnjHCdNn3rO4jLTjvjiEgPCfz1gEH0SpnM+G1K5svKsstBCZIzv2N97Fyegu8gETr8saLfqbz
0UXg4VsomtybykVmyIlaRYbLUCMrvdli+3jx6gdnJl85C4jK03ZSCcKxD1S3jMmPBBqef3h5oGPW
DHWgnPbj4m3KA3g9QRqE4eV0g6Os8t8cidqkdneQFu03zaL8ahQt5kH87Hgh9P06KcfmNCdvrY0m
ePRidBvbj75Rh1INrbsI8C6xqmh460qKjgyA/lvZaNdGcT3WZ9Jz5qDYVwT1HnM9d22T96+NFbAM
Ob1ZvTW1iMN3HBmLOcZwR62QDDzmU2++ikZ97MrCSqPVSJhCb7EG3CEwSjywHNVlIgNPv00yLyYn
y14T8WyDR2ulv/BDi5oZg78oZ4djG/iQLObmNNHkIG/TQH5ShjVjx7MlJAvUxj+iSQUPb7dUkJXO
1+RJTZFubGfFc7Si79aQEWwT/9K7u4gnFIX8F3TYE/leX85WzBgcs1tnAIw/HFbamMtrgt1C5KK0
qCKyITrhwJgzLI9M8+UZdyUvqxZtlQzIbg0mYS6yWb7ES08l8py3uknd79LcowGlt6tjQgqf0B3R
dCuyqEtr0zi4dFu+P11Pla9vhZWkqiQd5yqUOpETDW/6jewo+APSQeHNwfFfD4nxkWAy1s1qO6wv
Lcy1kcX3X4N0eQ42U3hYkX/Rod0yvPfx6D+wn9D/TNrjOSli6YITwWVusG73w7PZ8vzNmBtUhWIy
OkKh/Q2hVnA+oh+zOk0dMGssQUS1YWlcLKVsjfkQmUN/DrTSuAGwgc+XWUxUNxv3FJobwfnOkmuI
s0qrly0tcXq7CFiVVBJa74BgL9awpldi3MgJjO4ueZKbptUvf2/FkZXZL/L5Em2i2+JdqgDpZ+de
4U7ZvXBxyzMb7xA0g6KIX15iaebVSCsMTJtsZcwYt1dv9uocAjl0jvLKAxAJ4r116jmyFNjSHHGx
fKFr3wHrY2mmE6RtIwk3JxPE/9hD/mTDnboYPC7sME5/fIeLre3lH17omiRHiElsEJcLYTPlU6bx
AOmXm6A+wQuFT0fvwxxjdRUrRG+APxKglJ4TycBFjt8OmiSeGhOF2XF1KxeB7GMK4RARk3E71fpd
guR8Qz4jM8vR5aIBkmI5kXg4hoWhORaa+EC1xGeCIk1D2p2SU+AqjNNYnJPQFlshRSnkfK/pu+of
G+WN08CEx9feLvxLmO0OKHMcnU2+dr72/8mLuWcyhIIggdfvaQ2eFZloLm6zVTsJIeyyrKkIGT2V
YAHrdD9Ab2s6E3+Ir4eVZIuKdj+ZPZHnvqX8UnGXDjhmeaT1KnafMChmXD9KRZlIFpYsG5Z8PTzN
BnNAtZxqbV+DJVeG+wHCH+7ZrGSPH9e3xFdBDr5+sQrgRWLHDRIHxIqLwd9mb2VpquHdwohGTBzu
OgmkoNNwubHrf9WlP+8P1RJAvqBNsS8X1CH1SfTqcOzEW+KMj7t6O7zY/4rgwzw/lb4WIM0nThEa
Ep8cZFdx4rj/s76sQV99eeYd6ACtMJYdr8/TIlmw7c34zyZTI3G8RxFLVAfXp9ygSii4WEPkuvTl
vM+tGOZs23s4hNIhq+daamxDwgBJqA2ac4rmiCEaC7Ew93vSmJa3xATeX3SsoBOEgMWXwtY/rMaW
uzCTcnnCOWCymwhq1TYXBt4MtLDeMAh5zuCM7rg0pE1BaVZuM9fAR4tVhImAQNfDF6unXv2xa6V4
6Cu5/gEAx249itZpdGp8tiRKCgKcO3ggDi89mu/vz+f/VUA123ZM2yjlCMf6kX+2CY8rgtTfWwuq
VdzoMgH2hDgcvXibF7qpJNofPVCpLHiyvxiTXZUXg7sOYgdEwJUaXKJ2fdV7QWGwEm3hSXGDHJTb
Ibw1IrcaHx7EZqYMFJLoZSxhvLL3yyFOCl7faQzmbFtLgGBWSUmW4/YQXc1vw29Ae73xzvgrjTA6
/qSAk/KVfskLA74r/s5VK6ayAt20aVLwc0qyY1s/7/kb0LQfPhFMLfcQ3kQX4jGLleIW3C/JbPAu
wffM2KnXdlrJkvsB9l5eU0SNAsHhpq05imUBXRDbKyj+4oJsKCuv9PlO9jJ4hqWRJNLLVcrhBOyQ
dIibkwC+rrA+oFRxQ2LNMIggjAxQTRV23zFE7G3MH6IPCQDnPd6/Fiz21pTRAemj9nlx9p3gIPNI
GVGjJJLAbFDIUtpgYAJ2aM6I4PI7OBzzUVHLHrwhLID//KeppMZRgxmwuc6qVxCh9H1Kaak7sR26
VxBaRj1e5NVDch59VOU0Yzq2oBj3cGYF3ENomli6+ySdTyVqUxzkJZ7gQg5uNtJUto0K7VAXwGt9
/GpC/4t3x+BQIlTnFNUJdO40AWaw+0VFv2eCiKr+1lMKV7NSkqDktSNRUt3aLu8Dh2Klm7CAA9el
qTYzgn1HCUPJRM/aCgq1rnYy/5uSGIdxr3IR+x3fojJzHpkcwfVYJfE8kqJkxdoiPK1Z8AY0nthC
sgo+PFKyYgNh3KcFWGWWuFbkT4IW0SDYPyKNXpwblY1wdBW5aXwQpyVovZWQrpYNmzybhOQKBlgK
hJWdhiUUuEnQphmAdi2rkeIKjrb4B0/oXgjKTYny9re4krNwQcnhhvED7JAVJi0JF1r6DpLyF1Xn
CQpurVxu8JXqQJ4eKjT1vugJRQ27FauWZBo/BlsYGbCvSclBNXgo037hb3ry4tOEClW2lqTYFeSw
14QWBe2nHxjKHkNRNS4NmqOxGm4I6S05p+KX1hOmAZShIOn9bAVNlk3/5C2sEBST82tjvsmi/3v2
H5nCsnzD8shN3gluYb8PjwVc9VBDhEqbeL3hOF+Ivo1pPdIhEIE0afSFBp+BhrsPSE6OBTlYmgi9
6NNtlqbA6PTvu1jKPv4ogp1pzubTZvubCbEEaos8f7a+pcWasNW6YCHEkwOuRN3T/vX61l5J6gnH
FzuWiKDKBi2VIRK6sKLmC4batx9mDO2o+RdX14VfNMMbgOiKgkiKxLte4IgQ3STbi57XTdadORTf
c7NuKMgjR7hdBvu6GMgF3KIUxPuPPM4x0OTmxnCfVOZwDu7pOVMCQmAcWAQOsQduHQSeHX1srzr8
ZDi+yCeT5l3VqW4up2+9Gea+S5DOhuUnSbYRXxKYDZy8As1YUV7ZL/O/J9yYINKkSOTV6S1fL+XQ
OUdMB57RiEmKKAeR2g3nN+9kpo6c0EoYIAV/utPyEKu8s40zN99qh91FdJ0Il2ZvMlpAYlBlEQaq
7FTLWq9eQWLpCAXURQdHhS6RUkFwFLjmOozfi2FQYsp+KShVHpppMEL4EHFQFkXDVto5dMOYGCat
w45D3QCV30D9xc7CJDHgnpVZvxwwpuRLzc1iGBXxed8k8dOVMwh6xpn1WNsxM3SDJNyGqyjAaeoi
UqkRmIPn4GNFBRRm1zfrrY9eZds+cfQ+ue2ll0hfQQ26SCuQjOjSTHTiIOUOI/oxd+FWBjz3D1Wm
Mh5vOJIbOOhZd/Jodl4qcfUFdtcoRiDGGAkAMGdgyeAiDhZ3bgs0o0nLJU+b1dtsgrciNe5ItLdm
xsh9RU6mdslieeG+r5gnAAysZDOPDZKVzhGLxxH7k31+6KEfnpuSfqJ8yrhjkIYnN9DOwAHxWhsO
GRmRrTTkOX1D2Obhoe5vonuMe5OxRXkQek0Y0ZGjhopOufqOwNa7CPu4lgAT/HCe/khPlV37ojaS
Blhl+3y7k6jDKRZ9vOsfQ/NV3TiUVH5MEsiV1S4nEvvhAiwB6apYI0IL7P/odOMu8q90AKHDrrZ8
56FTfKeA4VLEbfR0AqJ4vPM8B74Qmj6mxAAWmWT5TJUXee01p327UyKJyH+vu3dC9EEz7AEXq0or
sYmTQ9jIY/aZRaImhEwtRvz48MYsc5rMI+6AMmL/a7UeqDuRNm3dqdbYH6trckXN6785hqCprUVb
VAvsFpqkmLUHFJH425SC6zfPMG3zyOOon9a3tnbM0SS7sARY6GhsvXIxLAlg9O4UOVhnaLMUvVlq
m4Q9/0Ol2R/71EWRX/7QWq/krz5q1C+9eKOP6nN4Pahil1QAtPTjetdnRtsvQrvYK+uiQh3Ra4wI
d74lB25Ikh9inLYP/Man50su0nIw2aww3KpsW8qDlG2Eqwv5U29+2IcAyOmy+HaN4yR5cjtNv3xk
0YrbbqCQ+UUMpV/3IBDM8Ph3kXkcQAYBzxaNwYG2rynL+5+ZLLqj8lHa9Q7OCwj5wf8yDk00N8qC
rjoEQiwV7eurayASqkRETJAd5fWMI4nuduJ7fnYkw56cvj8n+4PaPQwQgAn4MC7MXd/hjnG7tcsL
k9+mDqmtkyDbgUkKyseKvGoTF+SeyXGHtSRzWxFYumm2K0P1oTp8LW3F5nFD7hzOB8j6H5OFkoca
rnlZJRQdCuBKf7WMHZT7oZDb1ZCtjzQ/q/WaBOJGZw+zZizRr51DNEtkVFD6OaSq6145DA6SqZEk
1PMyEdbPFW4JYhJjueg7ZMiZMZrvUGmC6+yXgJbwHMXV1sAZe5N7RW9jAX8ASMbT9eJmQcjlqyW1
zaOz2HqmICAPBaSluurHTv4MMOx+esoWvJ+9XTsLqFhCwKCkhgpOLGzVSpns/j6ciB9KKShAI+/A
tUl873pSF/EXkaSY6pp71+d29UVkJGTVdudmfvSUZ20TDklkicCTc4u5/jEMYFqmJf1WlGKml89M
RKZrQGn0Pvvt95UTTSrFrZnklR8064FpfcFVZWf9JEKIJf8ZMmxk5YLYifZxN9eV0waVHCjSzsVP
fi0quliAe5MVX/tcmmLdKY4vqHn3y/tm/OOcy6KTO+GTQ7RtkFzYOQhTrJYtgRlTNtEbwCtiI/OT
kSOfUkDtk4X1dDjtZqXSrpC2f+askftlXsO9QnRExNzyTgIc7pK/Ka1x7zbhldPaFA6Bu9l72TGd
OkdEuLjmBcjtpdn/g1kjcmjmbrugppk1q/cqoZagO6B4UxFfljDIU4ZXlyRCgWamTYMMMxsdpPDs
3B0bKo1n12lh+HTyj8aIR0uXRlQQhHZdQBgEycTK4JjZZ0QOMGYxpaViop7fVFZ0s/m7DfHcDKDz
jQrKWgrLEW5i3+64OpZ36wDk8uTGs5AOletJee3sY161AFVuwBjllZOlfq/bWuesxg9YSNllz9eX
Ds78+pbJk5KMyZjRAy4bAlUobQ0jlgozaO7Dyb60yHz6FxHTM8kuA4S3AhDXn7+hMJ6+zJUI5FvD
h3uS7MucrAJgIdORVULOB6CBx8IUGnOUp7DwAUlk3jmTRpFVFaZuXU0R/9OL0Ky2jNzwi4HJy2YH
AX43PfLQ9NdK+IaV1W6b4AcmAjEbZaBgayPjaU9HpGq7Ls/Uckn08Dtd2fG1g0rp/ZIjbiRxtcBH
4T+g1zzA/St6TRd50dzwa8XkWi50bJ9zoMKkmD2k5cqb7EuAZVCGiXa6DTms+4k5R+gthxhIirgy
BL2v3sEgiPJLQEGyrNwhU3GHCPjD7SBlwtI9E+qclYN4hZdsfUbNNAndpYkLb27xV67tGJi/Uc6Y
cMiP5LtO6IlLETKhpwo5X4Ixz/X8VChnn5tOCMG6QX8CFqUbTc4iwvsBxYLYSwlULR+MyvnVXN9F
vFtzDjVzF/3nllfPJ7WvGCOwaVwr7338/iwBx85uGgxoxxIoI1BxcLYM0Kt9wQDBDFkEIqePDDGj
+1utUIOpwMMXnWlVG8cGUhGP9m+ZVpSEPtMw0MbuB1WlBh3B3TvF7RKXEvknF7NK6Cr31Tcr8I0n
GD12sl7XKGKCyGy96S5HmqNNbTBfWIviMlb5fpv5CNOW6sOwGRKccG7y5cuRSryHK4MoLI9s2Smu
2y4b/zndaVQED8GatBLUty9k+lXoKcxEdkFTMiBbd0bsFWgAbtgiOaqm6DIeuPBPKZ2Wcp3EaEBN
xcCOZI3sYNGUILijLfwCMoMuFbpF+8IgRmzWzoxmc5KizulM3QR1OZ0bNbBKs9mMMhQQsYDUkcvW
1nuHZ/QUHZIETfnMzc7zudAw5Hpne301qeMIpMvJZx9vMO4jgUgNplvPZJxolKzkjXBVHZ+qNlXb
o6r/CjH+Tv9AxLRGtI6HXmEUW0MkpnR27FXHc9cBrn5qY8eTo/Mbx9e2GB5NP4Yk248r4LKxujK9
4x+K8Zx4mRzU4f0LP2uRz9Oy73GNAULNBxQ0Y0Nk+jNpQeOQa4gaya8hJURvWFtt/a55rCBpzom+
lSnI8Dk8IcwzDLD4RKigQpc82ya92VFGNpzVsevCmPGuohLozBjLIyJ/2C4FvR5+mjzMH/SZgm9k
hzyQlyZOKZCo+up5g5obw/3sxrZr4pdDfOQok6aDRmWtZcxOq/lURlL6apCTRch0RrGNNCd3l1Wz
PRhXUnVE9sHcNXBUM+J4+WWHoqGIf69C7AuauLDytXmGwpiY64Lr/8BmRlOAng+bQ/jjPCDXNAMx
j+OLU1AB1+1Dg6CT6DZCVJxOOAhv5/wf8g5odSmqPS2aXOzEORSxQFw5z+f5KWgrhE67yFI8QGYr
Xe/NmUHIqAm8bUe6r/71TmGTOhR7mRB1UdPncng+39V7VHZOMTGBr2Av1JGlU6Rc3G9BnSJSCQlT
/ztCjUwAMrs9lhOBZin01TStABK+RAJ6Btr9deYsoRJeNbAxwidQoPwh1IhQhlIgxM56BWS3yjsq
QzktYXUslVYka99XkYZwFG3WKUF3e529yrMG4hJC6V1HybfbVK1OtUTd8BIXkEPxqt4MAuCl/CeK
9+WA2kmQptGWEKrxesXWsNWFC4mUZ/Fjk7+NhvZ9ZMe/4duU2LmIExyGX4cBsEASw8MKgxVy6V6/
bsYO1g8TNdL4/Efujl8z+5N4cdbB91CGla90/myhxXi6Q4jDnroacgJL5jTHIesSNcxLuGlghQDZ
199lTkEazRjNNhO7yC1lnxT8XRr0rxM6R6alqqMI0eM3/fY3jD5dFJo853zao18xq8sOKntePhZ9
lFrkagyM8Q/bkuUloi7yZRmJvtl5x00jyYf5GhjUcD/6FTi3liF8kdKbOg6SdGRhwY2bAHQVH2x4
F+l4+JEGOZ/d+CThpmw3Yfb9ZOoS3qGX73gvXGA85Khe852GNK2tIDr8OHjjm6YCmNsDgKcr2u+3
tcWxV2ivHltuUJcLOzxdzBJ72Zlls74FEKulPL/cgPkDhxwvoevqEAEJWqjQgfn0DPlI0RUjlusY
lKCvkYI3oxHOvahSQKBuRrd4NJJS9yuG8Zd5aWnO4Yu5BMzMntMd+HHYsyS6tCzFSI2FBLzYrCF7
t/cAXfhk01cDIgNQ1Y7XTUG+4AtTR0jYXott2eeFw3pMqGQ7BwFBzBiqUuYt6ZeNWgQejmYwSrUC
0zbaGXvXGoiYFG/76U9UdBDSZwvjP0O+JKDF7O9CBibDCYs0TFw0go/3RMrw0RSlNVcgo0D5Wjb7
xtUT3kQP3RkYAr1rUycmCoWKCTH1SGQaI0XI4tcUcjcjn68QgxStvEdtvlYCXjAe/ZijTSvICGJL
rAw0oMwG3837zizrV6Dhhh9ON+hZ/c6zwym1eYcgjTHG12/rIYmENwnY+wUw/BDrcaQ3oS+Chbi+
yPrCpPPUlcerDVrwRfAq6jkWyplTIARO/04fgSUfN1qIE2f+vb6czwUKdb2wnpNhPfFkh9BTBbrk
+Iu6iCxczbxMyxlfZNKrYuL7NjeNGOtbbNbgXOpvAOP8u4z++N6OJ9fgV5izTw1fToGBir9Gavoz
BO8g609+gYBa0/sj8qfSM6iCgMcCJoH7wHx3XNlRDuYUhBXCweOTqPMVd7K0zXql/JHVjvAV+bH7
1lyAcKae73MVlkpSxn3CO7BUiXV/o6obMRlO3N1A6B29ChN61n87wkwhuQ1xu7IQ8PjhFkmPKiE4
x+ER56W4eCUa50nYm5cE0IrTscq6OERfLw9Omh0C3+gQzBW9+s6R44VQgwTFdAg2FwScoY8s4flS
3BNbA1Wqw/PNzwgOflF0A6kzvipOm47YlpvX0E4D91W+BFX4Hq+bJ7Kv7Cj5EciJ/sSCXqt88DLI
rciG8DM7fjptTbv/rzSizfMoEozWTwffpHFVbzOQjrGbTjOByOLuVShkD9NCp8x9fPhcS35qVrh+
kEVGgN+rAaZGyKFC+/bOv9/u+IHYhhpQlSty2J1cD0JB/teR2lUx/JLu9bwPs44ttEJ4sIavcPVG
pdONpAyoZLJw66/nv/ZHeHulnfUwvcpt6Yz70xwe450dpoie1axeQClIezXkLgxzayKJwCDqMpGL
zUDdO/mWmaAn2eHYWHiTEcm0OJjYQzzp9qfdO5ibLl9H5ONCz4a3hy57r42MXZTPdWbYfbDGftfh
/ZXG/43j/KCxBjUEf22Vjw9ce1+p+0xlPqbOiXn8SCM2UDVpqOB6yWe6MAegt2HuRczq4LETWa7z
De7IKdhnXbCQI7/vbjbQYHG0krDdBrpleafuIbFODuNOPd67Qdk/aDSe5ehtBm06J/G2dqMdQZYf
k3tovjG0gsU2VPdylxP2p82I2GvZWLHpZmZkPA13fMG8IGrhkN3df80BoNgHvBRsGro9/M49pZrU
hHrm1tnb5FlzWpk2C8RTwXs36+ozgEto2maUjznj6+8PLPDsu1uv/NgQzzZKFgTE5LqRQdSWhqry
ywNqsJgU/FKD5nssNy1GjiIX/BnJZVpC1KHu5o4Sl4bHzBT4fy8BgQYkEwiX0r+uF0Uyhivju8Rz
yRObNwGDYsCrDsSKxZYxIGP/MmkaD9f+W/R2bfFt63/gr7ZSj2wg69Lbt+sxRyi71amyb2kQ4QzU
OH2qbB70k/JaTfkJQIFxr0MQDnHD/wc8VXHC2NfOnY4jjiVIqQT/dYRqmV+1w6hM7M4qHb1QuxFS
xVJFxhjqVTUP1sztK1huD+mYd13OzkfoOaFDvojMkdYO8ABdCauRx1FtaHJNHsBET8vhAcp3J9Hl
1IH0tTyPT0bz6VizEyJH8EuUulH1q8azU89gCRvShPM6x0cqDnz2WI4nBszqmt8dDS7JEkJVeLD5
QerebVmMCEhYr/X41vzCgRT5La5LxyZWqZbxt9vb+NltkWxz300yJOvChZuhEX+bQOzVuc90k62l
fdudBBkCJ2pTL13OWOKkmhiwx9ySJP+HeaTSsbRP7XG45dY1b6RUlnw5Kvp+7zCUqb+iUWOjBVSG
qmmDB83AypFSHZg3SXm2XaH45blnZYVgI8i628xy8psDUugXuFWI08MqdOjF5+dD8gV8IltNOrUW
9Hyv+Gqnvo4Jkxt3/OtUmmAjXope0ubGTJhtix24KKDierTEgeWo89/LzIPmzPquz45exPsFUBdf
IXergNHaO3oHqR12qhQR7gFwth1m35lABF2rnEGo9WOwEalo4QqmDFUZUC5OGFkL4h7NcoCOGsM0
byMOfeMIqoTqcNwTCTa/dVlVqPFppuidz1ODIWAclegZoJJSw1X4SVnvDAeeZOC5xlTDzvoKBU7i
pm9FP5QazgnK6KiBPwG3lM19ViGOtBP8QzbRdvhykLWVs0Fw8RpPGESPY1F5dGSP4KzX9htklwqn
zvMx5WhQa3yzPVk3BpAK8B1xM3pG5OYfhjFDnPSu4kCh3iiRB7TDuPHtjAJUi1DtYPnQE3iV3p1o
0b8+/zojhbTIBLy6DBJB1tL1rCtOQJLNZbSFFeX39lh79R0LmtBBm+oUgCf4Za97FAU0dZIIlYQu
oXzQ3Wf4KADwC8MQLYXesHyLBAapHB+E2KXsubGHrI/ao5cA3VGBQ3PhTxUSA6LFXAtk8gGDFydW
SXr5tm70MsuYohONsyl9CD8eErReINnGu8SR8V4QdTK65AZa9YpSmYzmbPx5+Qc7WmHptVZUTrTt
RWM/aXSz7Yi5ycLD+Zzn4IkoQv3iVX0Xu0qaApbgGNxFx64IK34JfyDfvDvZhTkWCeCTeXtP90o4
JGLSSDRAkPHGKT2bVkmshxTSKxL1f/qtTmXhcX9yPjJ0v5rntenTNPOXGz2l3BKGheTQzc6ZuvsQ
IqqYAv89NMJ81GNwtF+1RSbFKMPPAn7AHGqfof8x19M1wcksmNzSTFaW7RK+1JgnYfVJMuoDx7DZ
54JgdeWpvtQhviS3xmmofuxye1hyivDh7QWTzG7wojlDjWdXMdHfZUjH8K8oIxx43s7eNHMPjZvT
eFGrfAapDr5mu4Iy3E58YR/9YBw20kzydJUwC8PJVE4eKurmjxmtfzE6eHusMBmyb2qPQQ+5ASIF
qStU9E8j/6NjxR9TytpUGMSsMOjMHYHhWfzoJvwdMQEnxvqxXtWnVTMEle4NiycNxl/eiuyH29/e
zBCcLtrGfh79WGm0y9T8BG6whaZHXd/2xezLk4n91i6X9/+4qOXtchJtC2mtg/bwbw5nkAYGyZ+/
IoIrWNiJKHIBYmaCbkoSMXqa3mKrhavuhwW72L+Zb8I58yrU+970ZIjD6YEpjM+jimGo5i/5omRB
LduD8BqYlL17MGryk2P9KY+wsb+Rz2iBpA1HELqmNwSjyEN9PzOeJW2mRH6p3HCeEGr/L7bFxuf7
rVqpyTV3sc6+vQcutI5aBUj6W0bPDdHsyhipK5mqcBC5LE+aLQI2bS0tsLVZCJT3zMrVNa8FTiWS
QdPswRlaNw+3Od+AGd90lyYzS6M67i5MhCb3yeH3ZE42N6FCeXXSYcAcuLaZ1yVuBlAJ+LMeG51l
ysBXEURIvk9JyzWmcftNJ8a1ikJJDsAnUFYuonbiNGUNa5w+fjnNAneUF1tPk01+VmJJJ0S0qBUx
XyBpX6NKdvpZdkGeyrikhy/JZ9BINhnIBxjrhODTflVpoY7myJgJFqf0SjY98nhLxCiGHd6FNod3
i1v7LaJ3Ug4hEcQ1U1K8+hSXuMEnlR2tVaK0TCUV7vCjWsdp7Anf+7x4eqU2Fq6Csbjs2//+DmeX
8HCbEY1Kt+5ukdZAh/VuYmeZAFGsXBcIT7SNmIoefn2rS6+e7/qwXR+razL8YQg7ufHBlNmWUC5k
+5yYWCBV3nDssX5fwOo3f5/po1igHo/9fnfTffwnIGGxrLjjax9Tu9gU3ETtuJy77dGlMuDKFJ1j
XvBREi0Uc5CIXerRIofwDhakyMgGkdjQn0RV7GzAMG2hB0Rl+cM2imYm07zk0te552jXWNlU+YS5
dgIe9AtapzbYO7QUAREVB4Vma/vl/Lh83ZYxJ5rEQS4pZbzESZZZaDq6KrQUYKCspJzSga81C1I4
dLA2J6L89QDMYT0Q/DDdZ7gFCf+XwEE4Fa1oEe95HJ5H6RSHWNM8t3w7CEmHf8PFIe9rHWQBHiCW
9a+StzXgTX4ATQS13TOlr+uouIsCmgKIfSRJTAsiXn5ozNYeVtDV7829lTkY3RKRGWXJRzfuDYxQ
XeYOXjsr4SqaoZ6tCljPP9umX+zh/sACU/9rJ/mGy6Ee82TH766SQGBpy1yoCM3jGKveTtuf179d
0cdVF+8pGPnpElfQUqcrczk3GE8vUf9cr4KGN4s84Asc+uDR1RVd8VLaM4ZJOdgaMTi2SeHczAXF
ahwOJFUqBXK4z0PaIFwnMDhniLm9eYMIs8eKBwIxCvlWe6uFFaTbe9gcsq4h8MVrm1InVZyvPoKS
1UEv4bKWZtVJ1khTsMap/x/a1vrRlkPpKaW6zRP4y+C4g3zcRdtFXfZ2XV2in+Nb4YsDyaTtSzX4
pEwMygU3aQi0TrTufIQrS4nBYpJMEz9kj/iErFYqzB6JAWfyMbX1iY4xcPpENKxKbqnxiPGlDhhV
t3E+xaiFazSg6qNMFRfeZeEl4wHu5fuEgtEfO1UL+Gr3le4vmjJv3kbDODGJrSvPUgRsA6dKqlq7
MFXzuHVGRyYK5BtedLoHTtUDVk7zzqiBUwkx5GylGCR9XiXTNV49ynkH5o0u1aDkQMqWzoM1JPIt
KIbtLco+FhUJZdYIY/MZ7zk8+uHZslKs4fOUrH9KmH6U4bytVwg/qFCmlxQhTUKfzCyNY2kyWggv
N2W62/6UZ9qHTIWiKNoLVqSduMd64qDLEDBRQNzVQx0K7V9rmkV6pzi9j/r1j8Ct9bqodLFuNo3f
Ieurme0p669l1nLu9yIlzVFz9aU3FizTbzyU+zOWJMg7z1mRAuO4kSua53TFbNvvA3gXTVX51mJL
vflMs2qt3KVg6uqREDV+O72oKMY9eZqcmzFfe08JzqJhfYFVJF8Ftp598gaf3xRdJqgERlTAwUta
5w75Ze3Wamzh6XwUFL3cxOJM1NmS6eXASi0SRjMHOjFX6zb+90uXJwTwdNZ5zA5I5ePLYhnEX5fK
KG0JC9sUlt53M6ugNRlPD79e28vS6U6hcLKRQgcPBBQxcJPi6mcH5uaEbUgxR2FvcBQDMbgqaIQq
72kn9AqMEdu4yLOqJaLrj/DIhDgr0X/e4a3p5he+hVabCv/xrgzMgF9KKfYzwJlsZL2bi7+Me8WU
3o1ZWOeZj27z8FALRtGSwmb0vWHULgTdSVvhOvIJoGSNiJb2a22kj3/AmHp/OvUHa401qEcJVmZ/
iDahM+zH2oQu2bLY4rqMHGWZ3jQiGXARPTqnRZtC26CorSootnc9S2AaaPn5Zrb0koMUQYN8j71o
HeJfW0Z4XwvCQtnfDzBO9eTttUH3/qmXR79jH7+3sZM8YK1+ON7SvmB4Jf5JS/ggvBwtvqKMbfXr
WvnwssOBo1SvSWgyOda08oG+J2T/yaaf5RHNBX/kgWwmRy22fTTRRQBky8Pb7y9V7jKSFjdi3SEM
z5cXaDQGi1xfVTUt8EmgNVlf89sbdJ1JkNyUzNfiwGazPt7JZZ14WBTa+wXoK31DTaTlqHjbD+IY
jlB31NRUVdewOkw/TrsUMCX1V1N9ypSdGp7wWAqnDDCgP071S4O4tu30fpxwkK50Ie7c37gl8ZwT
PRnQdI8zUNvYNmO03nDTxs07X6evkt+dy0M0Lh7CqVPNXAYiYbQ48WAfmAeFfikbTyc9zD5rw5ol
7yCOyGott4R6UySosf0QJtdVWGhYoEZ5coauXZMifx0hb6i3JllBVvUn6qplWI1cmX1/UmU0XBUw
NKgGaFJTCRhnzvVCLoGi50UgAeQTsA01MWm+eTG/SZ+bQUFAhrZUIAa5ApS95pVoWlZppzcdviK8
obM8aOBA2J66yzFICuG3x6b95jhtGUPi8ndwW5tRHLTMSUMIOrpItjAMviDUvHC2cBx/BHkh9Md0
0P9EkOYKcrPmvR0zjOYj2+44qXh/WREhDO5sf9PkGYyqbrFvHwjPGtehaMLoXR1qTVu6MTeYbASD
QYrK10xIG6KMqwlDPxX5UsTzG+X2WVUHPskubJgojJEJrtCv1lUpi+foh9s9BgjMPWUpg9Q3f8q+
T5qetjFWWLqq2H2yhI3ZSaa9FWNoHTKfPuQpDzZS9hA9ksip3+K2N17KC3rVBtweDi9rMdJq66a4
ZIeQo9hz30CqNWQ80niw24zUyO+LdEI/ZT1yjk8Y/rTS7La3L2rMRB/wLrNxjXoTH+LcH4m7g+rS
ATM7vSzz6Wh9xYXWfBxxbQBmpb0tMnKSCbKAfCXK/Hl8hW7m9Va1UMoajKKcxdCSgzQmE3rlSw7i
VWw+EwlcZil2gksjnl7IFcXjgzEuTyEOmUMA/PSTp9iA8lUTQ36zaANZKIXWOs+HruFXtJTkfhbW
LnaH0viZC2xAXqe3DIYLM1SuxWHAjja0pBHpNY1bY0U6WoILAEwxP12MEzx6Q9wrNUyOWWikYOGN
ctgZ9o90fp0MIzs7uG1yAuTuO+QjbQLhuCX3GJSQlk+p3qoEacjYasbV5gW7B8wkGZNp+AQ6qK3s
WO9lQ4mX1lIyZLmv2EExCj/a+GQStOVwDgTKkBDPiwzMDwI76uNDlUGRLCZDZ2aCJbqjFsEj/K0x
txt/K+Q4dm95gjYFcjr7nHg+B0Xhs+1knOjY09K+Yx2va3fPj7XIqegheNlsxnYLSWpZUBR/qq2m
LFFzyoYA/yAjtODIxLZRg6BrxFDFeVUG6xyl3NI12xl80PfYmw7QjENvKofBbfgq9toHyyPmaMUC
JgR3lzhXt8Ys/Mw6K1eTjIGgV/wsSFRLA2uu/AfDfw4MNkiPGnaOdwL1BXf8TJuELP6MUaTEYz7Y
0+yFAsrikrslco4j0OslmatBGDJIrYmqVeBUVhZpW/ipnX7JhITu9brRacdOvrsVTQlUmUHl3M16
q6hDYdXONKRS+m0F4Ozul+9oRkeIObtT4rhXOvR3Sa5dqd4qPbuDDhD6U3dE8fNJlLFN1P/k8jBK
Fzvz8oo1yZntOEgFZEa6Yk0ALMEGdS/JVaPKFVrLfb+Hu9PMp8+wrUCw4cHm0ijjRi7N7/4008hd
y6XxuCF+ie/fCb/ZeZ+k1tpIR3U91v6TNF7N86eUEF5PL1YF31gwhqL0zwTMm+ASAY7tr+oh0EvP
K5x3iFi2PooulKbtjZqJZWwFJVVZAIoE9x3DhC6W2ujnT7sq73g+suqszC/YHWxLUdzUM1G0+q/c
fvFoyOpSDpcYIhgDtekLfItz1W3XjCM4CN/R2p4j4dGgU9TNiLjg/zlglLHXqnubgo99cp/iqjp1
M1qANVu06zltOtzJEW4PjccGfQf/9lY13kFp2Hadtz5oHBUZoktARbdSlS9aBgP81slbHdagPXhD
AVb0/Kz8ELfmbc//7uJCKA7MnkjuSTcfZBMjQSS+qmssftHuQZeEFSMJhusrTXK6T55a25d12O5P
V1PQfORe9b7BoaR+dGqGYi3wtBfNdo6Hvqb2yzQl0ubGt17/l7mEzNicoFUSwoVS3d2GFfV2/kWO
3PBKb5H5vLbmkQG8kQNizv79yoS6LOd3QXrYcyT/wcVk51iC0mlt1sivONX3JZYS7gNWEaygrTUF
LOWcVPRHtcljn+qcpVcd8cVozDtngcSyBVFggL63aOO+Vy8/EYPIuHWG3NyGR11vU2udCsT4xeng
osuayQFl/+LpLWrGLL8OCBcv1oyPjSQTpwiUFeZ6PyoL43x/zRrG3diTNvLJalWoImHVfU8X4gAz
amT+3DhRCk/r0KTFl0T0WlrI3uAatvtghhjZFCZHA4SzO6jVJQjgRHNFgp1Xs9oCETSOf5PnnaR2
7ZrvXqbh0terc8yPqfUQwjVUq4s/vZkqRp1q9ZWYACnUfA9iyHB4gQe7XYKLxuhqkUc6UheNSHNc
+jKnx+/iXGVObvcZQto5+aezxfHv8+yVSxwIi6JdHhBUPUD8eIWiYi7BEIAfDS3d+Z1en4XIyfKq
cW0IEEo0BLJkljAk76RAOmzYQy+/gA58iugrdTCYQHlTEQB/xeJRxaniBlNmWXMaowUBnM4rBNZo
5orw6uLP8UL3V1h7XrGywpZvHTO2Nz7Jubp8vCF7FKBeCHO9fBI1e2BhHChzqZy+YYu1+Qvi3ey+
tNypIvfE6ggOSTEQaO2d2XU090lKzayfPHniyWlbLQ6fzKAWmKoroVfS/Y4RpG+g0pDSFLw5ZT9O
sEswy18bpiAhW1R1Vlcg9Fs7tiNYVxf27ZGVwGKLSPdmGrv5qCX62fpKuXtM8IkKSlLjmY+7H0Mz
afoYB5OwCa0S1YMEKN5g4L7eLTiIleuLdHCsJI4R1rnfcUKKTt82X8Q64sxtow69rIfxBIq0q0ay
LGwSEDlcc0sWsxIiaBdp2lTQdF/909q+zJJzf1G8oXoRTglua4v+IMg14lroestCFSSsMGG5qziv
wyexp9yBhe/bBZVI4tSDZetPFRREUNltUAox2N7hXZxsWkZ1qcKOkiMg15BZu5cur0jdU0LRbj5P
2SA0ZeoTUy7aOFj1jKYocC2nLxeog0AyNSx7HH3sBL/T9HN0OyjPjfnldkQ78NVloeoVSWMdHF/k
ElUYLN8FR4uSIAtYPnEB3UQsZ/EvMkRbGa+jb3q7BVmYd2kComBjo3UYzl/NkHYPjfduD9JL/HYL
tss4z+ckXuXlkNKDPBZ18oqPLDZ7cztUKRtvv4HCK41kEmWW6CyaMksjQgwPV3NXOPVOsmh08Ppo
39ruQVXyuIyyho/wWSZ5FXecnMQlQwBb9y4VGZjsy574l33v5Pv2O5tvGtDU8YdqubxmFxuG/Mrx
2XV19ohOJHFIeA9QPR8dG46g58wjc8Iz8bmdDYVRQlfii3EHRHSlSzu148dXBObxgo6m1hW7tDXB
q4E7RPfAK6eFEM7DpkRkgU5qjD+/Pf/kOPa95NbqbpmikIiBJSmhdhw9p9S85VaueVE9PxkW/fJ/
rVMgTCIzVxEjcWOeeOwVHlp12c6j+BhguWdyPhUsNHDxCBApIwxJPvVT3frJutvgCv/eYAjuMYt6
30YC5ewYVCEtp01B+qKlONFcKD9fuu2dwj8pM+FwAtV0Efs3WFsGpiI8be/+wFTF0nCU8ps4ozUh
YWIlvzaKC2X71GqmaHyLjnhqaJCSXQ4iZl+wsJwYQQCxxaemzvP2hZJ4H5mc8b1ISbipD2r8a6SQ
NalbLxkIGdOTNmdsUPtGNU3CDYy/IFOYDHds8Ae2hr8DS5ZHHWKl5dYGm7jupjGknddxPxEWVSWz
47pQLbepw9NIhB86fCbyok5ovU+wtot05XzfNyz7YfIbuClGZkQLli/r6grnRPzmJF+w5npQbnIm
Y1X3Vq3YED75psQvq5p+98urt6z0YBlf0NkdBEuH5hozYUk1HBnKFVILj5pi78+EpAKWeouXrQ2u
wzYBlytL+CcjPm0tmEL85rk7slT13fyhGsCLlg2F4FyLGXKwLLqp4VHIzLWuCXJIv53k4ad+TWUH
S70eLh/Zt95rATE+7xmt6O6XHHOmCCxI+mcRwyaWJUljgt33DczeGwYsTOv6au5LBVvGknB7bqbH
WGHG44tYEERK3k66QHq2h360zJ2pRorYvxWk9uigCCIDUR7f1uvBuMNBgrsM/mRpmHjPRKxMZ28h
ddm8rnRiRCMWK0awVzLXAePwoLzoK07afSo7cr0uMKV9XRpvO36y3ysFTMWN+gquCrZ5OfrIIthV
JRcb1xnYIuKw44AsgGmLn36L5ZKFcGkUMTA1Z66RJIw7BBKhzjgiHY0LvgQakyNnC/fXbQMSitto
vLkiKEaqcDdeR3RG8qN/6NS/HmKpx8r2Q86ThYp6TBFJBghI9S691r6R1LQ64nwOrp4UaNoaHkxT
5V7JVEBWG+rO26cTeP8QnvOA3Icw80eLNl0ooI7gnDhjZd+1akJQmaS0Qi0/qTt4V/0rPLrQ0zuG
35iLg9E+aB3hFR69+8Ux3P6oJWyX2aFATyCDKpQ6s5gP2Xgb+NbAjWl1R+x6eZYp4r7wXFsi7F9L
WFvFK9+P3ikNFhPmwcXIvEHSYa/AcfgiVx+EJRJSTatV5etMigPQ2k0DzlYdo5zYEV3+n5T0syHi
j5tcl44iv2r13XLebswO8H5sUrpw4TPQRwkyC07T7L97yeD1Sx4DkFTlLmYwof/hhKoC8L0uHv25
LCtrTL64ZLPOiflEx2BUbTf41/U32Amsg0dmViwbA1JKm71k322PAtafSG9hAPgDo9f4APKAl5Q1
XWT1gDtspIFGy/MUJHX7To0Tp1Etj7maNsBY27H6HJucEbAoabIW4/fkRt6MLnmosZMMh3oUolar
dcYKxrkdo0OGsb+w8+8kDEKdQdMCeAs9o8tQ1U0nxmzjmxjyQvPh5e+/wD/XT5ZFS2VQkAUk1ucq
ZyFdoXDHjm25YQSLshywNdMZ+Ip0gQO+GfTgtp33qdD2wONZry8xeL6AaNhOxhXwcFI6Hjs3pkR1
mvp6S6f7mIbt2udfITsBI76PFdjzpy8Vc59UXV+EanG/YI3J4bGFrCZ9btqjPGx1A5qLXETpbFkb
Bx1A1cNZ12BHyg8eiyO7U8H88BopU1DtyqEWBgCeZUBReTRp3QVq8Y7GOJrLCNqVVRp0xKKDTwVR
Da8i/AsPbn3mdPaLgbXpuhs6I6UPnSp0eM9P0Q5MoFVo71ktsQZqQA/CFlPq+LPwCcNjGmW4vgFP
wtYVa5RRHqv6zr5ACWlN/56d+0PvNKfUieJLCV4TehQjRojxpKae2A/Voqhybz7x/dZ+EsUCiz2W
/2R3M9ED8YX2j7p+m8tM9DE8tR/i7FdANAgXVdoUOAd5k1IbSKItEBVHlftQBOZ5EBaiYbgWuhCo
Z1EfaXAKs5ixTegapv4/w3j9UwdoHrj1tvIsJoCDA/pQLV3QGKBi4OlI6b8MzLgZV+Ib6nz90fhO
/L6DZpzjQjljM56wDq5ukOT+kR/UWB6eHg/12EAUF5qGVtZEdEpd3VYwfATS/bNLzbghfvONbopk
pJ7x79Pdy9Gee6CVaqmKvaS85C2wETwzOg9R1qwW+CFsOFriRhapLVhopoRkgzROF/4wZEE/XjEO
zvPyOWD/xAqyRl3hhtBS6sSrpFzdFuL37LNb8LsSMU5SHC8G1ZaK9o+LshN+WFhxjY5VSHx+GVNI
e1YrIPBdjqlkRC/bBAlCT7xXh6MPpuxr0y7aKM0IgtseQdent7TzWZiIZVngobFGBvAZoIhEd+5O
PHV5aV0ptRdX1QHvveJGXXLHkJmLUfkM5rYcc534IlxRdpzwldsCsqSbT8ozeT6itfHw6KpYE8lV
lnqHFsZpljLVX3pzUz8RmVusq0iengoKoLM3/9kzaFx7dIAqTlmoi+DMadWzLpQ+2jKxNVwMg1lP
XdLvvkNypFJlerQCGPoTcHG3pRVIjO1nfLj7lBtwQde75NLd2kmf0UtOXjF03Z9I9fjb96vyNycw
9qxv2D61W1Mi+VSvIjf5FUVl0Rdirlb9cOX1+9VRawrg4R21fIsM8/7YV2QIU/lTZu7oCGDAiOvL
1ba6RM6Blvc3VKVUSD3Jn1o6ZNl3E1/jwQQ4JyBr7GAO+kbNoR/fGFfErhPA39egbJ8ZzM2hA1QY
XawpSOAcg5rW+p6xQ1B7xH+AztUIjCxBmXPEZDkgmtfQm+AJHLsWRivhOqhghrfzoDsBr9kI65oA
ttWYPnBoUG96dLuWexqbqLeQlUswXeJSrqoKSEQglO0XXKkGI0IV/icFRpjBvtQt6sbk/IkuY0d1
YN6pIT6I3y6SbcRyzmM8Xjn30NuZqpedNZZWS8d69/J67JaUA9vLuIPvGqBPLI6Y6KC+zIV17iue
rs04Owzj9KOMwVWmkgcrlAdteJQHeKN2/RpBj1wisUTVqcSCh3FiWC9N+r8y9BS+er2+v8DZOUSj
+f6gr5aDyVxYDhtnSnuRw9v3/KPl211KXoK8uilUadnRp9owruJhgx5m/GOqYWNjmOf/XZ0QYFvn
4alAa7S9EjdGzMLjvKjxgW33RtnTnyqG967ot9TKxGKSRZS5CkSXEZ7bJer5IrsyfjPFTbThx2h1
QsOUc+wFGqtk7LEU23+B0uEQwcKmQv8id4cIlFkqxPHCoF98xnKssjLH1UR/dThfRCmrF0JsGgrz
+9//BMARcyCN5iNLhJmRFgFXC/DYFTye66TahzV+6uR6Z1k709wPQKFXX8vdJzpn8013dHjhv9+T
g8BrBhISJva3Pdgnort/qW8miHNNXw8/FurLZOX5mmjIJytNvyPcyzSLubHLZTKz9J6l0rowwNl8
CZ/t5ez3l/uipInGGdwayBQ0ZhwmAXrbeHxxW84f0iP78UIC79shnw7hctQcGo1+vH4aIIwREYWq
ScRCtt///+vAzbdrd8a2cI9KToeZFanj64He/r0ZltG7eTpedMCLxwnmWIVgF9XOD95iFwI3KexA
r1plUdKPwbJ4PBswKWGLsGybQn6LkoxN5zM8rw+f+uvE/hjRZK9ycaBndNdIPA9RtL2zkd9rrxDS
XkomeN02Hx1O+0feb1K0Q4JxN1dYmJ42PInCJwznyDJVRbJ+AWllt9Yk4WRMXnZqjWxIKorUhUOf
u/M9WiQ/D7t7dTn40HR3HD8WCR66zl7KftR+yBTfWkycplonWE/cuQMDeEXoT0IdpwuQVm9cwAKQ
JjtAJJwn649h1lflQKjgxwraJlr5qlnc1IzA5hQQvzbU08ao5AwOjJcPOgbGUx7Rv8S4MkrYuHvU
G/pEE0mXYT5qQXTwJWI2so5HLHqpOMU1hj33rB5qeRqJlQuz5zF1TkTtl+nCy0yJ6APx4d8UYl+D
0708DDHJ4m4RacGaH3gd7ZwSyLa4xqaSVr/3SqdVTeJumBsy1RIoOw7Tr00yp+aNe9lt7Itfajhb
sUFowPbDdi/zXEB16ugP8BXcAIWajHh99dLaG0FUq24G8rAo0HP6hZKwfIqsB7mMTUGIX+b9Rl4I
yet9F8piMBc25P7YjDZCHmyx1yCY2p4TofuEHCUDyarbkKxrboOD7pZzRzE2Zj4E/4rAhm7dQARw
M0CnNDCkEIHfS3x3ldW9MmM0K597C0tJspIJJAvv2cUagIfbBAVogN3gwFIPCUgCQ76uavCHIOGQ
DQ+dNBSiFGm1B+XKpzrzCNvirYY9FmLEKaf8qOuKKfNwvkWCJ3Hy033BDwn716WaP55fKPa5MpYB
OTTYgF2kc46Vk/mW0Um5GUPVT7CNW58OGitYy+qnr9h6xg2FAF/3hMjrV6IjekWhsCude2NJNGYf
RT/z05xKifPQ68tl92dt9J0BSSFyhXd1UrY1DcA3oZeT3VdLDrnIJDF2rI9nkHXPtnqc67Xn8ozf
GHWmwRwakU7kzZldEFCajPRohi50CmIlqDfrZdvr7NCv1F8BB3M397YSK9U0Fp7g7s++a2oLWcjX
beRUXxpx/aIxbp1fuVKs2u43wKCjsJlOr272z1A/9jjq4JKk5zViAqdOczkf02+lhEp4iaTyOekf
al6Sx5XvqFe7GKxZefRebqASlCTB/XmWAnvAmvs2HfOc8R1iL0X7rxQ7xEQcyg29KXnG5AGYao7/
bWdAyAysgKcwscFhL6SYn65JI8X/ZrHIHSMyjoIWZeT6PPefctX5U7VeWDtprpBFwQJC6CRWugQr
Kg5RebpqGBQh40u/GQVg7eV0rU0DcA4LHRVrsEFJIpsFcOfNTpktTLMBxHOOKUDMU6MusaAQylv0
CBadrwFukAuRZwro2JKfr5h9ipy8FRi8B8RC3gaVdpPztCnJU8QQoD6N3Gvvgb6ZN8EEKW7qUHIP
yvNOL6fQPa218ubfZEDq7HuTArYEs1lu2y4ZbnTWqeA4njDbflS7La/BC0iFGma0/W4cN/LnbQxj
zTjJkrh7TxogAHhEZMiHjUBVppWd4D8jbg8jlMagiKkYU7NQsmpdUh2fnXHxKykhgXwWnr0QQm5J
Z5/Rra6H+nxxmJPAMK7DWhfO7yrDmj0p0JYQfGmvgaTyjT6DY031DOuFIxDjRMicQPrn5gh+sAKJ
lezXYtjUnME4MXiSmYuqTbENRGjM3NoX8Hwt0/BrA7LLF7GVnxYksNt2W4IeCk4U/BgWcmoBs6ll
RhUJkXDjRZOcrxQQj1bnwHj6rpOL5FMWQRvZC2o96AGF7Nl7BnwunSX2v/Cz0j0Pc3N+gJhVhT61
9ZqtgY8gbB876eZjbTMbV11CuBzi2jgyvXz5h9YtUDnvu9j0UiyWtMbot1q6vM6SuLFX9AoH1MVY
oExI6v5XNOtqb49hP83tKfEskpQ+ZlfF/XORPZUL2/86UAf3FFM6dmD4rKCthEi1tRsPDingQaba
CrcJZa3jaRvB/mlc7Ml2nZJI8cvQn4JXL+r5hMi1jPPakHjzTka6ZXMZRzGxXK6TPkjEgBSk4EMn
G6sDN/j9Oggh7bOJ6PTRD8eI3HdjG/pAHTOWsGW6ZS1lLv8OMtLDMNDOkDTEyZdAZV/1kDKEYdPl
dpe8YvqXZN6Tx7zLGc4hBXpfvOEMgCrgvaIikAczlvnKJNnge/KSTAMdYgCQWRkhfmK3wSBsqoF2
yDd+5Np4JO2Uk2WtTWnfB2QTVBscq6ttfP9iuQ5esisezyxCXrtPXgAJJjBO9Kh2RyrIum51qt9j
72alcjtli9mxrmLLc3myusApW8wzYDIjIIHZzO1ltqK3+QRe8e2mMb8a68PCFWBnWwLRYBGnYlia
LqzFdKgAyDoPe4pp1zQO12aBbkDraJRCDyB9AGvX0F5S+SLQ94ROiFAVpmV92Rzjmrxc/Ri7NBPm
JcB6R0aRLpetCxXgU4BxuTmK076K2VwtihL9OQwH04Cm/dxg2UNXSiUdSZcoF/eP9KT6sOtrT8O0
4Kfe6yeUokuZJ43UTB5m1rPlcbI+Zzna044SAIzaHrC+zGSt3BuY54yQgN6oLDYJjJWqzoJLQPo/
xz1zUAnW3wBRspLhXQ/kA9+c8hsVi/uO31wLYYF0s8jE6WXf3onH3BV/LrQnKQU85Ibgdpgj1YPk
dW9Cv3/tZo3aCdVwXcYBREktYm0WzXctdrSKX1S+A1NHkvubQg6oINMCXsoy/w7OZ76aWwVgCNci
Vr00kY3TahJ3kPirmG5e9ScagMKDK9k+3PHQ9hsLA6SWuIMODlDZkcBcd9PN5CuD9l6qcT24HZfQ
dx0u8rTshlnk4JnSd9FdRkshUAJOcJK2q13dH/IXkutYfsI1gEtB8tvVj5wJVeuhWxKsN46YBCo3
/Z+0BptBQBedyUiOLLPNtnQYJ9HptX8RXqPGvmThZHLd/tY5wJSygs6XTfcjuP3YIgj3LoUc0loV
qRUKJzRMjT167+6j57vnyUohgRjKQfRmsttoALbx51uL2UnajOuXUtdPaAqY4mUuQqSUokGbDcWJ
qBAtOpMbl6ZMYGlxl1YvsuhRZhe74Glu0rCriEIwMzHesbQ4RPbFjbI6WvNIsWEZay1oqXGcVIWw
Ka6dgTKGj0oj7dYQ3v6o3o11UCeGivjYejWxSqyK+xga1NcGepcWjuFj5Jkc4HKUlGEF4zLofjB2
hh1z9eW/drVqv9TB4Mm08bAVVd67WhRob5V7Y8z05VY/UgD7A4OUrUfnf+1VN3jl3oKPPQnEE/5V
zllBKwkJ6cMBX9CnYCDxskSfItiLe4Ud/OxPmJLe+pLvFpBSVF1sVz0kTKCkt6BWbdBC4CYy6Fkf
0APQpHb2HdUWQ5zgkomms/7udPINY3CxbHiJFchDnVCUopyNS8gPL0CzXypbTb7Az3ZQWQJgJT3w
ys7aA0nd9RrGKV5aHZihHLWlNMZ6OjkHFKLy5sYzxXdgahaOchpZpFFA8CcmrNGuDMqCuC9EeYvJ
XViQe0fnftRBr17tfA4El+vHpQAele+TJp2EtJiOO2/Sz5olKXf0HLPwCxm0j8xtSknXOhXeAzrm
LNMGdRRcIs9T/OMj/5LXiQJ/7LfpxhKMAlqusL14MMMPnZftB85b+1CYEnZMTD67uVLUDnSmApB7
RgwxzfiEh/g4sYkGzLmwmkOgM5FayUIFi7YBR3ZlBJSiWgZpxv1EOL5VdHYwvo0q/udLZDWZ6pIg
7Jb+SX8BL6MsmCTtT2sAdc7UbevOdqXEFYGgq6ZknYqUOZIqHyTLX16loRC+ezxhn0/KfOAzPccr
DnoW8XsVkOPftag0n5MuBk8i2jxhZK9LVDbOXAxgaHKeQ5PsbX41B+V4++/44qg85HkqI9xPW8VN
DEOMQRBf5qMcl3tmXTLm+hkGw2whvLuALkwi3LLzYH7HEdDQo69rFhMHHNojUX6mknYMuHKbMHHw
H5Y0df4EAni/PdqbzMMQ+pzsYJG9tjl9UPwcav1Vxbzueabeg8JyI4ybQe60V1fZnUFI4euSS/gg
dHHToXLVCb5iJp8uJtBZ24YzP5JBjTOwMyXUhob1SLVrfMqgYV6yEeFCU6o3qyS5g8gC2JHa2Uf3
YzsZfJ+ZaHqnXYWgZEyejEnvg/B7Y/NagOc5NAFzAlGHykDGvBfqrZkzLtEGjqA/p7/B/bK57EVT
GjmjFpKvAkr2KiXjsYAvfvCKQWYyn5tWyCBg3amukxCgWYSZkju+rV1v6tNdSd7e86yYu/n+JY/b
xu3TVblTb5DO0ZLi016jp4LPBx1vwM0ecLShAPrnWTUqoAyyva5O3XeZ8AYg1F9MxrHEqlgtGheT
1TrdjW/q8x7bL/yebPsi1uKW5cdQV4ePt0fiocTfBmi/UVjuDKhvJJV2CpKVhPmKYmbJIEi6fpLA
oMLLQ+Jvpw9uAW5GO9nDtnBUubMiNUMzpxheNUQyBBr5I+34Fv7lW41apXe7wE2sAAGcn/PAWGBM
GnSC4ufwNk1ahDnIRIBrFMDxlO0aw+herHNVNi6D7jLyw5zCNvgcgDKj0oaqwr2Rx35vMRJOdswK
jb+0WbH3/Ys1JI9ipuNF5vfmDEbiYnD2KuOxsj91x9EPqd7u97rqnoFmXHW1gwEIxmdFR7uGZtWs
xp9UQmzoqD0fkvbYV74S6zjxbx5eQYs31K1VAoCiW7KLQh0eiEY8aGXb5Z/sdfp1wsEu9nMkysqv
xI1Eq+KQPlIze+rCfUmCJNNxATiophCJ7xGTEU60/9qcjMNk/f6q2ocwmRlLebzJcCx0/ocuQKA1
b13Yf4ZHrvFX9Z5fosSsu6Tzk8uIruPnAETKbg3YtZzb9LRUvDyLGkfc1+MmWcX7JX2msLnQhphY
2HZ2FCqPrwGXEIfgg/x0mlmhqeKH6Zqmb/lSDUVgVQLojogk/BZP3liixttZDl4D9vHy9JmNY7yK
NDkY6RRgrFsq1DKfEC2hWp482pN3AZ6l3zzKyPdv7oNOYJTPPo0foTaOomI0OTHg7zxeKYSWWGbG
w5/pXW+RdZx7//fmTKh3qAsr7INfWA5tVS+MdkLTAm9ENjsBkgtGsfpel8Ovs4nfphFK9qtXqnV8
JXwHNBb/A9isSjz7zbvveoU+eDzANeluEU+bERuTvBc2nhd6YkLNt2ByNjdj0R9WZ/1cI/i4BYKO
0ioD/liY3XiTKIUl3o4SczleIcLSB2GFBFgQQyXFE7s//bnsJzLnutdePooqQQuKDUn+ANqb8bKp
JbwGyosaGIZSfNR0JClxBMobyVBNEA4irP6aLGj+l5Gv3No0tRiTWGYdyo6f4G66vaKp4c2CVBHt
yQjld01GobV3NUMTj60+0rz/TiU7aQzhAA3D94fNqpk468umiqvutqa18vvjzrqmUWp+d1e08TAb
48GyStLvEO1AdNpaddGmyqOHGTpvbfWGwpk1soxeIDjKtYS3lzzhikyMwr93ZFdfLmpiByJGU5Qt
Ug4RmT+j8ugnsRLUZECQ/Td1406TiwhALSgM+mStnPT2fCFBVEOyVanTAmkTwq6dqqh6vdgUwJYx
qpTwqH490vkzDssYzZJgWfiaWmX0o0BKSNU4D5VsFG2v7Tk5+WNa0VxSfBg04twDHnM4+g4JPB9y
AB/xgIjV95tC3LPBRSUTwfAuAK3xVL1sVD5PhUugZbtUnNfc/UDFGEL3dzaHjHpE5RD6jUHO9Nqi
T9tDYkOTQbIH3NoMuuSGKkEFUICN9cLj5AaSFy/IrB31jtm/lyQsF2Z0YpwzxTp4/iIO1u64h+3A
WITgNfMM5XB3z+XV5ZXXWaiESttH3tFqga3NwIBvEk9LIfmJ4HRKRTkY7oekN9rtUS0A7IUKVy/D
gPP7OU04GT7cPj3Dcwey/Rw3OPVa5F1C9XivYsz8ruJzNYZ115g4K3LSqA0dFr8UbxUM1J1Ux/oV
+vxAnExGZPbguwakDYigzBcwHjxi4kFINbMr/S45kXzPpIf5EKJnmx3qtIOHjfFgAe6JtBQSznvn
gKW0CBOYXcemqwW04tPajFcEU8S8cTL3kjcMQpzb+Z0b+5J40bJBONxEDkRtMmv8wSE+bno2btoa
CMbZbDJDqppFCHB/Ck2nIMydcraSEIiHXVV3RXB6EoYorZRxZanp6STxkdo9qPdU7NwAQ8yXvIpb
mkLqKydSl2xs36u8bo72c4ByGZ2zGLPG2rM0WP+aSzXc4RCxURg1S38W41gj/m0GZGboYFs3qK0w
igQL3UHf1vFm9KnBcTqHtwr/GnwV3TxJPIZHNwnDG9Gzcrvz8Ee8IGjHSoZYCa/r9OoaMz+BMmUL
YJO3kBwWErkC2m+VW1U4aNQ38LGKBoGxpqwaPqeqz6VFtGtxpNxg86vaJ0B3K0SMX7BYgzdW6WP6
VtkG4om3T9mwCKprwfEfxjKEZNvrk/KlDwdnP8C80Gv77/zGWO15qWVElLaqBxi0/Nd0MmNZ0F1G
AkJeRVjyqVTSvVe2FRP0gXIlAib7eRYzPaayYaOme/2KXsncAKCN8bKVG7qWTP/bEUf/u5liFeWq
gFbegIhktvO3qcd3BqjA6/wbiTiuo+gol1FH6z0WCqDsien1UfDL9lY85yh+K2zM2cCuH0UkODZI
HHNYzM+3tZsrrCFCA49UFrmcbtMhH1vTB6hag0SbXajMWQSArbNBjAXgMkvD+CAVS+Vom0pt5qcS
D80wms63AeyhSpoykuXxdhMNvuZQQFQGB9ClAl9YQVHdoBKGQiQk0Syigg7Mdc3eFxh581x4zQ3g
Ou0S3mibeUdJL2oat+0wLqn3FN3rzRTmcaV4Bkq9xIl/Yq8jg3e/saq8k32WQPySbnw6hczCxX3c
00bIAlKS3/KXXj+kqi/sb7peJ/Tvzfz8uaRgQZk0O/tdomn3OvGMPYII6DQmCYf39B0tuXj/JXS3
uorKJXH+4qCPAMo2YtGZHHgrKa/YB++Yc0cmyxRKhpiLv2x5ai7xAq/96g8JnOlB6g8kLw5yeziH
ORuasZZB2oD1VxQp1p8tv0FaXyk0Mpp0bTYt3TkycvnaEOJ8Ph6NRRZx2ekBx6bBnNeeEIxduHVw
c1/qZ4vI0GeOxov6O7whWHFOnWOVWFIYxFEp6MgsjBwQhM0UCiBbXHPCyvyNzo5fYcVQRKXRlVxV
J5Fblw2gCY24+o2NrjL7oZzh0IaEkyCfbbGMK8r4wivJ5Bhvk3f0dbdNGf0ekAG9I44S6g+XB2fP
Z0Y2oqgP86ZI8QgmlHNQ8bxQqPRPsjfTp80zYWiabLKkIStshigDyykaUAUaA3utO8Dgab4bohup
SiRoVuADGLbnn3TMeQiE4Ekd05zu2oNO1u0/XXRG9vuhYG5/rnLDBH3ghsMXMxCxOk+HTHqKTTua
IG9wTLKc2+2uXXU4sxDo/iXwkZgUH/YwUwoUb99K4ZS3ofladZdaLBwyy6Jjt+H61XrT7Cx3vpWo
N+0pP7p2REnHiLxIx4bbpqnSG1QefcBn4qOVNUSrWS06Idu6zRkF4k/QQUTtMtbY3/Wr18QRa4uT
hCdFujgG9o8sE3jpt1XfwiHD/psq7BiF91mZ3C+ZGPxk9IyIcgCSDIgMCZF9AtyO7HVjhWxpitfO
Uumj7hJrPCEBSYlvy2NtYNlYM9z6vu7uA31EXoBUnsjab00FKXnhdytewPkJSvltl8Av8BurQsx0
QhnEfyIZrYKoDe8zrfWfWT4I9ZlbTL/JxP4fHBaEbe7Fk7ekFmOs6qb91doQDAXmCWYRFLyMXAyZ
EtKuPbLgQrNcZA3LAjQlkVGyLgRpBnb0cLQ9YKIP2J90T/sXhP8PxQdRtcvRs40XVTLAqotPi2rH
eX8NbVAA+FvxLdiVoupGi6gQ41NgXONoAj70L+YPNIBcIjz9McXQNeCSRFtsK7G2dAV/iaqA3BUv
V4tObbB/WwJR1nSKr9urSgEdbQm6Ut7qCborIWVQCAKtytT8edLCeTKvlmzYSOX8ajKwmKTYqpmW
/G7B0D4FnEAso3wDpXIoS+G8ZoBXGGnhXnjT9/YTlEX/v6KiTtjUk5OqEKLLhl12Xi/baFqqMsfB
L0CIiGqQWTTMf6hwWeqzUwnJUtGoUyfb+YJ5GZMXKDHIF0Zyd+qcdckoB2Z8G9q5M+pNGPq+cDtX
aVMhI6p7fuaZMM0nqITyUYaROlwQWB251YJgvVeEXvD74IGhI+g5Io6oQqbdAk/ZreiD1EH2FYwL
Wsiqb4IcLmQfJCOvvD7q3k55gvu13h9kuLWFSEImDRwAXEp3nIY+lr3qWxyWnmsEU3dLeofkkh5I
zvAtM8f9gYZ7YtOwRPH+Z7g9kSIMc3fae8gb+Pxqh+tX9l9XIwIfaN9guAVII/1rYFnWys7cqaHF
I2tvnfrUmSQAfpm4fSdTndq4xh7o01ZmiihqHWdUCDAHMjNZj3bgiGBxBPExgWQ606FaPfZ/ydSL
BBIFbwNbq5tXoh4Z70GwHIrBoz0YDZA5zAMES8tq2+fJS6NdaL9SAFaOaJc0CaBd78CIkI5phkgd
mPxTnJN9/5o40J/ivxGwF1oII1Bq7O0cZNU+tY6PwPjzPeaqddL+eTUIisUpFOfS0wTaXoedlhUl
Oo9gAHF2B1/dOZq01MTbpTCzJNTR3ZZPeNk9/Ig/zLIhQlEbnbJc1ILzO1ClaeGpruYzacdvvGeD
+XDC99K6CAKodgaefR4AMP6hHwe9HDWT0dKvby0rJMwnoDC0Kgo430JQdN5cclneaxM6RIYIpQnh
SVcM/xmIBmBkF9096avo4Ow3rciLXXvHaHF7qHSvtvks6zjSREzAOJbNh1qjd1JXV74cSilsfE3w
0NRN56eN4yeim7mrYkNPuCFYEgFFuG/B/Z+unFGsstn+qtZaSabOSjmeXWOmQFCOlBmXB4yG3UKn
M2o1dDbmVCzu1SuvTNj0VKAXaABZTqdTipWwGFNOI+WMPHjtzyFAkvCxlFQiFdkCPrBWlNs4Yssv
earL0e8ii9wJN5Wb0G26WGAH2TUQEKfXZVTEhiOYb7cnZ7/8dChPAOZdyyw/wVfQBYBn+dx07GRr
kraD4i4ntKa3bFNwBxvoWUVynwRsvGe41D8+LnEebREwUu7rXI2t0tRzcuj9IXNF3FiLuEkfXFJ5
ZpIbFxziNbAd2k9LnO7Sre6TjbXEMZRvtKfkC6YIp5JVc1X6ITGIUIAbVDygmdipJ0x1T6yxRrdT
NE7m0LxDKfGfWDmwR5cywx5fGLx1C4y6eMtfUqOMWHWx0p34DIThmA+iRj/EOb1/6HvWjfrXH1ci
6zFBtctX0lliX7R4petkDHa9oZ8dtsTFviIyFk/QYdasXm9mE2DgAkXUjAhsljmxhRqpW/yq1Sd2
oJO9Gv/bTIZG15lRuazLPGKUgzvtRUFqbmURoKhOL0puoTKfiWCGczp3wo2h0VdS58Ou/47Ty5JB
yQN7M2T2gCulGtSqjWgqVk2Q6W2vWrhZJV35sb8IxO4OMdJldVshL8PHNXY2Yc/uVoAZkfP3AWxN
FwosWLVnYKqeFVon/m2igzvPatYUGmihzSRCx7uehDN06acjn6qu1kB1ez/35j6W1eu+kF+z/wCt
I1PIq3aHT7FMxdCTC2HlFBT+li3zp+qZAlxVV06oMcnVD8KwrgQEbPAhzAF08j4upVt4Iep/noMl
5cl0/uoBlH4PVVO1sYAfMAog4K3OL4UZ3nQAUa1ZP7YU0ZgCnM0DYwGCockvsz8+PJeYIgMGl5J9
/1ZCP0/fcJe/2f2Xf2MFcOAd0OrpNZZ2Rtu/ts0kl6RJ2rYBcvmV2M76eN9N03do6HHoeRBOlDXA
L0mJ+4V/x0u/4sVUNXrthX7J64UJQfdnCEVTBVDErW5SZULMiTkufrNZuVugjt/oi9pg4Gd/qSlP
fZBaeW+TXp48VkHMaX1aT8RYE0lKXVaNldGsZfF4VgGsrizYhyHnU7wFeyofyWXLVIwPmdYLeUPW
VsDBg/NiJJ0zmtayWQw4Dkk1uSYsra8QmCR6vBuntUs5P7jJ1xU3AODV1/6K3J35MFPSkavUs4Mu
3g4uHtpKIYNncPVEikhJW2TN0BaHufL0y+An8AON1yHwdJdqP+fVtjRKuRbi3KqgCjhILS+YfsTc
04ob4IHh8RH9TNe3mFOumG05r2m83YAWQ8tMtWkS5FbVs+8ckjBqDo9+QGkCr/yg4uQvPliOkb/Z
iLI0BzgMXFbzUyNroUiScNEXdFgvP/e7HRqvr/xlUUag4Wysmjnvaki1rTwDPchyTKlrA0hBJob7
cQjPk8EMnK4J7kK1LZRtbm40Njk/ZBOwRVOZX5ZIxr10UMs4L9F3lGnEpF4WSA/aDg7uRsQ6c4CF
eBQ6FWCnRD6w+pEEa4tYt2ZJKXVW2qHP7Rq8trDMbYR8dIReb27gpzxA72vM1uitqNBnzSz3a7Hp
0Ee0kjQFwoawzyNzYMQlYEj1Uf5rj143KVy66asTN5VIGVSrBxWY/V7dcQ8ctHRxgtTAhJlKh5hS
TROpBKajyuOkSeBfMqm61MFzMP4WCd9X8nqNSuGtFr3lwLnArBLcJuM0F/ReiNv99zyOJpvsJPzq
7oW2j1YsxVWsp0ZKTAc/BDDItCeGTQrYiXYCh+FXkHU/G2ul6Ul9oZx6zMg7bEFvNkw7SSmWZAHg
BBhTu4oQuZD1mb1tGb1vGUATwymqCUTwR72iBoqQPDCnX8cAY9TJlZR8GOpOQ90wtI5mGunQQD7y
FcDFQVzcM4fwIE3UbNfH3vMCuPyJIde6fn/GAc8kdompaa2uTJCoXMIjIgg91RV62XVFexPpxcvy
6/LXtiehvF3mhubmTkb9xF7XyA25r/5nqi9rIBIIqbbAH3WQtVdJMcIknj3Aq1wRmoyCVVlTGRLT
ITU0/jlVp4I4d0f+rtCC+3VXmhDdZZ3DF6byuYsGqy5UPHLD7DW3DV2+kYqfRfLHbBbgJfCxWumR
FS18SzwjbKCaaB3cjqsMCQIupjOoSBIixu5bpV53nlmy6GmfZ3i2VqufgKu4xTZVtP2EJUgPlqvF
D5W6gueL8+c55HfYrgljZrzsG+IZZjbWST9TRLxZ6RcrtN5/U2hqb3fHG/WqXKvTsEF3Xqqz1aCF
zHHqH9C6aEyCJkNNxWA+o0O2CVi4WbVaSVnGfUybzPy4AHGTGSiFHNR1TqMit5UFO0Tn8HCrQLGk
pg92srtybKragx2bIshxkzwLuaV+bX4P0O1rK6VHbECoW2lCVShjgW3lQO7URC1xQtDbBVPPrpM4
+RsFj/zKcMMBDwRK2ftU77OhBIbOtnuZ5N49+xt3te/5uMTVnoRDUVUPalrR5nPcgfpO8HlS8mWR
Apqa9j/wypVPpKYp+xNqlhinnY4UMPkTasU+79b2V4l5oDPdVmyPuCS3jw62xBj5/OaNZi8yxhol
xFmVZEBXcK55qQ+GMsxp+URSj3CecQEKfeSBA91ul5+uk+I8VrBbWR10rmrYppxX4eb4MJ87dKXR
lLK0F5dDziZdx9NaVESXzJJEtguwtaB5i5fXLYBAs7bAHw+qoOEVZyi45hLuL/FLS9BH3iwQlVS4
abx1rSUemjB3rrMOxeEZKFLBN9MhI5iLlygpHIWnhRsEcKg7kFEYS6vd/uKighZUCoQVHr3TPlfS
z2hD9kozwyKo46LRDekj+wgIrIgHh4WzRfOCM9+D+yJHPcxTeODgI7YWprn99p3lM9BinM/2/xqy
aqyB3k3kF3GDsLJHxU8Q4lZxzzuNNLjQOMpvtsuYCVb5kd++jeswxId3bjcrongabR6s4lKl6umk
pIU1cXD8d21J54tNR5wl/bYcSQQgph3hjTzTsAi6PfLLbZicpeiyrkKDvzk4bZK4EICmX6wQYlWZ
qdNxw3sqZryPh0XoNkePBZ5htCk8B+T+js8cDa8X8I1Wz28eJdd3hFEl4baz5i67x2ZT1ihLI/z/
WCmpjGQ/J5x0RPuUISve6cTkR5LJ06FhXhvSEzZ2dQq8Fo0egJlJZaTIwI2Z6UaZfV+g/ivTKr0n
KkYg3azs0NixukAmD/l6Yc21z+iW7cmSm4DfQPWuRHxW74LOjhb6M6BDdhSpL5xstuzHDwkg0Awe
ioPannMc84K9zB9uR29+5lsCm5XviIkI7TaYY8MBivafzXZRyfCgeBgfp2VI9aUMvY6/SiZ7nO4N
WhLkIf0DXztshL3U+iVh60ZtIMroOeArWNnjOD0+PvjcS1/xYPVpYJsDswxp6LmK5KUM3NCJPr+7
pEcE6ZtYVB98LfwDRJ/+5rQAgrRP7KWGGstfv7MTr5Z2neDup0c0lafau0GfcNtf6Hb+aJtRaukD
1HsEF29bxHfxh2Lc1QiOl2nSaNMJPs2gR7uzun/JRD8QFSgVhU+NZODvRXNH1sK0JJmmNbnZh/Eu
73tF8M1uDV+hproGPq/ycTlPXyWD/8yNsxMHDOXfbx2lJlf506hXXrAUocHPte6iBnGVbeT9ElkP
KWzpHxvvY6j+NuqkRV1dtu1V+8Xpsm9lb1QUTMHGNu0eqhA0+WXTp9N2P8+PE+IF8EpMX/a7Kq72
pq5KhjjU+BmGdAASrLM7i3ExM1ngXaF3iCdzmdmYnssObHsbYCgmnbVfu/nOQjBM33BsRZrf1RRR
o4jncphKi/Jq73a0yGGmNBCNAAYY4agSMeQfKbG23MXI2NlUkY1Q2qliV5jtv+I4U1ce2lrkelSH
sqlBoeFQtfK5wY3RJlcHED30CUkVE0DVfr7F1g0JH1+LigDdl9DQ8lqKkL01jofrW3P1jFRr4AiM
X4ATHg0fIL4EMIljSnwwieXMVrw6hjHGDXuY4FRD99tHdbW6ckrcTd2XdoZXd+UVwHjBVd8SpT6C
AJh76sjj32wvQ9gjPDyMaFd+kHuGGYESr7WoaSEs+haGEyrHuKjFq6IQ33H8Pnngr1MnFPndHAA6
GO8UsDn139KWWNEZZs5E/v9p9zsadYxnn1GNeD7l2ATtdN7nrBxn76Fp4umb6Di1yM86Gfem3hfN
2DJ2Lw9AfisMli+fiM/UkbC8gajf6a0wxotdgIO42gJxZi9PQs/PkQIXJRhz5Xc9K2qGj6lTzQ8U
9wxsplQnV5GcAeJpwSBCMkKqRezbx42CyalP1buVygr6uggJpg7bRPMot8zbeg1iqnarhQxVpDRg
H89lebSp+izF/DEvJrSjv2SVZ5Qn6Zpl6lemSXlyMqu343bKmWDbjweQ60OMpj35sBg8qE/rkKGv
gczf97d0vUsxg7CcSULCcdoSXmtYboy2Fm1ViM4KxvgXbW4y5fC3B5e+NI4az1CFDKnLgGYmItuq
Cux85sRAzwTm75LwXjpD60SjVdIY94hSyCiimH6GhATQqGqLY1jigSbPb1fhvvaBq8Bz2d4K3AXJ
9smBN70vTd5ELED7FL2uvm2ZLoo+O7EI3ci5UZ1qS8ulEzX0mWVwQSPX/mbZnzKM9hmbec2HvRoM
xVbOtDo+G+SNQk0mSr27Q8WkeCC6Y/bvxttgM3Yl7qO7LZz5jl3JxWd2dwP75HT/ZwZNxwuB54C6
3DdNYar+vudZWad8DfhTiHcsrghNh83TvDvBLvLd23Ud5jGVCyVPuT6+LNbx6kGBdGZTx/2CtnVZ
N4+0E8gVrUeI7/zsPZ61LddlttJAtc95e20AY/OTDzS+GKwDyL4N4nDchG5/LZFTaQGBvXGVsiLX
MaJmNcBC/6XUytOGhRWqmbU1ZK/a+9sXxDvuUwRDIEkF9RKk9FhO/rBdhERSK8dVl5lyjUejSo1l
nbA/V0CFbSZzpEed3l68T8rukmpyRRPtLxNJMBzjmNx2lOZbYgy6EW75KixYMqovODoflBdweVWD
4Zj6VqEoRwdYbORpNSHRQt2PlicQy3+SvDsalV3Ecp1cVe33tpUWM4JBCrg87DDAXs2fuawNqJOJ
IUo2BJ4LSnIbeDqDu57UQ/na3oZ/CHNo9cAWpbidjkbo//YAsHCz4P/nVrIvYuFWiPEe2Yq4b0ak
FbixeIElk2bqJOW4DKQMwN+WGlB3wsE98eeGBX8X9jCZ0+dH72HclMQ84VW1pBF1dKIyNY/FpwMj
PMgAjwCZBIOXKBU2LLCNnLGUeJNop5gZ/EiKfUxH3fU1CFN46KhYR1maP8c11qMkiWkknn3G+peO
Yo++pVkBGINDYYZOADOpKM1hkgtupZ+q2asNRhy2qcH4/wcJHGni0tkyeztRNU9UwDXmwVw/2C2U
pvuYHekR05xq+FL+YOTfx4YbKGV+OjtRQyVbLZVP3jiDUb8N0PHHwh9phToOSA00NmkT6QeiltTr
icsiG0fdMpzichSjTERaBfKmkOO9IagzChFu97Y1Tr5iIMD8spIq02nPQo/dJeaXQ3Xh6bAZm3ee
As4gYd0kgCeq2yJRJ8sRl0noEPdSR0PyiuqEzk+6lQzHEZluMjiHJlrcCHmh0zTtiI8gjtef76zv
Nlggs+m8DldMwAUMB7UnDFerq7WC4cLHX0fCW735gullAMBsEAwC2uMgpiG+BMRIk1pI0cR51BO7
Bufg/PLcGkNFXLkUtGpo2gXGT6nNWcC/E66LSFGTEuq6cvrTc2kPb0CXyJ3joCXiJpRmLBXquKby
5hTOZPPsHO6EScj0QmQeq7V9kUnvCAMZ+J2WFIn2WjAoVwnK+u17bjJUPqownRHCzMazGga90q7k
buPoFJSZadqBnJzCuvXBhT/FSd+2m+9ZB176OLP2/9TvNBv6rDspJ6v1uKS0eIMMtx6cj0EnoAKi
v+quuGoxpbPtzlYsshRz9Ct7PENAxD+BVkk7ddj6cxzH9R6p8GEn+3gMq6zSWXrszw5maWglhXnE
LJO8LLfSyCVgclket5d5/py11nrk+EgPHUyrHaku0QDka/bP4dI3UWNoKcn1gUwL+KzgqGNkYR9K
cz7EJvV6Adhg8YQ6XeqfRFu/Phf7xlsaTwhWCSeH+XJ7Qd7IeCmx5MfjBcHTZgTNF7oWBDmX3oxc
EqsZ/G0z2Mv1jzvxNJT6fGAqb3hQJMm3TDtwgYaE3/Nr5/ruJPI+TusCWrZqpDhNjOBTMcow8BZv
pMbP98XPrfcqpo8nJtZRndXXrGka/xhPykZALIqZbvjyHjYP+5LbuS1VNpuUE52gF7cLdJzn/yDt
ZC2BEfNriRH1uWmSMxsDwIGamsmE98tSvaQcOk2+7iR9mcxPUJkUlr20JpMYyhpeYotH5ZtjmRw8
2dxbP5j8McSf7RddVHs7K26AQcZHY6m0sDfw8gkm6t5afsUaEodDsUD4w8XYcV6EQE24BUJPae5f
hG0s4FQPg6ZUtJtFiKqNC8cxSJgyGFZHHFaUQJ/xDTXjdTGdfCyEftI2Yv16y+LUq1pEXuVBSsj6
exLiilt+oaAsAy6TzCM++q32ZXicLgOr3ZR7hZWdjlDIZ4I4J9PRhohHMJKPf+fRb5r/nneQv+0i
HblOuE83Q8Jend7zI0tLaN7NGUCGCIxbDnar9MZ5WWEmMaAqjJoMi2sRAz8O9aOQpejgfLe+XKYj
qAL7LLTVjmpp908WFwdxtSQQltdnOIyRrobzXgFRWVeIO2jZhNC1eNra0+WcUTnxgZaUaLNEsKPk
c5YopqiEI6mYQNrjbUetxSfHt6QVit/M/Amwr+hfkA5qFZ4rwIovDQvaOLxYP3eHuUJg/6EDi/Bk
7l7cCkk0V4/k63+q8/OSj4UTRCOtnNV6kCxUNef59U8GdhVZhZnCiGg2yiMD2CWy8kfxZy1W2I5e
G+QtbicLT0Hwy8wu6pI9nKe/gKJa1EAoHpIZcJg6KP78LJ0GNCNsPgaDp0nJj653/Hi4T+fOxHD5
oEGSXG5HqFjN5xYpTpTb4afREuEHOXaWh8yJh2RG8I8TIH7Iw1+k6YrO2J3d/mbBjoOdB7WgBAV1
Qe70uIcAHWEY2HqadFWLWuo+C2M8UxN4FwOTqB5Es0CmiRgp1zcLLjcgM7gbJmiCsZs2XcEZMETy
hKWWCKyMlZka0/xxngh8Jr86shJf5UniIm1N3hujk5XLeaPPwxHITxqoq6D39r0TAGzt9g/P3YcG
Oy6TEKsycNmc+O4OoItWimjZbM8K6KaNaksjjZJ7GybbRtV8sBof5LPPlyigmNfmVpRLwC1w+Zja
78HjODR31xbnOiZ5Ql1WLJOv/YGJrbgjb4EgZt0mRLvjtpNBe3KlacZeCX081yS/Sm18HxGNNoJF
KTXe1KWkEy7BztwvLqoqSgJtmHPlRtNh+shHxjnFDmFH4OnBvio/kaoadmHAwTCSrkqOG1uLMz38
LA5FxbdN3fsymOUGdWygD037J3M+aEJwei5BpudFinQVdQKitgb3i8+dnEEeGZQ5c5NEZlJNB5+/
n0DgkisITizxlU/oKdVIZATpz12J9UlN8rmxAoT4pczVckidSLq75folaVQZOfsiJgRUY04vMkTV
wI3QnAW98KKrYaymwMP9SKEhUCg1r8kDdfa90fCRNobo8c8A/oiR+rjq5JClfbLAdWfw9DmAh6gw
N29Y3lZFi3EH3YaXIVBLW5VN5Bbqs50hW/BX1jJJ5ElG1PSw3fY3KAsMFQGhscS3Fgex27ptcPTm
fH6V7EedpnBktcz/zMiokkSwfTqGnMJUrdQ3emHse6omp7jFiIHMKa5vSCmd0yNkOFzg6t3qRCwg
+69OARZqB6AHKpOlRZApEQ4qDTbb+lRzBa5N3teSEGhOmkExTcNjtZd/vEXmaWLmMmhXTA8wuRhj
kHnqmydpo5+znGlj1UnExXjAqpePDgtfS/JaQXrTj2S6YGyfn2ohZbjN0/kyWCk1f2wP2d2SVMN1
/fMDhz7wcWln8unsD85c05TgGI7V0YNwM/2Z5ai7K1AU+lVV7O3x2BDyeqH8UWp86b8Y4ZefsptE
07/+wsdBhSMXi45COeZnTx1hfBoRJjczcfgnJ8XcsgY2si7jZWNJWjNc211vjQHVRwWE/7xYkn3P
vbT4pq025AOTkuauPjjZN43KfgjBA4pjNjp+oYdDGUADpPE65CY8C9Tfo+4g5jN0h152kDYhxm7r
MFnmqXpA4s3yt8YX692xidtjKILBHNwu8K3ZCa+XQhVOLGBclaP6VEcz9k7VYTbsDndNX8yXNUuy
/4PFGmFxu5Kn/FTANXtnhAQ8UdgXlf8VSCBRtdVVpgJW4KasEwCQYTdybglBlTf4P9npm9oIC6o7
2v6uR3+09ZNWUeTp1YU+Q+xEvqHZALloYvwNJesUAg/Mb1xbpNB2tYHxDeekv1R3grMeI0CAqJ3J
vO9YlJtaTvVjkWLTc1mtbTXIC8ZCu23UUG1VwOBms4ZTUYxcFR02C5zjppb4rauLgTzv8/kqX18/
21yFJtQIwyettkml0a+SvLSrgOtf0y+mX+210DyQ6v1rRFlzVXuWki90GZLOgH1d500yAbeIzFOg
Nrllk9RM4SP9QB+i6DeCAbWlHnp5zqAeZsl6uVRBQUWR/CO03xUo/RtEAaigWcHRD3jVBp/ZutAf
HmISDg6EUqjxQCZWhICk+ds2M74gRlckcEvDNoil6t8Kjq/MBlFyDbfZOpw/nrMPQr3NnYoYdXyw
N1rfD3vh4+CPaOLk7SL2YT9xspCP+KL78T++r1a8+OehtW4NOAEy829+etee+TqMcxePyrCqKgJg
xp0VqPUOt4g79ecpmvF7LLPa7U1rtyMorXf9MbUfdNspBxyRHYZ2+L4KkV0VCvjjYaFcXaxG4koV
DC1y/VNX/3EbSmpFKFBYtzDqZo15OlUaZjAzNLMb0bwyc4Frrwxz2wTmEHzzT1WAvA2UAlMMB4s/
IHb5l0Rdvc3QpR6SPBRjJLFkcakNzLioWmL3kPxp4Yj5e8hv+VdNkctTtxiQmZIKB0eE7ZZId13O
cb3+39vhWTfaqmUGMC5Bxfxc0iyRul+jAOwunWSh444VwzMbuBvaIPNgTPzYffhWV4yiKjTwSiOW
q89+MXKWvH6tAN8g2mE2kHXzlyCXm5jiddTzJVP833Z9mvULBpJtidxQ5afOrJxBOFFGWgLK6Q0b
+j5qo9LY9zbJ9TDRKf2kdpgW12G0KTGANZac/JTk914zawYl1BTSL6LefPnrPW8PbiSi0p/DVfs4
sdvWULcYyyLKlCaLsHNyVb9FQDt39YaaT+diTACs+qg2CZut0uRxtuCMT4zn+CkPrayqWSPQ0GVz
H/sYgj4goANF94Mttzm/vkLG/ckwhTLqJDRasHqZiZNv0mrRhOyGb3idjXbW+wHeEVWrz8Rbe9Ov
7IBWgFA6dsENYQMX/lDV79QP/GXFoBH9NlnG3XvOd/Ymz2uFCc+s3tksjiePltmbLqSgtWlz6lwG
WwlrPEZ8HDSYqjm0ZK7W9pc9O67jd7GzHV5EJ09qeOEXyJCJWuwhcVX8mJfRkLxeT0IZkQqFb52v
NVk6r1CVFesq6z4BVPXPLCySBPdU1mZeyZ1K2c6KkE1vSn4J7ryVFxiYNHeHjF9PeLO6Y3+3LMR2
4NRqUF0KlYTMh/3+OvSW+5ty3PdTRqH47QyNMeda7e4RvJgncgw2T+uQf0MaKa0o43BcYfEaWnMT
5EF4oaG+dyNZBRMSmoTxgMRjJLR4z9aP1i2MduDc/O/GlSDjsTR53IXfsPzv3l1zsgy+v2VfW17R
cEvuH1VvVXGmCvCwHyNPJu+8HpCgGy81B9m1vEujeq5dYGZhOqLKI7Lj4aUQrp/OpOyikNQKtM9y
qEnSnkDDGICV21etRZ83C6QJ1rT84VFZyTxspE5A6UA5hI0XnmFd3Pdh7YF1OSsd/TVFl3TuN4te
TPRmPaUEPMVGjkQlqaQo07/ZS9xSIgwTXKVPvaKwvn3sGD/SE4H4J77M34zwwxlXfbZs9aeZGGks
paCIdwfIkk26y7ESKOIUYJD3npdoGxVS9E+HQ+fEZw31DrKPPF+VGAFbZraX9W+Grrdd3CJyN+RQ
mnjiY9VUQX8qOjoQvpYmBxQMRxl2JrBGXgmrPoWvDUCxH4n1RTOSPJZexsumIdsVgOIjV9UNjTJE
PVFwtOoIgr+3dMDwSPSk8TD31HbIsTWn6IyFgXcrAyv9fRqr64VsYb7Vjq9WSh/mN+sSb1TbiTo8
/N7RUZsCPJnsGHx0uOrCsZdwthO5mfGNfkK0riVnzIsuaRRBgF4pD9xbvd/C1utq/7AoK6IjEDew
oYhC3dOgSe4wbF8bS7iFU6zxo/6sqJ+z4Dcp87IceCvumvalxIIHeqmbAF5SXXY5nBjOPHFU0drE
I7ygoJGSp3iseT3G59NIOJRzXXGbYscYi+AOSY4j/uqp0D4oHQHgIZBvTk3qFldKGOqxF3r083rg
QqXcwAzpQ/Wv6dvdeOJBKVcabtVYzWSHAXDU9jqdDfINJVBadg4CUQmX5kHEKQsP+BTwLn303tM/
th78spDU7gLDaP7JLz5a1tlfMFEyy2dgY4Y8Wp0BzsJ6c7a4cpL0IU/sQJYUebK245NngABBfS3w
ff2LOTih4ppjGmrYi5Q8OHyki6pf/negANMvgH/odGn4Qqc2hy6d6Kf9v7X6wVHCs5pyCi1adiEY
8rlWlSDIQJxWjLgGyx5ozduWKkXI/krtXT28nSXYUMtVDaUHYgQCi5MUDYz3hI+JtZjps+K4hvmG
+UJwBfb9ItwAzX/rIY2Bv8xJxPDtFynu89rphsE2aDq26eDJk7P/Izdu4M+4wNJA+yEssm9YcRAI
AJZDgkKyyjNg9mtem2tCCxyErG8/YQTsL1WRwgZtGsMpX1uKgWJEeOVQNbjbi4i6Iiko7BN5T9U8
jYw194nCXJ4sPhXyAoso9Ya0L9Tmq4jCTK02/ME8rW9lfioTkgLrdD87G5ATKd2Gb3CLynYbUR9v
0kD3aFdH5Gn0/z/gOv1/9tb42TsgaIOdv3t6mHXPUw+HVk1Zwo/FOMtlXWqSetZZde8bpVnFlSLL
Ot08Ujjv2wiVV2QUacRNw1HZJ2TJaIQRpTAeRessepprPuoSvBJfHrGl9kMNgY9SpIbXQhqfSWnT
Lo6PwORKFO5Xwpy5L37w3RiN1yamliZILnDjkrqz85YoJwzZN/wWkBcE6QmRyfPvAPUNVfGD8G2g
NPnO85gx9FKHrO+JqRNoFbkDj5Yg9HJpJu3ne0QNl1cNXBjWMcA4imuYzEPa21X52E+1sKqVCBqI
vM3UhO2ko1OU26UoS9FG8YzdMNC55T4lP6TNgYVcVN7YB/3Gq20mLiNJoRmLxgOUeZDMrah+LECK
vXOykC6VRL+djsWKGHQCZqCEurmA2FVRnDE4QAlc3L76sFnzfrJUTDEeqRdYXFluCtdBBHNxSgZb
9TAqB18E10TQ6D8Vrq/+SkHN5duEsqhEeflCE8pn5a6ytDKYlUdhq8Q86BOyFN49LDWSERig25Ki
Bj2i9Yo4xrkOuIPorYBWpq48EUd2YlUfdHOlTK1m8bUmTpDgbMFvIEZ/hYw7aTXtesW338GF83HZ
yxItTtUVVPoabojSe55rF5dZwHV8eWS4gXcuoIPLYZDRhfVR1qqhVHw+dQpZApxm+P3cGRlC6Tvs
Z9V3JQeAOMwWC/LmZA7QKTvmjC7hSfeOl2gktStk7bmy2Mqq55c7Wp01XLqs4rc+x2KUyggwZA7g
KHMwzixutHzO0BYF7p5nZ6lxYikPJJhtWpFfmdGqSHYb56ptZVpmPrimsG9CMQhYxfKtDmzcTW9V
G6j67SBe2EgzbvEM31phjqGIZdFO9d9Z6HvDJ3hLQVvQM5WYQOYUPlxf1ONhcFKJsngmbsGmNbSr
1+bkbYTDhnQRrT9nUSEh6iTsXko7ge3HZZdXIQzXSEgHsVlf9uwNvWdDHcT6dHJialW1ZIUzC/6I
njoQhRRkTYaEKatN7hYHa3+sBtrDyfEkDMdmXY3zC2wptR8G+0hF+g29R685Gz1sSfQgjkLTqzhL
7/ooJC2fTzWKt5AK6IigHoimNctBt2xqcEShAxdXBTPiILvcXyGis38op+W2uLcdYEDo4uTRLkEd
Qy6J/3110qlewgxBlMtF5iUNvB+QIjbf+ikgKzMfn8tXmmziN8wfh+yAD+KC854y95AIZBmDJGWm
QJL9zv9wr6mLy4Dcg26y//jyhT4tStX+dxCWoVXdizlXOeSQly26g3zXG/5kITPAuUdZNnydlzry
/OMzyJ4BDc/akTp+nMB+q5UNnH8q6pISznx7G8iKqYq2atr9WYhXZ6OEXaadNY8h9nuM2tHGpdB1
HqYg8WpInFcaWy43fQ9AXHi6ZUK5IryJgC3fIv7QlAmMyD+yTbddeaUEnSDsZorJw9CtZPZ2v4R0
4myEo5XU5RCQ8ZKQ2fBuYQ+JZGahv/mdNZzhwWw9XtRAD113UP6ajYVaWgrAmHEKVUluRnuE9pLG
37ncUZfnjAEPp59QUGDXkW1KeQ1ryr8/6wQoZ5HLs8bC70dyxYGEC/y27dLkJt51g6jv+g3uuaVZ
8lSw4FJGs+XgCRrsZYLZkr0l6n6bWP0rpYXuBqfGtUWGI9JsrJBBLioqWQTq1WSBs0zLwVxbnuTx
xUvkR6fnFM6U0vUC5TnHWY738KKhQHLMKqbrSYJ7j4WDRpUrLVCm9ykIg1aWlDCEirOZbFv1KdVr
rRYe917cjdlLQIfqXy1Eqm3d8yVRQTXl4Bqshw1sj/A5mMYu6DGy7F4Vj+l93Doz2LEEwFtotnPR
5Ke0FxnFOX20m3XvuqRLMglPb2B9QPtqle60wcFuHu4HG+ADS3J7doTvo6L3ehmGOdUM4jWg8rVP
WNLbBsK9SS5wFhvj8V/QHI/oSBoQRplF7HEYH6COEn6WFlnZcWGiRcomaA2gzhc5kdcqDhtm6uqu
a4AiXnpnqKrcYXI4gcQLoy+KzKIR/wMrr2KJx59eSpzumoTaHWGIQNYCkWjttUu9Y+EYklZNEujU
0X2SAAux1R0ZsLzxKXoPYO+g8+p28XgFq0wYE0f8b8D+0IDI8pKCEK83doPcdzENYLrkgPvjFrFR
LteNtBwRWqFELtvuOYbheBbT4qmqk8HDSEKJaJwesooNwCRVLZlnwKPYosJHFoFtCVMCtbmIPV9o
wQFftmoGw983S0u96PP9xD+op6GX7uKhv9kcT6Aq0wReaKBeLL2UokwmEq2P+7RKYapu5hVBE/wP
9Mn/wyq0mRvdtqZvLSCTP0RRP3L37QNfKUkt5RqXrN1iFPooG5kW1aD5d013b0vS1TAgJGSB3vet
zl/BvsMDdS3HrN/A59sKm3BZ3l1w4wD9i3gXuukGdv+h5dZyVnw6pJCaBwcG+YTzs8MxASV9hqFW
YrGeUHVB1EKXfQ+bPIZ2Ovy7dd0o5K+zyG60wvELzr/Dtf6biQHYC0NhraGiejsPGR0aOfI6sqm7
nLoIVU3OPWQemiZovTZyvtYg/EUMk8KRhbRGHwki106XJw7lfeuQUl5TFcNFuKbT5/zjnDV2gN7D
8C7KYc7UrS8FLx7YnPlsaZuJGvbKyfP9YbjAqv+sCEfQhaPyqAN4fmNa1qQ5GQbkT6kCTAXsZBSs
gAb83/kHkDiUVWv8WPseF4JYMM4HoSGSm/e5WOY3lLJ42Hv87CTBkX9a0AoMaVKzPKd5ioR19rjC
iqsmJZC4f2WDCBq8uMHs2aq94N4zcqRCgYi3qCIJgHjPMkCZOWexehPd4rKmooMeTV3eaq/qI1qY
XopcttMC0xK9lK5MgOnPNkBDhXsMZrSsqRGzwvdBObhrheRCcxfEWI4Eru1WtgUqcPNeKSOJhT+8
WyBijsgeqx0oZmqh4OG/NXIEZfViuU3BWLTpYZPgyK5uG0jRDGe1Z+xQ+fdE6XWi/aFoz27EGdLX
/JMsEh5/AK7acyx7bXm4CS2aAaoNvmYo9eIBI14K72EQuin+MaCQuMGrhTb/4tBoObQ0je4VHTXl
RihVAvOSm7Vf/1R7dFBqORh1dvq/oYvyDYauGHGjYeyG0VMuJfYB6puNPHrdHJeQi981VdbqO44b
MVXIjDjSWBvHHqnph3Zq9gey9PhCMkFV4XFFMoQNcMjZebp5gm+4XVwsGiSg7+Vw+0jk6g8YcDbh
/XkD+uuNgifI5Cak8uox4fiFMzbpDTxIpBO1eVhNM5lbcgswSfEOh9UUz7Fm26gXpWEFXBSEC1Or
nUFSvGRjy2aCXhDE7qGNC2w+M9UUJnehXcTgchNErAqWYhNWktv9QC6Zz8DJ5sGQTEw47Fc4r8AL
XlxZJAt0qLSqlBGFGxRTSLhIuVqsCOSQqs1evlMBEhK2IFimCsUowJSwJaR5jQorFoLkEQzH/UPK
2UUkTrSluuws8+S9F4mH4andvSxAMtHsE3uj1hOQxcbqk2JB1bSXELWbkdCbNs8UmIOEO7pRYQj6
gFwK2ZGQ/ng+A6mcgbcmY0bWNANHyUrWSzn1106+0TEoiWzyAfVOdVqf2NIANQ5045Lr6Jvy2sCc
KwwnlJHjG5XmaetyV8CrP8Pwow5W5iKWOX39/w4SsXKc5d6CoFQnInA2EmPTiY35hUYwPVTqy6M9
H02aLJdjO+yl//VLqR8MIx8wkcZlEUeeamW9F3Bn4swKtXz25NYS/uEf4IVSC49kPrPh7WMGBhr0
nXdf3IwAKvksvfJOjaf/udt+AjlV2UDNGTQou4KpSiEimR+qWvVoR5zlW6JDmrmMdKf0cnbvZZuj
+qOYmPmpXeGPn10609UiR05r2vCRVZv3ra7fWRXAor1boqsOncgGPiZ883/e0pZRTgKPS2vS8UtH
d8QzB2f9z40tngJFZMhn8xafqE1mwmjk5bRgIsbd09IQ7qBFSmsuebFZ3ZVciqi3vzHGpUPlSl2h
a5BKEWAcLrDCtIiDC7N2g5qp1i3f7xkuQPTUCQhHR432aDLb7lASYybqdOCEf147P5bVrn30l50/
uDLhqhgX8OLxVXq+8djIOsMPgdxYZG0hxSOUCSB3IKtp5ysolEKVylDd+7kZdJPDB1ZP84sWyQA/
ADpM4EbgwiBItCFLFYx+4ck6lXSEwpXPMQjqWAG9Q/TxwsIzmd5IhUbE4MOg3KPoCT7mPjik1otx
dEI5DTj8TEEasWcWK6xj/lamBZWkqWGYiGk9aoRX848qlXro5B6VqTfNtv4VQrnqA8/4mv8cmleT
MK7Ee10bG1fBhmRq6NZ82Ty/mCzWzvpzU3hBxzDcJwOfCXa4RYiTvO0DU7+4wX6seL7N8fgLs82K
GbYnoaH/2/u8t5T/vBMlAI4S9R3gWKGHBQShlN9UlScx2cX+OXPv1oRJLrYPGYIc9EfU299yeJXW
k6k7m3LyhPcH0QdRt/iKclZYauInjVUNucp04HXS89IHCJFwQ+BsNdQPy7V5Lpd671vpKmGtwtwk
lrNAgRCtrpx1vEr7DhwXHkzgc9b09qg0t7kZ2ieRTCVpIWbMyKjCeJLDmysysg2ARgyzRMiVddIN
CPJ2TOHmOH3kxW1WpdpsgtCjuHK3drX3dNXZKLw3Psk4HZvyvHdWx4JeoH7v5I9IgIep+kAUDRFB
HvWkIiY5CDx1EV1hTFgGWf/Sl/O8kB5rJ6e1j9ZhFbpBlDEdK/Utz8LuwIGA1KzkSSbqTq2i8lC5
uPl/7IV/fd3G51zmVDjvJ0wm5sqDNzfuJOBi8/BGG6PjkW1Z3cGEvVMwnhzMRuPe/Yz+xoLsTmlg
g3F3Ebn6Kb/+7LvkfIUGVse+Cw4SDjOHN4FSc9rm9DFILYQesaJX4Te4cR57hnIFMd9eTWARVr+1
Zb02YaJi9UVYN/qBoke9iRZy8TnxXMwpPJhVaiSSoVDQP94nGy3dX4pMU0T6zANMOLoiY2jGjW3K
t0Dhr8TfWKbvjcUqXCEeM4fWiye2Wy9BpdInzXs0szdBMggGoWu6BlxkYg34YF48ytYXGGWP/Qh0
pXECHNqaVbQKfFZ3WMOMEo6EsrpUE+4NmP0zsKy42FCTwoQRTj3v7PxyAAGZ6VIlPY2SxHzuTqTk
KGGpWQsEjEpyyXlK7dO/RaaMs0XrSez5x5cakETaoSsTdiL1pjs+EidmQljS0YyO1OyvuXGkU6RQ
zQGZv4okr2vIPuXK3H0NqemyPFnJ47NLXYZ2FNkmvvvpQD0zDWs9Bp3FbuUzC28iaOkBTIKOkvWB
Kcc5P1Xi+39LQoLc45KiDkK5M+kOJC1JY/O9P73+hGJaO6BP4yDjZkTieQ3N9QKgWoksO9MNjly1
wAYLAyjlkmBR9okNF0SurFrzk5m3Nos7Wj2jjaqOJnANHGPKn+YvV+Tz+RGhPUZpifDobXluQx0X
kT7CahUqJZJ069AFUEFTcOT6pesFjCKZc1O0IHThhh8VuTOgsVOQGhXNuMAxIQOnOMYtu31YSHzb
HuVx5afSxS0Xc0Nspk08kTl5XtdLFBaBduKZ3JO1qpP/dpJzsrIRMDqZTvxBDlnDHPweaG0jl6GI
fYrj+9NyvLEg9IGbMUV5VZsW5sQQK+CWt6dB7rsEkbUCfJf7rTHCPU8YIQ8AQW3+SBWeyr7MOrvk
uUxdlVtmqSf11+tsbEks8vJQpkKPGocM8xKyb3yhMIgNHwLu9tPORXtbbWBgBExUunrAjTs47yS9
ZuIRE27yGDMKSkH4OAkGvfi7xAFvIgVKPkpiwj5HjXsrGMCM3lDQ3id17q/VZhKr9LMwJE5nV8eH
21csYgNLUepPlMtXX0+58SEKXjMx57XRiFu+tsoBBSQ9IZNOisVx+0LOE1jf7XWsFaJ0F2A5MoiH
S6O5q2EMdvvXaus5uL7I0z2kcb58lq8TG9JVBpcIgg6/RlKpPwr1Z8SyB0lBIQYjMaC5CUUA7JDS
OUc7KLZmfYg81rQaXn8uQMjNmghKRJ628Cy268ZOcwn8RRK2w5h8SRrIf3L+v+OMEIOVx7frl6Zp
vMe+ugGchpKnU5mxsgQdOu8kgfwlYSOtg9SDR+pe+G+7Iz9acWMlROvti7wYzNKoqgCnU7ffxnUl
J+ZxkCJ4hJ55LgVggRZR0WOoYR33i0fcB9dCJ68hiZXi4nHQLYGy78Ue/xhA/boAoH2WgRL4SVMg
wYEKQgQzSOZkeGBrfF90eU2GMUDEg9fFkgM5cH43yqLIEfYxxqjTfw/dp7Ip5O/q9Ps3IGMyJ8QR
cv63QWN4Q79aDzf1ckaLmYp/g25YLRK68oQ94VphGf8liF6o7Y/K/JxF1K10PvgWGgLVDL28Wr6Z
VtaXrJOhd6F8emiPp0M5jQUpbwutHaSL00GgfAZc5U70LcncEUKU7hKu7gWyWUrqUiKWiRnRa0HE
GIgQqKWgSZY8m+fs50hKWCV0GpyfvfyQ/nwRPIZx2d/aL8Br4yDxq/+Bp02DwMtid7AtGC6/oZ17
3DQR6xP80JuUIvXynIX0OcRqNhQi3O6usoMrnGi9B/0hwgvkLbJnArhwP4v2SkW6n6hu7g+2/MJq
4AQ/tOSkOQMUz0CMKwdjnGTTwc500COIUFeZYNDS2qZE+sAiN+z2jnJNffXcfz5nkDZkYfJmzXNG
qal4uwyFvy6Qekb4cMSi06+Nltt3O5TxbT/c9ajbeShgCLOnnEvHCoKgO2+nVktETQSVPby4E0Ef
QKvYy1IFJMBRb4et5+S3ZW4N8p7Lt9skA3KUX0nbdLg2GlzBb4A0bc1ZkNh3T1tHc+y6Dyxohro2
kORtzdLSNtZQza6ojSx1P6Y3TMdz7z4HGJOoLRxcmzP0J8fMqD4J//UKZzBW7zISdjZ2qNdc3qNl
Gxe0Mnf3uAeM1sZ0Sv7jEFzUDkqK6OhqnAb6EG2Tcd8ldH5Ge6OhvtYDsO4jaHcoofGgtXPZ0b3a
3HcD4lenKwmEBOCyl8xwqu3j2Di+YwGM8UkDa/Wa5Ge9WkfDbCtH2PXeq2aE1w9Is8TeGbpYgtJi
ZswnbevzqzFd8zgCJzSRKczpvU1L6hbnQaVPY9zT0GAdnR79EW6cNX+Tzlt3GZ45q1C9Tkhtlunu
xGLxWfTTb3q7eDKg8xvt4W2n9ARleyv8X1qLZqDeeq0y4ODnO8hpSIojLAqdChsjE6H57PZU1uNp
EF2yjN2Ok4kusDJfWCG5zya7MRFf+6JsGtvB2vWkBQSQr9VKa/O4nstmVZ1M2d0DuF/HqPeNez6p
WX9N0DUZ17RBYbTQzBTF3xad3pjQJ28AGoMKMA/9Q7DkqREkb5ZkJBj6KA7uUHm7vWhEF6o9O9nr
KY8usAE/w95AuRGQy3do81mFOEQCf3hEY7Lj3hf3+cfEKnfR4VCC6fNtM2W/tBdCIVOkldNdqIin
8OaolVy0zmeM+WGsFVEypRMXl1jcBD7SnZxyZw1Qm5EYBOGq+TUPQXHTTkOMHsmdHRElN6MVgP7h
QTYaiwJprW4VfMFWgORLi+PBkcHTYWT9wMe8HJRetvYFroJOysEDIq8igvKLLEc2AC0DktjSyDpW
IKX5zqE6cW9zOdGraSmrVHa31Nqgcx8zbE8vFSX//TKg7E4qQAPODpc/d9ZvrVcnM082ILPcr0+m
YiCu5MwExxZ7Ekq/9lTIxLKEDYHtMLw7LW3BqaC/EUBBICvwQUPNrKXIeiw4fqdMlSpm2AclVger
W2iQAxG/PVoP+C5Av+MFSUk6X8FiC9WgdP/X/VlsVkp8dmY+NpjkZqJLproSKunxrMSknZ10Fblb
5ZvsBwWcwC2hGLVo1EUmr7RVfKGUJD5/ZzccsjikPO/8l2tJ0X+gPUUfvvXL2eBJl6Sr8e7MNKL5
TSTGDlbDIxtvpvcMxw0fi7N5B0o6QTrgnbsH6VC26Cy04z3Gam5cayA0yTW6G8TV8llXOlTe41Cz
KUROGBmAAyBrsNEsfajYSWJc2tYjlr/LF13550okSHdwUqCOBcn8l31kiPYlGG3ckjyYU/OQ2GTw
Iw5JftFGXbbMldkPqLEVnTsopC2m8w3mTqn7v3k5OxOCecAjfYU7fUUIH/CPEVXj6Qpben2rq/YY
jKM3LkDru8l+han10MXMdGyg+e2CCjBYXNBGjNbu28GNzbtzbXKIzsqEgvULrmrXwyreQA/hYnwG
yES6CsFvuocvfY1rX6XNpUFqxLMyv7gGl7pdogAm/qf3+Z/IVz/tKsWGUpAPfexIHSCHXiMORMuU
FqXW/qkJVYwAGulrd7c4hVHdcxAtxH+IVlCE+xVUWywAXUFg6f5lcBxZys6sPZ7HGhP1LtyMK2HR
c6Tz5omXalKWTdiyl5DWF3NLFmrTFo5iZkAoJp4b4nkcrHduw7yX3vDyU+UvR9vGSr9JWFVWFAJK
5piMUwmIkhyQo/NW3Ni5KBhun6L0/HeuDbhMb2hU7V6iczaVnvj65sj+gWGjjCNke84TmTHbk/2i
rjZbsGmYDSUiVxDNEjNCKPIvAXI1k07ErRFLTIH7buYDSy4r4LGRpgXH4NQoLnCKY95bRqmaWfMV
Xz/G2y4lx7NMzCdrJ8maPYpUJPaJN6EnpVAjb32kj0pgt9aY4hF2jN0Dss/uSfXlg/jUpOORttYA
cTvq7Cltlrv6mIs1Y0QChkDKJwl8x5OzNNoZ7mlAQeppRkLzFgraQg2ghnQzzG3DeOAxw/QDmkn8
RS5UDAdxosR/vofb6a6X808hJLfyZkQuwridQvBNZ9P9Wjh3vklkH8eFjN7uorvCy2lVvTAGlYHb
HU+6aqM/HxMAd11y4gpJ8DwD3wk8bbDd5I/afHS+ZX73uevknRYFSQfHJAkb45reLgzqet34OsDy
WZw1N7AXAy52S5/UaHRwzp3XqaKi/57laV4eyqyshuonYjLgXwT9sHcy/u08EJVPigvX5Svzry2f
roMtUnn3OF7O/DPr5Wufp+Ofuzq3tdtehyn0O0KowAh7gAddSEWZHS/rTMic4MPZRztF4baC21nw
B1E9kpxwoao2VX2h2DxgkUqICrtjcs9Hy8Tk1dNtZWWABfR8OKGjHDxpc7jzUNWozCOhIcrmTPVh
RqXODTorGVWLkQspjk7dP0eXRylOz8VLVl3mmet7mHarIJVGgoyHq7kOBafPGUrzVcGg4LGHK8Ou
BZt9hWLC4Wel8gaLotprVzRN9i06IkPpQr5+mu0TspGTP8sTQbbqjSVbRzl9WYBTG0J5Lq/chx15
G4a3/G61rfbwO2vR8zP7mM854iTM+TPkAW16RiQTsSuXCm1NF7DpNkBpoYsjdglgZlvji7fv+rGs
XZDnMra/fLvpBtH8+40rkusvitqar2KJI2vjxRsCL2iGGhkzs+kSHYRnpzLwhkK3+vm9inO0UvzU
hXjAAT8/Af7L5tjsxKaHan2F+WT1b5ndaEJDEPTFGEJuRo78JJT8EIrQNyacdHRUE7n2a22XRb+i
T07+FmN9IMRcLbtHsi4gYPm9jQ7+BpAAUpfMyCfhdcONl9NC4t7fRN+S9d2hCY2tdsobnGmhlou5
Fa/RN0ylpooO9PFHXw/iJfP7fJIZgOeih5p8dwLAW84ORY+63+7dSI3zLBiy+7oNjcUvFJ53L7OZ
wR+jC2AG7H732H5thB8CSih+qWA63R1k0/FRXF88LJKifxvOgrNJzkd01b3kGv2Gkk0W9iTF1qpG
bh8gL/VEiHDNY+CXpdgLTIBquriI7bKGzGh4N8WMR0vA4Jodhnllys1t+ejkfrD5kcdbRnhmi6XI
CtvlYJlRity00Mb38tx+dQ4c/H+M7O6lOl5J9oKnbrGuGwWRKPfCPflZpJbHMnWB0+Fp/szPU5xM
QdA+3YtwnjH7xPd+8gxvPPPAWZsjVuqpMWhir7j7DZ2SzjKE/LtM0AKFSnOO8j8xVhsz3YK5AO3Y
Rsdi+Zk6BEK+N0eR9N81bGTlRYKPYTAFcGmrzkSdqCqVfnhpqSDA/ZBD/trzyQlxDbshjsoDSLk9
EukaSQItqrGTmMdKvPfVc+jEOONjeoEW0l5UP+LNJScHXOGPaH7GkRymJX6bgNABbJ6z3Y/a308s
1XuXdU8CpCvmwN2ukTwhxH14NUQDeipZBW0qJ2X9LoEErHM8kKYAwB/yUiqFGzq5hdpSeB+Cq2cp
Xw7sgj5xsrFbkILaxO8iju/xYf+4biXZqctQhYLuKSP+4q5hJcHX1rGXiRsWp/uOFYtZX7ef4YXD
98z5lf4gBrK2FCXHEINB1dEL0keU0VwqtY2r3/IWwIeYbuvh0YXrI1AX5maYlXnNnsKS5XwJ2eMC
qjN8npG0WGqUQkUhreOikJuxkWpwg+lzzuC77dRR3RoD28ugPgss2Z/DsANpjcWbynk3k5kPjUF5
vAxHE7WoMCZDrJyuiwiacXkHbOLuUq5093ZTy1M6XWdBZC7e2tU8i14gHdr957UYhZG5L/o1cB0m
52qaX82FEcn4ppjC8YbFgAqn3oeOSfixo2/sYCRfz/9/pYu/c/WeLktVJ4tqOgNS2P/R+DHSh01y
NLM+1FXcQqRMDyr8Hps42Agk6Agk2m5KsjP3mcj34iUHALpSPRcbzeG7cyK5yuk7tYQf2a/LfJ/+
clzMaSPSHAxhXDjoEHfzBpxvh4oQ24/TybS6ieysWCCB7A2Hi0aCiI/uYyJ1tR+1tbWwfskDAfFN
PCbnpBfumfRGamnOSaWT3LuKn6mUnlzyrX73iSLAohQLIrGnGyCy3AfXoGazUcL5+CoRA5OTJVgJ
QC+IsSrfplEIpBEzI0RwQkgyjHjh02tfZNgT17wWuWeAgzKzwVhQKuIzwTjibbqpGe8sz5aHJyzA
FY6mq5c0Yw69xHM3vvnI2BIpxlH9G/UrVoAmjdsjSfkL73bT3ZcyS5j++ZAoj3PZ1S3wX2O7IB1+
4WZYH2bfWlDoJl0P2FLnVjy2ucdFOSI1U9xx92oiMZK/46cxO1FAMrEqFgdvT6swH4s9fGnV9U9Y
/CQLBrtAKXYD1pMoNo1V5Fiwbw9Hl4igvVcQcN4ujx16PYAWXsqSmLurf8E0VgfJ/foZq+KHllzH
eP/9ojJ/NTO3qdQVViGndgLjWRISkIlZ02yMLXYqtxSjEijeaekCCPoMnJ2167dxMyZb37VLZmek
PwR8f92sOgMflWRJ/r3boMCj0QL8iJpRRhLkTWNB6lRQTe7abzZ/w1+u1ky+F+ytuvCgQ4TIUUta
3ouZ+UMxMVGhaShxtiTVIjXy2LJLmNksHa1XSMZv+MjigsqOj9K4f6xJ1v/ddwFvj0sl/eiP9/6E
peqTOKoLFDA+RTseOetmzUuK0W7+Gna7v6KSLjeWd5vu63VSfqrSGvuJZ+SaeLC5rjhELGGbM62F
AaYm99gEppqcWAeBor8kkQlYEQWVGFjwjpt+Cn2Pti37ZGX7hhZXIgED+vXR0mD+mCQYGLBb1Z6X
8Xn/LvXLppURJhpeboioRVmw3Y/EJHhsS2tMmEIwJ5ut0FZ6HamuyNqRVlVaNkwUNfVX2gDuQWFU
nFGwNPK74L8KWtvI6QKGyqUS5IeBnnAB+87KowaLNtaLCeqW53bxQw79+U0Y15QnZPCu9LCoeAIr
prS/dLDt4quKAVhC41JUe3Xs1pP905bnhtLYl658voDaZc4HzhZW29Ukrqhty4a0VsgvAcGwAuCU
kESGAjW/17GnakwlCXX4j4mdZjJWgJNNAEaRXhbBUPXdzKYUWxsNvYMFj6jks9GQG7AHipXGnmZV
fYnTFT0Gnc674d/jRXjpZj11KJtsdpZ0V+Yqov1xsdmtpGPQHMrYEksqmYx/eUCQvboh5Qvw3j8q
TXhck3UScDLJIx0b2/11haCVNFKwNluCptmAuv2enx+Zcnl91R+O59k3yQE5MpbRjHTkfMgxdB83
L3ilHKpredBpdQJ7a4M/rb7tBcNKtMoUbKeByAR/W4I62UoT2OPt1yHu0K907H1G3QdxKRDtFP0u
LNHNYiGLpgnX6gwntrK9K6SZe0pLV1Qv23Ly3HwFX++SVfT9fLoe+vKbZGWcSk36RZGF3sWH3G4a
zgoF7z7fuqYa0Ws+z4LL1EaKFYuloUgxS2C0lzDmHCjXY21nZqXHXKRlOOZER6D4eHAzbbaXN+hU
2HayBfgh/s4q47LSAfeUNPHeIrncxYpMl+oEuj2TbLwGEwDmOMTzRW1h4w51KpN53RW8kBSRrk8l
980nDOry0Zoi2EL2Q6zqUQ7ShLSkJuTDEBADgaftwA7VC916lrlSiPwfZYB9nBEI0A17mZI9vSq7
P5bNCMuIdBQz3Lv+wl5vf20r1aTUgIrDFZT1TF4u5OOQ2LuvgqExpsl+6kmnIS4nw23IxO0uBvvW
FbLCW5cyF56aW1mtx5UkY70jVoKMO5SOnWXPEW2rGfAWwDVDRnvE+IBbqoIYJ8tLPP9j/OAXlNSW
3MPtT7g/9uvoT/wSq2son5N1eKqetH+/khd5s/3n9Yj7gsiXmSX656ch5r7YbQ7wEuKTXtn0G/6V
LugPCHW8l+Dqnt2ryP9Re3bCS5gNNJrg0742hBucLkT89t1qh1d7xn7DPqM1RRAYhVi68h5Bxvz4
u6XWqIesK4DVuM+/F0CEy4cD1pcvoyXIO5ZHWA5lNL/vtONi3f9BB3WcpxQniled89BXUzW5uNbT
MVxoCS5/cxnZpx5tfAdeGDJlDfdUYHAkuxOJUfuMd11pPTROgJn2K1HPVRpNTWwdD2GAXEliQaU+
QSu/5kh2B6pafXYO+7iZcpEAuDDWMSwhTgEtk4dFFnhEpYTbQTn6IB7yveB/kaJA7xSluWUE2iDz
btc2lxZlzr7Oq3442P5FNlhsL636ZmbiDLc8v9ilQuYBA21objzY1ajbfMn9T04OBfLqqig7k9Pq
EoEi7Ejcvbh3c7n5S1XJNqpkEoUuEWgKJPuMX/GPrcbEPmvHwd09gYN7fCOwiddN/WDCf4mWwte9
Poqk5TGihP0uyS//D9K5u9gPjVd6E+pILQYH/52mz7RFcp0HslWeeje7C1rXcEkDvmc25oWatNeo
0AdHbRdqXo9meMK1FrA9aySWKaXW9yFFj1BFr9Y9rsMlcO5kY0LjkNg8J24prXnX0im7kX6gvo0X
cAc+WsCYwWuBtBbNYjPNn8ZDB3hoVkOkcpDtIE0eaoWQXRs/xO7VOGldSPe6fpe+KazEQ51j/1Yx
dBTxEoZtnpXUucIO3TNmjPk5vG1pymiIBxtGkMt5Gak3zyVbkSA/2rzlomgd1pw587EGFO5aK5Kq
XO5bpIxmUOEW49lKkF3jwgNLwgwwNAUHVaG3nLEmu6w3cwuhYMwQGafjCiylO9V5NSDYN8kte3u6
YRRSMM9UNoLhKUcQe3fZOPEUqsQgVXAo3MkVWsHXlwrqS7P/2T8Im+idiqSnXzsWWzGdOl+Y3wJT
k1WGh9VVVbHSG63ktBMhRnwnawEUXVy187uJtpfQm7rxXBOpegp2twexbMMYlrsmcCxtLwXZCr27
WZjG9FuG9+mWCK1ZdI0xL8a/CJU9dgbxRS1s92w5RxJEF7SYssgTrY147Nam9LqsCRmxrf1guGxv
AZYJrKtUpXh2D/xDs8uueBKjx1689PGzF4oWx6H7DShgI9jCIwG7xjGGoTD1OCjAzOicgBOFeuvd
hXQeEzy3QjFqbOxXVHaGIJj5WX2SF4w/Wsshb2AOT8rF/yl4U2QNBacJVq7FRSzl7Ee0JttBOsHk
8ASa1oBu03GMl2BREuFuHd1iyZx97CUfY4a9AGZ/wIrx0tOckfI1gjYlb379z5qxrPwEBQyA5tPQ
iap6xtBNfmq3hyt8EoHU5dhZiWY40VrV3puBqJxFOPoeyxazWPLP2jBCpuw0T3YmqzIm2zOF7q1w
lXSfqvWeRlvLg1ISUw899kQ5oR7eBiPFowr+Wb+ylM91XDdYP8Tx4kx04QyWefhXkTCu8/E7HITi
BfG9uSnwFkcqnGX3OxnkyA6nQeoDJLRWiD0h+lQ0V6WV0KIFDNKAeAOwJSfnjQkemC/9b3gBqgH2
imwhvXrx666EXGwF3rtPGLPfjRKBooMfKUzvLAmwfSab4b8Qro8dvmcOtAwY9PA9Cctzp3UnvCfY
enkEum2op/Fxu5dZOFusklt6kRg9rfKkAu6I1kV3ggUPdnklOGBZEnkKs56yjFqKM9rDsRz73dMY
ybBPSrHEvvyhh25iAG4Y/1FNAfWDV5ozgmdlnaMjv2Kv6W4FOl6vmUSAYroG2Tw6FQGst+USUpnP
jF6w1yRiX96ZXmpwkgoSr3PaOZEHW7+qXxsSV9dHjpZaF2odWu/3CoS1etwFtq5/XrZkF/Yo9kBK
1k15YlFK+Tb8NJQygfN7Eb136aH6iD7FxZfmgPjOLKpINQnuNjyJRenZ9cYIu9IJGLLnWxWosyRf
HeIz79qruFPJc6HswfUgKpelbzp2WAllS1RS1vdxQaGD5i5mE4+R5xlSw6HSMLLaoPNxSRYOpTqi
KiGD8HWuRCwN7WfHhiMnzEgcTU7nLcVT6xERvm7Rvd/UPf+BlSEWSFeYA86dGUIw0rSdR+oLlgUi
exsdXspNfBtQc4Ay6o2/Aaq8UEE6oQvPQG8M49gUytP1VtqkWK6yBs805/FSyPCjxIDFPzBGqFrs
/0W+TAsXhlghQqTsTEu2CGy3ihToDlgdJrvS+8GctoDvieFtnrXCDLHKZuUXRPKdjstjTm4KUIf3
XMh/yejhCWvnotGn2VhSFEmEAosgxZR3IqgG2UJzGe9FZDvI5+oGAI/VLS9JDaTcFmNvCtMHKj95
5zinJlZcnAzD2D4jQfxwGnW/cffLnofWtPPrM9emSs2hlQE52BHjXAYWOKu4Zg76QsZO43Pr6NOi
UfwN9LPgJok5uVEP6ZudijCp0T2zN+suWMgjT4BxPyTSBXR5UFxhpHU8/uPQcgKy8+bjBhfyadLW
dDuECFjLEaTNmJ1NGHiAC8fjFysHrcWfr5B47vS+jT242qmlSgyKtptdU1A/Yq7xX1+jZnqlmhxT
ZaEv80/HHWE0lCy6p1u8RRS4O9iUiM7bnGnTwZw9osZMhX2a8DXOkcCvO+52ihhOWkjZnGy0A6Bc
bZsSsLMpkdN7/a7VIt/rmlrx0c22EBP1CwRjcVwGyP3pqRNxGdwtNWz5R1JYUqlVuy8c8iMey/MQ
ZTb3poOVbrg5wHoKLUXw6vX7tiIRKYMFK4R19ZsK4Y/uQ7uL0FXM+3b9UFcsgchOBYCGNwNRLe/R
LoFAwmYQh+P5sbHNuz7u0B1lbR5d9qFq5OlC2cg1iD8VVlePv7HazrFNRNn3oxr0g3Y3PKrKGRjh
SLvmqN9dpGuJjo460pNxwGRAJayq6XefOTAXLz6HlbB7n7sDkr8HARK9P88kRDJHpMLOYzsstykE
vTOxiim3hhO2VsDGBfJ1WBpz5QYOsKqnqxTNWbtERT4/O/daAyyzSHGkfvMIZJFm+UQSEDyJ6yZ3
qialakFvyLYfkUHgnVjIUrHmHgEwGWAekU9eNFhorXPT/f42QNoFPu3lbR+4kLx+Czktr2QodB9Q
uDn8ZnafCfZfjD+rwhjNAFgFxxUf3JripMSWCZ2zMXq7RwR3+0CUKbhXrenf+1I+vJfy+/4eKQoG
VC2StNVMflWoM0xxJbOybGVjAn1nhX/CLe4awbFeb0eiQ2z8qXIF0+ofJ+mO7H1OfsYqHfip3Ma3
xM7W/YIVLJPFF0LfxMqHKQ5Utu9SXnnvOaLDnEnT08d31JjNRFufYHKH5jASI6ZcLBRoRXCMWEPo
OrkBJdSWo66V63EHPCv1ly7wY6bvzHsO+AwaT0kX1Hym6gO/1NukXRRocaT0kFHJw8gcXilrsY+M
nriN5CcAS38SEdeACR4MbNHwJVggdRs0dRvZXEmEtOPKW/vMIX/YkWKicKuKFHEXOEbQxljX9V4L
vvaYBXXNl7hEkR3ucsjeZsbuKXTHVpxVcGEQgrwJ9hEtO1nkIi1j+9Mt63cR40X/yaq3mZjMgN2H
eZXCcWibQr4zeBz/psvJGt6D3rJUycDINqO3sURl+XmlLo6iQRm0otDDs6O0PKbbIfUIyJf/uQKa
/xtxShuu51NTMT55C6HB2Lp4Jkiqgs5o0XXfu4f86Dv26TPRs03k0WqqGlV6mJlLuJ9i9u9zqefd
b30S+WHJbIUvFHTpeRQTMN8LgWA1v2Jg5Trbn2H9ucbuyRdeVnymy3pucArYT7rYuhYdLbQZf6Up
YTA2Kj9neKJ6DRg03oGmx7yjR3DjJoEIc8WcYM2ixrjOrKNqbCudxwUfTQbQzDYLtsrh3HrUIXzL
t//cY+6XFf6dbgW3MDrKy42tPWOmGWmheU5Lf24JShQuWJjW3QD3y087yUk8dlbPBF15PuYYXkNg
4GjtnzOXdVV+z1DPatCr4sDRpr/2OFzfKPVpnDn+FxpnVN8iTuvXnWYTBFSo2ivkAJuCsZFdk+48
qP1nRBJ5AGxl0fiHIklYageerNv30U5+HgM/c2iptzMkfFVKjmyymvZM//bx3uMR6wPzDYfWicCI
pRaxId83rnbzO2bfBTCK5SfaqblnozkmH2ZB6BToLEy26jKf3PIvWx0Lkr2T8gFaVzDyj9EH7FNK
1M/2cNtOHs3QqMNlCrpeLMxREs2o+4KlRpOCxV84bpAZLfx3oy4Hg98gzzHcbHeuQ6beaxshKWhZ
RQEgiK9pIkJpKU60p+tnO0ASiYh9KTBU1TCkahd4bNcv4m9OYbP8aSi48Byq7YTdsT9Wjf8Woo2F
AJJjRI+TuHQc8exNJz+q1+h32gZ/UxgzPmIa9KfnHyzMU2/8u4k69VuQ7AlYm8OuEm/bFLQauPBA
vQVtiHjSZF07uNVBqatGgI1avF7dW+g3bN+GmMGZ4Ppm4fsS0tfhgulB4a2ILCJK5wKG5QeDkLTQ
mrTRmNACS5ZbiVH0GCiEzdpQ5HToEKk+tOKiFJOg1FuSFAFnfo5FqSUUekqinqEwxhEpMVt/btQb
m3+VN8l5PF92qD7laEhwrGAddOLWrr1xb2oe8yOlb54Rg3oyWB68NKIo5u5rX2lxuYHbOmpwgTLT
xZEqqNtf3mD84l32KMjK+JXfTfG8gruhDiPH+k6ghDiAVNCmHZph2dDwOxp5phiLpPEFzX6oVk7D
jsuFhCRsga+j9t1B/5DKEI9+imnJUo6ajE4gexkaqDj77cdnvcle54tRrHrmN7qGkspuHM/amFf4
80qD+zOpiJOTg2Rx8EVageDxW2iHeSag7BV93WvKB2ls25SnE+7m1y382N+y/vI9OhC2uSe8qfOQ
Ok06bG1zcevVGLOBE+NC6wFFiQY/HB1At+Uj3ZaFlVVcXObdcOTGYb+HjjzaoaLDEu4QwCdzLEYT
fLztxftbv3lO4ENTqCZsXxE0+ay9KyJud/XxrbEJidCd53kbSGQ9oPsJ+OBYGOXzr9WDIxqHETms
n6p+nFO/jlMoOgPqEOetdgma2xWixETK/OWRVMnW2dimAARYABIZ+QZhwxiD55usW6uAjGqey4Oo
urxXUyaU2CzD+2cnOvL+KIHLIIX9Xao84OjouP5MNtK9N5NLe+oFh+bZhf+KvmRr1Z3tVwfw42tF
iQW3WNiUqlTPdsr+YckRHDE+nP7vgq4tWf9CSIRy+PA9t94u/1PnuQ7T5DrFvp45veoGokvpgXax
JinEtboi+nbOl/r8gafq2jokfLnp0tAI1Vddgm1uGG3phtdlQXBkfcykSqAcyAoQTOyOFCUCeSKF
EiNFK656Bnc/xvNQOreDKYdx2/2YRmZY7K5w1ZfKsOFnLe9aciK1uDGGC5irIctQeI4P1djJ5E6q
9K5LJqvnlUMQNPlNnt30UKxmHCXFpdN04/6iN/QNoh0JegQmgZtOpfSw8NKkdPV0rhEoSahb/C+X
5kP3KtTXLm71d6vHRT9DYog6innH7uVtdgzY/xEdoubA7Fwrot5b5FRiFzDdnGYMthk+EEhZLp/8
zeiPjs44zIZlUlQigJOc8cN/3Sjf2CttQJ2ouyTBw0Ctyksb/uWR0K2p22LrkgQ1puepEcFvwoM7
Rh8M5YDpJ7RTVYvVVFRxFSPNfpg2jaY7SNdf1seSkOKVbIs7KTLndlvK3D4Q8iEG5t9c7Pad2qQf
e2hpIj9hKjaKNpRU88V7KOAcsHqMJgIrE+EjIlRiiZ2pZwVw5UdRtv9wONANkueIWcdYRzsTws0j
+17HLkdWf99NnlLy1z3E5i5jHt7tVQkNEslNPUxYOxbmd0e+rcuYv9fNsrojUlj1eehbSevIJSCp
jVhIv7jL2POpVPYYMoGOy1BaDA3nwOVyh8/T4nvez0gB+iOaNtZGLzvSpEfQ1551gCaAligsE3aC
Y/O10LAgF3ob1fKNfqbkW2XcIJvZb9p81okNy2cHq6jjjR0Ecp9cCcEifI8iJuFhNlOMpGfRoZ4t
2RlVtFcSTKoMbeg7c1snxND4vAPqru2HTopZ57Owte9NUfWbfaFYQOOsUEjRWtOjfBrM+Z6kCQzY
XYq1ByyJiXNgMoEwoFRkiixCKAYcGQMWrT19acbTQT03D9vtAVL1jVbNdFUG5gKdTkmn4NKLYUGD
Td6QWtYbcwVnr9prFMAjD7Bxf74ANH1au5W3Kf7qHRhpcCXmhjyRYopwwCL3Kv0AD8eJhKf7wEue
faAjla7PJWHXdjHLttHQRKRNWkjVd5F664VuoyGmiM4Ir1gqQ0G2jEzijlE678ESeNkh1Sg+r1bf
Lh8TRE/QtQpe7ws5LCAocwgpVaroR06QoOGCSyx+yL5TWyEOntPMYROi+Y52Geie3DDadzryqDqb
g6PnccnP7wvv9pdNQkB8r4l5OCA924iVHRxwmad5qdkkiJSEA092vCLT0NHWt74epE84/IE41K7G
U3+Rzy36aW9R/gNcKDdlF+oSq2wqOCq/rV3FCNcNUwf5dkeegDL4UzhQ41VCvALoIUMJIi8vqk1L
LaEM576LRLoSrbWiGCPVoqOEfeAleleUJp4bBUwK9BQUDckjil9Exe85xtMlrI0n5yGeCViGccnH
TL0iVAujf/2xC8SLcK8tkEZcfQC1rvnd6WMEQbgJ6Ko0hStvkHic+bAvtnrV4QD7gMx0t/yHhcGx
UAWVdrmb3T+Q054x66t3MrOG5s/HXa9LCP1uV3XdPH19dMgIVmUnrvr60NttMm+K4lV1kxTDHDDG
PPeET/iV8kDukpCfLfJgGo8cKG4rMrI6SGDzK2qVqsR8SiCel2cDYOFI9nxLhgZ4RkR1ZlCJJUU2
9W5lxQlWTlmWW1bnKTG+R0L0zMqcPBSZ+jBindF82SpzH6Gh0eM+sNk6jPPKsJTKoLAfds8mc2OI
mW857530c03u/+oLZcrLl3VNN/kM2nXiC27AmzbNdJ8tdEQLZbnTZwhSI9Qip8QpFkF3scJgkUxT
FKXWMw97NQj7cPrz4pF7uh5SR33X9h+AXO3Ml4bqdaOCm4EILiwtCBto2CifUCPThKBuXYf4TX2u
Cx3Q6D2zo6v6OO7p/aADMkSDoyhGHmZdFOZhFBaqLAX7o/8z4hdNvBPKULIW/N4gcNqhZySlvgcP
VdaLqxLGC1Pt+vS+O133GJtK/3eC8qb6MN6o0+11fO+i3NbNMDXkpSMMBcWrvecWioDe5FNTqHc7
27UWwu9V9RSmSE6zHTzmusLpTOhfMjT8RwRFnpwDUaTLjyZ0snGubCQBn0QQUURo5y073OvZiXb5
VQgXX9XF7/YSwnurWk2B3+Bp7oSQYlWnDxvBbAZm7X+JDy8cmlLl09KqsSJR4eGughfd06HP8LhO
LyJ85Sb80tlWbg/YOCZZCfdD1QyzFEFakfM5gBlsjdelB+v9/x6gjE7C1evJN6TSaJ19F12zxK8t
sujOC/mu567bzfCruOJtZifiiohDTNpdA5RyhT/16bJUCTvWhX7hPuKjPND50Pbp2UovfxpTBM83
ROkMUIXEPqr++lur4eNGlQoH6Ehw4fvDbrIjwDUVEOJwrcCSyYNP5Npd0f7Bq7+5GDSy67vdNb0N
fETyoIkyu4Eh7em8n6cer7nyi7FDjBUjqq8MwY8Zo3/2F840/VOKjZ6OzlKZhqCM1RhxrBperJuD
52201O9BnUKAFCKHbrHOcrZbjPZ+JrrZpSnEWRCDPtiKHC0yfB+Vqzx277J5dbaco+2lpGCKkbFR
p0SigvpG6V9D1rW0JDWN/g1neoQqlUs3cAzae4i0w2XLXI1H1BgkPoxPHMp3T8/azbz2wDnfQON+
cYcQvHr3Pvb4+ASavEWu2JiFQfxn0VX2TRKsqd6eAiYw8i7W0va7ofzTw/83A/PQ74zKgrlR6thv
5lJq64dNEc3j9hKNh0qMrJOY8ichpw9OdZEHoiYPomQ5CvXCekO+u/loiYA9bJqkNQEhcaTZBaC9
+Jfih20Yfn0GbuTvZwihFSlcb7q7Pi3FJQG97jw+0gflMm667OvuLbUH1lE8mxFHLv/ohsrfQIJy
krwoC154ZY0gNzYW58rmAUztTWur9rlMwckEEvEjpHHl4ydZG9AZxBr9BZVQTJpZJeD36eZ/yna9
Xv62croP8kDxwkOuzSsUmYdIkeNPBCHOypNr6P+JWfZcORCFqPWINC09rzBNABNZHZiOUqbm7vQ0
0nhKk/9em3hVvcCixEXgcYgpEWAAklJIxmZ9RCEYOxNW+x0sFQggqhIPhaiL8aNx5zjANc0xNwxI
WA1XL2CgyTdOeUvy7sdGmLBStmRalcSfsR9pe7cVDOYIbGhw37lRAuDU3I52T6TXtPOK6I7ndOrR
l7uUSeLS9z7W97MjBONqlBsJgBwyRbHAe+hrUKBC6JcdO5jD0QCepEjCuNf+cNyk3vxKrlcjxSj+
dkX46mpGyVfQD3QxI8ndSv6HJOD7hzCT/as2wKZGb7pu0p5/xLDGWhXi9c50Nj+t3wMdRkwcngTq
fK+tPU1jPlS9in/9JSgWKqzKfoRc0ZSOEGfwqE/Tvo/e3h8rH2N6igferJef6cwyr9AtMJtxOhwV
MXMpccT15kYc/zAzp5YtKYM8M1DpjUIrJD0uYK8FTtbCDt0dNpwBrMXctYM/TeJj60zs9/quxKD/
VGGqwNvhNdba/AKI8jzOKWUUBNxb8eTyvhqlyfQBiZrzq2OcED4G8ed1oMz7kLpF/qvIv6HraXLv
zQYVH9wRy+45Npx9ktSH2sh0YA8/vlM5ajXdMNYohgvSidIJ2H2Hc/o/myP6OlJZXMjnnOAey/aA
cNJUmcbl1szsleqLUprIr+bDhSAkT6u4aSTCon9cZ8hyxpWH1ag0OZPRuTHUO2FW6FydW0MuGgsc
X/9NP/5A865wOlZ8wl/AdiY8WLve2rp/+5OlLtTPpwxyzgJFlqIlAder3dqd5Jti+03y+8xJOItz
Y1iih8xw3kB5ufIIUNnyB2+BLquzuhlpfpn0MzLxJlSIk3K5ZXhIunvx6LU0HmCXJho9Th5+tHUx
DKiA6PfmYdzo8i71VGvkZK/iGMzscEB5rxm7vpj+wKuNWTSCEuyxJ8KP5WSw41LbBbQ69aihNMlE
igBnVFEx14Zn+VUDh/RIIGrZmv06NcYtOmugeM7KrPMz6ay8bI81fORfmReWMPPtD6Mgb/nNMb+g
pOK2GxkbiVcToz8BvpNy+j6l++PzXuVke3rXqGtTsggKXn+I14unDyxsH/J8ukvzN9XEy9LmEr9H
sUbhCRa1f9zYT36gFbIYsGriP7v3LbelZ/8jgY+1DGyvDEKsgrggqIinahyRVgvZDc9hhLpMvA8F
rN8i1mqdlGvPVZINoqRpryasBJCW1pkOspo/h3TPIJQ7yFSOJgn+o6Ri/3/K2iHjWcvTdBzFCDDb
nhU/30LbHKYMik2OQy8qYLjFP9fkKjuN2s7YVyrytql9HMwmvN44/HlYfhddB1EO+cHafr16Sf0V
xTnPuNxKNKGlYKNRW9TMufcaK/QI2kMkrCAs8JxQyhbNJIuOlsberYFxHEPyUOK5jpBal+jK8JdA
xV0nAw6SuabbBTWskxY3cVUGAueTQIwkANOA6FRSTzu0xL90XDWtTnRlpH30ma6o0hBBUA1fsY0Y
/5uJ+P95IMgKQ7OwD8jnpx6VsM0iNdjVdhPWBxiccWfjGO+u/gON5UZCqFnNATdwOSzUOQ7RjoE6
szeZKZopO7mIwNe10Qy+lemJ4KQPFrjmK++RMLEmwyvpPxtVJiGJIN0B/Uam7w9vH+v7XSObYyh2
9QnaWDC2p/lqV2C2yBgzLwBL235uy4dJv2334xjMPJo0F3+lhTBHnmShFy/7lxW5xapcOmuPpJCQ
V/Pg3JRBxa2zDrBZLRec4EJ57m1y5kLGDP8+fOQkIRZ764sy3K8nOIeg5HmD1BCRPPUjfM4w8iMz
04fp/3yxbVZdzhdXCvMmO7p6iRwO7iYl2Wzz74mdqHTg+vALQl/49LmuWfedrbiJxnBHO3kBHPKO
+jzi2o2rEK+SqV9pEvabB4x2NC5BrazwkXElI8qK+E2/fodv5YdaqTeUZsrxdT8gcietVJ0rw5r7
BXX9s9mOVJ1Agg56kKVaPet1fnAq+CxqVohYvuA5RD4sMeTXphittQM5EOyh6B4JyIwMNY8yecmU
kgxErN0jKtqqupbHzQtUpuDR6UP+rJjLrCvrQdLelmlGu0lXS48BLCkeTkQlh9cN/0N9jfRxgPS7
um9ckzVujv/qpncXdHoDLl/Xx9FhZLPp0SoOt0tXqhPrqrOYLWsMiSi3h2SigeHleCc5PHiXCMkK
0q4yTFc3FT4mnT8ao3Ys1uIztoXTPkJLkLI3dLA4URW1pNOd5Fd7UwxbCsP5F6eVwRBoHG2W8gIK
W6hunDwer/UcMHfXfEGZGzOB0Kz4n/An67v4W0+9wNx0mcKF/1qo6EommIIgR80T0he75TVrVNan
gXHQWqhrzrH/1NZ4KS6bpmgRK/ES2PIHFp5SUQrpjdpMrszQasDlXFGTpKcx8oiMhj4yEwPB9gU2
anV/RSkDHVisNkKez4cbO6GIH1QVj2MuE70in7oNiA+3SWpZGYkMswajquD3W+3qJdRDJqKVV3f0
tWBrivyYeSv2J6KSuFEk7w4BOUA1swNQ4pIBRp3qsuVoB6yLAEtA82aij0gEn7LP2xOEJC82k/CD
POMiBVDYNxLz2TfQGuRaRUkfNIhaiDz49c8cfXuPDnsJZxsEOvKNsZw2vo04fWl+wn5577R5S2NE
qlGTFx7rACyT5Zbwl2rJRRU7BIlZgDwLHrkQzpB4zfnOYhvD5dSyaW4tSQS6qjgISIugGF6XUBO9
LonljP9AsMAg/7REAFjt6m4qqf8rBKAgompZLsX72HQFh1enlathL/lNiw7UlzenrCLjvJQ3muFH
3s0YjEuCowFsvRfqJbKTEo7dYLFDp4b8sSy1RcWsT6eNP1WzMBvyKnEzyz6ILfTC6pn97TRhrHea
f6RWcEbgNud1xkJsygYeaR1eeRNdJttsW7zpwyAABbJt7Yu/HmbIugTGRsSrRer1cu1HAzfIrd3y
0CNSIsPAg1ckzUBbAkOGTCvTKaIgbS6EZ0oeJZiTovVEAvGM6p4mSaNR3zgs33ZO1FXFMqPB/P+t
5RmMnnC+rEmgc37jKQc684tVNUrt6tCpeMutvfwwlsVhpEc9M6SPiWf6rr9tMCSc9ku6n9WP8BqP
QRN/AFSa8QHRNh1IsqFpOB6DCWmCaSZD6MXwMW7Ku5g3dlCWUdeh8tBOEydHDjbZJ8L6BNDyJouG
PKUFzAI6ryolDt9rs2qjliLEVGw4fl5dZNraJmEElAvJWAdSI7b30zGLtdUTkqRSpDKgIPPLSX8O
aF7cHrEqgDgHcQDrh7XjkOHE6RNa9sOwCCPNYQu+VXFHr+9CYIS1HRRqFLwRRy/hjpst2ULOso7v
nL514u7QLMPPyCnU29+dmqHBoJHL49Ar5PVYDyDGf8bO/SiXaGC4xLVADPgRlFzXS46fSm6tHD8N
7FgPA0AWZ7nF9MJefDREj/Ru3UluA73G8YrWZj0GQJZWr64AzOlRQ7OvYUriVT93EJcflbeqC7D7
Fw7+5SL1ByUd97JhvCzzC8RqwzrB1CaFNgsaYK1XTsHhstp5m14r8Pf2OPUffgWoFK57C01o5aYv
791SDPvURTC0gEiK6nch6Cz3EMbvJBP9onSDOXkW89DHi3+lbf4bu8TwXhmP6VkfiSQ/PSGfRgWV
JkFWsA9FMe4JnNrfchG1dgLP5wRJdUaEC1GWyb0jHPpo4j0hU2YBDwsaFlDakkVslyrillHsCfSF
+ZFIJmF4Jf/YuYi6aawZilMl0h2dhCutOY9ET8NYFpnYTom+SsATusiLjW6PAJZ76H5G6oZUd3tH
5CIsUT1OPChwDmLxig4GfcBRSmQWYBkl+TyxhHha6i+glLMvxpIvI2nt8s9VRUAYXCPF3Umx/TJi
2DLfjI6MzHUzo4VguhHTtUi79XsrmoEPs2Ku+n3htqUT+4SyMntQJV+63CFzuGi0XRZDfpRYJ2hX
F8DD9GCqNFnWch2eP4q38j2jJLJ7xnKudWCblkH8HYgtg1FCblPa3NzaBqyy07YcRvEk9L6I/HWd
2gWZe4yguGlV56YH4U+M0DddLruhongxT0I/LIzvFKhS8kih9fYhqIzVl/U5dUBShNxqEg2r3qJd
tGvYPWWx4G2sg//IjDceJ9loqTc+ez4DtfRCEKLH/KSaeVNFUe/aVmJ9UPn8wS2kXiVnZziU37UA
ChDPSFdwGJA4UbB+NOxIrT/3Xgzwg0Q2kQ1Ga1Ob5fmVs9MVgIuExTP+cEqenW1qRa7IxYuwl/M9
RFrFytZOD4U8O3BNOtDakbN+r255bbiuj/jW+Cy1NVljXe02W9suhx3TwqP/PRX+aaAHnE4mfr3l
azxTjwvgcdBT1ELCntjmYIs9SBrWkfY4oKKu36X56AILNinoOw5KiGeqgZSPOuajnUGuQdMVxP1E
udZz+uYJkouELBFkwbWNeLgWd8RTq3qVSl3sdc80q4ooVvE/4eA1C+9ZPn0RRc76aPWKPih6Div2
Bppid0YQbHaksCMaAAqNzPf8n32FEYcLFN1T46fUiDF0nDrKsg7L652RFvx4d9gH4AktlWUlhkbR
U+PYQrLjRuiRpfOGaUEMtSynhSsodO8DqVengL9+I6W1jcB7KDLXxsb5F/0VIFv6XvilX5lvHDB9
NjC76y1IheRDL07SxtvIXeus6BAWf+X8CMNzpDb8Dycmn2WLL8blU5mlHOykaqtdkT8nMHk7kb6r
byOK5914f0PnqRgAuNdQrqfbWsj/LDoKMZqMjnzry/FOgFqVNCQEvG9BqP+xPVgexmg9IKmJMtnO
fVz0nu4+pquIb2U2JHePddbEgAy6TzGoqBRRXjnCkB7Sl3VvSijNGvmAmJU+9TzU/azi1L23tta2
//Xk4/uM2wSyFpDMCyPmxtxP8jTvK28mHiyVCkBS4aZ7xd7kSATj9P9PPd5T9OdY2ge/BBJY0T3q
UrUOw4b7MOwGSAucf8e4M9Apgfts7hK2jd0nREfO6YsnzjTPYXUb9UDhC92ssKBq2t6ZB1HANhBW
kUq9skOXjwBTKPzfvAL8iHOygBvpI9siq4Y3lJ0rf47vVrXu8W3qAgI/Al1oHxr37mcIAwj5+Sl+
Puop/Dn9IcUXvXKiTeOjqGPpEVkvrr8V6H/3Ptxf9rTRQI8Oo8BWZvOq00w21mhkwtgOrWEqeXax
zfeumrm9TLr2eEaKK+v8w5CVHcr0uMJLEV43OkgkjlhnS3RSpOg2eov8zjmSke/8F240vchqR1U1
akX37DyoM1STYjCC63BsBCkXGDpYrdn8upCdOszYPgHUusHRKoegav7NtxPeV93u+uC1PDdT9kki
DbwQLNJrxlv+exJtnCfa6UnJuEsjfXKG6VCJoxRVexm2kIC/ZSlfA44M3XAYw8+Db+icuZXJFypX
dGztJXDcKXM8VNVjsI19G1Aa5YzbZcLbUfOazhLlE/Qyx2bNiPJc0TkW69K4vm108GCN56IJJ41Z
VihHr8kx9davFkYuBB85HDbXjLg5cFqzg6g8JeRk0uOC22XLl+0nntO5VJesL1g952sgjwDbsP4v
OuskQLj6/sM3E4AsmLEMVDn1uvNH94vF7QW/YlMmt9/xKug7vRatzTIIOSGtJNCbAW9srZMFgesX
AHFq9K7WHBv3dJ5jMicHDMNJ4eedbhIetRbzU2HvybyAKFrq8SH3JZwAn+n+0NH4GKi6Sh9xJYuB
8h/n5gemdV6c7HriE1+uZJeTmh8iYYNOVgLeZR2DfQ93rc+nsj7hFS9+6xTePsG980kFRgO/s7vw
w/XTINfEqnbmEKkeAk1s9MkvgOE0DPM/+Q8KIBWVXSSE3JRnTSO83gO9YB3LKaYNqNCAV16Nr+lF
bUGhyPJeN42sZJbl3J+7m9muvvp0Qvqc4N/7+oXTHRBwjPvjj+pxIAK4W+CGYiCr9kxFIRrzf7ak
HAmk5p87cC9r3R0fh/UUfDtg6hKHVQJQhDOSvlb7+TlsRw/goTJ5Hf6ydYPqd9dvmx15oFAezIez
NVFeRRPRY0Ykk7ZsycJrpo2PP35qDoRQ9UNT/RJ/94jh1Wnml/FcNZZaIblR6moHl2O9YBMKQiAh
d7CmE4WTr+HnWZCjlxemqLkNV3m5T/3HMJ0hqqmeZryG2FlaY0xQveXumCRwYBVMNNUn6rlRvZ2h
+srwvLIRpSOLQJ4xhLLpz4j0cN2y63FtjtpxVVvRW5D+kffJiPKUZrf/Uyyi3GEPPe6tLEyG5G0a
yKAKiM4bAbjMocsYvI8yxJkW58nqN/rk6rmpTLXsni1UCEvX3EISXp0XRmsYZYTPOs58s3lrFPch
/r6s4J+4XjN/PFagfW99c8w2MIwUpdReV0XctwtsfNGOEdxCNnjslRYpsNVXAk3++285LgGaI8tP
xxAnqh/6pWoWE/uQC2x4v3oYv+PMOgvMVh+Qgi+xPeiOKFRMgCGT5+JGB0xJDzIyGoLVCt2xxSjV
1vLPPXkOpyvi5KmROyy/QlleOoZ41m4ilf7DcwnDZ3fO2ac1Vnxsh0j6RFjTkeuVnhGp2ZiLxPaF
JMOhNaDtjFfhOfkH6GNC8mWd4cmKIswGGscag7HvmMIy/AaWWmwaqHduGkK3H09fxydBg3Lurl3Q
hYq1yXkuDWsT2sBlmP2vTWpg82pJLZistsKB11qFYcobh7YkbCAW9ochqGy3cUY5FhUcm/a2CGqr
p/QB7yUVe7LGeAPJIhZNFp1yVR7WgvQOnKjvyhAFsrVVPGYW3szgmkfPNosPmjoS+s0twidnHQc2
Kfi4S9fpv+bQ+KqBMOM5h3Oh+r1vZp2sJa2h2yb8rb1hO47MgroLirh93xaa4ySJ8SKh42XgpnJK
SMhcJmy8KzyFMkAS9c0bexBxj2wBNk2V9YqJdCIEX+jgcox9PTb36cnbIbx0+/OxJFznixII9LRm
+CA7jjkFHSL08r23K6oGp/GrRUymOIuc56f+ZDkWyCWmjn9ShQB5znCiKtulHfarxaEZq1R4pTxw
oWjpwwI24pQwF7yWCuRlix3KJqjGXfSXpuJMUzjOzfuVDbPin8mGS9YtXUs6XuIbGAZsergmE8VG
fmAZT36PAcq+gU7nss22yaDX+11+B90T9GtOnhgbrZ+AWqraTNR50H02jJRXNJ93wJ4oiwGrRXDC
26epygDqPg2Yur73125tfaM29Tw30d+mLj2IcrpJnvpaItD/mDKPlnAAKKtZo0y+j+e0R/Q+53M7
08hWO7fb2cbJ3PUTkgqeEMKJShq0BaYOr2l1WMTeYrke/PUn/tuZoisDAfAiJU8Zg9ev5pDL0sIT
lMmoA+i95wrZCqCaUJ0q0oV0VcltMf9SlVNzz8sl9Dq0eDycg5AcSa0wFWrxj3aPwUNHh1XUVG3E
YeqL/Ugc9Nya3hPESC4mBNbb8mXKFkx0RquqmzrIDYZXnxVW0bJdni9VDROSFT3D4W7zNQlkIFbh
SEG2/IbZLgyQ+42f3uWol4Rmd1ko2D5qLnku0eMmoJAaMhTjhuVPCRsdsSt6NQk0+0T4olPtq2Fm
sNYo6e/AkCyQKwOR3hXFLy4aQUGJMgqh7dtuWlQmvWa3S0XJ+m9PLArzLfB7wC51xaDYT6pOloFZ
V5pXkHGdxvKXi0awFEu4sk72fXxWuhuDPccV27ybUAs49WliYPVhAd0XhVZH2WNOIxyf/awpJHcj
asuKGWHlkQAw/yDxFudX2aFnxStEas/t0VT8W+k8d8P7EiCo+McCIqM56h9OkG1OSZokcoqsxw/R
8yQGziI2wOWFLMj128wPLilaqvLxsWoBWfB2S9ddRoRIVSoYTJ5TLRizVobEe/HGIjXqERjI0ucC
u2f+CUhVBePywwcqEIoyokkOSECWBrNQ80Bh9iZrKsHA7+WF+CEIFmnAfIkhay/u/epRdEMTx42a
Z4UroUd7qiCR10+0bTB0pFj8Z5IeqcHC5S88oaxZ1F+bB3KH6C3X57kKHaMIraeNE68SOdGGmaPf
DFTNsx+wwOKShwq7YCMsdWaWM2cjbaHpA9e0TxcUzMeCF8wRk+2T9b/ZsVVMQcRffPTircvOeWNv
YnlEp81rrHc8WTKQi+K2DFLr+hIj8oLLxdAaNyiC9OUWrfp5rFWMvBpResmpYGGdMPRBRSAZ7CcV
nj8TibnWbKTxKOPI8dvuioGtg/AAHuSNNKg6Fbp00tUrMWJyAJeS5H+pU5p0mnDcudlPARbr1HHN
O+cnz03bdf8q4INVxGgzx/gMvoclXAUloa3CH3iHPwsKAD5hNhWz0HvHNjwQBVPatXMlUpro7nvB
yK+Uk+QXt8SpWIoSZdBpclge3X4YOcyx3zMa+2g/OW5oX4rJ4AL4hKpoa+SjtSMggIv9pv9MyJyR
4B2cZR8lKSPydHsVBAjgRcJG4E/Bb4wQ5Qufuv+XQ644r2jQ97NHWkdq/vDhthmCfjJwaWu8CWXl
X/dL9fAgLa0Fmrkp6jkFZc5q/v9kRwqp+uiq9qL9hKJb+xiJCTkPBx43e3sZVSUJhK2ge1Xfld3r
YCd9jBikxWwM5D+iVpIu7Zu4ENdwzpdqEd+ddS5/azitdIGYm4pODWe8m+Z5ed7UP0jOFS4Fdebd
o0X3nexe2/OOMtD/fylyhWC+23iMDZvXSpu1snmgGccGNx/ohLblGiFxldScqR+dXwaZQQHxtmOB
zdXJc+ufoRegATQt9zuCLhBDpKtOM8GovHxO5jBDZV3JLVjjobYLqiu/X842Rb04UnN3zgWbg9cL
8oJ9q0YpmvtLhMy+PlPR0pFD1s4U0meLr4ha5SfvrZNpLS93slUgyovHc/gTFW9K8l7IK1Yw7pv5
25vm95UNUfW83QrqEbYfVIEH26MU9pSGGMDBO1VpGbUdxs1uttySYxCNFEO/+9gFOPt90gCEbY5O
S/4U3gAoPwpf4gYLNl9jnAinvtm/3Z8B1waG7EYX4vw+ZX/MmlcaEulKYxmL0yg6SPRpuAEevTDP
cFQOjXiNP6/wJHZudRWWHX6rnUOXgnYNuGcKibZFbR+pnJA1nDVW8t7zNuWgHis1K6dnBiqWoDBL
2p3NBcj8UxUeSfA6BN873pWG9HzLx0TUasT9cToFDnehg3GNRw0Fa1VgMWeZ1WxTTV8SIcn8CV9B
kTkczo/ZvMAhw4g7nMKJUjINyNLyTRSp2c6H2292K3u7drTnrKGAr8sRjfS0MfXd2PcacM2Cx/4t
rKhBQtcQ7YNle1Cpk2S2hQIHCWNk+x4UMQjg9pYNQDa61n3yO6dKUkyx76kL2oPE63tIlrP6pile
zTRqKh0c2A1AiAMbMuH9lYWheALMYkAUEHLwsD+dZIEMQvuClytBE6qRvoekFqxd0T0gcFt4MuKe
Wegtm5KWRAs0CO9irzDTNNISMf0NDETP40W3a1ofN7DmU9jMH2zOWjAe2aME+BEKlhuQXNF5G4CO
189NwMDD2pJs+VGyY0FmI42mmeasRew135c10rO84hmjpACCyhV3m7GrVvEnP+M4zflpae1n2dHV
D6y/zxMUJi+L3HZKQu+Q6PGhNO5DtNgbkwrHiEAREIHmV/ZZtNQixmNdABAygR3jJ7Bauu3wrheG
E+mrsjsYi+iY9EXo7TLixWtLVaEud3m1XjGLg7hhwv0N7qqC4WWvgCXq1x3vBMNBBuPc/HsZMqii
0GAD9cmjKCFcZX6o29e5jMvJNEIYPhMXMjNPjKHLKWXjjj2uC/hPpB0k/Z13+LxUlHY65GZyhy2F
U6l2OE1r9/0rfXwjbA84adzIsLR9n/lMjA40THkZXlT8FP1kxmtfk4Ho98CyXZ3OhnQT6vVhLXBJ
ctEoAgMngXUB9XY7kA5ZQgycsDPnz0G8UWnYmb/eOzrWSRJ0/oj/jWP3PLTbeWUZT05iJ56KFww+
vKw6mzco/xVH7uUoP6lEuFnaid8+Y6irLCXY/VXOOxjcPobJWecQ48tGWraVLpLSA3TT1HAY7Ra1
KHh6/5HHY6WDEaHuRJ+/NaZZFMQ29HqEyzwFU+UL8yR8kZ+a81e+DqJkltpYWF5aZiBS56LaAIG5
+Z9S8MJXdiwBnqtdYMI42alpBedbZzXdvlzOZnT89Xe/KelcFHAvZ7qKITpjRM9a7T5YvQ4U3wp6
FatSJ0YI6yyqMezdoTfHQQgt+w018YFkxHiGtT090+vJjps9Y6dKVljBbN8sOKVt3UuMhXx3kvdO
QHIE2knBNHk9pA6YV1cYqRZSj+8sRzQniL3Nfqh8EjPMV26vzBh1c0UCufy81AZ50uSbknMkB7cq
9I6iWx7gmsKVrrQdorvvO4TIqVNqObImaR6Gi0KZZOOyhEXWyAbm/P/HbIAQa3e23/+uNit3fMuN
hrDP6TDZVHmRu0c9urcSO3xu9ibO8jry4yfO84BVbqxfAierepUa/+2x0Vspf/6NtqmPklBJL8S4
EO+FbwNl6eLCtnj85MPda5Fka3GID3qfWS95G8Sq7rnk6GSb/s1byy6WOjQWB3YRGiWX9jDz9Bwd
Qr6Q7vNqATUCIpwnH8sThKdin+LszaNnp0UgsiPEvWMvqZN1PBrI1wAkJZJJ9j1sBOH+4P0WEyFK
Jb3IwlPkDdsYzqWJZCJseKRBFYfuQ6oS3+OidXObpdb+Sy+Jfz+clBxooF2tfLYE2Ui9dy0tuLvb
PCNmkcfls8AyNdTGO/NTiRAGHZ+fWB2bOdX9fzxe/lwBx2LPTgEaH4NKUDPKsDX++bBUmQC2HNES
zwdTERIcSFdZqEdLxkM+pgyXsodRxsfpKtpSbmgUQ0M+ceBd1qG4RrcjDxtTItehIFlITIiEKwCP
+b4s32lJf/LveuryPPjXnEYokH4VYlzkNLa6RMqWDVmO7iPyMwcrr4PmpofnksjYmwUFMqjAs3F5
dao82IqAYfxr5wjMx1Si9SZzAYTDWQLRBoiAhRu9aS5mGIK2bQYatG0TDb8vKCFA5xi844/99W5j
wi+nIYt1SvlXVh+lJ934yd/AVHS6onXx/VwFk8yuO7ML3UOg4UQpk4L6T7gDijuHRCPsC4gT50L5
1P7DI1MzuYMrL/On8mbQYolUbZr6wl8M5AuDijQB+yuK1uKjzAu4MypsdhfCw1SPbPD965issePY
Jsjgy+XS2yogVauClvyS2T1GL5n7A9jgD+4gazW59oGfnllgsnb+Tfrn3s9jkLh5fod4Dj3JIe8U
cprjWVjzqYrdjwdXMQf8qwY2iWNQGSsIHDa4zytJmaxw/NYt/3Ct5p4iba8FamQHJ4gzmpcTmY2A
oC6xeyTIgjDtsI8p/655YXBZwawghci6h0S1sXa+CFDK46MN217vWMFfe7846cDtGVpkuN3hyf3a
dbe2QVlcUwtTr1qLnOV7dU2T4pLgoHaTrAyllZTYMJt2NK1JKqjyyBNjKCqIz4MNLtBcHwtF+lhm
PfbjU1AOI4Ny7n0bSO3TFyFGnaSb6DgAEFawqQJfoeRotvNei/8KiXlQKlzfgDmyWjUDuJOvpk9Y
e7Zowf61ASBTc3NY/hQtiiGLpCYLiGgJ7vP3JwkaaAzCCsV4yZk8nVF+kfqDvNqCDKkx2M8khuuc
h+cdD6sD66qBYbPPCTbkiMFrWeXfk6E+h3wr8lR1a307wCfxIzdnM812gQ6GJ7QGxJleeoZb02J+
442ZSty6P7jiOOdDSUK9gByyKlRYU6mAEb6tsRbS9PCbq+cflGfG0bCPOk2+veobDPbyOHRrHw+a
d+EbXQI8uVpBJpefD/w6fNQ35upgjeKIvHQp9TRxOAJiOyztHv55MfcsZqeAyJtdbyo6wrt7G+gD
OSqR12pNGPR1S6yDoKMU5QbN4/n0K4pIGenDUXqU5S4BjGtFhx7i0VWjfkeM+RUHq7a9XTV6CQlz
gjggk4BSVDw6KwtsB51DeK/DrOU1HJdPl/ic5TuauuuKTrGMWh7UwI/pQnXLIwhnsG2ElPU36QqH
/vetxAaalwbzUjvRYjWP5bJVa8lKH+iseya5y7lL9zRrPXwKbJQOSC2M1dM8FRx6F1OLOfGcxLDE
z5rMoy4CjTbwH4N92+y2GuVSgQ+SWJ2pVFRzxyb5XGeWn9MeRMo6tkVLC3cQYQvia4NqP3Ld568b
78QT/UY8BZhA18+lM+ED6O5+PqXIb/6U3PpoWzPozEMPHCwgpVG3DcmamWpU9sMToUtdGZMluFnR
WkUtGJ74ieVf7deCVlDo31dTuXjrmR3LCxyL348lOS32rtQZs/KUJS3KArT+6UHEhysiQ1v6Z9Nf
hi4po4xLfesu2OgaBPFa/n8aqcM+6PU/8lE7CjDfFImFPyTuA/FiHj+seqTfAmL7Hn+sxQAPucyA
O27DNoDSWUvjDHDnbpgcIHq1UbZwn6LmxKoxHoAp7M8+ABQHdipXttjtNgYWMAwrLleSg0m/cK1r
sadxY/rzb4hZqy65AdVz3UxWFudB9TLPc24sYoCjOujJZ18T0heDhPfLYtiktrax8wYYsPUurBaW
Rj4Od42l4joCvVjmTlnHeNb7TmwFuS3ffMsdQ/uncJABGApYm4Gosvd47jRN0+/sZRBZpG6gd/uX
OX7cIFEQQW1uq8aNX7NEq0rKp4P42jYefcYaIYyw3XxBazJrWPX/1vHev+RCUJbzMW/ZKSwstmll
HdezTZvREtMSMFSvVIH+oH+TA2nJj4gj1RVe/iDzaWmr0lSsMpzvlRTog/nJf8/E1GSTF/XDe6Ln
4u+fxFViJ5wu7T/2dfUdBNJ/Bp4YJszazDv0q5qLLI8Ay3lq7c0WUzVsqzJx0zNNMYSYmY0aRBcE
dDZmlU1Y+SKa0RLYJCBMsHNvCKcOc+N/3r3Lpy0uAeBey35ofrEr/x6cCbHnvGi6CftUhoegHDb8
8iCf9wYHw41mA8QUBqHSfgK4fJVwDfON7ULHpbenWZlm66d22duly4N4xSA7M7/PxCkyxiL1RXZ5
3dqE1/BJQBxKCJyKTFvGwQodMSL+3K7yBrw39rMJN71DcxWZ54G1qdGbB0wjd9DBbVokNcgxaQep
HN8slQUA5+d5tqbnqnafpCFpN6SLVUpK9gyQZKAphl3IvXR84ujsXdg5Fu7sBBhAi01FrYWumdWA
ZEtgdBvMRnPGJi6t9oMOTcUeW33lDDW2rcLO0yJKtuKfR1cCuazBPwT9yQVNyDWEyouqM2bUuGif
FtHbF08ECyccKn2LK4YE0IwXn4Ukug6K2DGaPs29vK7xy11Wou3U3/v6PBpZJ0uXJVEjGizP66wD
RIeMoCvgW5HT/mJ54BXrnbV9ZQMJhiXJGByCZCLFeabXc274PKJj0qKwTbbjpxSnmuXk6Gp2WK64
RDQ0hwyH6GnIxVnE2uQ9iyLBDfonwb73gVqtdyNLRNBxpfXgcA+6f/cLFRje987FWdz6ROVAklK7
npii3er17WxWwbJYPolgAOGyqGtv2nlMG0CHwNcN3mPTfr3aKDlyGMmGFcOzGpGi/IxmAbdeOXlc
1gwmuATBW+DINxQMKj2PyXAeyLQ+Pgwyfy4ZciB7P2S3OOyACwNkp1kjf+KbQWmPsikJXnbB1oX5
NO6MolJ5ycQrjUipi5DGbDdb8bfKLA7Q7tTo1HDlLsdBPI78OmOXedhsT1u6uM1h4WB+KfTscZYn
5gUDcpuixrJFYeBRexT+dBBnY8IcSlo+qCQRx+WmDvZqNzZH+a95HTE6JpsGnlhTRgf9KG3s0t76
tqWb44OtVhHAwJfGmJ+FCYQkBfLXUygVir287kQvhToE6ZQN3iClQ+jFsTTQx1aOZUUJPWfmZ+oq
nqBd4qj7W9VFqRz0WX1IFzZPjJCWCY68kAe/MMpNjtVPudxlRRRptGpOehiRldh5QM4N5+Af6Cwn
qZFdXuctxkmD4Q7FgbFZKv8RID4+D7UoAOaQnRVRZlsLt92918n8UFtqdyrqO68H3R6pkTABb2rR
8rMzvGR1ZyesDgp/zhQd+1bfBuT8jM/2HXg7B5Jkf0ehADouB1q+lZv5v+JjIdKK0JftPScwuy99
Hq2jXr2eCqwr5GXuouGN5Pycl0Cq0VH7q+cbN5M2xU7ebmJxLsVyPtSWn/HHF9NXhc1UeL8Fk+1I
ZOZyxW88VUYQrGrCUxauyiHoyGXINVIGL2cHg105vebkk+plTxFgON32v1LoE1I6+95g+PJ9mpBB
LUFg22F0Hn+OE7PXQ+9faA0jHVcJEN3U0vHYdcAj1YDDGR7QhEufl5EYZztOPcbKCP/D3EPDyTHa
rfZWhaplDck+VwwJOmcbq0tBCmcpj3uKgBY58w+4QUMAOXtqVGpxIsXz36DF0kPm5N801dexF/yA
P6K0BdW0qhr9fbvdXbSS9cZNko8Fe1n356MdkrRG63Gx6mcG8uc155Hn+RXXwc+Mle4EzPErrgGj
YQNi2hs3FQOoR9b4Fr6HgSxxUgpctQwr7af4LCg1FTI3PednstraKG906V0T8ZxaebmlEeva/5f1
jwJXM1km4Lx8NWX7yhpgQCyMk5boB0o/6EloeDPFaViO3ubIwsC8JB9Oy7FR3XTjUpPZWFInS5r7
p6UIRG8nfwi0WJV6R5nB6YNkyF4i+mYX2/tPfIHbqdEo2wFkhIcq/VvJE9SHFXSFHfPheG9VTo25
S81mGoKZjrZlrGyp7MOYOAB0n6C/W0QUHo0L/GdAj0VmMTNm+XIP99w2lo6Iqi9tzSJqD3zVr7/n
1qkhc+TGT7i19LXXrFJ2y3N4tGIPMf8w3KRHRh6NSDDWHfJEUQweyQMEMfgFNQcMNa78sjtc4dJs
R8IMkuInSiLq9Ye/Y095l7PZQJAxH6nd+IsJSWTxwRexaZj+aUbrJ65nRQHrLb5jGwaYFK2cpzQD
EaUGJDmtUYaXvbE6DKjTgmosq8u/EOWJSvJ81xTf1jOxAajANFpezCKyMxPEsf0F+Oqo2nXPfG4n
l4VmTmMspOajdQRRPcBWbCTCdvWhg0H8Cgmu7uXHHSMonO2kubv7OOCC5wUXP+VL7dcSXoc8Px+/
Brn48QLcJuqyqt2JETIYoRhaQvx3fvgruKFesx3JNxlDI5RnWRbjONZ/8+3YwUKBGPP8QeS7geD+
+xiD3I+AYggJYWJj667Rj9/sbtGUVn+2LaGRr9ShDi37vQp5e1puW3+P+y5mtBgeJ8xXYHS1CFXM
Q6xWc+BXQ7wqYlQ75Zv31DhAziiDatk1NAPXu/nDXecOoKsaxkxPFJJBkddLb2SMA2rTAp6huC1d
Lfnihl3VWRjAMQK/QgjvF/uTez5JZsc1BFbdgaAVYXmxok9r7nVPx6YxcgIGZ80b+tQ+T97hBn9Y
tvtfWD1Jsl5pzOY/wdzde4nTvKa4a7NTiS7Yz8ihKdh08jI3du7Xi8cy3nowwsgsNRBAFG6/uBsM
3RNAihE1qofxSFyG1FAgC8qTSOoweiW5RKqiLLMZsEED0Rkhnw4RW17eA/zbmkLeHnSFMirG/T2G
XP3oryMVXyDpKuvasFfb5fpAnzurRy8xqDGTmlWawyHk+y2iPFlf2OlMaMODAamOHYC0J048J14P
biExuKFIalq+3GX6h1AwR0NXXG1BjLutTXO1refrruD02tFM8UUxrgtM/chbm5AWCHbRGOFWbqMf
sGSpNF91Bxe/hH1DsQbU5gLBJCh3abvML7L7irzHdr+kzJHfCFq+zi5JQ4ptB9/iIWBdp1wxxy+3
FCEMcp+9ArPBRyvhM1ITkP9qtnMdret4wmsXTH3Tpk9lNLrG+SOJMdvNZLyZgW1x9Zv1x9daaOJg
zjbw59hHGu/gDAxw4d2hoQUcC5Gm3sqt9v1PmhD1uCsyv299o54W/TDG5b88EBwW37ZiG34AkPe7
boGBEgvY1p2EgvchjMV5Lw9axYSZP1tZ+4k/i7Ksl3yYURWplRIk0+rmRPHirNfRPqtaLXBTa3Bl
UdgzOo57Y54LAmHlyPEJ1gYh2utVOg0W7lPLyUF733RLT3z9VOvrKQhHqx9zEu2sfrVeY9a+gS/4
5LArXMKDa789gSXVBmGFNYAIaCh+2a5a8o0cTXVWur7gIhETtmrfGQYUoODKraXa2OGfNEr61ehP
OzTZrLN4TPuTarH6N1OTEx0QgRoPxgQHyQwYuFHaN8Eb6KBDVuwcda1nMaZEYMYku5+pbBmgUaUQ
VHKkrqQhdfQLKEFGmTHAL0B8+5gjqVXwtKrPJYYFQTv5r8YgwLj5RZ1UObtV8O5Lp0fx+D4t5ch2
OYvBmyLLc8yhvrmAxtEAWv2+VvtmvT3Ch0ubLoWqWcVlwWig5KWkmtbCADBFAd+rq21oePzWiYOI
iCZ5eX/9s5UvLx47ZmFT0/KrtnM8zc+3QhIqbHw4Y2TskWMP9scZX4UhcOt2RutRzGGJqQRnC5Zb
WXuWThrhbgr25tJFnf1bRWZjDlpVI9PrafmQhrWQJYWEj1SPqrhH7upDQy4mw43ZE0lMO+yBkHbO
IkCQjNPFNQK0rn/YYJZhVYOccaGpBFuq9UtWm5V0DLqpOo/fgSQHRSKZ7M2RLinOYdKNaNgTefQA
Bq0m157E4yywa9hjWcPdhQN1K3TGJZE0Fn0+oKxNaN14xZhgStN61Z8i9YEwRgj2PVlYyawC1DV+
87xlIQIe7DccsiGY/LgJVgVFBhFPyoKQRzwCzpb4nbLctpg/6JYCpvk2zohDw14bUXsKmKkEervy
Jqq/JbJNRdHxDBCcuWYJkcU0rHjwIvdDjgcycVI3hHyL4CzKUIrnH+NB+WJSApdHKH8NJTBf6VXJ
7V2pjKbQ8vKZZm0yWqAB1SNERV8UCHr72Z4hHSM2WpgWvHR3QMsxsrz9QwhJ9RXd72AYwb6qZl+V
End64ibPHjQz/cA64eh0N+Ycf1L4J/vUnK1PODyCVNFVO/S230h9ekaCvif2yf+ltT7xWzaIUDU5
RCjR7A0+06515k5VoFQTZO/1HFMUirrlZRZ/KElcPY/ENQ6SX7fxxfL6tjQN4BlExcia+BTBwK/j
YFm8tfqCTVmgcJxdz2t4c+3VP6IhLOm1gKb3ouL941t4HdsDMEHmyFIlflxZPb6+KOb4h5iq+4cE
9/OfIkzM0mcIyaNdMPftkSAXiZ58V4PibCAbMAFSqFnHzE70JVl96d2RFM4D+MgQhP1nrx7JX41+
DGUGbMQfrZFlSrqoCNRvrDQN+7iYcyM5CLFKQaftMpCm6QhG5QR1saptyDD6SJ8kQNGsjgbz0lEo
rIUoLfta6mzaL9g40KZsMu86s/GZ51lvDquAc+vXvyDKSD3ANBRZevV2kslMCyqSyfae6gG7Yozf
q/kcqXbqKp+0SxtaLroBwvApnNrOZUWAJFJG+WbASV/W9Ct3726FvE44xQvQoftL5z43MrYb86ML
2Dg0W4m5Q3VLhPGJ42NichYgv4t00+YvRi/6kH5erGddpNQxGf3RGkwvu7nqFXzNvGI8AS3KUFnz
7MT8Hd7xTdD1XKEyEceNBn1//HME3Roq4BlqNVS8C11AkhXMV++CRBJRgFrO8VqeCDfhxp+kTkYf
Zgf/REeLDKOB5RgaxXgbrvEpPKPyJMQ13fP4sK1YpqLzu6YGvZyzZn6zPLKCTZlmmemuGB4oqeH6
tbSmoddGA++dc41Yx23XyhChN1Yr0CD7cFjdNTNQ3R+mqJvZrgBMZ1y3uT7AufuXKzDIeJSeF6AF
oCV4i03Z0s9KsWWbSqwd8/xTtvrS/+a+sFI7jZpZWn3kQm+z9MaL5rpQUju0mRmDuNCDOSwzs0VH
zqUcSpV/YitxlTJGBlb6/QbA6eRUmdsmNRl6giH6mPDmYkF0Vmdt0e3Q+PFkjlDu7LFjs4RwnUGk
SsE/LKu4fS1RoaOclzxOVYBQ7msEydDhgeLo+tInE5wttQ4yk6Wy/ULibPmQDcDzaW4tjQBMbu/7
hus+7rQ99CsH2r3qF2EvzkPe9CApIqD7IdjLhen/8A/wY0mUZ4zMAoKnGG+h+5Q+6nMneMHWogFd
+EyB+GhbqtwrMKHH9/vfTt87yXuGTFpaZkVpaVtR8t1B5f6MGUD77lV+vrwZr4j2C7yW18Mv5ftd
e/UehLANRHtDRJSC1yfAJQMVkz1jzmOSae12w8joch+vjbq+A0OOPdpYvuGb6SziRn+yAym+3LPE
tnrByrlvfBUGBs+rAHItoxFyfjrn2YONyKypmRGIv7ncPGa6wVHIVibEpjxD9qP4NaWlatlV9ZKt
gLvS2Ywq9TD+cKj7QGCK7hidd+i5qeByo+SthTFenPMT0PzkiRT+LH1zMFWA/PI/CbPVRrYDQyoT
mxYz6r//f45xg1Ee7XUYcI7wv607hGwmgCx0hmtiShejIeQXQMt/XWjg5IUzC+JSVXg8PLWQzmMp
px+wO/yjR/K4lqXrfr2LG677SIb0xNpuxv0Sf8v6afyowdfrWua6oLzTH70VSxTXPnge4qgUFlm0
XrGb7WBDrpdqcRxWHR5Xw9PlF4va2Q8MWgJTMDTdC2KGG7JU9/Fs/ARY6ynCnwD5RUo8uXUaa7Bm
MdkYOpF9uD44KVOSWCd/5kPS/3DkcEAGiv5SLncTNRPq26HhzVDKb3J98sp69RCffcDBceGDIlMO
bI1rMmrxzEp4znQtyB8RmWzoB6OQuXSm8p7K51JG4eYs3zbgMs2KsRf6yFaqacAHd9e2WLM1FmIw
urTgg5UR1zOYxRBOqwmV7m1TKZOG/FQfa9vcY4B0GJE+LuQkg6vBKdjTh/BZYXYOzuLETGKbV+n0
6eidEeMM236XZOkXeONYskil2iR7ygifiORW2wSx4mOb7WTMMjpPY0iVQ9WXAXYezoFQms1F7wWX
ZjNgcnk02etfb9YIiOsuuk1Ox3zCJctbb4IQ7pQ7FLVeoqW2m8fWNEdnVQe473MkyzgzhRRVUSPk
WOanjKAtKUbzTrRioRt5tV5FlMrLwYr5kBXLtYTnOqL5b5Z9IsmwzDPk9HCidY/zqrIHczqbHCMr
5AoGl1RCSS37PzKYha01p3PZZyV+0+6IAq2UA0yAgWqk2Jf1mYlbia+KSGAulR1OwkkGhdjoUdkw
3UwtriPkaGf8oty3DbUxYyeHe7VVGuMaWJ0EwMT60HmViEy9hKnt9uF/fK3VVuloHcrQ420FvGvW
ahiKWhG2nCGSJ7YptY6ogNDNFuoaSdU03vAPSF16pvuV9kHRQetX/WQRHukI2B3y5BqM42Zmk4GP
XHonrxcGhFHyG54uvgubL03E5+2i8TlkFMheqG/SCBnLlPmVelUXTQmw7ROW9cVyZ7bHMiAb/Fgl
4tcb/88DSj+FhG1YZ0spFHVPqnsFBUkCibShJdm15FZXEeWA/Vr7N0Pf53RW+QyVY9V9uVCb2w2z
ffeShEiTLg1j9NYbAQ2Y50wL72PsOaXwDF/jUT8TLAGIy4adZZQNfQO+ezSlcAstNry/ScuS2/Fe
gf6pVxZhZiB8/FVKwEsaf0EK2S7xfjD9uBvBBooxJJBgTH88nv+h1SU9EwhLGiNLrteuxfkC30qv
Cm0zNTMSuoCdPWD81nTNsTP0skhgRrM2leUHoHgA1fab1YnBQfBWzn3pnvW2+77qgujWEc8mjuLo
A4gm0Xe5mAgXFFD2kN9iKDdwz1XrnpnYSjuXi4MgkhUPTWv05n2dJqR8cgHd9wKs0B9Pzs0LXBxA
qPXnC1+4HZqsmB8KuXQ7LTIfNaWkwuB55xm9WcelSsxqIxh1qEJcvknqxdJLJB2pkZqNHcErA07T
K1EocF70mOw023p6l0eUDCB3E8uvogfOIUxY2FzjrrwP+FvzW2jed4vHNelNh04yVjxmDlTqR6UE
ynSrxj1gfx2gom+wdKgU9OvPs1/Qq079diKxVLyA+wnUHH0z2U1JQge5VfCGr4Um/BiRHS3u6YrL
Hilu9gbaEDuVUFMAORx48rbRNGFqyYzFOhbfJltq+MGJ2taiVO6XVI9Lvy9PLsq8Y6/teW5Ld2Xa
jm023c4cQOYfWrudP2U26LsAyqCZuWovJw+oVn9tE6e6C0G77MYe68aCoL3YCFnUOItR9JIy5jbY
WJ5aYbOkwL1P2P7Z6KG3sE9gIf/Cu2LlzoEfYwWLNf8QDHO47cyA0QgrtO5lD1ff/hBOTySM4xFV
gfS8NIB8lpR34LJHhWyxmNxS7LwMaqP4LYeEqJKnfHRrheQLPA73hsur0vMcw9X3DgTB25vGr8Dk
GPu2cMPouoOHGE83jg6ME4s2eL9yNLmyb6gTNiUkP283CaA169gHRq/hyCDj0EZAPknT6kLGkKGh
F3QEEhKr1Xu64H5jCEQxENq2b1g0xc6NP4Q5QyW/S3lNXBgvac0CuuPIZ5xi1OmPppI0d9DmHkZM
kvy8VfYCizva1NxDELPG1jNbPF8TPXS8f3lvEWiKVoA4WPIAldxJslxF9fEfOojwgYZxcwvgCVe1
y9qOntNbvtCLRTTVwrU0PUuTCFk5k6rHZ99E0Ca4WzODJu/imn5zUCGDjEf0zZ4GJ1ylDchRDi9H
fA3s/By0YnK8zoVrPsh0Tx9TkV9bB8U6vtQlIe8yFMV8OtOBSqmuUIf2m8JF2bYjHznIX3SyTrSx
LV3530HDMVNyZn8uLAnDnpkE22DDDNqD+aHMU+Z3GY9ddBx66ri3cXgkfFKZ8O+Yw+FemSQmNFuF
M8mDd6bC1wCGa4FlmXnH7TXko9NGdK1+JrMztEML0LNWlbhLdk/aNhWsFDaWY57tcc9qsnP94B+b
QGco85YxebqQ4vZrI3WLRR+lwt0SSN5sZ2Drwb8AG/HKFS8PV0bGhQL2+x2jsl2vyLXjmuf6mr+F
nKozIEH/vZ4AFetBmTV1ESggkqp2OeDbJUgitRcYmmjghY88xIigjQFDHY5wWi7Cm4YSbC28VWCL
4KNzbqOlf1rkKXAA90Sz3ms6dB9ovPkwjiIikv0VpUC/CuRoQk3asCNi0gmw+MDKFEP7natrWrTW
l6fvABYKFbKaJBRgzSSfT37u+pje82QdUwUMJqvozfzoNI/xbewHAdqJUI20elwvG0NMqT3Glr9c
3Mi2Ygk/j6RAmywmSzya/FPo4kEnsLYSKTxWdRCxBg2V2YL6RK8TXHSJTxCm9JK6sdiCsXZ0EO3R
8ok1lcYQQ6QFd4tMmuXZtb1w7dVNecYk+6yqrhIml8sRIJWFMDQhWLudRzbwT6qSKBYmGSl2Uldk
C7CD2cE01LzfsTlFs6PSJ0AyOTL0WzQEPoRpts3kaYjHHoE7F1/8y8UaoOn7w7pXLep2NYAYVpO1
qaUJCoYqQV51QW+MP83/bzB/84e4obLGFmoQAunJ4XEyV0iBKf+2PNoKeFUKmTG4qtUgzKm9mWmV
bNiHIA4QarQLBzgwAiWJrjOMBvXqQhsOhZHXBwREtkkT1NO2V94KEPlyXYxCDjEsYcTMcGOTwZLT
JcZs9m60etIiD0shCarP4rytOGxFEzLEsTYeRY1Ki4KfnAjFvf6SMRAr3pJYLFS4/rh90GTwq4OH
16APKFJAJDxg5ycwF2WSfpguHrXXv/C5Tu4fIjCST4wi4uQvMAjpWguoHbPnnOxeVJkf2qH2230E
QjBPLV+i0CoLBLH5ymB52WWyKkeUhNuHArnVWGcQw4HiWVczvxKEo3kgppFU4AGdnWHywq2eocTi
hVxdgN/puoSg0A5AjqjJg6fp9whi6/87OvG3NvNWyshQEapD3scdVIdezcpiwB+L2rxMdRsjaiCx
kHTnFeM4oQAYCHipMgOjUvYBH30MpjNVegjP3+tGfxX0YhFk5mEityVz/VKtPG8cv9O6se9EaFrW
vAgsK6Mt6HI1jhn9b8JbauKMmW5rbTFCZXJdXAai+/4P87cPTAkX0yG/RUIrBGZeF1QTZU5HYFWY
Lp25H+M6m6C8GFEPCk3+AP3mgc1iqrHhLxXEnQzhnD3AIHzkewRW2zpd2ZAFZIiVHuX0bLJA8xti
YOj9lRMa5lJ5AuZC9Gq0X9/h8EReh2BAxtz5YW2UG4tYF0H22RXYix/qT1bRBg3/3T4ey3nyCmcH
7OD/mLtY4YgFRJxkeRC8rmwTGRVaz4FTzmgW5uhzIx5uIbbIMzQ6WA7dDFu7u4GARmIwZnlom5mv
uYP6wsQn23BVtA3lSXzE1HyIgXOMigqLJSd+ZRbwOf9HhHEONMW1ZRWtZIfKcnpOaopO5v/yckES
0ZUki3ym72I8DxkORCbO/BTKBuzWFhrPNFmAiDdiVGRwh7DtAa5rr1JZT/uNmbxyQVKRpKlkz/yf
1J44/GPmyCYlAHPonA8AgDCqlNYKmER/ZXJP2vOQWDBxnFtCO2NecsxRULvsWzaRO7ErwfAIaLqx
O0mdgvNA6bCWDHNltiupY9kMHSP6gmD7UTG3xpa/9BxTmVeKtfvs446det/4LEQdYucqQhb6lVMD
cRGTJuqnaVjOUxnHLswTzo0L3Udo8PXZGlg0u43sICh8KzFMHxXV67y1Rc/SlUEFy4SKBPk+nYUt
AkoXIyG+oz68KUf12u/BEtEHh3qVgUqnamoYET35oP6LfNW6qU6+JlbJuHRn3URY9kHQ0xYLcgV6
uQkVsurR8EaONs5Ic+3k1oCJhQVHIzOgsAJJlEMZ+BwhmfeQGVPNxrEv3JlV8+DbGCiFyibN6G5P
j6WwZa5flzakrXxn+776CGptJdME0bm32Sl2Gh8mLyoTyLUdFj4Z3DmOR+IaCcdjNXruSzT0X/Nm
VBNv0he/83xyL0byxKBSMom3A51L9ySW5RI5MxqWxMeZYXLYu2B48X1OB5kxcrlCLThMgUN3jLlX
gVuTxYifOW6O1e82DLG/lbIo5YFmRHVygoYP3VUtoZYqhhzfs9yc0SXxWphNu/gGEfUsOGnRKWoB
RM6WpNcyo0Uvbq6mqNyz77X4Dq3jalsT/rU+sm/yDP0g4XfH6g87dqSwuMCJ3u+nB5nG3E+zs3xe
k6d9Ilg2pFTOAnBrN+Pkxy4x8F1w01RhMCxQbKzEI0p+tMZ+LmesfwZ/5eg68aJl1WWviMchfQZ5
FW297ADipIqRLlyQiICjw5xkqb5s2geaIVL/QPoq2bVdHR9WJZebH5mNfttzno+b9qBNPr9MifQx
7IdBOI2i+iuDZvgEmPNT/YqAUN31qWg8fNGhJET+jVIlFkWLF8nJh5fBuZb57LFsq4W7hXEBmGzX
3JwJ/YPlWYeLqubsXlYDclu3YdGVRSxSbBEVvZlK1JVE6mAun+ZYQKph8WzDVbBgeEut0sQd+RTe
v+n+m7d7jcVF9uDKx04CMjtDSB7xs9dtdpuz0LH3m0dbKzixojejBacDZV6iD4nI+3TS/L330TC+
nO+93r+3Z910KiAwuesPtfI3RcEFmszOXHxJ1z0mmb3Mx1SnmgtLYt5OzZbLEiTXkCcknqEBJs8d
Ks9zBgqotmJZfhYuQRPE+GBRdi+plFibovHVd1KuEIIC9c9OdYz+Esy8atcbFcVoshTJev4i4gQn
9TOXOgtsnyOJZ0o3sw4T7oYCsNTfd7nmpzGdEBReR6XeOsgS+oSjCrqvRcqBZ28ir/BEA+bPCbI4
GKxW/17HSn9KH1wi0or9Zr3uMgFamz56nr0ZKqT9OpSGWWOZxZYTKiOgIuw2lRm0mq9FXVo4BDVF
bb/Nvo50agoI9GyePktTAAS5V9r//I51T6LWduOpZnknkE75wODGXqyq+wlYSU3liwqWmEXDym0f
+011QIZYMO9WiKAjt0aKs2cdNGlvWIlJ3fLN3+K1o3gOfJizcw3GRobU8s8HCgw5Cm5H0RY1xS3+
e5Eg4zcDk4iP9ifxbnu8mEWZeVng0MiqwVv7Lmq7zyFp3l31D8QVHnwQIp5aYnHq5joW+eoZluu9
dQjWkOTVsunM1IlSgl7jzm2FJmVa11a2qS7Kbf8Y3AjqkAR8D4+T8V6yJx/ACOjBl67hXgblBQ8V
Bq46OTH8r5QsSlUQsO35Mhmct/ivjKjun0gHqlovqoY2UUzjuIJAoeesaGNZbKqqBcB8dGGhcCKN
bwN4iosPlfnII8WjujUs9ezamyxlrA8/eYyNybygrKTm1GxvUqL/2CKLAz92FMEgDd34C4paw9f4
9gcIa4w0U4vQ5/cZ+eFNPcyCgWOzQKJVnm000ozqDp48ELNAaTy9V2yfns43/wUZkqWDJGnfA5re
SOuP3OaK2kaPQU3jp4Q/xQBETpjpCEmRgx+Cws2aUle5lmaBdQpKDZIaJN9Wmhb5MnNytwVIPSw4
BuTHpMmNED8QjX/R8j1Km1g/5nPvoe2muN90siq5UuGTTZIrol539i0JYVH/VNWlSW5MMtTKGyvf
TQ3exHwFCpgcpfg7AmPEXhwxEQR1Ilgp547kiio+CubhHTlmmXmpji6Y/5ZzS1vzKG9OKxsKOtYD
UCPBuNitqBb+arhlQkA1pZG7ltYQkvbFZyu+1Qs21LsFFTOqdP8QsowK8pJmx1nqRxfNylvvT/Bz
5lKcW8L4abwjzI2rq0Mni2i74SlMU0kh9OIv/YkNCr0M3FE2qNukbhwHtSwPdl2PwzHXii9TIY6m
qk6yXxHqNH3B6l0HTlRFtdWJU0v+dt9OdMIkibSCJaHCiXSlACfcxmvJGnX7ChwPFdmXtmuorVjq
G8a8PPtoN5flX4cSSNsSInh/Csv6sp+JMMLjk/Ov079fU62ucPJu+ze3YTJqusxZ8sw6O1M2yBgI
UoCqZGC61aMyXgyNffzHmzJpOEK61hy+Sv/sqdqhanvKbzseM6VeytywbiS2CxE3LW4Y7R/OVi/y
JYIY0iFU+tAeCvdLqTv/SpmEzUhUUaVe/NLWAjrOOKHJ8PjLJw+N/aASkf+4Lzzi0yN2CSGCzc6O
gA2Gxl/Ti6humCVold/qbLS9Uxj3ap5DaC4jRLOSIX73dIejIW7DqQ94eedb3G+C0SzlEjn00B34
SsAIwaqSPmuDd/47iZvrw4TIHTj0L1ds9FaOa8DQEmDSmPkxPGfsyuL5hjU4eudt0Je9CLjXyvi7
yatZk6Q8bQgMGOqzzIev7/qm6TpnLxV+z1fBkegr2SkA4o1zKjvZcqqWuayJ2+ybU016VP8x5yyU
wc6y72ExwmfG7rDXczb3VfgTRNGOnwmtp8UdJH0dv/fm+GHXgz7yQfTvUs6g8Sv0aiF/TgSof1x3
kZ3sI55i2kqbReDCuWju4Wz4UShqh/p2zKd65EX3Z5wR34An+/XKybGWA30uhH+QcTU9l03Ny4nt
mQoA46U5v3/5WWfDj3YC9DXb6BznJg2B2kFagzf/kJQiZnm1gg/HHfhl78fdR+pLi65dvhV0scKA
iCkm7feOOq4tLKDhkIliVo58nmA7ncGdvlntNJunDpvbn1HQXmFbqBPhSX6GzOHlwmFWdMT/h72p
zICti9b7c3s/zgvfgkO0UAOyBJ5JR+ugZf66mAzTIqKG79oDaCsZH0LyNhpuCmVFUa/3S8eonhvX
9VTJ1NNoHtEee1iKVwi1fp07CtD1Tbe/ktgfk6hWw8eGO2ewtoK0u1nHoWliCt1/YOpbiUeMB1GM
ISBxiKeMws8pkw2cVvuEl8RoFRfzKhWYlWjAAwDNyq4Co55HK7SFoBAiJdatTyibgmEqxeLkA9m0
jY1CQyv9tsCeu5/3M+TsiP0i60zyKqLBKGuZsK4oV7IBLXpi7e3o+SYilh5iCxz4iVGCsu5Kw9WF
BxpEiCtkVbB9QsmvcIMo5VTJBzSRVvdWSyRKMzBjHfi+Hk456nDFncxFB+/36THB94NsLiwn2tX8
6ztPfy/Ij1Qc3RNprD2H/jdY8I7QsJoxdaaX9pTiv4PHEpuSOsYK7b7SfcbmOZADYE2/d/3YOKar
ZkEm/wkmN5dB80AFVEOT6YPxq0SyfMJdsa2c32JCBSPnXa3o+U5A0Pohj9/gc7OYJpNEoPM/SMAp
gjz6zuHFZZPZTr++J3o1uQzwmVojDacZRaz7qWfuGaVaClHmaS9RyeyE1Dy4wWqCIxwfSndvS+B+
d8uPMcF/Ki4zhYg82lxl6DMLaZiJaQN7p2arHB03GtgKBRkpSBMbECPylpRUl2yrD4mGbCj7bW4M
FF5INyDhlUgfOG+aNRC25WzlkhJzESrdUFB0xaP/1UI74r90ZxDjj7B+DiNtmfAsZPfRBkIEwIWH
Bjta3q1Qp27ymwQRuaTM/BgFrmOkx2lKXZCqMWTipeuCMJI7hp29C6zd2Ef6q7OELmmmUGDh52JN
IjfUGBC9Cwx23HY+NBrnwY88yK3sjzZn7+jlneguI8BdBLgRwp7tDryRt8HsIkpb1dVHuxwJpCus
9Q/HLHmHwv/mRvvSPM0mQzjEi0R+ZglKZ7KmqSVZKpMIScz8RzfHsZFZDX4/8Gh1o60osNrSvz1/
R6kbs8eTOOt7L8iIYIVwcl7faAkms3YlXbOboDZK4EMk8g4sHNQINDNLsqqhODRl7H3yzjtYOrmJ
d/9HuNG/+qv9hPpW8RyEAgte6JIXh6FQNB7Sl42utNLtG6x0ee7QreNWgf6FyPMH2tFmrZQ9Efii
8+M8lJtxJRQvnEw+9fL7Z8sCisLk046wAAZcrgcYjn3Es6lWblqwB/qig2r5U4izO1C6GH7K/DYt
7T7KDdv6BaUVbmbv+MTBYZ1Bq5natVXistULLe8DdwVao8+aVzBMzknCi7d43LclVkI1HhDGMct1
IJ6WM3+mZuo25WaSiv4zjX4+dDwmkM298PHOPrJEriovgaHbI3WeURMovtPZVFz2PYgBYyW8G5XV
+UsRDEc4EtFItDpTTctJ6Gqp1ysrHDOMws8FsYhsTeNtZDCcFsjLyE8EMMr2U65SWNkum+25gQWh
wa1qY2PZUfa5rPhf5BpiWdAaV704meu862b8iI+PlfMZR5hEC+dmtvhmfTY9ke2RhyImoqYCrfmy
wGGMS/AgRjCPRJdGMwu08ADZwtPlu2S9rSE7fF3i2l58lFeB0lojF+zIsfstw1UBwF879TYL/Hqf
ZSsslsZ020OXTXODd/vIUa+Gs4HIr83fJ8m6lqT8it8wzo419HOFAigZsLZiBqJPOHwggJTfJZZV
aCDoeOc2PGdfHI/IdVKP26l384kpzjbLkR3020NzD57NVizFrYdLoNz1p6HZ/ZyPrP00GASsKZrZ
1D6XzjUjN42MFG2XxIQ2Ism7yykBvKgpVRQ+fJZM9LvT1AxZBshm3mp5OI85AjvN1yx0KeDuVERI
gMhw/UzepksJX0fxJET1Ha8Abw/UzZm33wR2vMiUlsOjp9zjUExQ9pyPEbjj1aSfmah1YrWkNCAh
wPS/SfpJJ9XCpCleL4dZzy7zQFT8Zf77+cJ8aYPzy6eNeAGzT5K1UrxL38VSGaKvyA45uoTAH9dU
8tZZn35lAasJpwvKNntlk5egm2aPhDUultS5siPXWObYL/FZfK8jkZW0jbYQxDYlhKtikfzHDIzg
IoKPdRMW/1iTCmStn472zoqVzxCKNAJVAUu6jsKqgaBa28DEqECi4V2I3VHhaF7Dwr61GfW987hH
bpjv4XcnXVbsPiwYN5W83903qzgS+Ihs679+E+vkHqc1mOK4+A1tFnMvU8aeWFKw8ddzgmnMGnQ1
iMkPk0ObZHKLUu/NyLAZ6EKN5uqDsvL6AOBRCtSU5QIZDvM7Cts3Vz+mm8ITTwamUCwT0XDR2LAG
2y0JREDj47fJj/uzAgV+uxEDN3q5NgxuO3VcvA5XilUYarNO8vn367KMXeP3eHQGJBMO7DUb8+OB
Z4DiwXuEbXw62kROw9F232AJoIh/QSn59orKT65NKYu9CSijElOzgTocE5p2ELXY2X1nGPEdWDhx
kJcWVoeTXcur2Ans13MyN/aNzxsToqc8JfQn0E80mSk/Op9j0t2rWt9+YBllTAM52cTXc3i181b+
azml4purWDO4EN10hUCnhJD9K7h1X4hFX2/o3wj/fclztdhR72LtNFdDsUqV4eyfCP8TJSx8MZNJ
1DBLzPrV1rR0iUuAJ4465uwxv26Dh2ksbmHANTufvbfVSBX1lIxWCJ+KKUOlntKjTdOgSUrNGZm3
S6d+VprVB+9VzSDXkkFDRB4JmWRuCVLqFYS8U9r1c01drR8IWemxwlVtkaWARRa/5P/mTeHG7hIE
KJzDcUuTu+llq1RhhPPhzYjW7RwN4fs6FhVR8sdFwnxMzPOi+GYLNO7tH9NONJGRhgEOLjwcwYCj
2xleSY/IKZUW+rYjkPk9jzMsxmUWKcufQ1fJDdSvlvcKpKM6DoXztwBiz9rStv1Z/N95eeHJjT+s
OIaR6bZEDI0BiJEO9WnBjnsOOQfdA4JLs5Kmi5tfQsCv9rpndnsB3ejv/VrRBOM5nKQGRao9oCNy
XMs9ShTB1ouT3MhwaTvz1hEKXhXDQqvRSgYx77TgrKq25gK3hpCK4nVqHpgzn9eKAnpqbN4Xj2ZC
jJ14wQScGAlrGtnMle/tcnMXSOinfxoLg6/n6du2Iis4XnFe4u6LTWW6XBan3ju4dBeAnAikBV5z
LhGB7fwj/1ZXBOv0XwrGAb5tee2CBqcC9Xk7EeRoClpgH2GBf5aheEikCvmW5zQa7lMasKETcWa7
r5CmDI9YsjS3jCuSBPhDrTpQg0gi3j8TTp1DBE/Qrxg7+8OntAcFhU67yBr1l82DMF+3m96RHV34
s5uWx23ZeIu+U55XAkohDOQCFfASPe1T4znPK8yCpMcKHWnijn8MoOxNqJh0E0UTzuIoM6vDiAfg
84vbL//yt7g6UoqcVixw0bezEGTtEvuWOwJQ2IbzTWO6MJg5DdGigSdSfmqmqDLVW+bL7rPCpMDl
UONPpDRCG/zYNYypNqFylgz78G5juH+1gJ5PKn/uENyscAxjTopP7K3kVgN6h3f6Lqcm2JCRXUv9
yC/jjzji13OScRard4p39KtAhpd8kcgVyVf5Vp9mzKquFuxSvGM9vk8aGFNVumArNikNvo5UmP6+
k0L3eK/Cfv14CalzuuI8iFQo5/3I94Lsao85kM/9XR/dAuLnhFxOyg5mg5oGDigKYNJegxFRbFqc
Pz9AUqtDzQR+C+NznKQhbMQLPrspjFqrRSsPgdm5VmwM9wNaH+Nwh/pS+q1q4HY1x86jqFu6iJJs
6C98+pG/M5JcGGbT2UJwRDW2x8wLxKe9jyf4qoV//tduklb6I7PYkil22H0IjKtFvsm4YuYxFWX+
dHMX8rZHQUT/rtchspSk9Uoe+zbpLQ26RRToxjNdumn6+cgkBmMYUNePQ/pUBJr5pEnfuI0rHB+m
CXWwX0OJTRFn303UNUOS1V2QF9KNTckdJGAaS9cKJvXDVyJtkAb32Bc9wQK1LTFWfC8DvwakyYub
SafIygo2GJDb7srlk+Np5n9E3UZChPOpD7wQ83EiwSdwaaoWtUKsNM01bruBR/x5pNuhRkzS+Bx8
aoYazCzbg8K9SU1bsZKFkkV0CTlT2B6bkhaQEOA1bhInRnguur5H9fGTzoXtk8RbNnfcMc7baSmc
oTIpzdkzATXuTr8xF4iV6UhZeyryie7FSSsrJLXkTT/rAwdgI8AxE2PsgCkHp1Ow5s4x5UNBxQu0
s6L8IN9ybq8QPIGoE7khp3TE7Ss1OPWVpStm8t9T0POKJejNxMFhfIKa5zzgCJQ4pob7zU5I63RC
SPEpSduCxo4MpHEK8BQwrS5nPgshJLomGvkm5VrwyzWqLt+Zncx8b4kXkj8d6WWNBkAGhr/JN5WJ
hL/uZS5xd93E5Lv8XL6JKNCvIwGwC7qWiS8GXzt1NilIoSQX2HnuZDXPc33KKLu1fHrKkv2jxKTp
7a0f3IKl/8RpTXwyYl7KqLe4rzFVXuEYKA9LV+oRmmTRtvu0LSj+3/QzEyNkFxOlzsJJ+lwhYxvN
KZP6tSzxbO1yoOURjqtW1wYG2ohT6pR+vHybZJeKOsdBF3Y+7TWew1OChlP9hQt7X2+JwYZTFfk8
xvl8/S+UZN4lcCne9oVqgrHXhGQKujWAQ190n39Q0cFOWI1V15Ky8sD9a3x1r5O5AOWWUfGscqUM
jbudoLtaXLKDw1zg18KUQFetKvSvFsjpXagCD3Sg753+3zwJreIdnTaNrM/rDbjEXapEE2WHMVVD
opux1DY5ns7rcLihH6gSNGBOUz1BiYgkOO2PuvFBD1VymkARh6+dpcxsMqfVfMoY1VRFYl+trV00
6tprKdXlLkYv8r/Mo3w3HXG/41Cz/ZUa0O/Kcsz0tWlmQEvGZ43ID+/4V3CRC31o0anD48qoOa6H
+7j8IGt79pqIh+VQEJOHgwX47JjclimRBoTmA0piB6XH2G2VVWrvX4xpBEe19pW6JRF5zlJkdQFw
9QGohmBd5Axfra8S3GQhIA+01CNAO1dhfT0qivksaFcnnshcxAV40KqAdMiuJrBu0OmfYEJ6P4n9
GmUQVPsgGipdZDEJ7JojWN+U6KEu+sEC51KXrothl+mLPGQCPessse4E+b3qqcuERE9k3X2NvGMv
ExqHsl3kiwS7oJ091UkOF91bsUKVJD7Py5GEbvp7tRFZHTBbhT+3YPAqHBvZ85k8tFRL6VNudOrU
0+orKt5yj9X0NWavQMl70gIMIDyROZ/YsrtCcXn5z9A7SSl0RdgEnH7LGkosEB8Us1CfdItRanfo
KxgP0gm2Qkj5JrEzwOiGJHEhl4a66HBgVC/wgu4s9c8uJjPllwhrziO6kVdKgVFTtYqO+kGIXLAk
eNnwrEn0NVArAHs/po7Ezls4t3i1SO7R7+xsyL+7jnpNdG6mArs5QfQLculESVjtvzbrHDwJE4jx
vXyHAVNCODhuZZ4bCwLu2cAXqUogA4JJvU+oEP3s77JrlMfBfTmSCSl5vGG1L0md1oImCjLJCWop
y62dnjmXcH9cm/OMiSdRiMUWaUY93UQ6jrOsZfuTNtJLkHWZXLLjCk8f0gPAxHGOjknoTI5JXv68
X7/22RnoN7vvTLFRBthpPypDhtMLdtzEBS3Q0f9ize0ibPOXTnvxnACSgP5ULj7KzGPnV+uyM7YA
3GjJPPI4UVZdv3yzCaVP1l2lH3lRpFd+QTc1g9zzBt29XZvbc3in4pVbetJdxQHwnph65nuM64jd
2RXlMMMj+6rBUwHfIsEtWwViCZ5hvbHmnLqHo81d6ZF2/b1AgdsizCThFdpWKBd9mmQDOJlk+SAP
T66mS6jd5hO5Ee+7MkAKE9R/ASpSa6p/XbgoVQ5YripA3i1VUmhM9y3JBu/nxpIwPxzTPMeHYBYu
1mxfcIIldK7+jpFKNA5uTSbV3VkWi3VpEU/0ANIbnuYwif6w0mRrUjbiJi8N9FFpm/g/uC4B2TCv
UxgB83/v4rvI7GHyICj8b/jFZ0stY26wuFj9Xv2ddp8j5AKe5FoRvXULNcj6kXVQEDZ/Ri2nnukA
Vk7DArwHylvKDFYCG/XFFAjedqm9bXf3fxdgCrnuXVRe5CyjXX/HLBhJC+sI9qJ2RG8P3oiN5ZGo
v7q5xJfwqY2+f9o1EAy5Yi46oRnCKdEmwgavKhSj/cYYnZ4Hu+iTJ/4URoNUE1ZEAsSZifNL0RNM
8eAhyG8BaxCtWOPoyvjFAl5MS+tJUFgYVFTxKki13HYO6b5YAQangFcup4FC1B2gtv0p42pmpMqi
BiReIg24jqOc8o5G83GSXvQokg1uJegFTrGmF/XA+ngWhuTOZfNWs/lmbc324jEgxFi+p4gqGJSX
fEgv9sVP8CaEwlLvXagb2It6i0/UzjQpg9rQ24wzPbFvpIVFdsAn/yf3ToZZqve3QON5tyn2uCa4
y2rI1jHTtEL5zJdoqmpII84aKTJwhZDTQN5x1e1z8O0PY0o3YM/QAsfnmlwFXG5oDirpv45xgMS4
Sehse69BYpRplh/7xC25kinm9pr+zjClItD4BQHoX5peXelz9itlwYJGoOIGAV0WIrQz3kVst51g
CZCxH6PhFGpHwJVHLPPNUaz76RTtOKXeVFw6/GYe3jD0VUxCxF7QTcY2wtLVCeo4uJ/hMB2atE5d
aqqiimgyqZx9fbCRxtiqShSjujdBXzv/YHjdWfP23rPtceSIzdJeaTn/fD3OgZLB8B4t1kjsWGsr
GD5oLGkUEt0XA0IOMbYJ3NaHKI1nGu62yrMdVw8K3IBryOmGNF4YC3eavWz8NQpin8XFgmroEC/b
5uFfdD/O3PjgQBF/Moqel9mhfAEeXXj/DsK7dHG058ZtaqmvwYT+yuZMs7zKi/Li6TMFLvQP8RYb
cojCqV9bQg1JKwB7cz3FbpFIZ+D+mh7ppJLHXBvuuxi2PpwUKXznBqjBMzWPvKJYkZvv0QlnaRfl
HTrZKIC0yNsNILekSk8NHSJ63dbGB3l5TpDx2fUigCKdlvEx3OPM13W/8lrdBxCL1SplcrsfSSy2
TMy8qEc0Thpvour0R4R9w4IwlSdgl9wqjB9M0Hu9bogmrmPkz/w6inCcnqCK2Bp5VokoMfGBB58W
z75KXeqdITNRQu9WX1klHyvwgOCsRPQSsyI1sJmVx5a3DY9yicFlxtBBud5c+zbripXhS8u85c6O
mTKJsv/0RwuJe/kC/SFba7fnEmEFE3JG5qA6LBzcT/+zB6ZzTTuY7eFOfIid+IX9EImJe1PAAHG0
lB2hMYf6kEzxAAb2UqhnAHDk8/YgyqOIAcBXCtknWZUTO6I32h4gNzGoqC+nT4Gtm+93yx/DDlBX
oBNsufVl4wBA0H3+ESC7RYUzMf2in56EvY7uwjXIdKeq0g5OsnIsu0z2f4VbH1Be4VB5bWtcRHxk
QKU7bkcub61uKkEcPfmHl48NN96JVUtVMaB/5zOp5+kyVeRWCJrI/+Z215t7yM7NMy4o8d+LeU5a
5+uMRxF/oitNsX5rBKImgmSss43bbaTdmr7+ACl/f/5KSovkCFiUvW3u0BD6SNZqxB+4Hbs9kFiO
A0Mw75sjaOyOeKS6CyUGOxIJPC/btxuPO4NsiY4AbzJLE6ANQXg2I/aIxtfBCPI/spEdD7fCwnjY
6NtIvmxr3IYpmh4eR8HWWDlW2GHx8BtE/luXMW/YCKCgB1oADSNQQb5ji8X3cYMdmvGKxCGTQs06
EEuO4cK0PF6hv4TyDRVbUFRLNVom4dZwq7wRithLXDFnz3nRYPnL2SrTR/go68gKA62BbFzZrvtY
xxV2GhbNYEUCt7szXQh6RovMuZ/7r5+lBkYyHepc3XutiYjTW1C2FfA2UzHGIAZCZut2O4M/ft0F
IU7jDs2yPaJBjF9k4ICZJcbTp0YuXOYiD4iJDFZE8MDpCLRAw51YkQT6XfWtzNBkFkgtBnYiE8gz
32AMSvcLchymqrQNPlOH9PscOf8fQ6LZ8Bur1o2k3EtoGssKkfeea865QSLqcLYH3x6CnR1I/nnY
wpkHfEOZasDgjbQGb7HYcn2d+DVi6Ryl2lT8r1nhCtBEpRELnHtc+eoPpjT3wfJt9veIpWLZzh71
z/wuV4SMLW71vYvesfdAAqzOEL9VU7IlvxgI3wLQRPtRdc466IE5F1be/vwEdZe9KJvN3uX/7pDt
S9J3AiRLAc8W9l2aajrsmScBQ11/AFQBEn8ajI2hC+lg3OyK0ar9bqtTUD+PVupdpXc00X0YSDlC
Q7I+5FgXSwLfzFRjrb4SDevHP0i6aMEcw8AUx0AOi89vPzaCq5pY9QI1BiS3Kap7dSmbMQKoL3KC
aEi13MuFsLe7gPHWjia/JAURi05mo93p/1hY3qzolHIADZM8ELJSfsCRTwBhnYfFLa7lXooBJv8G
qYzJAhvwT76KIf8tOOcWkAVqj+3n5lqTZzPp9m0O8L5HvnA2a8/qNqqTUTJhddMP9V134GzndFyx
kUJ/I7LPWzOVsTHwu7AhgIbCb9HqVZsKEo1iYRVMam/P7FoimNS0cbxpAmqjoQ3Tgh9wCWCE6Bkf
4IGoOslQbIbqSB5v6qCQLaGNL4nyDyKQ45cH8qxE04diKNTADhf142+66wpnq1HFBRS0xzC8mO6j
GJfqUFEgh/Mu5YjbcBfek1dO8CQArviZQ8Qy+2yc88RixjTR8TTBj6nTKXLHGclORkgqwMkV6XHd
0uipkaIJ/FtdCAHfxOxBZHlEYric1LX1THvEn4odADXOynqaQs1QSqV3BxaDJdbU8uFQ43CFp2n2
6TzAJqxxXcpk/YID34PftfWblM3mPMCQL7vrrGOm/b496KlqpxkyTi7CcySdZAk7XLVbiDIJrw26
OeZOWFHi2PR4TbFD8Vl4SKgVJZqwBwMizs/aM+zYhh7COuHhQiYlh2fCKfNyJsSEGe6GgTOWYti1
Iy20VPILg4iinwGQpMqpMYtN5oqYIgqH7Km///EM6DJvqvx4paH93H9dENgC+G4qhtVp0qW7tfuU
BsZ+Bpc4uiEp3H6SJdlj6aazL2IiAjOd/alOXqWyFWHF0LQ6q5MxL7FVV6BpaykadawVF3a/tv3Y
YofcWAMD1MQsfD61C+DaAB8Qjache8koTHGcKKFPYyuGbWQmO3UFpmf8juzGrnlcVoHHYqqZe+pj
jpZvjzUHlTAMkSjMj1/3mnsOuX6h0qUVCP1synjke5J6G1GvmbbhZ6vYghLw0awId/ScBCdn4EQS
7urReWM+9oGWb6J8PO+kRMwmujxQceHxKPsPuO50odgHI6LArrFM5VGS1PkL5dITGRcPQb+dLImJ
AYb0TX0IouLcy3HFa5MeN/fRpRd39Wykq5iHQutHfXTBtaf/uE02R1+I1loNrM2EPm5IlrxMnYQ8
/Z4DLHhkDjzN01NmVDzDIZ1TWbiSNaruCZ9vUDIMyb7N11MyQqaE5r26UguF/9eBh4OOUhNAMEZB
Vod3fXnlGvySevexSn7gVu4CZBAAXO3qScJFAuOc4bOOv6cCz2bTj9vGvK6iDRbnDpJum78CwqRZ
CmAu8kmdRHXPr8lWmQz1AdliiJYP/LxLvzXK9fAZjfb+OPGkry1T0aeppslNeCyhgAOv0XGr9uXg
aDnKIvMvyaotxAshufOvQ/6TlV3gVBKvEWVV5z4iJRctMGRNI3rRL5ijvv2bnG1iFq9K1uv3g2t1
cmzOpKlRgSG7S0WraoTl7AEa1yOUELZzPTFGinkHxyC0AyvWMMkB7UrfHKlQK4/jGFlhanvOqZ5I
ydXj4c412xjwGOo3F9CMZDvFD6+QNjqmsd6qfcWiCzCioQmdA6zRs+ucycF64vgalkK8vJywajzz
wsEZjR35WnWLgYJSu6lImfJVSWZDZb2zK6sQjBlcYhLSwOvcrK86C5KcNAiK01mnRGLsIpw/zkxl
jbH5rh6ob0lelgOjjHMfGxaly9iCc8wTX9mTCVH8CSnmFAKgQKyzvG2hzhHe8cJ86sl0+UftWPRH
gRVGn10PvGAcG/OHq/pA26xqTQm2Rse4RNwdfDu37qbq2HBJBFp59bFwB8sZNKbLwNyPNwlJmvAt
rYmOZsjWDzCxFXFUVWqeIWwkFbs5a5sbkg0ZaDXkGk/7dYpTtObzQLJMedk8mD+qf+fhqpuddUI2
mmJPPURZMsQIno7vZA9FYPz6+TaGlOIQz7l+gPJ8zOQP6cp26ZcP1QZnUb6yvfJ7KsL3fVpxoRJN
fBtf8XfTdU06gBRlqpx55DQTBGuxDmF/AxbQhNW512vYdOa+zlzkWePEC3YUTGURz2Oe9vl/gIUs
4H+Hb4FL/2RcaWyPbrLruLmLI329MOFOSBJi0shfcDYG5pLkQGeRYIID7IKqRNPf07HawCUPuhBW
R2a4PYnZtUWCfPe4TAojf2XpOYvQDjRxrkM8aCNxVW44dDSlBEVuK9/7OqRliJMpzUzP4b8g2HeM
AT7j7DqUpYrIUt3+6wKMHxwG6stLwFdPv8KT52hUrRke85UNKtVsHNEDdcB6hYnYensW+UefownR
T4rh4ij24O3UZwvXwsHDMQfDZprAoayn1ppM8aTaYtY5NpoLHb8NBBYR++q7K7I+vEetatXnZDbq
ZtpJz2WhoeIxgj7nQrVHORXbPOpHbrCXmk0L6VUIJCpimDaKvd8DtzXaHNWy5Xx6a3OxbpZA+rAs
/avBQa767QKDRWtEM1mFVu9jf7YbqO8cbN0zRjpbGPbXLUW6D6BI443CasvUjALxxU0N2IaJ8hXw
76CWtS5Nb28X25zZY3J6kExOBI66lfm1vwsoWZMVjZifySRmv5jir0bloBpU0ebdvDg+M8x8Qa0S
qvfam1I+EjiC9VOoPKGznprSeJHvV9rswHwyUiHMQSfFWbGOAP9sgyC3B0oF6hSYJ8hBms0bqTWT
vwbqu3mwfDzNdMpyARIyqBuZ/GSM2zHQ8VWupixsyq2aPA8Ugma+1mnNnkiKS94Kn+q0GdW7z6Dc
PjwE4Pf78Bo2xp/bEAOsZyYeAcYSrlaCNMQ5cYBvKPWYpsXG0CclK7StgBDGk66wIAWQvmnI3/SG
5/XRW9ma8a906QvE5GaEfv5TA7CpLYDH0AkNsHaZTp7fye/wkFSTpLDmN/mT4uNyy2e1oLH4gi7X
qQH0NZ7sVlGOW0rSmpm7W+l7/Qa5LKKwlc5KU3g8j4DYSCGCoMCFbaBk0zjdhSA+LN6Ds6n1EKg/
PI0eYEDkfikj/m/k9h7lHaj7LK6DEnyY5wuohvceTqYkf7mRFryG6jcvgN4xiHHhxFaIRGBfdEfJ
NX/6D3fjBpcBNFJjMuRCmDRQ6G/L7avygm/0QxuUWZKBAzATmHihBbocn7oNGk+8XkfS6K4Qbw+E
3YwE/q6N8d/gJF69dd1AiLDTbtfYE6vNF2P/Mj9fhu60zE+2GSmzv8Lm1N0fuwdP+tYwuUvvj4rc
biT5aMaVa9RTtmVMOBPQJYXeXi9Ww8oNj/FcM38MXIShBS7Yu+UzmumFFKIEaMvzfJZ6hv9E9XUi
VJnBUVgrDOZnqziJnMEecJdC7iKWUso6CNK2R1RXSJyyNyKTDc24A3svV6f7tpCNeI5A6euQhKyO
5r1hwmQTJlQCGwvKd4KS+40Q6HmoQVwGw73rLsXCkhmFdH2W2tLos6N4xiHuvQ/fVbhBVGPWrk2y
Q/Swv+KH7waOHqfOTTebj+PpweaTdQyCeduSDZ0j7c1AVbFaMXAx0eB4V/DxFkS6c+tl9NXhta2j
5Fvzjl7gIK7Svg9EuX+AbVpU1bLnTmA3ou7QQ4Pip3SXBAqZkD9Q7DwffvREuOF/N6OWdBQGGQZG
JK0Js9cdGCLvPOAN+bTOQJq4A8zlIouyPPrs8LpNCOy432HwUfJ9qq3TtyW+r5Y/3K6/trvYuczC
rVgirHvmTJ6lkZL5NoooOG7aJOjLk+MyzzQ0K2PhCceqF7m2UeZRgybFmLnLusxdnHZ0YWuvU97C
vyQpeEMdDBvVNctLQaQXVcP5ef10BYzhaXs/dwjerZODjcJcz3mk5tp0L2xoKT19Af2fpuuVhuST
Hk97ON/F8dLTue/HxXRdnkmxVOn78SLCNTBIfmaTNmgf4Li2PrtlsgIUxKR84/eLKMPvC9FxeTVe
JxZ/V3DWCUEOQsahqOuBpk7x3DaJ2UatXdRNUmMiHgmRp4BnNTv5fgQgfQiFcct2TBC5eiOra1sc
tRpz2B5qGhrE8YZzgiUJuEDaOo99mB6J7N0kfZB2eSs1zenmrYxdJTrlIHftNLqLV9i1BrLt8cr0
Gq985Nl4Wm9rOw9ljNk2ME8Df/0B8nvUF9lMjp+MJgcur9gk8pP+h55Uzi1dO4TSP2tqgddowvbb
OZaGCJ11zvHGkeIxrFqvGPMO7CIRpu39cjYxbNZUwpSk0/MyOQIhJaZMIQDLMPT/l3Gj3qNbQqB9
X4rAtOwOS2tXcA8svzauUaJWt/Gie87ZHJSNdSzUeT8SwwEIEojqRgDYqJ+IiWE7pEGuOhaJWMil
eWS6KnY+f3tkKzv/yAvgzeIIvDQC2ZuP7LjgvvFhCvVa8T2cpbGxMUBm8AMQGBUziNkIxfLdhGA8
Po7199Rx86tM9eM3sR8uqLa23OCzop6J1FcLyfxPeuDl34ECkeF5emmOUPOVOdv3Cuyy3LCVI++3
21KmSapLNaDroXV6Ae8cOU3yIuV7W9C+L+aWMD+5+T+WQYI7t3oh2upyeD/IbxJ6FgjhANgnbmEV
XeXuufDlaXufML7OuIIrLzxz9rxImlM3LWmcQdn2hxPkJjHrERCVcQnxFXOTlmgLavUNVMGKUG/a
UFezO+eCZq/fWU+4XqfZvpg7GaXaz/rs05pVNr35xUb71CCL5tgBVbHCTtWojdYFjEDT1JjzB1kt
yOHsr16Y8maIqk9hhboGw9bPgzmjz4nN+qjKlzhblYZkqmsRfC8xKvu503nO57/KwmFHQ7uhsTG5
7sIdlsdx6l+9qP/AsXzSmCESxoIoIL79dwYvFLkEJs9Qmbu8CVtM9HmLXaoD4eE322kJmmA+kLlV
2nslFx9TjJAPifnhequZGI6BOh4yYAuoNubk7Nto/8pEtk+gPDkVfeDTbP7vXrqTW9dlM3VeLXCe
Ai9stbbOzacNqHyD+anLK4N7Pk2jeMHxcB0RFkQQ4DuD3RTEcL3NOQKFEO5IMU1RZIXf4Nd3E1Y7
Lz0yveEgSJFF0PMt2S1J1usTGLZEB+x6L0+CMpxCub9atXCUKmiMHdrJU1bjkanHkt4IMJ3nk1Md
2TAWkr9/s71utyInbHhJPbhHSP/U7jYprTCgqwTIy7tOKk8MXx5dt4duPr1UsfBBgLOcD20utIYS
IM8rdyxEurAJriJ0m280kKosunzNcezT+Wz+3WTsc+Lk5HVJydpdrclrSqzG6VZLyS2MZrHLXXky
BSe3s2pfcXLIIkL/bqGU40YQREvzCjHihW1Sl5USgp3Ro3LnTFnPYl4/3rsXL5YEMJVibtJoTSvf
eNalP2aTV/WnTXW4vI7aL10RbQZzkAP3zHZx9MiO5QNBIg0p3yLmluN15btovAwWNR66RrlgbIoI
MnbzT3AkF8lshVnO4VvFf+fgxwiugyoEFTFHGxXb0n4zYxY21+3RKSZpR2cRDT3dm7CLk21uYzqm
kcupUYk+GxEeJnQVEcvlDiJmXbBECcb5PekLpxgHLE6sGAsIUfyg1L0qdVAeKt5X68nV24YPSaAW
D9aifxjztNpei/oTgUBQpj5/S4xuhSli5OBCMofV/EYM8bnRzR3gtjL+PAF9MZ+c9w7q7P8oNv+Y
nLDvZoocjshuA1Z36F3VTkMDE8QVb8Aorf5BQZfguo0RLu6A3t46//MirSaKGhlCox/0IgmwOusn
p1NQF67q96ouVH63SexoVew3tO/iVdbIYRGY02nBZ8FwoRtg05BMW5h7isNI5BCs2RZdmxISCVH/
Bs5+ZEgXRnJLc7Eawqw1VoIAFwwQj/wM5ZIy/8/hfhEpXmv43RG7QSDdj2ym5+WQqZ14yPhWA20R
LeozHpf+bdmU/bF9XfVvV4lf9ShzlQbzIKuvSadGqky1dYtkZRfOp+rdN13BJdOhzEh137ljWG3Y
5S6w+oFJtEWQ5DFpgmdTaZS5fnki6IQh4LOs49Y5MUOJOEd5krND3KfowOVWr2rhK1VTw4P8pYSX
7aKPj9h5aSr1jyRp/YzNBcqzVc/Twgc3ATFmhg/3vjG4nsmn/+Zq/7Rb1i5BfNg0gNb5piUZWqCL
mb6MjHxVJr9Tu5W6LTMc/0c5R47KwW7zs+rCVm5Q4XmWOaAlKKh7JjzkwG9mgwjLuAK50dwu3vY+
6oaeOa7+JSZqCGS6aDzWOilvm7VRQNd36RzjvheC3Y7vVnk1Dl28UmXAFpFrfKVznek16Fpx4oAK
3Gln5EyRKYAYxGAMpqEsOptswHm3C5rX1eLU8wJvmIbLczH3SxjqiUza925/z1fl0TL5YgF1yw1j
yD4KiPDoKQkBw/X+3B0bw6ytNAN+2tvSd4tkrI6kKCU3IiupCGmNVpB/ML4iylAWnUwLKxcRrybv
mLmmLqOrmrwvOXO9Qku0TtJp/vQQ9eiQ3zyN1uGl/bLjCL0eLeZZj+dkq1UZzG+cBcLf2hM/uxSm
2HB7bzMEuCIeRV5cebSI+McXPZkwaDoMeeQqyAh9reT4jOJ9JwRF259tUNSfrxoWI0zDGx19cB/y
e9nEScYxMay+us60sHJvj50qLXxuVLqmbVF+FVSKRtlj+Z5wqtuEBX1LazZkIYQoPcCjl5OHlTWN
/6ryHsPqV5FOYoKXpNGCThJCfjVv+zyj6/PSS19dWMJVgdOeC9oV3oRHxP5gAb+Nn/ksysaLtrCW
ArXveHGvvPgjH9JOcIInHTFPPBnoxVDiWHSHA9r97itQcD19N+5hQw+kGHF552MFPgbygc/plqKa
UxfcI06gElLUYzOt3tI/Ew+5XIqLNitkOFDvEFWt0jQzq1mz3cNHJhfR67fRQ63pMGNQUOmS7rwM
UMJssrjrU8W3jCSRqOQYutlbeqrwGVM+LP3NntjqSsZA48XZOXeUaKg5IRbRyiZ6+1gSnpMOtEDS
8pbACb7yYI894lSfeivFFp4LAoVFUslP1Amp8+NSAb007elJOZPNDCm9O9RuF7ef4sWViDOqlVaE
q7H8X+r7YtzDRHCX3v0iruTEMxyEiWQOJKc94Pr20Dg6OOGyttnH1bhdlF84yyw5qSuiOtbfc+Ai
cQVMgmRD7hMWZHhQ10sILcUsc7iWTgJofT2Uc8dFvmyN9OBi7BWyT3uBQYm5KMgcvjcjCglNjqe9
tLELOBWc6zwRY+DcSv6hAgtN09kbKMmQqjN55A68k95mf7Pg90c/LLW/7WaQh1c7SnW8KpldGjHr
8eLe5IolkaG/Df9nXXwUGH2QkiK+UcsSCwQ3xPRgaFRIVDchLnOHz/3Q0WRZ5QuCYa5xj/tI3fNv
ZM1gjCRSaTogGkYKQxK/EBy0VwDklmnXYacX31X4YKgcHVEzb0A+LzpiNd+HZZn6stuFna3+FoGn
2Na7JOmrGb4zbNo385RWmxwB1uK7WwtdkLxm1Wn6j3Ajn6ATDGDR90xgjvI22mBqtC4GGnBgkfCw
UkwUeQOYO0+177JYS22omhZFL3f+Vn9reYTnhiNwo+MHdxc6W7bqPUpOuBQRDfv6WtO7I2WooapM
VN14uxjh6MhPpSptk9mvogIlEAZLkHtPYSiZLg27/rydeO1y78qjF4kgAL23fjzrEzsyVlIFvOcD
4t+Eh7FocG3OfqQjd+bbPG0U2tLe4LJRNLHn00v3dWrQsQPDP517OXKotJM/+vhFivGihzDoQ2f/
ZDwOkgqbqOx93Ovd3JRByvCZQ/rbCHdlDBbpISZ+mV8LGcxUdW6hhEs84WonJsFWjoCaKh1qyF4X
q8W0j90c8fzmf2hZCqzkbC+bd7nZtjt1SR/Tw79ni/sy0SiET+Vv4DStqfcakeRIdoi8wXASH/ps
KS/g8H4HPbA6kjBWp8JSJ2DoBeTxCtF3Axsg5T+7TU1kNHwDyJ5kvAsiWZT4KwjhczYetcBEJOLM
D1PnAzGsY6KLladd6ohmelM6rB90IfSVyqaGJVxMXcV6hBZtxpakkzPQVuI4cODBduuAvclEz6tI
RW4YzECjoFg+3c/YKWOhIjHoBJ9yFh0+ZtjWLtasWd6Dc9MtqS609+VfSFWFbPmkR6XVHKD7idlt
++wMkFlpvWSIPVgu6VSzqCyUTUAqD5ES3pEow9F3Zzc566+7OcCY4ubKOKRrPHYqW8iXC+i2b16/
nt+ySvVor70sgsBkmqztT1EowLZIG+rY+SumtOpT5P02nmf0y4oQrz3FkEZaqedUmV39J3+0gk7H
FZnm0QIXFv3WUvhBpB5LmrpOQdjbbVG5ajla3JdGD8zP3RfekTguLJ5AkucEN9moa1pR2qdKK6/8
i+FWjAo1ltvl9XT2osX5EVuz8PI2YzAPjywRpMQmkdECCkuJxDsNp8CP8vdQ5VcCcSuYaZgWta8b
iSpYX0ywdffQWD2KHDmAHQifeE+8c/DKrt9v1kp+1EDcaQqqGEXluU+2ZLfRBfG5mOMbbT6nVAaI
rMLEE1Iwg7O4NnV7ulVICMqh2mdsom9CgNh/Vzrj3x9xE4Xwb9KvnJU72mDqf8JASAFsBnBuW7KS
BZPbQQZwWeenDmf66BbBtrzTUzEQ4YzrJJjaVy2oor9PM3UoLnQfjzZZsv/MLv+f3s4fyL7xmzE9
9+6i1fYYvibIQp6UjNr0uEubaXMqY7Ld/HG8dYrP8cjUNxMz0T1wmn2JWY4QpgGdnYVmUBolnH/d
LFei/OGnkaJsXJHxGPh5ILphvrKLZhjHtxYuaeAPOeQtQ/nUZRXhakZT55PTi0CydnWG3+XYJw3S
sDJvbLm15KmoXe2SUSnUze4B6PkZ2q4PmArO5wWokbjEMoZck+TIAtODGvpqLS4ijib49JGEqPDA
GEEakNFUMMoyTBI1sry171xUGJD4c3GleZoYGJR0G9Hmc7VEerw6w1ql+zKmtfQE9ouiVtfN186h
n4MqPmFdyro1rYTWAZ4kZL9j9KqwCo7jXnF02vlglfaXnO99rWfC8FKjwF6bDCSxyLXyDHAtD4/7
NBpLShNQBvovEMF13m38e0vSf9EvTmL6qM5ZmduA6fN/W/gZO3klHAhbx+fZjziVHueemRE/I95U
d/C9NFk0CpurBSCU8+Z5gqkoVEZjkFpmuj6pKgIhY2t9RlkKMG57wzrEyo8daEFK5veHXS6Pgt3e
/ravStPXJ1YG543C1siTsCTzBtZ0rSMaUqIJFvcaN6fWjR3AqXORYLNACHIaW1f0rEdohQjunjfy
Oaq7WUN7NlRapPbnnSRO1/gaDfw8dO37HIlEYDE4x+YUGOBVUKv+b8d01/PxArrOWslwkeqpw0/J
NMd0Qo4LrUo/pPkHRo02E7SkpUcvND3NzOQ/y47VS4UZYEG8li0aZWzXKVhfDSKj7uq4L4d2cl5f
2zQyU/Ea1iWXovoqtJdAIbXkcTiuTgCsuFMXBKGXiqsPCyIbto7BDMLSlncGzgiHHhUSnbOKkN4h
BgsS2ueaduv3aVFEd3QWcjhWyk0WGlioIXKApJserexALDAXCZXmpLNGdeVGZu5/Ds40CHxsrlkq
sjE05uxRREtzOAUnKD56nkF7mEj/nPcpkGSWeoWQQPGxTo/1fIVSfxwVUODrH00ER9PbwkS4XGQE
KINzzNpDfLYQTPp82l9EPqSaOFYGg1f+EJu6RsLuiMY4P/7pOPFRT2AYqeoDa8qoyPtEF77qYx66
TtWomq6Ox7CmY6gWGD2sNhWpvPB2DD0EDPRxP+tjqpH/hnNF21NVZ6OEuZ/TewU0L5aHJvx+dGZq
pBAm/HUy5k8W+QuAYGlSluPwwxhCAEUccVQiI7kf7SR69gahLPpoNm8FQuo7woCAxqDDU5a0OHtt
JhrIwd0EfSzJ6J16ly4JE3dIEL0fr8l8AqCjQ7xFUSrfineHpZjjYw5Hoey4JYSyN3cJ7cgUhLog
uPDrrbwhw437/GfHSIlGavjO5c5Cp6Ln6rXqk4HID7mO5FwuwkV+13rMRIcgMrEOL6ApJpDYsOrU
fHuLQcfBSN6jHQl3Nu8PQK2wX2IxLlxhZEzsLZpCsSHhMJb0dp/CfMkE47WJVEdVVKjzFwYMdAJ1
vo2+jnX2XDG4kyZ2jEaY9Vm2H7vgNd1031GK/Cf5LRHv+51muSPPD80qjqjOUSh53IojxhQh5IQg
UD2yTsMuMCufj+puypmyh+Q2PDNnDLXrwCMZh7U+gHkG/e1aE0FEOgjpVs2y4U8Sun+KRzBH50w9
9YF8PMNVuNZ8tipIfd1YFXyB6fOp5AGb3Z9d4qA97M91zD6vggbIt+s8g/McxCJ81X3TgbbdWYpt
EbwCuff+UGKftc9nij3SIytYw4fGZQViZjkI+/XQ42rxeLcERcTZiB/gWgd3wwZ/CyosrJ0czCEZ
Y8NKkc0W3d0ffTBZipzbXDuBo1RawGisPunocQ87Ug+zI2B+hTObFya71DobtjxQJ7GkDlv4KAt6
J1831OG05pPOMA6wZGnPscXbhk/TssUJqf0AU2RoDROWuDdTgTfNMHAb6/j2rMmg9i+f7MeXkeSz
YcNvYxk0BuWm+gizVREivJIFSV3Hu56wkAzv+lycnN9CVowk46mZO8FVmtBedaKIIbBLLb16K1qA
V9bU94xZ8wYG/xWlVXrhSPFap7VY51BLVn6VHaLIWNfJZ/4EhTV0VrzfPsKN399gJfDgpuKNAq8q
B2i26z46grQ2Fp7fIpu/BONuOl8Cf+no4qwa1VuIUDYao7k1UUuw+g+BQQabHKnSGLfRb8vCPG63
IAliWPl6TmYmQu2GkDieWM0kTD0kqtctmrQS53fab3dFgJT2jQGtYuutzqKZ4h/KngdmpxELEvFq
/azH/LVVvYmlZHki0TY1z5K27NEfee+NXTtwPx85VFTzipkl7qIpk4yJ9gPRvQlltZkAbx1XtRbd
2vodMwY6ik3WBuz32XXptFWK/r+BVSDATUDZDdrmJ1lqkf/21rijnMu/D3GE+0Sh+rYZB9x5SZ87
X0Ck5YBT7pb3uIuijrjX9uSC8PMIJgoVqjKjqhKES1XSfEjeaL8VUmKwWDNcqvtzGth7Zln0PNHD
YUEAwX0dLHq6CHfEMqQvL30poQ1l8eRULMRFdcMqySdFz4frRNCB7+CTyIvmiI7u1o28vrTmPuPU
dIWpj+w296qk7GCO14V/GXPf1wNfit3D4+lNTf3QvWqTBkmbm3hfgshCUoaCwDBUHydKHrlgAn8h
zdD2QqrWdtcK494iJC6P2tKrvFIRbBSkWtsAktECjjtuZr/zjQhtU/CfxlFp2AHqPksn52+DF+/f
cZytaHO5AKBWkVluWTITXR8968DdJnDrJQe0VfSc8Q9erFx0hLxxDfj1ZldhDbUJDVX5Zr/iDcrw
2GnMJhMxTza6bAcMAlxcwISf3ddTKn7Gu9vZFWIv4B0sFCU6iIvHSH04U78fsoXjwRUVMoY5Bjvu
RlcoOQYvrJU9idIOqi2alotZjZ3fIJes3lA8Sm11sB2AniNIjEX3C/N2IPcZXOMN92fophLxg3Ph
vJ1+U8/pFtzxtQDimWQ+MC+zwEi3dH3O7V8vM/2A9/FJfQv0a/c1mqzvmk/aBnGT0zmF19qqUKgF
WgpdAKIbLQR19ZIWyxauCXr1ZSbx1ozkyNHuN7L7dKNK1cHM4+1cUY4Qfl1oZdAwr9+hIsORn/BJ
XK5Edkou399kUvSuB2MPBAeSb3pI67rnyThx4LDg/Yzw7yR9P1l2iILu5cScYHCZ9LaAAFMq1KTO
pslG/GxcUsDGrn+anuibwUG4yjsJXJ4L+DfdZ7gqQxajPRsqhEh4XQ5YIXDq6/QtkV0//FisT831
QlrIg3cxptGS4RxeydR+w0c+AhkiLGBf6j/9IX2R9QrfKZg0sZOrMupl6P88X2MEX1REq/ochti0
MPjWrLa8+L7x4AUFXLtCBhmX5H5yG2vwXguaZaswBXi91O/Q3XH4rNoJSpc7NV4nH3W/2XmzHazZ
LQPArxdxAdRTGZQqhlLmpg==
`protect end_protected
