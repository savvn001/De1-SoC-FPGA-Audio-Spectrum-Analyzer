-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AQ7fLj5DgqPbXmYGhE1QmF6FLyIfzSH3lVlqe3+4yoEmNqdAfcj1FYCuXQj0reWvDDhAcPhETqZd
GMMK5+IUz6IMK/ApC5cGzaztc9iErPrLoYiAhNOyZ4OwLeM7oBnN3IFjYXqicFpbyMf4OC5p5WcL
fcJdYmIHH2jNYxkVqwEl4nGBFwg2DxA5azEavZSlQXe2o2L18mTofifBi+528CXKl8Wfnjb3mtbi
hKml1pN9xn0C2fUCx1INBbs/PNUaUbRK8Mlg/YdbQKwFXYTCWlEkdr6j54syLmx/o0UYRzPgxBHp
BxzvoK3X7vVr12Y4SwcMaxg0HcAZE5vZ2Zfi2A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
RB1EgtF1+RZpOpYpLrQd6yANzlddQ7UDirlhHFVcn/v0t4Io52/+2HICiKvGcI4Hzesr1qsS9aD7
YMxFox2rkSxm4kGun9uUcqWvOBXMmxNUvRirtMZf0Wfdis+qHr+6r7s9z5AizQ2FL4Lu7t30/rjU
5FOLjZF7hSIQ1PEOGU69BWQwSeYkH2rkCSU03j3jonlRc0+ky+QBIagwO8Ey2EY0kh3hRm5NlkcN
s5OcSES/ZxOwR7DZpNUfw5u3gLVz5avPRv7M0twiI7G6SRDwuKdtjaWsfslgndEw/4lP9/776atB
bk0yI9m+BepRsT4Y0Lj6ul85C8sq3ElodyUzulm/vP4wkpQvEL2kQ94p1pUp1fdhJt++uvXH9eIE
lfqANQJTkD2Tk+KOulcGld+SsdZWyyArrvgt/ZSIDVJNxcpTIuOHWyaSTWBhzrxK5CU8Vj9R3W4T
x8AgR2kwVJozUGoT0/zO5g6jet4Bdoq0+nCKtwp5HRw2jodtiAufqoBNCJwlxVVCnq80uLRqPKuo
aAS9MyQxwsIKBkhc6Bc1tMx5oMfDIThYo8McFH/p3DTETDh8JzB5HFwWZ6Tn8pzC3Bnp+yqc3hXb
vG72HHxnemaKEozDqmJT4n0d8tpHd5kCbUCH34wW18ZDcQv9+GvLGDotg1n6uen7+g8gMX/Mg3UJ
yAN73Q3CKpSN6IC8eSes4eMtB/zpJC0pQm4VdRH2BGdrwTb2GghzaH0+L9W7NhHiGt2vgIZa0W8f
ag7UnTP7k3X372yklhesV/jNSVvuMuA7W1rVm9PsFRrnChFPYOjuHwFtEcpg6RUYqhre2xUdWH0a
abQR+yznJ9xcQb7HLwxK38WTrSWW553WDISmWX+65IK0SAhzb3Gbi8/grNV0jbxdF7NF/49jK0tC
ovTCUWH6KXA6EcNbnUOoqMKp92RdKvdVAiKRJsq8vcsLrJKWP4ITMmQlVoxBqL6rBWaQ7icjdxCz
aPvv4Cfdf+7FluFkt0B5BMCfqN/WBoQNYtja1GZfI31WdqYifgcBhlrCI6vTxCrFOqgPoLsCTvS7
MSjL9psYlbfqEeNk2skZxJtzzf5wpv/Ql0THKkKVlwfar9bjiXkTUw8qRhZguD9ddwXh2Bv7OXPn
hGEDmcm/6KyYdVysfl5GtYdIQEjfT8kBSwJaE5JBa31rfpPIm6s0jcjXfAxQWGRPvf5Sed8tt0FF
WJG3p0yGgNttOcaYG7s0i/0yQg3zGxHUmk2mCBA94DMxaHTNaMBXjlDn+eWkpVwtmpr8MopJ9ipG
+Z0uRatfLkQ2w48/2EO7IHnBB4SVNAtoXt362AAi6UgpdOPxQbfX0nXeZexYYcrciy0OLt//Ame2
ubddGhG4pU2zj3mYOQAnUhUHPF8QtzrcOHMgxOIM7xdE/bBAfiLoT1Cza/8pBnXLNzMmqUokajc1
blK8UAnSoNMK23dLy0d7Ao8kJRkkRgiIL0pRPVHXCI5TrqkGitrTeCHlzENNi7WG+rDmTbW4I40i
4VUTKdhd9DfpbVJDPVNm+HIBh9+aqoP52N5g+eIyG6c9+HYRSyVnMcT2VieBxzcPRAaE0xYOt8wX
62ZwuLnV5b34fzHrf5DG9uk/EWChN4gsAcc7CBllREIHt+VffNP9COesnGg6pFuInxomjvI6n6aH
xM7R8d1WU07NzxsFM4z4RsF1UpH3qSDwQ5vdpl9s1zPA4xU6iOX9uqy7mqXWIW3Ss06d8mI0ET0k
mWx/8J+HDujueLkz+O7+kXkAYxte75ZA+tqTmWrK0WBodaRUlY4YHVnutQuOg2Nav2xa0sdEqZgq
Aj4TXJKT17fNurQmwyDBetnEwrilox9kBHtVGlpmLc05LwgK31FqYtlJQs56/he/pcZbb8c/5Xw5
shcYIr3kz9FezjZ+zbIMCtocLhszl1+CNAK3z2WOuh7PKCr3LXtWJzyOvXOPSNgb0B81KBkSDnDG
Ncmb+r00xuTnKM0ftSRaZrMADxswme0dxEM0JCIwy9D9orpN9x+p4kMQ3zHSmIkMrxHz+hvBGKWB
zQ5bH5dn5YCrTXThGODglvOvgy0bkm3SigNcPPB6q999n/w6On9DBx0wDOk0fADOId6ZM6cZ0mO/
I1uBPWjXu5I97KYuwAxPmm3eGhP9/rYA9Q+NTFPwvmkH0HhgSRkj0C+QjW4f4hQI2GRh+OZ2IslQ
4MoLa0ehik02qfuvLAQcawq4nDOFsNLBMzOg6zzvV4R6ooGvreDP3n87Ih+A4dxnczB06euuUztt
qlGCjXZjmkr1eJxUP8IsLiGEYOK0T4zeXKwATuf+haVapmNWiFODYT3GKN6OvPAardJSp8cJApDg
hcBuxJZJP3vMETK0nvJBdSFDSSLL0rka4Az83V809F423TBBNnX/SsqYpEOkqwi9D9A2w9n8l4/i
ULt80CDPx/MYagKVYfsrBBlrX0f7kG97JMeeDdckvhZty3hrwL7j6L7bSpn+WqrV+FV0XteS9M6R
vX0r0kExTomKbFjKXx/mfAf5CDLujiE4MWBeaYnypKrHoqITU7Vm/JD/3RsphkBn8KyFysCo0w90
9VjGgD68RyTXOv86r2OQXYMIOfYJOaYeGxSeo/TTcjsk/C6GUHB9hH8emU8J5AYYZo3q3ZdSJx5l
jqtjfg7ATpEsKQVO5Mnu9pqSCRRcRYAX9WY3ToYYhyPhcZEegR/oLkFxDX6E+7sxhb4ZjKMleIcc
vR/vpk0vt/vmvozweUZJxmeWF1u0GW3OuVbRHI94cZh3Bzpmdhr0XlGrSNV/mYFmQcC5jzdyxR1j
nVWGpGbAkpgOZT4/w6kWV7k5HB2qVkWxNYlZxE1s7XHYxcLsXArmsTLKwf4NYpRix9i6frs+PCxx
MiWYSJZOJYJwMqjJVutX8BARSIuOAQSUiparbk+Xn6wJTlBf1AL/ow4ENlycYDbo723HGZXVeAwJ
MlsVQYKWmgff8TIyoLSdWkgY14v4MCPlDx65FpG05HQJLnHvD9xfiYJVK69UrrAK28ImpBCR2Ory
z/nSp5S/raZSCMbxLMK2YBsDPbucjnfJqt2kMEe5ME+Mtr254haA5r2U3iFSAq2lME+vg7qI8Mvu
NfuEkLopDLyRkFaz7UfsdbOKiZRVnkJLXGbUFZOSsbPLMWLD+WgOuBv+1BXIbsqGLd+t0P2TAw+V
EdUWkwExxzIPzZzpJthX73MygCxlVG1mKwProSN+Roc3qAdgWkXeCGj2MSJ40J+HPO/NCybn1OA6
ERYMO11Dh74L+gAS6iBuf8EzVACLG1QkI5KhNEKEvTn5hJZq9ZD7zKaRPIk71h7lI9t8SRzmwC0F
z9nWA11/RQDbyBrItjVcAFTWO6S+vEsuZDFlvfXjK4RR4/MPb6NlU/QefcKb/A7FkUiCso837MYp
DQ42ustsdaJON4DddJDYVpVDGsguxuuIw430UnLAx2G6qjL+VOPywvfP7k1lBLVzvsJPfJP9oUuK
SCAXlbVddQlRQABWvJZI1KaUnQP7/cGYYZGnG5ZSkLUKzaFVIXxI0U4qaaQ+VbXH4Nri6OKk1oIu
tvcZdJFirOpZwGOL/3Bvs4CzdpECycx/4spFVgSbXJTnLfyvu89ecd/oABTPOcxM/MK0IDdydJnM
7Gu7A4SzdB4fUCUIVSEmKEP0FxKQ+lmKSxrGJPFzppZdAO62XBw0E2TEiOTz7we4WfPLoWQer8+o
Etfi0VlfYeEK1AAmhi+a0olxFQleg31kcV+D3a5RS2UIZIkqigXMD1pepl31q8QytvaZIdojM3vK
Q2dNz/nq/fE21kAjP1H7YxxKi8R7TZ9M0KJ9hKFp7UpdQvRpRUX+OpxFM+WeBV/nC5kl56zxofP8
0XjWsjn6vSjxTCnslrTj2cw5SR3O2NrJTNwp6PWA6DnAsa53Q5M8CrkeVZlsW2gay5F+pjL1VLAC
cg0ZVAjd46MVoXlSYm4oWfzuEzFyw34tcYZBFAOvyR0BQpL6Ws9tSGQja0KdpWt5C2I+nflPzNVC
qsXw4wCkEVmXfPvPZfY+VqM1jJ32o/H7f4eFxqWqYzsP6z3RT9pdaUg+ZaDJFc+JkpX7MrEVNstd
cP0mJ0euw4jY8uAjLXZDC0S0hFcv2yeJA7c0ISjKlV/Dr4t1tGj6x2lFAAXQL55LSWVcVNoI0p1v
Uq5WlWNDuWqZlTGl9ojLJ/pn2Q3GvK4bgx88CgDO7UVkifKKuEVW1Xxen4u3Y8xc6uvxR6VWTW+Q
drH5/eyVAHbWJL0oG3+SaJoYpfOCZhZA8XphdcrFqg8a3RGjavJRo30psj44LCFQPRD/J5HWYaRv
zUG9U37IGSv0yGR7ze+eynY/e8UpaXcwNsMHvrGDrHAIE9vjk6sJ+jL4621dj7mS9m6S+yak8vaj
FpFeo+xYmHoVNoDplQQkZmaxEXeI+VhuLNk651LPcvxiHgt0KqXKis0dxo8ZAT0l8EJKonVhIAig
2L1VRaUFud8hf7wjxsXWNhhjL9g+OL2/XvLZL+ky04SPSDw1siBTH7VvTQUN6hbQMUOVXabfDOpm
k0BbS2xRk37et5dIkuJbN2de/X7GmtOD3odK9uGoD7wdhIkBBN6g0De+hYY9LavUUxRtXKjZCNXM
szedpy+oQ9gef5YxJcPuaju9Plk4gSXp0/19zt2N6ITOp/ga3+Lx3DOQ5YHMk6bGi9LqpIypnQDa
At3ntT/CaDIsAos2+4LA/fg3XJQN4lhCPXOGnSx3M1IS8mKxtMBDLw5G6g0tpfCJCJH5AOWonsrC
7ALBp8SSpQ5/s82wzmI2mrYnvMAUrnkH29wD6Ygpj8iaWyQ2BRozL5Hx73vQCcEKjJC7L5iZmcRX
yQOb2xlmXcg6EYtx5OcUwzf/udYTedad1cdm6qvX/odSks4dkK6stK6caVvf46MAevFSao43FfTG
mXveeDfauX2OaDLMNihVFC7CrOPdMz98HUB2Bd9Kv/Biut8nMTUCspn4NDskCppFNN6OdLFFlqBW
R0ohFlvu9HqsN8RUA+TzqNKUDrUdxpFb1o27mOSi8EHP7axZaxUXqn2SaMLpIaD6E4gIqi6zj9la
87qEISexZGH7P+rw7EvfcHugx/eWlwT7Un4u16EPaG3GLqltuOXmLqBj5iTUmz1hEA8pPLwM2eBD
/4NBXIGlvicVuIChgs/NxihRPNdcWVXOby/rmutCkRHnIXc4RPVwMuAhxGIrp/rrE2U6xU2tb/bY
kBItQ0BnXP+tdQ0Ol7Xwvs+AaJqbewMVxUHKOYp05uX/fkiJuFwNTYyeceP4FsrHhhRpu1VV4mkw
6vpDEr15Q7AFoj5z4Lle8owCH5+uWN4gi8PqaXrZp6xMUJQ+HHwBixvq4ldqM2U1G5yZw3k1Ciho
yRGDlFstLxAQlUpZxfMwIQ7JzuS0Y/cKAKpAIk6QHor5/153bF2JlPCbq97uhXxfvpO+dmZi84bT
dFQN6KukRV6lUAm+dFvjvJw6JvwZue2nGSmFB7sjmS6jJI29q3o/pEYh6+h+qSfYHDxoZ31PSH2G
W9R1IU634UUicZTBgvL6RLByNwF1VBZDuiZv59u+94e0Bj+d8dQK6uGKnhW6XjKnYIY0qc5VwlZa
SbP8FcDJ4Q+U/3XEGaFDTfk5j/MjIFwbXvH2NzgNusPGwIYSK4/k+DzvMnf/3yNJ3x91SwN4gVa7
Wn3I968Bd5r83bDFyvhgbnR792PC9OaXh2Q7JRC2Ybg10122hSZHN/AdYEGRcmBqmRlAyX40h3uc
H7uykF+OCEYPzqIuaStbItIWllRUC8YFKwYFChm1c6XO+I1xd6sFs88iPxDS5Vbp+apItsM8WlFH
7DWr8gRLtMezSoV8wDuFq+9roex0POcvBNRqTPA18+3oeMrpxlQdj/lsvNYWuiNbk3fbZTI8mWVP
lWMo11y3Rp0gnKjlOx/GvTpSlzNHQZaqZKb1Y8iIZhozUICOrVfjwPGX2hY40whArSEeWTa+qoj9
CXwNTLyTYQX/8thlM2I+TrmSqZs51JBRSrgxKXUEzYo3G7wa2t4HQTtGOn5zXnWk4TqmY9j4WyKr
Toj6RIyIslVgS2Vc+lP2kwRZtyqHpvhhhN9dOorGB5tBidqtnXfSZpRfRNTVRg9EG/rGFUSahCkx
y4OQ2ywPD24P36uAlu2pHD+4Q5WYDCGk+J2eHJfnXxB6fxlHc9Z7zdG9ezCDHj2jwos9NF3l45oe
phTRutA1mrDKwm4ZxMbHMB5tjKY53fBgeWIzuJ3hwKeADEdgYj9jDukiNXqm2Bnp8frmQZ0Z/os7
ikrJ81r84AorzP38+J15g+q/BTC/qH3VdggOSY3T9kH12C2PWMiVT/+olS1a9N1XWt2jcxGcVi1V
ce8dcuCIrM6Ip800AHQ12/8ptNCOsGAAbmcF7GpmeA37tM94+FUwXlrSX1+Wb7y/6QU1GxD/BvBN
YJGarkB8zpkA5cGZCwy6WkiLIBXX87YGNx6vjWJVhAKAvHyseNa2RFz5U9aU1SeOJbNl4/ipBqpx
ZqyrnrSyWYU00cvNLcmhAjJJlC//X6L+sslqezrD8ivO+i53JjFJYnjaX5AgwL+BdwQfYdoCHk5C
U0YDBp1TucM6G+W+RA9JvJNCV9OQQmgkDNU67KrC/7xInWd1aS01PFOSSLjVaZ4EyzYLvQiMuV8Y
nQEAB8h9BH7PGwSH9OtQexYgHs8TqTjhYH6QhgKX9SQBFE/8PVTZrSkoHyZ0SFK2sLArhDm3Td6b
qS6eGzVcYbK7ehiaEmXCk1ciKgo+I02jZz6Y8KO4zL38SX2sAr1TwdrGli/8/oxXuctEbhX9w6FY
j85aH4nsDnXWYY+Fd+uU3jQJTzRTEyS3ID30jvzl5/D3m9JDy6MDz76LO+552jN8sS2Dak/XvVWy
jNgLGgYqyvmmYDS3henNncu+uhqvqaVVY9Lnu1P1WwaBMnhtZcayGZ7byZTMqhSqYuQKHXxX+yc1
3F1e5u+YX5zLmn6NQFV6Azwyz0yBND1GEbAa/DmNbVjDedMb5kDW/0fvtf+I3mwWEFaYCkCzcUJY
7RZtpJaSEwlPFz7wq33L6P/w64TBCM9eMb+aib7jdEk/9mTqPMGlJMYMv02QKmxNius2S8mTQgJm
RqwrUomcA0Kheif8Hqr/DJ9lyzF3XqOsWzrApDTobs8DVi29uYLQE4XZBWRwAv5CecAxRVVNoYQG
X6lARnqTX3O0pKqX106YPRMgyLvpLLmfqwzXuMG2MeV81hEx3R95W+uWG2Es3fTPfHcSWz3561R1
sa6SwEwJYW8ybykXsSZQ5pq6wsfczMcEGpvEy7lApy1izq6tf168tgUx3k6EWNbeq24wjDqMj5sI
bm6L52y47usUDbv4RcxWVyjEEnH6UBXAJWPOnN0KAJ9PSMBowRwxUWOdW4hJSJknN/8+TddXFpjX
4HuTPWcmJR5LBNt5q2DkhtACrvjZFP3SB/BGzq92mUwvQbXReOE0LcUXf4XAmyFI26mMQJcDm5t/
QCdR0IP8yfHEQQXvYGlM5FtlUsVV8lXA98QnNSR8jGQnRg137Tzo/rW6JD9nbmmYevkJkjif6mAH
9YHIOPP8IDXaM7QW3gMcSmVEub9GrsT2bYxAaEPkhHUKHT1pFMTdOA6Q7/RcoD3SCMIP3YLL/aS1
9fmKh/tY4ldJ6ptRqtTA80FCoxB0SNoWDDRzVd47ij3GJf9jHg4P6av4byn5zgjrMp5OOfJqzYDB
VogZFybZJ9sDC5xfq1g86Dz86AVrYeJiBj+B9Zl/s3uGIr5qnT7WOGWflVP4MS+8sbc+eWRvktNn
0QNllKvyfx1oJ3kvhQhpgkpU5HpfaUhlea+gO6ulQGMaLATE5JenqGMyiEVKz5e62VXaAjpQsA6Q
tBS28UIBwsqu1wsRGjlJGdzrlhXz69s6wx2U/PjN53StCi39xDGcQJAgkxqZ58OweNaS9Sv/rJFV
3VamGHZSCikL+DOZ6m4as+QA8XVYppwA4CYdebZ00bPsi/0wXHEviPbCz+sfHGCpDf+McZRoEVIm
zKdNogZHY6pKCojILAshNdxEjHvVOXlAR0zxK2oSWDUAPMdFZI4yNEhP4zBB6KvxD9tma+2byLLv
I0GHQQjAtBgWWL46JWOdKN/yYEnpjZkRu4KUJLlDZvCgnB82fqBeSkzJQvtwozX+oBwC8tVr++ti
BK6qhFNxtdCG30vzmfmQ2KAnXdM/YZRDzqlmBjaV4ZY1lBMEhXry2DKlMmikTxS1yUpjzebGkrKq
qNSxmMhpkwyNvYa2Ok+aGRsrSyw7oxBEF90AgTzW1sz+1N8FgHdOX4lWCHh8lpnLP26Wd1pjtdaX
/aYkJKoQQoTI4j4WykbURxI+r6ja1BgxmSbezLX08CwhMc5dWQc2VTpQXCb5mqAMnl5VPozQXCyF
32jak0j54P7gCP8Q8FiuqDeOrfGk6B/5Z449ZKcHHU6ZX3Vpkg1HQ/x21OKN3fpWJBCkDI5l1i6D
+v7jhVng9jR8/Xxy3zA77/RMWXBc0bOVGbqcnF3DEwYMJiP/cSMEYqBy1XS6351tZCAY/tV25+mq
2f/jnfjZCzhgSLup32BL7NwoiwUG7u6KoOEgKRodwV/22xd3iFMLdBPwRodb40RIKEaV5igZOEL+
wAVshdYPrIEXPOXlfoehyIb5vRuFsi7RMIM7kUi4lRa0YXWHDlNONTWzicljs0Amc5WY/afORiuF
qcCEoAgGJflGZKD2sXZPAev+k6eOSU+4RaHCqD/dvga1dDyfhIvFA+WtaxUMFThvnLfRTtCsDaMp
GYyhszgP1EgweNFpLPxwzwPRgxzppB4vj8T6oKKO+NdoLbTWApDpB4EjXA6+cys2JF/WvaDn9ROb
mMXC37qVWW0c/jtMtwxfHnHCmxJrr84jFYgbfU1dOCq5ue6ggLIcFdO0kugyGogQDySXM7v3MBRM
wJmGcGcNw5X/hjOFEMVORip8tzE9Mu9mq/BNwHcNVPcxBSF/+PaZ1myN0YJO45TuuIhL9FgI1e3V
Qg==
`protect end_protected
