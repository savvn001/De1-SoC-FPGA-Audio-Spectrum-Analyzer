��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O� ʂ�U
$�PZ�,犯h� �I+�kod������ݰ��l��K%�4�ɹ��KK]!c�ЂN��c�Y��{ĕۨ��Y�K�d�:3RL�hx���p�g�A�R>�)v�h�MeG( @F2��aJ�i�m������<�H�*�/.`�L�9����V*(��$6P��Cؕ�f';�CWg�����7�'I�rNO�
 �|�����콒���fK�W��Լ��O�3��Ȁ�e���u��y��)ܸ�D=<nʘ��9"}��i�!S"��&�Æ@`�]����U
�J��e���T��v��{@&vXK1(Ո���	r����	�b�Cn�:��$&��1���'�v�wO\l�ɺ&@?���}��=�W2��9�a�
�����s[+��?�[�I���Gq _��I�+:QA�����Z��	$�W�g��Ѱ��%�</�S���~�6��S�+w�P&����Zp�����������HUgWv��M�����ez�+X���Z�V.���F���u;a�/�i��������(�L@TDD��r�pP�T��E��Jf��	9��Pݺto�zQ_J�`s����s����+��N�OS�K�-X-��b�E��6�
�Ŵ|����!p��/n-�LnGe�<�2�ގ~�Y�W~��3�84A��B��h�B��:ގ���־�b�$l�̼ܴ��lp�i)w^�ޢ����%�ީ	v%{��/��*J�N�GG���
��U�Y���~�"�xsc5��nJ��0��HC	�^;'صq�� ���:��1} ;�B���3��?�>�N�&�3犧���e��Y%@�H�Z�;(��+�k�t�⟌��� �kɇ������Bu\�]6*�2{EAQ���-kZ��a�(�.8�X��h��VTo����忲�h������n���nJ�C�#��jX��%�ч�p��̮��n/P��@q2���.�0�KFE��}vP�q���xg�h
|��� �᷁l��Ug��HX��*kQI��n��$�@��HO`���\Vԍ�Zadi���6�DX�~�s�:��\��#k���)K�(+���K�<�bXqQL��O�M�{%��e��Z7��Xc\�����ܾ)�u��Z�fC�}=z��L/X�ٶ��M]F�s$x�օ����3NsF����?k�h���li��!�$�E�O/Li�̶I�'?8u@��	 i{mJ@p����g,�/ +�}�K�b��=:Q~��y�{\ϵx��˛���_Ю�7,��m��xOݡ1h�AaR�࣓����ZX�i�L0�@Y9扃0�����OA��#F��4L��	���ӈd�#��� m[(��3(����Vi{��<=t�#466� 3�^jy:�݁}����Ku�A��$�1#�j�`���(�O�1+~sx>`��ߣ5S�q��>UD�ʹaR2��2�yb�@}WD(�̈��cR���?Y��7���@��b��_[L�]k�8g_�Zw��"��֤��$�A�C��P�<�Pĉ�pq(:Lk.%�Un]�ٵ5�~�e������_h0��9��3�v[���s��W�Z�Vf�\��2ERh#gU��qEN�:w�\���s��٥op)}�-?�`l	�rFA���/�9�,��c?ߙ�-5��z
r��@�!�J�Gۏ�B���tK����!i���rd���e	�*���mi��s����w@SY��OO��K�|>7��ll����� iK#��?�:j�����;�^=Z8��bQ���� �a��%�D?�c¹�ė:Z��P��c:��	������UT��z�f�DZl���\��k�86�Vn� �T�>A_�����p.�1L4��ֆ�]`���7Ķ;�#B��)m�_vV]��'�E�A���y|�:~{#��+��n�͹��d�Fx��Dz�U?>�� ,��bfx�d>����ĸ� M/t	�f}<�Y��ڂ��f|2e6��q>���md��e�����׭�7�U�9�2�{�����&Tɰh�uQ��UXj�q�ϭV�X��3�U�5ib���!��붨PT��H���D�3>��i�t�����
�d���x������O�EA��O!FP⼗8<���dB���XvM�\�J�U���&�st�Ҧ�p��TIA�,T3�` �<���X�f>��,䇿���%�iQ�?wka�`��a�8�L�̆ob��G�:E���)	Ƌ���fG7(ɤ
:�����$��a������h;E��ow�f.�`�ul�'
�j�f5�@�z���=���$�4)@TU����J���8�����h���-�/�iDƧRq�\���D��C.铉���i��ɿj!��Rg�
��d�=7[�J���ޖ~]*�,��<?z�����ȹ�l���W�s	)P� ��_��jtrp�Cf	Sōhh�ƯAn	����%uۛ���M#�m똿���l�����T�-"�[�ƕ�Z��P�9{bZ|8l2����
���Vl���1��j%�^A���v�u����Ɖ~}d��N{�Ě��ڴ���%�Y�_����-��Rq7��*�����<�<%�kI&>lVn��X�%�e��0Xa�O%O����$�G��oǺ1�(�cI��g��`����#�j�;���-��/*�&Ä8�	����S��'u	���ː`�����e�����Z�"i7��4`�*�s�L�M��TA^A��X{��7w.���z��\����i�k[H=���k-���n6}���း�镼?1����O�������:�V�1���ʥe��d+B�A dv���D(��P�s�?����x4�Օ���$��a�Prg�W7����M��jQ�J��ʫte�G����4�̊�EN( ,OW58���̨^8�i�^(����	4j�n��(jN��J����w�#b��<���`���	��W���.�M�u���]��4U�+��D��J��-��|R����X�gs�V�s]V���:�6���&�]G`5��ʵ�
�=�ܕ����M�q�/��8����=�7y ���VyiJ4�� q.��z�U�Y���!d!�>@�Һ���n�p&(� �j��@�[tLǒD�-�l\�H��H�1@�i�j�\d������]q]4c��)�{5ߴ%�bi0�C�S384+��D-Ot�����U�78@�d�.���[q��¤)�`c*X����SZ���p[V2�5�S�{�X*����� �oa�!�RFWJ6 A(.�;�C'��/�F�9߳�𺿡}�����A�3�gt��.�F�rq��Uyr=�m��Z�r
0�]qD��tJ|=ws�r2Ql�eJ��;�	�w�SE��ǹ`�^��=$8�!=�/�<�%�g�����11%KO�[���)�@.n���ϳ���g�L��q�1�pB���"���E(�p��jf��N� ����ťFgL�M!8�y�EG�����=a�X9R��L��2m�T�:�f<�#�k�5 @�X�M�ȡ�G������z�X�<�Ѵ!������&�Ҵ��S9��s�u���6��ٕRW���� �z(�z2���SVSnA��_č��=��%8�dWm��Ht6��H������{�d���i<AbU��/*',�ٱp�Ά7��~�����Ee�[�a�Yd�6�5�W�֣.�^�Ι�f1v?�K�b���C&��2�R�I�|B���e �4/�X�5{E���W�b�l3��t%_Lk6���q�;�P'�'T��F��Z>��$���u��,Sjk���ֽ�� �Å�CD�Z�����~ЭSI����F���^���>pRҿӒS
G�g��xI���]/���HPyc�����M� ����K�S]V4*����v��>ny�}�,�ʎ���M���k���`#eXI�5>�;)O�p�鍺Ӓ�hrq}��ݺ<ي�4ƞ��F��@��WV�N,t�[�^���v�Klh����Į�{�j�@hA�R,���L�=�*�2�'(ON�P�J+Ĺǂ0���l	�����\iK� ��깗�R������a��*>�:�t�ίs/�v�Wg���}�â��Ǵ�E���J�F?��8�9�����m�P��[�����o��i�!Vh�c�Y� 3��o���*ﾨ�!��^���yZ*{S��0�\MD�{tW�8����z���ֵ� �Bƌ�yy�)�Rf�~6Jw���o����dK��v�<y�(f� >y���'m������b����V�˂__��--��?�N�#t�kD��s��ǆ�G��hM/�:�Q_K05�4Af���(ϰz�����X�4l|��{c�h��YP��-�6�$��̋�2�!�8y�9�����y���r��7(��6~6[?t%�m���G��HY[1�p%Q����X�ޛP�EHLk�>!���d�7���=�/D�bI��Up���݀��[a@��sn0*}���&�G����}ز�3��Fk�$��e���4m�;��ݕi�=�E|f������#ރg힤 q ]����vh�Ev�<��.��W<G0k�o6�u�#Na~Rp���/\U�"��~ݗb�[?V��Y�cHG�qP��p��:�i�eє|�PY'�0���H��,�L�~x� �?���,I�DB�E����G/�r��!g�P�Q0j��V���m\�[��s���>�	2ζ�&�
V�z*x�5T`�
�ZS5'IZ�h]"��tHhw���n��f�(W�c�Fw�-�L�0?�K4q�r��O�@5�"��ˁ4���}BP#��#L_��^�J��]��`�H�IJ��ᬙZ�tl�h���
n�c2[ӈ��R Ŗ������a"���R_!w͑~�^�rz�O=iH=�<@ƙ'����	����X���7�2���WS�{iK���Yj���	����፜D�;���賲��)|�����i<��tg��~�8dEd����ǐ9�:���;���ŗP��sr%�B*�\f�e�7�׊��o���d*���0JX3��P�Cΰ��Xi�a�Vߝ�kTvg���Rͦ�K�8��)��+03jك�	�-����p1���uز�r�],(�d�Տ����鈎��خ!�@��JM~V���.��r�R��;^f)����P3�J-�o��R������'{�53�'^8���S.-�{�u�3��a�����\`A�D����[Q���w��# �a��W.���J[��Uˇ`���q@�08�N.L߱��§���TK�Pto��U��<G�j�|��R�'@�xV�㐇a�ahP�C��Hw�#i�;�C��S/���+ep�pg���
pv&��N�Y��K�ጵ=��%POf|M���B�&nL�gr�g�6f�i�+��$�8|��7�=EC���-[�߄�9�[%^(.."e�28���܏�%!�k;��EP�|�cZ����ê,�ʵ�Q��*��h_C�I�lE���hu'���8���=O~��Pp~t�I�s���{���\�V��ڨ\���Af=2���-"pH.�P�t��H�^��W"���tYk:��u���"g����yY�
C�F�jy�c�,?��(`��k���Y�hO��U_Av�4J�r�]Lm�X��o��^��H����<������Z0�?Ǵ.,���h��R�+�)�O��Ȧ�����T#U�{LY�ex�p��Sz��:�4X"y�y��儥��&�7n�cTJ1���]��ʗ���зP�RQ��̦�@�0KT�?����<C�+�M�z� +��\�V���ŘZ%Q�wL�K��̺��h��u�i^�	O�iN<|�����"��๲2$�9���j�8e�����)S����]�1 i �7Fc"`X���B�y��u4�b3��˞�va��{�6��d�(�z���׍/�|Z9Ƚ;�JC��kY�̀�>$�o�Ip&���.����e�y���t���-�����l5�V�n#���Pqo�g(��u�>�1ֲ������
��V�v���LP[�����t�5̾���a 8�+]¬
JCF�p����d*W��M9��XUE�/�A״[���E]�[O}��e���$�F�����{�2j�B\����v��ka�2� ˵�CcA�²(� ��%��~���pI,ID6����9���.JI2QZè�
���%�")h��i9�����H�6��'�s<��2Mg�|�./�!���迒�)AN�����ŏcl��0�5������R,r��C�}o�T�Y���AB$��YG���>ڊ��� �TZ-y썩o�p.`ƆӬ+�B(�"I�D��X�V��ܜޘ�H1�1F諥�,(�J+�V�B^����ʘJ�p�[i�}�kR��s�0������s�S=
�g͹��Om�����Wց?[ҳ���N�E�Nm��j�9�ˁY�~����W�R]��Is~���b����.����V�Ul���":pW �0���h�eï������r@�b�7{�!��u�<�)��yUɳD���m�(x�K��x�P
�hka���rk�I1��-?�7F�xu@�=:D�$��c�g��t�Q��Q�[��w/�����h:|/t�?���	���ۖ�B�����Z)�x֝���(B:�|���s�O��8y�L��M0|;�Z�r����YyD�ye>��Y�v5 gፘS�����v*�ө>W}������tzm�1�SE�K�?
�xeݭ��|b��B��]kvAC�H��`�(�Z�S(l3����Ddk�Bz����>�*���r�-����B�>�n����:������AX���������=�&�"���������
�A�蓱��B��!��A j��A�҉f�t����[H=�Y�b�	(g���|�8|��mv��1s>I��T 2H.�̉��K�l�B�{�����c�b��V8��W���WB3�޺g��I�_@�?Jw,������R������r�S��S������g�h��6�2X`t�60N|
�Tr��N+�.��1�`Ph���U�#��"M;�5�~�'8�Q��Q�m�I!F[��$>/t�%wLC\&�|���c�
0�Y.�R�
���c�b�9��&��)����mK#E5�}��ml���^�J��2)�� k!Q��O���~)��}��	X9�9�6Ŷ}X��}�C�l�mDq��G�%�6UM�+�BR.�PiL��n�o�>$G����i5nN��XH�/�K�Lx���с�<	�uŘ�ĺ��}�����*jd�~�;�`/h���6��J4A�nͰQnj߰�Y��(��y�ؕdA��}��Ds8}9������ ���r���|��\�h%[�c=F����1��Yq6���a7�hR'�����¨�"J�X����8Y3�b�<
��F�3'��3Imݘ����rX^`ј)����Ӧ��C�}U��{���H�ݒd�����h�q�ub>�������ܠZF��g*jq�#�*�i"��2����vQQ1u�ugy�.����g0Qg��#0�(c�?�̜�g���Q�z�\�e�#S���{c͘�*�lT��������3���'vA��bbqp8���_z3^Y>"�����n�E|���ߩ������6ɾWN�����e�������r`*���̿#L���.3W㪦3S-�n'�Y��	I��a�������l�6�+S��)_ր���/e����{�����ĩ+�jJZ����3IȨ��EO��lr�.դg"�Yil!��6��Fk��3�i�_?7�����"w�>/�%��h���
4��{@fO�v��i�/��+D�e+4�~骠� fR�t�n �'��L��{[#�`A�_y��hqs���z��5L�<�+H\e�/��d04J`���$�C���t�q�
�'�0ԟ�����СS�@e�#�3T�Ε�*6�H�iD��MA`ۘ�P�d'9�k��m������ma�;&�{�5�Xĺ�7��a� B[�03����m��;&��P]H|�9�qP�o�EQi,��Y�oA��1c�G���#ذrOA�R8��A�ܷ%�u(*dA���Y*+��8�.�V�����+�Pkc�"laa.w<Qq󕷄�48��ݜ~�)���N���N�M�?�0ꭑ�d������t�JY��} �	r��*��n%)Uؑ�Nψ,U�l�
�<	�]:��]�kKđH�`k�|g39`��o�@�}2��/�����k�Z;��ʎ���]��8Xy�<�͑Ry�r:�߂#���6�|�
>�5�wU�w�t3���;��5m$($fI �QY�{��el����-&B+��+��'�>��ky�6�����gM@���	�Cr� ��ދH��4��"��ЧH��X���}3�v+<�¼� P����G_���,�i�Q �sD��ϣ����S4�5�|�oh#*}^sQ�B8���I�����[��5�]$Qd�����҅j�"J���kR;� '��ۋe?�9f�:���*z�-*�2�+�z��Dr��D�[[11����M1
��T鏜��40>��jC��d��3C\}�y��������]�8�� m��K����K]���m���l�햮�2ŀ�_�~�&t2��
-a5���o�>|u^8O7D�5�?>\ȃZ�9=�g����k�4�L���$�B��;�x�\�j���@5 �5��5���+%���5@��YR�Q*߻\�ݙ�&X���DL$���鰒%uq �8���F�4�S��߮d0&yO�@�ل(a1N)���F��$���0��zńK�&@]f��Kq�?�"� �_8���r_�Y΄i4�d�ZW�c{�������p8�@ �:s�Eݽ>��`a<M��<6�M��<���u6�ܙ��T��A����E�����?n����6eU����㠴����R��52نG0nTIX~յ�Ү�"��J&sA٥r����5��.d�:b}��'�#q���̥�=v#UvE���5	��ë|T��_��Ia�?��������8���BHE��J�WjNi��^����-Ԁ��uQT..|9˱,���_sw�0n��Ǫ�o��T���w	�#m���YI�p@m;��z ����g�Xq�|������s�؆ vr"�R+��GC0��;7$kg�sI�n9�-ơbFgh�	7Zr�l�EXc_p���/;r��>�?ȃ~m���oN9�(,����l��8�H_g��Rѫ�{�T4�%D�;�¦^�
�շ�Mm�C��;�Ъ�"ȗ�љ��n������}\0��Z�K�L}���N p�F{6��yY��!|�ݚ �|��
Y�g�M5����%�*��1]0������-#
t5�(?���=?��\]ލ�@*���Zzs���nն�����}�]Gy�����~�J.m��M���K�P@B� �	�Z�5\-�y:��ϩ�����(u�/@�tb@�O��_��F�a��V�t�����c]ڞ�0�|��<���ȥ���	�~��pw�gqBf��ys]�Q �6b�q�Y�Kٱ�=!�m�̊hE%K���a��7۷��d���Öq/����R�����n��ل�8��WI�1y���,�W+F�yV�b� �J \OA�ߑ�d�䁉yk�|�zc�g�m&���:��vd���oS��3����E������3�h%��iӘ���8����sӗa�l�u�=�'f(�L�aTB<���U���4k����jn̘��m\���`, �k���B̜����s�Y���&��� ���W��u�r]�e�5�Hǩb�{���ф����
'����<�S�ڨUD�B�P�z���")1�W��R����cf^���
�J�	�{�wvv]AhM��~�M���₽�Z7@�X08`��&����4�;t��`[���G���-�%�ڤ��/��Gw�͹�X7���$�P�y�if�ߝ͓��>���b
r�=��`��NϚ�滏%�A��K���/�mʢ��}��A����?C�bL�9Z�ڨ���Toe��24v�&$>��D��]z���
h�$����)�x֓m�N���X��Ƙ��;iaRuj����l|ƚ���߬QQ��-8'�OQjG=���{5/��)R3B�q�=1k��nZ� )1eq4��hܶ���i{.Z ����}�$I�B��$!$ʘ����p0��%n�m0�|�0}��<9��.p9b�	peڼ3���]�oy������1�f�?@���:s1q�G��@���f3G�� A�=��z'��RP'U�J���n-
W�=���+�ׇl*��EL�x4�F)��Tq~�UZ��+G{v(-�����ݡ���W�Mse�HQ 
&N� �6�@}��hd�p������~��52�>쯗3-_bB0!��q��b���sR���:���zP����r�4�9hB�Hp&��w����#�%�<G�7����I��ip�*�[��B��Μ��N��Zztm�>�
Ԩ��w1�b�����h:\?��0����I��J������t�R�k/�w{qə;���s��9V���/ّh�pb��B/np�\�Ũ�3ז����Xe66t�Y=$}6�_��0K���)�e�Xȓrè�^��k�P�c��s�-�.�k;q��M���_�۳i�w,����dq�8�:+��(ޭl��n��&M�3�H|��r"�?�OuB}�� �b��U�_� wC?Q�u-�J�*���"��F�rw8�pęMT�܋W�}��Qs��~���RU�
.���{�Ri`��$l~�����A)
4n��xR�E=��rX=Ң�_�����z�GE�Ȫo�d@�?Y:�2�t���v�;.���1oޢ�\�S����>�(Njz�oγ�s��<G~b�*so+���΀&wqI�y�M\�aMc�+5���H�N�8���){nڇolz\�+Mx��G��QǶض�У$��&`�3��l�f&,Tv���T/�9 �.iv�&v#7��g�s#���:����~���L�:�%��߲;����-(���%��`����8b�Lj@���u~�%!?$-@�jm� ��	l�O+��G$���\�t�kU��G�Z<���!��z�i�Ǹt<��'b	n�7mV�1���jG⍯hP����ώ���6�cHQô%���3l��z�\Л��(o(�t���T�\$��{���3�د���bE{�2��ne�����t��U�OB1�6Vq��5��C���!1��i��A����؈�6���0�;� �~�	�Ӆ�2Vj��X|��A�l~Q��c���!��j{);�9!9���,�
���,�	��7�'"��@y�ν����f~��i�}��y������#4��v���%� ���Ty��0�mU���J��>'���dKA�է!w"�ߝ���O��k�Ε���z\x�Kϔ�5�x�M"�Ū�]n�M�;-�KB� Ǩ�[���m��c�����+��~���{/-ԧ&�$aq&�M9�E<V���nl�h�1��J���rK=@f2IP{������͸E�3���f,�@�mW�ª�	����5}w�JH�Of�UI0� ~����l3bO��i�2?�����O������JɻK9鷒��$r��JoM�ҭ��L)гNR��ډFmd?8�r�ɹW���3[��������i��R1�IL�1߽t�a8�uG]���@��ן9����/�'���YK/�)d��U�O�-55H'O1s�wmE��7��`�Q�1d�����}Y�|#�!�/zu�W��ڥ�s���z<LX{.7x�ZKQ0�I`&z�:�e���s��� �*S dҏ�AT<�y5lt�����Q��3�P�qNK��_���j�C��vLy0ћ�T/��^X��k��Q��F.�-�|Ս����çG���E2`�t c�L֡�&�0/���S�!���`Yy�U������T5���7=�r7aWUgӲ��QZB6��}��g�� UY�E �=��S0��:o�e�|��>�ڠG����^��E!�Zgm�ȍ����}��Sn�L��0Z�k򎰴�Ό���}4�F��j	Q&E{���ǆ�p�;�[n�p^׍6Ь@�N�Z��}{�����1��Ǉ��#�m��(�H��8&C�g�&;"K�I�PnJ+����*��S�����B��[J�x�In�o��<��zj|�i�C��c0��2�T�]�]ul��c#T��	qf����'MAt�"�5'f�?륱�H=��� [��)��qrl�8�~�}��6�4����塎��d�(�o�5�w ]�G��b�@Ly̙���I5�&�)���.��.��1�ֻ�,:�4���O�3�����ȋ6�Z�l����\]ڝ�J�b��4�un�_6 �'��A8?��n���N�Չ�'w(�z��c������OmS�����vD]-Z�r�k!��f�_�<sC�F	
�k���7��
n8x���gT�ll�1 k�93��u,]�nPx���ǸAC+�:��x���n���vĭ2N��)�&؇H/�[$���}�?e���`7��⣑ׅﮍ�Q@��a�ʻ�(/^�;��*'�G�Hq��5���0��$m��ڭ�U`}��峀#ar3��F��@5*K[4������QO���mw�H�0n�Wp^�����LRr{j�B�ɷ����X	���J�؆����+74X
�����j�9]`m	ގ�ϱ��\^:[�z�ϣ��:	�ި���a�Ж>[�������6����J�D�^�U���}C�m�s: �f;ȣ�x���B����ȗ��Fn���c�v�?ө[ܽ��(���E-��h�!��M�)S��Q��S��f��3�k��
#`Ci�wK8��I{�$=Å$�)�Ԫ��SG�Q~'�RK�%����B,J�1QI�/6�6A5���c����:�����+g��&qn:�ɀ-"����	zߴ�ښ<a#�G0@K��O�Ѥ��������Q_�q�N�'���1�I��l �5ű=�Ȳ>�c�h�\*��G#G���R��-F��3+7"�
ݭX5���s�v�yD}�hޕ_h�{�h��ddqj�ʩ[��G:�<�CD|	��
f=0�J�䖂����^�?.�?�*�,���xJ=�A@�h��e�e�.�nS�D(: �W�d��U���=<'�N����HżcZ�G�=KlV�W�\��A�U�0s�[M$�H��U�dU��g͇�$����#�,��E�#�{�� ����9M�A%K�gf�|8��5K�Կ�?����� u�J���b/����%rC��.w����d+
���O!�9i��hO���9P�y�����>�h�F�Mc-��}-�X؀�-ܤ�h/�~؛I�^);�9�{Pc����;�#K��)���*L
�w���i�7OwI��g�d�y��Vh������^��FYZs�p捠��R�X�"I�Ρ0(�D�*�sz�DS�V7��o�������V'���m�\��7�̲l��[L�Y�o��f v(:��:�i�I���,8a�۰��]���o+1�Ϻ�-��SVd֐;�5� �I�X�=���jŖ��W��&B�����L#��>ÎO z����_6h�����j�y$�����$y�@�]�)�v\h�� '�rzX�a�� �8vG�ι�MG=�kS���p����>o���lbd�8�T,����R�f`��{O�Dޯb�G��(�ȻT�������0p��Zz[_�
Rr%J��U�~M,����n���7��ߊ-�X�v1�HdL�!�z�3P8HT���V���q�.v���4��.B��s��A�!1��y42�����I:=wL_����1#�4��a���Ш�#�G&�G�x
FM+��cB"�;�4Li��N��H�'��
��"�/l�����3��p*����k�i�ڨn������M�i���"Me�f@������k;s�j����m������>di��׮
�Ţ��F����X���!��#�]�[�e�##�=hs��B��v�My4޽/#s@�k�M�$���(���?��Һ�}����G(��������ws�;^}��<���A�b8���d���2����D <m�`*MQɀg"�©%����/�C�1��>_�Ȑ�k�X�3l薙r6ZZ�6*��U �>�N+�$���ɪ!D!B9�5���ߵ2���c1`=Vp�}�����1~�S��Dސ�X=,�ƓSa�=���YJ�^��( &NF���^��ś�� ��kS17!�Q��f��8;~9˓���&i\O� �db�_�a^�An��T��ζ����W���wa4������j�^�����%����U��pV�x1T��be�ОO��N�#e���{�U`#�2r���y��MO�.���L�������/������U w�����S�՜I�ޥM�/:�xva�av�n,�m�=(#��,��w�qF�	����<-����n���v���zlO��W�m�YA�~��[8���(�UQ������"x�M�>s0��6Bt��0�ڹ&,DS�v�F��h�5�W��q�ئx�T��M&s*�Y�}a���שy燧�5SyW�]qB�޺��
��i��REl'|���;�p�Pz�>lO�% x�9(�DT��y�ۿ��#��������_��K�0R"���~�ن����*�GR깁�%*��7@�	g��P�a|���?ieGP�y��u���^AI�M�s٦(oV�|s�U~r�<Ur��Ns.9�z���rz�D�.J��u���m��+`��W;����]EQ� jN�~���ꚾ7ѣ�\@�<����yR��L)�-Ĉ����"�����f��d�;���I�)��ֿD3Q؄��|�1l���ۂk&�:�L�n$�n�R^�K&\��0k0��@ܡ.��HhCV�ŉ���?��
Iѽ㠆+L�+\[��:5̷���#����:N��3�)��+v����C4��+x�h�� ��t5 zt[F;�qK�?��{���|%ܧs��)�گ ��g�����������ͅ�[g�u��B\�t���oJeF}��O��Ҭ��_�^�%S�QwB��HF��$�\B��ul�s��g$;k6��i%\�#4�֣sY@� ����"�j��yp���$��������<�LB�xb&s�f���E���Q,~l���/�C�s��ˋ��4(kLj	-{�B�?"]Q���w�9��gʼ��߫0o����^�^6D���S	��_��:���0Y�JN
�G���~�ܭ�������[�#���7 k�Id�{f��]*g���4]�eQ fP�l�bd� T��]��
�(|�����#3���%�{�/��d{Z�+� ��SL-��|���2����H��C+�j<��8g��[)2Z��Cn�����2�֝R0GyX�68?����N������8�F�ui���	X��X������%
c1�S��-;�t�w�/ oD=(6E"`�᭽�}=(���7{DRG��:Z4�P`Fa�B���I�`'���������g�W��k����㲰�]��CT�V75@53)��ٟ�3^/���)��ʗC#�J�U��jY;:k,�F	9�!��Y��<X{["�����W��j!��Ř��k�R��,n�}M�,�X�ԽD�(��׳�b�8WJ��)=�XF��@+;�Gu��;ޛr��,�U(>�w�nLi����-v˨/У
���0�Dc��
N���嚆U[�GU��	F�e`&sbE4�d��h��5��L��� v������!~�7X:W]yA-*Q ��Wz�9�X#h	K(�;��7a���FK��-r=cꌿ?Xo�5����m�5&*��z,=s��͐��
���`�r�5҇�����Z�'|�7����&���h��x��5��LSZ&��Q�^N᠂$ҭ�B;'�������&��4�$).mB2�n�P�E@�.�Q�	 VUa��A�� �Kv��I����<�Y'�|��o"��9Q���l��� �٥�`�C1bn���1BFd..�BIa�D�Ы��\��^Ş&>�v��c5aߞ�^�*��6w?lm 5`�O�=%�΂QF��jI���Z�[&�[s��1��t� n��R��u�m���˄]�ތ� I�7$�"V���Pr�0�&��k;�z��r;=����T�!���0%��!�}E�]�k��]R�yE!<~U6��æ[iD٢�^yG4�|SH�%NE�^�)t�mP��:G�������S�ĩ]_�9�F+��}��Vڏ���Z��y�o�/��^X�]���W۔�<�]���_w�� �}�v#v_��n�u���L��<�觝�t���cN�<��bXM�DܛIׂF]�NjD]�c��z����Q2��_��5nN��|�D�;p�^��Q�Ð	������ :�$���F��kA��_�Ju�k��ޑ�"�*}��ֵ�xT|IΊ�R�j��H��l5�;М�f����0��|��W�k��on���F�S;��X!-����Z�yF��m�tv���2Ӧ��,מaBo�>�:A�OQ�To�Ƥ2�Sѫ��2dVj�|;��[-�oyH\�k�(<�-��� �I� (���Ak��W�I�I���~���5����%�2a%���r~�w�bX����Ob�~�]~�`la�Ez��lyG�U�VR����׭Q�e�H_�����y.��M�L������bK�Q�YZ '�!������tQ����бs��<:z8ꆸjTP�q1v	�����֎(�s�/�*FEI�w���5,�� �ž�}#��ؖ��s�ѷM�'�IEG�qaK���0m'	���;A}�+�[����^!�K 4`���h⇙�YǄ���zb
+^����U�h�C.ʩ�	b�B�:s-�DuÒ�����?fs��,��<�Fc�8joq���t)�͵U�E�Z����ݣ	>Lִ�?�@γM�����+�u�*�<�C%~V�,���rkza�`��]��۲��l<����g��Kz=���	�T]���$�2����
$�$��Rgm*�,�{����ږ��]�G�Hn
x���r��Bӿo�ic�����y��\(p�,�gcc
���G��Ɲy��@�����Ǜ7hj��b�u���[���`8\˺��h�V���]r�@�Kx�h=�r��:6dM~��Ó���>���J��o��1��q����!�a���]���Yw�E�`�d	VH����&�+�l��w��C������CT�N7����SnWϸG��t,�_pwǑ>&^jԻ"�vA]@XO���C�N5C����"�ɀK�θ2�u��:�)��~�?&m��� Tt�����S0�L��E*��7ά��F:��.nHDB�7n��&�.<eHUC�����ħ�=l�~�J,���dT�⁚�H�mQk��R�f;8[�|�������V&xI�c���Y�7�U���t=pz�)@{�]ľ�Ho&�H�"Y��9x3���P';��ǯ�������x����b��L����e~3�Y>[�����b��Q���`B���w�@T����C��~p���*���D��D�,t�`���a��l�Q>|���@�"����m�^�p�6�)�F�{�{��0�O�����=����?-`�jf�����,���^���v��6�w<od����^�' ��	YZ�o�h^1�����iȚ��o�l)'��(���zf.,c��1���:L"ճ�ra+Í�/�8y�]�[��i7,�Jݟ2j���@&{�&���_����ڙ$B��$��@���W5�/ӟ�oG��#�sk}YtO~�z9*5X^���t"�����ΙO��OY���sM��ؾ ���H?�w���P6��i��:��a"��\p �%v+y�wP_��dٍj��9��N�[44�0�U�[��ԅ�Z�N����f�Ÿ�Ot�f=�eA��o�a��2�.˫�����Q$'�;^Lo����0��
�?(���.[�S`N#�Ϸw��	k�ӝ��{�z��Պn� rnԵ`��� =��
#�&�
��7lߋ�e`�}h��6�-��;����d�fj��I���̵��{<Z��yE΢��R/C{F3�C��3,�DD>�����Z�3m+<�8a�R�1��P����5"p6LFfԆYB1�9��� U�T�����n�o�9p�|�Ay��$��U��P�9��7YF"�u��2u�����6��D�uE/-��ה��ɵ��lJ�I� u��j�zQ���j��K2}!K�e=:['��ĜkG�7W��J�3��1\	������e"��4��l�8����̡;z�k��.r���!{@|��'�˴
:��4��٥�ɼ6��e�^;0�ךg��#,0� Bl����W8i�ñ�7�
ZhA���:�H�ֿӵ�
0jD�qB�B�ǵ����7P��ށ�(-L`�r��q9dᡎ�B�s-���:�*DĳT98.�X]�������� ��:~
�܆on�u<�����4*%�u;�y�ǌ�r��y�I��ڿ����c%(f����\���ޖ7��u��{�s��a=9w�W�|)o�Z1i�Ď���u��ם1(u���?��$��(�Ph_�T~i7�4��P�C��:k�D��E��r��T�1�h�.�:�����|�����ʐ�O�x>�������7�ώM�,���#�/ȣ����K<V��ף����#_6�û�W:.}���8�߭�YGH��EQ�9�++RCG2(T���,o�h0��܂�:q����
C|��0r�t_����StJ�U�VL:JQ}���c��mO%��(q��]�"�%l��ѭ.l4���ts��@k:L�QɊ��)8G�-T3*"mԧjWI��ڤ�!1�fW�.�-\��I�҇��gJy`�8���u�_��n:����)�v�T��m��8G9����[�Bh�.S[��;�Q�����5X����+̩��8�c�j��6AH�jAs:k_�et��-}laˉ���y.��`>`a1صq��-x�=Nw٤u}�l�7����ܝg��3�0��bt�@�g���*b�cO�F�R�s
r�,�v����^����@~�i�.��m�nE�/�KGX���GN�����F����!�+I��.���w{v"�Ӄn��y���d�̴�Pߠ���gu�Yv�y��Lq���d�I�O!!U��L��� ߾�`�63���PT�=Du���8K��=��^/1��g �`���c)�T:�Vm�fe��q��v��C*qU^����J��i���f;���Nj$����|˙b��
�*{�^����z]p�,�9�7��%q���[���s4)�������gq,!ww���/^s�5:Dd0�j7�?�L|+��"GѦ-��`w�5����-�S,�C��A)R�,aK"�grh���|�eÞbʶl�c"�_ܗ��-�Y��oA��x�N�+	�W��#�g;�(*7�u�ϕ@�=���-�Z�S&'W�����eQ+�*���^E�w5�|a�� ����O����־��Z��&m� �٨
��ʪ���D�~
�農��jJ�>�T�Iwd�@2Ǆ_�v^�e4�p� ��T�i�*�� ��;�4m׍�4���5}���`�WM4��W�kT
'��x�uX�/0�f�E�%����t�1�*f�b襌^�YȄ�b݇������ ���S�{���+9:��vZB�By}}�X	�v��S�#v��w���v����#a/Yη3d��:�"���F9���x�ow���٥-��"Pٝ%��'t8�5�}Y�~i�K�C��gc�<U/��T�Xp "]��l՛z+�Ռ$v�Z�c�>oՓQ-Xd�Ȋ���{�b;�L�#���?�ޓ/��� 燥�����Y�b�[�.�7D&�Ͽ�
�����!�|��e��I�L���zmBDg�U�ȅ�^#$,Sj��	���� G&��R]��9\I#� �@R/�L��o����7�dщ��Tz.�p�z_�:$ނێ`�����$.	)��_�-��0.T�3��S�Qe���:ֺ�,�%f(ZYDؗc�� L��^6>�s#��R�H�U=W����~v��'�}��B���}wOFt�b/s�a퉑 ��̄@��b1)Bk�St�MEL�'ZB�c�9#^iw�=��������M���XQX[�dSF�ˤg4�p��f�)�*.�HA�6!Ǔ��[9�ʜ˲A�s�T͸��R��%�f̆]Uu٬8-��;kD�է�.�w�Eg�����:gC��Ȣ��N��)��晵���۬*�f����$��D���Vo�8bY�q�b��6�H����B�BOG�W[T���Jxm
��a��(�/��պ!�퓁�u��M=Q�P�f���u� 6�c<g����aa��@��Ջ�J�3~�m��t�㩭Glϴ;4uk���+\@ޤ�l
R�!����+9J)ꝃi��2�F�ڱ���������+��tC���ɽQ��n��[qCАe���|z��X�����U�G� ѧJ�e��B(Y�F�����-�����+�7D>�ob�$.���:�F�y��2ga@�w���jd�O��\J�Bmf�Lr	�X��6ò�,U�T���<ʨҘ�2�v�.$�)������ 
w��^mE6W�~�93����tc�;�$
ϏO���X��� G���2ƶIh�A|���m%�-Pƽ����L�\���@a	%Q>���x�HR�U��Էt�9S�C��>�X������B����j���]'e�٨�!Yͼ���x�ds>_Q�[���hÝ'M�林L�r�px�*PP:p���Ӹ���jLw�r��f�ư�n���c���m�eoI\V_y��H?�ګ�{�-�Q�E:�K�6z�c��qiPPxz �"s��N-�����M��	��(��pw�����'T	!�I��}�@҉l##)��3�S�+�/�����i'q@X�Le�w��2��{}��T̖Pr%?��6���ė1��Y`�|�Y2��X-2j�����1�nvl܉DUa�����ߎ�֛ԢwB�0�tQ�'io%@�w� ��S�E�#l�Y�^�& W\vA7NkdH*�H�f�����3��y�����v�Jnf�v-�1�e���%?��bj�"g��rq������X8�xl��BC��u$�-���/E&y��p�N����nxlF�厰���%�9P?�YSٗ`2)+g�!�G���})�I��/��L����	�R:���'f��m:�Eʜ������؏Η/�b�S7!��nU�~il��:�)�y���|>�{�������,��$��\d
-N_k�(:g���%C�3:VgN`̩����Y!�#$�L�~p��4�� �F�/���z}9�3�����F&�%���y��S�yTϮe���ֿ��M��n+��ԚAG��,��=X镱�[�?�ϱS��uռ2�;�:�(�oE��~lHP��������������~�_�:A��|j)z��D�,3W���2�2).7WI�N�?&�01?z�[�MD��]x,�`��8���
j�C�#}z��$NH/�`����p!�j,x�m�MB��'�J����@��7+TMÊ�r�ק݇��siv�</��)s�z���`(O�s��7쾏SA�ݏ�N�����'��y�oI��3\ʗ�s�����%�6�{@�$.rQ>vN�����~�JF�������� ��sB�et�ly���R0Z�<�f�^Ο���j��xB4���S;�{�:��X�Ix�U�?��?�Ŵ&��%ٕ��=س��r7�S��/��Jk���'l/D�T�C��8�E�1�,�����	�oqs]��nE���.�%�<�
�w�3��d��ݟ��$	+ ��f�4��a�N0Z�ar��\.V.~Tfڤ���>�潕�4��cΛ���a=޿���]�ϋ[�Q��f'��qT�(B�:6��{(��Fҿ��j��V�4� ��"^MmZfى�<��e�"�����	�37e��NK��/<s�Ե{>hY|/Z6�˖�je�Gd1v����}_nȌ��*&���۞���~A�{^`<�HT���0M�?p��0nr�R�0��샦Z �\�j��D�����<WQ�u���T��?�U��u�>��Qդ(�o�e���?
�Kתo�y �%���<E���W)�D�+R�/�6l�S^$١���2u�������F����O^E���rp��݄������BX`%h�X�츮���~=4�ȳ�̀�HhLTC.�z��Җqʫf���k2]=�9f��){�f~Y�5�|���kSY�b6��Q���K8��ަ�)���)"G�!��_)��a�,�b���Ųj(i�e?�~<�{5=OE�LB��4 ����7���ޘ�/����P@��) (
�1P/u�D`�醸\N't�yQ6F ��wC�\
�/��}_�����|�o�1*i0�,ܩ'�2#ؗ�K��/��@gD���	��iyV�boH���j�~���àM7c}$,���i{#@k<�o����k�&�]��] X;A@`�b�{�	\@h:��+��oQ,.Zl=vڞ��p��������>5a�(��'�w���x�	� ����<Tw���B��ъ���вnS�Y,��Y3l�\��&(�	��fD��v��0�������OB�L��7���C�T�)PX�̑���*҇����Q����d�B�g��e％��R��r�79���`�������b
*���)�y���J󋛂L7[7��5!�s�g�q?��*��1V
���~����x+��ZC^�-�đ.kڄ����f�v䑠p�Ӱm{Ov/�X�W�w�6���5�g��a��0a$�L�陻# �ꞗm�]��
Y����j;?�K ieTR+h�û�;d��@ܫ2+�)�ٞj�A(��,��5��l�����h�g�3 }mѲ�"�}��iSs1�⬺Q��� ��Df+u
�Z�[4�5�&�A���7_~ ~q�(`P���$E�8�~y�����U^�߀��¹,�L�a�9�%?��i�s:y�kj�
�6�B���I`����Y5!����fڅ��dg��W�s\����q�Z=$�E�%�0�㩷k�����QT/�k#Ŧ����V�F �QoAa(g#�e*C��ŜD[���~��.M5L[r�Z���VZ9�2��!�5�?�'��1�g�Rc�*��d~�,���o���)5E�1�tfcAy����uz�0;7O�l���3L��Ņa(�7_���z�o�U!̺�i��n�J~���)��q9\oe�`J=�ec�'"]��5�x�*(�Vo��y.;����r��j��yn
��ߒ���8Ϋ�@���$�wWMn�O�a]<:2�zǃ��������g` �da�^+$f:��.�+�c���E���i�p�j��بW�$�`c)J�z����3���.�t��RǬ�g d��vޞ���s�1��hk�Sp��\~�Eѹ��df��	��"b���x�b;���3� �	&�1@�mBaR�%��+k�u�j�Qt�N�"�"� �Y�A���?YD�yr�~��*U�z�����vիIj̜���)�B�����h.�(��q_��h�GݜQ�I�%C�)�=�K��[K�_�Q�]xGtm}�%<'ށ�ƞs{	�UN
C��e6Yq�Øh����ݟ�,�W1G^�l�O��O��q#����Ih��6�v�V?:2�����3* �,�.��"H}�u}���Hܔ���){�<�Ev����'��&�IB��u�v�#E^���2l��"*c��<ksZ����ޓ8T�@��!7�� �b����`�+EL�-SI$�i-��wf��o��?��kj�p��O���ijk�}>��
���_� ������!ץ�ǋ2m���ݷX*ʅ�v�y�J����V��>�U�m\�#vf�D�\A!���}�i<����ڢZ�Z@�gF�16+8��C����Ԙ�P/�$Y�ԑ��i~�!�}�F\�s_�
ZR-+aἽh�\nV�w4��( ܴ���e�A"<����AEZ�_���/u�P_uy�.�t�֔�8@/�^ϵ}�g| �
|aجuwu�2]b�ݔf�nȺ�ߪ��N�ݟ;��~/�����@�+zP'��eR��p�p4D�R�G�B�b;���K���d���3��Ϯ̏���S��~�>�}6���  �Z��ξS@g�;t�J.�b{z�)0ӑA��0jd�j�5�\�=j�����DN�E�
u� �6f��\�.S�uknS]��Yl��FL��l2E�\�,���U�~dwU��ޠ���Rw��a�#j����V}a��l:w���;fMi/'E�c�!a�J�x��l)��Ų\L�A"d�&��+����}��9ȹg���E���H���i�����|h�D`'�<�W(H�󠔐٘� o �cn�4�� u���SĐ��9U�,��9����pl�QR$}w@�`��+B��$�5��L�W��x"q]�R�%�/q��������
��ⷊҳY�tK��0ȴ|?EV��˧7����HYTr	�B�o��:��~��~�W�Y_Θ�̗+Q�QҞ�Xi��a��n�TŲ�^�Rz���HY(�u<���'��a[�1��=<Ŷ&T��8�j����.�ro<���!N`�!x�h��@�LW'B�\�Ű��b0s2ܝ���|�].�u������^5X����1Y�8P@sͧ�8RYz >?���%,��*�L_�K?�K20�B2����t��rڿ1$qQm�0;��) f�K.��4�nC��L'��
nr�S]�����'����_ζ�2�SЅ��g�/{1�)�>.!���05�>���*�EEa���)ym�ݔ�÷SL�\b��(#�����ਭh|��D�ǜWmU�Yh{�\�@����Γ��_��0�o'(�AvDT1�섑�Zr��������3���g�6P�ܤ=�J���
@&�����@�,'w�Ǳ	���=�@-�rڄ���m��-5,T3�B0���H��~��T�rY.�td�6	���)#|C�q6���_���|�ۮ�f{�w�GP��(�B�7�L�I~/��3ʲ�o�����1��b+,NZ���L�"{����xu��ވ+>DCʠ�D΍5�W>���̽�.�A��'LuE�
�WS�!�v�Z��ݼ�FB���� I�};j��;�9k2�zӌ�^�*�(���T�|��^i�)�{k�.��w�MW�f� ��HnX]L�F99"�+¶mϘ��@1~3�������)d����~��R*_�\����NY��R���}k 3�����!c`�r���������Æ*�m�n�3ίPү�j`|�YJ��B?,��>��9�j
���.a
�AUD�D��/�#��"���@�������(�}��q\Y��h�}[M�+
��^���֫�F0i�;m�i�ܕ��@����I���m����1t
f�"}�|_i��ce�m�݇��{�3�v"�>�������B�F�ox]��W1��,�Nw��Rx��;2*$�b�R5P�1�n��Y$0[���TvU���9q�ٷ�W����Lp-(�'���=��T�8cTB:5Kl��)�uf�B��������2DS�,.���S7�E��A*�W1�FM���d�P^��,�#��}��e��@(��}���}Ǯ,�27܋���%�
����,��&ھ��p-Ҹ�\L�'��u��'���o_d/Xľ��$�oiᠰ�
q-dG���8S�d/{��� 59l��
�D����k�r-Q?��� M(eT|�S���D_�3�i�Q(�p�~n�J����g�'�m�n�rM�	��Z��VcW���ecA?�"�9�Y�8t@/Ry��q�u%����A�&q�s�*@��i��(,ٞ
g�þ`�wQ�=�\Isь�2*Xg
R��y����y'�cO�9�3a� �Ao+��E���pdV�sJ�Z½��S�������}���}
��P�;=���t�FqU1��Xq�b�#p����32$`m񽟎s0K���� ��-(8x���{�t��FnC��q�P>"�ZS��A���5椘����6�����	�����*i	@�q�)��&�u�drn�|u�!��ܷ+"�T� 
տ|e'�   @���6��T5��'�[�ݭ�;��m[T���Dg�.��,�Ts����,QS�Ж>?�-�Jh6��u�\�UG�./h"��q�U����<��C93.�����i[��f�"��b�D���a����m�����.�'L��M�WW��Rb~y1��U���D^]�s�b�+���R��xV|̻��M�lT�N��6�*��K$�5�C�T=�꜊�%�����oy�-Rv��ʻ@�^]����͑��&�p�Pd�����ȮR=�	r��ː;��C�`�ru������g1I<�N����Ҕ����ڡ_4[[���Q�iZր�D|F����	Wb��~;�\!��F*SkR"�95�E|7:�#X�?$0#kP��^��y~)�~�S�����',��JZ���ЬJ�	Z���A^Z��e�" ΐ\S�-h`����U6�W�u�'R}�AK��O໛J+_����8��ߊp/��
�y�\� �;��4A�ȩE����!��W�A�.�fpRX�>���b�r�ߠ829��}�K��d~Z�_�C���`�B��h+��^t1ٰA��ҝ�9o�g}�~֗eD�C|JA�x��P9@9��=ȹ����x)ɸ:R;���¦
C$�);�ؤCz*�t��ā�m�ȯ����"���:�J�K����O�~CP3q`3�w�N�qdq����j��C0����Eep�~�Dx5�EYB?]�,G0��q2G��S
���e/���۠��|6>G.�Cp��u#�0����ʿ+YX$�����J�O\���Whl��������Ѥ��	{-+)GE9�2ӕ~�<���2��IgXa}��6̣'���)�g�&��'W5x֣_�ɶ�<lcƵ����(5؞����T=_���n��̋�f��&�+��5sf���M��X��8��O1��Pԝ-B�$��߷:�=(D��o���o��TF�{���h��L��1uZW��m�\����6�~��c��l?�H�v�	�^�2��߿�H�>��#��V�Gl�׎�X�5�~7�S+Eտ0� f�\;�a���WP��֛CEU �[u����j�U�|�$N�{�+%��G���/�łR��<���>0P�`���!��}ݤ}"~l��]Y��(�@�_����ʚa�~����! ��w����u_��MW �f����'��%@0�NU�YW̔�DA������w���ĚG'��ʭi�
e;B�L%����<]��-4.��[�J��;۳̸5& �fS�(�`S%��n��!kͥ���9�r�1p��#�����NLQ���ֿD��Z�%���MOd�'`x��	A(@�:�[2�k-�Fc��O���L�f�M<�f&I�m�Pa��M4}@�"�
�7A�V����{)����p����{OP���Im��gh�	V�|aM��Ü�Ԅ72���5�!Q5����svP��`�)BI�����7����`���_^�^����a�͆�x:ۜ��^��1SQ��v,H��8�~�h�{/����UUv7�Q=��0:$.�Rġ�ͰU���Uy|��4��w�x��{~���B�a4� <k���D�(3�uOm��9~=2��8[����hj��C����� ��8;�ćctu�Aa��8�x'��n����!���=#�
��cI���R��7"=�TJ��Ľ%5 ��&A�Ƀ�J�	$�wg"�Pj�V�:PLF��`�S���U��d�A_�6��?�0���+���b���x׋�h�EǼ�-Ec��?����f�&�ن��wp������ri`߬�