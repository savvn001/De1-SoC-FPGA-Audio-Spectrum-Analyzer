��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	G&7~�?2[@�x���"��y�l������>:�S�����ׁN��)%���s�VK�� � >�w��9����y�w(/�O0!J�ZQ�%5PRr,8mҩ$/��ܵ���UB̲,R��	�}��g�n���y��x{�D��O���b���*(�^C�sN���[�-G��� ��C��ֻ.�Si}�_�,Sw�(�(n$��'Q�ҍ �}�[���;7�)	�.ZH�<��6^��hɉ����M[����5���:m�t̍;^M\%TH:@F�/bkO�U�h����,���_�ս)��:��z�{�+:V�2E:��?��@y�@����`���`��4rp��6|��5�D]=�h(��!��������Ff�� �f��ʃH��j�I���@�r\e��.^�X+��h�)̿X��u���NJX�P{�n��%�5iO�Ss��m��b�O{�}AS��h�#�g�M��P�y��YB�Ϧ��/��b�������"�]���Q����K���b��(��Vg������]�&�y;+SPV�E,�g3iB�>�{_�m,Ci	J!|�%�A�
P��=���G�{�	�c#�(
�-,F���+BpZ�n?՘�jw�|C͸���³u1����Q̕�r��F[�C14ө������I���Kn%׬���Hw��<묱@�{K�x�QL5�/1F��-���",v��=�|5!�k��R�ᅥ��-X�;���X�!��>�	��_�`���B�yS�*={�,�3T�B{�+�	�a[�r�p�O�t�qǁw�e��ܱ��_�ԃo��2�:��1"YtTG����O��n���Y��_3��^��L�[ǔ$Ȓg�wP�;e `.<�����j˕�2��d�XY^���ۣ<ü�AN��fmI<N<�t��|� @�n��gz�%~r}�?�9�	 iA\�(X�S�f��n���v�p��j�'MgXx
���af�~�����2 ��}�.����8
i��q���A�Ȭ91bg��9'�l���{im��Kf�$�m�c2���2�i�b�Z�b��.�%�l�`l�]�*&q���J�Q���"%��*�ha9��xd^Y:q��ם���ju�{z�����St���q���+�������U�����4������0u:IT�*>�M�?!����0<i�eL6��y���@����A����00c��*�-R��>R$f49��{W��_Y͈�4�� �j??`ڢ|�&��K~J�b�.ȯ�
�L3�0	�����j0����}�#Ԗ^{[�`{�`��Z�S��5�-o�U����A�%2'�!��Ε�φew�?U�:�绔'ޣ�s��N|q�1���g�]Ǎ�˒A�Nm�G�W���C�,�=�#�ЮE�+Z|&��x�;�K~0�W�K�A�1�C,lu�9�D2Ͽ����]ǌ}3�DqϬ	������޼"�����w�����9���xd\��� ���9��p�ˢ��`]��!�`��PL�*'>��}!�Fc��C�ے��L6ɣ����J����H7B4I�y�6hA���)�[˴�E�Pfઞ�B-[��EPj,��Z���7t��C��-n�<��\?�:#��P?T%+�X���w�Z6Ej,ba:H�Z��sh�t��Fа�'@-��w�*���v��f���a
��B��U�%[�.+27y0��{�H��s_��C���:f�s��V�D �a��J�}3��3h�ZDqn!�9�Kk8��O����K(�y�`������c�ڍV���pZ�a�_~�ՒE��7໐�|z�έ���Ў��L�io,yE��lVӐl+xd{�R
���j�p�p���e*W#��@�I	B`	Rh�F���X}�s��o.9�5�+���d�٫	,�Zs�r��Ќ/m>��>}c�����E�Q e�KPsI@����8���G ��v�U���5�=A�c�B�L��n~��r����()���4b<��d�B���c��[a꫗���|�3UAR���?X�M�\�O�����3��u��$.׼Sۿ�@6�}�TU��ܫh[;�%��Y��$̔ڍ>�9�
�^��K��buQS�߭Ҹ��_� �ӟ��`��&A�.�x�yz�X�)6q�����G,ŏ9֥O6=�y^�h^�!Y+����r�����p�:���J�q��[o�%I�y�BX3l�?������bƮ�w�jܛ�(�Vf3V�JFl`	�T���X�`؅�)�{ןa�Vĕ}���\�о��}�I�F��� �Q��vf�o'q�O�;�A.�u��@E�_X�n��P!2���\��Qԃ�LC���y��%�u��9�>v�.b�㧹"D맄�Nt׮�汖�b�w������`:f��F�^(5�����K��D|I��|��R�[a��I��-2Z�s���x���}6=�qM>��RDO� k8�qsz�?���c7O�F�^~ᏮȘ$������>}7崪4���������B�Z��t�[Ȼ �W=�6sn�Io;�� ���!�²~��η{�3D{���F��6	�Vÿ��0ԝj*GIM����A�Lo5�8)^�ɶ�T�,����k����\6^2�p���iƆ�V�1b�J5�7Z2�h������s�{��"Z>�T�H���G��S�$�l(T5�����ʂ�CM�`U�z�"�p�nzS���i#Xz����/��6.̺�/�u���U�[4r��<�v���]�=XH�|�{��?"p7��e�g���vt�����:�a'C�걁����aA.�+ؖ��CTHw��#�.��gL�*.\�d��O.��ಧ�B�g"�M�l�Sۧ����1�G���\4�ٵC^[��+T��N�ؐߡp4�	X�/�Lv�������m��eZܗR|��'F��Ÿ���������h�\~����?;���avF�ך���D�*9j\������J��]f���on}A�c�'ʣ��{zW6�i|�����9u�_6(v-�8�mMF�l�ۼx�
2C*��so�Dӎxl_y��P�u� �%���Hp
�ʝ��s�]�g4�<,N%��1)�.{�}V�;ET{!�'�wZڸ�d'f����_�]�3TЃ�g�ÍjH3�;!��N+b/oDO���ظQ'lJRK����L�p�(lʅ߰c����K �c�5��0�%����[4� �­g�R����0�z�Ro�&���8w%���B	/�ܟ���v���?^C�2/kG�TU�<򨊚X�b#��R�-��B%���#�¤���J��H���4�]ID7~?});��)��cYt̕�~��������#��	�'X���iuߟwK�ٸUV�ŘH!QI�Q����j�+~�mC+���0�m>��%єn��<z�R¡�)Yv9��.��B�y=L4wXj>��4P�?˲����j��|�'��3��|���$�	Xd}��@��U���<�����wߊ�h�;+X��맕'_�A�["���#��;����ɼ[B���l������{�[;z�JL���]�ߗ��c��G��J���ǧ�G���2��	B�f�e�����O���D�P�W�)����[���As����Ǧ��v��o��@�<v�k�>!���Nhg8�(�����Փ�Id,�i,�����d7���<���X�{�BH��@��"�7^��J�1�b9�d������[3*)�K���n,�,�$V�w�����SᄼA%����!�l�&����>���7�&grRƮ��2�n>9Y�B@Dr��f��=�{"�|��NNN���uo^L3��͹ô�����$-����2�#;���0� 0 ~�_��K!��pIy%)�:c�c�V�ȳ�y�������l��Y�"���Up$*�Ju��j[<���	�t'��1��	9��˅��Ihj�T�����z�x{#~툽,���#�Q(�L�X�,��3_w%����q7�LN]���%�iK�U�~W�[��&�"lkUdmo\%��?+F���S~�5�B\>�B$_P�؟���i-�����3u�&~�amΟMa���Y���,[/@�� �IϺ5�
�A���X9��Hv��@��	{����U�0��̞܋-��wl��Dg-�o{�e��l�	�A��K/Km=�i����o �����0����np�7Z[�i5�:�j��6H��vYvX0:@(t�
MM�H8���E�y��U���O��P��e�7?���=N����\rId��+��� �=9\�؄�܆A�ʎ˹���_y�K�tu�lk%�?����걒G�`Ż��B��޼�픯��t�<:}|��e��)��d�pR���ޭ�[c��Ի����"�>�F�1~���>�uHkX'K/@�O�3�>;��r���l�o@����pC�?�#�/Z��s'�Oރ)���I��$}f���pF&2	��`����M��w��K��S�Mǋl��|�tچ� U����\�)f'y:z�ϙt�ج��(_����n��i/����3�ĺE_m���U�+R!�n�xC�$�o�s�'Lăy~����ɉ�5b��A�+t^q��lr}uħ#�߉jv�@6�K�Op�L��w(W�F��'�	�S�&���Yy}]��-�D�P%�X���	#��Wz���T=Y�vwad� fԭY9B�f
���?_�FuK�]^� \}�b\Q9e��ۓՎć: _����5���bnl@��7<\���"�Q]�9:��6x�T�m��2�@ �wW1U!�A���y�J���L�Z�����G������/W��t��:,^΃� J;�V�:��pFGI�ڄCN���k_߽-]��q�6����g-h��}*"J6�f�oKlg��������,Y}g�RW��_�<?6,�T��Z�!�kxB&�6l�,{��G��,x�|��p��;�x�;
��� @�'�Br����f�m,��Ny���|���f�>{�X���� -t?Kf�M&��;-ܸ�.��w�;Z�֜kѮ���&UȈ�����p	�zX�Lfi��f�L�%���3{�էaU�-�v�ն�x�lj�M��7Z�`ϖ�'Y?c|�xŨ����c����ψ
K>*.����vE�f��L�����{��`�"�|��Q���~����SC�ܩ��ר�6���(c �#~���qԁ�Z+3�Z@3��S���0��o�!� �l+���hT�h^���.g5�GxM��F[gL���Sr)�e)�%^}��Z2�W|�=����%�SZ�׶��"yS���'��]9���ARX�'�x����I�C�J!4[ց-2��z$,�hض���4�*�����m5���3,��e�f��o>�8���J���:0���e�a�x����ܣĩy}Q�$�?��~��I9Q5�))�KO ����9�7�;�t��-Dd����7���n������Z��(q���w�C˘>�G�Z�O��X��~hy��<�~��ٶմߡ��N�o��	��&F�-�d�Fl��hvW���ژ��������Z,����cG���:,��e^3ߣy=&�_p3�W���_=h{m��`7��aXI�Yz;p��y�	�������;�ݍP������}70�-U��ET����ː�_Dй,%2͕��w����ק��?अ���HhQ[��ғeֿ������D0#y��ZpQ��	Dm�3�o>���4a�����]�97�f�RZ����50�&k�/kY�W��r`��׋y�ȕ}��Z6���Z�0�e'�0��gf������zɻ�ܖ������/����5,����l��7'RPXG\�٥O������HU��������y�\�hjp�Ev(�X�qsH�n�R�V�e/Qo09���,���	���_��6�v�}���jp6G�����`���GW \��uvwŒ\�-�g�3����t�Tl\��]��K�MP!)�s +6~�\,��EQ<�ş��@܁�^i���4yV�酬<n-x{�,����מ��d�x�.<2��?��0X[<x���� }|�3����A�:������i��I%%o�<ErQZ7a�c��t�b#��'�3�G�j�*�q�/~�U��=���U�T�Z�0�IlA����H���fn��G)�R
�� w4Ճ_��E��2g�Ri�ظ��̯�ȧ辒�O�d�;S�h���ջ�o��`]00���@��^���T[q�튵���T��Y0����6���; �9�as�m|�
$i�k��=M�,�!_���J�R�'��Z�8�c���x�:�*���G3v\׶�� NmMK�?�G��jU�%�H�Z�F9�
�Ma0N-0D�ČĜ/,��CC}������>����,Yeo�=X�_�,�r�>�O�Eg�g��X�1�t(���PŔ��[U]]����lV{ZV{���V�����?�ٕ��	b�~%���R�Cc�)���F�&R�l*ܶ(,_N�z\�a�<s�]�7��װ��-����odW����'�U�c�c��l�.Ϛs$��� �8��&���x����KxlA�t��]�7 g�夠�Pc�L��`y#��RM�n7�in@����=�