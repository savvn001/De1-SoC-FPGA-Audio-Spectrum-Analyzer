��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	���)R"�=�"6FH����
���v�;?��V���G������nk�U��ۓ/����e�3F�K�}����'��O`޸��؋���e�n�P�.`��������~�ޒ�o���P�Y���.W����L��+����+��Qq��:!�:} ℾ�޵�� �"��4�m6�u$�5������n��=�32[ij)�=i�w�s�T��QNĽT��ZSrա���ܿo����>8F�/�Ez�6_d5�#t1)5��cl'qX��i��3��nb{���p���U{�[A�YUq��ϋ�j�E��f��3#`��'��rԺڶ3F��u���'�,[�B�S�E�V&�j��?+sX�W$ů�������@�c��^/�5횈��8V4��ad��(���e�/����9TXP�[�<x�G��Ѓ%މ�_�@�M�%_�e�>�	�	-�&ل����FD�/(JQ�Ё���s睄�ƺ�J�|Qk�[��Ǜ�6}�H���6�	��VQ����+��a͸�R�z���ݧ��t�n�QL�*�@ʇ�_��F�G���^��*x����>Xv7���g������Zbb���D��Ɗ�<��T����y.Y�|��o`�w�[L Kz6Т�)��þt�z�-�2M��`E��w�a]�V�;NF��[����˺P��P [H�;t�U�Vh���g"���I��[Ώ~�u� �����<��@
��P��o4�a���d�;�Ƣǈj"�ats��l[G��r6Y�+�<~C��G`���|+�\w�y�@��Tsړ����.B%񱲵uew��T�;<a�nX����f�J3�ɼ��@N�<�T�:��}<����;~�D���m���n�S�,8�鲨��������[���ύE6��2O�;���(m��J;&�b���0ד*�����}��I@#��a\PHsv �8%k�ٍ��URs�X~�!+���tl�L�Z��ܑP�K��؆ׂ���^��b�,��3��8;ҽf=1�%�ε-���̄$��T:}��}m]�U�[Qn`���g��B�8<���A���YoP#$�w�oM��`樤�������/�V�{��Ѥ�L'S��3s���kɈ���A@Vk<:c�Fx$b�"Y`�vf4�]N�(~D�l������Lǈ%i�{��j)�U+�ے��έi1���+��}�:T������E�ߞ�៯j�Z��gQ�0�d{m���BO����T1���v�\
G�`=?R4�O#�	����}�(bn��i���:��r�4�!�R�9�P/�Ȣ!��i�k�����.W�4����Z,ŗ��[Jہ���ɞ����A�T..�Bf+���Ft��;��ð��½P�7��*�5�u���{6\��"_��N5$M�Â��]"�:��"%O0�:�}��^�cJ-}1��i�%�ЋN*p��?򖻶S`����ap������:��v�_�2�����@Ft�rE�B�la	Z� )~���]�J-~4آ�8�иW�׏ө��"k<��
�_��m��6���؟A	C.�<u��	�B�����*�]�:�ܯ/������]�H�{�1�@$;Gʚ�]k�7<�	T�Qy�B���5g�?L�2��;d� "{��ܰl��5�֠�K���Kך_��RR��|��::'�,����vgV:�>��b�L;����c���P�C�����+D����Jʥ��������0�]�<�V���碶'@�{�T���p:�]GH�]'ߒ}�iUiD3���2�O�TO�OH�P�����S�6n���l��J?A2II��=В���-Z[Q��fNQ�u����e��b5E��F�SA��!wH��emq���ch�¾?k^�`\k��xZ=J8��:����@��n���?�S�hϐ<:�aU��`�\iu�����V&�d��@��ps�|��N�X]*��Y�$�>[G'���}�ͱ�-�A8P�T'�J�pV
�*K��n#T��+�i��±�`��@9%.l�~����R:�?y-+NݓW���y`��r��Β����1FK� #��9Rƥ.^�R�6ɀ$�c�H���x��?jz/�̱��R5��iH�]����5��ʍG�w���2G�\k:FjW<E�l�cG܃�41���(�O��x�1M����q_����Vf�9�+�y>��M�)q-��jq%<�$N��8���
z)a๿�����Wu@M
���Wa�Ol�&��
�X��X'jq뻨�{�`S�<�h:'�P!dl�����vh��Ы*�<GD@M;��*��y��e%Ou���,�(��v,zY�<^SCF�):��;�N�=s�P{�ٻ���3�J���]����츽���7��I��$S*�uR7)lV�@Օ�E�F��T��r��7ښ8˥�X2��� ���b�X3�0�K��~��taY�_PѢ�}@v� &B��+�h�J&9��'��u^��vE�����S�����0��#M��+7&o���Fk[�EGB��Wη*U6_�}ҽ��Id5��F�)��od�,p�Q� �q��kE,j�����AI��1R^^IP�e�#˺�˒�^��Jk�a�wQ�p���Vƹa�%��PP����i/���;�>��Yo0�m>���5=M�c=�T�P�I!�ɂT	Ϟ�.�;�(I�Y�^a�>��<X0�����*8�D����K��.~\��F�N=֚DAO�v	�w]��D޺���(T� ]`xN[���� ����1�!�[BƎ�����_�&�����PA:��"�bۉO?}��,�B�Q���A/����!KY��K��]�j\����~�iB�p��V<Z����K��_��|E2�F����_Ηh�щ�2����J�v��+0$�ҽ\dYg�+��#�iO�ƫL��EPQ�U�S�%�~�s=�_���� z�83�[-��n녈�%>V�Ln[�al.|��>)٦��57��h�%�e��(�+��n��R��#�ef��qm��z���s�uݩ�,8�'G�R������ #�v��:�U�)�����\,9Kb��M����v|��4ͦD�N���0?A=ݞ,���[{����X82�0{�.����q��v��8��a��5�T^�+2�F�:�9l�o�*b\��X���7����Q�Nji�"V@s��R����:�6������.���5֫"}xF'A�٪vD���Yz��M�	��k6Ț�=��`3�n��g���b�3ڒ̏���]l2�.i���µ����$���}�L[����,D���í�3��B8�d�&/�������� =S���Ѩ�a ǥ:��SK-�r�0p���h剑0\��f2���
e1�ة
b|��}�����R1�Zb��`J�۰�n� >�'۴�]92�v]X��;uy�X�n֕Id9�n�p�w	���<GS±�xr]t�v���'��.v�6{�]`�±ݨv���4Rڼ��o��)����,0��)�C�8��+�U�))��>L��B�����l�$�¼K1=
�-,/�1`H��v�e�P�H�V�BEe�����>t���,��G�͘��v��.�\q���j�<|��iP�~E����i��D��0���EU&�w���ZT��L�G~��̗E7R=�2碷g����s�V���cg|�W�[�1O��r
KXV�hϻ�w����24�S��`�P�i�d��z����Q��5PL��z��h���7��~���̈́f�:�N�A&<ҽ�o�h���Ъ�*J	�Y�c�5"�D����3��?�M�
J4�u�����OR3��䭚�����D�pZ7��\�c��h��8��8��<���ݲ��V9��ǫ�^�I��;	�F!�C���]\����n�RZ�]� �����a'R���c ��q��}�(F��]�_ީ�������c?Y�=�B������y>�k�TX�&	�Z-��wn0R@g��꣫��X�����6�',�«E�
��C9<q"n����mIv��X�Q��N���?���_*琡{�lՏ���9I���U���6����z�#�i1���d8U��Y���a2l�lN���:��Ɲa�?��*��\޴�
"�۽�l<��>TG4#V�`u�]^;uu���V$;�M.�p�چ���E��;��&(�t4r���QRc�@.����]P�ڬV�x��#HlR'?A��^�En�(���L�J��.��Ua��>n��OOk<���c��8=樭�T٬���J1y��ҫ��R���'�zY� *��>0��/���h����~�C����v��0a1nlG�I�J���$}m[����sb<)&T�(��m�"�F=f7��d�W�O�Ώ���5�,#�׀F+C=\�N��E膍��� )K* ��d�y��P΂��#�=��$O!�0���-@W�YVa����Tx�Ë�oFs���t>�����"��\���ƒvЗ�)�z(<�$�ҠAN�s����8/��S_(����\��ٌ��pafIu�T���4�,�w�Mލ�^�������0�ex�$v.���xu�tѱ�o��=�;E�՗��7E�c�)X#�J}a�~n|�%E���*n�0�G������>s��y�ڗ�)���ʉ��Y�:C}�����4b���>��gM7�V��!��c��/D��~	q+�t�]�䳿���)@��P���������N�Bsc��|�]t�)ate��j�Z�c�>�@ ��[R�|�5��R?3!Q���8y!���N������\��x̏fH��3�;�,,� �kh@��u�Y")�L���ق6^�7�,ZG����jYqw2ˈꋣ�6ͤ��kG)��fБ�D�PRE�����F�=G����/8�]�Q�؈&�c�d`�[�����arMͥ��@�4�U��ȒHM0L\*�W|�I~��W��1�3�Gʮۄ.�����3��Ъm��D���H�
�mgr��^h9��'g�"7Q�����6NL�*ok�����#]�WW�E�D�`Q?M3�jlBۛG3\c�94^�u��.H� �'��I�0p��Ks���"5~���i� $����'&��q��K@���	v(~��P3��]�����Hp�3�|>!�UQ�ދq�odVA����'�@z���P�{��V� �u���˨�m��:�#6�0	���-Ŀ��c1}T�ߚ�(��BN'��7nP1�G�K#9�&Uܫ^�ϡ���b5]@B��ZB�8{�F���_L��6;����
�U3{*��ב	��X�� =GƷ�n�/s��m<d| �u _i�bq1&����D�Cm@��� �T�g�@+��@�#v������6g��b�d�O�O���L4x�)��743��N	OڀcNO�'--������� -۰�yN�|��H�12Z���R$ ������xG��H+,�k(����א�yo_Kg���\d��k|8i�y�!�� �5~��� 9#�vh���)}�JҼ��1���z��
�(	��7X�Oo�><R�h5&����L���jL�t*3k>�d�J��S����<�K�۫׺ƞ$?8�[��� ?���uF�P,����\��O��w�_-ѾZ��"(��|ĉ��0Q�Et@ ����ƅJ���b�$籯t�6�}��8�����l�g9q��F������.[��V�Y�W���Bx�``�g6��~7ʈ����$5Rg ��ĳ�L�_{����\�ZP�$���-#��#߰9�WK|;@�غ�#�/3���`��>�lFa1�&���F��B]c��AU���'�k[a�1.p���Ё�"�$�qk�0�b�S�O+l����x��KmvӦk�L|����e �F�yh����5s
$�F�&`���σZ�����t���n7���;'%? &/j_"B�5{�c��A�-A�������"�5�l�����f����N?|���>�XŚ�V��Z:�?&��	�On���������J�P���t{���䰽* ��{$9�����:!�d�
�9��!�&��l��F��ʮ��|�٢c����y�₈j��ټ#���k�5�.�G�8��x>ΰm��YO�����@�_�2D�{��-h.�׀�yO/��A�.ݦ+j�'t]*�Ž���NiAV�}�.�;ouT9j;��*8�ȴ-��6���	i_m���Q^>�bNB42�ΒQx�׌%tق���n�Y5�n	�$��J�jN&��{; (`���s�m����m������3��4�~���+�Y{���`(E�����m[��$<K%x���W�v|�������� Q_���ڀ���hm���!��Y����|�o��2O�[^N1�5���%V�<Jŋ�f,��>�=O�s]�>Zw��3����=�k��^�4���i�������v}P�C�Wi f�� p)S�J��~����Ho\p�����+��%��-*��p�a�:!��Q�R��~�_q�p��MQj�*�O���M��:��bW#*D��>�«R�^��j�yHh`/HPa�$R�^�F��4��WaR)�G�M�|�M��!FA���]��~�f��[Uw��Bq�9������a�|�R��H���E���XU�j��lL0f����`G?���H	(����ӂ֋���{���}�-��+��?�ĸ6�Ѿ*�I[��$�� dn4
�:�h8)�=�$,4��c��1�F=� l}¿�T���rAbjꇻ�Y��z=�KV讳�YK�R�'���6ޯ��(�{�H~�6�-�a ���O�
6�l{[�T'4�4Ωy2���eQ�h�T`���I	�#D7��>����AB<��.`�O��2AZL*=ZT7~�p����A�����1�.�q=T��S���>�l��V��^)��r����F2�_��rqG�r��bv����� `�v""ah�ky5wD������y�6�q��=�p1d�Î�#A}S2a�]4+B�.�G����2V|l���R}�G���jXp %�6ZLm�g���;��n,H�/�p�#)���.��=1�]ȡ�)n��p�]���|ά��<;X�aH7@�[�����<�H��z>�GWM��Ve[Q5���0�*Qs7%��,Uo��}<�ʱZ�$��b�!���-W����9�I�h��4����?.�*Ťp&^h΅��b��>af��8��e�7�Y���2���4n�]���n��wrO�Z����
=ͫW�����%0_
{�Dr����`=��Dm�YX�8q�O���<'��f�J�_��Z������>wb)Տ�-ж���j��*z���Q>Ȓ��
`+e"�ւ�\g&�t��m��ф����$i1�w�6�evh�M����o�8	��2雌���["~j8��|�!P��x.��6z���*�}yOO�^6)�89G�7G���j�l��B ���h��Wzŵ���!2&��0p�c�D� �O�6R��0!�n�U�CMt������1A J��������1�Cxë��i��`��۴z8�#S�q�����9p�9�?q��w�VD�8�e=W= �ÒDSP�)J �7��ut�����?3*D�6+�k��cZm��B�C|)>�ti�[4���� L�(K�a���~�~��Wͼ3u�F(�m�Z��>�N;1����(s|h��V3�����In����%���h���v�]s�����
T���?N�k�T~�v'	�vQ6��*��̲<��fBg�'����
���Q����*��J��Ku��{E���!͐z6ӷ������E��ث8��f���� I�K�|Q�m���<7��|֙F���0�o�g�o� S~Ϯ!��zIG�L����x�qr����ϱQ��3�#����{�i�%@��W�E��<ux�U�]���ؗƉ\6m�B�5�}'`� ����>o5K�2���Z	��Q�X1��m���5��h����pm����2ǋ��CH�炐DP�@�=���~ɿMZ*pm��_�}JvQ��Q�Х _����>�&#��Zȭq�	+��ǌQE�6Cq���E�S	�F^l�;08�\�&����g�^]褃��Q�s-]������̉l���ݔ�Ŕ�'��Xp�����J��Q��"Q%&�<6���:v��j9��§��N�z�d�ˊ����gT1��|t��Rd�i�e@��D$�-��c�=BKk���V墥.i�Q�S}�fg�F[�H8�/C���7-�ĉpD��Jn�FD�_-!Fh���Ug/�(	��ͫ	%�'��:'�'7��o�\"�N��纍�U�g�.�T�T�����'8�����������{c��zDY�n����"�$I�S`����|�RHS�b�J;����l/�iTU$q�j#�	G};7k/؋}���//n\�˪VB	n�|�7"�6�Mn�f=cfgGaI��9��DJe.L8άv����S>�+���s�|cn)K�`��}a��� gvY��� G �4a�G��v�Ac����Du cb(�>��{�	H*�X��|5!�'0Sa�q��C2��� Zl�}5K5M1c��J=f�P�Q˷S$�e]���Z�Q�ؐ56c?
�!�6k�̔Y�