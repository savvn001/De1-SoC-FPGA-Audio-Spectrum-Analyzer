-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eIybL2A7eZo8wSwNn/nSblw4XlzvFReJyV7k1JBegpB3Tn5iQ8Mdeb1KtXlA1/ZhTh8sJfutu7qR
uFQ1i4yGi7bvKennqPNS5aSZr8zMYKb/yVdyOsJhhhbX4XhDbLf9iOZ+oL7vWdsnVU9ry3Dhlsrx
jzd1w56+QDGaeps1zokYkDMKk5aock6fbL2QtWuqDTwXWK740DfIyJF/cdSHV2A+E7sgmDevKCUr
bZ3dUd6BkKB6HUopYYcu00ISmCVmeOIQdBzWF1n4sdm3H+9T3+TE6pW4ncG9X3b1ulIQ/lgrH8T4
fwoe98M36Fj6QS+3tFeujoHLqWHk0Dq+TLiDcQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
T3/8WLgSVXQYyfOkE/ES8XZkmHPYyjPbXDH9zSOIvSEyCVZgCdNgWt+zY5YEbt7t9ooRyx/Hn8uB
SYvOBpPUyvK6LKG/TjpFpzxiqV/27W/8zjTidnwsvdo7z+ifUGUB/JIeYetUaZMQpJPZuCxHk1gV
sOuLqlG3QWfMbviM2yZRv/78w5TwmSo85gT6FeQ1+V1joGuUp8YlO2aQPRrEsaLPeRwEz3uEn4ak
DN1x/JHbHhL0b+EOJRX8yElRrJ9DGPJmf6rVWyWlMZ8PJ1Cj6YJ2ElT0pK+oZ+7/cPDalf6SXvFz
bCq4qEcTEUL+tiK6O6zB41KfzujtnMFLoJB/X9tHSimpuWtqnyu+G+J0cZc8lT0wg2LQxGEhIcJ1
tWIk19L4SgXZo04asajk2rgSloByzdEGXh8fy0bj+h5GIRckvfZ6V5rNcQUJsNhWZuoLFroXReNw
ZLF6ZZ/LXZn0unK2JP7GrGWUxAf1wdk1VkkXBgEALF2zQ07WK1unMZMsZliCmlF4m4BaXPspA+pM
AxBodpJFXX3DfigQFbBPK3AaY/soQtMWkmH4wOuRC5lgpgxpg6OCJ1v+e/+49h38qDlvH0+pFX3o
+PG6YyfyYgZ1i3LdoameYVU/B8PmfZ6ztn9qgWSdseOfkMp+60W6YyA9ifkKljiB+1a6f5IMPLI4
xAUyoELY2C/h0d4KVohxz0dn1H5vgiSpLgjKXPpjituItMJLmtxMaFrs8TvmWkS7HAkUZdV7U15Q
qbzj8UfjBLic9vNeprZ2BA2sd5jV5bZOdsTjEj5YZePz+sbQZEKyNji5APsOhnfAVCiias98u8P+
tAaGcVK7dEtpDXRmI2f6Uxz7fOWvlQhDfqExc/FgpTm2z0aT98+Tr3tkex+CL4HPUKv1Xq+PvsX9
B85x8kXfB+m0TTC1Bur6fU9a4kthLgYygoCtbTSW8V0TQxj5rGRvgBQdSdcWxZeFh9LfXTXOpnQk
r382nGMwavPO+15TL1C29ReYPyxJFow3b5DmZU1oN45Ua60qTh5KznnL99AI0naxBOIm2nWyW6Oy
tgPY2DQXX8bFnH+KwpaOR28BhNCRg4x9IUsB4sbMWiouUQqB4d2Y0s+8yk+0cpksM9PfqUeYxfKd
JEFWImr4RDWjkiLNqBVW4mKd7xtr2B3YcaitD0UmRD5Tb7s+/IYcEc4fKM976g3SxuCDdmuZGeug
LYIw0uELl4WTKxnfdJyj/acgjPFEZdaicZn8AD7ObufKGu35j5IESUaCq6CGym1LkXMr3nb4D5U9
QvXj2ueja1KPUMbQxwF8mrygicpDvZed207HSd+4g92VKSSn+JqjOoCIH3bXtONo6kQXUEbkSkfA
wI0EOK07LXEE/wNFArH34RM149U3M6g3RSJF6j2EVvgorcBDfgx8URJ3hYXfJbdLD+xWoV/QKwmI
MyEa31kb5AZNfTXeZz2rmrnJBaBkcp3JtikuTEN2GyIVPJ4YFIaBFpmTHYnM6bHAcAhBbds28Yam
3ZibynbGKs5+wVEJl9COu7s/DokTABKIXNbKBw/sCKKkqXPeGA5pseObIHHc9fehZ/N462TrFevG
juhvmzYAOfB1Yjnr0khybvsfCExRTH2ipP6m+nlJQa+vEGLdHT/O1Wud5tAKuaGUM+BFh1nYVJ9O
J8goVktElCpk6sqv9xD86KDXSsHN3rAZ+bIanSYS+gBLuagz6IupNUDyChX0B1XhqvPF2JZx6iEj
JylUue66QNl/Hv9kLo7MDKLvCkikPR8WVw6oec1YjcydnpTx1TQ5S6SuCNl0JH9vB+GzOG+BsTHd
ICAKEju2Y45xxcvXMwKa7HnTm6KOJxMPBJy1nXAC6RYEYJs86/i5OpwRhYeUrSAQwT9WFale8kq4
Ewfb6c6J55bUHHUIrfYJ5gHu+gpMZi3VXlh43nNDKpeS98bu72xE2z+eBf73VwMEF+O/nxPOCOmB
y6eUi1mFrWondB/7wasZBhPgVaz56YIQKt0W4qXgEQntMNJ7jqzEIKnONMfw6qEsmSW4t+8zIuVP
68FRmoOp0sgiAf0myi6COLgu1EthhlwgBSLSjbCssZSuUPMVpwfoBYtwm7UZfbrcKJAo5JqrVp80
Sxf+L8tfjxPl8Pf5GbrWdLPfkCBON5NbpvDAA83ldoRXfmGrUp4XbLFHDfRfBa/bDfG/GAlsaso0
jpMC0oBYDXsDyo7GFmt9HMvmqL5aDK3caKiA8ObxC10mcm2klj328k3aALrroGjPjXNk7JOYBNqm
TZ8QJA3AZ6sn78C+6VopDqeDUCCq012USHN7xOf7S0qXZDH1cwwWUm+Q5/FFGCflZoPU/bf0Aree
iMCA+AbqGc2Lm71gUEF6XlmgVmqG3q2e+4tUEUMguMCoV72VJvzH9QDsv/LJds1543abPd+cGu/Z
zbzc+HQHpHAQwgaP6reRrnvdPCi672qkQnk6CbG8jcrc9HAIomH25+wz62EJ20jyKQRSlk7QWz6e
KCLHx4WO0EtMN86IdmyOKGGFbXH/0hjrkXp7J2aL+QE3iiIwonSxEXVAekhx3HjcNpqRDJ3X2OQJ
qUN8d2jXptXpK00FoP+sUSt8x/OConc5FdNgo8Lu9cji6wpKFgBZP7aUwjBIO0zuMwJzuO8YJPcf
CG84gKFJyLG1FD2SqWV7k1Dt120H3A3I2L9Bvl8nywmNERW/QI0rGQxiiad0+4ltuhv3PTC6c8vl
GS8lKrjHeYc/xAxSz0OQVUD0651FwOn3Pv0zumF9S0mDeMHQooRC0sal+D+6yCS9hJRuoTs7WZUy
9DBAjtqe/j1QPWqgOW4aLWEVLD/EhoZO7oM0k+oBvUkoi7s3TPPwDREm2ykeEAWmLfux9sPVHEsJ
AOz1TG/ZeYvnHGMqsjdwY+1NwxP3uNGPsFGSIm4UkURqddTZbpPRwXnXvfWU5E319xeVrdIGmhlD
AJNTZ4dPKt+QxkSqLKCU4G/cg61JlnSmJLL9Odk2HjLI8qPOWqs5auCmH471Vn6A9Mepdai6r2d4
sPGfsUEuSS4JfHBdesgrqyzJLIc9jRtIw5F74k5q5864Lag29ER3rK1cmf7Syol7r0UZynPvcMxl
5py2I1Nlen0rCIdIYdEAok85Qs6vkJT3ecZwtknnI8SVOcy8kdmaY2zijD8JkpqtbVjPE9T3O88o
suLTgOqDUbQSjUYQwYxog4uRVGHm0GvWNtlIMA6nAB2yKQ2ANceW1Nc+NibmjkB8qRwB6Qt6avAp
RLBi67qf77Ty9J6Em9ujGZsXqq7w1SfJ0rt22iu85pskH77Z8B+2zcNX2DI5BUPzWfLft9Ir3RA1
OwZShUQUJJkqMQChenPRW1B5UonDuzRDJWA341golkZn/gOgT6RK+MorlvgFnc94Ee1QFLSCy+tw
rFkKHsuHrrde/rtSz3nBOgwkSIEcqb0sTp1swHEF3Md9OOa2TH9h7wA3OSea+z8ahFGSQk85Dbnj
eVSHGXkc5mVWQOKWV2G79v2Ya1Sh206ZoJf/KytHn58tI+UTCyP0cp4x92gdM4wVhoBFTRsQFEUv
k8atFgk8euThWezSyvnCzht2EguT6/Ea47BFSWRcET1srGehejULAQ27wREEHWgqglZBhadtRpMS
k7PHrvlcs+By+ncfL/xjv0DdneIF0k23VwNo0yq6iI5jtjYnisWYEc+0PzXuyRu+WIJlkPBM488n
aQ/Srvib8lf4H4bmBdXYbaNpzTS9XepvsiYrCk7iko67P+PP+Wi9kX0zqr2gBmggUFS5Bgy0Pif/
vLY70r2frmWp8Fnuoldg9SbIhCkozLJg/z2getRF1+SVJeRuScwJM6BY3RRkZLzxzzSY4sQS7O9S
Nxk8rM6tNWKiS2wRl/rufEqGI9cykdzWf4SBT33JttTW9WT5xjd/T9ih6FJaBFdZrKFtlGG+NAQe
yPm3kEcxvllQ3qdmxETFT5de8pMV5q9bbgy9e5kB3dX/3pSFhxs2BlaC20I/n6dDkmL5Q0vh1Akp
yM8/fHy/SZU8S+baD96qbtyotl88nAN4FRdzMuMwMwe2p7ab3eFyt3o7ikm7IJIkhFRstZgsbM21
bg8HwNfyL6G60qXGCIjr6gbRUj/fCteBYvOx8/J9g0Q1upXiJ/qEf9gdfFIS5wzeIy+MySPGl+A7
ZTeOiIVgFKR685yAQaGTDErRnaLTuU4CIM8H9d0YNJv4i62VAVFzpoQkCTq3PfAwj1eLscGSI4/Q
O167ExNtQHu2j30pRc4wq9nKrcp3qAI6+pw1iCdWJ7BUtebbQQPGXKu2c+87fIHJaMtefGKBlOcl
jK41dJjOe8HTwQDXujaqvn7Vf4Knp7HspfJs7R0TQXJVXbp8+bsPvWCkszX/1J+SGqQosZiwyHtL
UYpdGu6ekDHIisQchTGeBjtHuM5jx0SBxkEqa0CxLc+Tx/calXytUjhYRn41OJKlPvKoYTd+ZlgM
CoHCF9ZK40gZ7L7OU/0sxtoUXddVWHpEYy8GDdN7/nPKKwbDN2y5kH1z/X7a8m2XQE6J1ZI3pvu9
VJi1gbKpOuHOKmQrHkfP4sOvlafm+w8QC/hOuEcRYrShqBlZ1gtfGpOKpZylTqxjotFzIwsZueKo
SV1uCTDnaF3BpIMgWwOCcQL54DjtrXnpLxlLSiJyKBtg1gJ1MfHW3wHklunJxS4lpoMBpK2OSue4
6JbG/Crc3n7PckjVF9g8ZQnNu2I7rPHgmjPtmhHdibv5xpfPesAwX3DFBEkpyHcTPXzNrdrYQdSe
QzAM5AIb442tMAJslApfHNyx6C42UUP/LfziyxYdb8AQjlN4PD/pypnqC6hHm5UHBBMBWq4H0Wyk
llXM1cCIavIXhx6N44GCai8qs3Siu3WRbYAx+4cf2wwN9yENNMPMshzCrsMLe/A3L+LVfXtSP0qI
db1sJJye+7z10Cy+enu1nrTxd+C1mZfECrurE3jMH9AchF0lPxK2FImIDB9OWpvLsFYP3IccdhHA
wDew3wYhU+s5zin4Wawd6zw8iRhMuJuTbTdv3DZlZWLI4+6f3EQur/hQDLWzQuELPe9O66Rh6xfO
AdKY9dDzDbq7HiVAjqXu3nva8XfK1fIb+eA+utl/WId6ryF+CPx0poJZ0xshlODVbh3/Umf07BN/
CTgxMIheQcVDNNgQ/6FYE+jR/UOMRnmKD1pm/2SlOHufE+I+woaUaC/MwJOwqgOztlwprmpD+LkW
mlCRZXBFFfE7hf9xFoW9pUwrfQ4lbRiuQ8OlCms93jlDsF9ljZUMSZVetIzo3nsXjQJrmrUAhn1I
YI4dr7ZBJVKzaLDvaA7LYzvZNaNBf3d27FKEaZ+jBPWhzgITxmw/zfDh/P0TiybOnvHwtVpJBXC3
nsoPlMgKznR6UxShu5FDgKaPsgJT5Qc4eSjXLJUJf5kVCGeBASGPHkxPtAkx64eXjVvZKjxHJb+M
2YRyl+ntx2Yh+FfxrQs1riR63eGL7svr5k8UC5Rs8iXXQMWQsUEB6qU3BJhyYIjf0fQhxWgwT0Uc
0d5+bO6jnTXu27H3qqvzyCNL3+AH6GAcR86fK+BtN7k7SKIKLoaGKSngev190+J3bWwEpf1uCFX3
UFLF6Xo49YmzMcFGAGaDfxtZN5iXgxXEdyqahF1GczJpgL9jb2KJh5y00lyMvLqf/wEs3DAbLyCG
vXlAb/tlc8Ba2bh9wDMezkX5MxI4FQ96IRhkM3UIH6iEJfCYT9Sp31LLgsVtckCE0SpEgEz3unrI
WM6aBpVZ29ZbeVpNq4AN6hhhUzIuzEvBYgepugxZwulrCdgE75g+K83fIKdlxYT1t1WZJdWB2cCs
Jo7kVJcdagCmw+tlY+gOArXsN3+f7aNEKXtSD0iEYBy4VE4BpwS64kc9uNrQ8krtPLeDxl4gxKZS
7FOfia75eoIEpag8XrYeK5QcZaa3qkwxFxnqlKc1OdbyD3jn4Tse9VIpx6gBGjYYXtqKE06I+WGw
5Jl+7kZ8FVWVQli4bKb37rRCxKbb14M1bN2kDYbpGAYtddezZaHYXyp+wNuJ0Ma7eBKHuiSDRrmF
cKGwwsLH34EN5415euoJfCJRX/vs+zfG9lO6PZIAKvw2SefT1Imppr5gLbEk3vTwyeAW9nNxBKao
39awqLfKtWl0hGE670ejDPyUFY80fQ+U0rDIp4QlXKm8H14CYn2q2vvKu5lI9hLc0e0krxBvyH7C
3ZQzwLCr4N7qAKj2u64WTBQ6Z5InmgP6/YDOf+oeqq0W6X7VoS3TS+XKDmvVK3T575NZmoyRXHro
FRcaPnq+GNtyc4khA0cL4l4/XL5V4Dv4qCEU0cvocWIkZRd8Yy6RUDgBdZZArc3MbYg1qQCoS37L
7e/wriN4+fTMXIVWwPIo4sP5JaRzs8FPHLdWIv8DlLvimM/UI86J5jpqImGOX23ijOb0O1kte2wg
klHnvtOLbhjNynlf2Snm1tRaqxC7MPXEDMsg9RsBTXdBebXSvfvOmBlfHozSJ1TkcWdk5Vi7bJRd
U1eimym4vu6MCv3h174CZ/U26TTtPUD5hwcGgd9oZWMempPNZkvPt7m0fJgdhur3XsWHS9fwknjC
/pYEPEvawOQGgDT/NIPdVWYeSpqDV1zEN0pv7Wpj0IFV+zE/1earCNwd67dgvw1icyG3t8Gqe1Hn
J/zXwkg/JrD5QKAFVPnQp68B2fm5T8S+Jdq1IShZgyXLFWiQc+iJVv5BmpX99FXh6mb6zrI1SG3U
ySA0CtD9Hjfnl5jBzZYuvI0sOReYUOGW9cZax65RPFWqefwDcY2fgwxGqAk81FKBr/4yOyHa6XvG
nLkoZW267a13CV+l2WaZZHhv28bmIvvQHtMFZBqX2PcRVIKj8HQxDgjTM5GPDxJpDbWWEsdzEpMB
9MeMXPweODDmr2du5JbnFdBOi4dEeRFsXPMDzm5p7Cu0gE5mItNv1mah4GHeqpXAGX7EPGTU0HtA
3PU2i7MoIrwDRIFXvFZDoCHfPMQmry7sKVRcBH16bhCjo01y9Ro1B+phFKY42IrAleS3YT06o97h
fAFi/kHiEk9sCfjap2l6ODIvCA9AA/c5fLlflK+NrUJni2zVBm5TBTX4DeIINOUfbB1uhD2j604d
uf19VhSQqgm5c0nnHcSZG5dZLSi+OGleHSNjvC1hwTZg3pHy0xAOpG20F4F4nOOj7b0iaQATZFQs
jC5wJxhVnjqG6D5BGfr6/OtbhFKr3zLPBGLBDXq5fN8aw23eLWQ1WSgWkewf0e0aYkNbN984Wyfu
LIc+jXzKuim37qbYlHGQTBPGp0mzWoUXdiUh6AhjAHJ2QmiyR26TI4CE3J3v3i8pVHLIx3RSBM1l
NLq8jFV2OO/2aNfpvt7tjhZtB4amuivhT0KCFj7OmeqFXNjmcLKv0Ar1KnZhGnROskVfzwzw3snv
PmwucKjDffpHdMN8nVTHI/L2K5ES2YkKKtZaWj6KeSCpoCPdMQY7l3WJ8TMJIIdWaid7jyiEr/+2
MWZ0TZSJXH/oGoKrfwiQ0RuxOHeBV4SOcyB0fIYto+HTiiUG73hlhhlRFKT4awOXUZ/NCfj4r2vO
sfb1cvKwzhXXrRC1bCFxVUuXonY8jjIaLYw/BeBdB33OJett83F4c3t448bBWE2bKMcvNpqX9m7Y
fsV/4h9WTZ81T5r/eLSUYkJWToysICxTfO+T3spJGBNJcUj9kG05DHV7So/rv25wDWdIB2+l6YfK
QtkOh4OSY51cbjzE775PYz4zVb6rcUs9cR9G+SPcmMBR4vlA6xLtiRHKaSZnNvds6qywZRQdmwqf
FPul5QB8e18UxE2S7erqaVKy4AU/A+AoAX8fHeQdGLhq3tWNyaeJThQEWEOBaeHbBhVCBPXJoNki
z5Q27QWWPmdOR8acD/F7YNpC5kOUiNnRv5zoOlfr0ddX23UR57c3IHdKeGtFAOOQYLNwBGqa/T2P
jNUEbOpsqswwtVIfYlXoIivzagfA8KWBFK88/rgl45RMybXuvcEdH6AQRwhh/9RroV35LsB9m41R
+8BTSsMluLEWsQwvVP85YExGuAFEIGIrWUAh6NGkKVwsq6Il3+0DGvGQB9CGCzVLo5KwOBL5iwx+
fLYQtu/pjG3nAX07CGo7SlwaH3sIQb1VxRsJtAiEiXHqtM5wEjfJRcstVKuUiJGNLBVzzj1F3PKW
0OJv3OeoIQXehe2+iRy57QYHPPBFh/55ORa8QDelGk0g/INv5xl8nRiIo657cAvAZaWWHHbgMELJ
hseobieMPLFrrNzj397KaTCArxTPaQEK9VOvBLN1qOTocjqUiGta0CAY17q6IlpS83z55JRvlJ2H
ur7cCqVq1zdAQBXzH+oec/2a8J7X1ZQLlMb/8jwTDTNE/TwU8sbcgL1vaAHzs22AE+ZJQRK/Kydx
Il/XuNn8jdTrpHodZDz0m8hsZ97YXkEnQyWg9yRyIi6z78h8pfjRCfHgrGDKR8ds9o9LU//liMrg
vu4LOv5eICuPmyRfrq9+x8wRv8Xe0Bvgmkzbjhuu5TLopNXiw85EnpNZ0pG1YbXkg64aaHmTxEjz
2Wsd7GasPzPWMgykseAalMT4OKxI64E5yoY0tSvqT754drJXIuSoOsvRt0OP7/7A8FPCg5fWorGh
dnVlGRH+LxSXeh2aPM+3OydHP3u7cfXHPcklnTqr3PX+b0Zha7eLyWmAfWA5yEA+TBTmoLBZqzFo
PZWBxbSDwB4eG4/KS/WDhMRfH0gaSZe5m3LuZ1Yhnvfye1WtDLim2GMZOxGQQXYtm7TDG61EDEEb
kjvTG/sgkPm35EpHQEVMTR/EgX78UIiMScm6ta5nLVJdbXpDBLEA/x5+c9b7yH+fhFtR4KJySo9N
rG+kjzn7vVlDD0cQWjQTflCk3M2u1DCNs1Ok7UNV7k6Jftt22sHS2JPIYGOGFEl3X6lAHp7oNRsM
B7r0Z8vJZk2+EW/ibC5JwmiQRh6Sm7gH3DleVlB7TGACL3/fd1ZBU6ClJmyTnEjDlHK9Gz4qqLDt
0W3HC6yf3HalYNHW8Hfqh/Nu6P5GrrAkgVoxH/UhdH2vbv9BWzdx69FP1TrkwstTG4idxBfUhQH7
ud5MxnQnr4OTCcfL6vRMJqPmmVMeXcWEqcjrkm4+QIIpbO1h9pFhGiz5f/HZsi62MbizYV612pwE
A/Nor86U2zJwIMzZmZyzNK+Wv2UkPeOs1KOMLtkxPz76R2tNKVYYc55mDjfxzic97De3qEupZYsK
k7m6IDW2rFNjvnjNQkI+c6rtdsiqQGu8RTNKxCfjl0VQwhcCSppYX1SNVa4GWNg2CEEV/tzYK0Pa
2cU36WiMoBJCOjPGyvK1Qde+54RsHYwau0mivaW3NxbUeIfyaDT0cbMeEqALJGOhZzq8WHhSvzwX
yElMbLE1C5uE7gRAXYEWG1WtYZI6IraeWkL66HB4ofKoZX2Lchg5D2DLhAa/WIpKtXUaZY52WtYr
Km2nABd4AazokqbcS+NDHOWhfRNXdLw4sy2J0v4x6VVibzVWrqaU3x+oBjyx8kFY//rdKQmfFWHt
GIkf7CQrfsB+HjDbaoeNy6Zo51DdQJt5dGJ4vE+z5rWahiMKIvaAor/C50tA8JV+PyzTK4FpsQrA
FPnvUDdmAmOJmRkXfWZRAEv641ChfU2rv/4Zyl+JilhOgJfZyDCWtpH0QFZ+2gmLKmuFsqSo9k8M
C4E5SzwA0u9LHwFJEQKhxn/8oCq2sDFyEom00exQ9PRoEOVhB7z5l3qB+sCD33AqGcrSkFpwkBdG
TMh5dNu5aay7p3PtN+AgZV/nZ15ffLlPJqePuCM6dDGt2aXtOWH3dT+TmKd5JcA43mcFlOSrEk7K
6ZVYP2kuzvCrJsrpz6liko5Pn1n1LHdQJm2dwkpKuIVgCQcaaw5fMrbuWGbH0zLehYlHUgtXxnH4
1RkCcpwHuW1c4KyUGGLd3In8DCe8bgh1bQzZvqekkU+BY0GbtqECjyQGvCRepJbK9NvAhGxtYZiX
TaqGvwLCOgWmMBMeY6AZpoS79qG+P9QWSPzd0NdYuXzT2Mrg6tqsU01EwJQ3CAkJNn5S95p2+++a
qDYjrayiSKyRMgiBhV5bXG/w+FvBm/O7uhEXDkfuAgme/M7o9I02KeOWQ9g/8ZgEnPURkziHBgzV
I0gCpKhWmt2hU8A1Ltmt01aloqJMcJYoirBYcQkz6/wz24uld3ZtD9kp7dE2kSYod/K9lymtsERy
AQaRTLvbxwOGvVOcj0AFeAY4fP44kcnzhZq4+udAxn9uiHMlMEuPgaHBdmZTph+F/En7DVuUbQCk
zUzdRfxKAy2bTWjpH9GT3s0xKK16Vs3RT4uIeO3jrFQVDb3RQY/MrnrYtbrON4ieivM2OC/t1LLf
ya2Xoy50rfOoqxRsfUQBYiaw2TrQEAwlgx4nZ0WFfTcnGh5f6DwNQR0DmOvA56rtKk7qXRimaF6o
iKXhow2/qrPqM9rF2p0Bm0c7qNKkEgOQ4ZD7hgugGWqHxFLOCnGHdJj9NK7rxyb6N7tSFESD3KZf
abhrPhfpM4tWr9+DWy6LGC3CF1pX4XCQaFupmjP7OQJ4L6Xu9rJRDNurOFTy0p+JaRVwx7NtKJev
qYkAA7uD4Yl1Hx3aRA9DULD9tHCUc2jsdhRZS3PCeLLLLei/aJwB3TuWO0wcy1J9Rfn074nmW7BF
EFZpQGlGhr937hDDFf4MiYel7tw/rQ6V079W0vyte+5OasO8K12mJyRiRUlblvA9DuTLtVv+Vwmt
OQZzDGDvy80b0DlGBPDZ6xGJhLuNJMPFmDr+oFtS8TzvcGYUAYS6keT2rHJ7u0mqyaAAn9w7++bp
IAZsQsRTo9yQTC7wfVqkDYErcC0PH4RGMOn/X9jdZYnzHdFYjzNJIy3PGYgSSWEFpMRlvOGYeO4G
Hl3uoRyx7WfugwUZono8m5OPTpXxOVUqvV7eyk+eoTHUUJTcU6SNB0jt8QQiQHmpZGWjldbIR7aT
I+QdA8rzzDWlrnarzER5ZN/0Pb1cx9UJUnuDX9zIrip8lsRTXVBJBtIls/GyvLpxpUXybxBunaqh
6pFj/JKpSklT48RPrJoXCvXf+dWvOTKBEHFHoUyt/WuKr9cCTBcu3eDFT/bYebELVNjNxtblC9je
QwnEY/ejiFAes/1wPbnnGl6IwyP0pAQsWpBwZx+f8XRJoSOl3xa4UK3eINi5ShIMOZnnPtLo59V9
b8xiqk5a1nPjnktLf0h9+ku38HIG1BGscKv59N9RD4crwHfIgY9AuyM7jYRWGZttILsH9O4xcEiq
dAUymF85FeCymVnMKJGvEaZEAXOyZcY3NDGFnsUxzuNNeauU9ls8EAC4URjaxSYWCJG0r/Oaz7kg
TIIiHGSD+u43WBhAzQQEUQ0j3WeEOJZXQHBmANzGDTUNU+lZ7NKKdc4M6nDR5nI2ClUegbJbodBV
ou7tu8dy0g3ZzrNc20oR2CUqE+Im2zxvmrpyRgztF8HwaNFoMWTheG0WlXB/SgiG3ZWuDyWpb2pN
5CQkYwQ2rHHMAu+/PgyDv4D3SrOXv7e1NDaZkakTw4T2aM96L6/bNDSfop47OvLJGMH7bCaJ3JDc
iV7kjewc+Bg+3es1BGJ14KK8YQrnHDM128WCyCjOQRGB1199n90L2RwZwAkhny019KojvTteMNPa
NzKarnaIAu9h4hsiVHII0YgoS8xxVjj1ClNyem/E2fOqJv9FZ9IJxCVbirOPy+GxLT/sEz1u0wrf
cdUEq7ugRUAENGmS2a/PCAg3WBXj4c/vPfbkwjTlItscoUqGh7dy2kC/421AW4LOUla51hconzXD
k051hgxYAr8Z/XARuKH2Ig/FP/4z9NztzvUIqO6FBLqxrYXzDxPEYBFvctSFpJ+bjDfIWkRqGp26
IO5L5mFkSCeNp0HWbG8v6qbelEFr9h2rrpP2Fjg8t8pC+A9NzXPlxkyMuo7HSPGjNSexhUEstObu
X8jtQTRoBtkcpA6+VpsuP0isE0hMwCZfHwhU1qi5abFT+butofzPjojixXlje/2bJBAUvFa+exlj
n4tkuxxooJBeHckdfOk8kbv4JJRvJH/LDmHTVrVRyd7/8n5Pia54XTTTUY0KKtMAGmRchuXR0ROG
oHJkc8yXy8NrKFSndb4z4TuTc1Oh79FN2J0XYo5k3dS2031+VNFtWptTMRbBen7PQuo7m3x49BNd
mzMsIIodcsP2HGaNye16DDUG7FQDKt0NuT0LwMfEo8fAOX7bqaebeNAnes+Gt8EWqor8dBbSTrKW
rgjQAlON5r8tk8aOSfrcWuCM1uGARCZ/Z9Ux5iQbhaGjh/oJMqoZu6G2644tEJN+erR13Uhpd9rO
awIAGAl5bl1L8iudQC89YuyPefs8R6tWYBNd8RUyAMv1/W4Y+7hh2FYDBzHo64XegAdPM1XzwFcC
l6i4QvlqQ09xe0TTYkhh+uog3cx2niJnCzOrn/7/Ta6QiNqOkgrNhttFMuKeXkFPQUXks9Mi9PXa
gD7pGV6OryjPenm397ZKNM9qMfdjYlsfdKB4zBqR26f4gYfnbRGG1L7AQBb9m8G+Us8IY2pqTt7K
xTrZh4EGKPCvi4iGc5ztCgPEDXfLErQQ9pxTldlrGKaT6C3yStbg0860Tg8sZ+vvJQPpgTAM9Bqp
eGIXJ1mrHLiQeB9ydjTqZHZMXScXfGc5WBJfLm/i488ZoDqm/BX7MkAu8WwraQhUOjDIRfdR/9BZ
RAXvGDI7FS9jBL0EMi+Po3WKsmk06+fbldWhAYPUMbYznDBgDpU+hHUnt/93refpIa4vz4eMsEw/
xFld1xAPKfUvJ25kuh8y/6KJEYHUv1V/vdrGlZ17QI+UAUL/gK+N4HiuwfSwaVyKm++QnYLerQi1
JqSX0VCNgsxfJ4jsiyRGcC39jtTadlego7N/XK7pRxYkszYyvXfTEVxSmG809eIHpHYaeJWP5Ikb
uZTSJduoZL9hhJIaTayo1PM0xYYN2MSODNU6aiHoS645ScXV8FInpHhQZn2qQXW+rIBfCKEbAG3A
DSR9DssbcglvY5clqyVsPrIuzzgjqhaBedN6sMyASwqfpW3qBmDTOX5k9xxVf2ebp63KDfI+THqF
zPJjTwFv2cYaCVS/auvjXIQ3gCzitT8ePdtqKbaezNbY65o/ws67w/Oo+9DdE99fL5588/pR4Qam
+fsH63CI2AeAaBH0gY+LeK0Vdrsfw7ZvQi2cSJrj0WLXjUhp1h29o9op3jDnduyCEHXisfVv1WOK
iGO6X23G3SIzWAZZhvMnVopMkjoT1meaYSy14JTueodp1TrtDWYaJYOPyEFses2cMJfBcA7xxmtM
dm3AntYP3CzumrFCZBTzyFY/AnveAdAFvZeNLEDBEjLkfkMl+7qgvk/7W9toYXKEmmm+YmFzO9fC
N65ep/ogmuFpSOa84G0PEZOM4yd8C8Z/VA8TaNr4G9kW6isb1TfFc09BNKpmDQO5Ec/NUMIc0lJS
Dk+nlFTKJZdUkUhCtCj823qVOBNj0PzSm9o+6yHfFLs8u7EaYvqSEvZeWzv6ya2pWDiXHmOwM3VD
WzR8BhIq1DAvqCy3slmZf+YiuioZVl93xrDjAmLIpSTaRX+WBLvrf0S55KLvncmL5c1+uPAZXrZ9
Xw2IcZH4Gs0RnsmR/dFCh3e3w/GOavBx6htOm2PX8t7NgydTrdWNweoVw1vURYK7hQxk5hsSBkkj
JOoUdSBMA9UPSKLXjWBfoqUEbkaj+f8HLpcuFVqmvvaP54hVhuAgSAFbjJtFmq42uHM9IBOxpSVc
5zgXowKHIuczQmrlVcBsccnK1Ya+UcX0zEnzrpVFYsehiVLaBuHF7RB/M2IwPDuOHtHdzaOQGhPV
5eVtlksSnbCF7ZXY8AXS+dJjLTZ1+QqsER1PJCHy5Y1qb6AXudgSZKyuHCYe49KdOCmVL0nmfFS0
lH0409HfUaWZ20IUIpKKFFPOoEm78R1s+FZRRqO2ySw0AtgNAqV/X/hoAZyUZ+iegdeOYnTP/qx6
uuUkbk20/RHrzqx5cscfAoPAKrmEq+IwIJiQZzE2HxBgRe/xefs5oPCEkuI3ACSbmRvza/LGR+xB
ci6WJmAkwL1fqGWGRCScRgCnLxQCDq5baKqi3KJAz8hg9Ts/FAcBRjubIEUy00wPkhIgk9qFjF4W
1/Lfip/ksJDzb/0ziTj8P3y8DqE4Ebp17JanJrEqSQaeOn/a6SVitpC4E1tMo5SR5fvDIDjFGtMx
qd9fp6gqvvZgO1bTkVST0cB5Ge7V0SmJN5zvf1Fmh1qljcAeSsdZ2NXjMt1IsWididhiAt4xAkho
rsQSLp+u0N5TEcbPUZlUjUFAZkswbD7NaNezdNvS1HAJB5zxxWG6nkvhIbcC6RueHv39e9Fhmewu
Vq9KSJSBHRUwf2qmxpdgDaAzuXsgSb/aoXZRg39hOK3rNtpnYBVIPuqfja/57e5ah8Bo97yzD2FE
eef935j+ZyGnF7oXcuMSAjkYAZlNLgOXePfDQj8Nrcczoam8KDn02TNvx7uK0n6gDO7PeDv1hS1G
AgfKLLS491JcS8n7QKNniW1xAr6vV0uNQMBlZTxPowhF4g3xIuV0Y7fSdaH/WBIoFO86FTUjEIot
MAWSKCm+Fmu75mcBH8oRYwwb67DA1Nd9msnzJqNRh4yUSqUgHXQ0ulWh2YcGhxNcQFkRUaRjAn2w
0ZieK62n+tCzBDqYWu9EPJPbtFnSxxGMGhERVOTY+kU9OU9D0jevVL+ERrxXWamvslI9irN0rbVL
nLJImrLtAIgQltVQwp5mT/ljTfVkDVJaXZ1xbDJh9kAkJ4rqT+A2vhDjUjZOjk/bx4st6a7SmayQ
Uuurv5rgW4NlkirbTR2nHamNSPbAv1Gw1fNJpkMoeDGd59RahmwQNNSwlASwQAGXzVNyR9rHjhVB
vk/PU7YueieGqJTz4Od5S3MA3dmkm1gLaI+NYRHgO/5ACj3gLnxtlP7WVoMHwYSbHFmor9k9vZuT
UAmEgarFm61+xvqPcgfRz07N5KYsSB9W9Kc0S6mHwUP0j8OAi6Bwe/9R2qZ/RtDLYl69YM2SssHT
AugjyOMYeHbUqXx8L6JHrqOP4++QYpr8+z8nJjAwZlEQJvFfe6F7Mhnfk9zGJjnbO1fkMrJK56tR
Pjs154Hy1HihDW1yAJDJzx9Jm1M93RAXfx5eWNlE98KraLLt3lA65COna2KJuOC2UlzyMd9UUipL
z+T2LwAS4zatrZSMc+dGHN+L3dw2G7ONE2lwrB8WiA4kWhHNO0d4r7PKetH/Wr9zVgfNxlVdniaF
328wfupJWqNWfB7hqZw5nec7nMtycz6sadehJ3t/ldSggX41z8m0HYfl7MnOQXhKUxZ93GrL7LXS
2MiyCVpyrV4hlozxtmVKLX9/3fSsQe9DZlfLnjuVYn7+sfrJHEcNjQYVnp+WDYGblEZ5/ubk4pXU
enTM54oPwPLyIYFiXqgzPJg2wjiP5REt9rH0E9edGrxFBeIAA4R+79o3eaa4kNBZw6YxIXP9g/i4
Zs4qkNviR/5J9B8GVkAVY1JlzP3cTAK1LoYCbY44o/3cON1im2KRrU9dJyuca7fV+kh1pw/p9xm7
41veyEoSyMd9ZejQ/Hxxbw43xAOJJ9X/InQAfdnU0HhSHQnzmyCQA8xjDkPST5qJx/Ls5ah/mCB2
e6xhctahcB0aFngEFJoCnyRf1Um/SVxEr/ywlswAtZYI+1QDdHiEqTHXpLKWI2MTjQr0lS9zeoJ3
TjZLqI/h6QSEPJlWzuhIwA6UKrin+I0meGsufpa1+I/JY6mpeKt9GF9+DMw6u9B09DFo/fYhl/Hj
JmGYj8GVM56BPSxF5Z80xd1hSh2HzsJerZfG1NOPcYFYG16XLhW1CTWKXOGvMXS6Wsf3WXfAg/OJ
uv38TavMLlxydvwxokVrld54oyD9hzRtmETijHGzIGxTROxU+Z6SyIl5q1td3R2kZ/l82+ZG7DIJ
btLQX8DdGBKhyoUEkJC+iVKEYGmLlSsLqu9UiVZE2lgjPHXGF+ZAo49GWUJZAdsRCyy8S9TZPS7g
0ag+VHF/h0YhdEHm2hFT2ZRGZdpgkzmDtYU46+fHl+E1hA/zN3J17iTU/Enx5gtkmGNyR24OmhPE
SpXN9g7BayILIpL6Ubug5D2xoSNS35ndQ+hwRS7YYAIxjnu5k0rAr+iBeUpZyb/yKDt+X1KlXWCO
Ta5GIK2alve/LLQwJoAGR69gZu2Hnt05GAH6RTlfQOgC7hF5ppfYDhuesTAO3YRfJTRKfUj5r2aD
dN/jUqjPbpUH0gJq3UPGXxGNevj0gH1OBCZy+GUJUs/269+kykJeA/aCFe972Z1Zz5BGB6Hom8wF
n9e0RLu8KNKWNlzueNdTjF/PxqkLvhi8xxqbxdeYQnFVyiJR0/+tdxPTTY2Kul8o9VqxCgVFEDOL
vQBKNKXETfMvNSIe8vFGqSjBveyk2S3SgYIfh5C5sJCzxtIXNeNzmRDCQSITelN7Tj5nDeGdocJL
v2dtsYFxWgLe1fy3t9pb5XZpPyTTfG7ZoLFOjeyvaOYjDWLdC+FbwMlLjPQAkmWvmPcmK2seOFRj
xR4DbeDFjT8LwdcDS2xvgqxcOYN1OOGn1J9+H23ifCin///n6iOoJrA6mRsmkSkb6G+QKdf9JEJG
4z/WCqqSX29ZWITED0WzL1xUaYdnrCe8Ovx2AuUopzzuV4pa0VW4EA6MoRa+LRcB+4reL4CI+QDz
fhvhpBO10yA61w9M6xnblSZc6jl9oZcwG2DL08gfsEsyyoYwGVDtZmviAOXceHZqvOCIC3tnjBg2
NRYbkuQg+Z/BDVfhQM3/BEt0eC2zOIkwfqPyph71ZOJTue3alzIaUPJn4o+DJtkOyBTvF5v4s8Ju
5ijALawMMLoUtRKmvbX/k4BeZ5VzcLpW0oJ/WBOltuthl5wlx/0fmFj48wDn38hwZTIWpmIfHFo2
1cTN0WTiomoaYLIExmi3acTWWArWDY3spyr3vBmnoiS+1RFrdK15AX/aTw1KKYMe9PUQK/IGp+mx
m/ZEHbSi9+DtWUv2og6Ri+MMv2Mo8crYG9EqQpSTOoeJZ7nB4GUZDO0kGPQ+fxDVr5ZXpmL2Y4+D
06c3QSIq5FKdzaHE9sLT31sDMO6F+Ib7JHAiWgIL5Ob4B0jiRpQejuXZYbDh7qfN6fpK+H2jiRpF
H/ySHRN9oWrIcCk7+PB7iH7etoFhW4dd4Z6VG5m+d4dQllX5q00Mj6BSeomUdL6V7xh2AeTbPfe6
G0UruyhuVX5g/ux8Hl3R/smeUE1zhhNACh/vp409ythb4T+KwJ1tckx9L155F2i5FMY8TneMB0O4
OnPs+c+nXsqgoI/8diOpgb+kUPqk+ZSFlCI5CJKUJxPr7VNdFL9vQcobs3BgP9D6aXU5yYkQoljZ
CIVqslRnshHItjS0dGoe5ZUCYPQ73o6gZ6hZUtZ4xX68M7DLJAQUavNkgeQbwx49jNiezT03CbCb
CIuxFUIg0qKixwp5Yt4/u/9ggeVuz/sD6lbXz0FOLaAYm6MgfwMQEQyAxs+7DbqFRxYTDWc7PTl9
G2kg6X/Ik8fUpLQkVRomKkavGJXVyV92AQn49wNDVq3SPQaDsSVTu3i4rZpCOp9qa+puAeAOOP9z
ThSFHZZT9I2sbmZsS+COXmT3W/EZMk0aHS9R7GuqwD9To/xg8sOhfHZn0mZiY0dLWcpHuT3sykSM
pKxU0aQt811LghwTh9Gyj+fLD8z1qOCDrLniV3+BTtA3quOZAHCoKV8YKTYkbF3FNj58Ik67sfTH
9LFgHQmS7XSj7VHlAHj/qlxy1ehoertxUbQFh0wIVV7nlqsYF5g4z5+hU8CWQD6KLBiBYiGr2ReQ
0k1K4AzoOvJKWru1zAzNAd1Gz1LBOXoKcTlQ8ouDOHhwzEcwCLy2kPP2Mm5cnK+xH00nDND7TlMs
zB0cCcMmsg3JJsGDBsskz80PIBIY6AgNEjViPx08zZ5MvIxhH54xUzZqd1lKTNfmSTgPmc7oMzNU
i4vRFRsaZ0Yy8nmAWqkH/g77WUzdktepy7rhYfnPoylM5edpWskPIq0nda/oUWQSjkUGdpevAIuv
xc4HnbcHFAquuize73xCtJFsxABSs96IvndcqxTcqIu/Ej3Gk1bh8iNnvhYr0FnDehRV6PwqXHDV
41LO4dX7QCrqVQEisFg3O553AmK0CgW1hWZ+ZnwGLjAQxCjEWm8lUVxCG2y/B32Ao+5f8TAxMovQ
gS6cbfrXvzadwkSMh5sHn1m/LEwOL35VY29kNNcIoYIlGN0TWEeyZLmUSFCeEklgM1cF9/qSLe9q
MeHwAfzl8oRaEZZsOiZ8+lpXsC1mry06tMmtOvZnscGLRqeFMXzVSCQprePy66Oc8vK0qit81V0H
8fsMq1oILzdZBNng9G9yhxjHEdAB0J4npGPIX52ENnotHaRfHeAwDHxZyHzDU9OOUZukoqwQn/uU
Me9MDrX6bs0yGMxW1HTMOxySMh5U/RChFoIjYacdt8Xf3/QBawZg57yVEFszN5866A6zhMlo7rgo
gj4SSAuP16YxGoxTfQclqUmVylHmbs6PgOmBDXRFy+f7dWmWcUxSvx4zAEh/ejoXg8FwbDKf8nTj
a/gCQzz8viN+CdFqCt8MdOIN1QEL7Mic2Uovg9PjCRP3VmrK2L1T7Iag6NcKCisPzG49fft0KcER
Zx9je+LC3YM21QCaJlDg/eAqID/QhyfD6ISBJrV+mDOJG3yWndLv3NGbmStb5lZs650SyK4Kv/tf
VsBzllDV1sVSALxergmG3mTZVFkaQ0UcONapuZngmASMyOX7U/FdNu/eRgJPnZRrtBU4mIckJ6AO
vVJEqWRQjCqpWf3IlKpx7ObfedXu9yrwGEsLQz1ZwmEKrCTziHnhjOyQsPrsN2IhGI9rMacyH1/D
mUeomnsyGjKPYvjrYhB4RPuJcmI7V6smgEX1QUvC3zmLxBGPXy+Am1zH9hp4VaDexCuj8ryaGL4f
HMrTDYHFYorRrKWdl2Z7ayiguDvD3Uo3YI8+PDJxVnm/HklvYRlEluKEJLsp9X9/oV/cQr0+/Ov2
WgI29bXBgYucUsRgdXKk0rNN3gOA5YP+UyzttxB0TRCKm6rUJJhfZUaHz/bbrFpz6Dc/K7M88HQc
zj2bAuvgq5hdGW6rRC5xvK5SMZCHjSTBZQDP/7KkG+3PEmcMki9B6UR/gemXmpLVRsNWlOByH06l
8SK2dmtiLEjGWF4CMpHpHSkuvVAOVS7f5E7ruKSPg5EpeZx620uHqK8Aw2Pm441qun6duMIqeL/t
I3TjDKyOxz/tpwaHn4J3Xu4v0FUmrBnnQAfHzfKYJAIvdGGwRWL0oUkyInWBNkozxin3MTN3s94H
lKt3MZRQA0b6p/naTGZywIsvHXOsP9RcS6BQjTGwepSRMjAJK0OhttEzvWUJoPrCNucz7/Axdcxg
iMQYnJqzYTfYOt/1cO0iyr6usaHJMnqvzMvbG8JEVtDTvbIe+uJn5dyzljEELYGTaOHAi5jHBl7/
OxHlfFLu2q95SUKxsRf4MyqK3/74ySrw8IpuRGgYWR/1m8fydl/WlhXEUDqcq0RAB5ejCLCu/lzF
Ok/6gCdHkekGnbGJec9/uqSpAtnGhn3jpwelvod8lNhy6Mbq7PhkNHyK1eS4G/YMbRC4lI5SEL9B
9/UON8msXQ4C+pM/vrUhaA1Kr4ACCIzadU/Wr1DC5pe0YzcEP0hR/u/YwKRzUuza03mnbK0rsoCV
Phn6FOi/0CZtenMFMY2UfbuwKpnRXbRKGcqUf92l3z5WEF+fjbcoaDzNJNXlUjTDxMOOtXOaHiAJ
FtfdczYhvJACSzy7OdHViT912zBgJ+b9XOLKAo7F3SuLlPJ8zz3u5OhMxRn/gOm+CPOBRSSf4WNJ
xBxAKS8LbXrwRvl/6IGd8LY6ZHPK45RzsdLAPMS/cgnWbvcV2WedCioaeUAh+iEQMBMBOAjKtA9z
Q2iAd8oSE15rkjfrN87nZnVV5iw4a6qnOS/b+uC6pC0wjDMQ41rh5ygxzU33WP0p6h+qjvJ/Zf8+
7FED5/orb4wxvEozNirScYRmBqfaqDbO5Tb8uDIKPQczAneamlH3zURwcGGxkm9SYeqcMbkNLPRr
83IVMkWxjAvOB93FJIbN8/prhHJZmN7oTpR3fgEKK9ZZGRM7iwIqp6NCQdL8JVmEAqNUw1SWhP2x
itnd01dvLQNL8OfgCaNpiMPia09VNUti5CiLrOUBupgWwZZOguoLbTo1aTMcBwl4dBMJM9a57qIt
YxDz/1UtuIN5xfXHKTMjfMm7gQawGHKWuSLFN0/CBP5ovLClf1ipeTUAvkN2q1zWh+EenmCOk6d0
z+Y1feDOz0AQjzgqLrJBcgmGuBuqH8FjCvBimtI2WqVMsiyrP/pKXu2jvUVxGX2kx5I/JCSmP2VP
EdI2X4SyrtgaQcGPdYxY25WiTlbpvUqlzNCYG7AV3AeUhA7RbyI8/tIuiPKIE53s5axmxUNXXdIC
IiIViUxzoVR+OphzVUnm+e21mjY1HpSbHGKxzOniofeMgW+sZC7Y1oZJR9pfUXx5dOHDuTt/KJH/
HnEsyGExYUmDui0kqFagAkI6CaD6SdpnyvDLQkU5XmlfKAD6P/C6SODikwfLRikdeLBT70isRXz8
zz0CyxXGupx227oifvBRy2Mg8vlITFkqckS0nHamyS1N4MZpVr2QM2Rif1njYE+3FPr+Z2g3J2J4
c9L3oeSZW5+0PBilqjrulX/BpSb7MHU9LOhOHnPxk+u3T/s8dFS58uXWz2Qmkgt7eQ5N74Ww8Gba
fbOijlfPjUjhGVVww5SagJJqsZqKG5CCPDbNSXCOldOmicH+5gh7rS6Syg/ioIqvyFtf4p8sbUM/
xxPsz63PmuZCkh/fHyUXVZIDHhft0OpbV+a9RuXinomPlpP7m9geR3CelOycG+xa9AG1BLEzQlZr
gmrn/QxdT1zV/S8YuH/5vnvOPZuzh/8dhu4F8dQiVL3/mdLTiypKfp/jylLrvPmsSLvbyC5xel5Z
Qedss2TDg90YRwnHzBlexxTm4mspGQmHYrQQabJw3XyVnJ2B1WyvPhZMQh06zSjfJnRqUaj/4SSd
BWx4T7UCzF3VTbXFdPb6+g0UksvbjOaY1k213xU/F8mwzGok4h7E8mx9KFpB9anZCSCkCaM/UArV
wMd757LDFb+AsqLHjg3idGcO5FAPnpN20tZywl18kZ+1hDRbvnIUK1pf0ZYEAWavGSs9WSpX3nSe
Kw2VtKRjwnfKA0EPb9RevfbQzUBWXEk7RKfYKgWBp4XnpEKXiYK3h77UYbXLW8DLiQg2R8Hb7Inu
gTxPtQdyZRiQ9DoHBGifWtPvZTLAbiGsoFqJ9UnMhQGOpgWHLfaN/GWLlR8s2broKq3wSKomok2N
r0tEVBPs3+rKeu3RdxLEWdkthP0H86vsWzyMc7pvqhcmOTJXOlR+J2pYp4rvPNgXCAnTNVvyYW/0
siGvdcTT+Btpif8VHD+kUB5LdK2Zw936kcLxP2K50L1Rho2uCa8EEBAKOnnr1V7Qw0Agv8Btv4wG
IKfXAa1HUSVt3SGqehBPmdfJ6fGqyU1Kki1nsufvjHjeCPh2YegarSUYQJTzDxRyRxKtFUtzwM3i
LrUOCbRc6HSAadz5FZKQuY1MQ0DuxJp2pfEnuwukSgR6BvJNOyl9BWdKpzTOJU6ITjgdqzEbullj
bkpAy7QWZeEklBu1Jr2wGwS8G5hND3pUAk6rUied0YXhRzath4NqCYKarPEwGaiuhW8KYQUDG3rR
kSpUQ/kz2qnIJHQ+OSklBcXJUNnh4BCUOnFZKprQzlpcb6qyskfgGWbg42itCSoypgYjvC6PlHjb
msxbAhCR+VNOdvaMuWFavqoXJmSaUwyszA9LMNp1MWoU61Mg6yt5bYYeoXDeIsSMKliReQroi5IF
Dng5xlmvM97JpgYHf8qgEG/t/uS97HBnU5pKqAHEkRnr0mbexYXnmufB403jfkHjZip3DA64AUCR
kPMB+KnkMzaX6FkCWoYFhD8g8GlO8YObCf9JliWJCN8EPQ+wHvXUj4BvEGGrHgSjKuIqCoyBp1lK
iF7NywlVf7Pt7Eu4aKri6wIjcxlry5/8f0giMI8A1CyCQ8Gr8FQVQmWLh6rwdHNuLP86/237wiT+
8zbThDvbsOV8PJoeKJaRq60qiPIYyoO9fzlF/JXcg96ElxN8eJYePzslnucR0wTMVBHTyRjzmGPE
4oRHIRFWFyioPTgBAYKTs1Zf9b2M7UuRIU2120t5FrZ7uQWZjrcPuw2Vp0HnBRI5V4JsgeAiRzFO
wSjDNMrP69JRMErBwgXHMGGoUa9sJG/omTueem0pR4PaIueduZ6kNxu2MfVMfDklmCdIL8BPEUBi
FQLl6jOPMe1klNLcqJ1hAfKnlLiEkc84D5OoorMiiIlG+BnqQZPds/u6GqVpRCkn/+ISw2Itduq2
q88Dj/jFu7DMHo5wugL/Yr/rd/kDom2HJTz1GW4vMLBIHSYNF92KoWr91emKRIy/sDNMxbkaxGHi
zjyE5N2u0c7DZ65UQCoU9Ky8QXlRUvpSSbA4hmY8SByze4f5IlRzanIeQI+jp7gnf+61+De16fBq
Z7e2r605tmY7YId6Bp4ndTjZ4ie2GlUcMXHvb6aWKoJ1PdiP1YLu8nt78xEd3xKE8ogmsmd8D3kS
5N6IFpkH0m8jnHV8wviVdZpdY/LVSFII9hCsE8JksTgwwjXk1XFF+SQMRgB0Y4wnnZGFqpf1Z8GK
nvUOt8ikD0sh+x1CdKH9XLt8ssUqieEvuhHKk76fvEZJEpSXfFB1Kwnes72SWnONJHstZjbKtxBU
rjDOjUBceQnPhybCvlKyukzdHsCVoy7OlGVUha5InBCYZr62SO4DBPWnEPXPg/P2Hs/2EGUhWFE4
YSOn6zX9rzEHA8AB54PYuZ5eolhoJ43uE1tHhO7ZWlWmXsrOxBH5k8S0bgzISmmlrAcuZAlyS+sW
SGnIxLSR+BYMYC/bZXi75OUV1sOspal3fs19NptKNBQLyqG9mLYir10EWTnZkRYXRlAXKARCC/fU
Ii7i/pXJo/3hgqzr66HBBrP2lNFI0+leqOSSXZanqZDGMIA7AIjedPynHxeUz1oKllYYkIk6g07i
flmljwvTUQ6XozT6qu0tUPNmMcuyCsyULCHZZvhSMOcEjPZ0MOUF3RW++Ad+9nNzIv+k0BdDp5Jr
PeyRU0ehwo5+y2t1xZpdGCoAvJjKntuVG8t0zSzCeHLHlGU3zc5a/v6oagd41H//h5WfaXz633jP
9TacfH9HvmM8GKzOvRWPTpGrIKiPgGGD9C0tMVBZDG3iSCKeEfO+fTV4ePJpCFfXkzMdG5k/cWCi
88lo3WGrEcH8zjTfdhpoVyGbkyGRg2gQaeitdRkwHVVieW0O2A18rHl1A4QLxVWY1QVXFfjX/0Ih
pcWcdfbCCgvAto2EOrZxATX/3WwC1U037dW+aV1Ra+j6Cduw+V20koTFHFzQbpda0cb1+mOWYGjZ
CviIfs28lS+hNhZ3E47W06+AY8KFsv6ssUta4MOdyhA1HIjHRnUJoccLdvkt0+UJ8wwzEb4wToI2
803CI1bo84n/35IKojaP0eVuD5h9cH+iHVtlyogH2lwvC5Vh7/XeSb9UAgG17CpIx+B0m4HnBlJZ
ym4P2wg/zi3xLVViADUzMhyYPAAFg1w7wIe/VO4KpS9/S+BmnqSYRcTN5jfh4nyu7WDsGTHKwCkV
YcCrdzQfDy2qiHq4vKKFpyBOgZlKiqol1JWYPD7A+dFG/1i4gX/+v18J5QVJ+Jsev17ppXisuw/a
bfwfCeg8TAIV68FZB3nSawcr76gYwSL8GDRiMdOnr/4Unbz68F8Gn/L2Leb/87So+CB1LaWlobZ0
KTQ4m++ahsUIjmMKfJbp7YtdcK+nFIrn2KP8lHxvct9K327FN1k/T1tB0+cLqtPqVp12L1EWCqhQ
uFP21/7WSHkG1gNkmJYVVSh7PRsTcfeI7lqWutXVeRM15IIPKTiN/qTz8vJB4li/kB0iAulBv5I2
chE31J5ud0os+a/h4XVj7gjtBsPmc3/lvE72flYEop0jqffcpZpHzkz3f40TQo5UuK/yJ4ZLAz8W
jXnKV0usUToblChsxcNOOIMQiEezrfhtD/Hlx5VIACPSvWMaReD6STYW3JvfWYHLmyHFMcAQXGqF
28XvciBvrmmNk6xprfjDSDFkrzr/qCPq4Q43igD3wwhe8xTpWMpF09MXn+or5+2UxA8FiNgBtmhp
K0JU1ql+bhOm9+C0hjWABaIMaK8UemIPrp0+SNah16rsISzreL+2g6Ui1TL9vDId1qMGzMqFGIX0
LEPy1xApCM2ZgtHOfLBdeSQuY2z6EDGvyGtyKgBNIB445RYGVPUHdPVJpGkusgCss7wqF3S0AW5g
kxAJxhi/rN6iMkqJLn+mcJp2qItkdi+HvnkeuF73UkIuKJy+nE2uIyZ6MROL3opQ1ZRYK1Q9dsdc
myCc8NlUNgQP5B1g1tT+CO9ECysOwWZZ/aHxxhXaOLN1yrO58bNA4qCSqdkt7IaScZ3VGn0+iUxV
O8yNIwggPft3x2nhpAbnSk3kzJuOFyGnTIIfzAA6WDbONN0QfyxZC6vSTrkkrfsXocQCv6mV0uO0
kEgzn11Sb8UTM59pg7XaCTbiHGQ1Cx4BgpWJRMNvlkHcQ/Hnn4T86eEl5ylFRkp6Sxq62mFaGWfV
IY63JsyGUq+4sRtdUiwN7x9bGmKiPbXgYdKZbRrdDo9YPyfp1jk/ASgWSTzXxqAKMx5SY4OSyn2z
8ri3lyp440dE5CbbLuW6g3Bvpl5kKsCjK5qO0+IF1Xz1FAv8QLMYrgyhG4NDu+s3iobeOeyaUUQh
5lmTL7Nv7S4BEEIDKbBTCaEHpRGVPrFCYvJrzMSQKsmwDI+Xwl29qxRzYMfKCujzBVfC4hF63POt
5zysCV4ccIO2sdUvjZUjND4KQRiRfMVoWcbLN2dSk+TNFChqaCbcHvC1aOTnkbdZYeFErPuwI3dE
dcy6sSsQfe7w4iOA5sdDippcq+607aqziRXfTqFWTiJOEXwWl7+MS4sA/QQ9M+wUAE/ZvcbTMZ+J
ZGMtbzzM4vbmxC36tCLHcvJSI4e8Err/479xVzJ/RbcmOsZ7wutQTx6r0a5XAe6uq0CTnsnF/HB2
mpLFVv9ocrrUrUB5qXkzD9QaaD7DxW6evPTugXypOrgJSTfeDvhHf6bpyn/HwdEeoL0bEIsEMM+s
WxSJsaM81w8zSS0gB7zxXHd1iGk2fPtW5aqE1gGcBWMLwuWFoaCYp0Q7Hkbz19Wz8jRTjg+Kp3H2
pM/SewySb1kOpYCLE+gCcJYXlkYqA1yr3lxxDf6gWzZLThPsR9JUuaLsMLQp8erlWB/pVvhPc7rn
RrZDOsUctf6e+SevFKS3H0eVLXr2smBlSzeyBe3yRaJgRuN5gghEaJJ1lNDSNdtZV/bL/VnCeDCK
r0c173y0exYloPSqrMlZMYDJmgZJwU3rLYFgCTGCUXVVFhvYnh45Bm7McS1PmTwVVljh0i/IK2GA
5r76iI1U2lho21o+uwIdobn3vn+Fe1VPHJrqsWARiUznTLhdHnGlpVISbQObCDXE0OTX413YIk9G
8uch0NYVDHjAuW77vEtc3SqUOlWbszr+Iiekc78X1BPb7V0Qp1lzbFj1zggnFtt3XZ5yGBQysCTD
5miH3/2/kA7G/IpmH2X/xAvLSXMB/AsrsvcTFu5ZBc0NC50P+FUreg7FsXUFtUySBCqUeBlD9cr7
WftNgdm2yQfD1nrb9TzYoFpHhffnyZzJjirZqtLf1Z0qSNrnUNqV/u2C1VUgv5R089QGZPlo8Jr9
4vg/R4d03PbpwwK+XsyF91Zqf4MLlyYSRZBagSao1GbK6VH+8SgWra2z21UFLiRwutJIr15f0vmg
PjdL/kgRhUAcjKiVNPTeDxkn+udqqb1vHlzdv1P6IROgkOvluGxNyk6XElCuvUWfx14deZE9iwpZ
8XpugA8e/rRkuVjI5Rip5SAX6Yxw4p9LUlsVjD7t0js6kuuJ6D1O3MWKyEzZ3dbrmIk2dmTZWjst
NPQ61JnRu0BnQxLaaCrhdw6It9SNcuZBFAtI+Fc3LJVRRiF9uWHAgBMjivUeO9HCJoQO424m/0Xw
6S+sSriCSDDt28exAc7Iz+3TzdirVbz11OJA4oSgUGQWRbTxkjR5riCHlzg/q9gfx8MreRBCizw3
0RSeCGo8y3ktLkM5yAxNNG7qehTQeVeNZnAMinSoubxVXbBAoHnLijJjgrvIBRUphxRuUIUXNyVz
RhI93x5PZrYGkQ1jfPX7da/E1lHgrgEl6SC9b/F3AEYrVHwXO7xGBxR8kML0lMMukR1uzHLe4rYJ
2F+j80EetVJB0TlEYgE4cKX56x8WV9c9c0ePh/ntJRlFsP7UCkzzKIimyFjqbVotgK6+llFC+Fgb
ggnZC00Iuj5n0wPYycgCUP680949oT/Cum49/O+w0qqeEzSXIhhYJKtBglT7uTPNqgzmBT/1DuAs
6OWSv5YylKCnAyJ8EDNHdYF2m2TAcXjhcmzj5sAaNivTCK4bGtt4q4tq0Xc6dMGgUUgYxGC8a4EI
+HA5ZSt/wgd5zsdvMwdNHfWgndlfZSZlkH5Tn2FIkj3fp9RFuJx4VkSmHv/6FfcLaTsAzFfRAror
PIlTBgmtLje+qTo8ycCm6J69If1sVfqC6Lt4w7gLvsmi94ISkYnD3XxwLDMRs3RgROpMNPBJ9TiE
KDY6hc1ZmbzLa8fl8A9P9KYrAXfyKBdjaDqzXjhulgud9Uso1NURoheTvMCizW3OcOHK9mBWQ3G5
DOH7HIgd6ymL1Jln2ZlS3D9SdPIdIfF5uZeka+FCoIK4VSVshrz4vAZ/TMjGhYzbW33cEI3q7dEM
7XdNmQR5JJXqiPN1grGCoGLb/IWtaAMUSXpmGcateQJhIFvG3dkzcIbqvnfQ8ybAL8O3GzFlsXpq
/0yyOiI9N5nAHnE6MvYOwNbDuslv6OdkFcsAEkEGZIKaEyKRJLuUvZP/sejbpQ2U5+mMCoeJ3eYI
K3i6OBxBefNRjm23vAj9wKipttzFuPdvr1tOjfmyLQLdxt2eBaRkV+1yFx8bhTLytzG24iBHfWAF
q5ALQ73hIMc97He0x+YvPsIQkEC4XPJXZyA4psJJXz/FHrtqJU/42jfY/XgYFN6io2qZyhi2535D
ZkimLPyeZ95RLcvJDa8cSbsRhRsUC7GFaAOeogyEkK+KIeTAsS5Soe0/0kduiVoB4YjZggly0eA/
Q9g/o5Tqw/86kCFSdtZ+O+1ZL6g/pXSJgTbVlvg4cPhKpjfzHR3rHKeW1sKEG9+92aIWHtZ0xAoi
SJen73obAvZdXELMRYPDZOti1pqBK3obUvBpO3S8yCoh4VuE95JkHuAN+jYnmaTnUcIAmJjKWQgh
8pSBeMOWR4yLH4XO6681gUfo21MZ/yzuPQN4YQs/H3D2vTRvo752hlHXdB4KSXPbGh7pqBqv3mGn
iu3p7YOg2jsTp6e2uKj5QXA6P/3XgKbm0ZpknxDOsa9+CpHlXvNqTW0kU5/Uc09smdjZvjRlBkXb
Pi+gh0mEx+OT9b5Gv3HI0JmdicQhmQIzS0g1Oui7aXGHobQo94rkmfo6bvUF3lWsnyi9muX/JFX8
IUk3f+E/mwtWZ1+VzJSuVux3PD58Zx+rSRFUlt+2rMhXDilUJGbM3XPm7ddProP1lyfpd3VaNxDc
wIlaTeK79HUKDiNZKANX+nLENemJa06LNu/dwcaa6bq5BZqw37XdcyaBQSsmac+BZL8rGODAakyo
qdWC/PqbeDh1TTRNEaN1mukKdpvBqohJF6fN89CJ3s6ke0o3M9PZXn+XF7/UYSkxj9pVSSDkfZkE
iddkabCNSEjNYlrTogiHJATPhzIat4j3x+Clg3k+XMHb+c8En8J5hyUx050Uxt5v5tu8IiX6MB9s
DMZiANQtknICyORE66aBYAaPNQzmWmj3GXSmZZy8v8k53G9olFJiC9cY8OOKnFSJ0rWbDRHZUdnM
OUy2LjyGos4FrX/w/2gaANAgTs/AsVDtPi3N5iQXUh8tm8sV8juyDToRfFu4SEGS4YuKiC+w/OQr
MsPMeB1b2mSXLaGakObChrEsuVtgOxoM4DaXteNWSlRGU0F5CayvrWK0PSo0x0iqTOvOVf2DeUy2
gxcqkeeaJLbel8hQUiVodbvVSLwuxAC9u2+6m/6yu4033tVzr5DzRsPc9ApU/i9YcD6+UgAgY5zk
OGlarZ4iZjH0mUzwL2rAXwFgjJ7bfHm6cVUg6wl2kbyWRBmds1f4FhvHtmdyI9n1pTRo71JcHHsP
ntmR4GgM1kdbPpE+IjI+lkWVhbX66aYk+dFy5n27IMFvOHaNePljwD8lZ8k1/jsF2En2vh8sXx8W
QEqJRejkYRzZfUCPFKfF/u6WCYYeC6H+2lNeOnhwGAhDKI8RsaWBeJr8aL9QSu4NOKLVXQ+lquAB
37ky/YgGoJSZ/er3BaSzISybuoGfPwnxvpu+DGxR2AdLPOl0hfTH+/bCpv0ZDzyVG7nRDvpQGyQC
iMOHWlUyYeqBy51gLA5vlSwPkgbZ+KfanbZhluykLzBHXDmUJaJAUr1SCpRa9JwS5gsusQ9oo+zU
mA4ksfM7BDdB1L5lfGuq1TLBlTjlwK3Hs4lSZAJLzOOQh2K3SU5n71eHYE/gXcL8z+gj1hGVm/DN
gQo+GSZ42vVXYZnTLAN+oRMekn+oohAcsv8eq/vP+tPl2LfCstcVYfEOGKI5FjPyrchrNw7bSOBe
ijOaBaI73K3RWuMQkW3BZU/p/VYd0BIww8+r9sQXFLyi0lOCmdMTIKfBlZ30eNjLrvd9Qgf3OZdf
AuGa5QBvbrgEPFnlxXuaI3q/Kx+fB0Acg5x9giTa8wjtAbp8BIhj/0OTSWqR+AiD45KC2iRmrur/
0z3+pWfaGhH9SQn6I3Cx7oDK5cI8BcAUnokb56mqrALqu0sDo72h4HhvgmG/SfWIEFBLJgym3k9O
f112Zk9U+74js6ksNOUzL28NRmlSPVfSe+vXXnqRRDKq6HDdVT3ys58CghP/k9WKLG+koC2LcPkK
ANKbzVYW2SeNgVR+m6YTo5aRxP1PRlCDjma63ItEYER3GzkvdIjpgPHoS/DRwQH14mzH7Hl9QyYq
ha6ICRMpYrm/mtFYX3YvUcMKKej3YHLRuaoP182wxbUcmzS9IFBG/V1OYwMhEIO49XNCk10PGEQW
hHDuTEMODA/3z7eObzqbSXysQGnZkYL1EVS5aA20M0I6n2+k4EnhRmZu8aOrKkBQWtBsy+SjegG4
UeW7cYhWk0jQhMfA6M5ysfn8RsxfvQF6SkA/z//yawfTRspJ2FZh4dtr8duYMc2oV6EOuhafqf+j
nQoncVcK+EvaKNYP2+vP9qm2DdyjNYxviukfLblN1QBVzpr3OG47qdPhyP5jSA0YkF7RDOyd6FQL
82L8IDSdNZ2qbyIV6xvsyWc4aVUWnrNUYaivLlW+1QLfxdQEp+EijhC3xlEVLMyb/AvviSt4d4xc
L5QF7CeBcN5i8PK25HY5iuWTKZFtoHhCOvfsvgUUiNTqX2BaERcUBcErtuYDZ+Q+bvAZvKZLW/N2
q7+EHH9Vf1er5PkzQ3xtiQNhyULxeNNeKQ75LmmwVvwcy1/21qhK3q/zE7TlKezZguY2cWPTjKco
9+pXFU14Xw5csuZ6gk7bR7hJeqpyMusvHMGo4s5ec4n7PaFzh4okLLa+Loix5UEjaUVhI5cXoD3+
y8glAtPWuN/R1JJatjF2+YhYzJlJPsQ30D5OuWrf+GCZrRLKxjO164xW3HqUC6cUOhxfCNIRaWzy
4Y42aEhTp+dfoyVaoC2k28CT6Ugd761XgLFaVZrd5Ctm8VNFyCbrzWjF9c4BLHw5rotgoD58HDeC
naMH1501ng5RNm1FF2z58t7mVV+/IDI7QJplNvWCUe2gbmJvVZAXB4fXgDYQkkifCZm2deQHAz+T
15X7UgTdajFDPklxON7uAZ6ohE3+WQABdDGAkjdQ+ot2JdTg7rfmGxL1UQ+nM5VnitpS67umxRPz
blOuJxJvJqEi1U4CkgvgR7nhAenJNgpUWIw3jWQKO0HYDjeq75SlKToPRpwjafl4oKjt8nOlSSoj
pHb3CjNfdxQ7P7eJBR7D2WZRXVF1txXiG8uqr1ca4IisBdHCXijd4kMbUDUAkU5c0T4rmIAvuRZ0
MG09U8ycrtBdRrkIzsSFVtVeRgJPe5t/QG2ccgnIWY88fLspTpfLPLtvdoEP1e5JmAdHTY/pEsqA
3KAeLHHtzvUz+X/zuUTSHLA2dN1sAAP0pA59utpOKemon7H3pBmVF6lQF3A7rXwP3kFzHOKuhIr8
Ki6JVvAt2xqMCzkktghWQqBWDPUbUrOBLTXb9fZzy2AJ5SITCAhT7Jz6HSaayP/1Eq09boViIrww
KDkd1aPxPPVpuig9l7bPHuxBLNhRMdvIcuWyEN+hqX2XfWLrZNx5RsbMavUlgE3W43731xZ/qG1l
TIjqks6sU0QVuaRiodjiS8Sh+3nJ+LgcJYZaMLKMGKZhQmq6w6k0UdoYXxQSSBuGc4qCQG0SFgaB
jtFK4e62cNB8QjEXLH0L04E1gckR752X1cRaYlnNIHw4ic91uN5NACXFT+qI8jDTrh1FAzjKVALu
Yb+h1j/jOBRKstWxFdcdxHxe9pRRX5O6y+spnueDVT/mGGMiXoA3MocTFxH5vYEMAClXMwTnKEQe
YWXhfzQLhufcCN3yR4hH+TrbFDRdf+OVYLCGiX49q+KYQg/AiZc2Oj4okI2p6iMZbUN9A+gP7rQm
9KwY2t8JrHf1ndiMsAfDKRqFBJO93LpNnvZ3lk2wazlX4X6vj/W3/XO9XVN62c0xZNcvIyiuXW0y
3TLdZdo2Xmh4vSDjIcXKK8GROm3H7fmNTwhEuPpjrbqFmw960XBbvIiCRApZKW15CvQzMdSrjNH8
cjzeXCDQ3ReORoGjGXYXxYUKS/IqTm37O2Zu5nYhXJK+zmCMsglnBlaK/d8ICAIQ0D66IZT6t7Bw
ohr75ouyf/SuqkTS+s8ZxLlVPzgHOCNM/DIpjQXAeXuFZilUD96wIhUOIupTgNXsPbTXsvcW5bUb
h4SSoFc1PAGD8AsFuIoBG2YBwZLUJVf3AMkzV39AXHJbHtSHuei0sbLUufCdp5BMZFW2kdH3xXgH
D9CRNi60eSjDPHV0guHQfcDBF/w8ZR2lJkNnk31jIlGNa/FOkvfKbGb4FLJVoF8/cxwEcuyxzzga
StqET9FS5AJGFmHuXCeJsGqJwUNWTBzS6tV4j+XMAmG2xaJ5wlW79sSn8kIQlyqQLBosP9aiRIIZ
F5QYnKTICopT1OPwvxG+e06tl2Zp6InN1UIUTTy7ZURabTJFhFlV+olBzD2j447R6LJ4VxIS9TU8
HBTs/+Hy2aKWaQ0QumcuOoHpZKXLUrMpOerdw0TYGQheokqRclzDAmYEf56uqtfDb5RPqlQRO9mt
grkcDshxtaHVnnjSDNm/AEPlp0dRr1kbh81i/4tPRSZUAqb+z/5vI2UIxSIoLrn4Krh4+BH6cqZj
G51Wkhm1k1V8U2/4GYplzhdVf2MlZNhM1o7ZnYggsMZheiR/t3Y4Z5AR6Ph8nKVoMVJ5tXmHM9ZI
zP+WxwmnYp2jvmuMdRVeGaqWlsbpGpozbOIrOSU7xgidmGrCVivzlSWl31EJ+EciJKG8vygUEMcG
WmSLgS920dMfcKfEDn65guDsldDP5FlgOhSibSEBqJhOjXK3kgGxKkT7xkXqsP09rONvuxXnOKIH
nyP+WGf5PBLHaI35fHzFQakT9vVg8l9SD38SUqyZsiWbpvwWPWflFiei0YOHAgWE5+Ghrb7cgevW
hk9pXokuBK2PjevDUTjpuVhgkVtdj6asf4fExLL3ORE6bkq0lhmu4DPRjaEqcULEjbm5y8CBDvN+
0EoEefTyfQ1huvE13bDZtn40BCVNzRHUe8gGYHl3PDuUkFmKuO91ovocUEo99SieXO96RUEAKZAa
h4p+W4dzIoK+iGhKZniopDouOAL4ebxwuTcKFFx/kUFUoa/Jrs3kEZ2iqnxp9uC6YkPYNgo+yaS0
nCoI5+lQ5jwVYQjilunrdUEJHM/Ke2BqZWVYGwK5T1NwNVmgfRSzCHatEJ+Gnpmx2gX/tIW5Cp6U
DIJfYdO9NPoD4EpmLe+50UPDGQQHSnmrk5AaY/ff8vdUCWQaWtXJzfQRWmtTyQRTHNXnyeAc1HBg
lrm5HBmlfUjw1YE4eV+n+8ouFxhm6H/3fcReM7AynT5uWZ28rfaSaVMHBor39DIqXBJJpBCw88V3
P14d7gPlR+3Vw+HLpD5np3IR9F4mpHicM0m1IBZQJwdqgc41ci5ximh7DyEFE9toXwLjmKQAwv+W
tnHfyW6FJY2WomjKD1hdmFCTtWCGv6jan7Oe0++6ArKSqaEol7DW2orsjgGf5Z4cDRucuhmD/E/v
lS5wfi0Rq6n1ppoMvJaY7f1glz1UNHkoj3JAO+/2yCDjmnCX/uGIZsozOfe1Prf1XuY0aBELyVJM
rKqdWmn7ZCkKHebSHbVqUvJSePjxe1UoIoNF5pqzFtOQaDfE5YRJNJeof4FTleZZ+A9wJUFt4GVs
wLlBp53PaJAIooT6t2sfGIESuOruWvihHvxipBfHQQi8dLwNspQJMLIOva55EA2XJDa8FdR8Y9e6
5xFrXw8vTV/iYLC251KBcrtvDvHVXkscEDQdEPHDenlHwU8QNso6FVBxKQ1pu1mktBPoWyJDvfbe
o9xqppUgj0KV49y8fU9kZUSduMBogBp7BcUsHTLXde/yqsvhOMEv6FN6bFMZJJEh4O47IF5FHKpW
cgUV7SwoTgP/QrQ8b3hcR37E05QffR27Fr4d7HdHFKo4K88QbxjCUpwxa3Ub2b/Mvc6HF2WVY3Cc
1NFgMV25pws/dc1gQF3IUJvRur0ss2hNTM2CZV25aJo23CDSZMpLT+5TVEdbtBz+uU1Tl5/GwLlK
WFFg4/gIgmLoAuverbVAlqRgu+SOPHf/i9QG68g/I6kmxVbhQoJimRoko249BjhT9K+hip3V9VWf
gHPmxXoOtxfu2bbiYeH6YG2POHlzHSidzysHWF7Cyekr+pv/kCbm7QO4gWn6NzQXJ95yPigCdpI1
JfPa39/Qc3HnToGijeZvMKnbupqY3tICJQk2kb1atHQBisvOUtW80+Vw4Rhhb7YWwv7HcIR3i9xn
osxRonmUkeOm+BcPSDNrc3hjXCSObT9ydUjsm0x7pR/385jHiyFEr5wJGGreEyrz+TNTyTZUKklJ
WcQCGYLxwLyOJliz2wrtnz11Zw56574ihlJQeCG637AfwHOrJdvWBiiF97STMhwFDoIEfUk43bl/
RwJS4tuhy+iYhCQu6/7kLDOrqzLodwM3YcZXkdNPQmJIpm0qwJj/yjU9WAtGKhXXWGT8DLRTAjqi
BNN/MeKgw5pk0kwdCo55L8MnVJBVDlLwjj0+q+4R15WdQsen1CEUC827byOzsaeW6w/3ocBcJmR1
WR7bxZM5twpYWlvIn/5MfJTnhCUIbXAnmQpvAjUlOZnVkT0YFSpxg2LWxdUfTkKdtbKv7efR+pWz
aH1S+yLtrDaFP3VAFZeYoOdiH1wQwNSDHnLbhgBYgIsHXprB6Hlg2P9wDDvJPAhLFuo9V20JLyw6
judTUDvAYWKjm4zsi0OwtIwXbj1wXpRWZdTo8HJUx0V60Hs2QnwNsHkbNMwlBQhVl9u8vsRWoIpw
8j8ppb5fvo4TARIsiNIfSeZM678hQGC+ooMezdnwra0/WaarOzAjxxrkpIluD6bLMQGtq/5RlzUx
ldrCdsTjnp+AayX7KO4iAmxaoc7e4PhzofY/GevB13w7XboRKbZyfxRR/6Rjt1JDwHTz1SM7AlqN
USirkAzzTtz8TkKBSIHPgzS403YZUOoPUPRP2sMjnuKXlLL0A7/8eIWses0g3bRI0IDb8OOPLjcZ
xcamJiVaA4B/x5Sicio7XTNZ827EEgsezhnyqMZhdktgaNve++gDw7Pv3tGyKpxz8cdHKgIKlFOo
nH39XIhIafNrm+tWDvb0zt/DTzT44Gib0jwu22rJE9MfV8cHykPa4b1PMiEZGsDg/fYaKzhXsLwm
hMT+sQr/ZtYvhTj0YaYqUbUYt4O3UcWTkOdclkZz8ar+XrSk/Iw6D6fEfVNK0XaO2e0QbByC729F
6Z6R1Zi/IU9p8S5Bg9UJ0B3lD6UTV6Uv1o4zGbXbgsx1Dqi6JSd4xVe3UKzNZXOv8gGGMCfyxJzs
4MMOBYuOdKbhH5wgdkNxV3NsWTq8Xvx0Wmpg0LiT6nLoI6I+RLrvRuopnKO/WJ189xSX5TKEXsY1
LWbfDocZX7oDNiga5/AyNoR3DV/ZKU3ZWl6ghc17OCOxgfD96HWROXZGStsnCw0o+e4IqOPPHr/z
BWbXhLtzr3qfu7bmaoMK4/1FC9Uyy5K+45MVWvBQeQ7RkBMqLXohmcebWXtsvXPbGcrCaOGFIDQc
GZqfBXOMSWPIc2of7DmdUHb7+IhNYmUduZ2U66woaW8i8AApUT4gJIT0FHOGecx3KU6age0zcr6S
EZXyKnJyNPa0zHY5TjCQ9XBxYM+QLGpiYSKDxKWaqHi3zruWKMW/XbdmaB9xpjtJ3ICBE2cJDk8t
zriEHo5mTldEvZTSVTc64F5jqsRpcTL30qZQSztsxQISOHyOLGMlaob8ByW002s0g4xpdiu7JC/5
yCbcSdZQsbIfd2QmudCGwyta0jJjHqSUbF9LigX/ycN4sBZY24z8KsvPqwFzmkRN3QxUq3SFsmyw
e0ZzsEdxuE2lmPVu0V6Y3b3sFs70wpgq47jd4uqTdb6FywJ/Jq+lZncrpzGhHu/dKYSO/yIse40Q
NFDWjlepuM8Y2E1oOPfNikMTskOw/cwW1n+G0pz11uTAJk2K7wPSsaJmqkTQPsXfMPRV/usUsWn8
45lzi78/b9YPr7z0hQk0hDO3tLZpzhGiOzlb0Xs7aABQE8BalSk+87yHxXVHQr36x17Y6o06NmsE
BT6qPhebS2MVdIUHDJOyJ9B6rASiiQyPx0Fle6YJzmVO378fdtThd9oReyiMAh7OWhCX1mlxONmC
w4eul76HgNhNLgZUnUAwfBx2/UC2pd6IMB9t4xkQKp+u9dza6xJiXezqGVoa6KDrwDkt2h1LaEtf
f6xwN2b/ezOHncNZc/WW6IYkS0wjYga7tvJcAGkB0no1Rfw+6Mo9ZMkXQuWDzAbxV96whUA9b3Gu
YuAT69V8O77yk+VVLpOvYhtwzy4PAKjIX3avIslkjXTkGeu962jL+hQNB2+7BxuJqHp6xEzDW7Rn
4nOsP8N16HCSmHYV6huLNx98CNSA9qinaFzVv/LYAgw96Rc0gmy8LyoQy1z2aq7XbeTzGwRfqPp9
dpQHZ0G+C4q0OVGMw7Cm1M2LaiWj67O94kvWaGg+9wj0MPjrjx3wRyQzu3PnmbgiPkcHOS3NWrSw
hQQtlR3VsJb309TB5etYYRf/cCVCFNdtdTsu/en2s6w6M+7MICoFeDxhdFbbU6hjrnZ5gWVkQUH9
strBKRDdH8lw3YUapQ0oP9t+SJ0aZoH8dA0KZS/egg2X4XmwIV7R/gmUPU6yJgoK3t3fzfAzZQGI
ezOoeulPE/qNe/K6dRPpHHwfidyUyYAkoStSOGtdjv6CAngPV/R5BSgRC7KPYjDe0KF1eRfMu+pe
+5oT3Ap8OG8uE8IvkyJx6N8ZES20I/3ZN+ZQSbKsne+pKp9o+mHgzzZLGePTbuoN1aluat41EOrz
5dXQDCncXlUI/jNLuslVhdk8iZJ7vT+vTJwcqL4iyK1Fi0KEeKW7vmEusMhHxddYTBaSnOcz7OXw
qrTV6HxqW3GlKCQq/f4mEMTSGhWfKuI7A83suCnXDhM1Gr0zYSeTM5g4aSSDVxv9EfeMBmV4Clx+
ibAi1VZIe7J1xQT8tt5tQPziKNHLTnN5k6aLpe36NQtbnKd0e6xy4GvcyjuAxCE5AbrXVDgW/51x
nZ2D7XmrIm4RlNOH4y2XoD420ywfvpu8rLkQ++C3Zt9hOUZKE919VN+vznUJGwiM7+WK0c2ayRW+
jRwo5/lg/jaHkncQo7G/7F4GvqNrhfEREk0DiJQfxWBXRCJvQluD153UTxE8G3wGrt4sXtF3DiRA
2J5T/UbbdxNmFTOI4bNe/wAlD+bacV2YzsbIFg2rgiwW3c0KpmS8Tfm4H8Lrf72WRLCWPu1L7HuD
FMLY9h/GAH2ll/kfyA+Dz22cW95VfT4Tq+J+J9puO5AoOCuSuxRxrY0qO6LVDxVOHRHPBVgUi6hK
WVz1UHwzCAeSszIdf8mErfX10cmN9qAEjmCcvvFXc2zVBnCsUVq3JW3BRtBN9NxWnXa3iITn3pmz
BhY6R4NaAknJaFp0dvJYOGDQiuNzI5aDNpDEFlSydDu0P3OgAcnSlvpdS0ryEq7MuINx4SjYgVnB
E0ZCK9KpPJFanyj7/+oswWcwgWXmg6BP/Z7FrHJnmny1mLFQYLD4BuRyGz89jceTwY2HARIJdFMa
18T6AORprPcgRUmx6MjgJIMK393I76nyXJBgS2tVMXTeKr6/RkaRUyvzU6WRwsNj6KEJHRmtVGa3
e4vyz1ZytS6EwCCAnrpG5pbjAWbOIcaZXSGi4Xww9b1Lo4sUOE+8991AQmRPkahyQhulr5RvY5Vz
LZcsfbInNSz/MhKq2fse/j+dHQsVNMwt9UCV+bVXT0RIqpLD7Fb89R+3Bi1WAORxpALREmAIXRmY
NZjTQT2/qxi83rflfpfAl6i2lymMCl/78Mj69BbzFiu2Qwp9MujhVCaW+VZ2W7/KAgn9u6RCS6Tq
8o0zPnxriuMqLjA6M4x70bmzLHjSvX253zLQvKh2vIUySt4k2vMUf5rYpz1G7m07A0ZLkktbm3uU
JPH/R5QWuQGF/S0YiXBRBTQ9NUTNiyNykbsfE2BBo6IrlEx6IeYmyA/Om4Ge2EKE2yMSd9ENULES
zxJGqTb8HiaOIWR9Mbqz4cLFwELl91QqsACxkzHrdurTQLgvPY97ICQy3aZnxrZYOGh1Ejqg2Acp
Dpbc/pKjpSyXlOvgmMDhO1F/cjGs4UCWc7Ab5MmrC1TD2fOPsh+xTSjErOF/uk1RLrznj9FZbO9t
6Ho7MTCNqT6QGwgSKHrJiJB2JhCUzzfZ3XqUhDhh0HMvXT/JZYG+syX/D5k4pQFxvmXcSZ3DANh9
2lQ/zp6bKsani8cQ6lL/6fhwQmq7I4+dGIIg2yc7LfAG2Ba45hiczluBYZoMhiMCFlykKxG0Cx/4
G2m/FEZA6Z3o31X05IWlAyJ+yY0QRfF5SUQKfUvt5x5bSwu2CPOdMAV8168Y7oEgXW4yR3RBNk4l
XHFmGw5C8zgk/YT0aXBV9IFg02NOt+urWnBdu21ou2t/p/5P8cN63NxWCDnyaDQNcvQzBbqdeRZN
sNxsxb5lJzCNzFFj8nBh7+54WVP4wUbO6fjTluzqKZjfhTiTdHTQgbYhhA23Qszms2Q1gZVSlhqZ
5mW0Z8w0UzZr6H7I7Z3sCJc3g2K82gnilYAD8KPdakaQd2jpqNj0IQJuKULw9webLvdkyfV4uwjZ
is0uaEYV9oHzuo0gRCVbpRgTkuLnUqzpXtFh+/Q7hKN8m1AgLGj+QLOLFJGCE4sN4mPN5mxJ/Sk0
/c35a22+mqEBJD6tbhs99y+HlAAifa1Nf5BlD0oLaSqWzlBeUfyVmhXTJ1zO1XsziKY2pIOPvhY2
iVkM95tAcAfmfevMCC5+a/IPM5IaZIWF+NHTT/PnACQcgNANhO0ScLcbLvksv1BO8UxgZBXoWg2z
xMKzglaNa9ciOtewaWr8NFzGbPsILybz+EhodM9RJXqur8lx2ZErE6SWKFLdqerAvH35gdh/cutH
oyZPEqKqqS8G9YM2nDG+ohsc92s/ZJsf071nG6LBkEDjOn20RbvZNE5m/J/drfceXXjtUmEptW9T
Y4Nj9wzlBlu8+IS6EoQmWZVicT+8TJN42oRFss45RJY64+MuEO42Q44zi674TXNqWjOld2M0Rahc
tHM/hjiHsPg0SX+G5YUhq5S81cVzR2eL0yrrvZ+32bPJmPXiVG9QRfz7eWQWmtg1a5okD4SMph2a
awA8Q9Szss7QrNMQrft3dsxUu16bdBjHQIAJnBnTwyFtl16oBbINz8LAjjEiHLYHB0dfcUZHQGkO
kggzBoba13QW/gDAo2W/BpVJ8VTZt34UlZMVXbyBM+PB2aZ9wmWV4cyTdGDNUkvbvCFAp+P0HH7W
XJtLzYEl2MVpvkdMl5V2KSX3q18bWFMretAtCRwJ8nutVk+loZO8mVflP2f+B+Kf8X1jnudFFL8z
YxoiQXqJtS5Xg0aU45+aqy50fKgEz0Nw/cTcZX5bfh8tZqBgeMghsyuaYW+tk5fKSigZ0+yx5t7b
RtbCffXAQVknEFZiscZE2JXgRYP6gHbqCt2VsffeTe+rdWhvIz5wQAuq4fjJo14/uAtIxswZYyCF
8ytGncQgrj86DUWFxL4iQump0aAW4ILwLaEApCaXAXIwvS9SMZNY+/Y9hni7dDDRpkxZ254BX70P
Xq99y8BDMaHO0zt0Rps2xFaYM/S4CwTIm42TtsgA4E1UEPPozwreJbyKLTMn4EEG4HZmQgjB5qs4
pA1+BeVJBJZM7KddRlOdf7LWrik1b+mqQh1pEEmDhDP7/5RdFDJfDqfS5qExAeC5ZfBfNfWxNtv8
Qxfbzi/qyk2IGf7fs76CcAi5M10mvtTtG1uJkMIbJDZ/mDCasHHeaqpubG6ls7CghoauEqZOWR52
MktjePb4RG1L0FM/pfDSLS+7597FgTrrey4wcfPsrV41T46cWm8mxaKt57tMm3C2+7YFebRTlnxr
Y/nyTGWGBB4S0zHd/IoJqBmNa+lLUX3WjvZaXeYa9uujovTVp08m3uwC95W2FiuuQ3p0w6B3m6IW
mHd1mfIrl2GcLcPsav4CZr/7SSg44SevZ7hgZgmpFIhPwndz+3RyjIdwYMAjkyMZjnNhETHF9NYr
Y+9kbcyhTVv9WYrMzI/SSuSPXq9f9vRUFcgfmm6rfHyTeTsxBpF0QzEDxGRAq6Gy7IcdmKxMNqMD
58JQ3MzguJTf8m3iucpe5QWnoP7zKgzVX1O6pbeJLBvxLQNTs5ygo4S9oPMkHBYKlc3w4hX2eCj0
Lkz0AIXJ9GFa3P8TF1eJ1qo6z/bg03LqCRox3HxcV6PMpcDbS+Z1NAjrX0BGvSCLY4Vs6CjcmEeU
16DPvuOBHEyGKR5IfxTVK9zx9ZccoeLWXK7iP+D1AhcOBKz3UXmoE/hEs/yK9uIEw00EYHTFR8m6
lXLXuJQPHRHAwsVlwGoyRBz2ddxq5dGVzN59ZzvPLcVt+G/LTq3DtypECE7l/vbC9i+yvaJod3MR
JBBFsdd5ohweAnrExSbmituYA64maZ7T6xyyk5cjJPqW+206/asvRUZlYeu+ddX5Z/+GFs1PiIx6
S2LATOvVQQ9+5o+Vp0zdBtFAlvTyOvYtcf9FeB38Y5l71eevRrESyEyNXsmQN4W6lTT7uxc0bigh
kGgXsWwT/rnicXj2USME3TTNlzzIFD9AZJBUHJvKt1uEBWLNwxaRvbxEmrae7ClG32+ypiTR0G6L
RX1JpM5YoJWPWbxSj7OH9XM1mMplw6DyHWtR8wDvdooPYhK/H1IwznTuBhmABGB2DBrmlheGPHPM
2+EZ6LpBArnZGkEuVAP1k1OSDGqi9LgjfMQDm/bqmaj5kv0Fz1ryWfGHVfBKZ0gnyQ4UHmAcbnjR
d163yobMimOEohxm/P0lFB9JQFV77wowfLLzeO4J4DsnP7mUfK3iDwQyAYWOW8XPrLt7jOAkOMkF
UAfD9XRfROumDnuC/GMz4aPYV4WGLmS0HSMAwl+pl+N560g9HTJ61oQwP14Owz0fTWXHWJFJ8jvz
3zE8Ze557Qc1YEiddFgO6ILV9uZOwBf8jA7nlNF+6j5QHhmcLBHBKaKCQTCOGeyklor1ierU1L4p
vDYyhTz/HBEgsRASVPxFyCLcGB+OhPX3MKRuBeGj3JuOs7oBa/MWdIBFggpfofFL697lk0I244gR
clnUj5TqaZTMIbaJf0j76yVcKUE4aykbyrA+jKM6QFuAhhozHKUDMvz/A5YYI+l/BnK+8E9NTtKB
n2RnxRas2w85zGkb7ynsqd/Dqlhlbpm+m9315lTQOrplPbMHP2urouxM9xpyzXkEpMAmjofdxJvv
jdriD1PDV0yFQRybz0Q9sFNO3pAfko5iP0xCFTjauFiTURxud6MYFxSnwWJBbR4IiLvssvSkPNBU
2sq9FwCMlQFsEkZOoNZo/Em/v082Jj+E+mex8a0KHujEGoDPWroO4AYKBWgNLIK872ZHTaD9UdFE
PKoV9GzIun1UbPhNNVBYu9j1tfew/sMNK+5HrL2uL43az3PkFbvDNIf6+08l1FyCR90H7a4+N6xQ
4F/xYsq+pTdI3Dr0CCcchCtAucXMwBCrplig9qZcfIEVHZQCRfdoiYdWABUvzSI3EtRTkI7a3cxZ
YJ0I7YuSxM4KQaEw10/CJ8A6/kwZBiIZrWbczAHLUi+NaGgKxSuZTWNyVMazTMZ6LTSUJL3gIWdO
9hAtlLu2wEoQa0PnHNCcDTtlGPWQWzSaU87eV6u49FUFgtMeTpbOg0qeqQ3PCDTyTeqCOkvm5316
vyU3FR0BWCzxutjlPhEcOwF7ta0X2KpTZh+/+MtZk4wUudatk8kQx76CKN7hYKXA8FJ/252nBXr2
G3LeiBHF/aaotG/NTxKXZaxuwAD19I5uZaV+7A/7mxuj09VygqjrOb6PWYwh+15HQ0b6EmhgmAQf
Hof2RVMp1g/CWZ8IzZ8Uy01k1U2++9BYh1wpD0w9kHwiIbXpJrMyY2scL0gLL86nPtKJZQ/1nzSG
MVw9LkOkhi2x6zwvD/gb5ruhU333U5F98tPL4Qp2/jtXqG1ZKGaERS31BPxFA5ul09+WVISiVF0h
GT7blWBOe6UmmVcgUxoNSWdykKpgrlx71pIH5Jw7pXxBZ8IZmbSt48cIjMdusD4Z50SqensM73ae
8VUMYXRfTBFlL+YCkS0hRif5n8b3Jcs/QJwrOut0GHhRG/1WmyobURE9yrTP2Pwy5VetVTjl5lR3
fo6x6fMsLb9VpVjh1nKv9UGVQfpwvs9l00wfvePRnqbcPTIKP8Po7qRlvPlj6P6wLyZyxfb8GVlR
Ywjr4JtDFRd+WQGvXNJj8pzE3KIvwLnQPn0tgtXNVlRITOob+UVFko4ehPttEknTykr9apBOX+7U
T/iRknC7oppO6cI74KdUQvfd+CeEXWrS7oMop5jgGZ4Hv2ko5FKW56axy23pVR5guPGn3BVMCCrk
GCKKFjfYc17wzcF9gQrnmtvtWRvszg+l5G7JaEtxIcOVZOV+wXQ6wCT287yAFlhBeWzTtJmvITYd
xHjXIrOLF/IK4QWmjhBnVuvbAU7Xj74E0HgIIMUy4YRCKfMcADTH9lvkvEdQ3MRxZueIxSa7ZUtb
dlYT3XRZgNOGg/frw+qtaqO5Eu3R3CqgJxZVpNCc0WW4mTLqQYwaQF98TkkQLV+VdVujBFLL0m1g
J6nQABRYgRyIzFMlPHqmqNj/fj0LuB7+puOaogwvtYTB9eGGmoroSSO+efrpp4CSVEqb6euJoIap
CE+cHuBzwc9CcIzrz3O3BfotJc4/M+Czlc/a7Nfb8VxTCbtj0BFXSuSUaJROc9Nzn+WN6pQQSyIT
wTEbyKMkk2frzMzXT+KMS2YGuMwuQH3x/mh6azSCQNGz+94lnk9mD5xRQyVc8nCgNTTW6XG0tmVo
llc78HM6FJWkkQlrolBB8sDwiUjYnC7TWhFEfmIEjjH5CJbxvpk5xcW9i/lvwHVYQXdBWfMLw2aL
IUf0MQ5k1Jyp8w0X4qeWcoLfHQk+bj9hbERvPtHIa92rusp+g1TAgUK1xOG7eIK0pG5km079n0yr
SWBPs4qmBwD6WaShNX9EJUvceBdNFgui2WRDrO7EZmQN/idYMix8FXCcWdS5lwCm3WkrbdsYSXwl
RjUP7h6xnNAoOBOxI3zE9F/yhYlDNGEbIBblq9UPfsJ8kZslqTE7ZS1VhiQOu6GKeR7vPhCgKSmC
0eNzxGNf3Ga8rFB6r8iVz8WXc+zFFGLy/iMzUVPrZcP/9ZihIXgY0CHhDllsX6DMVCSDf3wwMoqX
pAR9syUEVKC0aVGQlVsPaSJvL6/M2f1VNeJsvtuyi1DEZm+I/oK03MYhrW1H6v8kmhcfAQsz83Cy
Z/kQ5GM34cz583uX8n0NPudnCqB4HYDsEvhgRFDq3mId9CG9fFNEO/ijVk1xRv66Fnz9FrKa2N0H
cnF+9aQPOIm9OLClDTKp7u73kxvdzP+Mls9MValXO/0ARy192dv60QbODX5E7JfEFIGTprhhV+/E
5wKLazz1mY3NFGD7hrNr5mhBrFG4eGaM2l7LQxJYYLsTLgTBWnhBHQAeLTupEgh6vFNEDILaFzz2
qdEFlQCxAiSSa6KxRPqddJMC+5V9/exHNrpkM8J0PnoyDiwOxXCEIAjWUTmOXLytPfOWOZL23P8n
hdVbwmvIx9y9iQk9aMJZTj1yE9IRO7lxRYjn+AOlGmpb+rz/p/tY+MwRCymqV3QidOxni3GXyfrb
dx8zR7dE1Z0Heuf5imKUGgfLyix39zBfCSf5g9c96B9thk6e6Tmg2Y7INHCXkJsGzUt7aCrvBMsx
ZwSdFnQBwACRJFuPCM/bRTGTh59E9f8ovC4SrCpgFMUuh2bLNClhciLylnS5m9h5o2GjYXSA+ME6
ELyd5U6iHPMc0Sh2wMkOpagzs+wgrB/0PAH39VhT6OYSo1fu5oFWX0dLOO3bzahquYohrWrJE10h
nwwAW87/+q30Cv/gwNhUmtjQ9IRka3q8WBGwIJibY2BjY9N/NJHYEwpTtYfO8Ii05JdUD+/W4R6o
fAgRFP+bSUy8Q5pykSPzAL5lLE1+eZhw/7Ba1epzid+k3A9lbQAED79S0YnLM3Ob8GBWPdM9FCat
2WuMSAK+5TTy1GklvAUR3FLRVJgtjdgwjrxeCoDdOWTLIdgzyA1pOg/9aL7Y2wZHrmIELClAvY0R
kiXnGkf0CDh8Y9SBSlrzNcqwKr5K/HAptOfNatfLGcK7PEYgt88rTdR1PL2pHgZKDWXzp4yRJo8T
h36PfH2n4/UuN7hgHsnNxfElsa3j81tvq5CqY285a3A2umxNnZ3KplOCy7A07JriKSNVQUMm1ilp
aaSV8pqTlugQYc4xFg/zfjynFP0ibzNbQFBNU6NdC7UXLHzWV/6xdH2FX7PoR1eXF+eQabYyDNvM
EaAMXRuiQsrCQ8Bafg0atlNMwtVhK16ljbzx+GrBNyvoJim0tk9HqPBBhvTc+eK0HAicqzIc+HZe
y8lfTuzXbn6fs5RNFeIoRN7ms+cZljCEJIb2VWgU7qHUYx4cZCaEW55V185llZ7lHcDITGVUT402
7yvorh5AyFpBmQowm6fLwjrd0uSzu2UfEMF9SEDQbgA7iUQWtC/Im3EJyeoiLkeGhGXxbp09LpuL
+wqj5mycXKnpZNw0rIxAIXqSZ+3srLNtLLYG2AYQNHtn/Rai1kxIXd+FqrNrrShVXB+bhzJoXWkD
kBJqN7UAuLfH96K92gs7od+K+3VO1+XuLqy+D/gHIs/kfFhlNv3OdOm8s/1OiCkEQfTwc06IWM88
hDMhhoy+U9vBUFBU3mzJxhCCARbUtHAT8P9AwRhmggqNsO5I+ghrxQaP5mTpWwS9AJpcLlppEE6o
xSMzRXDuvbsjdqCSdpIAF/pD8igXQ3p7Q5pHqJxko9wKJlrDQxd1779Rc4VDfV8qHuk3ccYniYlc
m/+iSvI9Uq4kgXeb6hsKmfl3XC2QlaZK6cLZGTJFVCcbyaKPR1kGAIE55/XdZNkGEs7EqOl0ZZwR
b+UC04ur/7V/UKW0xlZ4ZFJpU2/ACRVL5NsTySiLi9IFzsMUGd81DhAYksFtLKRclzcm31bAYk2u
Evf1MsU1+dBgIMwJHiybjP7/vuJqx8wvq2h6uS5a7bmiiQ+/GYW9SYGou4dN5f6q1YyJRUju9xuu
UmQe/2u0yh35Uwmpwyu1ihHRb0FCGUC6ofaF9Tjs8S0bX0M30whAiWvxVm3eeobZItqNo0phOJ+M
r26jkIWUIirxZFKSO3rN4996f7TntjzvEUdgQMPCyln7lIAews8uZhwsPHScMN8HaVUHu+46Yh9C
EvQRVuKOhfC/Dv1mnlMt6ypY+yF1zCVOXLz/Y5GVXBzDcazCRDlEnYf3Qeu3619wF6hzxw6Tt062
pn0trE480nnlcooPN3EjgNwuzDX4DUjzFo4z04IFgzfglXWr66AHafZdRjJtUNr1LagTVGZ4vJCd
wLAJNiR5xJxAFyZAYJv5Uq2R+Pa8YdNQPhOinVPG8xG4+7LG6jrUQaoCRby4LvcSna3Ihvl0QYUc
knmByqzYg6i62V6fOl2scs5+Sp3Lo1E3QsJyXncTszoDuIlSCDToTxpJ3O/Jxer1ZJuDBOJ5dHFP
0+KNzbi5t3Bjg0sxo3RNcUD0QF6mhvLu3rejHFDyPwyFPT4NYChabq3RV5TaBZD3hz3hqDC8DJh4
P9PQZszPIZhmQ9xR7vckb/ql4b1jf17ebstabnUTsekdkNxXUyY1BzbAJaVX8hOPm3FyoR9KpKtF
OZV6nxaAw8yF/SqI76yqG4JhHuy0XSWYA1u3GBDYbnXSH9Ut9lCZxGEc7YM2lveQ9ZdsXIWNnrDN
yTk690rvPV1UT1s8uUsvfBlWv51Yg3saVY/au9m9ghpBYESFq9C4pRL89q3UXqWR+AZ8/tGUMkoF
IA0UcO7moeA+n9ICfgZSVJ4kSf3pdM7bwRs7ffBTufxWugZR8Q05+vZxL6GYTdN4UlDff9Y8/Hqm
haurWIdQQqa+sPgOBBC7x11l712Xophpa/sCZI422vew31TP+UXqkHj37B4Lm1CxScCLocGWUiIO
XscS+04GX9/gIs8U8w6aeFtfu2hO+uKpqgBJuzJn3QvDEa5Ce6FMemPuqiXp8QiEoOOtyfxBJAnf
jwF71F+Opio4mF4ecYGt0MLQRO331PSO4+xjk2NbbDH6Qt+cCGOr1zd/WYR117PmGDz1/vtVbH9F
Ym8WG0sBdH96hotIOI5wtJVAqL67nUeeOKva61h1tOi0YodWlNJOOauWqsjn9mpDyHFgv2EXKTZc
78RVfdHaP3+t7Ay56Vu1//7cBh/f6g8r0YcWBiL88MZr1d/afvtGaKeBrHieZESq9vo4hOb4DRB6
fCo9hyG2xQGKOYeNGR9vmYSujjRpFOcgwbwg2YTr9WQaFuYEzWTQFwlH0120O1Fr83fCX+G2Y2gp
vD7amc07UXQ6gEdmHSVcMy4LKdxXzt/fYmGh43o/f+IShn6u0aiHC3ZkDKrqty57avr1Zbd3zb1L
DSIuAsQhdwRY1XzdGk0O4irhralaG934ZkNkklZbICWMAWoKdxe7QnUogWJid31A4jULklhrKj8D
ZfYp12U6oc4bXon/r9DEGogFUDTFdEhveBQJZZ6FVhBzpvFBkVDLfUYrTLPh/35BJL+CbUlaC6zl
2+PrXE6zZFr+oxyR9Fesxp98Ne5poARFlQrdEvZX3SlFVnNtYPuX/oPM8elDJK1/h5XA7s7hh6cY
3omSXZ3Alv1r+UPmNkjnyDIjzPTQQ08qw4IlglSXYRxm5712eUJsRwbvJ3QCPHuIJ8mUul3oFEhH
qxX1mY51iq1tKoCVhEwPuVTaOrfwiLGhSJpuDXUUL2Exfc8kxibRvPiWcdZpNv3BTYEu6TZJy8SB
HHLBY1gWOR4YdE4iwy+ge4JCGIlUXkbBQh0oHoP89m5xk9adOdvBHxFl+vexIdN95bktMa+J0+BV
NRnZ0NPksyQwd21+28RVT4ga+FnGztRySYN/qgdXgMoTHuuqUx4HHBY8EmEgLN51SzIkPN8fz64P
UWLy3sikpZ3pNeltbuQVlAYpCChWS7BEl6zHc55ySfZpAPb2zcjYHAn/6HT66UMjgyJpTrUzQvej
x24I9gV5Qx8hE1jrs7dT5VahJPYKlQwqdgc46qVG9UxWCTSGvBQMZR8Jf9wo1nLDB64Rt483havK
Csot+VHqQy2U/UateyTaPDIN9ItBDUKQL7T4Uj/v16AXnl/qQmyirkdSlHeKuF/oNyuZm60K5VBi
fhasIDNW2T+xsYWb4YSFCY51RlS6R8fFSm9aplpMCzxT4+4yNjUsGsG0CekQqY8KRu1QkXnfT5g5
dyqLS+tJ7sZVVT9Lzw8sWXkgRa0M39Recemc0jQIYw8cBc8fQnfboMub64ldbU8r8Un441Y4yq+5
vLSoVLw7t4Z0Wtp6hNGBy/8CKL+Nqf5udL8RseOVG3vfrRN/WOBn5hcFRwJZh2FkZczX+QFjyIwT
E2t+ADHiMKsSXtWuM0SWh/UFkX4Lkl5xl7MJ0OfDdZDgNE/H/ceT7Qq/wkDNsW/1xMJewoDIT0H/
fkrkrN8uba3yiNDDoBmloJK7fMakicWxT8fpPJET8/QRBeZfihUOFGb43ypQyDiQBUvUS3bdNlbX
gWGXtnlzpUIqMWEfmIK32coXRgVddwjvPhrzrgcmgcsvAvXM2Q/iqZgm9LcacvAY/Ww36IGk8UTD
BUAVdhkrx7AKTTUhRoyryZ8GUY9au8XVhGSX2N1LJ7xqqW8c4//89KyPtS4hR7zeG6ob8x7zPOrV
ifWS0vggTzVkeSfZw/fZ0V2X/p9+f7Iw7vk2gZ5XCblU3SpQEQKmReo4jyI3dlaxXvtvo+ldQ1Fd
HjfH8mUwIVPgQ0LrIOMAiLtRxbBNhnA29RQkMU9nBgcm3JxYwrVK0SC88oHkdn7I4yMb3h3b/flg
ioSkOYP3DRQWeEWWHXlGahZaAfVUEDzCNGjT4i7Xg+SV3vgOhXiAKf+qUC7u00Ry8sTmYV9eVK9/
saWZC335auo4okajtFgYSLS43x7vaKJKNoGHfag0VHmqisWzyZrEKnVB9eLfrc1ylEJF9Nz4iz/f
Uuf5EjojpcFWL2MXu4dmAMXJLDfhI3LUbaPHs3/ZGIFKRovnfGUa5jEPj191zwMe2752gqt+PAHV
34qyxBMphm8NLG2iJQP7LcJkh8y4VI1xWTdb2ia05IkhXlu0T2Jd1ZpoaD4iYlEAKnz9woOjJDmw
m345exQ//0BGJOBhJqGN0z63lSeZf4tLlkVPf8EVXRxLgUzhMcewlybZl6IaXA/5iVN6TpX6Drzl
ddiOhUbcM6/f+W1ZT0U+yayaySgPAmIN9QiR2AWHF/6NHIyRmV1VqqRW/Lft2EVEa8LG8AlkYpLR
kiX8HJMo07hJPwzP8Rk/s9mOGb+/8TMksHhdM6oHb2NY2n35kzOHtb81+CND6lDEumJgPqMk7SrD
XJNd6AQYzZXaCUKjYRbQv7i6jhEc5jCbpONH4cavEl0Rnlt3dWyMXyCRxmOAgI3rWbBJsqyQ0O01
fEYr4k+a/4zCWqpOAQqL+BONiGlPM4SBFattWGjdMdNVuhtTeuNWCTYlcVJY86MudSpqdwdD6Mg4
SjMEyuIbHEV5xWkNHg0688JE/vo0oeEf/foCe23BfT1UlZ+YZ3gqJsAaUxJGiB85E5y23fTLt69f
KqV2j9s8lfH73HfVcYUaqwLqlBskjInBN/Hn3cWUELFB8UlnRqEy5GXjEKtzJQiemoRKiyjjFIWz
GoscZccZHFV/wf2FSdbO4L66AxrnCdE0oZU2uxTY+eVhhkLJXjKazN7h2BWY9/8eEbPaAkcvEU/A
ob7j55Ctr6IOZLS805TFVA5oKFTr6Evz6zWtOjfsomB9xUOJ7oif1Vo6jS6fGHvJN/ovOFPsmx2Y
EQmDYZzssjf36k+/BeY/l3ChTDVxDIUzVV3PVdIyZPBB4fLzWyoQgVW/RwYxRg4EMMhF0xvk1+w2
Amwcmszx3JYmB1IJHOwYDK2jMihvHhhnlNC3vAdVL0brpuelOZ6RnKAAA7cdbr9gWMDLtmIhMPJ7
DoCa2q+Fwq4c8rlxeB98pOAbzNO1WXX2/uETTG3Bv4gCM0ic02ESWkBzOctLtj5D1PC0Hn00Ijur
XAayLa1lgdfecmj4w7V+o6dWhN15bXR2gnHxSXy+Qnln68w9HNNzlZxUdJ3eZItMl8QhAR8uk5Eo
zbxc4Za+795AzRJE6INjstQsF35+db+o7lUnuK3K740rXBR7YRyxVSw7xrGKKl89AjardEx9GQe+
VCa36MPdmUd4qzldQ4gnS8D54DAtyGjRNv6bnxTPnAb3B4yhIyy8OTQb0wulgfLsFbVE7oiXEzNV
aBNpppH3aqx6LZwu7W9LyxC39orrioTGRCJAgs0gtLB6tOCzViZOKrxAdKRO28NjDxMJ6sTVmqsB
53uhEKsOzcblvpiGuKF7lwDOSYxfFN9q5yVTfQL6fMunu1v7RAV5MkxGxG1GL5XnNpmg5+tpA0uP
rr2zC406lGuXFpiu80bkv0oIsTP07+/Y0D6NLVVkLvCXXCn/Ou+QoeDDyIsyQWLrHF3A/wnDDbjh
8Ih08Afxkj6gJKTtk4VC5kLowPGMOcFSQj1GmxKouNcFyRxEzLGxInGcnsjjI0fO+FF3NzdGmzLm
YbfsF1557p3giM1eeMe7IvGu+Q5zosOvT95vC108t6sSIiKQtk8rVpFqLoDCunOw2IKsbOtFI9VJ
IEq0Pn99WErJX+VO7rkdVjALZcFRske77jATfbVi+viLzETO6Cah8B9wS04AZOHAdEVdFoI4d2Es
9YdmuiHeR6wq8zXEWU2nu1c9O5FP9ZelO9LseNBCNOcVfKd+boV6JCQSPILUexq7/pGQXDSOP68p
BKBE6TaiejsyZc5T1eUBKFR1o+JJsdcL5hJPZwQSAIW4Muc6QbaBClejPebyzsTS9Ciw4jbBMxXq
Lra3+y3FCTunAJVDBrRmGu8Qv6a56nSUER/wsKT429g4yVQ8sgMkD1Os4NWE2/e4gcHbY4UZitgg
uGcpqUdZB/3dLqG0hRoKmTH6h/Ens3npYdgYMvSSi+YSjifjvUjZZukEc/8xqh730YEtKJElzFHA
Fau5+pm1A0J0s79dheyy9KM+JwoBg4/64rlj5fM3qVT+pyY91NGh4MFPofLt4cOM6Agr+2YX7X3o
hY4fVMBG6qGRE2oRElCLthd2gxcfx9u8KRSPgHBsIBIW0Xr+/yWK+0hV8HWsIJqqbIoLmx3LAIOg
Br7s3Tv1BhOOHFi8iAGeT6N3kCHv02krCzrmxkvVvQjusNiPSV57Lx5yniYu4lIwYu6Jl4M2Oepe
v2bsefXbxJ2u3MQBBaHM0P/zZ/iglZuM2dVnGOTYbvaBpfxLvviDNB/41MOmUG1BcezAQohGHorV
MS6kjKW2FAgJsdDKoW8YKP5+AeFWj66PTVyxZRv9HtBZ9LaO2G+VsojN+1LqLfsPSrKCDJUSo/8S
rGOj159KP2IH8Of/1ijIZilotazxl4fb3yzJUvfxWO79sPN3gmA4hxO8fz/DuexHam/jE5Y4ZjdW
f/iN9xFz1ME+Zo3SoKxn5BFUhEWA40W4G7UCfPe3V1r73hPdxS6BI3V06SsM4rp8V4DnAGA9aJOh
DU6ZUDoOghn2oysyj+5HD320QZNu4S4lbBTgIU/DEmWgV0lDS+g82KQSeBhXFtjK6n4UGxWXw9JV
7OVD6TqlB9i+QXFjP1aHz1+AGS6PCPsC7TPMZg8L2typMUCPjhpDDH2uNq5hyQD7TCkonCxvzrSX
in2+8uqxNqElTVEFU+pNd8zvUMpBmnfswV0D0mF8K+zQOFwC/hdVYTiN1LYXDP6Q88YL0btlK+DI
oJu4AdhAoAqQaSeQUrhraBRjqXy9SjIZwDwhZPLUYJrupusf44wgBWgIdzjjIGhKIGjIE0oIOiqe
7mcIO+WaI3rylyPnYjO5EFmgzICtOIttqnH9jVjijiJ7tiWI1YumOIzMaPUiJMi58LcYJV1UotYG
kllDuvHtjxR53y5uR6m5NlOkiNfajihqoRJDmuajzmYbq24SJLUAyTOpWBAfUx9kE668B5MltFfG
qb+WVOsX/U/1ha18YxSRk0V4kURkC17KNrBQsxZrDNTKoTm53Kfng5MRGjcX9B2KHNo4MvE2weQC
4B0bvjI8VysyLN1HQoh06gcr5oTl45R7DHh+ZAfjCgs3+EYI3K5V+UOaAUMy0SFLOKn7J80ndHBv
M51PlqB/kJRwT+QhJphCcLKhr3M+FCmHv7kyisxyiVqH5KvaV2H87ypAXsEvm+Jlb1nTpumdxjvB
yS/E2/6qdvZAMjSpeqXlAbA78IAqJPQ5efIwEbcInmJ072JxmjEU6StKONwcOZcmRlWKnjXQ/zSU
XvfmDamUgkZOaKMmbrL3xNOoiGMereo5uAxy70Hojvn1zkb059+xQtk3Kw5YgXg5ZYq5f/jYC+lT
aL+l7OZY1WjyN216WWu9XHXikVDF6buIfJAPnA9ybvusIClywbDr6sBuk0KyMol4clBpbGSGltiY
CIEkikpbtJ3CtDQLm8KuJj2CiT94vVVEYoOSyKegm18SVamm3zicsRfTS+huTktVh2qTZAuWXxXd
Duqu7qojXO32bpvb5Kmin69IK+qgFJGAY76Ei6tG3Y/KY145d6JdrHtAbikZLTsX2zbc64BzYOrZ
trQgdocEIZpJQ1KM0VXTkZAwCvIGUsY/f1WYIdTOA0fSoRJ6uHp5Wte8RWXtXrJ3xr2hQQANMJx9
1NmL+K5oKdM8NG+54KO27N4NnaHnwc4HizlSMHvEJUHeQjypuOokTNIEFo/gB/dKgpb8IWnBGa63
jgKqqPM4Mm/TcyYyxwEjq2KKzv/7qBGh0KsjhSQbiXm/8HaTl7H6l/OQos95d9u1tUV++oElYgmN
0pOffkQrP/V8xzo6r8jldKFIZB006yp8YxGdZHrLJWLVJNjaOZzSXChkhVLwVlHl/yUZION1bKAH
y5n2it+yiPT38fPuP9Buyjh3eGwPUpSQ0DT2eJMcW22KYrgVdkFKCXpTCsawmQ9ifaY5pUKySs8G
6XNjY6Wvqkn4+sqguDUJ80ICpI/yIqmCW/htQBqUAAyYf9MYkp0ab/9sGtrWOLUsSZwHiZ69vmSd
JPA3UQhaJsaNrfw3h7FN+9lSP+xDDEJsIIQqO2dv+ep88Bqh4EkR/01OG7XVHETtCAGyS4P8sYLl
33A2Xy1E4QnRv5cmVFg9s5oxrNPct/N68mf0+S1m2zG/e6BUUtJ4DikATZYI/KuHvoMXrNYuiyWB
WDa2ysuosKQHpg50GeRq3BZNRla5cqVStPDrXu+xXEnA0Q/G0T+nyfIIJ166r4bxA94rNwCCtv7/
7fjavRV9scXOPzm2bQ3C0DpvAfoEOxw2ENwJ3VElVGezb1qzWJfifKyppaOuswP6X+Qj8OZ4nYZK
yqdblfP4bsm8NEcCE0UO84SVlyoi6BuM4g0h3fx1VdDHiWIhCHpKhskzZlylmoy9Ag+RZ+zFFCXO
gXl+UcIeJYlmtDWUxVxvCsDcq4+0hviRjohc5/iSMeVReKZ6rEBezjslCHD68nSm5+KZi/AkRIyM
heda8wstEGhveiE8FclC9Qd/ysxLZWWyLAmbWHyiw+A1+U8cZU7vq041KqtksVuXpG4GJfrrkzSD
TDRO2OpCUHiYbBlyXVc7bxFhAi0VkuPluPGkuBSyoC8zWLmNwjfVePdvkeqJjEY3vc7ad1q+Fwlc
ZM7Vei97+FXTOlCCWU3HvJqr7/7Q2ha9VSC95jeYP2WRqH8QF18Gtd+cbvoZB5cB9WWHSx+OvwGH
wzkZxTxHtpCOhlr7C070+sQA+JgJDTisdVt3S+zbOAPGBAAYN/g7tEeWFxZ0Hh/ZJXl2V1cuQw+T
4PXDk8EpMVwv3ReZ/LKIhyVOWRUfyjZR2pDqv18Y6FdU3d3fQzueCW62DLPuWfDFSz5nC6AJkuWn
10uEUawSEFDp01vvUj7zH/HbgzYxdxJ2ylOv52kA6gAfMaCZePihXfe0dWO7ZDXhpZy9nuu/fEAp
3RaAiIinIbqHoXwHkGUW+hioVu6dXD72srX0svvQSLl/QeMkRgCJIQAqR0EFSr08hFyqcqqiwy1r
kdCMixUZpcjEr6Dp57d3As9WIcXUrBpqZaph7STpC+gIM5mdHv9jA0ex04/OGobHxDrVIc7mmlVb
BvTa0yyumfZI8EbQl+XDNxKHatk7DDNDgVSx+eQXTHVfTlaaciZwrfaNP3z0+o2t1BoBJBwoPU4i
7Uv9f6sMTkFsiw6/9JOnODgChr8XRCJP8obZxX9oeYcKTjbQSpTqiDrAOyUTY+AB+xsloqXT/qHA
WFfuiWd0DCZp95xBiS66f0iTpKRS/8unXsS2tUS2EB17fLcTSpr+46OnnU1NuuXD+DIea8ryBxBe
eFRCC+WBd7hbrWIWKnRQjyQVVhQzFjjGjWz/qut41WWh8MjFVlSBbtKoKOTo39W4FPlerh1r7r4f
pM/cblPkWDvlem8ZnkBYE/l0gOBa3WqzP0wY7SwBHtEovxhE+VlUjh5X1kq12YF+BPUjIVzOZPko
yCvRhqvyHWrL51HToKmpFAKl6i5FXWwNmPBIB5QDHA8GNiD3d1UWu4z1jlsS4df8zS0iPoBHICQR
eCeDQz6cHJIxOVZS2jeux84i94DsqKMvR9f4rnO1hT0P8r9ZwitOxM9NIkALh3zw8/YzAL1TPo+D
qRnQwxjLenRBsD1i7FSkPP4oJFOipbsf7BnkpQ7OPNNQJQTBEV9Ph+YTs2p0EoF4rNzIkBPAQ8yO
gBPE9nwrQWebHXufr1h0rzJGmT6G3Z5p+xTyLaF6Psq9pH/ACUPSQErURd8vwfU4e/21ydg9Ac87
zRADSqYVxFEWxSuj2fpYaazRLdvfuPnX0Rjj+nVuWnppUeZ2iwlgNJHWhKfJfG+y5z+MFYQkVrXX
tlSN3/iT70qNlrLtK3uJnqrYbpht1Ts3hg/UCk0TqtSF/FzPAjjbAqWDlekFktMTcupbrYJvBxjn
3Y+jG/NV5YFiZTlMC/FEnwXsmNiq8RNMZdo3LSRk7TOs94cA/Cp1UfnGFBxcKB4Q26+rIu/3q0+C
qKWPEwNY0fxYNvrRsxuBf2/RUmh9s6hfrQAnRhaUhzEIAG7ihPscCJPfA1Ij9pT8wfCGWLnxLvTD
bSQXNvGNpwfz4MT2EGZsvnbS6dIm0OFaIUGPHLjbPZjPpZ/WyFy4m04dbfDfi5xUZ4Y5FnsiGgTv
imPeABPn/lGNUaHXNqxJ4Z7otpcnflae3/78JDdMn8jF+VnwaBmGylkMeu3QfUt75CXL5kOVzH1Q
dJSJ/AcxhAme/Cv0157XDN2n25PjimxDsVsryLpuijQY/F6Elyn/inJP5NG2UsvPFu0hHVqy1APG
ySgNpkH+Rxi8iz4JO/EVOQ3e2m4djLDDzGXWV+VsDur+FGk2w1qKvAIwDzY5hlHH/nyk+Ff4NNqn
y2Zd2ILsxucQVPl8AUFnq/Ku0CXR7Wk9qvz8bqE6lPETHkPZwow6loNvgg3utDjteJ1TFiFv/cB5
Tfx9wEHzfqJ2o3yoIm6Aeu9eC2XUc6GzIuHb1F7KPC48fGd1VVzvtJlycjNgxhNjOEkdbWmRKjiC
AMUcUfxTZSdRurrB0cB9/PPnFkXCNAqiAh/lIwRwpdzXqPQ/17C42WPg1WD5s7/OYxVyOq47/jBl
4bqsenrbZIWkVfAS2bmi3tZD1ZSYtzqBL51c+we5D2JhwLew7uOL7OHSoutua9gm16piDuxUXDKj
GhGw/eXDnmeEP3+oveNmbDpK6IlfaPYEn5z81wqkSBwzE8fXG9WdKmWdbUOpi9Uw6kmrztX13iFH
eYSoe9tDUcUlf+iap6rf10oXFD7StOMvNbm3m8jlR8l3fakN/N+jrO9mQowsena/h/cOeVx+xszt
FZqYR/hA7D7kYPTZoyTmHFpKZgDb8BcClFvbE8x/dKOd4iNDlhI+GGnUpogH6QMfDg2I56Qx4cSD
hDeGRKqMtlvj3Jk4dr4Z0oJLfeBKlwXBEWlaP+QA0QgGLiDFeXH4ShecqnUkZ/nsKHKiAubWclqM
02urVTTQuBf5ePgzrdY7XEC6g2Ymb0iq146JDhJaWClNBYrYdb2KqTthhDo0r1aWZhcfd6Ac4PHT
uoald+l1QPdnHT3hdyuzV5LW9CXRucs44LL5uftGi2dAnvemv2bjkfCXwKspz/H8hTcAgQ5Cr5m3
kbY0u4FKRsXt5oFGnyTIucs5hCIUyY+dDhwcPufRz6ytlZF/azmedUCxx9jfywVyMLqCjDSy5l3r
r7Vf+IbVhf+V+wMnwkTYDjXCOSYK49JectmLfzWkabOclAS3MA/mAWmbzeAj8lyZI/nV/woyLDSg
Pktr6kvQ0a2IMhoQHUAdPK+H2mtBErc8pKISGl8LNnJ32espPgGiFuvtB8x92tMNmkwOpy2yAU+o
T9gxhV4G4LP5ifu5nwhGZvbzblYdwlYpydswTCxkkDFd6IJN9BFw+BWYMEWZixRQDqUFxyXu9h54
PutimOZ8HM2BjZzqKgMZgynLcrCR67zh1HGNNCFCCEhrbYz5oof9tl11VVXgptlA8mg7MYO9rJmw
F6tmSWBh5+NQiAGi9z9QtLGaizpG/CgdFceZhHE/eq+Wi/hijEKnvRgUIwQU69YsIcgA6HTkg/Ey
YJzDtW6TmZ9wxlZ6GZUo6MrLpG5lozsW+KWNQd/eIyPaTOsqy/sfxToV1ltg8KSswCaWj1BrQAIj
n7oPindsNsQ1Vo2cp+2g9j4QYPxXp2fTwJvsUkcNVZ5SrcV8KHvxIYKhMB5CSaZoQYhLWIkHMaya
yXntzzlDgXPz7vLCPOj8U8mEBjivDiU7L7Hwm1PBKHIY/pGrvCU0bj3oJsqnadiUn8WdHNWMd5Wb
vrsggTcvdMFarTJP+Ox6xpeasKVnzM9bpXe6xSXgyd5ZG9qcGSUpygYO0Ovp6ByYveUd3Os4ojpT
03xM5vu/fJgaJYejl1ItMo2ObvY24kd2O65l4cyKOPSXaB8vipBtu+UzUUUbqICZlr7uzBCjJjKC
rAjs+wr9LeZyCsoLudmHcahu7++MVPjh/r/9gd8yMd1YMlgh+dBeUU0uBnVHKvf9izFj7RJUc7Lk
AxOQEaa3Y6EBcvuDe6K7/tqwm0C1UwPoRMTO4C2r2/OYj5C1oTi+JYkxPmJV+Rfh/GXxEwwaAF4i
ImxQzt92mfxSaJC3U/AI6YO4r7kDTBf0B03RWu3u/ARJOLLQbrG3ovApI/8LbgYlShaAZr1RBHgg
xGhsGb7iQswngJeWaWenPLwjG5YD7zbUoWphn5i78ZbM4o3PdLRQOBpbOzseg4FHDSaU4iswTlJd
oehj1OInI0Wki7GoM9UJ+SgBrdKvEl+MMZKzOHCqMQv/PbRUIF1KqD3TnM7LlUjnJ4djJ47KDJNq
GIyXRV21Xl+TOthO8JdcRo5uzRf7Rpz5GP56sKm1lLEDLADChNSWWQdG3CHTMQuF14W5+HAXer1d
+0pyakpnD6e8HlZrDv66Lg5IKiOMJH2HofxKbu4ixVc0yDKDFVcN4lw0tO+JehKhwUCWyPX6X1Jc
CNYV3rU0yj1wj6yx5PsQm40q8l0mAV27ymMU3Po/WdMhqRKtlKLrGDMjmaONlmQ5qbJR/hm4WLI8
Ok96kEUsRBNX+HswH0hAAJmI0llX1FYVEdDPEbUgdIu4jSJZJAU78JBhPsw7ypT5P4CsFngxq60m
m8plksZ6DegyeD6gg8vVCHHzTlBpa0tTOYCxeKzpZOx3+zVSYtr0hAb9UXfnO+mwUXUbCyzVjtbq
WYo4qaLYi8D/fofEYbr2bhjW+tP2Pb59dajMjkZVZVKON5lZNTsEDAg/NAvF6eZ7duQAqOzo7jeX
zZuiONZ5fCcAsB0ovZj6bsiPr0phkPeWjhDnQMCruke13qR4x/KnMcFm13dj9EqBGwLxMc8lxpys
VFerz0JT84Jzg2UroAErpspkB4Rh0G9F8AWxhUkGAkqxVfceprl5DaRjqaqfS3IOMlH/fxsoaTb8
CkVnaJKEAFgilW0It7AyymHLxIcUwV4crKdke5LMG/ETF4dmzo1LokOS81pZvnSK7iCDVPgQUmVl
SUquc09Fx/8TDnTisUF45CC2VU0YmDKJ8U+NxXzkwy8MdLY+jl0gknpHiKBPkKXIBmUwG57462tH
T4IW9FI4XDUmaiBfVRaiilGN7d2pu8hZ91TwyIwn2r6i3+v4t0UkyK7CeKpwXJOrqmXrNuwfI2xJ
jJA3lvhHq4fqQIfCuTe7BHrca+1NV2Xg5U3WgAJFqPTRmdkLDnmYZznaDqH/9zBh0V5rSnidHoYx
9GDl+1gzrH8r0Q2KbgCKgDCgcZ/iM4FX69FEKtjMahX4GMbqNoRCM1ElW9oqn7zG8zbk4PJ1u3sO
IastZObmq/VkaeXhEHjzAPNpLzG9YEmOMBpW0w9WXOSIWShXe66hy18imfIKEEXVMOR4Y7feTzWd
yk1g2d4bZqTpldNdgVX4hWNu45uwXKYNi4qOLqRnTuLnOza56RNsxX7w3GGGqvTbQI+tWZcrca5N
/fexI3DzuIPp704Ykj5TJzbTlTY4pjU7plhSbQnYW+/jVMxucvX3I+UYs8o3OioJ0Tu2SX3+1Yv1
TWP0jDbfR6VVKlIe1ulqbM9mvfuMrgQMysGeyWaRd/RmS+mRL2MQAEJdP0EDgsW6uorZjXsmsyts
P10u7hD9GpCD7UIHSlKXgDUm/uVXTMKU51KCCDqo5nw7o9l8DWPCW1u4HvDapUbY29LpoAQPNrc0
sant5+iH+5v8jOmVTd1U8U4JpHF0NbRqC3QkzdKp6oVGVFm6OrG5lpeMIJhKyFl0Njit/9fAXJs6
07eYfI51h771wHg5iHMSYtvOoC35pSVeHXhDlGlXoYYVgSqIcNlKahDAolihmffnDyG/eM5bdbet
/xRgs9kliN1OfKD5wVzzXRagcshPUwA/q2kjlWp3aV9tM31iWP6KT9xRGhiYVbe9kt30T4Yqpa7j
Ff6o6NPQu2rtl/VnEcCAeS/vfWvvUb5gGZPZYpmcFLZSmpOf2HgB7bLwGDGyicrgZ6wPLb01OTFO
UxBKXr38gveu/PaD4S7BYAkiBBv929zXp2aJR0kUe6b+WoO57x86oVf1lziW5upRUVvfmEbsi406
/OTGDpnCjcqqQLY3EpraTj3ewhbZ7iT404LyEp4OBcdgn3tlaE8wcQtgml0bMCoO8zyy33cMJ9KH
u9arPh8EarlVo+qD/3XIiOhLTN0r2otXdKFSrztzxrAjR2efR/jZWcQ9hoRd4Yn9cnpTeWMCA6Fv
HIdJ1TP3P8pY/+Uu+cGbmNE+PSjIzaU7ThzpJ2ysYm4T17GBm5cpi1EpEf+QAKhuQkLK3uKUSOBi
QhVNGkylgxdxrzMdppv5O7rUWrCEHFyaxvwurMeNOvD2Bfm/jTmmR4c+HcMlNuRzdk9fpvcn5Drq
7NQ33wxf7bQn8zA/XPSkrYKQTyeEaclZpqc9sOxQnoWJOw0MmmM5MCD2NEItx409EJgN7eUYnLzK
t3X3CT/5r0aRfWmZG7OMTacqiFkAoyXuG5Gimkr0hg6u9SyMbk5gWHdXDvGQNUwYDbcA5/PSJieV
G9Dw86ODaQBsAwL4ctTdTBxKe8RXmkRmAa8WA+PFpuRAtkBkz2ShUWPag2K0LldeSl4mNdfWe0kt
Gz5C9kp4WbP/dlkXMypj9KYpDvPGBG88QF6D4XOODRFmt8xivMu4NOaqg8VAndrxX33A2pKlAJn4
Oc3RNp0GS9DI10JomCBaKD7E78a7V2vAjH9Lg5kNy5c2ReBIUjp6yC6SoToS3yV0TfNXnkBVdxJI
DydaCjn+Wqew3iK8Q23Pjgjs5TbDf80HQ9dCh97Xg5Jff8bZyci9o/QymbOy46V9hw0v2RAw+b0I
pjCbU3llZHzMxI9rCkpZvoDQPYpY41ktl1520cKY8ffOcqr9iYSVH7iLkH2w0QPqcCLFfhpiDoq2
hM3fFXPpFNBMkTjYGbcIqCufaBCGoh5qlo9y6+b9G2MKD0mcYNr1HRzBVEs+VniJv2GZMC/stY3k
KbRq30IWHGmr+mXD/3Ssg6MeMruT2V1SD7LHiSZQ9Nph2RMQ/Z9pLY+NlgCJP5RkmJPQlwv9Mgp8
OXM+msBpsyZOegstkebovkkhaLpxHiN+LtFysCRaThpdb7CmHSoT/wRRYWvMkhcUNpK6P93cgrQi
bHAiUpyUGi262KpTeV/qZqOaqYj/HEIzdUJPz+C5wa+1Ljbu377KEaTXbOcdaag/1PgJSWn4r17C
EY7fs+U8L2bwhd32AAnq3KLJfHMniUJjh/l6oGK+PRMKQvrh4YKZZyL001vTN8ALuyTuOFF5LIKl
PY/GE8djI3dKIny6oOvt/Jzq9cJsZYv5QprvsiRrkntqxaZXoy/aBbxZr/450ejf0vdaIYj07Q6s
biJVq0GkajuNeeCM/JfSm6tYUmLzKPYerkPAjGYb1+j5ueY/kZaT8ypMa9lFIsxcqe5rk3cUQXbB
imiDqMeIXDlJOkPcoZSvR+lxt2n7RDeJuINz3J6VV13fkdhNR/lPSoRcl4+pAGXzJvJs8fGo73RU
x/TeTN5TK8OgOt9S83zUh3AhBop8eZlvvnNi0c1JtX6Ne1pxAuHF1b86wnjSIE//KzoQosHkDcWi
EF5yUtN6rS4vuB6ePpmNsBQcfUmQ7nqKLeUByW01YtLMDFEd0+m10U1pOHrdaKHAb90ssQYgYxFU
iSGDNj4vkTpW/zfYfQ8tBhKen22rSCBsqespp06NvFNlIOyFGiaZARXy6Yax36ETAzwT6K6nWFVA
YXNWxPuWHuh1woXwYedbx0bde4VhaKTzlZEqgtDScTSO+374fd1/rZGYh3gr6AJ6XlZK+8G4A0BR
wEKPH1+WoPMUZQHh8+8oN44pxUktcoJyav54GOGqfFrC2a4JShx5sESB1EsgtRQh8VVoJGbNMglk
DuRQEqXsvkdnamnbrL7HPLurhTZE/4XrB5Fbi7CPxaAMMWmWquseahe6fVWg1ub+C/HpBrguJSGP
KuslclCixNx8Cal4ifHuw3BhbyZFRCKjJEP51zPippo3t+KhhVATwe8SjLjj3JliI0R7k3QG5xEo
Z1goNnzfYzktApLKcq4WG90UBdj0+WdXAVh++mHkXLE1/wqoDuJgAKOmnrN/gbPJ0N/EZf0x0JV7
cbE/MCP6g5qyXHj+DTOcu+cxqgGxTYIrkcYkw0/HAA2tVfSsIP2blSmY/j4T2IiSjkaZ3n3mLQs1
j3PR3jiPU1MseDPv7MmLJFGO5A6hEIrae9c1+N8Vwv7AYYwCfr0wOlKBizIpAywTUdnjLZVMOH8T
gfw9fau9MBh1MFGorr4Vqw2e0FVWyJRqkbm4sO8AnBuDKbs3yEbxocEjtmIOF2+pEyv1vyBfr+Jw
RZ2AwrpljhDs4TBWz9JauLuqI0R9WsULQzaMCXUzNKGXlt0pxmIbvZtVSiaKhsRinaxGHYMi2HF6
nNHinXbDac6Yp/bfQ2mnZaIGejdhPlekQMOStElXpREk+P3xWnTWMF6x7upzBICYEQ1a7BoPUaOj
qLmkE0HrS4ZFZwTKOD8Lbp1IpWsz7y9QXlQkxkzs+mrThzTP2Ox8mJGRFl51E3L/YdhUk5DeEmIe
vceRm4GF9YU0/1bsIb8QXxnJs6eBExFpPtCKE0anxZWXob7mSencs6W0BCf6mE897VnYNSe/qkp6
1UQIS8FRzVhQA46o2mae9DXenssXaYEA57F6AWVDRf9RAaMeFIId47ozUli6nyeAYtFglHmG25wA
IqlsgBDBomMc9j2jKGY4XBYpzjguPoZZRT/wyZTHONYxrCrywZK4jyULZ9hEYvylTEgulOcgUyDf
I0CaY3kuZg9Vu7FXOSXr+abZEyWtRIlhEQE+VTew8dqIjvDTsSm7KYLH+RJKKBC2pHQ7DHF5fX2c
SagFmRkeuQzmQo/44zK9hiEfrsFCq2q88o3wDCFw+IL+9RKmyJ3Wdt+sqg/Y9D1Xy9AZW4sNxUZK
Wlhjmn0hYjWAOR58zYFoHYN9Tcsy5fWaEs68ANAM5TYU16GJdG6sAq7AszZMuRPSBCE94kqWfVok
q5wKzjcTrG7pwFD0MlMir8qih4wmu6lHma9fECKfpzo2hJ9EzMBGiaObNniVu6YrmCBT1NA7O1bj
RvxOG2RYPCmSesGmEFfkEfE6jrpxgQI7xVfzPdLHTpG+pts+7r9GrORNQ8YF0hSQxCpKXKIx4OZC
Pg9UAGRrKMTMdLiiAqlj/+1furL4+vdukKqPsgSE3up6zJSawHu3ZYD2uY4p5e0jyVlyUlMJTjP+
8BYb2qs98U7fadh5KtcFC/YohtMPmAiXlkY0G4jWSM2E14xfQxff/Ln1IPQysBmNBSvqdfc6JGS9
6a23LC2pJOR10bV/PqfJIHU7gbfB1r2iy/q5el0gPHBEIHF9rTfz1vp80yGoRWFBQ6VfOIBGDclP
W3ij9p8isPlkRkT3lkezlq6ddoNyu2+X9nAsuy4eWWGeyuGYBFJV1tsb3G/51SNFB9IGCH8s7l2b
GP3Habnp1ByWkavtgB9KProgVIQhayhJK1i65T3qJCT7QAb24Ntq7gnaOveLggalJDmf8VtmcOMp
Jvpi6dr4fmAErewqdg3jg5EfJv7HcSmf568OoWXlaCFL84F6YfMy/4imZg8i1Kr5OXwGVkT+177C
dHwgBO20k3B/hyP577XQCb0iwtFsfrXWq86+90PtPwxsHZNXKRQk2NbzNne8WwZq77trlC2GJFsc
t2PCkic5/yk6IQzwCgBhEAA4K4JwQMSr/fSyoj+TBUf5oGieF/EwxjFEjyRjT3jkez+qLSqGJjp5
GweUDywxdDrqaK6xgjbA2WRZ4023mtqSEsghnQLSzXmprR2qLT+DehBjRR5gX9N0VrnDY2AVoFcE
rvslix1RQSYrkZijFLKWTyoBgA17xSTDGYDW+OIB2PqPBM57HpdsjuSRETTq9f7ZVYkMEtZWUIRQ
lbj2iUdDCKWiKgDeQz3BOqzqxZMijLf5P+u0VkGZ1zgFASDgGD/BSWeT4bvcoaIBNV+vJsYs6V8j
ME2TjWXmU8u1NxEHx5FHb6WvSIp4gXvyVPTZzUYkMtABGQ1q+Eubt+f7pBAr5knsYdHsBmfaUnUW
NJz+3HXjMLM7HNEwTD6yoioWDVzQXZCQUDiTOmsU5LKTkCvla3+LylSkcDXgqdt/gGH9zs5ozrc7
hlrE0F4bTUbyJ9UzGot6g7E8EDQqvykrL62mft61QTBSRMayzeG7T90UkdCA2T6wTYWk4DawmVdS
RGKF0sv03jIVT9UY3B1seuoG4LWvWRMGtbrmNPkI/pjVaYP6t/gJnz7h38aemY1MpnCpmWAFELy2
srE3zGU8VnRlf2+lGhUED4HuLw/wQJUzd5+KiWzWq3CrVFGMJ8Wn7mhO69xjD+yHAEtLsTABMUaO
4MxLgs4U0p8EtIBISdx2FPfyZN/tQmn+dRql3teeE317RPmKBV5QRwLRfiRl+SkYxN0Aur770ezq
wFIM7V6Y/hUJTCZB3Ocgs7zwwxXoP/fpuVG4GbSelbls3crRNR54xmK2RYP0Rw73QX5fh7djZY/h
WcGtaGJOp0+l7Hr1bk6RY5k4pj3dPtnGHmknORjbS6e0fj6M1hNdeCIomS4QtDgLbGzkWLO37im0
7jiVMYQ1iJl8a+cf7C+Ka+DrH1YEsuBm/BGold+vOjWOMd1XcL93Bzigk96vsgoFxXecxupBSk/M
nolbOI7d+KL9NXPQN456ODj0SiCMg6SS/9p2gLSdePQSYCD6JVz9BgdGbjAIP+PEj4v+KFXbFlXX
37Jof4CF07HGcvWqxq6XIkd/0O6HkgUD1ee4tfBUfpSNzhm/uqe8BUG61Y7WWNEAxLtPYP1IDdmG
m5a6N8TBo17u57V+VgdersG3I9kVtoDqogu1CqXiE0TSej0Eaa/OjaQ/w+Xjeqcn8yZnyoyXepHO
5DgnZ4yEDlXeNmKKw9toPc6AqZJC8X+Q28OJ91iIGF2UEnUB7kHuM+w90zpnGIDR199n6Dj8ckBN
6Ww4RpTwiHVuYA5iCPngGdNQAlIWipy0+wqs5HrX966B2zPXLdKGmrCz2nExGDq/fTRHpL/zrUWd
digAGXO+ipkOj1co35XomWO8vRush+zazbvRWzrUEzUwSM2r+uiz3mdP3RsFRe0tFWEmM6nCueBV
OuNfqs+RfbdKa0DYYSBejz4XdM9JTCG8ooKGWWRyzzqy5CXuYSOIDbdAJTuEl/+haceb0UezaD77
/g/qfzz0b5OZ/61w1jMQz6jD4f7Q8rCsMFAAIzh3rJ/b/odhwCy/GgFKfibs0yh4QVlTm74/UR1S
cBSWMp4unBZp16oCye6TZ/hg2swa9hTeYR8XwthSh1nOMVpJDe4E/yXzOHzFzNkzxxCWGQrcoh2t
f0TQUSAQoSkL82fSwRRAFLfDO+Pl+aq2qKkWt8C2qKTpH5FuG2sdwu58+RpzIs16tbKi/LhXaUOB
wJRh2Js6GD3bZSD+EfnH10anry/2jeTeriuOGt6KZ5dOq+/OXRkYCIFtOtd/RPaYch7bixBmWvHL
tIHsLRaIVRZ2i4ipBCRv1qptd7D4G7HqCKKRyjlki64eTh4ZQIMPMDK+IIDaK6/L3CY7X3SE0jgr
KLvTeNAdYbAT1kY6sB8wMQPCRp4y/JQK9KzGilpWAw/pP6c8TxsD4q/c0y6qdrRsBv0Fp6cpm+5o
wBzKiwY48KBzVy6d4p9bfPVxZdPH9qM6hsgorBbyfr9ds1TFUH+h1SG4ugtqMYouGpOLF0K0TF8D
wEd2/K8axQh+16PDBjwqn//LL1RCcPeDiM8dBg6dfYxIAgY35Gz4swcKtVTZoeeK9III53NWGzXD
/F9yRdyHoEuOVLvkTJGHMDdIJN3wctQcEIVOsC3cUnBWheNk187jh16r5wOKzA7s6UBDSljN6FPR
HLYAV+xsgIj6h82SJ8lhGnakRxyqJ/4xG/YsKsTtUxqxUJ04dgrbHzTVvSzWBVDm9xe3KnZBkSn0
KUNeuQtgGhG6rNwcGfMkWtBdQjepJRBmiAQJ/YjVvisHcES8Hol7XT7yqDseMsUkM7UrlageDQgP
Xh+fASv7pF5tTLiddrPMejaGcdJo5TpPor2xXAvX6F8adcK4v1EuWOnBJ0V6YjZGU2t2qxzs7fs9
os2x3N3DpHNytFwGdg415b/lOmlbtEKj5oYbstnm5teABB6OWXlugm16CpGbcvS/BYkTjhF/z3OF
EPm69iNLeC3hg9eB1m2EHZ1wUbN6wtUhj2eGE5YkBUQMlPgVRvd4jzke8cjhl2vc1A4iuDk6xPis
BNLYoZ0zkFaF3SLtoOglcwFQfPophFqSF7Bpj6C45scAmSckmYccrfqA/Okl3kaZHYOLn6S4tty7
iB2vR3mT7j+KE2zbOFw4GICrg2q2l/a8T8wyGPig2vhTwWIqHCja10b3xaObjENKOFrPhawWtqjq
UEaHgzp6uNOnce0Vmk8cVQwHMsyvT8eQbd49wRT1waZykIAlVus3oih/vsLpODA8hCNyNmm6kzae
3z1N3GhZ+3O6sfsU+MnMqL1qxYQowUFOGWjTRx10l1W5ggriP+v8kIP3IWrroaJPFMcbtuUwyXJr
1wUbnoLvkcA1jSk/cdh1jvIHzDhUFvOMfjqhg296lF6MTnpbzOxW8prPG4huTrToyrP+UEJR6c2P
z6vh4WN3tqHOu7Zr4MXDF0Nom1PtRfpAljVNgGqCIaLitwg2RmZ8B/vQcuOn9PiiBMCM2RtiBaAw
PI5vPN+Mz1EEb5LMwKdtFRn0rJRtVEXCSehphExOGyEwHslJACeSGenkxP+41QfGHjYSqOqic6bL
nvLKOMPuypSYKNzOWN78Cyf6nUt9duW7mF9bBNihoZt8NBCtLJ3Tg/5p60/tYg+DVcFQFqhEzkmL
SYHiQfhMR3Rbm5jOeIXUk0/b9hUvRf64T2c5LiD8Jhs2tdckYkQqxcExDW8azXLrU3p1jHjnMy5J
H26lujijSmGtKYUF3R8GE/urNEK6/flkxTfDkf5Lxim4In5jC90W/PFZ2cmu2FEX2UwpeSDjmMo5
+AmdIjhFRyrPBTlaORNAAebuJ3mvgZkUMXYYql087jbf366sUuV7xxU8nc8dyKvBq1kWHAGspVKj
xn7elk7XOa9JNulcf8UkI7KIkcav93Nj8x3nbZwDfN7SE+GGKEhYDOlAwqs2tjBEIolKUkUoSaNT
yBq2QYD+WTHTY1bmbtI5Z/36SwflMFnwOq1VOEHuuTLq0EZb4FzqoJOR5ENBz96kY3IJqaZMQOP0
pKhedUBbWUTGdw0bOPph1waXWmsmEJ5fj00DSxsEec8uJ2HmcrPfze/B1uGIbFJp0KWFEkB34rMA
xu+adDU6HwqhahgkREPgc37DDhn+zw3hx77TsK5attGY2nvs3TrZssj3tjg0HC8GWdlzBFVC1OoJ
x2hqc+adX6QDj3+IoqbdBIrwLEqEvFt7FDe4cZr+JwSjL8nBXSmTrS5ah+pSMSnM4mMN6ZfCjDfX
vwiB1yeHwIbUtJb8m4cZD+6SUX7PjtWUkvpjXyGwaST7q++IW+RRsUSom8Y0pV+j0SlHPbVyi1K2
NZNJzqQzwAY0dn11LpiqLguJ2gqkQcqEnkcgZwv3yExylGmcteSlyYN3tSys0pOgkOEZ/Zbb0rLc
5V7GhPRP+zZ4elFDRd2OnY12aMWHUMviKk6cgO9YTMDKV/Pa9z01rqZjaA77octWSHnQ00yLIqRg
rBH08RYem2DwRcUysYgJ5dyZnz6tyERYkMMfLddsAsB4INC3Zc+6l76+niCkjvbiRpaCrRYZTK4f
ASNxgm/jC/wQnp4/MJsIwuCl7uWl69lu4BPATpgWIsr78UlUInWYALbVqv7Sk7DP9h0DpKscvEsp
RDGWrQ5HAgEgLDz3M2lWmKxNlgYiUdnKsXSx5mcgiw36G+juVQOok5JDmEzxwlVc+3RS5jSLUpWZ
Eh5ikDMGtwFQj3FV8p9I0E80pRuYdWyRVRHZ4psqIXhCYKvlu1LhgtEqt7JltjunYvTzqJ1t1G0J
nPXVxgMO15Sn6B08VInsUvzUWjgIH5GK+vx2hEh93UqC45VE6eXldatrRY8OZHhQHEoi8d/PB2jh
jfiIZzAngSf0YbFsOCVVZa9VRaGNazwkApTsrwYCOG6n/HCEXX+EarJQR85eKaQrDBKiCm/VHaQ3
6NjPnu8h1KwvUumzZC4guyjpYPjVpWmIyfGD4WC24HI338SxmCKqf7UwoaL7NvrQGb14TR4mGh8D
59WcdXB4hwJaspIqf5XVWTYgR9t21zTMuqLjxCs0lTlAhf8mRTGiz1OLS8uotuoo2ekZOLmkfgT1
D2cBJiOrPDfW+cQynw4OvXYRbKkYp199BkjJb3+zQ4H5vV6pbt7V5cvJ/EDMykbd1Mzk/gnyrUSQ
atFVApRdLFUmsIFPoQZ3lgGCaJtO4+MiSOBpK8PScG+o0Zl42sdlX3/k4ORSUSwSqjffNcTlQWxV
vHSVOyhDuC9P9fAhHJw50q9Thl2SfTTN2fN/CF/m1QjJXIpbwSIE9HmzMyWAlDL+/rPSgGKuZ1kx
NHJQG78FaYm2lt6Xn/Ho3bfZRdK1oKehCs2ULc4wZ99UBtLvPw8OLIaGUe6g4EJH0dvB2icWekUD
ZzuZZc3XSzWevHSIrzxM90G1WgecuRyxPq3lmUtuEMic064xVlG8ZLpdtliW5kBoehbNsebJrZyV
tqVTzTYwnx+iEXZyCNpJKuG3Z7ITMMObc+vPQFcLqifEfP3/GE4euO4Lh2jt0yvhChXc9qI7msm0
Qf2AX9zKjNEC50MQIj9Ppf/uXYs/Qrk68EAkEitcKgjwe+aqPUvs3Q40cJrp68f3P7oFtDTIgvet
0v8JoISsEBwpxXyI3kNb7vnKoIKuLSTcFvoJUUD14gmbSQ5D7NCe1hnbw5smmG0Zs9pFC2nXnNfZ
CLybvdQleAJSYABseUuRSh89DoSdnEnp6GnmKxMibgjryKNdMbsF/+C46i3k9jDRCBN2uBksy0tJ
0NHRIyKymty3auKUHtBovxlk52CELxfX9UIf2X4D09NLQKztDCxOpB0M6kJFBmeLdydbLwnTafLC
Ax3jli3pPMRw20LGdnK3OzDru7IG6OSAqnnu1HDhjHXGW/GSOTgBMAzs94//wWuq7oFXMb4HX1kH
eiDnkpXYY4t7L+rHTlO5XJUjbemqWMYyauPlApBkFQhWZexg081vBPQRqZS3JUAZKx/aEc8z8cxy
OYws1hJMW5SIyrFV3ZMyyabdUWQb5xfCubSpBBIUzaRYJzzf8y3Wit5uBbX0wU5G+IULnoQmWivo
u5TStEEE2FfpsjbWegzwqQ++z+qeXoT6iaoM/nGhe21/cls45+QFrzb4kSw2n4b2YZZjTNk//bie
1QKfSTUZ2vWMKupZl0jhxbMhfgvMfpMrkgnlXq7ZcoCIgOWClCft8It/ua6NtM2irohT9hMNuyNO
WII1Em5j4ED5Fu32wqodJ44qVD7vDVA9NEeYRAMEYsvDzvhhNVZQJRn29oegF5B3cLYVAXY9S5Sr
HxkwWL6xtRW+SbK7bFePe7bK68jK4j2vB0qvNy8lhqX+BrMhVDG8CXW9JVtHoRnuyrhdgOyDH6B/
Rp2Ky/Xtjxvnkw/IatkDp/m3AxwImBUNuLFLRPV/KljjBSLgaVN4QrzIAEsQDlzRItje78eZ3jFD
8NQcrDE49JkgrvcA27u3hINkvdNqP6T6QRG0L+yzSlCDf/QFTvlwiMCBWZ312XMARAz9ZJCSE4Xd
nhoOZrSBLTHZkLFXHj3eT00+z7bUnPcVKvx3MuGgnhoy2mIoPsE8vIxL850u7af5qZvpMfSYG7ps
Q6jNf1nZb/P3n39pclJ3e1SxeKV8tlhj5JqDqbybgz9+AgIfHjokSl4Yq7OiLFvT3O5ADWu+Pa6T
neB0WHuPNb0ZDJW/nkww5RCa6jvbr6Nslc2yreSMvkWyOqw0wHG+LhWlGs2ENWJL/jg9phLQMpgZ
jcdbq6NJdbkkqhx/y/FAhRu+HVNnwn6CsWsgl2p/TWNjkEuuZlAkgqcTE3HgSVgZL5R4Bd7rwzh3
fA97Bc4tcxj6z7r7GZxy3wWa0Ft9WgCpg5XDolNefgeuIpk9jLW7SyU2nS6MQOFIznvUNbOvsq6g
LAeOytNeXWN/Jf8Tyg5BJq4o8GTavMmbifWHbj8kLDHVnv2BUMMFZ0KAj9A49leiuZz0H8Hq70km
7gGUMuL7vW4qHZat9oaOd4djjTtvqYMK1LJPjnnMiPDwI4ymPDZ9d96tJMyIOhPRIeSz8ASolU8H
VZBHaxD1FBTC2dNJlM1xuHFzbLwME+Q7hhVOu/xWvyv2qom4Cy140eyiOE/plgYqzAqt0W2isETW
UMPYpguhf3VDFVcsMqI/XT5vtXo4S1QCP3c7AAPtOx5DQV8AGMFxCLF8m08YuZLM6b+F7HvdKDyc
06ClwSPhmyHMBpCaIXQ9avVU5+hI4mkOArJ1u2nDxoOPIZk1l9TEAMHcHtd4YAAzbRW5bAa3QcaT
14PfTSomaX1GQq560RF9YFH7DhIC0sDneqiqGRi/2zuRCCy5+zVZhsolkTL+VgvV1Q6nZm3wiDii
ePoJgRwu5O6JPS5AmA3efteTpTHO2oGlx9rLKpygWdFvw7wIrHBrBQNDrf0l20FiqwCMjx2fkWsM
hgctHLnzWpC5FatpPtlF4IZyMDd2oZV9FgfOwnPBp5FhDifhuCl/KU0sSK+VKag6B8pzbf1ky5Am
Brtlz5jYuA9ze8A9VaYuP+KaRvU8Y6Sb7sR3/f0vMGXoQO6+zmnsbJbGQXfTnqzP3Yvq/PAjvYNT
GYPQjGsq8SePP9KI9lC9Cu6qqVqVUuza+lozxltxSggH6ySOSXERAZ33eIeSheJ8UUKLekMavf5C
KpUQDeccp/blRjM560mer3EQ2hafrPukAfAc/gU8mYlUH5paQEayiRfhh5ufJrnGxYLDQEz/GSCK
j2wCv0J6icsgDjuv8rpa4qws50paGjigKex8wI/KIBkgXjn0STClDdOiRY1/shUFh8ImeSXSpjbX
OrHvrSL18j/WBlldZXcTS/JhO+T2wdqtqbAkp3nhmHEbKDM7zYJobafeJ1RojcOAzfSuGRS5O/8E
hllRZ8KvwYdXjFNwIPgRN2NISfryPAbOYPwX5Z2qPm/hU4PucN/+vepBlaaHyRb4bQC2rxaRfMPi
4rVCLK4QKIS4OeUqILNwyNyF6Fb3aPBdvvOLrWmiIYmtwcEjzu9I/Ci6MW4LC8QYrQM57wvF97D9
ZlA+hWEy/Gv4Pgqe7FZaOB6IkNF0D+mBpbYessmdMC/3x9IvSnmStWeib1SzZzY8xYoj1wUVg/59
mF6ZTnBE94ZYPEHoQd/mVT/mhNgcxcGhCrC5zta31PDuClNR8xGiQKGaj1iPu0stJu911yF1UXhL
4z0EuHWajsiipl0fwUJezKuUf2WZhUnjnzUPMNt76TibsX+1WgSELsWYVJ+sGubI2SA8gGhVoSiT
nUFqJZ1XTxIhSKkA8/FVzyfY9rsy+1qMSQfyT3k0/cCYQ7kxSZwp9f2zltgv4rvbQiPEaPdiT6lw
ZQWBirMm9HD8EzlIzE3/4jd/d/TgHLtto/S3jNviJJMjRkNyaQSKnvQWoguH7yMHoMkLQPBUPwLy
Sxi5BFSrKq0sIPx+EAeQd2gFPcOEDeqNoPBf55Gu9zvMrjaSHkjbkFmzDJhXCIf06ClyvbQ2kFlA
RW8oU9Y5JTUJoTl0rrb0EDH/hBokcrFBLSFbCuskgq6k4auxtuAJKGgaTW9TcYi4Ntq1oqkxg8VJ
SDRlUM+VHcZLgFhdNzc2kp1MmepBNrH+pRFgxJcISa9gXvYkZTYGlL5YEXjpLELxJLj2+UUMr+Cl
71MAYQPrctfCZWKyorKuy1WQpjmLWMZx1RC1vRNJ+xi35WTmia89L1vLL7f0xaimxD/wGL39ntrS
6be5YNaDjvwSe0irEdp8q7DZIXYehGGi7GUkEiuLNEr2k6Nph7Jmgr7GloX2s9P3uWm+DJFHyswE
mg3gzaJzDjPe8gpH4yOpqlwyETCW0UN3rr9VsB8jcFxcjJ1in06ytxrLfNT05iBvOefY0U2WvU68
qBMmuq+KN7YKgMBTSahEaDafMu50U9HcrP1r+WDloqVtgZEeqhKIkUBenq7ravu6OlYXSR8/gzhu
EuJK+nt72CdjLSlNntoL3iPR0sUxGH6z8K/QUmA49uQpXcXAaWtCH2vLQh9uWqpImEb/0aQQDJFJ
oM1Y2tQn+KP2nwOjVLlOroJNjyJjHHQVomZ6JHhJMGWEV0g/kfXcpPj3QFtLuAC22qfDw8FULM2O
xr5rKpd/qnKkMp2o2GudyLRfYGNSYmZYHi9Uh+eH2tyQg9OPyAyEUB4hGyNxtXPJZPjpAWxCNaAv
wJ6guulgz6NhBZ0hmmK5W7HSG8eusJUEWalfv1qccdFHUpHbRDsYuoUkGQvFWIcKBdh07BqamyL9
G2XOsYeuR+tURAeWTKmFnD64rf5nbsLAUPS4poSO3evte9mz5IQ7St2QjrhmD6oNetFCKEOkcp3U
flIlz++MjT3tCuNJ/CVvLoJI3zzMLyAmXCrjC4yLl992UXJ5ZdU0sjzT2s04QprsDpQz8Dxyr4g+
Lb7kBh9bHmmTjTJwoyFMu7L/yNcwCGIsz0Yw0Ba4R3HwVzdAMV3kQlXF+TIyS8Dj+ahy7bBZuVY/
09/ByVjW7WqPiYkXkyXJscAoGMBvOv7iBgucyMsrs/JTuALsWM4+e13zTRJ5UFBxqi2Y2o/Jd/FF
Q4aZOw1U1Bh3sRIG/kL0Ms6ZiclPhjHnyGeAdzTbHLCXqF3K4utSRq12B2qAQ48zZBEq0HW3AK59
Q2Xyu1P0nT1YkP9yBCSzI03rUhE7ekWqrUq121EqK+UuySYXpin9JZtz+whOJwHoVTSVd8ASZiOb
WEz5JrxMnaMBEvmdizDuRUtV29e2/AfqCeO9Wl0kiNgJoujMVNriiX2YyEFQ9AZCZUT5wkVpt875
qmPP57d2LO43yFJa0AZgsz/nlNXaHoJ5CZriqQxPb3P236W+KeYABWnFLRwQV6YkiFkqfDYY+vWI
apl6LvnRgD2qn+DH+M4Fs+PTZMRVeBv8wz5ih1MCAZBePwWg25EyxnhpV1DRjjnEqUT7uzyZrExx
ntRbNukV2Bn5Nq7Z1vMn/2CDaQj0v/e2rh8AM5X4mNzSllBKBWlz/PxXJ9C23+TYZwluickNXaI6
+oyn7BG322W0pzGobkkl6hURg/DQ6khwF6BVGzb+kM3W6xDvusk0AL1se5ShPAfA9HGRuVkSSALz
7zApNk/SWm7Pmqm+DoZ6Nh9i6hWvQWKOU/x8U2YN2L0DdQU6dRHPOdeC7mczLNoN5FMfyPlPTD0u
Xl+QGw2Kqfk2vLywIvLFKXBV3B1pgTlCyQUMDvk7vKr4oHDXRK+U8u34D8NlKNBpPcBLntN7I/WK
9tDRr76tdXDHZ7Sd9r0D0P4gjrj+cQVaoG8b+NpCSybzRjM3l7F01Y6DkdBZRBAv6cUQoUZoP79v
ZaIElArDfWHB+IP09hi/Sq3XZUGAQcmS27hfPeI2ZiLLeXBxWCEiiL5ARmZMZx0I6RQvc/iaHduv
9zOdhYMgvMBfLco0YX7//jQw85MjMpag8QkVkfL+kbBAhjjIUjLyzpYuYHfAaXD85wEG3RSvPpTw
VPhlQ8GYqzlYekiRTCkkKR/fiDGbK/1jQfxWq/Vab5IbnzMBDxMlneOKCHe5r2MphH7A3CwwZCt/
xRoEY5lH0LiliMNLuI1gfiuTW0koQm7xO1Yhqk8jRxS5OxPhR+H+0sufyqGm7I2fxUjRFCamEVG9
wP1nxXx/AQwFvrhQQBi14dGS7ikj49Wsic2v52BuGkL5gQOqWuRLEjYjD4BNIyhJNS8/hDBM5Hql
Tm0A7nuYt08MQjwR1X1r60wFnBYFISYSAjwG8n5ESVy170u1Fsu1yVehBKCyQg1pJxwl7L9lUhs1
ROsHWDwbJiYiB72QObswAM/2RkvL3aOZJxAqvlxc2Oql5IEjYd4mEf5GHt9lcq3U6/A73RxtuW1U
1DqUDZJ3Q5TdCu6vfqiAZRZtG/jl1ZwwAjAl5cvGpEBRUCabV/LSaQUphMGnv0CtOce1gzeP/PdE
BxQrgkYQ45DEsD2/3WnuV/juz4DkuAh+WXZFjSXjjva+2TZ0B3YQpRtujaQ3r6iPgXS8csPg6nS1
nz+R9bSkK/Y6klG4WiDHDGcsd4Z215nSZn4DGIxbb3tvg0stv4s5Gjbnlgn64Vo6a47KFY5jrO22
USDbSI+5HGQuHHdSAI84Aj+NsvzW8sFZjFtGuuz2z9GkmkPUY6vzjAB3Kchh164vdBheUTzulFkC
PJwH9lMNLChNwcqtcAOmrCxk2rBprBR1zPQvpecXePtij1vo/Y03dobROUCzwLV8OMmeSkxRsDMu
7FsxE2XsWMjmG2eieDu7E3XKJsCdoVCZnsR2IIXvChuvv9fak9mwsHxVAZXh/KSA5V4RtgdgFVzp
CLccOVXjEo9GFOMo5TjwRGRfNQGof79q44bV8rWSwUO7QNcQ2eD25WkrdqCjwPx7G/uO3kOY9Xgl
TxpuHH56lIA0XC+lwt7qUa523u5okztr6wMvS6oZRv8H0brtlOx4/7TQy6WtYUVESfxbRoIfRzea
lI+HUEUj+D66FIi2cdiw15YlFf1/NMJxzd6yM9b1eG6+EVC9itPpKO0YcvVyHnWWaWRP9zHsBhqB
P2mqxD57DBa3VVnyvnnEIYoedMKYsLv/2NTeW72pplXc081jT6x2TsHmGkdhSPN6ENxKRRMhy70k
uUSwKTChgI8aYhKlIlDfzBj/UGlyO9iAeH5sVZD140TaARCYWsR8GA/sUIa1lTER2Qgu/sJLHOeJ
KcTqK5CD6VIbxUh20mtJrCwWIajnOM8YSS8YW/VxhiocTnMc5KTF0UykmR9dWlTJp6rFtRPMjCRn
cIg/5Rx9rZuYLuoFLxgJDJUuifTU46cJJATlqwyYLkdGRwarSqPWVEKM0pYS82ywNsmPtve0Wyc8
w/bvvw2B4F5T9mrVHYwK2fHDZagJhUvK9v8lfhUvctvM+EYiBoCpE4dR3NRKs2BBMSs/2wpDO4N9
DcoJAyPuK5riHgIf7+S0CHfOb+D46iSF0Hrfrb9hUNz0VcylkV3A3bGO7re5Hg62a+LzvQ9/r8/M
6mm3IddUiUGgrEpM8jSDR7ZWs7WTxdoP/IQUdE2t3L0l2eqQMcSRVIniLfuxAWzwUf4aHqn7ZYrt
dCiab8pFsEEECMCAHIOrdA4Pgu4UWBjZCFmcTO2+W3dGlUqANEmIu7FvjpmsEnXGHMFHqVLTVNK2
GquXSCqzjWn6GFwX0C2SKXCMUwvhLs0cqWVbYLIcv0ZhcObRv55+ZLdrY+DjTMmDPMsKGm7VrWss
D0bSbeXgDuxTSbjDEimV8Y6gQ2ANHkLkZdxqZ9I4+RGK1vkgF3hGaD09ShSNZd1H4CqXRmvreITr
ZwV/vPBDwpyNBtNIYyFczoUp5Rkt1f2k2tY3P81oM1e6mKPy9e7WewzdBNPq2shaPTShVtzuXYzz
XX+js/4i1zqr6VZ9dldHxWKbgvweNI/W1ikweWN4GVMFkZxGADmv3TQ152zU2YHs8SFKYH03JeS6
/g40xE2NbiIj1W5b7kwCoHOlPt/h6/vc+mTEcr2iazDj+pFkJNbqoOORZezho7RSaT1pngb9IDea
Cfvj5BRMeAQflXrJ7Nc0B343rcpsxJso9Wu0bU863IhwNXw9/Wlu+yEC1IANb6ky+wTQbHhXCVI0
/5gskWA3ovKQMkTJVR6vKg7T4lZv83Mw5GXamCMSwHfQFmJGLJL0aZpecHTBx+bbK96KcHsKDj60
BjmSacY173RkpeIzhjkj7LRvi4W/P0GGNkI+1mjUKGnW8d9uNjYOQyV4iPJpjhJEonPu6aP7iEFH
ngfIGLINF49ix/oibPoKgy8e4Gneqwy6TBCwfkqialIpTtK6eM4aDxgLs51MKQlpBYbHhwPlmhKd
onnEbLaLdppBXm9i/t6P2MywRT6YxaxU8OVcKxWcka3CqyWou5yN+CT7f+hpd/rE9Z/A1UpzbaGz
oUDdJl50xGZteld/Msh4TDaAiv651mg5Bwr0tjeJoFFYGEb8rMOGtJ7HwRNcH3iLXs0d6WWYDCjV
N1zMXabePBSijH0BVMiM1DWW0tbcbb7Bcl8N26MDGW331gJNC9Es3kTH+f30OOCHJe6RKunNEryK
acON2nd96r2wAL3IfgTrVTVCpi3McJOgzXmyjsFOJCtVZDSb2VvN4U7veu5SnIVh8ouaiqdbT1qe
k+zJeUBNPpo3E/lAfmcUaw8IWbbQRkBr8Iw3kbOX9LvAb90WvZ0+6ssJsmixjf3ksz3JkEnKRGWC
yCKZ6qQnvSkG48kRmdC0QEpp+RGe+u9SOtHrDoON+BYo8t/wVqCb/GKpg9erWo1BZH3Hb8NiRjpd
AdGftizj9BVcwwbEkqSx9ilJR7GUZIRx6en5AThOzMWkE26IHONY+vPbTdxbMnL3F+vt/2XjHodw
dls4UGGKmJ3GmZHasbCp6cx82gwoXJIzs3I8oanjk5rEqD1QoDu05MXi0nQ1Jy1YxKc0DtH3u9tD
coYxiUzzn08FuPx+AVh6Bh1QS6KnqnmN62kwzMRYOkAwrj2ZeGuLXMK4PIZeLZbKM1P+pMK7ozZi
RPxOrFEiD5t5nm8qfNgZFmn3bT1RC8Joc1riCCPKqiDq2jBs4JxSEGtUnvXgyAUtb3WOh5A4i1F8
zRlGZJpOl0U/mJeViHHQN9+zv/wZ7H7ZoEVIQxBL8dNN+sbLIJuabfQlkksiiAlaaAIw2uorDD3t
lzBXclUiBECkV+qt/RQwghUaFnX2AzpOXD3AqbD8ADpq6LWNSlme1x+4+KuoWj5mBTLJbBBC8dS8
4xbDPkJBKRQ3zq6bl7P0SURaknax5gkPZ52eccYLdnR0AnMfXRE48JJ8hPvXwTInb+VxVVUACyLb
TI+TmvrAlE4VacscxpLkBpq35npPgl7rpVB6QiCDNyh3Gk4tfVVprtEZu+qOckLG31vUPOigDKA8
OvG+E4owRuY14rVxdYdCzovS8vdlTu7Ea/OdyFb09ZflLRE2Vbluro6VoaLvyXoa/UlqRgaX9F3L
0uN57e5+MtEQuIQZonqZK4laPcXTnmbrbHYFyakKgSgIUmbWheEut2yltGV1TSureEva+mHLsAJ8
T9sXfOo8Z+Fwin+nkvrUF8QzoZlFDoi/mA/rQaocIYnb4zWCZF680m3fAw9eHfrvMdqn5Gn2GX9M
+b5TYKE+OUrAvD8zNWbfJCL4WQklCxNG1H9o6BjoAvQnpXul0Wzxg08WF/4UC98l8GLqljSYB8DF
0lgFz6Oco0CbmxZYMCAOBY60FG3C0ohTqTdKt9dr3w+2kdt6545kGVnN5NhyvuI72hZryXmdfGHL
uTVo40Ys9Mo3qaW1Wy3ZwLgrOEdNJqTrmF7qqkQNfJYCK6lUXuy9TWtzCs6SPMMIN/zlWyBLFN5v
QbNKaln2t6qdx8gxFTb/LvC/bGJQi5p3I8bQrWTEF5J9tbhFBVmn+EXgx2x7JuCWIwGXmbhTgOH/
h/kV4ulUaJnQBeRs4niWnwc8tBpYSA/oZpAAj/1N+psQthbOciCqwyfVGClACJo04tmXxIptk1Rs
2oAcHe+pEozXEKrpM+nkaCGiDrDtzq2g/qbhSmJzyi2aQdn1fm2yzl5KM5us2qH3aXNAMh6it02v
fishJO14Ea3lJeiAYuEm9+Vy++xTKx3UeFzHDur92g24/XXYzO0FUqWH6aoHeUZX5oDibOjXmglF
maS/ceK+G3KCqNCjoQGhziZV7MdsY9nSWnmZyXvHuw/dVhJ2MKVzRoI9E3+0oUQm9jEf0Gp6H0pJ
7vRcGF/XF3rrltiS0bKYhrE0UfKMRzieylXsbjJar6iB0vRPktyKkKxSHEdAqFkvSLAkeWMaZ2X+
JNCFIRdQsXjgryCp5gwoOr+sq2PS5UlHI8k9x8PhYmq9d4pI1dSEmBn4fiKuVsACpEMabh0bpZr1
Cwz2RwGyULnfwan1jjTbWb2fL9o4OGj07YM6+f6522079+qBSllLxi/V9SAByIi2LHEv+ucGpw5S
lUuQRCsFWZypCXomLAXwJkz4/WGt/fqZhUkRKISyxTbiBJLENe0woPlEK6/7HVUuPYbU02Nv36VY
bGNi3sGRVQvTvi3uHbAViWXIzPz+4FguF59PgPEonnnYkn8C6RLeZ74XeHhr86DZG7O4dsxcLjoZ
kOne0ZjM1YZfNkCyoKZ4Zdx+ztYXk0l9LXA+0zGj9t+FmW4b4iLE/YANnEZEKMAYlpgEgESjOS4C
ZEFhbsYVeNnL5P1cKAkki4504DLW8DEW2wcjj28fmxUaqDpGNVQwXUZl2bdCVuxHP4HECsws/7gR
xsxZoHd/P3ZdwLHTEAO9xlNXh3DZOTpkBrCVbWT4r89UN3WK7zNUvPT0AWTFxmhTj3pgbCWOx+2N
hV1ILYSXFw15fqKQIzLgOZPF2j6oF/P2GzvnPJ7Iw6ZG/zwG8fiO4oZTyBlAzKfbZOXd4Fg7Wy4G
kVP624kNlGYmkqyYanMV9+fcg97F+cvSD/RomDNqUCnthdffVaM+kiNeEWkhS1f5fhMFvGRhFRZr
req03b/PIU8TV8mtL77ErNWK/D8m8pC8pBvBeb2OY2kq1/sqsTUeW/fVaIFymmYMXlUZwuTz25l8
y0OBijhvSnatJu7VHx5CBCnsxv2vFUhGcHQs3gNjU5qACGFyaOPGZ/dB263XPlho2Q9ABpMonPQ1
IGju0BOyA+B2O7pNn9hAVPgXjbz7KFz/miNvVqJ54lEZyiAuE97+EF5aekoW0SI3Ti+7NKyrWpVe
MOoy4IJNqk6AfvSe2dsfCrE5XtFAKCf+LilgmHd4DgqzcxR6BimDJn6F8Jwo5QFl2nafzLsXctRA
Z07A0+Zgj13xJRrtMNMK6RUNCpTEppntsMtNZZN03rTkWTCgrUw7SLIZBzunaQlTjs8620wgvDXp
kKd4+4EQj6MFxDQ5vThmRM6ZwKcjavLrlWRjnwo58DOQnBSS8M5uVC3mPl8y7BQBB2+xkVPDw1p0
JEuBQRxUwbMB5+VEWP4OGH8r1zYut/0eJPD2whJNu7HBvjj+aFs3BhhOMfgd8PVPRPJ4BLWj3/2B
X2zw9JreXr+9hFmjUV0KMu1JDgiRJ2A2Ohbs4uS+RCFMVBJk8EJSM32Ev3oEtPjwzSgehjIeMVih
xfv4g/Y+s31lYZ0WRpq//vJW60cWIjiI994Q3VMMai2i3WkzHool8UilI69r0BXSKZZuzOqrjo2n
b2VsxS/vIrb0yBhCyDeHldSLE9RbNiC6caAwQpElK3x7XvaNgH6IdEpi/QYBqz1g0z67AVoEO5sE
x9KyXgKo4H/7YnPWw7vcIMeJt+7Qc4nnJIT3iDUDAM04oYYVNUp6aXHkpc8STgljqZfxqKtrIZbY
louH+UbdBqx45zOe1TbKQ8cg73uLxPm6dFt6tWd3nUOAsi13K2+mnWM4GjnzUWTye6p0G4Yy5HZC
1irr2AOezHNQZwO2klwbt28TuLDujBG62dVOLQklo6MkwBLtzkkJ7Ikk3eLDqKstkonsnpgDeSQ0
elils8jTBjuLwCwEtIvuA02JPOLkxjD8uY91sGkX0bTY92yzPoMBh3TnnPIZXVpj4RDp4yp7Ma0b
yv1hiyJRSyf3cBsE4R3TRpz/1SMaLMp9qJ2Fsnlu953aaXSiuGNb3KGIZ5nehqRS1uDsFAcyoy+F
/SR1rwjFEXL13M+igAflJgR6e7zA9uFSNp5BAsokv6e9lwQqLFcCkOC5RI6gdqX3ethg+YcIcohd
iKWlN15/cN9NcmF21qeTgRqXcKRl8QTIDGeVno0QN5TG3MDrXxDvgIynkaKtdSW+c1vWVnmGyjcb
uZhFOVNLoPWSLjIOvkxMdxUTgciSYlMCdTBPJULnO1i/tyvU3sifhlJMdOlMWsCgpm5RThSCHlrf
6hyXHBfiumCyLKQbIOQhjXbUttZ8CUwFt5oqRORsdiJcaxEfiwksA9zzStVxxwHCIAHxOHj3RSaL
kQPP67ebotlB/U95f+n+j+M2LR3O8maKwTaLMcoKxdB/Epe7o/dAZfqUY8ixoOJIicQjISaiTbTP
MMmD/xmz2KOdJndBfRRQA5WAWWaXg/mTlKa8u4CXTIiI9chi72jY7LszIVtwy5IiOLb8JckiB5gs
aWq46RH9O61MHTyXHWDdyI3a1M/cMxmi/0b9sky2UN50qGQlO3myiEyhUN9L5QRabrqrQ8CZhVik
gzxTnfTgXmpcmpawCYrRUbwjVigHZUWSO7t8/YwIkJ6b6pXda+ov9KEEZek711tPTPvnSuxE8t/9
3UPDFirJYFEjE8tx0cog1ZFv/jLGE+Lh3kg5KDxEUI/RDVo5ZjFC+jPWagvku2gHqXdtIC2sNdX+
9szSutH+4LU9SgzYzaT5dCvKnwRBshXjTEP5nFYAU2jPnHhRn25ON3JitapouubJ23XGyK005oHO
JELK+7TjX/ONrU/NtbdKd712Kl41kEzxC9E4OQYPiC778PX/ODkLGm+D/iPSLxZLPPYyQNDb006T
XMN7WslxOvb1WirPBYI/OKgKd2LApU1E80N2topDtAkMJK2r/Pp3hQC6kzaZRcwker9nJC7OHJGV
fXDWRUixF61MfKuy90oRbKgqL297dm8AqvL1f662pj2yNHFNZi4ogEk33WR/C8ara4t8jtD7kKI5
pXdX9O1MJqA+QYSsaFEYiHG8lb38/CUGyDMALxZ4RSqyi+ZWo430cK1juurgxI7DFTu5LIBqSepF
dLrsSiyUWFhSlm9Cu3NqYGc8ObcOqAG4cwfG4uemfmO21it1933CJ+Z0QT6XVuyLoqtC/t1S42CT
02SWadchQSWgj5AGceRSi41xu6u+B5Iii2K+W8Ntsa9zWU6zFQdqwA2ue4L5d3/NedytLOeywAa1
F2zZKTte0VOzU296GQsNDJ9F9/hrciBlQ+JZiQW7aTLDFn1kdnnT4TOvh3EbiRiVdZBy+5BC7MXw
8b5+XY+VdW6PUlDtuENOt/9ws+sIH9vG9ag6j5VNLpuMN/XwYGDiFuAXrEUqspfBp+JdgcxfegEi
ZKYBG0ha9jsTUIsBUMvfxiPfYHK8wZ6mC2PjSgQK0QCbNElOsSR2vmTp715BCVATBliqmGjPaEDN
QBXaz5dMSEAoxYGuYSFgt4BpoFhwYaaQJbR1HpO2tZNZaMwLvbnFzotyDKNxwUzTCQhiTcjnKVht
AFU7XmZ/gkiPlyJ5UvpGx9KEBxWFUsHKLkMVHewpSqfRB7Rmdfvm+6nUFC2KoQw//KdQ+NEMdVpx
T2IuwKJU92ebnONunl2z9JiojCdicK5WaN/W/EJ+HHrbIBtkseIbUR6E/imKy1HO38dB0/W7Kjfl
tkfHQTjf3TbIgPYgIfbeUUNw6DaEvwCD/B5G2Fx095Ey+WEjYoczkkvBZrY4I0MGRBFKoMOaZeA9
uHtraxb/304zIBZ1Mpcf1XiNFhXq1TlM1BvK/+bf+ivgNFYGs0CbrO62E67GiZCplgD/KU6eMh2l
CiccNo0kgHlgtngKsA4eC9BviTfLvBN5ALCypDYYe4Y3eEX7Nwz2pr/LsJ6O3tp4s81ucELutBNy
ofOlwQLspSbUj0c7/nIbGz46mL0nBddMtnkwMfeSnWPfPNjW9qLlGDM4KGGYMAJMIpEyIJe68SZD
RFz/1ke8pzK9d27/g9Aj25Ulpoyt0qQqdx2paZCl2CmKLleYT0hXnpAvt7judNuEQ64hOjhhqmEV
NFkPROuOOa4rdl4vxNtNd1vYK+Vegott0KNGQKiAfOWV4SAS0UAFITiX2gQlnu08fgYezKSF5jeh
vSTZ3htVaQ4GVllYRmru4h8CdVcgEHTP8A/01kGlqYvOl34j8Wt14womX1lwv86JL7nxAdPuZZ/V
y1gLmizXiUiKRQZSswWL+kPVsM3UNMqeTu2KnaMf/0IKrIcV6myCaDVzZdwPnN3w0/6qYtmndaTG
enVUtfogXWNqw+0q1v8Ed8Ey2JeTbC/rIJfbzDsHn0SK4mVgtsVAFAklXV8YSQQ+0v9C4Ssd7j9h
OLbeRl4WaVZm1JQVLPqUJJ0mGtiTEVQJHhs6jNIPQKDg01bu0BKn2+lhb+55uEq5OEZk4ZsfL9AS
NBqbckNPdb/AsPd8Lxn2JyOBYiEF6Ee6bAq62MAGuxCmL+lEZ7uTNlsTN30iWJWwFFARE3eyyIi5
d3HDRnIL7GCIqYfdIBENW/c2p1sV5iPnW6+wH498iczoaFdYbg85r1pedlWiw/1WfCRTCSuB/ypI
Ij+B2CVqDVVM8fv6mX/fmVj+JvrCD40WX814NzWiCF+ByvhD+tVcm9hmRj2Sc9kBEvAP2TJc6aZw
4NtvXuJv2Y3z8S/Osqv03R/lKBXLmoUNMNLLsw0Ia6YaYCXsT2ZeSv52N4h995PPn9yIGG46JLU/
+1lQjQYsYz+gD7Y9vD8P5VjYtLvNScxLNnO/MWLmYBmm1mC2x3kS1hK4V17utSTTua4cYusKBYCK
GHeDSugCP+k8GIKBiTudtiD/SiwlAIZJTEz7tHgkYyPWkujL/4zIzYmwUQZfRpDeYbMLm6gynAZ9
hSapZkLg+XlfTqmR7Nm2Ct72enOatslLnsqK+mwvkdEk5q4VORdvonexF8kltDv87NaRc7/mq4Xl
iJRoD49qJF+Es/0s6CsRcFeynY0VQHlbtxvdHGm1Z7GEnCPhg0Kp3YMaSaUY+MyROkUhkySzwsd0
CZ2PqSL7TDQQodICFhSv6NeaLkPZSLAIRgAK6v9o9/0dAADWIjMwudwKhYCjlMwE1n19L66riSKO
g6FDqjE0VgrgUWP75xrj5G42XESbjNVFm15+h/SKkpL0C0TAzJBYtky6oXva7YEAmL6v/u/nZsYU
b0V6K57FQzbZR8+eehm6zlq+40mlJZlUccvAwA1HPk/vOh/dRv+0zTOKSMAsEgO+kSZL9h6vqHp0
lqeAeYuLYTDhIo6uBAXP+2zi+IP2FHOpubsXLlFwf4cjPfTIa8AZghbRaapRMz14co7UiX+2ArJ9
vvdgBFr7I82N35khO5dYcY79PBYXtreEky2ZvLzTo4UW/GlXvk3YAuBmdU84jsNvHefu+wB55Syq
vz7ko3BABXD2lmZx25D/FeCgZyXwmQrLItlufJzRDJ5wdM9J0XOx79n2PoJaWs1K3cgLCufdEIMQ
HzjClWbFdeNcDRHGvrw89TiPTLQXDet/rpoG/2LqIj7Ro5aP2lj6Qcnn0NHutY5xMvyxevFFk9iC
8JzvEGrSFLTgjTcBJocT3I4iLsqbAW14irf6wBf0Gg//lWfLPqVH29yOCeE0VxsQQ8VcSCGFMt/T
QrXG3EoX9Br/RduPq7mFcIIED38IRCfk9muq1wSskemz64dRRdwXkc6UJZP7Wo01tUByFUtRQMuF
AHum6Rj9v1C63RY9kErQxpdc/ZY1LybNzbsDB/GnABPoz0lqP2SmJsDDKyZS6SqMhMgPs3/SIx0V
1l6SNkNPz3vWpceYk3UliMlpZXC4YC1sTk5fa5E4mG74LdEs53efn6HAi4A0KEYPNtUQpNCB5TSS
Tsj8lLpPeolT4NBpFTFZY9Xv60naMdihI4sLt092b/6DwnDDvo68PoUdsvRfL12tAsh6MY1OSkkr
wX8kfUJV1efOWV9jYLhDYSMc07YLj/qE8NlOTDB0PDZ7IJHzkNbx3gyzDKBi6s+jYHE8474l5f9o
tU0a3lVnlxgqyTQ6D4FvzV9B5czW/gJx2OqZWNTyqe7MQHwDUjX697y84TVctDmDVKtobh0bf96o
cle9BTWa8bf/ofDcXfYUh1t2MOF9OrrD8Afmbblngx2k7z83Ls+dCgVGcxRfBcaAPE1z1hIss4Ph
FHIsDiEl8YAFA7T1jbMOp/uw9zzJqtASCSBKGSZ6oJJ0CC8gNVUM6gK3POpfaczPdODuj9sbkXf1
XZ4uv9+zICSvHnPPw1ec5WhCpnqEwjQpfDAvfyktfQ+1O2owD1npI86S5dVlaLiDtSJiZJDXsIUj
ZYo/B36JWAiCDfWTNrdXaStKwZdbSkTHk1mZ8lasln0Jnle0G/W2zu93IUZwdZ4JwkMILVTv7VhU
sVanq2eXhH9qHXWV5473XvBdYUAE0QEt9qltLoceo5CrFdJw/2dpYiG3ZTX+bew+ygaL4CYv1Hv2
m3gq9P4y6FXbZcYG5+b5gnUJmeDnGYZ8R786StPW5O9oXYVSh/GMlCHbBuD37TzZBjXiA95CKHKs
Fz5kbsf9SlnwRFrOuwlx+s+TKdN5UMs6EnqJ+RHUIGywPdv8V2aAaLB42kVGVlDBQ1IhSQu3M83w
91yb6hcnvNDfesxpnvwFSILCXQds2H69eWDTtGPNGqVYINNwn/PbZysx2BjJ8vVtPwq74E4Py2kS
9WRULQy4GLnh7O30EpKKXoFGJNm1Dm9leiNFq7CzAN5wHH8K4w+Sc3/z8/ldlki+SWregfHj6ozU
6DlDMrp2UJ7d3xc117v9tzGeZ+13T3xljE/Oou3EKzkj3Rq0SAKXPaTl2ZJRrBf8ULGXTo3Ptctq
oX1PwJUEnptxVVA9sWRvEk+c8XkcfjIJWnNhFjhF7803c8PM6poyZ0sJNL1TOQYi42P9zxVOiKFk
Y6yoTagYjmm1gL1MgLi+82oQyJh52obvRZg8qhXTPuNRTLFaxDkWlSVEvlT6NQpdcT8jU6C0Os7v
uYHUR5hGWxkdVdQLoBfl2kUcaUcx+PFHe1VQ3tNQlR/4jvEcUBTaDAScIJqwgfOQWhlCx/Zu611y
zihW87R5oWhirjmY80Rio4MMfXdPRL6H/FS0cIipdxSjqBG+VWz/dD0hTlyvpLzM++bLekSU9reW
SxU5metY99Y8rDn64TczzfnoEsobY5t7mdUMV5ebFQsFpf7LCaG36wAaUN+Z+7RoCIq7sk53L2wV
4TJkntAN24Xt9qFnekyl4OnhSGDLjaC9YpSIan2AMJfW4GvpJszizRi+Y/yFqoQ8h6DxtycI9SP0
8fzV7TXugd9yBV83AEB7ujLkATzXyOMs9j5+aS3chhHMh3mWLD3ZLJ4zYnuyfFL1JXkzihn3f73T
2bbaWmdWhAJcECrbgepe442P8WerrIframu6/NhFUreAhthhGWldNcg/tBSST+qwK36InVZBRsZ+
x8rufmdK5krGJnHVS3TIW0+gKhU8X8cbhZO91nGX4STGCxlOL/vz7YXKBiAZNo3Dvk1uajcxCz5i
4aUap7Yrh2qp+MsscE+y/mOthdQlXgSg81YvMbjIm3RiXAbHC9VSfR1E4+ujaeBCQ4vQusL+6PRL
D3zYGfIak8bWyfZeEam5vE8RqEWXaIJ2G+Tszxfqs35nhXr82zzMDo08E3jzRwY0WY8i1B2e+q7l
SoCIJUuBftzkge3rG0sWw+zrZGJ5LZfrnF1seWEEHMuyq+nMtgQlCo5VOY29It4wvfA72YCuYrir
245fAZONHQCRXQawmYuba89qmOoScmSFoMqOhf/A6TABoP9z64SXpvFPzqTqmuucppHQl/cQdP01
jMeDHECvN8zEZQ255/u+pJoXubt+4+VG1B4Za/poTPsnZXqtLnWbGziEfyg/E8j1yZedtS3RhK7S
x5kivPmTMxrW3R2jsuRhFP8KMkdNFe2djlwaARk8RKIeigDritcG1vlFlkrEcTyenprvBPdUlnZV
/E9pk17azb/KOPa+qku6d4FGBssdTlvkDBlE5F/J1U2NLrJ6cU9lIA/V9UiPqqNUeufBZqI7KFoz
/bS/drutgQuz+FmZZDjxmH9YKZaUbp1JyxVJo7ooUGTjPfEy2uHfwWKM3AwxqfAUfGmyoIvNj6tA
8C4M5AMiHrue82XaiYbTBd+oAOh9ZCbrTftBRiupea4/a7QQjMVtl0A4VlJBJhBb6qsC8Uflh/BD
NetpVfhyfettfcq9As2HYYR4IkzrPNTRUNL8gpD/zLUmDXY32CVv1nUFaplJL066RBqdYknVC//p
l9n58PAXQqx/CGcCZMCyh4CRHRo/0kI+YwKZX72JWI+HUPeQrmhVDKb7uWzob6YQQSn/3Ani2xyX
WKU4q2NFDBsFVwQvmpGMfmnaTcLjZA9Dx1deakwcDLWopOVUXEvDWQOFoJCzVAihyu/SuiCQ5jIH
nXamXdAX8MoRzEucI/D5EUzjm7EF8YRopEyakgL39MuAT4SP9RkZYrEFrp5yOK0Oqg0ak6Ax8Utj
Vs+DsDrPzUyfhy3qUfYc45ZLMrV8F0/iYLWA+GlxCd4muTZdhN71eY+zfU5GE9M0a0cfHrQS2/gU
8BRWpN20dlTeKJQh/nOz7HHFn8qYjVBmNrpQ6HtEV1p/yxM6Q1tibkkXmBswMfDEg0B9G/ro+USm
CZLq2vHRktBGfeCZU0WvbspMo7eta6MUNY0lbwoYaKxfTAVrbHu/nWfqeP/dmYcsv5ii4s1eKcCU
lueECkPgG+9Zc6hCUz8xvAGkUA9Mz6SopwdlZKZoton/LQ+OWaoco192vod2cZki4ILhQKMLOeOt
6U1e/IWi0ufd5yewt87NCo6/i0DQjUXHsPGNPjqlypBwoSajbD3AB1SZSeW8AgxT3q/dR7saL3w4
nUdpbEWgZ8HQOF1FqoQQoVbja16oiApkhxBRdzLBcop6ca9jq+uJlJAXdduuF2FUPCjM75QP//Pn
mEIkRIvFoTejJQFUlP1sJaU0OqKCdmhIGfRB6mJW/Q9691UWczQM3yebNDd4e1v4yu3Lk9XpbPUF
3l54Kg7txp+Mc8+aI4TFNwzgi5iKP3wDxNiQfYWAWCGb/QVsuXy9Qj7fD1xXrR6tZ5o88rtObdf6
kcqV/rnKjDTZNQwZQ/sBKm6B4qjSjlLgDcry28pbJ9wn6AydlpeWuYNjF06S/gXfLbKKxPzW7Yi8
pZU70AIsp8mfuhVBZJ5w7G9BdeP+3TS2xEOMEmIN7xaKfIFf5QjNrvv4SfC/FkyM7zfFwEpigQJe
lqaXi6msH3F0MxVwhVsW2A1SujXLFGrmWgCQZ0kE6iv/wscc5NXNsOvD62RY0nWjORuZyD7URnxB
Urmzz8364mkLsR2MIBp1bPQzXntIQGmcG11pOXOSpJAC51Qopd64wsSchgjBbSlivZGEg/A4Zv2D
6Zz/N0Pm8ZHS/+fLVsYEr7DKrFI1vCLYNDnRtRE80mxAubq30wCnBcUDqW2ifsZYvD+RU/tEWXmY
ovdAAiKLCRtT2pPPpbOzRcmStESoR+kOJlFdVM3+XhyRUPJmbOXJOD7V6wFJ4gjK+CksV8SctpAG
AqzeTcNmUFJ3fs0SOLk2z3ZPFHVc18D/iTq4kouJDKQA44jAbahkHEqJU4LIQDlZtz5Qo15NV794
qXQia6ejF6+2yNBQ/Jya0zqFes6fb3r2JX1sld1ym9wi6oEyfp6izM74nHvW5I7mBfEs2OiYiNQL
/+nPJ0WuxzrPa2GpDgfPdR0vYFFBJltfbQvDbbJV7z7Ox0CAsKgoKd00SB2mrR9wIkra7FdThXbq
BNc5NHbIZDh3nswuqKzrVJ6UXRSe12+wpH4+eJHxtPaBVl3SKjI4LYVxmk8XD1RWcZe5xOla5XbD
5AOWrprpXMpc2m+LEE1Hy3/D0gcOIPA0AggGvDcbVXN+C5r0qLOA3FNO9FkgaTGPbl9eKSysUmhA
9weJAETOgHR34qVa54ddSpe2TokxmM/3WuIZYK4MuHQeQCOS6z1rNk8bgEuIwUiqmqxHay5zf3a9
oT9w3kImJjbr978DrkLwaS9has1UudeTKa+QHehTl2xaTQ6QuqMhv1OC64VVvKlyMYdqWQV4sNgi
95YzJ/njSW/vEKfsCmYAuOIAukpQSh3R9yVuW0XybA3ObwxNAagJSVJhVPCZIjbE51cCMz7nc/K6
BscogtJoLNBzhQOHVApxu0jP1hXLyUG3KLu9j9kYyUJSDiS+E3R4ts5I3GYx370M3r8Hl8evvsP+
2N9IIhVhxdiIIweUW26avBkYmFlTi0yzlzr7M6HgW9QncFhYaQytyZkhJmi56eGZF4vfWuffNdsi
ep4uwsX3QZCbEFUzKiJljSZptQH+zWjuRjJH8SthJ5WOX87CPkxXOIl47pnnnchHug4kkPyniWFC
NZdnyPJyB7knfEnq5z61v41e4TIHFZpypWkiLdLBvqCEliYFqT2vokZrgNAVXAqamDBVLAONXkGQ
pTXmqDqMLUnPshi7tQSfrZ2k9Y2gdisvb2RnBRgiTQtra3IH4mEngOod5TT7tqfdTKBoVlXUW/Fs
8Z+YsDD8x7buuVndatp78zYH/buvOxrV2uLx/d1Wg5lAf1JZmrqjeFYenTz06uGVbQUtnzej45dF
BChiV7p6Yc1XVa0EFkGH9y37jfE6lByVyvVLtqgfzEuPS4noS2NZMeeGWJsitFB0uySS4zpguN9I
IW13fxzX1jPSr/+4DcvbHn3nEMwkX5Lsqu0uIMtVvM/FW/mlHStkzRmp/WwBaCLkbNeT2yHFF134
tGXA++TN1GaCMILzQesdqERulaC4ImDETSLuYymGhSV6TaLlWok58cpmVsyIPCx5edFu+I07a44u
0/JiUZqHGh6d1vkU4rmkmFLFncrhlgIwUREuPShe7kBErAfE8NOMm1vIq4ig92JYghStsP5LiY9w
h6dJTyV4UZhDM+H6wICI0nYViZhRx+7PnpT7slk27RrCc+z2rIDhAhoGJl7+tL/veaPirrvuUZ59
BhgaPpW27CRB/xqY6vvGyA38NpSCbKNEd3eUeDuk5XuoPgptORO8ubWdUQfyNsW8G+xZqB/ZaB38
hkxwPgSres6JQQOuIjulbkCj0OvU5HGq9EYyYtrtXq1jjPSgoSEkCt4yKlmV9MEYI2kx5BBf1jSE
bkVb/pGPUGwShvKzmoQM0s5R57BDdxi+vJMJecsr95pqo/CWbXK4EjcEAs71UFSLpaY/4izOMG0J
opw1m9PH6KzJu63o+f46WYwVq+a6Tl8hN5mOJ5uT2E7+YfGpU5o4fqbCREZAYWzpjoLCbAWkhT5t
E7y8oAeCx44RufGaOBTbLdJc3MRemc4KvKQhyXzRs1ngpR0vizmD4ZJNbd55YA3MIf3xCiWaPRZ5
RtAyF+smNajAZV+t7CIjSs6r8coEAigKx/ttsLgR/YeH4aB0ll205wS47Ew8mStKchwBRdPhS3ny
nCvhkwqFTd1ZEeI9X1+wZMQSlDbhU+qXxajhpTERYJfBT/Pr/WlbKzP5kHOZDbUCKEtJmR/r3pOL
ceBI2qSongf3VHhQzvejNMc0fnvwM4BDTQL7KbbGgH6pVrblQvg2gIl9a3mmliMbKmGCCL8qJ+1Y
IPCOJcP4rm7LoNq1R55+CBYgv0PiQA8TuzPTezVRmWvbo4gvoBqKqP8BJ2KbzQv5ccTugWUF5h4D
uZKyFhyJEhbuHrA3vtWreswEkjJ/gOUS97uCmKgaWxeC/JgdhJ+2QnL/M4emEA4GkmFZ17H+vMwM
Vr4jnP2oXgh97XUgLLQYeHM+1PC0jtaJTctz2CSfgZvi07+vDrqTMCl4f+SvkKdIYM/vrLNHaDJr
CvoYkMNEh+98B+7I1kXo5ply0le8OkWwUNTvrXp7FnywTxISszVjFkQkAb0/51yGQgMbVqkUJjH0
nzS6/xa0vW/wDBd3HtRKs25mIPCah6ly6Oz8rLuw6pTZ286mMNZp6f8Dum8UEQgdCpMJFw8LL7tU
aA0Fu+U0h2TyCQUUeRf6/mF1U4tMKw05Aa56lRM8j7VLvvruUwgDklDeqF9xK1AlmyVtBlhjLMZ1
jca8G8B95PrQADzge0v9jwYAMZVGeePX17HJahuweJRtIKmkYWp5uojP1kV6Gny8BabG4DWY7AW+
p0J3zLoiUbSyuSFveO5A3wwlC+/jhPzUrO8kPBY8OtKdGvH3BLRYLUf2cr6/+6BB4ILu+g0Gr4/s
ZDqLdx3jr2zp4kZxne+Zgm/AL2Sj4/8+wwf6J2fXD75qHbeYTwHWWBq2XZ0rJ/A+OfZpb8iAykXt
zNvcTDTOBwVR4SXnIpW4bPz6+invV0KA+l7zp9hMvsbLhcyk/Q1A+Fi9D8OhfmeflVKrgkAGoUp2
nOHcR0G2E64M9w+CWJ6zU4OOOcmIf+AsVO37TIPMM5PUsHosiHeYea3RNPMcykwhxqBXU690+bMV
Z6yVzEJKyVmQBE2L4TV4txTnzdU13tTPS43V0jNQ+m6ZeOFqbtYTF3hyH3fwIVTXrvi1yihQ0T0A
iQunw64/2GSC5CZGFR/3P5bIZxnqT3qXLUTMD1/bjOziYaBSKT4KH7o4CehQs+GH5WQx5muxjiAK
DnuKimK4ryRGUdKCLXIrw9iZ0+bQ1rbkdYxjyaNEXvy98pi7JXaToFB8SsEByZwTwMLOIkpHjrqm
FPi3ocYQ/TtSlIYmhThnqB5izumw55f0kPTSMX4iehZTKt9LYXxr2MuTSiSXeGwtxCQVQVR/vKvN
A0Q19hVv2Qupui+uQwh8LGQD0rMICVg6/GhA0iLeeNqt0p03JLE5rGM+liJdwQ82lXuxGpTSQv6x
dV1038+CxXZGURZyJy/qUWYfokn1up7UPxY3SUQ9Swq6Cc2YIliekRsxdM67l+oNgHcr8NfExBsJ
1RfoE+MrWbZpaI3wMq5FhTudRsyfHGHu4C6mvrEQqVzQIHl0/HQxetNU2HF4h1suSKb61p+zCwEw
WYQGOrvnS57ZHVhhneqkCXXBHQPYKZumBI2NnWs23t0esQQwETjXBQWTLkilE2pOQs1ds2QRn6xZ
W8rqcJh2Wz+aHYs+6vollQSM2WzK8AabBAyOOm0iEvaOQPO/fxnwertD+ueUR6GDLqcfjEcxiggV
oV0f1mdarKVgSrM8gXo9lYOty5er4DhNA/ebE2+NYim2WDAUFuzSv67abYt7BSuyYsBoZD5IdGNN
KCCHjJVZypXM0q21FaNPRkDt0kFh5zrmG+1DJT9zyKaFSvNaQldg57h5V7hltOkvIJVoBggclcIH
Z6LUfXCm+9FpKOZp+r0+m0fuJGVz/SjHHVvNyDLlkRq/SS6wI+8oF/I8RMoLrbLxfHE51XbrUc7E
SuxkKjJcp9uwb75CbZSErb0vtjiyKM9esTY0/sHtvA4lIDvCymlv12GYkpir3Oi0W3XixfWPr4lK
w14Ts5aTsxWVonEuscP0AdRI5UD+ynLPdXZKcQvHgUC8OD0VUDrzH/6hoIYKV/1KlXA8kwzBiCYN
zLwuz4vmkuf4n4HWFa1pWGEy85Supns4ROZ0fCuoEv4H4CumVVA046HxbzCVn/xUYhhwfPR92X9a
uqfVmlr7y2mSuFk11pKB0gBsW4DYdqDWDYHwER0f7MernjPu/TJvpH2B+KfKOfdq9Y5U3SVImqIV
v3nHLlesjnBjS37O8it0DGNx9+uh42btcGD1pZDXyvrXY6yIJYwnFA8gqTqTC0DE74SQHd92ckJ4
3cMAlZ18eSRrc4sa9y7ce7dUBh6LgcHBcFDhANxAHaFZfTWEyQD4ROLHlIYZ4fHc9JZ/ThZVyiyr
WWLfCFGohLmYt5ohXBCvvc1Q2YYMbTgCkcy47RIwrM7WqUzV0rmgmQvnbWl37Mz5mmAiexJf8xes
YZjoMqQlkmcaXkRQVB69txfTtBZHjrLlXpCsPxKRt1QOhyH24tRm5OrBIwUjnLungW5WwiFazcyI
ivcr3y+RKjQ0vJrzzJoxEviDweTjEVWpwraslOjddHbwd3lGO9/OLdh79zic6MJeRlVS7h8uw5uW
ScX2Pod6/IUigbinHYS9zaA/pPuoiDwQBvWv/lxZP06PcwPgfEqGpqfxk1b4J3EnPMldEdnx4cra
iDl41z9Y3VSkycPek/vxvmbOU/pkHz8gUprwi83EnozIWsSUO9eb2wQ9CyvCu/aIcOkp5zRDAiIV
/tuKDdg9kRkzgpcFLWxDyo9FhG63Wly3j/HcLLOSqngkqw30TsOaX4AMklRLU9g2jskRGNCzwcNV
MjcDMNO8xhsn1MEVTggsuQ9v+BncIm02ilSJSs5Zk8lmNEKRXW+OM1sjkm86eGJ77N0ifiuWbljY
Tvvw7xMwyBGZhpI8ASZuoqKUMn8HY65MDuJZQENEcgLFLgtuyz5A7cNKiGUkF0mILWiB5pgUcD4Q
XpIqUTW22D0quKfFJ9nqKBF2ajhuZ5YH8xigW1ojIKSszyzGDRT/fSyFBuCsxaUmrJtOYCij9uf8
cxecp0zbXhYDX/y6xjupTXGiK0VW+Ttwq4raH0Tleexg5ShWl8kTfY5Tdpd82L/RqU1ChCRTsYlu
PfpPZE1vaqIM4R7iqhKXww5hzl5kdYrjDTTU0ddAKecMgfhmYcXMLVj9ibfA2lfnPc2iEoetj/RG
Qbv4rwUDfhT9C/O4BL2DQoNQXaOymA+ebWszE6/71S6F8PcWqhlFsYp4mhvKWcfoapwS0uVbM7o8
xSqRqU+OSJND0JmrnkxgWcdH2bGBkUfh4UHydDJ726ebaehGaxaDiq5tQcC+f/ZbKaqAiCxb1Yfp
IrGkEAnXlaLFITgvUgqjd4/AbICdOav1Gb8c88aUduIvU/tru7K000as4HElJfEsp8M+icyx+UOY
lOchr7jGzeSUeeNwTbyc5NyYx7UEp8lj13KqFNF40j2P/u7ttPlNcBCaOelynxQiPLFIdOSu4q9G
j+xrOl4dh7GaIoFVSVI4VSopLfmrHZ0j0vvkvgvrJ9aAkglwFO45my4K1qB4demR0S4AKKQClTCd
4wKmxLwVYA9WDwtxYkQhYdUP/QKglU34P4uskmf6Ltdnqa6DrSjxOnXFCaJ13ps+RAl+VjhIMPZb
VnReT7xC+V2w43afMbakSaa/EkluUskte85fmEduUE2OtXl76y4HsGAZ8pVZbGhKiEGH7pkRsCLk
fGlYv5zJSd0b/4a3IuZULRIptRDdDiQA1Xk2K4aKgrgDyC4EiQTX6p0MTLO0NMQ1lAm0ikwxeKxq
+E2AsMYC8XIzbF+gthXJoZvSoZzyzvI6DnBJiZCHL9b+ctU+4jXB2Sv6ZA8IrcWJhsieTh0iK7UO
wRHz7aVJTeqMrT+YR/NsgGBlCUoU7f8EhduoC8qxDynn7GWyA0wKq4RhgGpRkKVM1JCxYdERRbU9
zuvWIioQ4nk3C+OhpvJnSyb2T3E4WlymbPIhS9LHMKYHfyHvUOmSXiwbwniAC1ac7MBbaTCVfK7u
LT1kMMgjymtvebaNQPmftzP+FqBfACh95OTOcl89wmsGw/iNtaAslI3kJ4Gr/0rQIorcOXkp7oVc
ujWp3+fHQyQG7vtm/74YfjufOFbavxwO8fsFFghb+vFOYPdDCMnE5yRTDdjHZL95khYuthlzyzG9
z+u7bArQs1zoKIP0jYhhpqKgaykSBmZu6X5ViBf59cviNPeOXCDVcFRAWN6CH/PsanBJQPJFQjl7
w5tBkdakrcs81JxHslJb0mzGX0U/IJF8LUrhwcjc/mLP8YFuBi1LjO58Lg6GXQa2ZglZkQs2LWSo
WSsya4ijvAn8VJuFhoYbYUGu0QGC8U7qR4VJK6fqfehJgcspRLHlSReJYwvZVyGKqsGo7xzmAmHq
gr8dipOtS0P6J+Zt5bhk0KNJWqtNJ2vld/nAln4haQgqyTdZfV+uunUrYvl0yVer4MxVRWWoJ19s
Gz3IMI9zcBsgHHEspqm8SI38AJCmTstwXSguUxwe4dCubt7azJg41itlsYuAcqXFXj1slaPte/dt
ly1KdPFQ1mrj9CSs9YfUiMCZnW1KGcBXXD/Qw3zD2YEjeGfKHPS28etyW3nyBcPi/Fr/fa6cdzOg
RSyleCExmSI31pyvuF025AMMXJodTZjDQ3lpO4DwpOVDRMKv18qPx/TydWEx0GAfxN1BHKtCcxyI
Es73Pa0TfjFpYC/upixdbN8iBN8qyfuphVOLys3Fu/ad98OsreQGLAI2XPreNg+ly8e8PcK+gdb0
/Mqcr0lVYsAlXdgs4uJFIScCxmLKiTzYegCbIIM1O4rg20DBVR7zErPtRdmWy3XFAyCAnYMQJeVB
Oot7s3nFLQXlWzBE13eTETfo6ZDK6Km3GLHWS0R5lKmN77AQZK5gIqCW1yRhg5245Q5dj9mCeMfR
aBMgptxCCPY/AAAShM+4IUJlBD9ZXfGR9D3YPlsintXKqJGwjAVBHXNkwCfB9Mt5lt6fYBQ9s1HK
/Ljt5OcBpIXAPRxBv9dS1M/3GrOFSMOjM2DR2PQMVHKcUDflQiZUvnHa+rSYiSe/cpl75VeOBitE
znM8Zzt5afowXlC37AeV3sthIqxKy1adI+389EAFpdabIcwVJqQk4YQ168Q6S4TBG4V/c+2Vs+F7
OVRj2qZC7eTfPn+Kcvhlk729eki3FzZ2xrtIsOOxvA6WlY+fRQz0gc1L4oTYQw+sjpNdHhMQf+4s
lFpgtPG6ZY5gnpH8wm6rEAGMj26tQHx4uxSiEDbRiaMGBO7StpFB3VGb1bjftVvpJKF56hpfhfhs
W6Z5MH3tspvFdLVzJfVy1o/9nIVbfQytqpN0MYDaDf7l6TWJq2B6dkU7zzvaBkmg7GSDfCI4bkgV
7UmD81j1aK9PiMAdQS35WWMypruPwYvrqr8WnJf2ZQDkhGd3uA0ck8ME0ksbMOmoQS83FJf8AbK4
VqnqzavXwqx1lgAu6hMgDQg9ABazzaeaLMNlMHJlPb2RP7Wzzi5HtRQIc1N8EmkkFYtNZv0zKxj7
81963Sa5XYEGB4LEHdq56jqbADrJao8LesUuFn4jM94jLpFKaKZ3DnbellOJI9jHmwCWC2GvsrtV
Eo12TyDnHJKj2vcFAzDrr9aVE93XqrgzwvXXvLlLxOGqZDBQyL6GNiiHDy2WWkI+69KZAr5BXDCo
v/9lBv38NAVlWGXPB/8kxsRNhEUqG3u9+KpyWmZjsQumJFtKGoNU28Q7mh/T61R7rnmdXY1n4vEW
j7qY3vOopaAD57DjWWxLOhsPLdVqw3LjxLpqH/cx9YsXXKFDzJeQs8mOmimAcVoGZm84Tf0the80
spPtvY5dW0Iv9cBV1Rox4JyH59y+vcKQVuZc7apXswb/nMPpQrhnIwa3LM27x+2ANRH2Pu7nJfOd
U7x21dT3FTDhHMEeESZMgXbJxf3kgZ3UJnGiTIizZzb+ruHqY837DLddmRIuESrux33EpXcUExkc
VZcVR9J939U4WYqHeYwFdbGBSZS8C0ElUoetQtHj9SMw6jcwd/t6y1HY3Z1IQDdhD+lmvRNTsiWX
tmXr4yfhjqFyT84u3cSbD0PT9RSL2chC0X5Bt0TYkqmucrRDv/epFYVva6T2gl0XKw6XjZHMOrNe
FMfrqL6NZm2jcBM+fVkCrSwzUYcBr0R3s17J5zTffDfTPnPQSlvExkZOhVwR1oQ/dSxHvqlaI2eq
5D26j6Q1VRcnMbVf0DOYcmBhw2QSh5isKINSPX0oah4RLOjaOwxGOxKTohhENPr/uG6kn6nCR0pd
ELL+61msCa0W6UKrKfayljVjIn98sWd0PVSI+lleCxiu3+rU0/fQYmS2ZmSTbxfJJuuJRVXJ9gwK
s83qmFSK1olc+F2reJVOKKAB+ocv9zAgIEoIeEu6S0y/+De0kEXhcgzGv23hR8XxBbvlcXptp8lI
uSx3LvRrHbqALF98F2F/GMlyef0z3AJ3NR5R5fecFBfLfJ9rbd18kuZKEb0ZvWIx6RzXaooPwYcs
qmpXrQPxdQTEV25S4LcaeNp3Rj22cMsC3BUqeANQac3utu4kRg3DNJb9YXu/hjpcJ6owhAYwLA2j
uqE/T2XJNQ56vNXg6Y4qoKc1ssKq/yerH5ddwT0Mv+TlSXSKSqdXiTmtumQjNJkFX+2MNsyuzj+N
JsgSjUoeJuZY7F4905sVdpSJxgV1u9roY8XtArdHXzJBdHYWWEDPbsRN71UU1/OBBD5lm23iIU+t
QiCZRANsWjKjAtwnVDHDzfeblWRVS+Da53ecCyRyb6Y0UWtLHj4mLE37TYZi5hYkJ/mrbb+AUhPv
ZKU+GELixOLYcBK8HO0+Kmj7lN4hcwISE4B213p96PZBqRtEcwJhxu/cBfURAul/rdGy8Ez8H96w
rduruYWsfljPHmtxPSt8FRasWpqPHQ7+z9y9ajySgFieTcfLyRvWLDeXG1yrf1jh80XZuPQvD/cO
05rEnirdl4LcOKiE88iFd35gW9YsHawnZFvFnhB5YBBiR9uWoOTCv/smZNmar59wMl8mGaNFNzIi
1iJEULpeibih/9lxnvqwN+EMJhhqQ1Q3wQ3NhT4kr3uVurrQqb2zO+jM7rXvU9Dw6AU8jGHv2cVz
IUV8uOwfycAyQJFSQNw9UQOE9E3tryVdrZmqipJI4oIYVM/5Uascmelo63gD/ISDX20wHGec+B0d
h4qqHMR8+qTSI2LLwu0ZlZ/YMrLKd/Ro5eF1YQV5u1ux+4u3ItEGXCaUeuOPxFEx/3FHicDrENaB
6oVK4cvJOUVsU1VCS2fPIF6QRkC56pK6F4PB4mwwJI54Go9wbuMZ4QjTgbcf6smGTccptY/KYP64
D9umXfBE+x/aiRrBrceoxKbL7lOrE19atrqGrQXQvXfkhl0TaFh663nc9t+3Xasir5BNYse9Cz2I
42vg6ZoXkPsI24oTdFd8SqZih/Xfc4dsRmDl6ZFgVcha5qbYXa3bHpcrVH59YCISV+dmQ6jjd4j0
AXZcGJKVHlNB2NOq0PtsVMMmkBs+x/SzX1/8wV9FBSCDkSQvrvPf1XxKPRSKt/m2lHtbC3vmCEHk
1nXwjCaFBSIvjXGywFYnNekozlqGuGeHnJVGy8KGNbgXO/+joarQM2qrZ+BKdAFGcmQN529GvPF0
04ts+IvUOxbrxdZNLGd38QePQn9k/kBZO1cmNDoKgaHoO80P98oGifI7wu7iRcfhWTXmtx8Xa7PQ
uecqOH19AxvxXhNgJbcOmJaEvB+MZ0bBKwmCeJr1LgxRUuVRZjZ+U9SAkaRY3nnP+zW5DHHl4Y+X
b8LvhthFdBHJyXVhCYuQ5A5T6lXfh/4YL7TweCcGjvaASfeZDSt0plKwSLOTgaIKXYZ1wfu2W9EB
r5bh801C4U53o3V51vwzn0IGgxzk0N2gUX0HVvYghZqu1d4tiL+rZgWIBLq0MXjKS7suCRlp54pF
cUN09LOdpDxAI9PEMywPvhvwhSynED35Zs0yh5PV32AzoH8uP521+mNwPXYYagmoU8Z8kRW2BJHf
JnUNK6vgQSQej1XXiKvmp6juYYJ76rveC5ImkP2R0C0L0pDdhhjHA+qQz3ltf4+IaAUe4+rjzeHl
/FI6e1YS4S/4ZhA8n/4g4nmRnPljzkCzX6j+MKu/wElrzwdINrdJAqwCSKmL37BVnN1HuEqaCbBn
Pj6Svp9GqgXLuNJF93qP6S0tt3zdHcFIwfYXi2XFJqO32OWAFrZyJrWciSUAP2Gw9UgO2TKfudAP
7R8pV4NsCWnBQaWPLlD60rtvHbLt77paMVM/1V1ODnoVnqZMwsjcCPTXXtaLJFyzAeTvHRBiSTSt
zeIa/7ftWn8KeDqbwuuNbRXdNuRXQ9Qgxmo/poiP9Pju6zuVwnbu02PJmHufvqkTzWs0zb//OSzp
Gukw7Qp/KrEs2P2trKat1O6sSsfH7rrrqU+/E6MhviMHZAhaUddJYZSEux+kWwN6M+FywwflwOIK
ha/1FLqGQk8VrW5Kio+2m7gRLP2oSmTPRsdsJth9WETj5mcckDHVwfLYWTFrUVdxL2/5molwOrIH
a4vPI9Z/BT+GVZYKXqUT8DkKlxEE7xsAcFVxzBhKCvB4j1ET1BlRYnEi9o6f7OR7Q0EQONGLUXXA
jhSaFIhAYci0rdp3PqyolVslkxMlBdt9ktS7qBfAdbPP/dNmXVXQ4JAl0miB78Thof4F0c5299Ej
3MZVvxzBSsj4kkdBVtkSLybievVVEMRq2ohNSmr7va3omA5+uJgiTsrAEcX6qRoaYdTdv3P58rmQ
O8ZZ3/ZQKG8OhSTbZq+i+6cVsB7Ti1XWoS9GEzJe6stFg6uUscutGOiJ5uhRsBRdRi50sUuJCUpF
2dDW34tfWHgx7StSaCjZafdnuxzd+mbKBVy2DZ6MCTPLP4GQO2eynPYO8WunenpXT0d74kcPai52
3e6okDraiYd9qhf4Sh/4BN23tM/IfslpStkqPlhG3fj+O5w5Xvb2eH6EKUI7vPt7eJSA+cS+0zZx
ynl6Rvxob/ZV+WOFueTKfxQDzlB3ii2TIjlkSXISPkH3/bCVWAw7XPU+p/gy7+svK3F3qTAkpmbs
vuoMTGp6FAHzsk0klGnMgOfNqfwHnYQnuTfgVr9DOUXXSaIoWA8UVSPzs4pE6NY6KpM5nljb4pmS
jhp3jl56CLEejdTv0q0h5lMJfRZ/tRek8M2yQL3Nxtc2IYhOQVRQGyAoXY/ny587jCO7QQR/17YS
yy/Glr1XaM2eVN1epLd/v+Kh04Vk/I8kyECSflQQfXudeTwvSdgLzc3FJeTtD1aoIRQmjV0KH//E
51tiW7ioIQesVRJihX5WoGtgwkdlq7N7I6LY/GA4ruHZnZjc9vnf59StWEg+LcJxPEReMcFTYru7
BSIUJufGwIYFg5jRshs8NLHiCChl9hTLzqsybaU0FstOd36SwfhGMMQnoKcFGiNCL+eyZngpJWpO
2z6l2D0rBEdUOlF2jDOTJj6Srzq2EM2pmwVWUWR1nIojL+hX037mrdlXY5pKIs5fCCo8FmYQHQJ+
VsSt4ulx1LLuokXeeesHVo2XAJVNSL6k8S9TZOM/+QxftrkHhX8ZHKgTbPJWmw4VuEMUlq41BHek
j84KJ/H0w5I02Ibe+BgQtj6JxbPB6EapODtbrj999d2Rd6k9TsmDTxl2MnFhYbaykG2qCAujudYp
Ltu9PPdsdvo/XUht87McJ4Tbcd32WJtLfAZcGGNyn/KsQQbr4Hy52F0bdn6lEmasX03oDhY+zto2
3WgCAPIn73kBedddU1EU449FG3ZIVfje3NQwrbd2zBRsFMCyPc/M4gXQSCx/OGvoiO7RR9jEecsV
t9bs/EMMO8VnoqHfNCzQ6Qb2OE7gyxIWFkQ+oqu89vkfp16Bykrey8pP36im6h62GYsx1z3SEvy3
yoa25aMdAzm0gbKQomKz9Q5HXHubdyuhNFSYyXfMmcEWCLVcJDwATIOv5pTxf6CB1eO2O9uaOkOQ
9+jqYs/GhrNe5Aypk0IpZ/Bl/oFQQY/UMr1pu09tn6sSG9idSHM8Il0BU/UD/sTruEDdXfKXLyLt
PVhTjhbCRZLToBqgxlEif2W6nFjKwKV1nwZu4K9TpNCBb0tj17y/XlcvynY+LAycsgE0EFK8/5lL
ie7/nNkHXgvjJBN76BATeuwykcaJenAyjKL1b2GsTwP1l44svKsRDeoZUa5ovhpispaGPzn0+3HN
08qfsqySLJitzTDL02VyChfRmEHIFmZZ+JCEI4lxyQ/pc2v9bU5Wao4z+E4DfWHL6IBYaHtDT5++
mrfiLzWebwMgnXbQpG9QfeEbqM3B2C5jldlFrRxpicIOKRo5PkHR/lS5g2jv0eCa+jvBiND4x7x1
NoKUS4t0kIpjtKm0pbWroYA/VKDSA3N7JrhInw7arKXrZ8xiNUYYzXiUffX9gZOrP0y4czuS67mP
eC6NnHrQZKPwfsh5dKU0P0rPzCPYbgp3Y2SDM3w/64d5KzfgkZ4Bt+aPqRjOhiBsqXr6gCEzsW8h
JBZ2/TUvBIEEKQ2c0Qh0/uTzlDvtMnN2YIvA4NeoRBEkX8xOkVIENiGJ4/mpSgjp2a3b8zS8CLTS
GAeC2BsYL0VgR5DovP6C7jfZLkxmNFL/PGeNLcDqtLp2aJO0f6+LvTn2LLcLqKejlNncgAoN2Mb9
KVrgFXzOK41CscrIZzVe7MA/UceSh/qG+P+Rv98aBxVNb/249Ph6VnmGfG5orCr/jCCZvZCb02wY
fdI5mLMOrmURcVuY6PtdIFvXVly7/gdoIle3V+dGca9YDOmW6RG/ueStvxBUythL3bokxjo5HLYn
MYiD3fHPyOdN0Ptsp0xCzu5bRkcXfE1JAdTMDyDo8i2VBVIhvGFL7GakzgtAJnt/k41gL2fEaTTT
JGJUW6l9MX3IuuzoEf0vkk3kjdJDWIp63iVKj48MupjTF6j+SuzB/VQ6tj5s41Mm+uG+C/d/CshI
cbjhYynJCaCfAe212pbQgQ5xFKEpiNIuoc7dB3QOtnQXt+9o8sstA0XSCB7tJekhGT/Krj5ZRETl
LYo/n9hr16kZkcLp7maB0FSYkIsEQMhUf2aVQbNYVSMIp02rPyDAV1pcDICoB6uSN8vpSY7VNVcB
T5ql8ZHuiy3+CxN0XkjBWOygUT0nd8lEdInR6FnyR5skcboAWuJfDrLIRFSX5yLl3gHrurJh56uB
hzbF2Bgf680DrExRQA4CVQQqJcfu50mNsjrylpI6ZDdB1FxUeF3+8mrMprjbVeL0dq71n2EuIIR+
rsEj1b9mMHuDHebsf5oV/lB0g75+kqmJQD3TcHxe8pd6Rputacs2qbOTDV6+2DC4uQIP+WTjklWb
/5VB4VEdZmWjqcH+judIJPeTtr9c3FPmAWzUOKnGE+lHBBJi/hQ70xbNmFc1dVh483dUkODIjUqN
U29bOf/tDhxuXT7pPM+mzgDJiabb42shT+gRCkLS10GhSyR86ZvB3HbZymjvboZvQVsM4hH8NZOu
rOJVgZnFAQEBqhjwFJQ1YiV86lxGY0iNRKmFfAYn4JYxFx2rk2L6VBxbwHl5oy76ZnB9rYSFYHJT
ogMdmfE2ktFvy7TBCFRd4qlfs9YnZXNaYtZwv2YmBTpLHvfvVlDqdT5PuOWNmuE3bIcfaMhwgh+Y
0oNqOSJMMbCLCOlUEYUXbW2FaoqZDP6AzNOttL+YE5Myhb1hSzDvpXozniuDEuY+3prVOdkXeajp
imOUxRYwQWQvdIFzLtRRUHIDTh+b45fUF2CmyGrZ7YqTQWHZSF3nyB6xsf6XmHuYTH7UfNfQkXls
hFckEvb+tcND4n17iA4CapYhzVMBdD9P+VW8mnpitfTge/57BOQJmZeWC+flv6So3AvPaxchBEqV
/6Vfk5k4D3GmMGp+acAW6J1nxd3iGGb42Dvv9IcnoQnHxPhDHyt7pM15WA+pRTg+Q0iiQIkyUbcB
90vIXbTCf+aA6B42iE+QQCq1FDvVWdnSCjC96jjeSrl67EZjxapBGxu5zvWTMFIzfdvzxIX5acX5
S8TcE2mKPXv1/GdoXgxICEQaebzTHCjwDOe3ea5RbPy1TOfX7JxQcEDeGpVzMvX5DDYjDFME0gjZ
7XUeQg3mMOMyWsVQREyVbgefu805OUGqogvc8fwbtaf9rE+SypNUZHGy+F+IWqbYxOAKvRYipHEc
Vm5WdLw6TQxoDX9+8qk9ddMwZPfmCnZXGwHDYuI+6c55x/J6y9qfjc4G2xBoDCndKvQ0h0UKpF7t
Oj82fiui+K2sUtjwTe3CQYhynHkgGtOFp1y6XUR1UPOHIO5mGeowAGHpehLRQ13elf5KGtcTykPI
J4cVGkwWLexoV7+dM5U8BiRWrGihgQ5KmMbFAUKIQP8iQQeygmIB1HULNwqtRU275dAQqw1k7neR
iA6NM3PclPFUF25RSntwYgyZrWFlYl8GQQsRkdAW8XzedrecG51hlUsFEonUglv8LBfSJ1XY8NO5
4v5Tho5YFPEVBo1g+Wh43LPlX/ZfI+0qizL8agW5q63vDs/zVzEMhSp70b0G1g3KzHG4/seU2xiJ
rVhbGOqhtiaB/dDSUz9pSa2eioq1AQA8FZpB/WF0TCHyflZ9SU+78euGwqf4+J0kaBVKulM29uY0
EhiBQYPAiM5PV7oAAOUY6dXd6SGO03A+I5muKbiIQROi3cv1cB/VXfWyWCttU3qaL1sdCpeL1Moy
DA2wRP9LygFoIMcnnJAgIFEo1D9nYHPd0Pj5F3CaP36mQR06srarV2KvEjhndL+3z4UZAIpoZ9Pj
wjtojBYP8EVP8A2vh6oxW9twsWc6e1j6oFG2pgo2zT/+G0mstoRxegUEU/wSEWtqL+pvBzrNb7Oo
83MqaIZTJZZHDcptSVmL3BFJE3rW4fPaoqsFESdtYjfgEdjaE5Zwp8yNokfiUC6r9dIits8rKrbP
GX8UGMuPdp1D4eGhov0vOfEEE4WxsCY5C6ABKA6v4bZbfk/qCN7dXjGqdGE76LxSp7d2lbrNyRfT
DPV1nel4iXyp8PH4aAz/qFUfzaq8FoYlSTprxO8JE2wGzOE0Yw7iuvqVK9eWl/nB8+0mysTdygOg
7M7YzdEHD+Qgmad4uDwT593fhuaclZ/tUJUw7yDTC7gzujJfQvawSkBr+pJwB7pDzQeBXezvFj5o
Ofqx9Ho5Jugm2IcySwPgHnCTHKKvrEQD2Zo19oFWl1Lq5HdYFlKXy7w6Mj6CRLkZcZA2a9nTAXA2
sfO7cJZk2ao80n9nEzOFmGbPilmM4xECPN2LsMyZ8mEo3VqJr3BnpdXVu58AM9KxsOQjqqFCTqXi
Flsu7HJ6+6S3e1sq9Uvph/h6af4Iq/Rip43wO5dQbOr3T6XONDmhcwZRcZFxNUefK6VFnjvKq7b9
rcufbk1qTTlWq6mDd/WbXiMQYm4vvwcdn4lYRNJB6CZYpGDb1WASH3bc6sJKo9TgU4G7jCPitLtm
RxfCfebVIKt3Nhv4KeWnaGULseWZNtK3BFQHsfdBw87I/eQqVnsQA1ofjTaNkVt3CM0ZA9hGnzLb
pG9DptcpWqIJOZuRW5RuwE/OMj9oNEInlFE5YeIxYxxvt9eJiACVm0r9E2fFkNldDQpvjpkRpMc+
muxW19RoV8k+uCvHtkuV/0iu7/C37+ZhOOPX5AijGzVkTPwofa1PxfppkpD+6XRP1jHmsUgtU093
72KeVQonFzOTKBq9gwBzJ7PbrrfSt6BXX5GvwYV49YfnZ7I044pr10CDdiEsOmgzGWNjXojKgGZt
6Ea9LHYKOysJm2DZsqSEPY4dqc1ehQk1dKwzHs+aVJ0u6pQP/s2gRpy74ZZ2tnXSwW6CPTXETqRc
PLwIFWFEWQrl2enIcHH8whhljLxgjvFWo5mObEIWYKnnjfnhyykESIh0gKSUgHgqbKUOHwonZq1c
F7WhRkBRIPVG2LmiXxQHvu317s6HvsvPdd3d+3VNADBY+SCsGdLxfHbzsCP5DYi+NJ3yycY79Tz9
vOK5aKu81zwgs7I6qKobh8WZBWCTYuSj1hXPOc2OOuFdzPHhWscZYJYZmDGQntbSGtqi5sOSgVj8
BvX9VV+rT5eI1iwtad8VqV8N1v45cJlg9kl/+o9cvs0FfL1NFRqw876VaRKMEOaM15Xp4JG2x579
yjt9357E2krunrIy6TW2SMUuI0K5QiREK9bgn74WgbKMwmuHZo435YHLi/rmcxwXoTi2ZCQb8BHE
yrHL2cUt+EtEBcffWRlu8ETfAS2r/NLBP3enC9mhmT2j+pBcGhIjFuTOC1I2qN7DKaxufu0KIQYW
208Bh1Fch3nLE+a7PvvbFKJHVSVYcSTXT9l5/WTlXuQiKOk1IC8Vb8Cm5DNOt8YFbTwbdMcAt1yr
Kvp8gOehy30TtDXBxbvaTOOYv+BVdd5nTtLreYbdveapCwqgvYT0sF1cnMOvGmqpgA5KhKdRZFax
BTwHONYeMAYO/M6B6BfwfEmkK9quqAKAGXBNryve6ZFopAGYTeC29n3qHgQHkvy8K3zerzEV/ReF
hjR/3pbG2UYgQbuf2W8aobX5WTtx+fj/0HRRivC0bg+wCmMmzNemJ6Opj/eMPnAJKg3Q2Jx6aHPL
2nSsXLU8+Ma/naqtnQ6uDCCwSr3hXnl+A6grNuhYCc6MPjXNVvSbFLDk94ZIu8U4CP2b107qA6l+
icFeEU5qfRUnyH/2DLriSAIoVeeVQdb3AQ3oSft6p6gb9D49bKkbzFH/MWO9xrfGj6Ga4l/RRIjW
2xEsUlEu99jduhpDkV2S4TSxv6b9H2bhTiCq+w2c+sFOevGzguQPMuBcRDfGg1ox19klJ+cxqRON
qCphHUoVmxApvvNQ4uqFmNid7htrsYxnhWCcE1+BEh/2ds9EBzOYUa9qa8D/cZpD1ckvxDnkO2x+
kYdvD2l6CWvxanAQa+PsNduAt5Q1vfIOx7K4OzZVfK2j6tuwDKuNFNiitWSd0+hpFQXjJMV0Lo+B
KYJI+8csa3l0CsZJlaf0jM/maEQRdIYWECWIz6FcXl4mKoR+rrE/eaVuwNKY5oGZvPWj0O27MdqH
/hmzRQOEVIW8Ow/jeQD7PVzYh4ftrEnU4MmsOBUUuhYnd73EvGfB+KjNqEAQ7aTTjEDFUbbBEt2S
M50QdaQUn2qjSFJTZfffGVOtzQn+2IoS1TP1AjhCUxTlOFOO1jPqsMa//PsECYkXdmaBTSShvNhC
AN1Zj9xl+kntgwI5aAEKAyK3RM93DOT4BeHhZ7vrhdZQaAvKIKnCYnt+Wdl8azIpxCy8s2B3pXBP
0sEEVRG9LwFs0D6foJgZveBz+EjNMjRUuUHWYI51MomA16XQx//359/x3PiU+hrA+4RV/sNetHwg
zr0DzvKz5OaYs+RE1LgY765apqyGR/bI3GlaVZ/jukh1xGJQc+B+B7bf8RIUQWPCjPKb375DJqQz
4QMb+fRVwsvKEgFMsZ9qCzfqK0z+2SDAINV//GoLA1Fe5Akb6M9RVS4kT20ETlw0twugYQH2ChFb
e1j8BDvNaShXXTazHLH0Pk7uf/v1gXmHioFu973PIU/KdrGIfKRFP5fhJAFGwHFBB8qMaTOfBLGx
tVBFdLZ+chStIqoCODgXBeC3EUMIGCsMny3rmT5YUdjsipKJqVGCKkmgGFTlNCqfnTkkq+UvuBVy
EQQ4lDHoXvlvpCctrc/vDbV6WZ0buHnI6JlQhk3jBFzk3YCTEnhPPSp9Y6HKW2TPzdfyp6QpEt9d
icHJzU5x3XNMpQ7G2hk4pgzjv7rnmVbt+0apYmhERL4Ir3j7gnkeNgY1LyTY8hgLgXMYpoyoYXk5
8oLliM1xnANGHmSHHOq1nokF1Ov3GoRlcd3ZoaJlwEjM6Yk5mSMZ/4f/0UUOc3HG0keTbF0g3EB2
9CYzvBQeGKzyyzeT8a5UHkfQS72T3czxS6d+NJ7xYMXuUXI5aL4NYZQGje6iABV1yWlra3k2ZOmX
QhL9zQa/QaE/sjk/IEjlD4uBSXHHng5yHTW9RSeqOFcm8582NbfMpxtHmEE+HStiIej3dShwnZng
lSf9lZMF7jIzAxnQ/7IPEUO2gPowDJ9Tdc7CLDAsGms5xFue8WDcEKhmUsPqCsbcxekKN2bOeWYJ
njmudX5XY9+YMfMyFivrLh0FT0JAb1a/sTRbiblTdAltDbTkgOKoQxVPRLsGZWeCy2CRetJHc1TU
FABX8rEvIc1r4aB98Sg+Ig5/mVzY00vov5PCcY+3yuQS5GLM7uNOgF+MCsjlECIkTT/9XtTcEs9I
CMIzbUZIvIpnUtQJqOvb0f/ANsp44vf60eY6zM4qf+62ahG5sTZzR8t7ag2tVq5W/YR6C1s3qCpM
1/R6dpc4ny2PbL1PeR7nHbPqHdmCyPPW//bvLaEt6jIsLHcyUd96VoPwOB3rLmRBjvGU1GlZ2AYJ
cZ3dazKeAgXxr8B0Ir9i3ROOYsbf0vR2pytbZnbaJJD5qr4szCpORd2zfmcf9wnEUSxvxrOzEzKs
EQLkkCnbYn+ToRGecncTstiBWSBVypKyBZLv2Qv+hJ9nS1m73YUDSN5R1d/7jDTdzjOkm6YoWn6K
te2kR5MqDdXzK+h3pLDTwB+ljZtf+7lO1a7tzpyYrCWdytcJVbCvZT5agsmTmz0SFsyhz83uJg9b
Q8r/35hb6U6eSvzRpBI3LUDVQsWFoKLux8EjQ05GVr0EjkHsdM5hWjksB4SYvnHveKHRmhO2zwD1
eo35gq3/facYAEHQ00ZWn+78TjjKt+HPog5MytKmgoEl7PDVtk4GvTblDrh87Lphbvz9bfbzmQEm
EX5Sqsd75LXhPz38O+gSSh6fkAa00QZtNsZYGdxbiWEciPCuB8y76ZloYrAqJ66cO3i7F1i4tRMZ
HuUWipCUlIxs022Iiv7IXUe5F6p2skXF4GaoO2bP+iK86xydzEMyHVP/krHrr8h4jrzgqt3kfKAs
YOHVoONLwlLdnJUrRc30AmbESoF6SPuJipdVyeMc/Wla+x48EtgXuiUFTHEzmMEcGIozCU6wlcWc
KuCVpdzNReM5Dx/dzLk/F/XV3SaGL4ylW8ApXEvStKVqzvoKyt8Mf3WUBx078klr81yvlUBqOI7D
CwsMWLlyVMIDIl2PphTmDnHOqZNIoso5dmvAqJwPYVixNzXOtSMx+sF/QI7fLlhlog9Lug3yKbnX
NQ91B5p3tZ0t8qewe9cGbwnf1dtMK/iZgori8URx2nyqQblOWBpswtZS4TeWZ9NKhP6taU9MtT/e
z3G3+oBNA4KBvDNXi9kR8RUHShXKiTFpC+NxX4SrhV2+DJp5AoG9MOkV/XEQfEcHc1+ERr7m2txo
K8wNUm7NHOgRcsSfajvJMDJImWpLpZFqZjPrVDXr2rXUAWmXw1K3ighTWVAuCALl0569/9FkkMsH
IqVxDPJo1s5lvtbOqsInrCyObIykUlf46uWZ7E6zZY9HhneuE3Z9p2Ex+lPhFCLDqpGyFyV0QFfn
J6WoBKgSIZzJWhA475GRE7KbFakB/FqBUyxVeguuqMluR7bMMpum4Uh3gQ5dgU/zpLIGZXOvaRNx
yRBZRDXAjMYT0zhSFz+G/k4dDUD9CKCp2eOQah2VqHfny+ilOo6C6fte+LL9aY2GV0YhKpiF/qZP
boaEcnHW4Oj0+P7r0jphg4CYgh/HgBOMupbwN1EHr2zQTzFI4ffzs8g1epvmC6MYpoS7cKdWm72S
WNRqzKY3dsPyCKzM5/VdWE4lDVP3TlDSDeCUiYLxko5fDhPbYccxt9rSFPWX3X8BpGkLhmnbYTHC
0T3BKHDIYnuSxvJIaVcQqhTOBXdx+Uwj9yKpWRb9Nl1rVVh7RAKH2cb8z69yu31Ww3HoBSYXNJ6j
KsRXKFpIOeHdy6+YGH5wZ1YEJMShVS1sdY1CpEPCiAaw8vN4W0YhpBBjSKuNkf5LP8/x7aDGGdl0
O5aj/UthgciyZrWaSMxYCEq7oOXsDiz4XbdRDN9QXknBdu5vl7DmhUBGZXKcP0rILZ/2xPOzN7o1
XthcW7CltJhUxvXkaPYd0m6F0dJPjKgazHJP4c6SoW120MNMoUL5wnODthH2FPu+PrYuFOVsizIM
fnTNprQWIherNZSc0qNmP7mFmgfM1yhFzpTUqqlrUP7/o8GBaqvsLnNJUL2EXAKGx+EhRjkX8sEv
3mQkXLSMlvjc04woRbLv8Eo++/dDZ1+jtRL7NDs433wtiWCa8+3lKajQmbuJBp0X10tqF+v3eZRx
zZDoY22gNd1ocL+4nGG2Vz1wi2Y+Lmc5WcLQNfwHP/GxzFLGG1XwjR5zePCQSxIx9NGVI/fn9/N8
61d7rmOOvYj4JEh0kkj93RY4y5Q3oyWaji8giTTjl3j8qvE4LT/Pwee4VkX0sfuZ788Bwk+kuWUd
z+kF3y9MTewgvBNGZfO84Eh8dkhU6L41ysrT7wo3y1UxU7SsISb5C7nmloPuZT5n71PxCHQn+HSe
yFkVh2dI5G2SzRk/FmyQu8f9Omdg8me8N5kDgC0Mz5dmy+4X9pV6vsHAt1C8mtTiWxdBHguvkunu
ksCh2FlJypO7fy5Nv28ptPNI63bBymfFHd8eS20W1rblHvC9HL1zgP0wExRYmCJnqmOaIRIIaf6Y
foSwNvpdcnUdV990BqbCglIZe9av/QYwPjWbpjaWFOuNMDJBOFxexevyjrEafFy4TbHN7c7JhrwZ
llyBh4DxKmIvBetw8Ohn+LyA4ufgk248YtN24TI9R8BsltGIiF8hbgS5HfVY2XG8JuFl4aJSKaUg
hvprTMZ6xj05DWgF4Q5aNlG4nrjec44709HLp4xhKbKwL16dp7eN+1s2Uo3JC2AK78+IiBX5uTNw
QkUvXrRS/QuKHXlbXjzx0MUuhYFDiL6dwOb9ZQqsMGNw4hsunaVnVeIcTQvtaagcn8BFhGG9Rg2N
FLhSWJSZwfx804C6Qu9q45WiDyhL77iej2DEiigqMPOfef/aEajzjLgSIaI7IwcBluOaqFJaYizz
5Wj8CwJCAZ+RFK0ZvA509HkdmZAn07/ZevObZRZ9/DbUkl7ReL+KApX4J5WirLBwMl1UUxIG8bMb
3c6JAo2eUVqhHr3aZhiMyaBgRb6v7MnK+7ozhGXl9aYZs5OUvIneouLA6IecwuS/Fb8XRSD4p7lX
/OHFJ5JvihKk1x5zu3a15NYGsSy89jek4NTrBv/T86Rc0jYY/hrpdZ7tO2L80+h+JOf85FOohGV6
2ShFHTNZGuN0IS5Prqrd1q6Sj2w1cKJR+AhapmoOEKTpjF0FxbZexYKZWFKbb0zqkDLFQcMISBYb
/6vq2h+2nCKwu9IPveXcr++V96CVfYN1RjVwkXC2RJb+9HxGzOuYebsp2MQSFgQu0nOr7HrFf8h8
TtFLc8LlgloOmixjKLlPN/RGJGHZjrAuPtxlmBXcR8Nwf7Dx092yrCn3Eu9Gp2/mOIHq1H/JP/wk
hz5tjUtq67uDFVMcYPCuqmWzbuJRRWjwXbxpSXYitGTKQKNt4GgHI53V0TQMowBtFvXkPb9yqSsf
lUoCp/bdeEZERiIywczr/xMqWzW9y16gZY7uEXenY0jtW4SdgtQM6Pc5OJz2vusDLGbJTAzbtEby
wkjID/xvZwdT4OrxBQjngLrr3LQdtb91LSBZLakSXb4v9AhMgzzBwgdXbNY2bJdKjbF8qCsogmes
BcTH+Dugb793VnsyK/OfkwSwxJVHkqr096vVk/SiCG7ANxnx5zrYudLwfivQf0mBJ15cx3gV9URl
37OVH4uo/Vq8dXQ5buz9BUPCbnoRKTpJkBZeADkctitjCExRZ3HZFIZKR4L2x/onrnfYiOsQqj8C
L+ZzYa010Po5s9m0CbAUh5/K3SEQxVfMuMmyB5aQzNLOcP+pVU8XHi/QKG1Lt8UgpvFgYTHVMkPK
fTFpmU/NYxPbSHprVCFT4cy8iEaWQLuA6LTNQu4XpCIgft1RSzhRakjl726r73ZHAfJmNvhRwCYw
zXxYBc/oU3ZfHxQxoPf1xjOeY1HOodO5pnu//MRX5rgkbEIS6UYE4iJ2uyZm6K+0DPHLoruYaPTZ
7gAoNTD/O+A3Dc748YCDJuvrNS7CkNhcLxuUucVwNIRjJORNKVyckWtr9tS/apNVreC47lue42K1
QMvPWB2aN6RoTmB1ufk7KiqBm0YOPs59MCTBlTCA+XBTN0vXWeC/+RkC3wR/OSKsFCXl6d5WWtOm
YQ8+WJwuaRMEgK7EU8ffZ3qAf6deQHKV6xy8MHresS6DEuH9BU248dvcP7uH/pBvzdiHTtM6zLO6
gg34H65ulnoPhdOF3bI9FautN9XEGN/4ERpiPgtWAjj+G6eZyDHY6fZwmvzOpz60uVxUexRkTaWQ
7CnJb0VviVsQJrrnXreQQTLKUgWmG5d53Q1IsTxKfPTVUDxrgr2JZQR7RoXCU5wxeehWmre0ec6n
kV6tmA4Qm9tMWFCcy7yLRq2P/ZJFL4E8XF4wMxjde4MRrp0hiIOEYfVzb29ONQeduvACx4yb//U3
dFKLwgfELEQMtcL21xLhwb3GyTKWOFx8Kf639tM5eBMyzSYLApkZkXS8KTfc+MT102Hw3cclTKh9
zWNhUao5lnVcfS8UCOJZ0gvRjTt82gFKpPCdIpNGME0XiwcBj2U1QiBBHRCZhvmOo5WkDjlTj6yL
8sF536ppLXGmQfzRMX9JagN8Ij5B1lln8uuRTNg5pXxQCnHsgVxhKySNI8I3+HrcBSz4C4x5Jh8/
6KAK8dM42XvttRdDYD31uwW+S1rHeDjWxD/AiT6UjiHaABmtlhN7gw5jKfu1bDmh1A5A/DJfPfsu
8DFA3kk6BoO4AZrh/VRubE4RS0VcxFi1IDkmTeEFKZTdvb0phzDSUwk7Js7+feC9NAyb17nme63U
lrwKSub1VPuQsZigc+FHeq7fWVf5FENVrhoL/tIJluSBXD3sdgjlyCW9MxjxTtGZABcu403hd4JT
MjCmnuHaXyINle5XhQET9gPTp+IGxiF6jg1Ib8pR4YL1LkoKGFwAVotovi/tvJlGEhiYnUx8sml4
rN/v7+kUD7WH9DelCK2zgqhUVQFj2oUrnDYjYyAdeTZF268OaEumsAb4ZWL41k35nHTxcLThYl1V
rvQzJeIngUvcq1eLCpOp0wEt43Z8zo3W0Y4M3LrfiID0CAZ6V4LjM1h5nzf0EabHyMnswCZYtkSG
pdxikuiWCrAYjBtWqazTmcs0JrpQg8sLveLLZk4MDLnOUgWgjRXLO+UNpZymEYoVdNGJImwM+NqR
ravpKO5XARGGFJkOYrLgQpSWFSUO1eCTdnr6R3THN3csEtGda6l/189WNULpIzRMi+GLAJ72P6zc
dXIsmaQdVik43jPaq1X0quWultJ5inK/Eq49Au3xapKqk0Y0h70e19M52KGcBSis0p9L3G9NrBRy
QZVygwuwGlF4H4T/iAyub4saN2bxHUsSOAG1X06fLnzzHxfOdDT+RSK/JfVNp0mTrw+b2dz7jPou
fwX7SarIEePmnvJpUHNW7BJh5kPXhqY30qtoYJSwOhTjKnhfsfk0yFzp2AjA8lGLGEJU3WAqMscL
YVOAQeWYD2hcaKeJF8tlxTjnXuEI+m5rKgkZjM/HuPeUA/anPshdRwFdGk7jUW3dp/YTCHkUjaxW
6o0uTo9/VJh2pvG1WLSFXCo/T4grxBLM69XK0yLg36ZgG9bc99QF2NQYidROI/+GrI7dYKm1WioI
CRTcRZ78FHzAVvn1WqB6cIhvcwxhK2hDa95lQhcBnUHcD6XhLp6clxiX0GqV9kDk5vwpjkmB4f5A
47RtfFAZpZOZtkf0wF0rvrT41Ha2WFYRVh2EGoYq7vy+eq2ZtC+Oxfcy1fIPXvMnGgLY7BBX4EXZ
kiXcDeg9gW+G672ayEn9HtmZxm8Jcnxp501Ojc1Yt1xgVy7b3k2p3dmVVjEZVM/uEWiQ9TMFtCOs
ySYVJoz0Kf+N88MlUzB++wGdHeoodNP7JkStg6YR/WaJEDJK3xfCa5W2xHrl+R4fd+Pz49ADZZq5
nxOu62QUHeIvIkIw8ECvC4bDvNxItvo4qSPuyoQ2zPzm+Wre3j4gimlD18/kvqhIRRKAT2ql8f/T
W5twVDTU60vuz+VZ6Og6anoOyydm/SagjfYP0uKNXnJyJckZlb8cgRfOAyvrLHM21bOcUpxxnpR6
Q6nHJH5i533PV/y7hnlD5+zoQjPxr80M8jZXkGCHMvck21NxpjeKGDXAhtu4CHiIFlOik0XAqLzN
Z7Das13REvktvfTXeTb7YFB4lb5DnE2OSnObR9+Ox9SoR5WyTd6Z15grpC7iQOfL12t7fByeXYMT
d/8cUv+xAEfXS8Dp4wByi43e0dbPNEG44x3ufstxk0GlgOyUS8nZpLqQi0C5AuZxyh1200yVhcDG
Y3TPF5RdZ8rY3LCfPyPANLpLkRQRMFqOk9LGbmz7S6uLFqM+AXILwL0giJATj/CoS1rAjC/z/QpG
hcQbZZRXxPYL0buwn9y1vm+Ltn0xEbKB2rnCUMT9FkiX4bmHdCHaGkQA6lPLugWQGa0SGAjk3Kfv
Zb7ZEuubzEQKsXPDnjZD3EU+eOHKEku+KvifJUjvnBZu5lv0OUhWrcSaLCWkBWYsKWqQBGymCaQ/
N0zLrkWALjYL1gBHv8pt359wNt/sr3TAtTcOQPgaf5nreo9dBvIKk7rjDZ7ERhUXkZrVBTgKnuwY
WJm7RN14jUWS6wk0/FGp54NxKWhuOcB8YdLr9O5UX80vHEWgcXSbZpEBrRG/Vpq8Df/Rdgfh37sE
CrnHVCsnzA4xmpJjPb08OizsypDdSUuYgeHSwcXCGdeIN/jGvOjE8TKFjpkw07I8JwSwdlTdyWm6
kRuXKzc2B3siDPseBTYs3s25KrO2Q8K50nBvrRU5U/6imhJGRR07wG/D+krHPNQsHHCJBaqyzG73
sF9r+whxcyQq5A9UA3c8Q6YHlYsYlCvuOr2i1K5TfC1Uy79CWtgR8Wm8V8Zc69GrxL9UzWRyyOZ4
7A17GnM8eejqhbk+nNcfeYTxYK+bxlB4sw195oDanlY262A/TC7IzeBoq5V+wdJbuUKl7oP6ABjY
Xk9NC52BQJGfRcLi3c9u9xGxJ5guy0XjiNkEaDoUFoxuvu9iAdKWVa/FmD0zvS846TMPELEkV4E8
WIXQnCGZofu0mVw7Kg1dcigs6OYJ1x6IzWKXbgJk/hBSnKFAQW8cqLjoOeb3B+OVfNfgUuOWxcRQ
Eznn7S38wajdoKOPEtW6xwy+nZcWhrwKO5t6D4KgNJTuY7WwPqNiXrpmIdZ4n5yQ/RYz/bfbg2I6
fnY7tJIqD56MO2kTPSXoLQEJZRa33zeHJzjXp0KC1UUOHyovROjnSf0QjbabsvAFQ6hotNkz5i75
AB5nJCopGswq8hZTe0xRzmuKvV3Ehr/WQnE34mk6rF3zBwHBIZ91GiSyR3Jn285wMIIHlznWsg81
yMUeSMgyONV3tsB/WtFJbwiD2fD8DwMDpnlP7aKAwGHido4vF5dFXKO+3UytOeXQE2FH/7SkBMGT
uXaUHM5TVhsa+jzxb7jjDT9P8EmGLC0iqssGkDxM+daMEWI610USM6upvz85ii37dIyUtTha//gG
qOIFs5XXjRHme6J8qJEzGEDXvfg/7wbqGcKQFOz8rqhUL8j6GxEZaKPCd1KCzu8YnHOVzMXmRgp8
IZ3ZYu5yufdnHYPaT7jZ05byTDTPBnSRJ2m48sJeDE7XlW4K4VFy9EHMoenA5LE+0pJ0fij7gM28
oB+0wS/tykBiW1GkEWDpxWr1aRcqziXpom7DbEHiC5SwV0TMbksbAOyWahCNmh/AeDDKm+UhPUww
dF2RGCmIEUInsHu9i1ar1DCYLFB64BqvFkqMhoAeNw9Gk4OlSngR77GF0NiHqgWpNtgUtaIsydHL
N7y7TiLOKe0ot/m+bsmUFMShqNSRpV39mjMCDFW26Ffvat5uISpXJZbPpyl89eEsXyduNUNXaShK
fLdJ+xfLoASoHpMEoYBgV8F9RihBw6h54/X9vyemraxUjg5ytJUJZPRTZjt43+emTSRFN0gJ6Aru
DtqGa053WJxkrFVAvPT3g0jVvyQWZZyfrE32Dltf70L/ZhlMb+H4dzNM5mX+YJ91FyR6VRmN3XNU
n6q8MPeh+iznzxVryp9DzIBT1y0Ndef/ds5B7zcGxRak5yJk5x+UQrY3+NJiOPYF2h0SKQMz1qZm
ba/3TelXVFckW8yDDWp6m5H1o7+5NOcqtMB6cmPPuvn45UVdWAIiv0Mn4bgpn9MOW5XTtofslShW
MFKfna4E84yh7lX0s8dRqhW/IK4cy1PKuYED0O/t25ZslHsXG1rxn7RxyUgMl07/H+zS6LFQhSSY
6bEEEWMEzauqLZ8ewSYbMBVa1o2sVuq0ONNsBvtko3VadehrG/of+tDCzq4MhTo3Fon1JZDphiMx
Vh7Gb0FKVgyOTnNtRwmKoR0apRV1VD7/fgJvHFLgF1E7T//7q8+cxqKNXrZkMcRbEoxK0b0Ylw/r
jmO3X9vvBiO9BZnID+dYP5sL6PI2hKnRLejLnncsMh7jjTli6z3M49yhO0asqyECeHzPZIFUQ6/j
tJJpgr2NyER+JfI6ceXrNkx8ETrnDqLsVZXq89Nzg7mU/hRNej0rpAD62H+HVeCamvB/ARYmQWyo
NYaQ6RWZnS1TcSS33xlyhszoByXnRlRYQCGa8/0gsZn/zJxorwMMMsi8jMCFWw8pSqgM0ViijtHX
tXfwSRZUuYKGFkfsrNw//D6j9IAFdi5pRPs5xu8h6I0vYzYkTcmerPIPI0kS+A5gAgfg+beidkRZ
hK4shU2+tLnbF7epv+sWGMIsnt0jDzDdh9KxEJbEYD5g3iAba/bgK1J+yJ+6o+U0WNU90TSSsHjw
me15u/GLYadigSAmXDGpo5aekTxndi7AnJXt+w3eHjEpjRTEJAdkoBnhAhjxzCHiTjCl5Hpnd4a1
a2eauUJcjuudgdGLyV4COu8dz8EGezkys72nfADt3DYSJS66usVcNMmKaV+Cnwv8/wRvkRYtv68Q
nRR9zvGGJ0E08PgSza4n/1dgA+egr02z6qa37avEtmNlmyI6TGl/PrkPrxMD2U6seZbmFO9Oe00g
VR2XrxiU2kuojtX5lOS2Nia49jPymeBrIKS2TWrg8dxjre7kj4Z8G7HUU7c3tTvy+s3vAHYkCGP+
hFeLai4DqyAJY68elwUGtdXY9YV1NDMcv1Djs5lWQQDTVGWdFldxvoIwHDrT8f5DxNsMX7wBf3lL
UhRKnAuDHLJAyCMwbSZ6PAiL8qH3iwqhTw/L0wbiXi5rRSn6lxG4xdkrIW/wPFZqQl/iJ1PAZOUV
/i4eGhklmbBddtRNyZ7oO+Kn9YTIsl4JO3P2wBdiP5q+b5rnEfAHf6Y75d+lrhIspT0jBOhFB2ck
D8rWFfQVhsW27PvHgCSZSXssHX5gGE4K+g/mLpHpdEUmdN/r0ErI4KcahVe0W6RBATJO+9Ir60mv
XwBITe52v5FYarpwLkoTvrdot5CANqqxZoUaIS/zpAkadRQ/2UiE/FRmysvp9b6u+v3oqSVKhyHm
ywsEB47XmAMwSbBuisUtgo1GvQ8NgPX/rs21vdmD/qWEYDPNO09i1BglHh2jOkM629dJcOu8P98I
czNXn15E8E0KIChNXUebA0KsFfOGcsFKSLLP7jYr2n2zvPPekDYhMeQZ2VL4mrBDRmJegUrq/3G4
MSSH+8qmlq4fNHOgy+mvOeb+RFqh4kA6cdnMvs/8XE9nExPmCDKB5JNZ/WS/45Re/GBXFpjo6cpG
FnRsCJj3Rkb803NSS4IGV8LJcTYh2gwJ1cWaPtlHaFKkI1nBTI759pLvjYshHPZ9Xs1lWGXhfTRH
Wut0N+7INZJSmk9A0jXsz2FvkiVDyuprqvMNhrSMr2oLidpru1pgQRurGP98aHX7kCyKAu3cXuOD
gTxSKVnzscfuxtA41p5OpkGFLryAig7siZPNvOpgWk/Gp3bp5/rzLwRqECsopv4ERr/NvWFzTb8K
toXQB5RBe7GN2gnv5t26f7b/XSJXF2RNca6szgUn2/Rey8My2WkNX7XTPk3RLmrKoVCcw42BK7hP
6a5yZtCk9HBssOs4FjMOa5rAJQg495dB3V9BGsUPgbOz+IoUPeTSaWVoU5S1jhxT9F2OTisk8uiZ
OjfzeyVk/eBDg7bQqyoVHeRmWFWE/UztTbbBxmiqld+WJECJ+pbInxfpo3lpHoQ5huhHqg3X4wqn
E9FoWqeP2A0WAaNAcevV27LJd/It2xxX9PM7MK0OSgMOT2AJgQ283b9i8fvPhL+8BU52wDBrpE2K
1mfGMxi1HwbGqHeXqP7HPBmO8ZMr5GtV7kQ9nsqzHAStOO5Ke2sm3rHVfMf9wwRQsb7Fca6BZE6R
YC+D1AO3qvoWguSBNliFRjahGW6y38ldxr6Yb8y1aO2huGw8SYf4Lu7nm8pdKsktW0O2H76llWKB
Cqgiq5zT17nTkFBzgh8c+pMepqB+76SwnWZ+GFcd4KJZW9xfUzaRpeURfQA2IXWjj3WLOjjx9N0d
5ROSwfIvYI79dnUPTXb18bUECm/0LzzlWUVSq16+2BUL2O3bEEg6WXO1i2w37r/i8x6m/9G1xzUL
H+pwWP0YpYsj+oimYgicDPkCVPku/wssdV8LGveTceRLuC3w/b3xhp1EfMD4Sb8gjb4E+88WBcc9
0tCiBfbxz4AMsKX9yUefoGYfuQe+WqVrk5lrzxfHs/gkhq3s4rNyIYChwsnB+74a2gMcBmuovBIu
oPxxY09FARYfKWynJ1i3I4BmBq01+CSKlu9UM5Rr1uT0wqoouMfkIHXR1RZRxdOJJna8LlDlKXVq
l+fhWlbRMoOXTCK2LkOMUKiDphf3cl5FjpfGQom5LdArW6yO4uYChT0DfEgaDxUjlysqMw7Gz76D
9DH8CZnMsKYuRmah4czegOZ7OaI25Z3xCPXR+OYkFWCXIrZAk+Z4mwP4K+z2oATVKZJinItTR0Ft
rAVuiBW1A45SBbK0aOBLNKBHzPJ3wx847CKrdTIjITKL4C85c6EYjXJCgtX/O7WOEbhvNsOgrOSx
KQL+5oooakwLgjnQATgmsWterOWhdl8mDSZbFQR9Jg/SM3OmbUgfsXT7CYhqINh+1e50Aei8MN9B
c2XbTqU2lTPZjaFrsaYzC7wk32D9TG2i3mITdsPI9j4Zv/PaRSS8WoUyciXLzkjU477p+Phmmgjb
iHkxJtEcrZfLu+hLj0rPU5oaaqsgmL9dEM5D2dvZsbF2umpmBliu/2OHNxRXdz1bEDhsBDjc8M3J
hINeXr6LBmT6WkaPfTZqzRvZHUT0ycdilSfRTUxiBNnuyG8mmTjPHbUVrzqBu+zA9GJZssgWiyXn
XJzP1Fm6H2Cvu2envQ18IBw3ET3fkfn9ZW4ZeojjzcmcQX/Isj1zmWjPB6S9a7OyGcpVrRbOOryl
NqtUkYpHvfVdFFL+hM0nVis5tUou5Fj/VY588nPbCJ6gndiD/Mt10C9bNOYmT7YKtWqtVaP1s1F2
3ejIoAziAahFNZwHd22DCpgOIC1TPyDzSo567oMi4dec4lonMQXiLf5Oa3SZNBe3KTKsaQXqlbFo
uU67CXEfkdsCJprxcT5UB2vlx0z1OxVYeqkN0ohEpY2NDiPBMF69QuwtRKRtt+Q1AXBB8ItIDEPC
Q71gpOywfj4oOR20gTFohL+pk1cXTCGkspBID0X5vpacgbiHscQfpAFZSskDMyEmuidEb69fRYCf
2uCQci87VLpB4Vn7TaY27JqaNGT8M2iLtbbKx7P6IWCvWVBnv/s39lgMd+HW9sz+W26WXwrm/ZVs
K4W2DAIDRQB3PavMg5NNnjBc3P2k7JKllSlv3rbucR+dlFqtFOvUdH+hojD91O1WcN28/UFYSJwX
yLs1NRmnQoflpLawoixcePlTW2YcRSM1iqLQO2hUMkijYO4sOy4yOvPmEFFMq0bJ3ceHEp9D/8NQ
BQf5KqVZWlLOb1ww5hPe3zjoYQ8H7wv4+XscFuknQq2Oc3UXLpck6f/xxzdiD8a3P1IWs6AWZSGA
1fBHQ58s+cc5WOFq9rw8bluVvx5J1Oqsh5Fqto9Yb/WYAGKwA/ac4h9VSUTDEvfl1uM/LMmJ3Zbc
k36f3BDootJdiyuxwUcjwgamOwy/Z6CbAAgm3tl8cu2ylzTibZkQerRmJYgjLoXrXINZTa9mDQ0g
aViYMksVLt7O9zqpLL4PafErIYI8ak5juVUT5iYq8coEBNTh+wtzysxNsovZT3czYisVO3g/Ldqx
Cd+6TQE0zWKsMe9jw58iRmUvmcQAAitWJuartCohlbA1hqE03D1RoLG7/4u8GEKJ/wSMmBWr61rX
uswKI097tgD7KfgYHt3wmjulg5Q6Qw8DJ2+qqtjb2H4bZdYPGqa++zcsk1Cdx+sgdzMc09OXsAOq
UJ8OTve5t+1RgVL2DGsy8pZarhpEO7Hg/V7/VMlUzCaGHAjmyksV2AYZggJJZ2nNIQU6hX/CEpcK
z9ESo6HT06z/xg4pWRpnDmyGsiRtasS5pePORjrJ5ytd/xbi593fwzEESLth77hvHpxKji8wADKU
C8EVcWEmMSixrSelp2MIGX2M6+e4nk0P7tCFITB4wdrCUd5d52pNov9PHkph35I5cMpftLwgD6nd
cB/4zcBAwnVCu2+Jetm5zcJuGinXY11R7akyeJNIiRmQmD4U2Dy0exCLdvri5SwtVzkd4wP6Yluc
k3iByaGleQaEaoy4fwGualY+vdd/2Ch4GqsrL9WiedCOr5nbXpZjlESNqIi4edSepgGhFfzSVVao
oNJ2jIbFgMeGk0btzzyviXY/4kPapebnFdJ0uFutHITXj/rqTz4LXZQkUQxqsoiuIa07KZdlcKfr
Hn39YbulidZuxZgiYEQKuleQPZlOghoe8qqL0suQ5/TwM+9U/NnCukLcbYkpSxpP/n5+rYg6yZ8d
Aw932PS/H8a86pgMWOutAy6DEwFbo18eYfZIU3lo2onRn8Pp3xeQT7Da13V1UOut/vEL7O3q27ef
ByNYSv1hdGpEhI4Jbq2bN5+Dwa6TPKV/y0MxmJJJp87P+cmVc/lG0pFc6uodyJwJEDTZqPPHw6Zr
5txoj44IA1FzMRlewUNJ9qMN59q22BTO8Eo+V3IV0bG8hALvrhu3jITJYZqTJllRYkCYzrjc+jnm
AivT+OjW/5emvCJ5mohlLq47S9lqs+AzkSuGI4vTMWo2Es4MR/WQueIC3Spjf+HBoPvUj6WOu5OL
DDgy3hWB3gSSZBaJL7FTpu26PXd+aThYDWY75FMIjzXl9HJZSn8kDKJH/KhKAmHdtBSqcdRKX9f8
KmzldTYRlrMoODKSVXGP/Q8NLFHWvg/zurNf8vB18dHFNkJufxLvfERhkVpuXDXysmW/FiTc65Bn
5hE/AvQ6eLRNE0qv/smUF8Ic/swy9dCXNTPoM7Ikw2zGjuM9XoY9JQBw+SIS/QjLBYZvpK5H2YYO
WdUvNjkFS3C7g+EQfTdWC7USkIOp8Z4krxZ/vgdYvDVu7BR9ie9OQPmSjPkGL9XyfGHPCbUvVzYm
wJyOhnF56sI21Uu6r2TWcu55tw6YDAH3EEUIbUN8xqTHwLkBORFubv592OvXq9VzGLfPC315eaxx
HEACx3qn936FvxrKWq48errbXwY5vmGeLE3zosdrlPvh2iL0FpZxGzJbJ50S3Jv7x811S6HwJr7L
OpZUH4tUao8Vn6H09KF1qPkAZkj3oKCfEtEeVWkwY162mPZMrXoFX6wZGBaR2Vc9ibrkacamvxlH
gI11sUa2g6f+Hu6No3ymPHK6vI6myoHfQaMSsWuy2aYIHQFpejZACq+QCDhFD54Kn6kUtnqHu8El
wkgazeXN2nsCi/6hTNw9Ly+I4aKKM9NQZJ0W8gGCheRWqSpneG8sApfjFyA+ve2irGAUGI9nR0qB
yioUFQVMTJjPOWdJu7SAzLPDO5ftbocEe2VhTSB+MF6SYh+W1eJI5/sRjkFrBMRGP6GO+y944dYV
Rc3u+0TYEhwc041WMabQZkN4KPI9qCkc2aMX47PfqkMR293RKZnKmruqtFd6c6XSbIEH1s9oCnQ9
zQNS3OXdqltPkhtByV8wOzALzNz0O7Bkin+VzKv/fZDGvjDtGVmMmb2xgIUVA/nnXI+z+KRmH7H0
uH8Fd+wKDVsjBx+HjFMOHiCieV+tazFmlgKnWRbN5vwNf9yt70u34vAg1+ZudBID0QAjw4EuJnag
9JgOWmZuDh3pLfJLcoJgKJK5mhtSii3Vh2iNcKiuDzym0aWribKvkIKZ2PxTMBig6TjOZ+Blo1zG
CLlhmzmW5hFtslm6z05Yk2lPr/5LyNhElNcPV6JEYmc9hpHVq5vnQmu0G/eHGmdCBOB6i9RBTZLF
VQO6y30po8H1TN1x6mIok3UVlJi90PXEfKH8rpvHMNJDZeXw61EV3NA3xAOTaFkjO8rbrSUCwM5X
rS0M3aEOs/iWOs936tZIYfwKAmLSzviRmi94cm92KUwjtvGI1L8n99lNYaZp/wvNaHdkRgaiCIro
eZNGelq27HXSnJ1kJPpX8W3kVg4pflGHW/2ywaa1aB/59AJfn8o9i1Jq6gRXPfEuuVuR5K75sYhL
DObpHJV95TCGjU4cxJi0kfaEw/2/yMDYTKOStxqtmKe7Molrp0EJsMJlOFT+hwM5mj3gV2fRAghP
74x41kD0H5wVjznjIJBeKtjtKbBUFg7/xugVrCxAdRNQ+OafFVsCl4HpN9/As6Pk7PDG2o1Ig3LT
zf6aar+Tl29NVm3wtXKD7KuLc5pM+AGZIxXRKe1FE5ATGBV+vI8BrDPwC6Ne4P0ACOzJYJVqUlL7
axJzW0DRqcQKQfd8ulDs4nRiVxNCe5wgOrowWi87Jl82QN0yuJqK4XYeKQFoms85s6N2n0V5XN9Z
/NKHcuRuJzAJl9lUgTx1vno9asXXHP/B1RxM4VnpGNaIhsfVmFCH8yhMa1DUx/Yt5qrZRafT1tEV
fla910Cw2M8gBIuVSHi4etMdF86s5f96qhkfqnh5pjr9cUsWjLWaXUAHZH13nbCQ8YmlWvMUnOEM
axkQMaOgdN+9QryHmvyEsdJfZJsHU4uifJFfChXpSQhud1W7AnAjt45FkiAxDUiUoHHC6hyi/Tdy
kSQ7wBDqZhmy8Mhpj7T5t9aLWFXSOBszoibVJO6prpjFSVyFCwutCkuOD8xZNutkscBPd9m2ZMfl
OPo4I5fK/hZzJ/vlNDGqXnGU/drIZNu06nUdABVKv4h0eLJzxQPc8cNGQdIBUrobCt1OoML/wwa7
+C1aQq3mV291xg6dwFaz2gYBE5P1vH79ln56e1IBcIj2j37eWwaSgohVMhp2+ySGFBahd2YKJtfs
ypb6BghFGz6drGLvx/6zFszSHOxO0qr6bGTzQqO07PTvWeDQyflt1urGedRBboWRmWNLIlCz1uBS
PCVMwLSLKHEj4wY++JWugfyIhg3qjQ5RxrzxceR9n/6smU4FTRKUKsYoNe+m4EQ/qhtsNmI3pBVp
EJZ5DhZUho+0TsdmnkFRsbRnQdB/6cNUmAVpz+NUwXCoHiEpv2m7imwf75F3JuOF1dyaQypAGF73
YySd8HYRjMGaHaoWQg9TWc6eJBSHbi2ZrmQGjl9ZUj149zA+Pd0NJ9oMv6pzz5WaIU8LyMJlM8bb
EDyYjErrPH/09R1Bb8ddNSIUAiLEBo+ciIgxRZ+pQ1Pky+NFo7VYa6el195Vw7CX++NwL0vVnkj5
eRlcEGlN5dpRiJvMu2DxGK8Qd05S9UTXznSILIoDpHUs0PPdnAEJTOKLJxSOoKNlcln2MeJI5wDa
IaRNjMBeFUAk0PzfxADTdh9fTQBS4h28U9hgPj9SVj5Jyroc6tHyYB9Ncd0qJM53+SP2ZZ06R4lV
IKfgz2R12E6+duffDH3PyDl+GOLhFUlpm160rSkFmXf4pCMypImsWTFobJc+Uzaqnsp9LTQtSBIR
bmtfBMIvrSRY5XkPEQdl5RyEQwSk3ClR1iVwbXIra8Ht1pjDkc4KJZRrr7d1pMvL+csQ6N2jsHEb
x1r+hI+jr4PMYB5LidcqsbjHZU3TtaODZQrBSiTNKDGn1Ri4WE60FOMfW4wYX+3dkS623nPCXJad
4Z4FKAYR8MnMV8017HWKGhW8rrr/wUoeyzV2M4EmkqHKZXbA31c2KbzDpMbQAzzVmkJEsa72z+8a
Lenx2pVDMHqIWETTAqbWqkmjoSF1yL40AoKg8GUF8fV3ked2Adg4kBt4TNdKCw+Al7/ySPETvkfq
BZfUCdBh8CY7j1lkx9xftvyCnvRID8HC7gxL1/+Y12uDXCFc+ZxWOQh6FY+XFal2foZcNtfmn/T7
qrp5Vj2BfDI/REz0Zha46t0IFbow1B3n5+rAC/LveofRUvwUaU4Nne0kakjrJPfYJDA12lq/N7mf
id/u5fo5JygT+xNGcwaLPvDAKZdFRHBfjhRRa/LzBkTmSy5pQ2LjVzUjbEB8PLaFWEWQQ+kGWOyI
6rD8YcajNccpYv4SkARfWifKInKw1uSW0e3KuVVy1SM25W5xAzubDE2FO3cYmchCy2T96OEEzZJk
4/CHnF87mJ1JWGKS0iKl55jw67Y7xt719tDcD9orkhYXBnNdam/NYQQLxNktWHNkGaL+Sz4TuAa/
0SuS2yLfDDT0xryBOFSGLwz0es0iIenkpJPm8uNHFTFayqWG/JfshiqthiATiFB9zBcCCNvCFJXw
W0JHuc80lHqcUX3wlKwhQgj9SqIZNhtw6QekPDMfDeXixBf83Gzry+EU2TqwZk8pzY24/UA3WmCm
yMG2GvACAun1dvycGDb/cc6VwZbyuvr021GBembXrcBLbZpvbqxgO9MxwSAHdu2yL1KvsVYEedx/
FYB3u3ZBIUl3M1iUdl72IwIVpZ3EP7ESOlbG+e5nkzH3tYOOeAmDdDc1JXjFCnlZVb51hol389fd
q7sa8AehkEIrc/JsBsKj/XlJ7+XPxXFPEF9sKWhBPRlN/yQtzAZQ3BVSGqv5E2khZk2sVqU1x33U
sfpS7RrsZAKw3bIOAnN0qTR2xrsbrdfmQXEVqBXw8t5/60l4URg5HicS9/aXP5P9Ng2i+1VBS025
YEdEYRMaK4BPtU2se/+zqGUWuj8fLY4cSW+CHnkzuLHCOYB0HenkdOZQJ2jB8OCcjVgbYrEXynFY
ql/adBo3lDqHRc4bYvOu97y2d9XWIQBq7u9UGRFHo6kPDpZPY+dTHQv+0Mei/0wbT4sXCHLlPyuy
aepKi10+EKoAv3v3lvQEEYGmrq90r+vpTA8KF/3gXFYHL8Mvfi6vqSSgD7N0k8tx8D6tO+giP9nB
0Rsy3T5xNbrfCBIS/8/+ajgOgwmkze1B/zAPbLb/Mj6DKVZQi3h0Si2xyqDYGL/vi6MawGlj7IoT
xQIYpJQnSHJ0LCA2q87m7lN9iatf6wbGrq+rZGNARZQhZULzm2fZMCoBVxJIQdbsOOSkAoDV1vvf
EyDSOr3a4oIzMYOpO9QzfkZUSeSxbT6HJAAzghCbiZeFcxsghF6GgT/HL/jvspvnFSWMBF2L/bbw
StNEEr4U2j+IXXLkG8IojBdVybf6hLPS0kkiNAgN7rOFmPjIBr+ezyB8fdX6NeK10nqInrjYiMov
otpzSOuPUv5u1Gj83z9aniJFY8lgahoW59UpKn1LNsNBoI8fHvaj9LF5+dvMFF7vUJcwMeSG4dPN
IUxhxQziJCNHn01sfGUYuIaR1AehwsQ45W+sd0DxILRTaqF9mN0AAuQ23waSZzPCpsjjgS88I6Tz
9HvRuzzd12qRygs3RXxWTSqC5u1f0Qu/OYI/9GUZl9rKAOr241NJn4+IgvOha0A9ixZ2R5WMDeaz
CeSQgs3Sf7BBAfpIu57pVPTuNPFFSh/mipTiT8Ggva3cnb4Ze3dri24FGt9y1zXkxEVZWVKnXsgL
oPVToo5k0o8iQEag0Y7lz9PesCasyYMYcICd5BYDb7/io0ucgTL6wwlS5HWRO2VctoxrX4rtPdgB
BT6zs8n0sz+Vj18UQ79LKdfzwSou2skp5RGwfKJpTvYuaWpQzdBlHDjaUQLx0s86Njnf2Q8w7QDU
kU7aGsg2g55NoJfoOKGz7dE6oWHqU5EV7eEZXFcolenb1nQ0LoWYeyc9rvRMcNxLFkbOrxChWwTV
qj2XKb+M+2xeRl8UjYSWvXTZmeR2Fs8Umwa8NRDA5Ljmt9wRw88/JxB0MSqYDKOGCX342PddjXHO
6E0UOQD3P+wrwP+fY4Wr4apibIoxJVWZC4xactrSyS5g6DZzreb7I7zRzxN1mqY7RvNBY7kDsjJi
iNdVuEgBixuC4M4+CNTD/qvf8i78B8yhcOQOSJb9q+4/QhUByQDNwMo3S6FlEUOaTZIKEaKeFAD0
61iSv9r8xJEjWKH91jPJTxIzkF1333So/+srwczNICRaHxUZjK9LBOCbkgysibSgirLRHLx8Wxn6
QCYDVNmybx6gwKypy3FzzqXGziqJZE18p1Yeg7lcvnzhyYjq+AEVwZWQAmZLx0GTr4tTROGQy2NN
V/LbQofuux80+/hDAhSpnD5qBDZcTHIbbI/gdHNnyxkB7qNRikW2u1FwREFocsMmnQdjtllNLSBD
c0iRp8tD8MhF7GxscD37PiMgCdDeZOJ/M7tjZRaMbFmODC4m1hskLU/kPSmcM4+abOq2ky0j4t/0
T5V0gum7ef/vwYYQv1cCO75JpZGzMaglNKEaDFj0Jf02fkYAjbY/qco3YNQb3WcG2WPLJG5u6ByO
kRxWAjRa0JB+1lPlPGZD/bb1SMu1IzL8SWyzJ45PIU1HZmHVhscciV2X5Ms+Cj9soBGh1nEOL4mK
SOu/PJMR3JiQyHzi45Mk48VqWO4RPQHMXq3jqE2/kxQwttEYwSimdO4ZqjHGRwH5shUzoKQGCj5G
1rCBWxa/MLa/Njk0sqyTYCe09P4qMSOCvC2GLFxQrbvUIprCvikDGXp1uAQGfeweHVh2DjsYp4nV
PUmCVmw9AOmAI0vNcThvRH5Ydwid5LIeM6BesokjfspuimPH5/3YMae4x9+Jlz3ppSzU0aPjdaHH
FSJb6ROrgxkvo05UEXWUZbUUVvidP8MBMcrM4UvwvHBjjr/AxZ1FuucmSYO+Jh33NdrVlBFlxABA
zrkuje4vkQCeQssRNnkNiY4Ma9AUm0lLEuVo5IHYEgfxqPqOECJBy2/PiOW1x0SmciDzO5AKtQrp
zeAekkyHmPOPq7L24kJpZy+6levZgoW8Kdafuhyv93OicjR/2W1WtHoAsSMTLVqZX+eNBkdQEPfu
EEHoxE0kqxkYkxcKEtYFUjA2I5eJp+INg1P8otBohYSwDl2UkR7gUkGZkdMoq4kEQopfxdM/GMiT
a6XSixVVmRSABILa8/tp7YcYP5S9Rge0+AUU1zcnSfuOxDVmeCpwgaI/xtloCyIhzYF5xMHdoDEf
q5snA8vQcTk1aM2Cr7jyzddA9Cg5+53l3ODSalqNFeoxvXOXP9XR2czIUuhjh/T6ixcUbfx/Tbe1
EttKxsLOlHNEwHJG4rftE2kXi4ZGY/yjy7WN+Mg7Ot/4p/CDLFXGoispXvcqyyGylIulJX+EIA+I
FyEWEamMQ/9p48Nh5VoWQFst2rV6748ILSvcXmPSPgFdES38tnuZiP49bzOSZA8NLLiRCTLQK9Mt
eC8FjcapYtekHc3ufqw8DZPnjGu3slu4MI1l1TqkYu4blHtjBLaRlkNe97gp/8oEbPMRqvbyeuq7
/r5s0LubJ5DPordz4myrQ9Ka+krCQvxfOGdrl8zvLbNo+HSB8YF/Y7F6CKtpPYBt85iV9xHV6fk8
g1PkMoCxP+aKHcff9JKsWG5z6fSFpS0PXIQeih+x8CJtPuSGkTF0RfLY//opAds/2SyXjZUVoB4y
6XWBDY29yAUtBMf9nPi926YcwlcoOqoQ1WKPe/5G0P82ONfcaHdSQNTqRhH81H5J2IUDtGXacQHc
OIpciY+3vcgPa3pU99kE5hFYur1ItuC6T9b72VR2ItA1MbqF1624rGNH9cYU2Domqzv2ysw8h4YR
tjEjHc0YxS8kPJe/CJ8gims0LyqOXo9zDmTk2WmNWAftGYtyIGfjhDPtWXl06dGeuWw+Cfom1o5R
zkC4VV+n74i9RUx8C8JHTXb1O0giFIUWrP39HCe0SHXXdAzfdqyWNcRegaMpdbVQxAlqXGOHHwFJ
lDPk/51I3y0m6Lol+zhPeyIbSDAcZyxiv7Z+VWrDslb2nPyOeFeYA0SmpSZdZ3jHr92FKtkYGlus
s1j9oQhjiHeZTuQWYUiFKMvFWdC/WOHaSvRNiVcPt0wsz+0g8fOwmrKrnRhYe2isOOF0ekgBT6Ts
TeYv8lA9EYxZU9bm9y0GAP0k5u1FJvIMIq1VEZ3uzFvhvDu6jvlQ4yt/jHv3I8a7qA/V8Te8UDX6
biO+Lq1ioCqifa6i/OHqsfHZ+XrhCsb6NF6zjmBmD45Up8yiP04KvRr2Z6KHt0RGi89SLoArkEtv
sJ/Fu1YY0MpWxDQeTHtAXbWJV/dYTCwPpdfHAQ6sUcM0RaKjPFTJAa16IYFuhMLnIA0v5hB9J1Kl
sl/veienDku1WLp2M+uOeSh80mh8FUJPt2joULMGf1+Pht8ShEoNOMnV/yvDagtghx/Y2wDpJe/H
cSKPnsOv5piJuAiI7h29yJyW52gMLIYFWWJ9OSIwJpA9w7BJfcvYp4ezEwe7xdL1uGBcPJRq9A6H
efWcgfKnFDB09rbwW2/mT+1WHuJ9NQnI/PeqmuKQlXhaXGINoki1KpQv40mBHkO1z9YHg6Jd+6yT
0VX4TXxAQh3uN+RKKOaDM56RIHaMJeJxeoQI6eV/oYbZxI/RGTowhkwHSOc7r3/7UiZTFxucdzZf
uFFbEPcyBbH6Xpuu3sOJ0E4drujTHh5NLFAefrQVqdPQ4FtGMd6g1jZdvI7b0KSIQa6Lea6Vzokq
pFQPlVzMqrg2snBjKo4PinIgEznAsMksP7WvNm8bbkfvVfEPtM1coBBUceZ7YkH9ZV5MYb5SfhxH
/B+s53djsIhmz4UEJa7TLTGYe4x6FMGWeKe0YRzPW7ZNjFZRlGEHAwqxkKTxXHj3mVrayueD6Tkm
wBLMTgNXcBamFhy1RxE6sjOrcM2kne6pSCadwCJYSW7TREYt6e+G1lamZBbtTJE+GH7cxmZCku6Y
t+G8SmiD4uE0lP/8iVrIZbOX+tAkoKAeH85Z48o7g2HqDoJnETyEC+P0QXzBGoQ6S8oOISarHzDK
An1DD+HdkVqOCyL9Pcd4ZeOdW+p6KjXKyhxdj42oAYHLgE5yLoKXdm07Ljtn1J6r75hKSIsL0qGS
GQ+BuSyPnYVWFP8oD9dtwWhM6CnQ+H/x3zAe59QQSj8DeN5K+SLpmyzSeaTbHUaC7gA84iBknZBh
3LFe/liX0Gg+uTUBiPX3ruRyMalkgbrWGgIDHOj5wepOqK8eGpn3DGiQDDYgX+nbLrh1dTivS/1x
QajkEBrQ2tW2kj6jyaVFAFhKODi2IvooWJemHa17/8PceqlEV/SW/3qXw2VbpUhabta4IAHAjkr3
Yk1uhMJFTrYOBZPbPBotn1zqxyHoZiSy5q6neSG+OiisCLVMEhJ7MfVSDWzkGtPgJcc2mOBJ9hIQ
eakkww2ZR/3FakcEU7z2C8DLxNpr3/H7XUYAVAn+1QP858BLTTY9YxNpGtqmnyyOc+56xWknarvY
Z+2b39sL7U2IdSdxQrTC9fnGvPdYs1tp9s/tqcqdW8BiQ6xpv9Rqt+GSglLbmFBfFHLfiSC6BQ4a
vAdSBY4/PmJCIkPEqg9ECeEVOdr1JyEDrQon6Ium7b0oPtbLs1fCq4jQ2wsd9ZIDm5Xo5QVA4VAF
Tkj4SZCSvrGqm0NNOavc+QSYxg0kA11d2IWsXtlU8k3zyWlIAhCdYrykehI109vDrb0l/3vnMNDv
VYTrS7e3/4SPaAhkgstJhwVzWVwWUwvTjs81sM2a/ywUw1iPNryjBb2o1gCuU6h2kTR+vaXJDvxP
34r+9qKDyagVVGtBfZwXfiHKKNYBfsIYcvjrVCxAqHi9/8sHUYYc61EuodBztzANU0fTtuEQ5iTY
mbkYM/qMd/p+BoeiA7EmGLv0EJzq0bO4R5i2aWmPZ173fwhNyARDKcx08L3DuG2GcLMuKTPG70cv
p0f2jVVeYTFS+lNpYRk+ER8ScTDz3xBG/iuK6AjPEm2Y94Lq2tlEFN/zJwmIAo3DndeG4iLlHGqX
ftHeLKEIOGWD+2JfYmHottuKNpQdyzvV8W9gt/LbW+5xBxeLMAqE7/Zf2r46FLuj6VXUQ5C/yC1r
d4YxiO/dKkk58mdGdeUzWyD70tydDV66XZ1nE9NW+yRys0F7EbCmbQSCo7VkX8R3+jQ5zz5iR1z8
ucgHnNMS1TppcgN0nTYXSnubNa5RHMuOxoXmapWE9wRZZJBaQKuYN3mnhey/9VtKUtilYLct9jXu
xcpjTLyOp1vUOscFW1/1Ve6J5j+rCTzWQ+HsTtE+br/22FKjabWvD0qfsszTWzh7NXSQoiEBRxbl
dtrp8kF90gO3T6tNAazw/gg9cCPcyAQSs5OOhz+7q7JVKI7nx8j0Oh5WzFdrScktyZdqX//sUVS/
i4jMSYcM0hkMZFbVKlSf1xTB76oCeJZic0iJun5ByzUK8EYtDENAre8hmMVfZnMe7bVXV7SgSf8Y
5jJKZfJlbHUmEQU2eHn0X8ualqzt785PPTUk8UYtx+2sHCUwTSDXKv6UUdEjlMcYXDNXZ/jJbuJk
WU4KkYfkoNKp3+MRLKnB7onixs6lwwbgiumoeJmcU+rlUwmmb3AbuPrKjZqIeWe9Y2OSJFXKiutI
Scvp11Vc1FR2YqR0E5qH8jcLme1/4wwmI6/s2Ax8b56c5k6OiMYp6mQlTOw0py+LoJhf1Dz0Zour
ecuAqpw+Mi/qQGTcY9J2OPzAEsWd4ywFMV9+Y3IoAqudB09XNKmLOhb/SNr27qKRj4zgltflhjVc
wTZM+1me/mccfDITB0Oc3E6c/MAMRu8vAvnLaMGe86Q9EMPdAxI+6rgZjv52wLNsMvvokuBTMBfH
kNrMN4UWQs4ynYiYBnsivKLXKrClA91r+/mP/4LJuNEENRTa6R7bQ5xzxnEvhtAYB2Q4QH9LnEOT
OVG3PSBTdS6HDFDOoAxklJiMJoxL17xkYnGYJkY+ZoK18TEeo2rXZpayFofpFOJpvxzu/wkmME6X
h8OlLLtVJBWUC8+WjYBL8uFBG33G3dL+FJLkwKYp5PgSGccocRT/+D68m6eEdmC7rNgjqR9CkP+S
pV2vSlHzTXKkir2C6hPs4HhsTX4de9nrjRZGkMoMwgi5CqoDa1rfsvhgume0TFpFSIvWrJT52zBr
1OGnYTjHdzJjkfrheVWA3sK6ecw+jcdRyFiViUx4IUQeJJbEGn//HpnaQXJNwwmrWscZxiMsdNw3
lKo050LhELzHSG1hIPFPIdJZgxQ8YfiP7AbN69rJFZah96XD2sz5gG5GEraONCfqhJXnY0ErOLLw
ojwz7/uywmYxgwxLXDmTq/xcezJCfV59eVU8T97rm5Darb+/O5ccKWhtxtFvifxn5uhS3Qke10Pe
euBn2DqWXXECB4i30xl6BMzj/Bsu27f5wM+iYFPF3/yNjJuKIZsZP0ffxHr6DHgFXD9CSfM0oOE3
c5lbWcH2UT2JWxlsoN7PEWukH2HQ0W1Em6F1lTtMCAS3eyJeIGpPDylS+eU8MyZL5ZzAcR3UuU0+
NUp8/A+ZGANouZVcYGG9DKjeKITjJTw/5zIJZVDFk++a+dVRqSRvr/hccoXoaAzJUb8Nk8gXOega
DyPpLouUu+BLlU4xA8hapeV4fL36bobXS4a7h9ocr7e+Yye4o/EWH4+7V0VxzvWHHhkD0Yo0Ykod
JztLwfZRf+4GdeyRqdu6CFgO4v0nMw7JyBg+94Mii7eTQz404AYetTa6SeAQkUIq+DG+ZEWQtu70
xbgKscPz1Txk5SB8u1XLsYMRfKTTWSTQqYrchlAcXEMJ1fqadeUyCyLHzYvhc4BpGk5NNia+z42C
RuL47cQiKpew26wMR6XHICmfKL3f7UuVq5yAhpUaiDWBgcQOAYp4bHUCxz0AWev/+hk84OIckLZ0
k0OtChYK8gHlsusuwrCM2ARa2WmF+USZtUb7oLSeC/uflBEU6EwZzBP4Kez1bLSEygI5xJSFowlM
vM3kZH+YMMkZzwpIQ8macMh3+xGFn2WF996Ea9DcPgndGe8Hd00nI4UFik7zH2aHyltxnQTHWIjx
9hbWJD9WgkqMY+0jcmMEIe79c8a+cdxnT3wCt/frmaSFcOHqBx3cx+yHvK5f9fl2a3Ln3hHgRrTH
qrvkp8jqbdJyKoo2BGFBvVmuNwWlJl5ek8wzZNu3NdDQ3MHdzL1oCaOCEydZr1TeazgvWY0Pn2bN
0Z60pSEmw6on/etoh8B1E7epQLoPaKviHWCR03ez1v4wT3GnvZ5TzC7D68HvXzUmYWduAhoPC4zu
A1JLZ9vmoLppIWpbgxob8kesbL9uFb3vOf8oItIt1JzbpUeJ1mH/el8DuA6bbGuPDRVyG6mThal3
tjJ+IAFm1Xk9bO2JiVyzM+wrXuPIvJ7mWZzdD1vm+MGgh5vvpc5N0xXAjizdKQ4w+SOwSPmvhZSl
Vcb30iykTT0sevDiYZBlwzQdVq0k4/LwXkdHLbCr+vicqbmUtTM1iCYzUuEEQT/P62aNo31s1GTu
FejSQkwYOQdvXCnCeT2St1KdajPAilwx/jFUEGr7Fm3SY6zOHIid8/GG0YgQjXa9yznZpqmcABdR
IyhB2834ZSCtt54SQXooOjhoDJgKH3/wGD0k9iFCCfJqQPInaMIRUX6kl639a3fHp5YnSXCxbwUh
iBMTl+NH4lUv+/io9fkyqlscdohm5U7bZCudcM+lVBrE5JvMQQd0GjyFeQmBRhGWhcu659czJLsJ
52nTRF+X66X5lKrgqauUyDP4cGXELTz3D5JGNQf6+NJI6h+BMQefPwLrOAUOGikVnyDCVpnGycJk
u7WE4b2HHaoQza2nXaC+0DYNtqrAIR+tc5q6ZA+8+y+Q16myv62B3iNCqGmECo85COoHgu4vOBGJ
C4j+6meIgS+MgJ9jxhxv9n3vHnYJmngp9FTJAeBlfUXUfnrIZ3EOwZIIpkebE2ZlC4qajR2H4tz0
HyOSxIHVLcX719sv6ZDfBe1OkMCEL04RO46XsTevMOF4btbwUGCkj3mc2WeVohJ2cg+v0lsFLe3N
1LzyrOX9VmXCRU4ZiOZ3jDHs87ImYwQYpWyQNH3Wn00JB/oVsl24U+cT4lovHG+UKYdtyb1NMeoN
cXi9aj3Nt4clalBx/w6aqqn6j5T1nyNWas+mhsNEXQgW/9JwSZzJRaRmmmI64biDbqnhNFdPUHg4
r4xF4ReVq+vfCN1NZEmkbP7A/lm9Q11SVDkoufWPFzTLdUwLbwVeCPEXojUuMCJ7gvGG5hGHjV4C
JflKt7Uaugjaks4W0hBPYxxfLszUnhk4+BFYXTzPcqq2y4nfwDm0Ezl6QJMfUnHUUZBwj8Ere4V/
vLVPZ7vmF4lmUo1nt2hOjIs+kQH/s/mx8NnsKxUQqdtvrfUQpVfX7dUICuc5jTsB4rS0p6SHpnmF
lTcoK5MWlJ5Xpii4c8H0g65CUp2Ho+lf+8EHg9Aa2jm+U9bP5elnh5Lav/MqALnySN3N95N02nsu
cVcnQia07xVWFzwQZc+aLZog2wU8f+fGHdR98ouQwMoO75xAXCTCXnHL+WyJ72p68AwWiulZXshy
QIeZ1IBL94rCKb0ZoJNsZY9m3u8/T/4pwbDju7WXLJ9W8IHXiTWtqx6RWSaYa8rrm7Xy5NYpIDBo
QZbh0wVJQZmdDGHbL2vxRznC4SmWyc8nUCa5zV+tTqPluj0+vOilgmyV+byTuKbzWr2aKSmuIHFl
Yb4QQTxbO+P8EXlersbcKjWaEqTCI0LYhK0GjVN32HOnZsZ5pB5j9h4BW7lGQ4RJlQpPP4V2FkwF
1ZxJsYJ1YS7fq98Ej4Tq51gD+2vADa48i71eG/vrSp3OKM4jPANACBAgKnxGoDR18A4dUpYEmoML
sSF/gzk94fePj4vxY7FQ5GPZuRXCcm33CG4cKZLG8Hm8CutB3lyQinPL1FJ8Hd4+/CVNJlGN6N7j
RofJBVAEc60XsKpJzvfSlSEf+S0KmKtmTRLs5FRXkrR1HKZ5ufMHZn5FupW3413z4hu+yKyHh4gG
VALcGEQHo70Fuzi6OSFtGa7lSC47RcaHJxD0GTjz+DcRLfXU/UplxrlcExNqAIov9TLVrjHCREP5
s05MVyI42SzY0PnVkv/tXFPa3QpGMPviRGznKfNvgp9B5EVSj2Esvr62uNklv7N8+Al7lTvRW6Gu
CzsjhljHBzHL28zgpbS0Dis+JohENlJ48iC3Z0voQ3RcfsYbv2hZ/bgGwnQ8qBwNQAcIhhqkV1ez
K9+/9lhCCrkBUkRZXeQ4QNKMyZt0M7HVoAdLpvguF4hwTdkp77701Uu8Q8CQEHLHXmuZ0pAkTTfS
QWnGOFCcx9VHRSh6IuiT47i9ghzosSBE6x2eOYSs9Mdr4mXHRdMWFOnMadps5sn6eu1+o5uPix3J
I/5Pj/9UASG/iqtIpVCL/QaCl5wVwzEMLZTXZkAsjADy2QVZ3/fdWamyJl7TYbyWGBd/ygeC+utr
VWkJgoGlb/eIFXXbip3QciQusrG0H/dU35NvUX63jMLLQku+TdTkY1PMZNrbq9Q9RyC9gqwAJnK2
V0zhChXiye3JuuEvHV4d4T9tWtJSkNg8xjfHoe8AD1BlPswXD8/qKAHdZvzDGm6J9QZYN+eCv8jN
Kjx1buO73nztQMiRRbyECcG7by5/WkqurRSAbB/mMAp5JBHH5Ge91ohiVg3ePd/vMtgGqXVIRapU
mgaAijRYJySZLBw3uuMvCyiyhgRKc9RdumGOOL401FWm7i1aI10nfRUWLqI5jt5yEPTD+j/pizDk
NmEKj64ZSEPCZSlAEb5zTPmJPaE2Vi2RL3u3TZEBwgsgcwpbtLiKLgZtCCSB9pyHUa7tdiu2iLgn
wLA6TN+3renQuSwGJYWJhoaaAu/KxdJpA2A6mTspCFSur9towCnKgSWXwh+MopGJCn+3gn3K6a92
jK68/d4HyxdBgGeCEzqFCId2fT4cchwRzQlngxoupznCVRqV8xpj0cC7H7RUBxJnOORRgfmEmO8j
GMSKyn33qQ7umrNUlUPOytCdTQkfiW12o+Hd5iZSOZcs98ka1bn4A1w9OHdM5epaXmezSDfFYuNI
Liz7UydA128EhfWFWzD+LKrasb8dd+jqeHx0vXqeMOI72I5N8Frc24CvoOWD8KJV6KcgFEve15me
kwnQcMxScBaG4PenMMzxXlIQoWQPVw/YLpvsRdeEhbXJLgmdkqatYPM8/+qcLCcquiY7lR0aFyq/
Kdae98xnmWhEYp5m8E9NP+SXyOJkdtxHzxR0kIq31mT+I/Kt7RGO/QAhkD1gcRNZbMFgKfYqT7wo
gCANUQNEsnKQqpoM9snUhneMaAsrNZgCXmOGYjtEHNUcmJ6zYICcWkDsWgcofAn+yfgEq2Iz+81y
MP29Xf3Ie4T3z+OU1oa5n67CSr0y6SEjzriMB6r4X1fFHD4dquRC4hXRH2fmZw4TncUo0TvwKNAJ
sQXrBwQcvsUem5Dlm/OyDXmyHExZpgcKkB01DK4UERcsxwztg2erDT5P7eUgz5ZyeyTmms6SYRDg
xXqb5txmhW4Jkz10wkxVYxfzCMBDwfaGOcq8xheNRuKS/hCMpjCca74R1uqHEf3OnW8XXttlZ3hW
UL9Q70CYnTXnXhZ+jjcRy5z+YwL/IXZaoAIvIJGZF6D9Ed47PZF16Ev7/AZICNCA9sKPsb9HzC1N
OqljSNPK2NwTPFwHsB+vB4sQhO4R0o7S5PqLiOGpl+KaAbfGhnxVOtA0Jk5m8l14nwHXSqwMq6fl
9isxSOKhKmnNViAeoMdw01b0NjaMMdHwpOV2j5PKw44YlXC/VKqcqmVj1qsCbWVPJGrm3+EVTOxK
oIl13fWL0qXDrdS1+X18rQUBZFK852x/iRcby7csMq2nv1y0T8cxmdmOG1eGExNBTPL4/7hkO+Aw
WxbEA0SKgOg7X23upJE9Y+FslUW/ysIedkBts+9cX98BSMavssx9+KQXq5nsPfrtGi0R8BPZJPDY
JnpbKIuAHus4ObSPSxn7KNtTC+nXJpkM3/PzxcCyWyLs87Z2ftqmtSXpO3zeWyX+TLuQ6e9ofk4O
AdaYqWELnV+P7BMLkIZvrQNaFqdGZYWtmEI11lvhYmpX6qwBwrpJim3wRgOJ5nbgQdpiysd32W11
FXpUM38ooNwtlJdpPy5bnh1gTDtpHheigG9FptQRb/+efaLfaoTdT/1B6KGoQVFk1bdhJKJ4Uyt+
eBauKbSqginBmiomrbJs4BJkSLacpQ/naAY7eIYTwhRm0sLDtHVGkfIZDKQCHZsNvW7O+HRH65Ak
5bGQ/SUZIl3JODjMgxKhG5eCGmcoT0JJthxsnu+OXD9CWdhnRk/yXqdPnX9EnoVy4eZKBwfgVvlQ
un3zjiZw1yoNxYSSU99AM1TDtUBGFU+viLLWycwHcsTPkcQXr9Oe4j/GvmhHrxCFS3w6fi/6IwdO
CprKTT0wZdvgJpRa1X11UilujFjqWTXpMTjX+rceDq7YfuT6V/UKwvhia0LMX2gcMZpdFmP2eYdy
MLUGaq5s0zPu3CUIdVLVbJTv2/wfYi1kQ0WX4PGkxXDErela94f0JMZ2ZaswRRCC8yU1Yx0UH6db
atTFU1aPlhzs7RB3I8C8uJAK1FSImSjo/lpbDiA0lE59Mmbb5QMrmwyee6dF/077Xk4pxTpSsFLz
Ug8P5VM1bx04PpwkOXZBL7fd2BYDi7o923CRMQ6h3H7h3z8+GhsA/3a1Gv1LpOkExcKx89FwbjEw
dkbVqhAut7cb+yj9ZrwQ4v3oMf+/k0+456hznLj6nh7Mhqxch9q9bIDDh9Yh+u31Wk7bn+Y7d29x
J4yK0lH6B9pPl0FgBc3DP9VKEvv+jk2McQNcCGD3fKkj101nr03CrCXPKI5VEMto9X+0o4BRZpzV
fA4KC9TyBIFXyqWX5Z0V9kel2bz2stJJTK/Y51jm80nVqvq/w//VpUZbskpS6H4LK6AYryCsKEZ0
Ud853dCIWTtIuvJliaQZI+9ouYEehEnsovp4Z6Ms3J4UBrevwz+tIOAQqMcc+4eIiyzKjwrf6XOq
ow+coPr97gQLxUl/UnSTY2aJmzCkeSLlZuxn1NJm4vCigEQG4pkIp0KlpJV1WBsMF4gTaLQqU+mU
efP6bRuORUPxaM6yZRg+g338FASIS9COLO1jZDII+kv0xbBxRitOcx814suequSr6Duqfs0ud2ih
1M4qWwSrX6w4gQpHOuadp0EKlrhaeEcWmTP0hD+ThnorlQ8OFvtMP6sWrfh0eBA61q5B943XSKwl
OXQu9ZWS2ar0ontISM573dYJsGfrYjuogTwnM+TfIjACJP/BXYk0yHi6zmHFZZelgoEWZtqaWYZ3
lu5mGTrldjO1AqCZYVV/Gfk+uIlGZzOaYmagYQcDjuE7Vr0FzdJ7e04mXJJuySIaOH5fFYQ0ky1P
3rnCRjSKxuQ9E/eYvjhK79HH6C/qelZROOGcqoa8mGe6NuVOcuJM8bAYuQfSNg9U+4EM2UC0ta3v
6Dcydug/nD2JnicT9WqjRkv0+1Q2TiVH8RNAYlfmCqsy1H7GITYErmnF6BWheLeLf6xATBy2om1o
kQxMTrYSFZbfoYM93n+6ctIJ2dtEeqNYzg24ti+OkHjqOe5+8voRTDeYubJNGFVVfuGLcu2a+9Y4
w9DgU55wmOlxjvVnWDBUP1nOZa6OD/teGrV+MbkHdsJDFc7VATOpsw8UvNLrfUqTKKg3v6DYNApD
7z/1BkQCwmhrUhdl0ts4X/v/yMxJpSB3BlQF9SAsnopFT6NefJ8LdHRyQXnbTBa51TNhZWWgxyDU
LDykXOAtFWBAQ17VhsnH1B4BZE+YCyfEBcf2sLvuBdMbF2QzLptfoS3Z0amffr5jf9Bvo6xrZtfO
vN5V5l75FhgFGTfmPRWeNNYLNGHC1LWBSW1B6TeiQ1xPzGV8aF9+hu/S6qTEPEySbOQd2lwHzCXE
1CvO90N5TYh7QPwwz2ROF1Cs3m9HGToFxIZ1octsxtP8IM0ALY8BFXRdVn6ZewSc0msRjuG4ABzm
+G7Xx17p+cC6WjhcF8+ESwB3UiKExOObRvyjY+dOWu4bKSvL1cuQT0jDlMhhaLbjU2qB0MWKmHTc
KbSTzxazIzLda5P3v9P8YPU0G0QSZ9cxYhXtXgCKhS1FmH9yMHmIcxJJtYGBVoNM8zX7+dl8qA/a
DX0qqBHIw2OFwF/e6mjdPMoCM2u2N3fp+nRYhYRmlaTDuiBBmaiRLnovRgoiTnwyuudwJF1WBkJM
1XOHpESXzZeABO2xmH42ofMANPRrPVYVfWMOZcjrcNR8CCmZXp/1CzBOmuapSHls8/9PXDjiSxaY
wfUCCDcRaoKyGz2usyqKiOvufACnvoXB4zANFlbgFFu28n5slg6E8zLSDfqIuQXEtWLxX0YkDZcj
oC8JP1yPXT0SX+M8yVHB5qcmW3K3fVs8fq1xsl7vgmvYba7TPqruvnpjV4xNLW67aWUMjmGYykqi
CSwhLYWplcLhVhOnzPLre2JRNXZqvZJv7MFJC6siq43xgdqgnUgn8IfPYdTq2U3Ao3Q6m84uGL9S
W5E87PAPJcqUoCVAvFVnuXVXvR1lLBKuUYpTCY91SQIwUBpBonGSdzZy4SuCSV4EVF2wqAlTT6QN
U3d5eP94RWF7/vAhfx1iF1zmiFCGDhff4AuYwSxMzYKOBoRd5aYHIjYrybJDaDp23gJj3RFMV5P/
R5wKEuBNyHgAPjYQjHne4ciNBoL9RbstCAsjctfNyVgiyGCux+prYP34ssVXuiOze9lsq46t2MBl
1pYQVj38TWcDM6Q23N9Qpc5Tu0ObDRmRIoFdhEz5XcpNK1A7hW5VAMgUKLG+cgbPm4giyGlRShqx
m4uNsy/VDkFSSj23bA8ywTpMPMfgt7OPcnailPE9o3AekjKQvpM20+zy4Qf4gqsbiCymRlJxRQCU
vnb8XHUn17b7nwJfkaY/X97CQJ2ndsFsI7oZk94i/tDx+8uPELj1Fz4EvAG0X2LUkHDgEHIkRafz
FqWMkMfr4ow7XQ3BwnNe1/Xho4U/CZCn0Jbe4u6O3HaB0DJ9rBHgr3pXA7Nq3+3XekfmWPk6pHjF
zbqc4hFBWd3wdhcWxwPr2zhE1bKG9oJQHnwV2aaHmjQfZU5AoQzqAOd+fTMzp3cY+hVxjd8U8JYU
j2xFZb/eFjWkQwTq4o3marw8gzT3X01qARxJqsF5nPsJJghaXloKlHg9nZgzNY6zO37hFZdfcJz9
5nNr8HRt5ZhjEjBR+DkAl/qURRnEAfsQ8QfJGAGXcSkKETZMQbR0k2/tlLcTTKat1jHrGbnaIqiy
h1hawTR20c5cY1rZsKYIV3OROahe+l2PrBTbXFUD/mBfm7tmfDoVpnpBnA3no6bV70MhRhuosd3y
B4kzYVuwUv9XntbFGS176cW6QyheKSvhVhGXF1/W0cQufTbXSgRzh89+shVd8z3QXY0MIAmbOrev
cZbt025sY6kb9oJd4hbnS2yN244fh5bnvO4bDD0R4cemwZgZtUNWwVywhyZLMmNHplCAanrzXX7h
08iXlP3pBlrAwObq8eidHORdW6rTslFFA4VgqflCIPpvDwpfqbCkwX1B4Gyj/gmwLlpaxTgZ/mpL
7S7OCbcP8vNXWjZjG0hC6/D+FoGiYMUz4AkMkRb1eZt6TgYLr7QZEiK1dyiPPnLA7xFLO8/Fs1A7
NUXZYF50LeaK9XJDdii/Xji4QAOT10GVGHyupVOF3a9RrVEprEDD295WZ9G1ijErrY975jMubSbg
wYD17VMr2jEZ1trI7NT/bfzPUalbAZJTZ9G3b6Z1K2BdYHK1yP2W/5sQfbqL0ZQre2tbtqsJNN+i
xT3FrTZFP67mSVBU82a6UBzIRAT0Kbm/Pm4fJl3SR1WLmiAxchHg8DSwh6Wfr1vE9xo1ereqh9qT
Kx9ZxSnA0aj3iyqscpzl0PGBHrhzzcM4iDL9MQVPVp1mtje1pbNf6bMUETGlDMkdL+e0CR4FWAnH
H+SLpYTxF8/taDxTTvd2l9n/AGUm+6lGNwS8y3gCEtxJ8NOaXOwrtUMgVaF4S5KoXrSGuKAsKkf3
TwVXflugUXeTLG/t5CMF/w/taXuki7hdJtFhSNNCAiDOxvRwxe5FalyDhWtrj67k/EMSqEKrMaSj
h4Q5zBW1L7zJa8pAH8UIegLUmxuLXZ8Ik+fE7yMAnMgkc5RIJLY0co/5d8AE0NhnONOf+VOO6RG4
O08N6DUNOE/n/XaC+gRUi36pERLfdu7Q/nibcDCExw/Pxpj10kddwuvHWBFM7SF6JW1hWUZv/LHz
xrbrZ6JXAowjLyTTmg/M8vRIg8l3OcrWrCyU8lx5Fh0S5B+cwigX/DCt0KhIrTlzgDXmTQNBr3h4
xv7m8reFMjhvNtZ6GBfMFy/+GSpIqB0I1lkMpDZgUzxlP/z7xefUOJ4alnviJACcfMmxeGct1Tsg
HEtgTNNzTOCs5+XpVxpI1h5BA01gdBwnaOmB4czYH6QpqEY60FDGm63ryPq1lj7kH2lQ+aPWbnLo
WqxAHHjLwtI3TsbxUPbcdTWDMEmn/u1yVi4EptOgYI7O+YqKpSKsfwFaOWsN946uYN4UPKrLFuov
yed6VllkCAwONaR9RJ9zVsLkp8YxxFL3gYyttbkuy2YlMFGtjm3I6olxXoEgt73jiKdERmA1M2is
hk0+6W3jRs4SlXFjLasnBhsE3no7/PqcvHYNoW/Nd2Nssz7fTxmTLL4N/Egb7zPJRAiyrEfnmrFm
tAcIeBrLiUV31+fNoiwLTHMYRQUwiOZfi6W/ZMvZZlkT3xpA9GCWVJA55L0anR6yu6cX9uindjpT
NZCcDfgll7VCsNXFhCNUrj/PZzcEIAxKoRKmFZZt3hVv2HLotmkioUmrcYjxz4SxrHRGI0M60YMU
oAz2K+4qT80e2dQuWY/zqxlwB35BXZ7rEgdUF6BHrU3zEQNlseqotALtfIr17rLHuJWKXIjectw5
YSbCAeFgh1sdsgFiIlnXWEkyaNtCD+4Dh8K9iUMNOoRTndvixm4c63HeYgzcKeH0MtngaTh2yXZb
EClKHGsh3jf1XapwlwweYO7n2oLvuimFUnY1UfDnoNAS19rbWMbAGiTqEoIevdoRip54XURj52lg
LoO0bRfgsw27GSIxsWmcaya4n+t4EdhYo4gxID23q+edeOniUqS1U6ez5txNBXBTBB7DxP+lq9Fq
4prhQPDJRp6/fJFLHKelzsLwWnUjHpzlm+jvztl4sE7C7CGfcVxooVPVBFr7yHvFaAF2dyEP5rQU
gIIjGgrY5GAC2ymzgTQ9I/Tq3IMZQNqiRzc3ayXiKt/hfo2/wMAaSexNo50OF4FF1ouHaHdatNML
PSUYmzElapeBnj4L6zaIp2HvhWoGIv2/yKtybGmG+rage5RIswOVcIfCQShSK/w0ujeH+HjYBi/0
dbH4Dn2t/eGkLTJNAXgMamQzXhmjnmJYzJsiBcLfLoPwGm9vu3/SbR7G5SyKqJ39CkRqZWgn9IqC
BDY9p35XwSkcWOJynZHGo70huzL8rFFiiOWmqnNtafUMilJ448kazbP7tzkCawVYjv0y4+0WUr1D
o2BpHSKvBX1nFlVVqnOBRnPTO1f8RVuYC6lJuouGtLO80S1v/wJ8+0UOoZ3EiJ9nqvSxJF7q/k9y
JFbk2uhSYMqjf/s/U42aQaUcuky8fcASBt+tYPZUj37vqgE8ij4I+GCwDjKzW0qYIcn63UrYGTNw
7aXZ8fcCSuF8aAKhPl2lf/rcFn1nKwP02VjtI359jlIL/U+lgkDzicCBs2ZkBbCn2aPxW/K8vkMk
9OelLFcNcjJIIg1y9no1qIMJZ/3watMWlZXbkFqySxttXdPt5kwiTCXnbZ8iR/GVp6+j9JzGRBgd
Pqfm/1/xDpaEQCs/IPGxvKWwYuj24Bgs360MwKoyh3eEDvg+o+rvxlw3CCbP923p3u8xR35qXgJT
L03340N3zP9hGvmUQL0E0T8ildTsDD+hImfIoOgA4vBXB7yEhsskOhwL3Kw7zvawKmnIhN4L50GS
326XKUO5OTe4Za4DTq/GP3jHAISxzxQkXCRrfrXouU+bUQdlhRE8ry4+fnEOAHL5UFd3OmQFAlfE
9WJCUvjITCfeMl1WTUbu/oMk/6iAvnhjDBsi8Ov4AfZRXFnZUppOxV31pY8/7PLRIg6qHtVLmCdK
DvjhMDTGrAwsJCy5bBN9v0lOls+6F5ZFsAgxYyf4A98NXXrQGjOScKx2jjrsJZnCAVxTz/GTN9d4
FRZm4OKqzBMd9EDwkGqf71cM1Vc5uaDu4dAOaiVz8JMWIniWaT8dW0mj13ODTSeGksC0lIi7YLs2
9wXGOXQFMaXN544/t8HnlWpReCxksdkWeUhVLCQrUuBhzZI3xnovMiA8GwGdH+1lr8cVNQc6H0gJ
+d7Ydkpe3NlmIP/34ibq2gmv36CgHGLeWJk+nis2md0XVP523V45oye+xVj8ieunrX4naMKSH8GE
mOCS2hm9f6WwD/HDPNqcZqvTEjfhmk4h+T1Y0tIlhA2Y/enRwkV0fVZPFEv9qqx0R4Nrp161KhpK
yr+bS9SzWakBwMtCf2ErX8pRWNimr6Kzi1zpiN3vNN16p9X37LyCqXiNml/wGBC3AIkWfnqcAjri
8ZKf2Or1tQQonyR1TKIg95/J93YFvhmj0dphg4MjKi8q3qY4WE/GhWAizCe9kIKHQBGiEGvy3f+Q
JF7MaYDlCJ3WwhMm/zZkNeBiiCBhCJCwzU2ZunqI2j26ZEPb6oBIb99y4QRIIk5e7fVkffitEAJn
uzyjFtOFwCx/lGnpKTlAFwXz9DZt8Gke3IfWbDIRjhmf3OOndaSHfCbiIhY5qrDQ6noNSR8Kz1ZT
vEVKQS7OdEUHaw5/LkIgnh57NP7FoP41bFULg4Ym3PrG7/eWS6cr3z9aax/A4Pkt0wxouBvHQ8zr
EDcrGjz3ukCHk0h/oH5yzOCRKtC/BcTBjkMfKPLVnIT6ByPBCHMtNBTvuhP4ehMyt0+RxroPHkT4
e9ygO/wI7jvrMcOTCHdeRQtwMp/MtYvZqthznmX9/m8EnBbtSnqRR2ATB3mm+eG+gwnqj+EvWBCW
oBMjkSSZZGkhdEihOMaec5W5uDkvptFebq0g2StxdHGbi9ttFmyjo70B6N5oub5vqvwg8cNpU461
jARMRxhEMTHDtNvS4FZh7qjXEslZpJoplB/aRqkamLFCISXVOIyzrAf1Ne/t1xNudigqojtV9ooQ
99LrvRFfATL21qhf588VyWKKfTUWgq2EDgaxzuoRlcOcYL5aYt3o5uID0YXq86qSi0vwfYHPSFQC
8yh44xkyndSFjzbDkMbe9QyzgLuhmstqnshFEpDHyQmVEnyLDJGxF61aB+4MsjHsVOcgqYjD1/Aq
bgcbjdxGNYVnwnX7t0ejUQcKWLiX3iHaR/hBdVF96VDXBWH0hhgF5q094Tjqy2J14WSXuBVo1Qqr
TrGUgCgBPxl7T7q9Q+0aLGyQSAdb30S5S18CgLXInlpI/oxcdrVPjknt3Iw+y43drr6X4jL3OuOb
/ZJw52fXVPDREkNQuQD1skAnfZrfpknDsDGvMdyuBhd/qK9Q6SrEtGPNHSWx2Se6g1WvkMqX6GIl
wRU/qV49PajwS/xH9to/ydyD0WAVK5Gc6JWuq+epYy/mwFY5fwvhIyK9+OKsUQNNtobdAEEmXKu9
fkT0xar2bIr4F66v9obFcQJcRaAo0f3kgfHckrXyH52688a6Ot+qUMTKutS6ZyY1gjVNXA0TiwCy
n324O/DjQ4Nc92huV2qnqZDrwBFsOoYuzEYvBcYpwwCBAONar7vqc4cC2bfvUTqDCsrR+1pOXcXE
IGAgGLILZw6uUNCOYcw2X0WBEfHD6yBMH9GV38g6211bvn0j3vMW0RtsWkYtqCP+Sps/VDK1RRxk
/U+NDi5fdQCP76UJJ3OrtMBicM+WdWuekeIyYhShf4wL4RYzZyqGvCGGaus+fZJjJM5teDeySSux
YcTNkk3Xzt1WlWpiQ+s7IXvgzsLwLJCk2lUh8MkEQPaRi/msjeUq2BeCaeXdyvUsW+s9oCstEV47
8UJ83L0URk5YAeyl6+liBDsT3gkuA4HTVUQYDjeAW/wkLjzta3B43OMLEPXrEaXN4cjwli5TlCha
n2qtg97Ppr45htJja+F+O+oVoHuBapzB4JC4r5gE2Kp9Ud9uhU/64Tw2OQk794nh//dO5FJ2U97O
qAjXH+NP9CCSsPIrhXJK15yZ+wVTXNNkCaOcO++jFd+05K7IdJ4s2eaTVyDfJkb0mkXvxxBpp3u5
RMXuj82kuvxH4lU3QdovP5sr60ut7y1+tNaaoemqZJizlBrYPSKIJYr734ZsXA4wT2ymf+mTcnEo
bM+ka2iqLMgHWDBeeBvIVmG53jkZW8IWDC3U9bq//dgIxrCiQ6B09AFaZkDpkXlqr2ip5rFkKUL6
q8lBmfu3kZxm36ur5lbpTpb0QvnubzQah+CyEPpeqLcYBwTCOLQGMeELxxV6ESy+7sDQU5q5GHy4
ge1Q7BT3vLpLU0PRZyoBMlsbPzz8+KvWZ5sM0hWL4fmia4698vLgBfPjh6iuUfxhL2xZ3BhQnbEI
Qwx4Vc+XEZ0JOylWXWp0yTELqM+DwvgKGqsAVVPGyvu6mnGWu9HLC4wbMclNyWyQrLNpwoEVftfd
SQaGI0+S9JFqg5z2pTzXzK0qL55X9chKKM/7t+6SNCYKHXcro2uLL4MscpAq/fQ5ZLCkfiu3e+rB
/PUSctpXSSiqIRK8D6qiBHaVI54lVtG5m8iZ0lM/TMcwgSKMfzc3k7IrzknlyZY7NEGQCUTwERg5
b0prx9O2WbmxGjuLLFOujVzSq2up5/ZfC0yJrAVkhxFi/T9hj2Q6JoSXRZeDvqHW/Vf93TzKwApJ
We8EqLZG4HKG1K4HLV/xkVrRHNQfly0A7mmG76MOrld24QvAU7w4TCC2EKovMxhYgNQM52kg6XIT
13G+NRvY0/vJaM0luCHVkuwCGfAzGVAP4BaI/BZAgUDYAUXN8u1oC3VbxNIwri8V9wT3LTLCkXM1
bX4QbWD6SuSNmKaWq6wYXKLLDZdho1MAJsslXvai19ChJAv6Z96wWOMkrAfj6kV1lAQZUTrggwuL
BwHKJ16RBp0SMEIxO5ibEHQyaAaSkPjtLwKM/KZKFLu6+y5tYA9doJa5n62uvu0g5TV8uUyKAkXZ
9+HcxK1w24d4apCG4y36r1j/kXN3SLvGTPxEuyLAplQDow02YaMofoa+80jjRbF0099wXcPDYkkP
kze/6xvSuPQmffnZQpiDpJIrpFtR+0GC+ej0lO+xbXvFJoDEtJz3B7nYRai00zucEiRYl48a/Ptn
59x4Nq9pDrdMKuPccwRtGjsp0ouOEz7eJKt/o/fU2zRNJnMa+vL+4goI7WGf1FTsmuAF1jTbLRGW
NmWSnv34V/bSdOLDssNrTaRNu9JTIVN6/CDj6x/2PSplZg5fu3uA5p9+qxscIpZp2rpOlQ8vJBsD
i+TfUvfrEhl6XCmEUdnsSwurk+YI4Z8A4N/NnF+34a+hr9vA/zdvK1O+dj2AUq6CmoG9tvAKeD71
aLXu0u0agplbBGEQMbTsOKRf/j/ZqNBhUyov9dXGDNcJqL2FVNiy9FFCnMrhsz8jBgxMQ/V0DHjw
y8ZHR/F160geu/1kOdJsORErgq0/qY2tfpB7+pOnu3kiTXkRoJaMCeElDkTLtLlaGEXKHUdmAoAb
/KCPGfV3hdjsRbbf89sPt54/+Fyla3XTTgednt6WgX3i/U0tk5/RQ2dKZbqHMl2lSTYTsa/Pokt0
wYZtYUfloURwXgf5C7e9XgAC0sxJkTQZW3/OZBIOXNTG3w5zCmGDYDlHy2anDOFNXYnWbAa5hZ3I
xc9JC9HqZG5kNtpCmsqlnnhEnsBMDLQ2F8XePJqxIK7X1/HTHsLUlKxmdQGGwSl2/Uuc9+Hu/Fq9
FaepKDsU/UHjGPTegnqbNhDWU82w1hvNFH92oKW7lMSK0Dt4Y2AcvA2uLF3HXKPbl0NpAUGdVkbk
RR/r7PfzOg/Ea67vwaH8T5ik5TJcNt5XR1OQIzFH8wQLlmTWn4fiotw0csxaz8Dt5b4MAw8KMid2
DelIohMV4uMMmgXwwC6DVwJcA/P3ammLKSwnF0vcWqFRfHswx2rgcW0Zg+KrRJjP2AkiYHYq0yaO
0xMb+F/X3KpLj9iurHpymtMOTZNuNu/LvbbFviFR2j5Ssfh/bDitOx4WDUT5MsrA5Db7hxdKQM/l
FxqQu2C0VZIpnXanjtGrfW58fbELrpvR3cg/1rxoCn+KkXwCulhglWGhhGMU5YkqMPGNWQY6ac4F
j8c31KkRjEdmIYsGVsHRxxNFnD7/zXpTyQlFn7lqnh5PuQoZkUtzN8wxFQGQRGisD6z0RN1/uvTg
EJ8rVjzY1/XhVDtPWSyO9fVm3Xp5B4/MYs5J7QGWnn4H84rmwfuobQ/W7tpT6X5BnBAoDKfrqzsq
jTv0ry5czKYgYhywysyBcxQBCue09ti38UtHSPdujIjt0aq2vZOl3GObmxUZ7jA9jRPxQgoizeTq
O4KjgGurqzONOpVb9YIcH25jKEbjFhPJYoW40f+qTFjPLl0KMx4dcqznnZteTlHjD9BgVuQO9eWP
+QOKgri9o0dxG7GUQO+a+qX7edhcmC2amUZwxo5+FEptHQ1QNlhgE86HUImevVfXughpnJ0ZpDUe
hpC4uJaj37qJqNwcf7revGr2l+x32rTv05g/cYSXYxYsKEQvqD1CE7LvtfP0nKBnPAd546OiodOv
uE9+jdclIVoFAWENht6YeUqEwK715kE6h4qa0jTXLtq6XLvWVrxfNPMrZjCwFqnkmSKUwYiRKyhH
UQw3XqjcPAk6sJjj/RFpIGgNkp8FKdfyg3W+U6X3PbUoUHC89IOmhC6JhOYU5pRvJGXjFvZ1TnVC
z0Pog61bN0sR7oPh2LBP0C5gRTxleQ7HfErIcVVydvLNqS2T4oNvkyDZISyt2Rdb/MKA+Ef3O5Wm
eXil7/GY69A70+flIXkYaxso44phW2IccUJAuqNP7DN6sK5Vgzx5JStBhN9TWyY3f174cgAXqdiW
RgYdxwKjFK8VkT8xKttbnb6XopP9fRv4TfMCH6rsgFnLK0xVihC68bFwcHINhaZnh1Jmic9KDHwd
f/ajJgl5a9gKyeZpqqdtfPmalQOZp5R+ng0Pml54G7tsuXKWNboHAZWf69288DZCvQwQXEBOzemY
LHROnQC771ln85f/sMC7aauZ5Mz3sopZ9BXrL5iXJZBW/Uc22TP7yf8Hlq33+pS2oaB0PBeesJsb
C4r7fwh6PvVfnJpz2fJYC3SwhPIzq9Nt2C9e4ZhQLyv8Q6mDz2VXmoAnkl0FKzf4wndUzd1bd0wu
1ypMVq5tNIuvRkTOBMsUwcznRcR7LxfuVRWcllZFm1miLXPwU9Gjka/jOV6h7E+SUXASNdBTEkQ6
54fE+W/WLakmt2oPYAh6M+sV4OeQ7yo6H7Ocrdz0KuSUXACAwXI1EkD7PcKT4vT117cmLnp5Eepw
wO33dwXJ+PW+KcSAeOiYPCWyGq4/5DJcIWOthDeDvr71j6LQXZKY1Gj7J7IfA4V69QSlaDX/uVkU
+D5puVeGj2Go7RWXvwbV/8DhwGEpC/WjPafugy1iAPQsI9N+MaFO/YcixMyA9OV8loUz0jGD36La
Zc6fxLJqk1xcisXxZ4SYTf8LOslEfNiLFxAiLn7efYfOR2A7LJvwmemr8H6tuZCSFrUQmlv7be2v
seKO1+uX2iFXKJpGdibhE7mU3f54cyeF77ah4obx+F4TwjcxL9lq7kv0FcX+ldy8KgB/Xrw+eLyY
wsfbZFTaJsEcsKYLYQ2khx8rMS9kNoNwO48l8akTDlAyT44iyzSHhRBcZ/Ghwf3wacVaQ/VdDqoM
MuciWf2+oh6e1qle9CSYdE+Vq28H1jkr80bBR9t3WRuJ5r1VCiGV3oLzxBbn/7mwV0L/Ug2Q+2U3
JHnmwOQs3U7Yzy+76m6iQMJoXCGXZruXbXyD1eEOkA+e2uzwosMASV4cuT669+JNYPyb1EdO65Uo
kECyPC3rnJyOsePrFnnVsiIUPm3NCbGaMgoHw/VoHnd7Yv1+36dFNUSm4MXH2+38xRIXJuxH+643
JDqEIO+c0CRxFSgnivNt8RaP2Bt0jQOU+yKmwxikdUKBHuqbdGs5d89Z1vGxlRAQS4U7Ws4taNXP
SmYsEnmxGsZc8Ruy+U9LfTHRPizqrN5dIkNV7Zx8tttL+xjPAQ4MzyJSJl4Cnysg4I4LeVMJHNac
GWofgQ2LbmWv33XjZndQKD+uR1akY2gOiMfOwVABNQsR/ZsouFciXswQPZWcOIMeb2gsQqyd9hIc
Ve6g3dUqmJyPHu8DgqrQaPGbkw2778YZMBjuzk1z7RHN/DVHEFwjuIcUjrZ1fYDbb7PH75PMks0U
Be+3qCxes5f90oAravUPc70Ce7faAX0fLlist4atcMeQNask4hmDpM0G0Dd7YYPFLlhhee6xooCE
E85hh6HkIHxMW5qeNdq/2MoByIT7rd7SRd3lmG04zKB4QYowwlIi9kePb2B3eD8BsU5UVHz57jPK
9KkVU9u7Gn1K0/1tBta9SnD+nlkqT0I1+DL+3ILKUrYvT9VkZ0zaBeqMNWkVkjsV6ksfcWQZ1UKL
Xdiu2nGq+oTHANaj8rPLnrk8BSdGo0GTglOZD15bHoqIcrknEwOFHl9LsFYluMTTxNP94JEkqhNV
P0KB0puULbO0fBanb3yo6bnRr8lSBwZlIxEw8dc+u7naFuSvxpAq6eWhzIrxb07cNYHgwpqBA0Q/
0CfEnb531De6J69GWpmILkEeKl8emREa6OFEY7RTQy90ATCQOANjIQHfQQKcI/pW+wIJntqOrnb9
ZPI9UXzzrCNdiK/gWZL4b4soO7TCyxsYtOPlDFmGEItnAmqZO2dV9TPsCbDQJU6hFZQDUI81akxC
622p6ia0NG+RtKMhAbpFp2AJeIKojrgq6/dEah9vDapO9UEI+IOcBGt1ZOweLtIk/lwpi5uyC6nF
DTPLCyV/BbsSSxou0Sb/NW0v3hrau8RD4/fo8dS5e2LWH4hIoGBuUgh3thDLz5oQn1lGGus1WA5Z
+ciXLVtsAM00l06opguoauOCJrgqXHWNkb9gUxi9Ph1yg7Nj1IK6dBI4FD8piG06vNNqss+80kca
g4yEDTRx3OXASdjebeiLo/FRLWF6jvldhav84oHoDH1X6v2Thq/aJUTQ2R+fIhcSw3XRgazpIVtb
Y2WWnO83MHjllztOWY/MtBhqM9SQa1rSvMGux/ZzHoUzRRW7W5kVsNlkliKmvYbySB45tGLKoFZS
zYz7sgebf+OW11zgv2n+GokQhCZ3H0fkLSALhWXKhhDyDFo54Y//t/2P/xhkHRLcX4b6LDfyca92
r+37hDChpqklOSGw5Btw46kWwdiFniiHyFVQloJkwIp9DlgrnFZRGDCF00nwujPYAl5Ys4cYIf/f
LmBQ3yr8SCBG+RvO7HOOjSklgdEJS1K+S9iL3GzPqQQO//rvXXo2/4gttJsjRmX+fqtJ0s+FMCof
7h3/fXTfW/ucu59JOSOkyF+e0ajcmzi6KGwWb3JZ9b3JLW689gNnben5SV11LgLH796orCgCTW8O
o8fihdEzQJN9vqAy4znaGP3dd9G+DysDW16emAVC5kgzHdaUd3p1zBsgyEBE3Or6nPGVX87kiBY5
3mKGPjKsGzAMFKFk11HJ6ixq2BjAQxqy+8Wo0jBywRB/az9UufWvvqCkiMVnIKQUaxwTayTyowzb
cL5A9qsMJS6dZZuUcdx0N0fhENx5PRwa3PU30fbus5bQJLUzkiN0ERbKbIJ4IcI+xfb2hIn8b0Bu
Y7eu5i4qMCZ0qVONsJ65uMOXiD11343358HDu6em1iAXibioo/DiN+0tnCu5j2cYfW0irQTqxkNb
UZuV/HSseRpPt9Y8FNqOcqlaTtZ1Jwjtdr4zYEjfoFjfjksl66ouQ/tRYT1Pz0MYOYEt7JkdAChb
mdM5Sqy73ZuqQqUuPWssJt3eCBEaxzgqhPFikK2tkZjWdUXdswqEHCtkabeVL7Mnl9oHrThqE6WQ
wR645GLQIXm+NQub6WdHW8V8XxZeSt3ULipfJv9nsEdKRjTD0gPmQVjyU+5WdDhVsFdfWwXdQ8yx
mWxttFsxuz+TuaYPBWdxziDTntl1uMzI71wiiCaEjGCDHQAFAgnCSxNzptVtAZ3T762tRl/d/0g1
sCdpa4+ndxZwj004WzGXKVaeGS0EOTEJxf3mDJu0bqgaC8pOsN0t9cmWicEXkjQAEiMLIb2+JLsN
Zt+9nT+5mpCTDg/ha/gDT9RCj6YBLdiqi4zXapp4BdEqpmmBdmLCH9E1uBWRixRjDp34x3jWLKdh
AWZEUpRm12yrZVdZYrvUW7x8l4PhYKv91B1y9FAzzGGFnLj3+n9jXQt3v33j9zgkcjo6JpQmNs6f
QsWAB0k5C1zCnoikjne1/WSlUxiHm/QLCRe/2YPp3QBxxGbm/bxSwC/cCQAZhCK+1EIxKcMyoZTn
c8HK2apw8aHOmhWBXYMdcYST0e3+LmgWvFQtBIqRA0llhNt8dxAlr3LxOrDe+5zuRgTUwsze89hv
etiszmznM+tjU4PMw4ZR9ZfDkDm+ItPJRF2nwdcPW4Tdo7LQK+ipJTa32gUSDMPZXp+58vIOd4Ky
aO+M7Hl7CjgnUhBTfKOdBj1uNretDRd2OBHz9r6nWkiPb0GEEWaus6AJZIIo3XIS3ovY46FCFjE4
ulEPeKONXxf5vc5NeUvGHv3u/JixEz67qDVGSgz3sMxZ46WhBhzl7PE4cnSSJZXoYZqqguOYyZfa
RNUrI3UspthzaDm4q8YM0r0AuPhYr2OEU92CxULyyz10v/yo8ajdYfNj1yr158XdpDrJsbf0ubLt
ghiMxx2V0HamC5OtL2/8aWjXDaLbPW8Vd5ZlkuTwjzoLJxy9NBGVRLjAJ9HwSN8wxGZsLnM12ucT
8FWtlUHA7Oa07xAog6Oq2R+PS++4JC1lGMliRjMSHGy0aliChre+yDzJcAn+9TiECwEa92tm4EmF
+Y2k8Qsk6Zge9epkK2hA/3NhBtwLKsBc+9C6UID0ET5VgGvSPlvHUljdSs4HU//JETXzOB6+aiIf
1lkdo6oXqnw4fz/u+onUeTUVif326K1Q9a1rg28Ma09j0kdVBEdna/gOiZPs1TMA/i/WxWZ8SqA6
44ZKnrdBNt0xXo/WSTXWDKakodX9sdAREAa2V2OVKfIYtC0zql0zZYgQcSp6loEDYXAba7JRno5G
sq5MTOLc1O7anM+GNOVCInwI0i7Kz5OyN23KGxTIdWlsam2+Pr60FYCPhMxmGEfAthxtdmbb5r6X
By21GcUqkM293zVG4j9xq4pfSGfWJvuzZfocN57+tY4MNnqZO92CxJP9E1Mw+pORYCHUgvaVPV0k
PXDv5GnstZnEIdrtEdCvH1x3vikv3IXQPUZJK45CwrQwHsSjRhv1YhQuVUl1dvvF05zVmZjFGNM3
ITuQwltBWLH3umUVyQya5DEqK7a1y8GXrOJVA/qjBZ+ctfMWC8E9vuwZpvt0eSCnV2fRhtePVLD9
8pLEFbx6wMfpBF0EKP4bDxGBCdyQ2tYgFdjfytXbvYvKidycqoKT/+UbhswN3QU+KpV8fXAhl+7/
lUtcaut+5d071u6SAk42O872Yj5C7ZAorpy9mVgWGa2o9NuMWgwR8936Dsi61FJOgHl3G8ywFCyi
PgNeze9s9H0o68NQZVhpHIXuhqVVVBs1rOCnPOwWOZP+h1IaUvJwNBZKgTlyuvpK23+tMp6E7Fgm
589H2eEBKBibdIezkg2EmqRLOWNSBn87RDwuAvy78YlCgnwAQNd7K8dx9TN69y4Cwax6WyJv0s82
SA2oT4MgmraixXwhnPRZ5G64a2v6zL3nXtJ9cQnc28H8wf1Oe1meXEOxNdn5Iuzfds4raqGpJwdL
IhH34JfQKWNkxDLWYt7PHguVtZaXqbHPJ/bSwnhFx/KcLKowxvYgsmBvAVepOh/XN7WyZBgWUF0x
xk78cF7XhrsuDJ75lKdN+te66qZt6E/vHV7ZIoDKOzZuHIGblyNX2sjIgdWEWn4fNMc00YP1ZAxP
KYu0eL+C94hi+dJ9sU1mkKV49UCI8k3vRlhbWjTnu5hAIct5rrxKW7HzhGy591h8x3ovp7utjhTq
JQhfAZ+a3Dm5CRd5+8T5cymuu+cmy/Qs+UGZXiebFiFdqFEDd/0OtzMGdCfWS8OtI6DpcuXDJtkr
NyYL8p4Il7Bx7ZryQWNH9r1YdOcugVLMjhXRqcnr0fQsubEb1jxtbW6HfEioRrB/DMmiIRyJ2qhm
LkObWDOmdh3aDnMHCvdq70SoxySeLliPmpp1LbC2RdJe614wY2DK3YUzRuQdRPOJnyz6u8LcdfEp
56owBPFvsoAOqQ/MiZZG14Gh7n3fdymtWFw/pDb44314aJ++Tdz276Hy3fQVjg9sztB4WHU5Lv8v
BeRS+CMiTCwOlSW1HlmcYoOgvjOcQ90lyXrna+Td/Nupjdh5DZ9BqM5T0OxhlX11R1kFy/MIVN5g
wqZXOXzQApJZEt2WM6hMgbqz5sXEjNMghkFwewPo49r4NhJ6/lYkKyHHg1rPyERjRlBWhPbgQnZ5
sHbemaDTf8aU8ZM4GA8kODrT4Wse/s5UQAAGEcV5vswT06x9PlUpRnpXo9xBKI56eBR/Kd9UXg5H
HKIoreemXywt7RAKfZeynweLzQc5qCBuog2yd5gtOD99avoVkhEwyeUjUh65yCFF4YhNfYPa8t9J
JD0rbBVUWklbn8om3cnEpYqA/DRQ9hl8H3O8aTmiV3az7YK+8JDZKTHPr42QPKeXnF6MX/x0Z7YQ
kiuq4oJsqJhoEXUnB5wPnFaB0ou9BgWbQgn9hlCKKDs8VHivVr5ccAih9wXX+F6wOfCb9ME4inuE
UHXPVojuhehkTgD3stdjBgW4y/XBPhzvGIZ/yU2/VzmBFzyk6yXJGgsA/vg9rrhM/64tdFreRZgX
KW3qNmCLk38KsDlDYaEAxKF+DEBDNyHXI1J7yzzvqMQOmcbazqiON7TipJY60aELd0KY0zOwkA+X
ouiujLPF+220RoGNteFkeEKDCcbVnHpY5EwwRaXL9qAyIf+uU4QHTXhiXQoDZgIRp0u+6VAK/GOZ
N8fDfQhpLuy2Og906bDycWJU/g+4ePx23kFwHZzhD1HNPVXsfqgWvurLVfiRYuFoDyOEyb5QJ+Ac
CMMIfSj/e8Is5VAYecG5Bcz58fvuj4ZkVWMr7LM+pXe2qUfAUH4/In1uyFLzpxgZ/zbxiNTnYDHV
EJO5S6bQO8AwWjeOZ6oef8PO1tYdqY0BOSie50AAcBDhwFZ2plMqBbp441eMERiIExrowaLUu6VT
+PXHzpejXEkxOyvoNLbC4SLCOe3P3AqBEWFFETkJp1gbpffBc8jfJIZA95sxvZj1NFLgKY6WLFwx
hUNrFOuEW2uNV7SfJGD+OBdV0X3gXqNDAT3RNTFNe0Z64MU0fYNd3ZAQO9TDyjDiE9f2eQmnhQZ3
/lrMv3ucnrWH5A7/mH4/aFC3qBSpcXND+xVGbT6ULkS4RQwG/8CQpz2AEM0clKXreGlfFy1i0fdZ
h+VxN4wEH8wjuTqz9J4RShV6mPwFuN5MaSvqVCBMU600yoSSLsvSEd5EdeHwkr7y64dAMbIU4uRH
Go5+goVjKL16K99Jcpdd1IQmXnQF9mMKh+5Afpurdq/Nth/QQKLiwyd3Y2HabnE837D3jWIHgHY1
CHA2tLeD2w2jH+W27Osf9rY392V6cp8MOvFGaUbz3eAsVBBQ0UXJ1rYRixT9AEGq3msqzPdsddqm
BC2YPDBOAcbQRSLoAh28//+eLihrGFrPJ6JR+XW3X+v6UqutqFWt7q5qFZ42mYzZBPnHohtJf9FE
3EXPDcWcC8cu0Ak9lWW8gufOg9izswgp2mybCh7viDHJuAHW291s+JERCTW+rhEcVs+fyG0/DTdN
H7h7vDHGpRxW12MY8G0Jqze+nIqrzacd4rneuunSMUrb2MYLVJnAE1ZTSas0SfsPzCTE9ovKUpOq
qkgle7xVxGCakvlNg+o3sHX+BU+3YikmcCXuCQRwiDE9wLOhwYMTMAFA55jJ8fXqKzcvah1LsdQf
LkaNPICXZAdkNPRmwwjUThcjqrml7bzboAPB21Ed+ECfYIMwwL0w7/A4S41GiBzQ0CyK1BwETI3S
qEEHElLHRGqMSLK6taLRy8hK5DOynTx9r8y/NhRV979nFtJ/YRn9roYOHQ+ZAX4k1LJ4729bpsy4
BopwbTkgjq8UM+WUeY5+Q0SufdbqpghOqSAvSAJBIepl72ScGVc+H7Cn1Z21/aVHiR0dD4ahowZ8
bOoZAnnNyct9wcIyuFiqaoxL3MzugyUD2jHFZa7JSqtu3i1QPqOYKoqGiyCU70Y72cAs5ad4kI1h
NMcc/GJLP0svtUHwiJL9JurmOo6iVeOChz+jxh+6yz7Y/aywrFWSbLjhNGwLquf3+8J3VL7b7T7W
loa3/WAPs97DmJerm/QkgAtAu//5iJqSvHpW1aP8J+Dm3VdeRVsoV2yTMzctcmFAN0kTcD5wWLAX
CYb5j26p3rQYoVMYgImnq7mdi5Jb7CbLNEjIk7Hk+8fCI40M/1xj1ZLpMnl7gSxUzx4u55rD9k4u
tQYtIufiF9moDMdJQ1Dt1R+ffIW7D/H1Y4bUy54hv5aEd4AFax/hv/ej1rhDn621eEJ4Tu97d8FT
vUhiwkMnzTmdpNGE7vxM3moOUp3hYzL4+ZrLJ1N+g+32JuecGkBajAb1xsVZlDyO46zI0IoAZAZ7
ueMSmtnIacY1BvJA+anD18cX2/FOi4kaKg4pvWl/GX9/je9ARFQbsF1tXHc1Vq9lyrvt6TiwDxuR
x9TpxBHm4f89AVv3UkH0HYQJ0yQ0DoHXgkyGXG+WgB96y7pdRpMQCoE3r9SZgFG2Ot2DMmLTtajT
3rHD0WcZWamiNwrnnevR4BRr73UAbLvGUPv/mENqA0pHMYBWnJ5cyivkZRK6m9LZjQ7lrdWDkhZe
y4J00BokzHqmX8FiWJtGCXJcKNGhjj2zA5CzvKKpk80QXfdbPV1H9v31AAm2AwPw4MlWra++KV16
DgdSbVDXYJz0E3R+3HHLtEDUXiMV9dvq4QpiZdkGAs4pYbTxjE8dzI3r2ubK635KdbhsO7Hw2sdx
CAR4bWI/LuQ8ufXe7o1y9cJ5E3tHdru2EQNdc1S6hwcgt0s8+xsJZAsEP4inbhH5xdc3l/cDPJLl
806PXCGFp3eNS4GfiGbIZ0V1c3MQplKR7A2ZAaQKsr/JFaXmi2o4/IeM5Np0LkzW7pJMLViZzQCp
KILEyQPe+5sqTEdupf5LI9Y88TmF2+8BYo4AA7TsWWIt+ncPk6OTK0gJx3dxM9hhpMDUqZMqy8Dy
WVLudHkUBd+FQIfUv2VVBEaKk7sSoHSfSYpMO2RNlmPWWX26BwaiprE1NnXayzB5uXbDgtAuq5hL
g5OmmWukxftJbWiyLVwFoOQF4qwt7Mzq2ASz4HCbIa9FIrqvx6Ym596ENuDi+bwJ5UXVfBiqKj0u
gN3k2a/ZhryxShgkqaxyvn1HBq+D7kLp28tSzctpIchsXcY6AZduHYx+crzPj4R6GWOp06xa+D74
VJ2eOsQzI3EsCEJKALcA3A+jSGg0rHPxmeCy/BleIsjhqd0NuA455Dsr7FCNrI5YKA/R3NNMuUw0
GBxAhdQHdXX38IJAUkj1mnatYUPyamKV14bRx5kTojYGCCtPmv8qmb4rvgCgYmkDhwIbdihYPeHp
pq+R9kUdrohXXS803dfkAsXzITzUnANqO7k757plqWrjWacQu0vP/ldaoLjdqFo7gW+waYwlHtP3
8O+DcTnh3DWov0Ryw7/lOaa9j5t40dn1iGN95hXDlbRGJ1dzWxdjr7Ul6wrKRcQpKwpdc3Srz6uT
XhgPfmmsiDhbVW0ObZEsBi92oRWStP+RNlHgRPMrVpQk+MJpo92EaWoeiE0u7SKDrcwkP97oWDLA
0zICAsG88CRKr4cB3DkbT6Whf+9poehh7zjCENUDSTdXThfsj4OiVzs7P4cWu8FV3n1pA2wtkUOo
+KetJZafGZ9yTMTvP87/tutlJ9ppg9zwNyNDr+4jnrl42CyB6998P1ckutw4AArbFz5pYTXaSjGJ
+34kmuqAW3+awtWAtCOgXHvm/KEdCrjS/25yq8R+lprs6GX3n7C15RCjX4gyn1PRxFYwl35QQZ5T
QqS+xG6WscZFiVg6ys6BWh5w0q8+xbUbhuZF0JjpQSAGriQvlXYQ9mE4n8cYdT4z8yHNQ5gahj/+
v3Gv8ZG2vzm8UUih7oS6CE1BTYdYhnG8UInXgsDdaT72HyUQk92IDeewG3zXwzpS0vQ+Nj0rC8w8
FpOTedlHIG9OsMlIvWLkEsVbqCixDFOKXi8sEwO8hC0WWoSD4HNnc1vcBMsBUqCu6trUGbmt3q3T
fczNJQxjQT79k1axlUtVwFjXNct1VfD/Hmvc2Ml1VthVL3dLGwEIEVaez1MRGI5uB9RibqTE8raQ
UAXWl2uLEnQ6WD+LTEE2H1FuKTUAU0ixqR2HCjKDsK3oVBrE0qbVnN4P2ikf31DWw4TmpSHcazfA
ecTYxf7S2tUzuiJxiGJIzXl8BbZfpoG1il7C55vGteSmmc6b5X4KZ+Ig9ZuIwy9d/PzURljCaYGn
uBpIPv3qhciespOXzgrZDGYFLtTWv36fduLuuTNwY+IpQtzTEhLs6f0ua+Vv44oTMOSm+RbpqekI
WPGOHn0dwilG5VrqRmLGB49DEpjNse2ANfOKADiygiXMix+o0hebV5iyFzwxlvYDu5Z5o8wK/Zi8
cIhSWflWAc60jAt7URkf4IUjKaudTHNTthoclT7XAEaW6K2RR4n2B6qWLrNGuQ5Y3EwUrtVkjN/q
EoTn8O3j3Mh3Px/3iKOsvtX/oMfeTPNFqMR7DhqQIGOVf7JCHBiNs9oSOCyhTZzcMvsqCkBnkKm/
0Vv9G3d+VxwCtud8FruAx93dvX+IQrR2MFDrt1TZApQFKXgzEwLZuCLd0wIiYkhNSspkldSP7zsf
QxdJc3pJVVymwVyu9Uni+hLeP/ja+RiBYxZGnJlP02l1pKitkRs+59ICwZXSwu6m3m6tuNJe5alJ
wcmdD48G73K5OS+N7SXH1XY7gHEOMwr6ulCxjD++lGGTIan+HsZvtZupUEmOefOn2NOlcCVwi2MY
M2VdtEyq5bZYzhGPa4/5REQ0jNsA6cHk9lOc0Zd4bCVjWRlRwH2WirrStyPEqj5S4T/7BJXXween
2a8Eo7BLF1xtt/iOlB7joUf97wCr4V559/sxMROTD7FRW+AqkXReZRNzUCQdgZLMjJK7BuEiKPpG
ukyoaShJSiE7SL5lZbQXRz8KDPzlSA3OUdix55x66quU+Is+HSbjs0pIpDLImdHg/98Uk+TYfSoV
pDpycrhNyCNNsEi+S0h6HTiN4dkx/cjQsHuQfRkNIYJ+b+hmRBbY9wv67s0+iXXXzYfG2Jw0+dZQ
1L9j6Z+FYWpPjlMfQMolWQfU/umb+hRStt6umckJNKWL/8oyonHlxOu6PxweACVjic8tVN6zsvam
ty6PvyHZ+cf9KtWp6uQTbuzJAIkg+8MkNMmsJKx5zQKSvrLS++QPDbpBh5TuSIkY0j/Dtiwzfzl3
0IHEOyiUCOC1Nfk8PXnQY3pu+GkO1HECmer2QrJ9XcQInqnSRMma32gX8cyHQn1DLuz7onU1q0EM
rEWgdvqsQnL7VlP5PoAOpnPk7bjwoiamdK3tFn4R6ICEmnVW75vc8X5M2JW1xMlIEIK2Xp+FPXNy
aAuqnplyHJWpA/MmwB8BGKsbM2E6taz80won92ztozd9uFIZ/SBg21iw2ocYwS+lbMw+eN689PoS
KveE4RWrJJoaormJXWGBF4Q252/axHbU4QzWZVzVRhB363Afb/BrUrIbe2bZKdWCcwmqqC5LIEP1
H/tW6l/0tfJ4g0qNuQ3GG+Z+SrtukCouApms99HbI7hXxO/FLeOdrqR5NpFbhKYoFnnP754BVNRw
umxK9TtMMBulKlxWX1s6kgPNb82Y/J2f9xRYUh0gscIksOXGUVQq3/lXB+8aISTEPVU6ndlwpQHk
g2l1+ZIVNpwQL6r/o2roujKdbCDAG0ALNTV7xIDBtTbWoUXrZ9WDEUrrEiHOzHnwMSxBzGg9DOf9
oYPdqYKscUsHTvAiQS7gGv9G/41jgLflzwfX4LJEWwgl+0U+oozFTnlrAbHJXv/y01BuPW9VSPc8
TWyt+udluIEuS0dFp1UmhU6hmmf4EzGJWFlPkiCqFYFYVHMkhWrO1xzqm4gs9xAb/k3ucSUx4Eii
QNMAQlwbUhLNAP9/hAuP0K0sln9pzVCH75G1hjpl1FWJmBrvEW2iQdl4OkeEekYVVYhpP1FnwHiX
04XkkjSxxrKcOhl/1+F0MLhW/HPpAoZjSdEh07kilgjDqqlkmIYP07khdMoYRfHZ0hgrTXpTxia8
WsHOS4lYKsU2iSlozVuC5egmZ77gm4PNxERwK3EsxDtJAzu1iQ84gLTBAR46Jb6t0ZQbIYP32YLG
9bAb3ftyP8Wr6q/ynQrRqc/vCB7PiAcdC4S3pO0uai4U1neT+TZCsGvh3LUpXi8w1636xfO6u/oe
2kiBfXTK6Fk7UYU808nC934E9VVdHJDo3cfQga8kllIpqxMmlabAh8MMKCi7G03TqzJl3kXvqKTO
hifm4wR505y/X6b5n0oeXp01/oGZ4XT3Nof2RiRm0PsJpyXc8zH1Q7nRfM0+7/XU63RDKwCYWa4n
CfIEMldn0rhzOyJA8Xtu4uFbHXGoN1Vy9G9QFUA2EfwfXvzQpzObE0wa6ytAQZR1bhNijai0bjYE
aNE5AbcBGCV7m0LEo+tKrxuTqg7/71DE36nZtN2SshRdCgdOspvqACeMehnUI7b/XBonfuPzp3aC
B9XI3ox5N2uY03eyL8zaiU3HiBqrH5rieWChOaIIYd2knbtjRoYfGXbe6sH+xhrBtFoSW5xCmww3
riwe1xWo9xUtsbQWifB1kIfLjllv/pLunO1QWwrYuY+JCqo+YU7SHJDN/0LpZb9YJTp2npf3yfGx
7fXb8qldMT1A4Pq5kclo7eNJtCKMuDHdpELezKvgWGo5f7cUZpilO6s1moZKkEqF2mTrxp3ep2sb
gNgl/SAoZPjOz6cOHqQmntCwyOsoXybfga48QJBxeyCYKrv1lW53NLIOsL8eCmKSYAImy7pOo/GO
wF8I33KLhuXDq0xEeMgjOiOBFrMHSBP42hDpCYr9EyDPxO/FwFxGp1Lhq2m4U+TtgXjT6o0LZ6Z6
DsmH5TSg/D5TqYQEha2yBCVigJFjrB9DXeb772o1vecRvIA0LCEqOt1pgSDOFwxR1PUcSPihMcDQ
3IqZZAoaRTBwmTpsin5z0FgR0ypTL37hXV96DspwRwhfsJt/K1FuJywF1t1ZkrbqMb4pVaebvPB3
sNeWaBlopUxJioUMdG/BRRGMNpS3Szpv9sDsFbV0LRUgDiJa0gAYWCJ1Yo0l5e/dJyH847DXQXOz
qZMf1tQYqcFSNMz8+Rs8APL++0Vqkw8iRFvNcgApd/cYZWFSvFYoJgSb+/x3/CkgQX0exPvPeLvg
tRK+tcmB1MpVDrkFHZyj6+B8L4Fua9N4srmoTd9D4sIQQa0ZBTnnp3NEDeGnqoRKoc0EysyIuaCQ
FyNGuv32aFd4F4ZvNK+HrVnvDw+hecCT4UstfxY9Te8bh337D1fKZ+Yiah604BHrmY+LJ3K0HTzK
PoYohj8ZhpRxA73CwVgNHYTUtA9SDBH+JSGWksNKl+3Htfg4tfCH6CInDticzodP8D7hAYoon/sc
GUm8BboaBfkIgj9mbouBX3Xi3kosj9jQhZ+fObA7g2oxfkhHYAj/81JePEYiz3h9RubzJ7rt9c9m
nRVxVmcanE8ggi2Ordx92Rgj4p3YlGaIcC+PEVNWEVRAdXOSP+YmAoEud0eeTjEOKH/f2ueaJQHq
L/Fha9OZq5sVn8cozI8Ru5/On55twrBznLCjDVKK82jG/Q2BNis1EVpHilX1W2m4Nl5+61EBJHFt
e9T0umVDt8fvj/SLStAAiVdym5tYF4DtXyg6qMkYkOtHovUF42tOyXxsNsnkyweuTm01hF3KCqRQ
pX5Ka2uzIuGq0iNGcpONckNTqnnUApP2sHTlXmP9AohRyu2epG6dKtsuuOueVUeAzuQsep7HEw60
WvI1ZvB3k+IkWlrFcrYLuRjX0OuF7gk8fmZ4NKSx0DYzXvYap2Dn5vLTGsVchCJXEbvk8ErWvlpy
F6w9qcGSASbEWCIKAHFXuP4BP4TKJqaTHxP1+zCHhn5WIR8ZMU0jRgTVN/xLRpNOYw5313jLhqCT
yrPENG399yxByojKXM2LR8IjKlxxaP2iJFHe81CG1Hdmg1DKcQjufmulwCZ8FG7x51u61E8jIA/L
V7ZOa+iIZdAicirZkQtwopgyJb0z8SD0Scw9r+usDZJOVc7yk4qvkYIPE/wQ0vHq15XOLtoQ1+3z
F+eyGwgl1zjGF9sbY8dFsZnBYXQQWfAj8vjbf2wi608AcgAudAHPsoSUzE9Od6xpm1XK5semmVFX
kf5MP+2ajhUHc6JQqKh6WqhJsw9JptOe70a6qFJPzU4eWxgcpIaJwR/OrV9dfDbKyA1037OUczZk
Lbe/LF6mP6e95iL69iyYvHOLiBfkQWgVVZVblSxWhYIoG2h9vL5frq8tTRO+rk69mJhsDMvpo400
OE/QmBNedBhILmT52yzVcS9HojM/BSnfAV3dJ8YlFSZLl1XdT3EU5EkmJmF2+cvpLtay1yg/IWsJ
q2L+gNNn1d617iSMdiiOjo6BNIqLvHOkxyBE0wU94zZszj0dSywqvJ1BfOVs59jaeElPBgQblPyZ
OZfPzdu9CIMofD620jeNBpLOqiyQntTCGCTsNm+lns/9Osqw7i9lpMkvVX/z6uYFS/kX8O4PDbdB
x0PVqtQi4jIrSG98wJxGBfxDemVf9Mugm/6HNHjxIiOrn6BuozPoCGGGEh+sS2f6r1VIhp+p2IJI
N8f2+ILHd2yGk1hb1gOgXIry5ukGf/cxGekw0elByqQqupE85UIsy8kLHU7IINPiGNsemmFFNZ5M
NS/05eT3We6QXVNBNrfOSXYQbrxO6fjXSRi/kdgGirlq4D5iLoKydzP2lWyrD+ToY/P8ebVjut9y
89y+josxUrAUNfnDX9MCmViE0pLzSBusknPeKqsTB/F5A+PHu5Id5nhDhUcCOBHX+GUNGlDjJX3G
dEs9yjlw+rr8m+b7BbXOn7DUr1xvZhCuEjq2XhtMVT1cTUfhks8Xi0kLG1QDHS2HEtfq34WtEP76
nHF8g+ISJWjV6uEo3I8SnIOt4qLvguysG2n6a7DibL0KOJWVmP3xjG/P+3Bxqk2Ere9Pps/BFoXo
Erog36tk4j5PY70fjOUQe4XnkmAQwvjIT8FigdXfs/TunTSRH/OHtI15pMVYU20erS1gvfNDYqz7
pFa2u+Ne4wpFk2IPDG8+Luz9vUOphiyzHh/iuz9ZhkjOQg04zdbSyGHkWNGtl/3X4kN64C0xO+qC
rGDixO2wM7SPBWXqWRo13rrEfRol8wRqaHm4j72UXA6SisnMYfOoNMbCgvtAmK2tu5Vds/u26zOT
os52H4n6KS5VZM0F4G4UaUUUiUyK2E7yY0RUoeRpErOCHrbF4mym9bQl4r6ifB/bCJ6cAZnzq3nj
6lts1ZPxYF0Lm7mUmhvmh5XGUhrCt2GhQ5D0MU2Ww8VI39WSJXwKPs4MOZN7iVSLXjlG/SsPV6jK
5jqZUuITAN0ooYtiM95Bb8sw98nwEPrfc0aSXP2RfYTdXfg7uUCs6Gd/rPZM3K6lEnVg1ZmeHdzm
YmfVL4t0NW+chzFEE9hrgKSMhepa7iMJS31Uv6deRvNZ4XG7aYWMlYKp5DOEWX8bGH4z9XU+UW8T
ou1dKzqBvvpFmOtURd5ESTTYI6deM3uiuIsOQP5RJ+XeXSO2DpM3VosBDtd9Huh5uwac1xL5fv1T
bQLK5cFILoOtufSPXdQ9022UiGVcJdNr1OhrP7mvDa/F5i+U6tbcur4SPAG7HpNSWwSddAJoz6vj
vCl7U/H9Ml7w/OPWvbZzLFaY8iAJRswXoe12QGvbrxWbxR2++R5ycs88SICf7CJXEtp/8bOYFAW7
4ILnVFxKoM7gAaYnm+gLVFCAaR6wBbf63lAugJXG4bv0bltiaxuLeL0K32R/Cs3TiIB91H+cM1uk
+cBpR6QHX1GkqcNSMusPmzRYGYCtjzAZRe4vDsRzimUtlr6EVqS+WE4xkorLP5BH7bLvXzXeZ7jh
D3cNXDt8A5AaT+tzfDpuFwLiG4YSiPBtVSPIqTKFMs6kdkiebMgMEBkpV6BZjruTiY3FDvEARU7V
Ocet8SS632iwEw/2breZt6wNfLmiEZswfnb9edojRItlqC6OVjk+K8ojFThMkhGpV3pLRxeAs418
PxoQdVZnDWq6MtAowQfSR70CS4+9thxQKBB/jK62bWDiGcYnikPXfh06C/Gvy3GVPOUi28Pmlwhe
UQgKwRWkOqV0vwcHTrE+0poOw2mZ37GcCK5LdjeT2CzqqwrDaxKNzqit74bo1NDJaqp2sn7rWAJZ
avzYoqYYiIPJIMtYKdosV6mH2fNQzBnPf1olaxCvI3yOBchLBpWi5ha8I3gLn3z39TZZCzLQE1Bu
5LBDaIht61/sghIY+3GwtKh5fYAMzLUsdA3K+358ADSQOCBTjAmleKezok4mgkyMTXepE41Of0MS
h8Yy0T03nCjY3rAt9ZyVY3R7pjUU5Di6F6as4n4lPTEFWr7TazsGiIRdguZeaIDipC8klTv++tDE
1iyTX1m0dyGVa5tZ4vrm0PbNeXfSy1EFWnNb/y+Y+NtBHK33VWvsMuouer8zwzfWSoRO/hadyh++
oNdVjkuMRv1ppuLUayb43jyN5z+Hlp/yVUemb1i/Z9C8irp39CRXxeWNpGeZ8QX+A4iDBGPDmbhu
lXB7qwY+AC/B1aA4HHnHlqd/F9V5HgSRJlJTijASA7MC82Gv8HbD4HZAjF4WqYetzkzuuaIIXTkS
uwvk968y48pSBZyWZ91iqVM66A0aojp1WmOtGcrciz3gjF9nW3VnZDE9/3u6rMeQt8xKWKX5N73K
5zB4Ss6motOq8hEF+ttvyCIo5PgaxGVYpGdTL0jfICsiTcSpO3fmUI8mmiUDI+PKxDhwew3Xa/zq
+ucuZySrIB2Myb+42unXNMhUh82PWqnXzBKs+AtiEI9fN4R+bLRr7VFa7EvTyivzeghhnlXgOJ2U
teg80juTQtATbrdGGpdBcprW/AABaNSX37HlxQ+T/YNoEH8FHU8EAnaBjztPT5XPDZdWjFJAEfAW
rF8pfFt3rYb3b/hJVKfTQqWTY3wNIk639ikBjCQxxSYZKanm+qH2vfMwQtmd0sVUBtytdPRCAekv
C9/qI6bSHNQiplthBW/RiQQ/7I/avJsyoL1I8rZuPFMgt8d/sVHF0CSeNP/I8YMJCP2k/uLX6Py2
wLkXGrhEBjbWSbWWSYJsDyn70yxxfs71Cv3EyF39YedFF5yaAtwC/noQ4zCAc+hllDsUjqWiASzR
CyxnfiFKirq6R5jX9FoUVAYKf8LiVFyC80zm8ZOAt8FOD0fYDfLAey6MkwYpscF87qEWIAIdpvHo
eOoNKzE0BnpWmOwgFwryeZmx/4YbiUQBwdo1yoyMy9WeNLrwi9BuSuqS/t8sab1wgHsFnx7lJDfJ
vuuBhqZOQvdMKfHyr1EEjTUSKPpJ0N+TYDWpSGQ7lWAThjWXriYLLofaXrTM2vGZgkzIJp7WXdRj
Q4XN4N7KVjVnzsmOp7fYQPe5V5BHvNntQ9Hrjc8jA5J8G29OdLe/38qEepC6fEJM2jQt1mvM3pW5
u9ErGGldR85ajMl9nL8ohPuZRTexChaa88SvSOkhyeex4PVeRVgRfjlcZRJSf0QE/UDFIpC1rCQE
a/CD1U0aCu+d86rAbZ0MmqTGqvqSoSfUx/4L4CROhbF3nH8BQjVD34T/11VothZUPngYUiqMXuIn
mKAo6n9nm8+viw6v9ZQBIfv+XLyrKCXudAmGDBcsBoOI+sthAoWvei+4hXyCc+mkwIRg33fMeGTf
qU50VNrnkS0llE4dx0tQQyAq1rj6nFuYUHLRYmV5FtekBCfCf8zqbZpMve3WCJZdSEP5L10iIEhA
Jwuel2Kpm17NpW/T9uA+dyg3fQ1JxNhIig1f/BIhEt/giv1MOXVRlWrk9NnKv982rglzH1/Y9/oF
VaqRhyCNfC5XvVgYmud/Zj3R+Qz8MeDlConrJAMiAywSm29b+mLi7mjJNaalkbWZnBp0+1gSNcCS
bdySxd5HiwC/2wVj2xarfPAgsy1bBwpms8TzfMngL3glQupytWYDS7ub3fO17qYhZbGyB8BcI8s1
uk0h/iFBo+L7CbPsAmvZIbOmTF785nZ/7Iu2PHpnUIxpFD9fLHjOdttw+7mSwtLou5+KyZwH0SlX
Hz6bpzPR7Ovl9X+KcoZA6bPiP5XeQS/UuLgfk4fmAYaTXV8avpS0lt2RkgwMdXHv9kCWSczDUa2N
7Jx2ALB0CfcocoYayeBjPujtD+7sjxNtpL2fBk+XqdLJM22kADHTOwybAOZQLhMECf3bn4IS/gNv
mbTAjdQ6GhAmBpzYEj3YXfHmHESLB2h3WtVoH1rWVmYXYKdobl+/AAO6EHnXdsKYaXS3bBdhreQk
gLaMaLwlYO2gfk1G5KXQidyPodg3tiiDX7fc0Nnw6hB00M+JrdDNYbg+PVELtERT44YRK5ku/qPg
bIJrrWWx7nNmvAQ+TNmJ0/Ynuks8eqveTNAhHd/9mpf+OEZnOa+EVeajQ7oIB79hytVFITuKlcSd
pZpcnloGYNHYibPAUVWgdu563h9j/1F55XnoXlEDgxgp987606LQICNvZByvv4zlYFtHQMom/g0i
nXtd/k6uC48dy3Uss7OtCKbQclGlg3z1SFkCRAx6LP8NAzizPgcW2BZfC8gdxuSbIu7ddje1nFJb
ItZB5/BAVzpllx32Hg3+gaFKchw4GDowj9eyOmCtWGvY03/2zGzOxQyBS6vID59iS4gYjkV7zeu/
lk/nAtIuq0RyoG9B5nUK/jHnZ3GY14UxvWJzg7Lasyo8OE2UF70W/ntDYFwFJo691kbEaVQmM4FX
Q2gMx4KM555Zc9fLZUcvGX328W/lngyF0sXTWHtZFYc01M6zurURZ1HeG/HGzOR1Xy5si7e9d070
LqqaA5efkLv3z1W5qHk+2xvI0eIA4YpoLnUyY6Jux+dxRwty2E2Wy/j7isQYDpUkdlK1YHG90z7U
TD5t9cwsPzbNzEH5HgR2qHbXpex8iwvAMl8WRpNpyjgpO7gw50i3roN5YMIrGIFotj5A7Z3liZLr
7ATiFuj46szchggIExp7Tj2FplVvKFhQMIPTwzi1Tbxjb0GWoyisBJXNpUKm8pJK/PpSL7cgor1f
f2jvq1zbSOMMQIxmbmDctkeR/ldCEzMbmP37PgEMTV2PhlagTUw+AauAP9v+BE+DmeUby/n2wWIJ
41L3XSxKL1AgJe6a/kdlIlZ7D0zAcci3qbiUW1xm9j6YQYHE+fQDYK2gN8TvS1LxDbRvBy6shOUj
YDjYUiWsMTlKu71oiSxIj7J34vEll9D1tzKwuojPlpqiN+nGMT7BSYT4+7tTtiJsnFtFCGydS48S
uPGGaTawyI+zez2pYe3pTRJ3TjXFBP0btAYl4uNEPdiB+t7tckKHy584Obz3+L/1uYJG+MSEFBuc
vjKCWti0zY6VeLo2Pr+04ofaXqzCIRDIJBmM05pAx9DqfBdIk7aeYh1+SQkHWHSGTOAtDnJkO1UH
da6L5Ww3FCC6R50JvzKYPbppdTyaUWn8rguQ5HN7++y8HYxNojelF9UgxE6vndFd9PuPYXZuquqK
nSrZM9cR2w+KwxcHDfMZIMTxPIdscgG+uL58JI2d3lIE8fZ35cplxFawlSb356Hv3SKcZK/32URn
P0Y1YaczKG/8IEovVNtD64IPj/Mo3OJHHlbJuVMn/TQf3k3QAnPfVqTYajmhkxoZvqA/dz3iLTTy
hUvHPaDrhY2e+i+eI1kWLgI9u2hrShN8Z5J8SCC/KcjJMVGk4rjwUZ+KRG6CWjxR0R7XvQThKRr0
wGnYDnNuxlOwZSObVTdTvBhteNnalTRMbGUYlJPveZqHzfUs3MVN+9wxDkKv+ek9k8M/7eJZMAIs
FGFkdGyLXqaSe0aGmP08Dal1rrIuIB4YM8HeqUay9QA75PQwKSjNfQ4mxFCHPutYZUrJo1TUlnj5
ZnL0jm0mUoUfkXkjSI/UWMN5Ms1DHkYy2G7j/jLyWZGNhh3sGXVm/ZVlDm8yjtHF9ZzKk0TkgUAu
qaAg9MrnTbmoWG26ctztp1bNfH/XyLp/X96Q8nHvfEDF6L4NVAc5XhnooBYu06uCZ8metuKuRNCz
up2WEOaZsLjV2DOXOAkb0s0NLGOY46T04bsKyu05Q6GOJeyeXEln1fp5mY2CGI4GH05yz6Bsi027
eAyVXUgqHyeVA7vE/+He9WX5w+3dMlHK7YAzaXmx4ojcc1jmYiqpw2yqISiqpLIN6u4bYb7HiAqN
mMVWhrP9t3I4a9W4tZrGerBWo4vZ6N3NkSUzEtYdfmmq4LEPOk4WsdCyP/la0fMngmjNC7Fk8UnL
2YESayCivFYn6Ds0OybyCIfhzjxP5Gvxpgox6WbG+LDek1mtoAksPb10LqoNxWFO/GCWTFxkUXnV
nt03vZ71FLUilmT2ryiXCtJwCyxNwVqCVk4GHfvRVQ0k4M0uBSFfjJVhFNJFTBvVJCw7LkSfZiiR
2+gnjhKS5MmY23gCN+j1T7v0Jw5Ni6EnhC5zGNVqCiZqNMgeGySK8mT3t47WDSJbKPaffEkWouWk
r7D5zP7sWIExLKA/eoFoVyr2NVcHebip5bVWRaG29FfMulQkcYz5SAA21XLmf+9fH3+XVFGetPBQ
k8MF/4uFKU7udi/eN3hiNk7sCfzFs+vVO1R/0F5lzZrTVRW6+CSugCBbllYZC8MgpLuW1dicYJoH
CyNWqyk2jG8WneAhzwgaSIFR15coB+S9jonmkp+oM2CxCwVrWNOKRH5pGNx5gzgspp+SMhgeZHbU
cDNTCocAFnxvFR6bArOvX/WIJWQNX5vUl8rT+0fIlzYNa312i2K7G6Ro5ABH+h6z+yRz2dfeMcdB
E/x8HnYoONe33qDOaNK4MkOj6WCJHH4pv47sQw2cepVdDM1v+5VWL5zWaf3xIEG4g8rBz3K3NrCY
oFxHQFaOB5oI3DDgjHhOBsK7ax86jRSQyO90edEsFZO0jHSntpS1QL7Y+XACr9psc3fkceomBgt+
GRbsIfJy3XeRrbfzak8jVycf1aarwIH7u/xpIKYuX8/d+AUyARXIXnndyZOkPdaR5Owq8BDnU9rf
uBb/Q73H9yMq6+YNNRi51FAvcS1HJ67PdwOv39zrIkDA0KQqbhi9JWKU7X1XRVZf7wrQT7zCY2wV
Iq2B75WhtNqQ6RJ7ESDc/dN9SMXs1IPG5vxpTnPK/hVyY219P3Rc/Y4P7z0fAy4o8nHoSsdz1mSy
Ss80nqmkn9eAx7SuLiK+OByeLG43KT8/lhsEBfbJeff7VZ23U5DkAUuqCMrV6Fd6AAcYKDA3U9u+
bgYoPL5y95TSGxJpDlMwR3p/dcITcQcEgUIPhdp/TjFFwTSSJnayjVOxFr/PeD4bCU99su3bPPlM
j54AzOwPwebedFmffUn0QzUMG76JVn2bsm4adBiNpYUSPCISKHSEMTjnVZ/34xe8WKXXBpAJoPRr
FPj0/pIyoea3b64/mRwbVfUaUVOyg359NOfkLPJOWxJBRkZfjLKd1N0gmSTQiCG5azkg3PideDQC
uf8ya5h3opqbsJk1DPJD3jRgd9Gu9ks+i4RK6rDZAxgX6faHM5kLDZghRGDpcUSa8y0jUMpIf1gI
jPuWJcmmU/zvb8/9fk75lakMsKstonTIvQU6bBnCqX/mtAEoHL79wvshhxKy9jBY+ADpgv3x6tYF
gsjLRFlbUgIguylBDo9Tm13/Wy+U6iqQLkIY5/ypUkf+HKMcasvCYTDFM6arhTOfbK1ph8IFTcxP
tojbZsuovKyMNZnVNyIwaAkQ15cArQ842qBriioUmHW39h81z2XJ9C6TlQzzWqTv36zDbHChZGVd
Zoya9iINNemMLg6K3jB1sB1vylYO5FXqXQHoqnrrgwt3OTPlzDlLYlnEs9icmfP+oAvKPifC0Gg4
bDJDVaHgIK+mRmj/a2L8UeGQmxlEuWeXzbOW5LClm8EdZ4H6gcQ1qSUlEl4FNmG6QcVjQBn/mS/V
TKMHSgwsvu/QMf19l67Vj+BFN+Lw4zMoqrIdeb4NXAli5Q9gTQMLTIQoX5TySG7YcqMm1Rr9ISpH
swSoeIyqwr7gZNCP3rA2WMrfRblylA1caCLA0ay3aSz3gLgEdPKCHRS34yswoc7ToRm0I8snXqB6
QFBEI10A+t6NaPYRYrjaY5MSNO5kh0EwGphIdN3N8jw/ukyFr1E0C668U9iH3rgaSq4wa6aosoLS
fUGK9R+McuNd4HCLCra7wXCrzepvQ0aj8CTSIGnotSgJUG0AVtWCqrxpg3zq7K4hp8uXETUrE24r
TkZytl+mARVFYXWrhA3kq4crbrAfhL0oLFwVTJ6fyR2iqz777+G+Pw968mjtCUX6fEDSHa4L9XZ0
WI3eZw5M196BLRj+GXnUuE1ffsksfpWaWBZF1xeaJkI29NQA1i42ZZRW5fdT9JzWnd07Oh4gE17A
8mUjt7ilyCvvuyoKskX/rNoL655mCwpPqgkqJYn8AbFE2XGD6NmYtuCyiCbdnJLZzfgMnoO1AjSc
55vlVa6ZT1t4UJqNnViK1eWkiaDmZrAFtqInwkvYD0EjRGpDDZjZe/tQAfGj/Tf1pe6E/EgcHKpX
0OPzDZvmbp5lrXYzls0wMItYVYWTqF0YDby8Lu+SAkZQBzAfoAIiaw/V8OmLHg9RRoAmzZlk2eJ4
r/3+NeConHloCk+wHOT72tLn2uFEsJd0D6+Cr/2vgO8sawys0xbwG7FtGy8FLvftD2ERaLLnVGRq
f+O/Kh0PdJ7rdsQw8kMS0vwnTiANJ5jIKiujxhRwzyza9dWUaJ7L0Ux9kFcOKMEY/aWVB4ypZ/8M
HcVoPUfi/G+K36VWHtCLg7H2O5TrybOIfX2ddjVtnILzwfOPKtQtUPTmdLTjhZwJLZK3fd5Rwiud
m6I7vBlcijLKRezMeUtf5ABhL27nKRzJ9bu9RVf5wBZliJCm/3qsORPZhkdM+AYnhxEVfJUh+6AT
/qupehzOIcUdHz955j1SEeTHUZKVTog9A+83I3SF5kjUUZbpDRNVeV9biq7LN9qDdMCp/6zfcBHo
XSmk7Fq65kC4xrVtzx5HwSoqK2JxmyiY0u4vUnJsKyU41Y7i8cPGixxgVH1G4qLh+mkGhp9AXL5X
zq4GcjDZvAzyj1zuTZD0QK0gEqnytYn5UmoDsLXPu0cQ7+dta/4BIuju2P5CovVlgFRPROzzL9cV
aWmuGUa85ZZvlXTxWpVJzkkHni71DHY89GwL7igJ3eCq3KxhA/OApjUrIUdx+E9GGLJPfNuG5UXN
gmPzBZ55gOd7K8eLSpsLZe3xzljG84IXhGrytS+f2L+yVDmx+bcCyoJPw6tf0jk6hXeYZCb4LjMm
9apK2XlgDNiDJYK8GGj4PM38CLNwvd15BwTdqGiEvdIB6y/bSPkPMKYMCKGghDqmEW+f5FAr1GIS
RzRGJeBm560aWM1z8I5dGekDOzo9ScAlVgYTeL2DGTK99Wr0YOlRvvlY6u7UVPHmoe0ZcRCSrosA
2EGSErpFOUbIlK+nE7Tg0XWmieIbvKwgf7Bxc+k9/IfV5Pgo2Yckout3vh6xUk79hTEuUPhq7uzA
G54+GsxP50Gx8X/whh9tMjjCVAc7a20RVVtB4Ax2pgaSkKSKyGsgNAuP4syNSqulMr+rc0W7tsFJ
nQy9Pci6sn6RWsod6IqrdJ8UQtFlJ2w3rHfB0GRc4+e796QyQMQg5PnaYsj7NSdfT5IQ7S1hoW4h
h8pP0qeRxLXYTxY0vKPKU/qPFlTV1qEkKR5Zp3+D6lSTGLSo3KhJhEWFvmR+XG5thgJejDAyczd5
Pxe7lhRpvwuKNUb21N9t2yXLf4diRiWPbM3j2XFO48Yw59sRHw6RyRzLHSQ05DUxzryremqINkIt
vRRFeSKnob8ectOHu0tKEs0tKoqN+JR5Y5+QrCRPHrGE5+28GVEiihlmdJfZk5teRK8EzbYYKcqF
DC+PAYoiT38ZDEeSu4hM5q5F7y8tP6cjOx8cTfP+9qO4S9Eov7KAhIaH8aQvA4e1lBAPGdp8wxyk
JVKayrjhbuUR/7tjUwPJtLAJiukK5LK0umOAR0HhTTGxTVjLJY4znH0xELNajbw8fYfdTx1mc7u/
X/KacJxLTkNXVf7Yh31Zx1E/F+JLJezLnFh2pCoS8FnaECJr8+Je0HWQSe1Hx7SbCU3nLtA8FZoM
ojlciyKTS33Fpv1aEcz/31L1hJ2nCMb/tLugbxHVTg6h27ihdJ0RBak9K60aO2G6MT0aQrh9YJEW
bOoBKBpMgyV7W6o0TiVIRfaarQhQt6jrwJ6TCTNV9+Vj3EhI6Wa2NE31bcNvSuqRHeZoI2KwVowa
JzUVB+799BT/LUiMjrmcLGtNWfwW84Ro8MCbHqGUZFgjM5g+/DAGtSg7Wn5kCy7WaVPlS9E6gdCX
ozXrUkOwpWli6/pBowqyARaelzMXf0VmuUcrKRis40D6Hx4SZ15SwH6Bf2WtoA8B3Z81+xsM3798
tl29QtTXc1Cn+sJohGCPmlVB/J/Z/V0LR4ZN21CrkYA6o82D49pyzYwPL8rjhjUAzqiV7x6b+M7e
AykbHWlIsNCFW7SGAl1nvVxrW/gFm5Pg5+g98DigqDH3SNvh4jXBLBepYtbWjOlt93+nboTAyqTF
/S+va8OvyPhS3vD1pBAzjjEDsNxy4yq59OE2sRlx4uwKgWDcq0EQw22s4C98odL7srDPLlxB3gmg
2y5gPpHN/gpnCzkVfyNNG1bKTs8SKOeTQvRth6P+kC/+ijQW8R5ThKWKQ6846W8OaAWDRa4Zxlso
bpmEKC2rB/Gx1LuO3z0/LsANChatA/nk3njIUBOTPJREnO25MEPGot4KgrGrRD7Qi0lN7ifrITd4
GfJCrsPrlc0a4H1JkxDk4Jl1MQxCPqg2AIJN4olFSqYv3f5FlsHsv/PDmdPc8c+d/lR4qB5USiCY
RQjKtm7+bHeb52h2YDrst+IZOmdLNsQy2PNgcgAv5ZUQerpW0e5Cyf1EBD3BSge8o3uW+XXogCzJ
zibGHgLtGoyhjcqbLp5ELFBdJPdhyHezDDKEjCmRk9u+MpJ5tdR6cUP6NTbSflVos6FFo8dZxr2z
/I+QQLtfirFhAJ2fBzHMn7s3eqQWJkBqgMaBqpdBm7XU0SunAitjLzngUGWHRC4CpQg7EidnUV8W
BX3kGvVyIpgPczac1NwTQNrxxyuTiN+iMJwD+mSFujZ/Nlgx6AvBgzSr/3x3cawYUJdmDw18c/E9
i3r4FH3LkT80oejC0drehiwkLZHvyu0A9JlAM3utH2aKVmTeCXEZxYVS82qRyKKzbdbrWld0+kcm
NSZBvVN8VImYtvS2dJpOaVMDN8T1zxPTg8UEiILxur7d3bs139BUC2OBgrlZVlDIw+CwGoAuJNSk
gpay8NfKfeBnqXiWnHBE67ueTNFkwksVzj9XOBesYlL/TIyfmE/Z7VhfA57U2Lyzu1fv4U86f/gW
HOd9t5VZ9sjFZkAqcKUhp3qjC5a4ztU4eIIcdkeKK2gWCoK6h8OGHkxaxqc7EdnQucfJaWyY3xiR
1/svs3GKxqsw54uCNZhQpwkOwwINEIf7f8psOPAfYdAQWLoYQs1hvRpppBVmqabeQ648T02iWTkz
KHEkkA23M2FhCGiB7AU9cKubvFR28qYnSpgbfkBScljOOt9mMQ3G7oUgrjBJn3ghkJjPRKrnNeHQ
mjnep1qU8bAC9njqkYhCDgwQQj8yMBvN6ObWyK7hZPYr9jsEjMg0heN+dlq3+O9Y7HH2QPDZa+Am
9oEoEFTACtyhpv5wVx7U0yP4jAKXSqgIzqCji7NTcaRCRB2DoNuLoCWXzdKo28CgK6/Ndzw0WvWN
1IY8zdTfjElypRwc7v2+BkpLdPzBCIdg5r/h1FWXeLAV9feScovpgxR7n1Zxxjv1Jptt7ZwT5bo1
9URYh47/MNXatxWrn0KLs5WbmY4nPal4FuhyPcc+WaoMv2C4KDhyUx+xeu8MLuGsRxaeZCWB5Kgw
QeBh+EhYgPOwGvBGAe8emoA/EW+oSJo1YEYmtSoeB8/NPSxUQAg6+J5btVCbzKMW+fqk6EOevTFx
MT9vs6oc7WvGANWAWtD/PqIWdfFUgJ976yXCACX2wdSZI6kLmWuid+03ahJowp0Dl86n94lVLvXN
Co96MZJoQXQ7Z5RMVOdJDavlwX1EkUx3JtzQI+D4pCMTFn0S+xu4ZwN4I6/r3ZhK2ah2LGrdmTgV
ffDU3AwEkXFaknMVkfRPWy9LohWKquIF9BhjIuhqk2XUkz3rBpK9fQT0UD5/MtWA/3WlaGPzK5Zl
4RzSvH62924BJSHKLlzIyLcLTa2hoEnzY95blkPx4JSBs+hJ4Kwdi89F47VFQlUYLJ1jMS5lesbF
Og/fNqSsE1APONoo3w+uKejzieWtXwkGQ5yI8YivczNfAFVMZf0pIJ0Z1sui62Diyk6eL3oftJr5
OeDI55WzWBiij2BhFT7qkqAjkft7Nm5OlYy8unHuuk2j+GCVefthyDBKU6d4JVTdl/GWPkyLCTBH
pmIhKaA0LrJ+fe2w1iuVaKl22Up8ia+N2SnSfSg2rF8QGRYavtgNrvlscJfjsB2dGkYuBqObqgWk
/RH12hCH6NQZnxXwezE4SHtgpo5mOo8zgn3PZIBU49wyrni1ZOWfFBst4IWsnkoUUrg8Hq98TBRw
pZaGBCPchHPgk1G229ZbWzmQguSPYqcbb+lih18t+7arWPZVJgNwu6A8Cz5V/wVKJak3yL5S7BsN
MWSk0ok/7SvwR9dXJYCpzaPy11cLaMstL9DM0of5TbbcRLZY4jK8p8zFGxuu7g5SfhwZOf4cgYwD
HECeQ2TlTVqLkZw5VvyvYQFpFCkgbVxEGJKsWFeS/+YYguCgEQNcpPYAUL60BzGjiAzDAr5wNy38
I/Si80k+ovpiaWiLED5NH1nTTlNJMoHr7W0rzvBCA8UgVAiaR/mTGB56DpEFY/3bi4VydhRpkK/G
3zaKM22OZVB0Sj7u2aZTfwl6Cl0QUu7ee7pJjtyRaKHIoq6I44Xxs/vjLzojgSHeb1GBTNERvfRh
nKUwKcmfAqBO4N1OqR+x1lbzkC+RH5MucV8KU3Od2LcwSXiyS/sNmwpXG4D9j6uuf+fRBhu/foAb
lO1Vb1m2GQaagkVLGuO3l1xcWYJJheacXbRQjsGqoST4ZgaIzKhNToVPAn508CiC8cV2yxlgPL4n
mXlwCr+nEFc3T/MO/n+oSe3RKINTcH118BEUOUlag6nXR98Xe0Zospa42kC6ng56BeUXxX7fcV0W
7JUHeoJ7KNWkI8DBYGXwUKTF3vG1CRgCTTr/3lWcGnFQu4Li7F+IBd00X238JsudB94J2LvQ7N/P
u8W0pan7FJr4hyygxZyUFPCeHqKdmlxkPVOdg1C3XHYcUgRSEeYGpwHjrTnM2ed0RG3gHvtpXqQM
BDd2pAziXWeMSxCNt99161hYk+EB7WW1qhpP6KqpTO5SwN/a4fmWP3Y0Bt69JNA6WJSF109wN/7W
PiTU1gMpXpWZJMIkNeJbEKB7HhzFV9QAIhpODxScwWuxb5E8t69Mzy+xooHdjHLKxON2BORxYfDL
NxIoMflayNA6Q4XVsHvLF+BuqHkhVGP2ru41HhNPbhYhtgjg3WgzMsdExu14B1bhSw+8vZX2iu/K
MJnMpjtSVo8CDhNEILX+/Y2BZupsP+vMKH6DwO1DyNkwyOS5PJMBYjoFh29utJ5WX/wyc52i47vM
Bsojc8WMN1jP4D4Yb5DHEavMo/F+typ7rUUcJpTLzNoyU6c+zlFzF1EtcdkUXx69excNrbXNJau3
hlm78AtZSbHVqv37Bst2qLOOiXFLGtjCFO4AYR9Xp2uRkBFi3RWh9AlpiAqf29bdSj5y6KYygE5D
XPAzQQdHlfuXmMBCFy+R62nDjM73YpW2EJY/MzP8oah1RHHF1KY69Nj4JNWfFy5KupzmYhCWbQuK
WTDYwmhr6cbHyU7JWjo7z49aBqHAEmknS2MYRbMjrbdyhZRBDrLeQLsu+vTYT72bNoq3zH91Esl8
TvGg0zOC4p2W2BKFwrs4bKdqbRnDzpAr+OmxwW2U3DygrgW9MPfSZ0kk83Z0/jszmtCrL5KMs2bP
4BNQiIydTmXlQj4jKozmDfc5DbO50FWY0zeprDzvoGe8xEK1X7u9WRg4nBV+mRVqv+xVP1Ax/q3S
OoiqYE54s8GVvhb5Gesg4GGuzgn1pqd0yfJh+zMtCQhYQanburVJD+SZKkad2Y2kObWCuWZz9HJk
drQjUBFcHowUQtBWBlXNtYcWXr+4TokUIbZ0VpWRi4vjBT7rdzyDHcm4ycqnh9F/ow6xyfDKgk/L
zyT8kxLbCSa3Cn5NtRW5eLwHt4hK4tysdFukG4asDrPembPDwyePfrmFqJ+f1hQhfzDCTf2HN8+A
1e62m6EXP1cY7UksSLC412savjvS7eeDJvJENy+H/6cos5B7qhZ3nBt5vx2OENgvdY1Y/FIHR1fK
wJJMKMuCn6G95U8B6zA2D+wRldwCNM2zvLGHetZ4JNciVTxZMRTJEx+9hsR6CF4KzBi5r6TCdryv
bF9f834Iqg4uskScRaOjplN4U3IpqszxpcoK4xVf2B8+IOAHSrIduh6LcVYH7mBNoe7VioFpjSC3
XjM1+wevlDzfSN9t3wVm9Bf29TgC7jkbVGZuc3wmmdTW3nuoJ+F9ajPbHxhepBBYD4O4IwaHy7wT
tY6GhqthLpvbdUK6lIe0DrRXQtfHUalnlxeQEFL8P+1UD400Tt1Exefpj69MkpY0GZQ20gtfRZ9K
D9Mwdoxp+z6wz6xyaQUCHlnrcAB7moN+cbawzSpdHjoOgmuPawnyqu2Jl+RPorIaXL4/viZVnXdg
w/3A+Qx11Ud9z1mmxU/LDHyZNpDaGhWQYOH6/O9rSj8KVM4d6FU8LmLZ2A/nGfzMUEDoYMahM13a
PpdqZ755V2XsI0zuh10k0FZKWuVLDfanGQ9IGKsgRAjgewJvDQAoAD0u8lstLKUk3k1/Gi1AnbVt
Ztf6PbVP/39RaNzsb0algs6GygtbHlwIW796XuCbtSrUNQBTO1QTIVeF/VAozK8mdeYvPlYIv2K0
5k6VMIZnNoLdLUA6SyDEg5EuHFf1ZxYW8B8BF1lZocrGFiOvNwe7QLFBzEwYpvGkVg5WEPMuxRaR
E/ovggX4DdOp0hyzIffxpfa0669UjvwXs8NT0v44pM9e+DBJQxPrSOqzLUYQjnhR3VJotLpkZpHr
4rbPvZR2pL6H9jJl286j5FFqtoEHuzTrlC7KHYcVFDc+fkgV79VeI/R5obeIzLI3d/Uv3/3JquSZ
o96ptU3+vmndXa55dhCPfjYxk3Jh8ZJKHztH366pBj2BZ3dm+u0mA6sENqoBYKrwdyCUWtE2g/x7
KVH0NEVBhd3ZTLyX9SzhGqpZXruVA/9mJJ90N67IxM1wa8bXwSwVOf/YGYacwkOLP7pG/sdrJtv+
M7VfCnn8SB5zPWUeGZFV2KvdXu2/fXiznHXIFK9AoY3Ap7QlNLr8174+WN6UhyGyiC/1E4+yD9Ig
BVDv67JUxd49H1Vqvxjv0b5OzIrGhdcMKdvcPwkHV+j/N3B+fe34yD0rKf2tY/o8KWbjLIOSGPAk
Y3VrOAqskscAwSWeZjzgTtQ2EdvWQspM7OYR1+FoVw3+XHx3dgzSgQc6f9CuRazyp6w2S5jZYYH8
nImmds/WRhH+hTKzWjBhXjxT2qVaVkF41OmFu6wTMaPZDalSk9eU21NMkaZuDuUBBfR94HkyUg5D
r60hSUC1wNohOqhFlWRLXGJGI9OmHh9Ix7jvqGHUJRujzvjHuPvXOLUYkqzyEQfyvHfcSgZ7L/2q
rWWR9zzwsiAULSzgQtOXRLxEXwGeyVNIy6OEvU6Y2xaeIGvN6RB0c6Hfd28HT2lCCFPXp8yOwzy7
Q53jYg55aYHmGmtmzo7Dd2AabRcUa3zGvuWsMqeMZMtlON76rLaH1xSHcebHAhIhYMITEmL4Qc7k
c0cP6dIfhF7JDrCghRP+iYVkqsN7CjSG2wkU7M37UpsUm6+0t9z5ofrLXyt9VetD0Kcmqm/6ilmM
AgXYRgD6G/VlNK4Ymn4GKVNEmJTkkPPJUA5AsigBxKwDVhA/OidEcbI6ouSM9OGg8neD1HknxO/n
ibbLrRcWA6fD/XK5YkgmVs39NvxOG3d1yhFPUwSkPPVLKkYg6uRnZo1vPF8vFaf93xHUxYWGAGxE
nrAwvx/vHVRttK9g5Ezwsr9qBEPdHVxBGmlXm3cs1FNlfAaTzP03ew9YRsW7Yc6Ecnh2y1O1NbYW
2+AEuZ9M6qVk8LBfkzNxjIdDr8I0DaFOXDwTbywlTuqxverdJlcF4mxm8OWUArYoxhGn7NYnxJtG
69TeNPDcI5Bg/WMN5stebWIi1ymJ53buIkxK47Zs3ND9Z9a7RkcPM/Dldpj8anWEV0xGTFcqauIP
PRLqz9Q1ZXQ09SALavQqa9FbapUB7m9g+yhZCsT7MsxxszCiG8sClU0anbSWFA8Zx7Qyvad4r6A/
H06N2JTT5Ts+DXvihMkedlFDsBjE4J6NXFdcm7zhKYJn08kvc5F0EjRd1WJ1aownM3nHH7WtkJMz
nNW1/DIBbhZpIs6ykPfq3nW8aAbcTD8LeZr1EC3a4aA2IdisETWT1eo3gEYgw/GmWHp/0U8tGbro
kzbWz47UMeYkRFzU8YlbYVTF9s7AHsoikJGiR5TSBDZE40D7KuxRUOhHZ0bK7l4TtQ6wwRrutLPH
vSzCJY3jNUoKNMSpWuS+3WNxPHTgc7E+6Rc+gQUKi1Zam7g9qmBVTlRSBEaegU2vAj4/Iu+XMG2S
71cjlJAx2v+s2LDOZE5JZ2NjhV9sKtnZvsT5URtBrIFYxMfkhVdFzZz6Ebqf/2fw9E7YFMF7R7jl
ppL9lRNaKMuY23QLHSsA4tcTCGdW72CEqWd/pSojGgK2una2fG3mEz/XRjJFdzCuCz27WaPd/pHX
4fU+RJHaFTfmRh1KwEmDbtKa20ICED3rfR6JdKeNn0f5hAhyIuqiauD0KA7a0DYARnDARhg/MMSF
AJI9JfSfMycLKfowrZD+nhIGo8jUxhXWfRHE3CRA+sLUDusvxzr4QTTp90uSKMdHZYnZg6VRFJYD
FzMoYLIbBctQ/aHd2Hi0MaCl1MszZwknoB+4AHQAUsgRti//Qh07+H79hNM5rUxNI7Ce8Aib3pk/
lS1ebdZ7g3DXKz+YwLKFWpeweJPpVV246AMam3SmXsGvEeit6eZMd8xmNMU3SdIsanOvPLdp/qtO
4Y26QRp16JZP4MH4tbDsRPVWllQjOgbzylY5UHNOlaXT8BZf85Dyy0sWLG9Qg4KNLUNYdL+zY+zq
YrQBl80ovyFHfxGfcJBhFyf0zSQpliI+hpKJwzJoyXOUiza2EPdmD8chzOzQyH/PMLdnteGpnD+o
SqTEeXR0cuQsiR0r8fKNVNEI28IqfC00aonLY1YUAOtRa3Voe63bKCnCd2pnvG+td7/BOkxBSmRS
kQPFWVCwdBpEANSP6kDsXuS+fOz4v5ym1d6Fay1VTn6g5s7jC9VRowbrMNZczB3IgD3E2GXoxdxU
UgVfbWYtmuviojCLGU5535YxAUbFGWui3H33TGjTWXxFLtj1F57xnsqo8tlel/f1PZmX4bhLr6NY
O9VvGYu7PwMZafuVOubzc8DzVuhc/N1f5WH8SsU68BBlk1YngYqdKBcgporyGNbrhGHKpgfW3ZhJ
h+jyAI/v+fdRJzabOshEMUfOGsjylcXRK/0y5zST1XBsW+IDmWiDqkn0Ic8no3TK8si6tBy+F4ye
WtBk4CwEaJRg1Ml2z2JnSqcrV/BWhSQIIuovUm1QXc+zP7MRLzybQshBVJzzOVFG2IkvjLO+SeMa
rrDf/S0oG++Eizb4+KA8sYhWBNA3K/BLXMeOswb7nb8aAEx+efBxcIAFREdJdVf+S50LyU8QCiRz
me0WlL6JDUh7Rvz/PfRY8yq66HeBafUODxCPImzKyVyHUcJNkAyw7pCu4RBBNU+6NzQtY6hC5rh8
QuQVTlDTWk4ociQFjnmrB0bNzo/YvOkBTvIN24KXPU3VZgpU/E1RYKv70NpPJnNJ3MO/gZmQCuCB
JSUbbeBXW5sHXB35RpyZQkKHCStmUBAZxi/xS9LXP8y7s9+XFj4tX6Q5phQUy7cwCnTczy0LKDOA
uV/6GgOTCW/KT1lH58BwEkgOY91TnSOaUnCHTcFyJTleFR+Vzy7TUMS3I+BdqYxL7/WDYywBZR0X
S5NgzeZykggy54AAAsldjUt8SnjnmSkRxs7+bfjk6XsRwypyIVFjKNRL1RaFY0IFIwWn2RVZGTA9
7qI4E4Pkz/pnLE6R14GOl4weP3W/32ZuBorzK9ksYzA9OHaWqhf0c1mIe+/ZbusOorrKajBg0foF
KE5VM/Ila/tkj+4DN4Ez4VSGnr+EOsI6Q+rjrweERE3dz3m5pvhm0wqNQAI8fqvtMKVQspYSKbB0
mUp/28UNsDHRAae9w8z9gTiscXTPO/ShQQNL3yGDmPrEWAcyOysPIrQ5eOlxoANi+7nP06uHtYnD
j0bkXsO4DFfmPJA4m/o2642HFgcnKWqIpjXumNcZv57/3gZ64UqgBhTrTVYCgVsHIQIcxPZ7sfJ2
eckbRPc6Nhf6xAUB8e2aSrH2VgW1zCXITztincXj3HU3X0Z4JvioNdGmXkpwEDpfr7oBm25dzZSd
cQK9OQtkgOb3i8tAaxspgaNwbg52JMtoqtBSNLGzsLHBw0LchrQhOoXextAwwRZdC9S80OkFW9PE
erKOYwLAjYaOQE0UrW50NiAUoHVX+j7f/w+EE57wq0Mjvq3/9gclDQK1/ZWnoCbQJK9qFH8KE5cA
nTqG5QA5uC3qg+AgvJRyPRWxexW9JO8EWH2NYigC+i1VC3LqnvVW+LzlWZFfQSo7DXx7Qzdjd7hm
uTMKYSvxljq2ambOmhZ04lEisGunpjt2twLzo1ELHiWv7iuzmeRYddKdkcir5c/0aqdyRSX5QlIE
p3Diazq9QSxmZky85zgb7FQOoGaU04OAuCCc3mA+JqsSqE0RaWKYCz+bFtyHwkR6PZd8pW8N90u6
dEZyPBgPB1U8Js/HPsE4AlKzxj3cZVjMT86RAbDSgG1EXwui9EIj0SQ//tyV8vocwGuVYCU612YN
nE7krDpMhCtwg8r2mc24Ei+2UCxvvMyKVydfk5bUBc9OtMsENQXNmCd7ubH1Rgt4HHeXOyrwacWC
yHLuNdbYAgnTFzDRpqWppmS9jPQjJ9Fbqv8gjblnhLqkFA70OLqIlWtqK7gr/klx/ItOItLc+tzq
ve5ma6drHEWYC/DwIPxmAWw5VT/pWGaaRcdRSUQKdcDvn6uXvwXQFAycnjWQh6lFb3mO4jFUN+Au
Agf6ulgI1EO1anuhx+cyCkyUmPIb4SN/ctGMBmlr5an5G1XjAPdNjUDosxhdJ6eIpXhzijbJusIQ
9zqrRTpGsgu3+ZrIUUkYVDaYkBNCp7DrqwaHJHlM1yEskXsP5ZYujvUtH3Fk8RhzhmJFK2xm9Ak3
qR1Cl55CMgQ0ju67bVHn8QTfcnwhFJcxvMWMGdW+5BUD/JNA4GUqZZKWiCU+pd/GvO1RgzLcnuRM
LFB/Qt4l1vlh0X0/2vEHnYTYbcwxvy9/XcyszppRi418NL3nfMEUGpsxIKH+8WXFZKLCfaStwjWD
Se5kIjKxFMghePM4PK67K5RVXk8iCh5asysYWh+A/GffJSELwWluYCtlZFt4uWzAxI+YBUrkhMXg
NnXY1sMw0knbb/b5M6TOZYx1FI8RX29XL7rRL8gHy3qqxE6lvVGiet127BmWN1CskX6oRTJdNX9D
o0Dt6iKd3Sz21lzoNT+YETWVEzfimC4/WnpXerheDrXbQw9b5zQ48r8ir5rNrV79fzYuhj++Rp8E
rLVbOJKe35/ZKPbtZI0KLQyey32vgJABhWpJRPig9u8Hs+yUjBB9Xvhrz/YG2o3IOU3foMxe0pjo
Sa4mm169MmiQd3jpS85gYPA3+w/Qe85URDrg0EcvB6uYu0n1D7FkMASBUdHdS8+Josy4P/XEwpC1
pFaYjSnqUDydiqcTNI5z3cjtuXfJK9WJWoKIFCh7M9/DFUgnWmGdk1OfdXy6RdDBc0Ehm/OWOgmz
YHxnPK2gaHvFgGGd1PzZ3jGLvfKxCLziSHaYsmIfjUR74EgQhxwJlzWPjV4b/PGGCwdLMyUDR27i
dd3PProZfG9c9OGGiTyIDcQPnP404DT1Azbm5LQxrCXndEzuZGupHvUMHZ14SATdoTxSXLHHBdB1
rwGXi9NiJLTsD8WvpoHkBcrGh+IgI1lefwnA5NS10oZdNpKWrHBf4Aeaen+cI2dg/aBl8pcBO6YL
mZazH5vqC1AfsjDAJsYBUax/8qPeRkzqE6wIasjFVdZV9DSvZNyjzTzHa5ylnxX7WkXj2WE8BN0e
RTBbQTIwF3T17QJPtgTSiBxh3y9bNstyCROQOJIVq83fae8XmJyogqA06xF0fKsOE/eSScpjLka3
/W2DR2wPZspEf8OWZVm84zRQ5ZSt8EPSfMCyhZaAZpjhph9x28nUUp67mFajPmlE919PpH9qk/MF
51YINFDXdzqZyfdc9WuVoEbWl2sIPlt0/gjPZQWZAQm6F814bmABFy2FyudXSdOHJXG1sFIevZUG
0BugE+THOPJbp7yRz4gITjLQ+XSfz6m7Qifo6rwQLs+cY4Di6GD5SuVUbg2hwtUdC7wEQGODCF+A
gRYnJNVcNVccHc/WUxq9dxm9Mu3+/Uv24XNT2TH22f9J0hzQdpNHQ9Gm1wzvaEJnSCDxxx6w6cbJ
lfPvxYm5l1gPzIIeeQP1jpoLFst8qb3VRzmp98/GQ0m2rPgKHSXNrI+k+AIgz4KvmvvaGJo75AJ/
RWeloNmUL5VstQmCos3epxbnz9En7OMziQ+XY5v4zMz4ib2rLvWujg3mqGQYTlIexP3h5zPpk9eh
G+VGdJjsgl50mWSCgNj18pjLNH8Is3PUu+TRZCHr3raihWwZ2yrI/UADMIvOJU7I5hG7JXqXzs0F
tljjbWRuAWIZFwC/Ncay3KM/HfyyVE1E3ksELr8f4iDw7khq7/Yse+ahxLqL6GB3UVBE/v6QtYlQ
4oeVM5d1rn1XK8MNOrboPYVJjD/Svbf+bu6ffel5ru/dEeRp+0R07nGEopwo/UeWeGzhRiwU9xDO
NOKazQMMyQMZPhidxz0r5SAAtESthacLOPyDUYjiCgrMRaYlQF+EnGt7XEgkFacBtBtAanKm9WOA
B1Ab//2jA5Z1/jLM+pI3RqCnqVQlx3sWtLnmmXSlekLX1fWq0N11ieLebnk8p4aLtxg/6IuhOa9E
1ZEHWlx5RocjmLgUTqLaa4S5vl9pl5uOxGYKrAKdu13JtKVURzjL9P32FxtTF+UJmIuSdH2jmYdX
vAOuHP2lCUJYnK8eUwqNsLmTZ/kLgyDFZynsu9uNsz/f/yhh011GA1/LV1RdpWo67s6yTEH+8hrx
TZ+G+2EXIP5iVkxHLiCoZPZZ+/wFT6FXZja9pNMlOHpXQFWf9Si1yrIPl+SSTlgTXmdPaE9CqIhk
bXQMogd+ijVntiSdjayVyzIvsYe95NyiN68HJISdbk5BxfA2ZJntv079XWD7VZNwW1vx96HE2q8s
jz3hwn5sCkPPz7yJnu/V9rA6aBbXFn6p67wpbw6bzdtuhIk/upqYsxFPAQGs1RTwUaNc/p4VhYtL
5tdXq/8nc6FgPFXcklZR5b+61qjhBSVHp1QeemGoSNsy0oUe8112gG8tXaqNddR2bUM2o7elUN/w
sFVHyrqVAJp19a5vyMt8jCmeyp3MJkFjpx6BrpwDNB8FfaIcTH1kVYFPQOUwApaXGxJ9MFCbwkns
jhDlyEXyeI9aFfbNdA6JYPsBeFCwWW1FD0v8paVufwAolUPDNG5QDc0FQ7WT18F6QhH0Tym/Cl6z
PZy4lWaz+wLnnqvpnQnQ9xvo80nfwse3zmIDouVy9MKVi6TQySPfFvk6+W2oE0GelvyYQeBVOUqf
izxqbsmecW8oKvlCCDg6sUOfeFjqKjio4VKwlMW3ziEzETl7M8M8Qi81JFEQZ19pk1aCzRuxmTL4
w4zGz+xuWZFBCIH9hPIq7dciLchp3rzVeJ1E+0+WFt6j4T43Xq/9dTPRObbwDihqWX7KqnahLsgF
JraFQNwlvMuUmXJaRI8tY9gdAjQBQVjcdJW5NJUS9BGVqkWtG8aIV4wPTY6f9rRT8U/FXOoNUIva
dMLlchUBmozfspB5Zp3ReB6rPFR9uFnMOJYyUXLdwo4V5TiVu1kNLwfkoDOR0vNOT2aKfab3D/UJ
NtVqcsmARGKacbEJxOYEJsfAw0Pb/KUc39MQS/h2CH675trporZrrlzYNO36zaJ/fZfFLecHVV0X
2/yifqECDyry9zKctqBp41WMwwUMur5bRD+VgouJ9u1McNEcZ1j9rBF1X0iNfsl0CSBlByLaasHq
oU+ELv0IecQ2lRB120q7bKLnn2xTbiLqWanGfutTZs0SiNb4MMStbtDRL66ZAk+X6eUrG1feoa9K
QJd6yOVLHRehm0ExoElv5Jx7LTSXXZS4QjMq4AWBSuKviwV+yg/3WI+zedv+OjX/AtyvNT+GW6ry
tc16o6TjZR396eOim1DN8VmbGHKZ+kmSOYjiAIrScTz2SJCIJrC2ZWv8qSYDiKlVhEjW0rtYcuN3
3tzdniRji7LJCd956O1q8R4tjf/MCOxlZ5zGQrgtugDLTg1iKGUoFmaR1v8XwzT1T451XX2zLxSR
+zcYlxYesgjHbKT9gh236cY/RH/KKvGEeRCqfILrqU7eQZ0COj+XP5C2ulm1Tee1FyiicK5L96OM
PCMnb2YHkszTwVGWQB3g+OUlBmDcfK0VyFek8/zblMxwMP5gBXxTMtc1YYLCRj5YabA5Q2oRNEwt
mB9JSsKD0F9ylzVT4HVNWWfxwg5afAFTlGjiuLTsZY8i0inMJqeeG+twjbIfSv5akEEo11fZqBlN
OZ/4v54wlIbJ2cHXnb9OVPJtqfji+Tq84t13h6pHQNwyVGk9bk8QBAUwjrfnVxrPdp311WsZOrQ8
jzkknudcsewb7ygSyFNXj0LERg7tyaWFKmeI1FYhWOWif4JGsL7KMSOVqv/W8dz4L5hQU12zYVlA
Pm/0ZpieUKLBmgUilAkhQSmawQcdtfJsYoUQfnA2d+MpzEywuE2lwNBJiC21hSO2oPs/gNHfRT8b
qm+2pllpSHI9AA2KEG1wlwGW7s0IGv3i/dYH0Suw5JlOr0bi5IURPS/kQ5DJN0/6pDqwCEX5NSq0
mamz0LBvCI88cPZlsNIIeDSGWpCZXJlPSdQWieo3K+XRyvo/ycDaA4mUc7/SdiJG8tLnauYQbMm7
W2M0BwMGZaELqPPjZbMoxnuKVjgrGr9/LrEkkC9vzrfEt7Z4VAIVsdGWKVBfEsRuaplsfr4jNsGu
GWF70oZJ0l/trMpuHXg+DAXK9iF/weCz1fQfTX7rES7IW9a5cAYA9A5YQwibZ0ejeni8sIVGQmsY
jo4Ao6iti749Dol0/LpRWBqCLBi2kL6+utXizmopBdxviocVrYg/nynot5+/11BrJ/Ew4u9Vg+z/
RCwoR3QuPc76Q0yh1lvvRPWJ+N4UzDjJjfIGWifU8oQko3UhADBt9RisLb/t3xrIRlPKnAU+P/kt
vG7dLMByRwQEkZPyuvm34SyHIQ22acOzrLS2qEAdiNnRCTvHAtx2ZtcNL9yWZDNbi3pqGdhqpBax
azBSZmXFbvEHoAKEmurJEID3oHT4ljxWU+9TyjB9rpXCBgaf3iV+XTGVwTDo/QXj64cO0AwS0zHr
dVfJItCVDgfkv0nS4OmWqhL2nXfBdGRZ/855eqkG7jXwMvEGZ1pZ1/EeCFeL39MGDyA9vQEfcaI6
rUQFR+Oy4kkxj8C+ubj7sh0md+CgJ+zWdfNG4jV+qDN8DARny3qJbDxE0i9bJcEVf/nthulMu0/9
nRx1+exO7xU9EI7NUXWL5x1J49IK0LOYxA8STIqTeUtX1ZMufU8cIlQ5Rhx8fE2kUtb697OwOTXj
xkoLp49zsq9F3Hi4ykNvT0PBgtfSTDtgWhZUU2UCr0B6CMZXg7vtsMrfudJkpydG0ier0pAHGQMM
dAyhNEQCnQNUy7OnQ41zTI9wCu2LPbZp2C2f8MEA5in+48QXd1Y3G3n0Np9o2oDt/kG61b4+KKcr
w7P4xOnfufCq9+LqKX92cS1SyC5Wj9jmQAZa5/4iViN+JxTBeD5/6OceIyFGn2CudA7kLptxXx+I
AbienAdRr9JfPoc6UQsqldTjHZxN23gdbi1WFn+Mi82HLmadKSwcNqXpNp0qi0y2EIdgyFncZTcL
ebHSQCJhZkEsXr5L3m6L+vzPWvDrHxGp2f7Z3/RgLX0h2Hi7Ivn7qT9ibtmNMv2lD2z42A4GMlIN
gm2dv0ivnyjd65QAFqC3Z6U8QJ4jLPq1Y4xmT3A97os3KU0U1AnUUOaLvOKTEew6+sbomPuWmgCh
5BKhkrEieevXO3yWeVvF7pZl6h3KFWeyOk33ikO61jY9C/lTq2njLiXHUXrr7/8UQDkxnnlrIGWA
pPMiBdkGMseJJPxH8WlmDeOcwFu7aG2cosRFjZfMq3doyp1Xj9mGQf2qgzY6XNfh912PelAuQAqO
MNsvPgEjfkPuDsEL0BK3ZPAyu/TtubR/5jSRkJh5A/Z7Hbd6qRLi1QKahEKxSEQz58FRqxh/yQ+M
dZQ4a5if054Os+70DFamkD4F40donhEHnDXc6HZO47TE95QZIKbd0JmTcKKF+TSUIZN3WeD7Lyj3
ZT48knBuDDAH2Tw08CgP9IPIJ1hKJKI20WfGOM3klp2BSrkzDK43iT0WlNqlm8EvkMo0SiQPJpg3
W+rYqYhENrAp+OpIAJ3LiS8PQH65rkm4DvKhbLrCygS3r2zTsL3s7b7FmdsAHVUQMjUI17yyzdl7
nh5W4SrrzWqXyQDoH+6Yx3Xjsh3A9R2CM73Oh2FlA/B+5+UjlR0HVtVYd1/4GBdC8MeK8jJ5jcmt
MC6haNtDXGHVPRdb8/J97Ut+8VgHLGateTIkCNUdaD/P6nUWMQqSgqqnPG5A+pmCJWVEogpRazWx
DUalhYLdO3tzqXdwJ4G3xUzNROglXd8qSrg0rxwoZZRdL1xADkJqcWaD1OsJI2h5ENctUY9cAf8F
jXKSM0V1VGILWaYkzDT3hb4KV1gcdnNKpM9CMQWc0OWg3aYZ3RZmRXNYv0RtD5yUFdNBAOPBCjtu
TJRFwEWMn1EiQc+m7RXSh9aWdsRmyxpJn85g4erg+HwYW62l1lCNLprG8KefIgHttKmHo3tnAtMO
rZG1x70DIFfZ2sE3VnXCat1SIm3ibBBZRRNpUpEn6XW5FUIcBXMKNzfNNIldzSugtmhkrTfoeUdC
BNTPvfojmlQapbZslC4it2eRy/qE8HvgM2g7W+IpNhsoa847i02/25FDHvsXHglH7ANafyRNIFCx
UNHMP/w38+7PWWQc10o5QlR+kb/267AoMWXTWzPJ99wdn6pT01yn8/hSFJv0i+bwqCqJSFNK0JQj
43ZsOaplkLb8IV/0WknApMIlb3JPJXz+Kegt89k9+eu03QY8P8UAZT91rPuHwXgW9Eh1oMOuDf9L
sU0UPZOnTKNK6ICyhDZ7BJze3ZCwBAuSevKx4VUZCwaOnwNcNpLDzaBLAhuYutjwbU3R8daigOpv
8WP8UCO9ur4DIcbntNyYKi1XeFUupzDyE5OYa3vV2ODJfG3lLUROWW4iT/recmPhfEMX9oBcsUTC
7v5GEEx80Om7a73D6on3Bbow5SXnZ782rIid4ekXUp7iWUy8/JArgdnjJNg1M9FVF8UfnVt4hkR1
MWbatqzb0S4vHacekbsg4qBvBhUCSa3gcXNwx2XFik4Mp2n6jM4cVAr9NsOdoUVzUSlQlzgg0jXq
qtdQLR0cFOzvni+o+CmPlryrd076hLZzP9MMOacd+A19dgz7Hhxu8/kfPbS8vg1lJQItoyv7PzBy
m0BEeRWHOOqPLsb0KUvJbi+uKN2PRfICIjgWbxUMjVnZpcrZ5p4g6QV6MZww4eKJDSwm8ga+C7qB
F/Z6sLUFWpB+owvf5HigVcfe8p3yPOkE61pgIITnydMi598Ge6AgvbrF4hpBcdYFnRH5iEBPVftF
pQMB27k/QIH6cvaa0qLOXawm98wGaXp1+0uK0ST5iXrKnOzRphF44oOvAqECmp7D5gZqy0Xw2E5U
YK6R0qNrOFvTytp3tJHUNLhO5JkAod05q+tYJ83C8/nrkjk5NmDaEBDI0X7qLYdE4hT10ObV0f+C
xJPWatJPRvviG1ObtLZGU9t6ugyLmbJSZWqVK7FceehBjDQnnWSwnh6tOboGQGuz8xBMlEVVB8TD
4c1Fwypo8Z6iIjdaATmo6pW7+cX62Z7sr0y98XQsIV9H72jqVZSCkiWx61KjRvM8+YjKJKNLOew+
SRahoOE6XHO6swVejM8Wv2J0gAHxfg+xN/1RBjPpdIdJaTdEStBDZpJT8l2NNgfGUgIjdDY7rCt7
WuwgHosNUWpmX4dXRDzNYd9GvOT6co+EMFxJ16ED69ueTsOEL3Vw1p3L0tWhuYlwQBA6HHu6LFOn
cxLeUlh++W4RKzsqVxTLzPPU0O7akXvPGVkl52kr3FvvGGu73JAHyJQunND0NEqdjjMB98EHXEvh
bKbbd7GYqklTnOBTih0Ozb/qfiOmnLpmWqogxdRRUFYmBWm4mc7Qa/x6BB7yl9vZYmrgkVg6FD/x
kvudKq9HG1vJkYAp6pJjyb9AVRPKJW1/WEJ8n+nL4OI0fmq+tR8b8B/r62NEG/eW9v5PDtaJnRXx
83qickaDJSfBKmNqwW/opTh0n190oXO3CCpZmRM0oCuFwbkvlvo6pFBfF3X4M0rf7AOqDJx5uxE5
A8Pa5DiOxRC10L1LPGTLZGDHpjfb8GPrtVIJmGGEXz7pJytNLaf5dsf8fdLfE7JSmPBx7ebQlUrv
22qneMYWq2L1jgevH+bZP/xH97Dardm9N302KJzEx8phHlwy2ZaK6IwwUFsoS+6kAE1d89QBfYfJ
J8z/1JYFu2NvnkG6uSFyWNfbS7u65UADKEIcF2vBfsmxBejdbynaEzfVjivXPTj6ZXgQft+WF6aC
EUwzcK29I4q/DGIeYEp9jBUPGrkBDGo9/KE6MZI9LwoCoOVrdb12yIgjmF1DGWQsl+dkRhv5q3w+
M2NI8nl36WLK4nzcgBL0HZwzOsI/TtD3KRR6EHaWrMMyfjrEKh04ppqtL1qCJ+zl7rXJPKi72dcp
0NT9yQK6Jd+tifUK/mnepsCgarkUh8GMc4seWajfOXGIOReEhNUmvbYYqgMRrJVnXE0/pUSCDkU3
dFabp3NNqkHO0oZdLl9PvUVSxdSupephDsJIyGwY2qyDcW7NJ/+Ne7B96wFhUH1cyZCAVPN+nXUI
COaAI4JmD8hVM2tOWIsuPc/ukySVSxWcV13cfUbYzpYGmna1OMZgDtNR9qvq2QxF8tmRrSiyBL4p
ds7WPXGwSjHus5eazTy8JZxFIjDa9DCx0t3Ot5kEd+HI2ykzVeD+3UjxewfXsHtRNF53eyWT3P0h
vEeqil64RVUEujL9DAZOkTkLlpEqmfkX5aJXcuxw/7uh9DaBW48gH0LiUxG0VJAdENUpBXqR/IP1
Jmwx69rahQjUa+CtAim0Ng7k2gIVkko30x3KtjOq8fKNhuPHplt0pZjFq3dBO+pkqdjFIzsUDNV2
6fptFvZ23zrgXDPej0/+0vWN+j9EJ0CR3c0btM9woI66154F+MSXYb+7YijsY8xI0gu1425+BQb9
MFQsoxaNkYk6sedorcKFL7VQJh0oL2khmVeCX2DqTEOWJ/eNgXtUeSJUwFX5nqq9cFpLGuSYYzPb
sCHdQ9cNeoiU8modGZtlw7NpiWXTkB5abt/IeSYCoA1csDBA3XRskiuKeLErluqvxAahpj8lVJSD
u/NYi74izFZzMI4Z9f2vlQToARuxa1Ev9LntG7EGSXaKylCcgPiQ045ke2hEmsKjeN4u3bzg4xjm
qZQqNTmYPm8VZ7/MkinnQ9VU2cH50/RNQnHTBv6e9yYnSEmSH9qWJJ3SKvKz3SPlCKaqQ8mKIjwK
pLouCoyL3vttXBF5+n3+Pm4ziws3gxCzgu/8qvTeEiG3QlSpn1Dc+D0TlP+TGzqfeVLEAJa8lvQv
HjiBIDqrKN6FV79yNjbJj9GJBVS0MpACQB2RdReB2DWXqD9U/ilOwnvV+DBuILslNiamzxIsd15n
ypSYd3FKZV+XKxC6q27znIJOiR/aFKMsMQ8a6Bhcwv6sGMRgsoAZ6/VzGFgogtuSksEvkHEI0caT
QJl6YIWpImO9f3Lht0JhGmUK7oVWgq+/jYhX4QBQaCj0Wa88XHHCW2KZ3K3UhtNfbBbSq5a/69AL
TX0A3QfOa6LIzUeGX7ekSTjbD0TKM4sQ7La1hhFuVGfAYPevwbUjTIYidlXRLJiW9qelmVaYmlz4
50FoV/yc38l7m6Vr4lw8JDXTTKHTp/t8A7rwUooq0idRg+m6hLtNtHTZ3j+CLxvZ+HjZeWE9KFQ7
q6i77LQ7nAFPGhXNnyyP1k2Bkhx+T4OZoJ1y96xNnCJfLunwbxu4EDVRxzoD9NgMfbKnLenWcZvH
P5SpmKz/TsXGT/4GLdMQxxkvWaVQQYcQtOQJOjTGh69KHogJEsIWUh7dqtqjNUNGrNdyotAhHrgK
uCYNZUocC0VO7rXuznqLrItKo/bZ1SyiRFIiznuUopf9vpyDjj1bSKeuP0PyFAQ5YC85Xo/UZu1o
7/CR8Ea8i3tqmjHD/Vk/e4XaG+vpR//k4dsL61RScJcvl2YUr1lzby/1PxBYYXopVeQx9EtyPvKI
HbMkzl7PEk6jT1cSFROBGM7cmUdDqLmAd8fA1ZDINkS+GPKvirlu1MngGhrAIyg4LhOIOw8+Q6na
livimiwcQ8skjVWf5plYJsRsb86kwwS2VabwFodvo6F4CKx96fZft4o23opsVDM0lofuw/6B6pSj
LxzR4rBMNzXeGNPEek0oqzsq4aGuwcZ5iefhukTYAKOS6UR14V5sHkstGkMyoVtawp+1ZOqLKbtE
ndxWQLnF1LxRmEmrkrBbUsPhfb1ZTXlaWW5G97Jrf4EutA8RHc2IdsvzNvaxIZTDh33TqJnR5yrF
n+EPV4dT8VbMXPOuA1rGAyROEoczWEQigm3c9AC4cO44KSHS5rGONOoV0FVUM4ZPbG4n9oQpUPVP
jzZd/sxPB0UcRisSb7I7UFlB3qGYhbTO0EhIjDkCunNd+8Zkzmwm+juQM79HnhLZ9G7DILFfs2AH
c7zOqtdA+icAk0hpSIKT5dPjQe+3GTGHiGB6WKFvpxZKN+1roR7FGWF8shZ6AC4Dd5LXElQeNCQY
i2e/EuidsOySgaA1UtsGmhlW/IVyPmvjMHYXVuB4Ab+H+wYNh02sl9j63uzqWy20ilZIq0mV/6Mz
xrABPVI0ZRXzbTwnIBudgKGwM+Wfut+D1aF5ZiR6gayIK8ucQP8xeUSQlkTqhOpt56c/+NSqkvL5
P1WR7903UJ/gZwiITGfT+9LGemsRSo9rGL9e3IktFoce5/Xe2TE/Nu8HvHE/DbR6FM1UcoFqxhm6
eg3MuSgRtsw/ihUm1djT2C3lqQAZjO1R/iM2PHa2TxHDKFoTADBOXiNfkubfb0kLsdyEc1AdDBGz
2oOeHlfgGE4YhkgO2gB1hWkZOToSsBZ8KIScocDQj40oXCI8LtPNjjeU21lU2vbin6HzunE189NG
+r6kCkFG/4nvJ35Orjv+0obaN2VpD4jhnN8CuLtwAY+Rj9d2vJAfljDUr1fT1fZRLqywnlGBsI6L
UKDJZKh6recQsqOonguGzC1QyLFk5rWn6NCj8zW0lVxLw0Cla1IHyTMBvHxcuUuAmaPhyI/UvWST
rWQJHats8AMxgZVQ1nLbcL1AfTAJVpN6QNJXYjcU4SHgI8ISL3eMgaCjkCV1oeBdTx1h3Ig32m2w
vi4sv/hKk0fMkkMoaMQFOt314qVLQhmTZ+yvmvbIq9TfJ/pv6qpd67qzNflOpAqmmWSpiMoodNdz
aMMZJSK47yT+x8iyDrglOQrBHJ67fEheTfQgxg2r0TlC2/rztL/q+rNb3uTXGCRqBMG87umxST5J
NUtSK2thIw0kBLVinEDQrz+vXlUgKjyYtgNLrccjlSfl/kE59HU29YfnKp0095O1YejEO7BGAf7o
7cVKnAAq4ME+Ea2fHDyQtDLqZTyQQEaTKNzlqfGtvpmnGSjW4yb4+bYSnhKZ4SffC+B6xGobqTdU
J8cYNSLr3T2UWtA4fSeqvEnyv13LWkZ+MBR6oCVUx+uHhGhXaRvvFiObygVOjkxShoJ5sfBUSiZl
GUblFahziRizaXDrQ7BjbY1OGBF1+5OIoI2rhDT2uhF/qA2S9a82WuGYSv3+eqXPgYL1UxHxZuDb
hs254Uk3KOVm2gIczrnc1mptkfHn+0pov6JXBFGjnI/xq4eMLhvpVBbwXDe4KOkSkBp+uCJkQ848
RV0IFJeWWybECrT5VWGExGcjrySp1cHCd+dTrspxhy2CipIzbYXih6OZ2PohxRKBi6iRYSeSt4p+
BGvDFR1WrvQkXSwJuAOhblIUCJk8pIU2JIW99CqyL9BQV9JHfbyAz6t1ecVJokYVHOSH4MUNp/P/
phPFKwVZLBZkKia06nCHFWgl7VaZ4+61ZWQvTxZq5mWVADiwq86XsAz+TuRkrlcWzuJnVDDAODBS
xdzh5a8u+AlpmyonpT20UJi7dGra6qHM8o5vTfJSjftj3F0rErqDSrpzcYl7JKpYNHLRb739JEal
0BQipGR43fQ0D0J4ue43ESiDqYXrLs039f/AzpSUkEr+9Fb0vZjtVKiPhGxMSMluuEWSfRbUX7T1
zW/bwZY16QB78/DdriT7R/cWflmdRzx5Je9HkOID01u10hP2zRiC7rOL8aMDIVvAO44cZjrUphC3
fKehRvEOFetowd+cuWa/yAxX5JgPXP/KjhT2uqFBHwnf1HSAUBmIIjrwxAD+0cGSxSHcRXlYz4Vs
E6vu1D+Bang5mJUeBmuR+qFuPKsy4bWfEHUh8+JGtxF9N6BWPvKEn7WKu22wve3eWYusAY3U0PKZ
6ieAKRNHYbLH9k9qb3xrsXD/0TNRWRNcVTd102QCcZaclxNfodmJRJwurt7ZsDPe1htQxhRq4bQ4
YAQkg+j31hrdjuyCNQfys+pby6lzz4mYfvmb+oPnatbCWqKEsraJlnTbSXKp6U3RNHeAmrAFtkVB
7GIIwbhk3Kw/HKuGzCG8kds8UUczPcR68JeyKCwj781+lI9DeOg9s6MN0/2UVyBXjyi6kuHVY9qS
NQcmxB/LwCXkQwb/3/RKqSm8fp1MJfuu34oVWkDX/593phz40K0Z5dXnwTiQKCe1xyyIt+PpLtni
daU5lMPVGoyDyQ4dETpOUwMP/TeiLb8ZLxRGT7wBocqz9k3k/ZHYFsU0MfoRHgB4WdJ03NUd8HsL
bRThpu7tRYesjfIdPj+sSJ0O6vGTFo+v3RgJ6aXr/SJ26UPDor/97pl8/ku8EjFxparIoxckZa3s
3I7rdkbnMIqOqWsnKQ+7LSuzCkoeAV+n1P3MZwUdc+UitV7rky5hkzLrOPh/yrgYdQJXjp2b+BpI
5rAXjr51bBnwhOwYfhWWfphF8JBnKWJEh1jiPprnoldSV7+UbJPFlvLFi9/ixRk5Y4YVdvBE9j4o
4RrYRbScoAXVjaORE+7xV6I/27XFS9RL5bH7j9Bl7WiOxm1cRWH1gGbTUG1a1UBAbDJvZTytgk6E
O+xB2V2ScAwTiEakJs/HeqPNuAEDML7GE1v5IIHuRk05YcyK2/HZC1M8MEIFznbW0fpDgNffiroW
e0uwZZdV/u8qNDL8lR46R94xBSSYxUTi0eYyWOHtbT6aRpjcLrm84RrmVVV9/8+7AJLANDlxm95R
8ueHzvM6oF6eVdRpvD1rf+QlM6M27FqPdcmwaqDj+xhbRLYNdI3TFpick4f/CbmbYMb93+ya4Bm0
oPwMdXZII4LvChGcYORVJnpOSPDmn//mwAKRt+PNG8DNWAhlug+9I/JPDgy7P2fnB20gZmYGStYq
O05b1vpChejDPiJvYm6vN85IMXlU9+F3G31Bu6IW2tKx+3xbDA2GOpZ/uD4t7qIPeI72Yls1Ndi/
ER1tgqWXynFIKUIZKhcGOCb0sCT/YFivgVSGdAB5xO2cZ5iEEi8YCF4ARGN9N+tBmoSAXHPx0Enl
r3NmdgtZxoPwoL0AOrjsK+aw1qOb6jtsm7mJZcTYSFZFF4fdWZEDS8+zyw3HL260U7VvBr6g2GCB
GqQj+NShj4D4E94ROZjDfOcpi5MdEGmXia44w7gcTFvtw8CvNRhh6uYNhj9De8Ny477z9vXVJ4mc
mRKZFlaCwmVuwzOcnachji9XndB0rJ4dFEIQc80E55VQhaq2qaJ8Mz4QTZXHm3gAPKg+yvSCjcqy
7y2JhVc6BLvDUswaeZCsCnrYospB4k62Aqo9qgr5OUvVemhZUV3ARatge0XjI533Oe4iNF4qbel0
wp9fmh9OFAmmA1apGWzK6qYljKWDHeEFys6V98phFSzz7IxSOTIAucMOZczsZ4NRFKw4cMe0zyFw
OAkUJ/o/+H+ZX/RdFgH2qVnYAkhLvNMlm8+LsihVJzK6QIjGBXt+1UbUCcB9o09+ZiMFGeVWOEKA
L6xljI99lGY2ZjMK5LR5lLQxHVyOP1gOjIMOwe5gJ7/lXoA12JMKTB16SVky6/sezpQJD/vOrPtV
zURzwHxWIYA1MtxW6+N31xWD0hMcqeUovNiiljprBv6+3uzSPW7mHKwbfYzB1F5ZQhcz5lysdJJ0
Jh5lvxIGpYngoOv+j+HnVmnKAsk8D0WaOMyVBXslENi3+/tYBxtDvGdWiGdkuku6q4viAqTdcBLZ
hnCSH3UOe1AfA6Hpr/QrPLAOiPOR3H+TSjaiEffxnu6TDhk+VM/WWwgswgXFImmpCP3ICX8eM7Qu
Oy05spY8xpkJGw4wX7PhTzGh18qzMxAu33xCevDUgS02r/o6f/OLVYAbpfeFOytBowzapcj7wYM1
2OA8mOGRlB7QAu4pyFUdw98BqJqaAQNx31cmPQOWJfKL4QAmIhqU6oSEAhfOSQph1SXQgSoSW99x
JAf5raQxy0oXu0rVdppUOKbAT9OshNagZCA0nnxZSjxRG5UR31BAWRjkGFxVq8EOXJqC7CE9RU1l
pR6qrwGhJ4xXrhTjxCiK4rXWUrElIw2a5dhEiRsGpaY0a68aQoahXioON0FpnsipI9vlFxl17mKa
pDlo6fGkDMJxDKpt63GCFIOoXDQ1DA3fW5iDpjDiEPii8vrswK97iBZk/7jPESoiKqypvbz8+YNF
TYGEu3LFa7GbpU+cOFPY8UTLcjNEkCy1A4OORkVyXUQIwbtA4WJgLYc3nAZrSAjPTmuUSKBr+9xQ
T1NVJogUJGwU1ffG0TgReo1hlGmRK/GySE8qoSreTxtoJNkzU+/aAwpcLx455lrcv3ovG0BAMuzX
2R6fQTqL81vg6VMg+dW22wmC67u/yqnDhoEVZJfGyKfV0fmAvlPglhcLsxabfBbssjFUE8rjtleI
mUwewsvwsnyumAA5FrJEHWJ82z5shO3SoGwXko+ZKeclnUz8NHvzVvYAFE5Kfrat4wNik932e51/
PLkJ1b3xAmiGZBBGiAsn2btKOIPAcs9evUqjZfrShrGgLLBWrUJKY086zA2eawCg2EB1UhFPaaiz
PUR1Eds+CLaDl1XeBMpR/EV3EeNum5aygFP5Thwm0nNrzSgrAIr/WkgaiaVoQe7waOi9MQbTEyVi
K5vZJ9tlEv2ahzgYIBekgeus3UapL86XQKXdVCIxaLlbHv7U4po3KXgLMaesSOtTGbW4hX7DxQRY
JY6XNZtjct2FCEVf6KlVNdfcFuwmyDf8ohIRpLyXiZpCdlmYwEFsTpDnpAlhIxNI7bb3v3Wv7Q5v
Ptfjs4t8FaRIZ3dPrB8v0yCJbr5ThnkoVZMM17IocBo/BONhVE7sdUE823ut7noZDQsEntcJh90N
MHoaiGOndsxUMXRmLiMmFXoVlb6VyWZHQQ8GsImn3EKugzSEPLLfBvi7Vq7LXlV5OIED0ETuh4Hs
+/Kd17dvloo1ClfQDJPKgo6GqrM1ay0xTgnL08vjvqVrzOnE5cT1RKvIrjlL2lfchtVMmSQx4aMM
FWksQGh2EJAfZ9jSTyMCrE8Qy59O6gEGPmhlMZcOFWVsQ3fOj/mXQ764qq1OJTzMHQ3dWawvinls
OhFvGaxOZE2sh70kCN0FlWKx/ULUKlLo4uQwZEstjQiGau7FGB9glJHVUHsbQLPW0TQjUs0cpE24
eII3lypreo8LdzUfdbulEaYteBBc8uy/ivsjBUq+sz275YnA5RO0HaShQyjjEM0slvY2NYq/QLrf
bQm62PQWwMiDQGLu+A20IxfYzid99oHKjXoWlSUxeRqaWTNpnvU3/DkA4IMBTuWDmLVx8kKpIkGb
sEysF4nZ1QmeHB78owT1nOo6kWAGl1P9SjhoqQDZ7kcKlAmKvzKOOisUFWmvFDpxikzMNjZ0z5UQ
V2pO4D9QkMBFX43Dq7axmMJ+qfLrk8Jp9zxUt72VyPZ/eDS/WR+bfe5flqZ2p57PL9sM7Xc3xUue
shwWDoQeFfeDhH+MHzAP8RQMNPFgw9N0r4A9wRobAetcfoHQg4rz8u8Jq8xBB4xYpsY5zkriiV5e
qNRZHFCvtXE1VLFq6IW37TCq9FRwCtYkLO8UVU1pgc24toBgaKyFULRGoOBIWKMSo14Hv5tm1dSM
dfCbHrxA8XNam5MGl0Tsf6eMBXp9ftifcWcsfKZMaDBiG8tV3va14SKRBGMsBRcsA2dqk2Q7Ogwx
b2BpYEirXNA/tKFAV38NN0jf1ANG6Ch1Uf4ehRpib1v0j5TX2gws+MlUGpw98rWocOcp8O1MFi30
n+JlwCDTY6gP5mqiyFsEeSAxxgi5UT62RKgRv9M4vlLJO+jzSb6N1cUu+te9Ac/BRyb1oYx0Q2yl
vGHQ/csh4anmJgG2azDMCoPyKcNAUkSStusy+yyfSPzwRvDfeWUUGTTfRE840FT8v+lAv9GWa+Zc
/9FiSRoSLKMYWuQiHdBdzi/5UPEEjMW+hkp9hv6F6Zf6vvF0/s5eQbT/d7lDeWXCJuqLW9qmhI5T
nIyWCxSULGgmG4lE7TCIdpYbR5/P6eRtmZmU97KjcOudTyd+tMDY+dwEEDaEIYddSZfQdI3jjy/L
PbWU8EHCQyIkDlmL1cC6kVFGP3G+ERBSLvlj9eHTfjS3YhHOK0AgfbZ6KENdCfldcuqlq8lZbutU
d9OAf9yNwh/DEo57JykJdfjH1r22v7AFdjBNkTqRNqBuApgeEVKKn2fV8h7cUnrFKsd7sEoDnANk
fQucb/pYVD3u5s/PBfJJAKnOdJsplKMH9Yaeb/clZo74KA5iqO7GtrySjXGl4p/1VK0e0GY+rNSa
6tbpvk5AutTsXm6JeEbl7cUxBN8FKtKD8/e1XLV+J2diB+Une1T4kEDi7vwBhX3NKQrq0Czp3E1W
vYKqADEW+a4jiIfXajjAIE0UbG3kIyLliwM0a99qi0M3B04KjDxIu6fZ4BCv3Vu4YxmI+UKqARMJ
4sjGhbHrZhOyoJLijKD4j4eQzgMixxcoTGJ+75qpZ2B18q6kWzIJ0balVZ0250omz3s+te23738t
XGEn7N2BzLUYOSOMgyxWHY1nfl2ZIYLaPVFjcJi/GbZV45n7hVw5IH6+pbJ8HwkTuHnsgNJ/I4gy
ss4n8hBL4/EwTH0wfIMzd83Jza7f5SLgR5BXpSEb1abCVnV9YYzGS1c+jLmhyKdH9tCu/D8jBK63
uJFszLtZjOjt51+IWZc3O9lfq5LKHSBJlNCknD0pD2r1P09+36eaGeO5ch9qJcZG4+zCU3B9hWaH
FfXOHjW8Y+LpKYzILmoCIETvMHdJOoRLgGyblAEgPSvas3ueC+czAaBDnanZjFiNwzsVrNj8kMuZ
cmRyF6ZoiLIEmapL4+TqGYBIPjaDapAvJxZVZvEP1rh1YE7aCPjJKwCGpzRvE7R/Sqfu3anTP1jw
M1RtvTMIYS6D/vlwGHUOXJQ/fGE6Fcs6njyVjmD9SM/6hhtskRaC6HDMIUpnIykeulmx1cM1c2Ro
W5gckR5hMnKFlfDpi3YpmQEuSTkNVbx2DwMLq1yyzIO5vhumqq/eag6AgOc3JNweLwqXNaAp3PyZ
zHUtpC384f59m9nUdci+IXB67/6gchmx9p59uGL0W2LIWrAzl6Z+H4r53ultFKuKlJePgkxdJ/89
rQxdohYxIGvw/V3uBMISLrXQpHxfgT9xZ8qCebS8IuS1XdRsyZeqCOL6/u/GVx2T20bwbXC5Bo6L
93lODMHUBJKH0Kb7hb7K5acGIsAnl74tnwprU1Kp2oEU3Jlur0dEL2pXq5T3Snb93LF0XkSl7tO/
KLFT0DPp1NRE1w055NcTwoWYsR7G08fy8A6faETE5XAKZtxeXLs4jWo035GvoBMMnwBPJcSJxMcB
CDJjDkYX/3t9pLC+jDAaXROvQTV4LxijJl6gF0d4GP1upPHXAfU1jGXE/ji6GuQPaAZkSlBdQ4le
kbNNoNxNFpkekyFNe8q9TUuAabd50WZmeUOi7WU56e4bx9qpZ1euQbalu4++Ii7ynhiRYUopOJny
7SSs+3PFfnfFj5JykUmXThmlAbQ0AzkGGk1R1vxoHcnHHsTPzJvqhrRpjd+4AoCwhkb8wZ4yd4Vc
QwKleIwMBm4D5hzX0oSRZi4hO8suprnjUyaih4NFQnCaNNvJ5rtZ9kcpQj6rMQRTkmZFMM1HIUQe
iqrRzyoeo/Yi2omxciTef27sXk251QImR5x2tZvXBQr5N0C9yzo8fVw78e0ffRNk3xXF/gIFO+Xn
O6RaMUKcZ8zZKhT/mjB7YlM9KU45TOCym9nOcf2KQxYGDJZdTqN4U2SMvXSoy1RE6qRcBlb9nPQQ
6Rpj3XEpkXowDaEPhuJjdLJo1MOwDjMFWvwLbGbHyY5OvBe25JwwtyqF0wdSVtnJ1BcSnMp7ue16
U+WoU8r0dSwJFkrFSC14H+48zCor6oBUol5U5susFjSthpZEsvgejoNFv0oVb9Sz+MMGstFz5X+b
1po+0Xq9+Ae2eSKQI4G+C/CSxbUyjylHYm9wiQfeJvlaef8HZ5il+0Wnz5zwubUaMWF890sOF6rs
oGFI0Y0o/TjT3tUzrrbCxidkxHkqbKF5r+NflhzPBFq4it3kZRGTbORDiOLNGzZlQnLUtKI1KxQV
A1iyOIbZm1HW5NY4u6prOhwMixZA2uBnjB46cV2Zhe/DIr9ib5Jo85ZsYdRMVF/OpQlg9Cyz0PWu
ckBNl+rLDIJpv3ytuAfLr49NbFTcb/LmgBvJgRtgPCzozhgwCXK2iLk1zmA81/L3FIgm/H+q2uxf
yyX09w5YtBphP/vr/OabQkprX1TOIQKMSpKQk6xGeSQMGBzkRjN0HPG9kJtPZGshGHFhpazhE2AI
mROlhlI+5DBTQFgrRc8BEqyQobCM7zpcJmJKuqwZT9KWziuObnunuEm55PiewkFyoEDK7dWHnhDq
tX3TlzkE8o/mESMO8TZ1CF+Q9P1rkM7PVGgvGAe5oXIJ0ywZgvuR6xXiihkoEYYQWrCFIIOYdkOR
iWnl06CwIQEZpbepeXX3XAbsNS0TvAnkioslWcN7XKuekajiWRrcg37v11ViAnBfmbsbFrooNSq5
zLj9vjM9alMqejlOgIrTuFAf1AnWou1ST/96Ym2pOJIUXhRTJ4TTjUchnZ1YDI8VwGsJ8O/Dn7Ec
vGqHBbulrXqufroAP9Uclpx6T+exS5CJoif3zq7DlPGhuC1QlqpUXxRyrqTJFbLGCr8TCT2N+pZP
FzZzW2i/r1a+mBpN64xUS8FAj+jFKw+FgeWb62Qzk+MFTQ9X/5KGWuB2fOXJDrYqAneQHxIH1C04
ifGfhcU5yoW0wpDWe6qyHJFCNUlSQakYslqFqioVulBtx0b1PDr2IePwaUBUR6tneD4VffUMdfZx
3wJaALP1GRZ3OUT8caHbNwggBwNfSHtJzKOunan8b0NtcDcaKYqcZAya41LvCLQItN1N5GeVQyL8
EYGFyp0NoqdRjAdeJeeTU5VooB6BJbpaf+pRGMu77FiIzI/fLz3uLFlBijYisTgcaO0B5U1fRHYg
wQK246VcKIr0Piv1RBBJBTsjjhqiZIS/3tHsFMKwX3qaDpM2GlsEu4SyGJNjnWbBdSwqI2m5bjXS
9qfsQj2pJeapM+FdpOuyrTvG5YEgPetbC4EfrAd9Q0HUIlz5gRuAwW2/tS8Hi+ckllTc8WBlJgpG
l2uNsYa1uvNbWlPbsom3zug9TjpI0mGetTDQsTmHYTmBDmUF4gNvoCDvSmUVzN/sUh1UFqCAE+3f
tOyTvsOKmCJjt0AAVo1PoZ9JPlFMlLk2Yl+2+j8ygVbmEi2N7F4hgUUhNVyGhPpduUwRcyVAK7hH
Qec8ouIoVkl/5tsUzCTN8nMo4UVb5/yDbCJIjwyPf7beWhQioKxTT3VlGCI+HZX9ctLFdJwuFNNX
8OC83nYFSUql+PypiaEVMNJBIykQW3g7SD8AvdxYmGDZLKJ41x2zgt3tRHCPbqOIUWu19jhjqqBZ
2beHMvcSNMg7ZopY04dqWtezA6B8sidH8/+k/4TstfZAZyNedP+KG3ng8ptuapbIIyTaMdovNOei
llUMvSOLNZ4llSVmaNnN5ur2WVTvbwyhPLFKnmJIJQyq8mfbwyaAi6Y7a89r3ODiOB+DBh/Km9ky
I/OvWRGFiHv3PDl5QzDBouYFCFH6FkYTbA3HhjxNAgWVqAYlQcsb46ScERZrDe68xZk+w3iK1e+9
NlbyuIC/SMcFMODe6luAJP6pjbBPhQnPAtoG7XyyVEIuJaItjtmLLg0oOjQu7n8rMpv2xDOU9jL8
ihu+MYi5f0vso0CA47B65RkiQA4HAYYySZ66C+J0HRxfcXfgW3cWWRK51WLBt2EI94NX8NT4L5it
q8Tdsm8F9C2ZlXz/q4UrNF7mZkjNaQk/6kIqHFrPiI1t+K62SSxnln8PgJtcNDOPP03L596NmhR/
z80b26TkQxkavpTlVipjhfvKmFb8VJ3+/944sgxwxyjM+Q5uXmdc1a/vZvDs3Qxnj+tgHLw5Md8d
1vRZnQVcOevAK//yTRVaksP7XG2DGfqTj4y9edAhyUZfdJFcjgYRh7yHZF85wytlpzwIWs2ii5Bq
CT/s+p5w3at8rULcSOXu+a1j1pvHdJI8Pmbi4YsphTP4NGi+p6AGjbgK8vGU531TGrU3XCB7aGjO
5BXSo9Y/W5jjplgJIcvG3zrSYKI8xkzvr5IpQjMLHATd/SPESIZLwpAR+JXNVRMQ9lJZ+So2Kh5E
le/kW2/9uIJr616an4O9OvwwSKtJOADLP3OM5ZGZe3ncbngc4WltiiX0npBjhWxsw3QQ3qqq+ZsW
ebhWDgn6dbpfyBVylieMT/FvYtucMwUfE51fm0ySBoA1OwC1mi4YQwougV76byS7wkT4gFrdtM5X
p8sGRqU1XXcQwWHbHImT0ee+YW6VwTp4Sh+kMZk5XY3gQQ52rtb8BW+cs8R84OXPT+X3NmlmSxHq
PESe4K0HDgXYA807X9hdnAE5PjBHiuBU0uHUAmZmE/sSV1w3cdHESWzVJyD53rgsY6G+5Onz9ivG
xILkUZTj1gl2aF2PSvB5RvdkP4Zf6CIEwizn9iAFjKFpjd4zp6PdEj/bqyi05jiODklkLHjSrpze
kEPkEYpeDX3udl0DCbxlfH18NX8jvsAoaSo74SogH9DFkzwX633bx+kdfqVlBLI+kWOiXtYL9OUf
pRU/wolsiTRCfOgBlXXkwo1WRsjMyVJ4Kg2Z3JEeiFcuWqjf7rsDGHMFvXknFi+9loT5p6vEd2/+
wRL6JJ/DBZ8X2xsbSqb8GIs1B+KR7pDp45KlGrTrlsNoIRheKTQbQEgaYMhgFwyCbO9btq3XR87c
sCJ7GuP5IE4DVSHfAXeDq6mRg8a0Jk2943E1ImKyZif025zUrkQNaTF7EuSexPLyaw+yKxjAKusd
rXctWZHAU/h5IY3CKCP5mWyWwQjLzTCCoEtKxnNSQc37shPpWphCnaCg5PzY5JBBwn9FOoIBCvJl
l2ETuR3Q7o9hYCEwb1WbBcxkcaXjxLJhH24KrUE6AQgSauqDflRioPHtqy8wQmh2fuoAxxZnR3pU
06ol2YdPEbDFJeA/REwMAxiF62Z9DOYOZMbBDyQt022Re96DmwpX02TMURaWxxRSAWfTDdO+qbKQ
wGH287UYTMSlkAYLPZk52s5hVD7dvwtsXZuURJlWEKAO1DzSwyIzZOpVGPw4a79hk/IdbVYFRrvw
/S2MTRWi7cGeenpChpuVTYkv4Gz/Hk2zSTt9zcLUL2efvWw+VjrSG6bZqqPd5B5lHzxyUObc4dwk
TFz7CdnN5Izob3yK8CVvJRGAeeR3B/VrydoR5GKe1zpDEPw7p+EJGsZY8boSQAHuPh6n1vVWMRnZ
MJMtthMbTAGAfVCmxlzGlso2EifBFIDCsKpHdhF6ifx1csGk0Tjj39gk7Aw/Ss1uemxB/DyN1Qa3
K/Y88EQpYNKbPDfXIW1S77RuH6Qd5VSJ8oL3kvThxgGDWv/nBWdBJPfTEBBCMkifW1xk1dPyodWM
vS8yKFvZyAIXFmUMJ7ZMXwIWmE85V1Wxwm7df653Ii3/ED/qTVlWQcDjxNzVhh2Gw6qvdUHDEB1w
PR/F+zHRmNIltSeYHSJN/SXCEpwV+nuaHONC5CXxkFqhizjbQclEkONmeJhq3W0/CQ5FTFMQicxq
AjFdJ5IHX7I2WnQT+WWA3vir28wCB6WrypnxQwgLQnWoj2jUQZcV3BQqORpVTNSnxwTVnsPWuAch
RYAz+K2rEFzeLTNEmg1MMyB2NPs/vPUnN8NFQaDNZtJRGFyK1XWCSqFVUpE54EMWdu3FiHfLpz2+
fT4XVIRsKGEsgqyp+S+jOKFqTdxhCrG7c3GnbsfAGKTy14IskvQ9ux0SBzUsNDhES0Bj8Wt6dMfy
/vIrmeTW7ta9dQjmfkeHirwxXQS7bEmJf7KjwLfhcNjbFYPctwLJLtXEqNE4pqD6X81vIlwoerxs
158qK/eC5zCQYcFAS5oGKmySnTMDr4xwOxM/y6TI5BG+o0m+FwmrsbI7EN6d+E5pfZBrvtyQZmVZ
oXzEJHS2K48lv2pqiygx1P9ntSWE7PH0jcF9m4qP9oXAlw3E5bgsVZmoGNyqey5LthJ7SCwHHHOx
+xnAnr3pYGzKoNOgmWJq0WtKi/xqNpeEzjEaGUiR8DQWut6UO6HpmH7CQ5NwHOJdPSipur3ZWkxv
BB441V7981L/U+mo2REV7e586Pi0OflUul0hy+a0KJzCGIhkSAUrjAUPWAWnVfGbG89DuycomBAs
/NTTf4ukwhUS/SY2lHaEz9sj4CT5NyGb7mOTg2SVpm1u/KJRzpTaxA7UrRnDhxj0tOr9V678kjZM
/OjUjyAP8HczRI8/jrtGcQNZmjy/pzlFg2HN6LO28DIHoblab3roOSIbBHftVJYRtXz8f2pWs817
bSwXPI6CldNUsXv+QPOzp+KU9+8Y3dl25in1mkFFb154f9yyLfmXU49vaaJL9ndXI4NSUY3ZfIZm
RgWe6mhi+vYYzevFSYfGnKp5BlVROosjOzBVW+dizvycmKxLPaksgHVEuzehlTcyh+vtRiiTRapo
jZrwrXRsdMY0lPVsjSWiCTGsOQ9NlEBHXx3UWjO21IiS8mjevgTf8smQa2+PUx+EYiSTug7a5ASU
ynzyCmUUf7sUF7nzyjNE1yl4YTGTyOWxICbl30raBHcR+yryhL1jLwlwnkWBCegsD1MZpeJAgbNK
TTaZKS7NEqcGxUcVq2Yfh2QGdbY7k9RAEpqM6ysmqJE+o9HRUTEV95u2qVz8JoeE8pyKe/hel350
wuHku+sbzRiLrV8fOE4+oOrP4O60SCy5VuQ7mzIR8w5mtdPcgUJacAdZAMRtaMV8whLWAXO50leg
tgOjhoqDuaoQNnUo3E7dDnlfEk2AOFl7vI5QOL0IUFU45BlbvFcF2Tj9AHZzAP0UtijokkomOEIu
iIxbvFNR1SIThCYQLWA4NOC9PCyD6bWWWLQrDcZND4XXZ57t2T0td221TvvzTu97e3CYtmKC2XQx
D3Jdmi+pl7wr2RIv8wpXUqfxopt3OdPwDLR0WBrLbK5aaXhtzam6mguvyVFOnuyykKZbxojvuc66
SWjGc4jW3v/xsn/LfI76OYKs9WJq0m8Jh03lBEndHPx1ZAhYAGf4Dgczaww3qRcceMV4Vr+Y2wt0
ynOveIzLJClwB0qCwEyrLXRxeOItahGSpkj3Rw/I091/0ktHnOfzhsN6yo+hvYWHqOnn2cYMhe8w
gUecBVPNnvvzYp1B1YfxyrrZck7yihYopl9q8569acNgPFWc5T/ZdXtQGQZ0C2AfbPrgRLyHdaJr
tcJil7iL/eRYyMjaVqzuOuGcpElFcOvb7RuQm4TOKFuJpug7DZlBzMOugzsV4w4yNBQxZvCtZYn3
rnlRu7/ItYoQYJdbhO/TlUYYx5S8yfNBxiszbM3PY5SkgIX/BueWcX0xM3Fjvv95fDFnWegbFSbU
NbXiRriZYItD6hN5IMjRrAmMLcshxlKraGeKjfusEzfkii8sV/+ZQ2FgWbhj1PgvVsFFOJWSsNvr
RAUCbFjk/BY3ZvfqTzQWekANRh5v13oDJUTOUzNwQbdtSp2Y12AhEtNYLDM74CMWMDHjzjYdit3s
JXu+D6yBDTVkG/dipJG4DHs5ezPyz31CWD+bL0C5ZNO9+HkaXX9EOJj/ehlvGnnQww7X2uqZcdoe
fRe3LO/PFIlWO/+/ndu0YSH9+rVKvBkjWzjwtXkInPgQk46ZGWXgLbzgPtKkRqIuBM3w8+AQDqpS
RL4COkL6AIUHUKevomsGStCdYv82aU1CngHxNuTKbxe++OsHXL6upQcqoAY4vW3uyoS6QQz0JtjW
V/BbxEHXLW8cySvDSwzGI8dknwiq7CETEs1k2zslNPjqBpDdKMfoOHASlS+3fvrtPbVwTAbPpYri
ksy9LVgqv750PWURhj2Nof1q06HtlMsS6MuLRY7Zwh03ujdlqJD1kT/ZtUjTLy2te8q4Ce1YFrBx
2VKGI0jYIFP9g+nalDQLyQaoM98QW2Wz/0S8wl3K+mQJs9tNDcwaLzcDjG3ISudt5/9vz+4XOjuB
TjdgPRguhsqlBIs5TlHX3mUD39XkhclCk5rRkq6GAu12dGTX8+9cxiYCbsHf38IMzABj1KXY9Ps7
zLVlrR9usWKqbHKowJrdRFsILxltkzO30f160m25667gguMZi98hBHrGsI9YyJm5ggVEADrMlHjw
oxIlL7JFfwjfallhEmluIeRMfImnAnubCzpOv8DLw4sO1WhPUcZNrlUNxgyUzJAmpyH9kQJxj8CT
ylYyEGCYqumzBlmSPfFBpNffSfsn7vJ+8up5OtYx60V6UJhni91aTzaywTsd11k+8RD/SGUlLQhW
24a7Ln1w9HJsXQbOLG2Z685/HAJGwnsL8oa1T+40ePwfSH19lech/GKq16gpI8v1REcpw3Upl44G
eRGlF+6qpXidfnIhbALn2XF0qOjOpWOK/8etrXW9H+/ZmNs+7EmEh2fb7QROKNqa3vyMMjeI0UGJ
4x3lw7NMKs8TzG6uQonmz+DJmpxZf2skar4LybyjA1+bozWTfW3E+WZkoA/8XaO4vmZOXOZcFYth
w1/TO874n45nTXgt1310qF45AgTCktWAQgv03XJNkFol2SE2xEkAIeE9AB5plZgaYKg3bG6L2CYn
9vK//Y1m+VCv6+DbvHOI5d3rVZ/yUvslr5QASf1KWqgu45PS6PqFk04RRTxskvaDFXWvYfJuOX2H
3PLR6NB2q8DbQakeEloeoWsX3fhQpLykszxSIQ9uGEWudiFyFVS3LWPpmL0ii8xlRXG3F41TuZaJ
W5ybA2tNu35K+2rr35ZtJpGzjaRXFsPCaf0XaM48DRqGj3NKqwzMKwMpF/gWgOFwbKuk6T7FF1Hc
3deNVNkejHV+0kT9nrLUZBv7+Sgu5p5KVrPPU5bNVyxINOK7aC8EESmv1+lJMNNV7vGi475+TSsi
4WpD66E740fK6kujVsLtOkAPHgJitkIOE9O+X+GwSHWhO6EOBl1shEyxncho7K9S53kIxqjojKYJ
UIJfv/16+nKF6uDYh9SQeV5gsyFXI2N0OS//1mW/1k1FNup+OwjCb7jzRhyzo+sI+XmTiMnWOnZa
F8tAolgPTUVANKgblWMX2MkGbXVq67RNNi6AD3MqYkPq8Zxa3UbVTIucpN8iNo6dGJdrZXxO7xpi
o869BRmDazbQG+kjRAwMjpTNFXSyJe3+ndsfAcrQnmkb5tVbnFacpNd+SHZAfOHWjvU2i62Nsnp3
fJ3oxPn6o/fXFOPO8FFN7uzay11hf61DLEp0YbfKDscNGNDQZ0rdVIuCZCiOwNSKPbUKdzVnqmTW
uJzcv9NOlRUubpVPQx7ujrE9ljpcMYorrTINozIUnz4hBm+tmgvRQa1W5IwyTdv9hFg53UlNueQ0
aA6xC7M/isCSSnvBw53XDP++fiZAg1E52hmkQpxgAW0p7wgr1sAIkAF47rYkuMGtJ1szYF1zAJHh
Drq4VLHeMm8GQk2vsRHOS3Gygaq7zAA7ZLq47n+jOrzTbAWi5Yk8GZLnMVMn7KgwkYN+cuLo9wVS
xPOF/Hu6okv5ZK81Jj/inznglFqbETndT2coMW64XI2x6HlHtsZ/5IcWdLHemw2bOx4R1n0SDT8I
0xpH0Al4Kwpm9tfJIoBlcimXeOWYujuk/vrY2XfFBeTs/Xliv+4QEZRRvdFbNL0/yFSJg7mYyavA
qp+hUGsxTZwhGintHszOfKhOmrn1aSJCoTdHa+bgT23BHO4FDajpDDgeO0XO0Yz2RHXunEsFrPWN
MeVl0W3VXuzYuIew+AyX8mz/38ebfqjr1n5c+rTIurv3fVhg0N4AzWSco8e6aCmifavvREk4KyGS
SHL0mjDSqHiGX6cvkvcziKzLzdgjcuMad7dweS3PvgF6qgo70dXkgjPaqoxFLwnSh8OUQGSPQ6xK
Iq/h1FzfaDCF7Y9gH5gIVzrV6jmcnH7Lu83OcPGVVJ3LamntY+IvAbxmWUQcTHOKaDCUeGRW6Jwj
ujJPHjrcIGSXRNJbiyvmAA6qNOZA8mSrJzXLiikI+snlP0fjrfZEVr+z/yl/ogNgAZQIyEaKqeAp
baagUoFaCqEGthPu7nSf45tmy6wzm/Sqn4X8cHqSrieMMb9bC1UEAjk+ee0sfe4mO0g2DFYLaxXp
ccL9NJgGoUgZm2c837tR93p31Pzv5Hmv1UBfLrkGUMnE7uebS50xLeHWbPrgiUQIb9HxV/PmcNMk
xB+6840IO92Bkvv6RFeOUdYvBQVRXtAWUB6YU1FjGiNhWQ3Yf76kg9vW0GiaAog5JxMCAvskcvp/
JzeUxPE8CCQxQ0M04BQtKP3DdHytYPVMiuj6eTaVxVGdQ5OutQPNmKtKonBUxDRzzjtJ+mwgJpi1
mWlKb/lrSiN/sm/S/ApJAnv93djMlffl4GDOhJASfryEuxH5cXKtLSFikz/pZwob06x2YAmRMJSm
YqHmyWWknXgJpOGDmdA8XfGq9FSCP+/fNmue/EMsRrksixliLpYfVYTGLQ2qgrOc+iW8IJd2jTCK
xrN3mtdpT/2nh5MH1vYgqtyIbzSXJKdaUMLloQQotIUoTVH6xQEVUWxSWibtTAXiJnLZqnsOcEDo
WYdQnRSeQiRtuvS7wt7BeYaPEIyadCcxpXS0I2Xg7xlcEoauE2b2ZuJslRudu631dxiIq0pSFPWl
ju33haKTStYRZRdrAymwCUaDjX+rf9dIvxBRG9V9kVQuVd1o8t+Vrr5WwsVBYzCulqJ8V4mKsQoe
2cimS7HvzkoBr7YZNvEjQr/+GIl0zYoZxuwNiY4vBO8ucv8VsKxWA7xSC1ukVfQNrTykX4YXSrDz
Y/L5LO7FMM+7jaCfRpubohCNMDIjyaNxc9gndWosEB6Tv5VnXixAmG7B9YFN88cBJ5ur3xZTElAL
G5Dl4qISnTU75aD2gKnuTUMPla0FbxTZGoXk4NoiZv+hrlPOJmD+PxjxvpRjo3JGRo9eoi/Rla49
JfbcveJaehQFAQy89PzSFF7UmnypvBBFPLsTKMBSTdcI3dgAPKS8FOHvdPrXAzIOGQBfSsZ0UaLH
1Zwc/2bqrsEN/JOk8DUAYa+u62U4KIRg+ARf7aZm9z3shInUK5tDN+BZ3qihktvYigEJXRzhUVf1
UyVJQa0ZYNuPAlXcZ2YD9X2iRMNjCN0U3A+pUvVzZ5DA0aNM9nMaOkFKkjdDDi/4jTsiv8ho7g4m
7lVfz7Cvig+t9nOmoRp7pTsM9sSy26LVkvhzmBc/HeDElNxpgWNE8dHAubUEsii/E4gUAUHS8fZJ
etzqxok356OYjISBJkyKCM7nQj4TLrzmjp5On+fhIVdqsZjg/xNb+7gjCUW372hQCMxnyuWhWAse
9ut9ztqP4jFlcuBAcrXEau1U18KdsYHpc0f1VQZck1eF1HvnSQsaxS17GUXDExZdf3msHbthNcvV
kQMDFyv1BvvrIJeySArqXlohrZRKKHOs65BUkxAJ+JZfAWfEJrnEpGfgySGe66cLsUHQZAYIh+yh
bYhcxy0vDufimZ6rWvSVGLFo17oeeC+OsaA74nq4ttRGne8+xJcufKWSn1cAcXh9GzZSdkHVI6Cj
FM8Ewxg1sIQKAKBmpKOXhleh4A0Yvm1MNiPtpBzJWhcrdkW2OeccyrrsgNs/KmreJd7fKRu/mPrW
h4KLqxcC4QI+p1XyVqqUeOZtSbCX/GQFwItgRYB8/QqvIj5q+wrcQ0qTGO8lrYy25VhajIMrwUHr
S79YQ7Ky3BdsrM0c70NhGQ7RVoK9cQt4qNsVDoCEehqhxZkO7dBLDj/Hsg8/jL7lSV7NW4cZH3mW
VcMWblf1Z3VY4PYEfMOzIcNCinKwqSnvYDEQgxD5vUwE9seBqngWIPVom7Md1IQC8ps/KgeqpvzK
wVmjIPMg7XjP5AwM2EJBgJPQoI54iY9tkRVoI5bNTze17I3RH9kbVhZBGyJY7Znkr4yQeCO9EAmE
70MJ3B5rIzVeD+Ng8soohHDQnrFmF8+3wI422zVgbk/AWDI+lqNbUa8ODD7j/VPSn1UpFSlW41PG
0ut/SbPDZj3i9L8OjQrVa5j154jlSF5DGXjfUg5jrYI1jkRyNsEbv3xur61mhZhVR3PplkJnC65r
EjoZWyKRtgZhVcQPjBhdQuEDvbLxriXRnOEhh8UBFJh6rPbTrPzlC3Bbwl9FII30EvIPXYwQ/Mpg
kEwSroaYWWriG+xvvpXZN+mDpuMr72Zg2HPgn8kVG5ugxqf9VDdsHxmnwX6aKIgq+4TGX/1rqovi
jRbpj4Tp7XJGflJpLnM4d9+iIKNeibtt8EHD89AaT2AwqxLQVbYvGnrJq65t9mxrqrYRoRpgEe/K
eMfZEgunT/n21JudZDo3CA5+qmCigNwHMlnUKiCyjosvE972XWIIG4v+2uJZ6sGfNSf7OtL8NRwH
z0haA1X1IR0pFv7l7xmV4/rjhFfyFn//8NaD9q3C9p9uJZ+SP50MKlexbwM+1z6xlz5zkJIE1kPx
8kuS5XwZcP4s8Njhk3eu1sUaoRsPpWRcda68C0aEg9sYlRvQZBciNHbfVwM7hMSAG+qE/NTzJik2
k6E+j0D1/iAxKUYh11kZGM40gbgClJBDM1oEe7dzplZnxxE+wQu/ef286lSZOSftO2QL+7yKKhIh
iJVBoU0rfS562egP/eY4Ycrnylryl4BHQDu40GwHAthZrFnSkP0LB1MYq0qyU3E+1tgLIiLbL6Nl
J4Kz+6RUAPC6ccy6MK8GNSJGq1ZGowb1jvXhFjMUMGO/9KSYXdjPoBItOy4uLBkeexjDuorhoPQ/
kr/R0eXNwkpcNB/8CjlyuiM5znvA++bfXoOyB2kVCg3srHsBJWtk+ty2p/scHwr11Vd2Nmfz7YmT
boRLhkGUGSsdqbu9zjkrqJZWSrb1Qvwh+o7CK/WyTHwb1jk72lpBdfbrKLz4kGouSom+j78tNpW8
sOG/NNLpU8nsAjilxIcLb69HjcCABgtj1o5PcGW/nsebhzaLpbwBuJYmRhm2uXVHtcNAQ3ld+rZY
iC4UWJ9YMkYICnsTtgMhotK3PJ+zfUtKJMgxrlQ4Lxxhvxt//IAY+AHKwPsQvVlQdqV9UMSRFlje
UbkBNH2Rni/l/qPbf8eZoyVora4pde66ovX1xlDCxbBVWM60dNTwIt5vEUJ/IcLe7GiQ/DGd08IC
nMf4qQSXQLtffDTkDuHChEiroLKrILccOumo64b4vOE+blRdQ3czkjdXLlA2ff0A0RHMke+urSP8
gXzUYd6L0jdxWgcnWm5+i23B/6CFUYDcoHpI6wYU8IvFtCsT/OynlqOr+hTopn7S0Vi/TTeCOKA/
7OzU9IxvnJ67aa1lna+aSWurOzt4FD1PgDP1hOMTSUddt3h2L3lNPy0eNnzenQ1wn+XCx+BBzoet
nLljWk1AxlhDpmQWsR2bpPNVBNOMdUP9iG323x1FxlrEYxbn3FlW0SaKyCJiR1LYQNKFGP6zwBYG
aIpoCsLTsaI2oseQKQQh+dh/EOtqq/n8gjWUElEwGXyGkGm7ucPRH3y8iljOfnNOaEc49NmgLB/E
VOH49MXooRvqZ0eSMGjtNKzkhmXBbAaN2JsitY6xvtqL3kmxn2SIN/yMFMwmHtpmWTA81tmemTlW
G9KjuKI+sceaYCyb7uBCNvNXXihzwvtQX9cWoP4zDmie2JTUh9ekwTRDjKOxLgDNqoY3c+FdCxVm
ZQep3T8L05L8wRfLafP0xOn3BVrOJ9qb4/r2Tweml/Bl2tYmXKfgIKaQQN1oqffoFK/dqNx8+6Bv
m5aRyCDc830RzXnBpZy7jDGWd1m5P1uYiYAPlXirliaPWBuj/xypH+Xzy0s8oUQDdTYWrE+3EQcb
hivijnBWrN8ZDXd66anmH/gHMCvL3ZHWRhbhrPUi+brgdQJ8hhTTBaE5YiMrS/IOPZLRYU1/6/3+
7kcgvaxpayq/+8sp+zjWDNsp31zocs7OpgGq77GsP1+57Hn88RsKE/OWfwTpDpI0YN6hJ6WCQ7hg
dilri9cMRD//GfeMyUMdWYBKBH8amb01pgNzeXK8+XjX7bKRlKBMJOmL0ytbcQv+hWLnM63f+UBE
ut1lW+DWBmPdDXSbIRM3qHEfu/Lm125rhul20UlJyQt/d/FcLJvtMdkt7s7kViTfVFs8IR64q9Oe
BrU7RCdzHA1fwnKxq1SbRop4l1/1iEKr+Nf/Gf+wbnDerVa58ZTMw5uAlTUi5RFL6pfQkceHD9wY
upzdHspwdDt+tjHR4YwDFgbghNE80XiS+lbHy+tnOttxEsw92KG9O4RYhEcJdvm25CjIzPTeboc3
QkcpYEZux3fGjjQaW5e4qP6LgkUtzwPjomaLqwn1pSUqOQ3srWfbqRqBoYe8/eDPvDNF1ds8qRpk
pVOanY2O/d1CIXiAsHo1mEN4pIcw/agFbh9AB1pfHjnDHuN8j+gYMc1DOjE7b8+BjesnKWSiUx8O
OYxT0xy5/pWOebmCAHc0skSNip7IrhOb1QTwI2gxsNDiIvlaKK3GRLEazkXwiAf8YgUUHH6Otmqf
gPKfhUEwOcFcD2N4xQhDPyjJjs/oxamEEpnhFII3HT+Zi5zXrPTZ+9bX/5MVVxqOrkU6G5I/w9No
k0vHjGdMlkZnNS/2Cs8s86Wp6xOl7YCocQSPvDo9aUBH1KDI9ZF3gezuEPMxLmt817VzYYC5DZpn
+fZjfWiV6f/BlxfIj1IIyOknsRJLsUz8RXjRiAwsGMlXIL0/ObtRZ9QaDzlXZPVlY6Qc4ordQhSp
V1H3bFGMcg91i6/T9u1a6guUuIr+Mq+OwQzTXIPsBG13h1qiZOsF1xJcgGvZ9mLCBHDQXnkM4OXn
jO1gyDDvl2Tmp6hcMmstVsTe+rUxjF5iHZOqOHsGis8gf4YT18tmgwkj3q3OqDdD+FFLcZE6fR4T
CQ4jg9y155SpbPyfnbpLj1ArN/pDy8kQOyK7NRZY33pXMyvlo+rt8zTLVstlY+LLmk4Ao1t5NtIG
lIwBDIvGMyKndwFhd8Iy035/ahvMmPiUN1GiBMjPvYMToZb1M5VMnPCi0AIZJSKnOFsJ99WOK4kh
iQLsyOC7m9u0b9lPrjoMcFtJRsuFibSbQWBBvBpDcB6htK8RJHB9+Ds9kML4l7O9FTcOymBn2Jdz
3RxkrJBBBpOQMQ79oyf27RocJ6SJcLYxdUrD9I85OdtgUfbRKcdeq6Qr0l/UWdDvUNCnzwxiI9rb
C22I96mGjTdaNqeiZeq60yqESn8Dgaq93t2BmgOFPBQuIJO1F/EW9zuuFaln+d3/rw+S8ppI4TjM
h9I+dLmjCuukl+Lf3eokBX9eB2VhYqSqQh4elN62ZbW/6aZdaq4nP8u11w6bmC8pffCLKhk0MZoh
4d1LqFzXsQP0LeVLFR9wSrGHfOUDip/3Dsx4aWR6AjVutdP7UfOoBqPXSi6SVMMMksxluQ/eOsaE
CwWRISM/23gxJ0oQjIK1Fev3nbUNWJXuubqwyoLIccON7tARLbFxLPj1aNn1oJ0WitOfH9djD5d4
aTrQ9wGt3gRoHqy1bm0aSAA0HAifbNvjE6AMoDxs5YOCGZIMSk0sZA04axWBAuXuCfhsNPLEDbvX
O/R0BDHSe8u+OxR98pQje7ROfeyk50XwEeL5sAXPWLiFqxbBj8GGRqhnwKpkWcpx/uIS9gpNGV69
BkkzAlPYbnnuiaeWw2ofIP6F/HP6MYJmtoxqoeDHREsZmmOcppGYS3ju4Rr6J5Oq88XxDohd4KpP
hCb8djcHabXZwdKCVHq2HX4r8zWA3N4Kz8hIQ8/DOa7VMai79kfm8TMoDxayKErrsES3J5koDNFv
xXNeQO2kpW4qi3sbdkKm7eZtiR/ApJYv2qWQfGbt0/A6XqwUFriRC66E/itgcAKXuBGgppCl+4IX
oeaMuRf5MYuCSOPSsDljx9qzosIhjaWK30ye/K/XdG6d7MCZeI0jfR3vXaWHZ/2WuddqYIFWM6/g
kqdnvrnT6Y33ziU9sauTW/XTXCqa8s8cTjK90uAdYmiu3J9CeidmQSwRbiXtrXCSInkyiT3oSH0M
mdvQmaGtD2lKtVGLKHb+1CPQrplJCl5fRlsz4VN9K4voESrYAmDnSagvrL4vkbLpck+5E3l03ZqQ
6jFOoqLciw5+m9PIaUI0g1w+9/TDOHvTLJka69vIKXbrN1YswMqrAUGlt93iBWletveeR+CoaDnl
EoV1Jy1X1yOMcunXzAlsYqg3WNX9Jy0/MF/zdXhaQBeX2qoKKxlIxoa0d3YWWWQlU5p0CwTi0cEO
rQmMbiw3fV8RL6FsVgctD+FiAZJrI18oGf9fjBCZ76/LDrRaauu6lDAecPMfGhWFIN8n4XXictsG
OqMeNCuVS13KA2cRhR3ZYbIjWyGmBapFSQ3rU6k2SQ7+0nsEkMfTwJ2wHmS6ULPiXwlFhqpSQImE
ak3vZpfTq8TMz6ch3JgZNfmyOoLYVl2v1M5iJ4pjH79pyG5Wb2DnsNUMZRZhaIPxPyWrfh4Rw2Tj
qKRAwBRWOOZEr478Mj2tF0nXYalFA+lVQDf2W5yQ+pOtsj5e2DS+Lq1xtWAcixXP9PsXIohCR6a1
F7p/uS+5VLHN8FyLlhPdeYTCVufhSXGHATDXoIfQm3Jdw12Ho4D8pO/gsTMnzW2im+QaxKvC+Jzf
h95FIm3xOuP86x553V2Zzp36QHSzeewf8/ajJJwXOqp4LhS1zC5QLAVqlRbhfThxnvIQQQNRXpvR
FUfezYnX93lKHSgY6Iwoo04r4gkvgmO60FJbOVcoFBHxHNilcs7QMlBOwxVvYDvdww7E2bPoTS29
VlZTj+30M0ONzEP1g7RZGRmlnMdsnMdq3uhAPC6HUzqvD9mfIu3rOq4C024g5geM75qJihKXjBLK
zZrotcEIvjBb4YfRrK160l9TLdrrUfwcu1/q1J44Kx/yRStkh1+zXqgrnwCDi8wEtNzryCJZFO94
DZ00D+ArCqFioYrPozw93GKWaVyig2u5WfPywV+zDwVl86hYQ63yMlb1quTwBo5+2RMS3ecQvxxL
NfPiGv2P5Gq5vZ9VfTI8eHlyYZStaGnQM8FTaEeGGdxM2VCuNbYyplZq4HDuHckYMspYuvrinysn
PdjwaE/Ubn3DNbqkSaqeLdJj0r95pj7gBRLePtaG0b/GTU02RKJNEyf7DwPUQRiy8u8pZ6dNdG73
TvKye8VmTNz8t0GjlEc+tejBl3FeV3qBqeuGhbg9gGjL+ZZPZQmmud/7iYaKDzYpF5zQ8bkah1hi
uNPtymOuqLKqJwrd8gR7ZEnDizlBY025DjJaZcB4stjJOF8EZhBa1aoGKOV5nebMeyiGX4BbTCFm
4BCTUUHTTryX3aL6CCthnFG+Z+S49bv6X2y7QxQQ8NPrQWiNHpTusg3mh5jwrgzEYyWSapAJNCHs
k3qi4W5u66qcOGBBYR3vf3Tnb6cu60qDbXsjGMrFo55DfyYhqEeBNzcRpSf1+DYzDx4EIvvtX8pF
q/Z2bgBlnSTDjF9SaK3FKgn4wRqQEi/3BW0NYocJtOmknGsjHtqTAbF+DK+foTALjRg68FovP985
5z6ckIlTQRYSxXOhJ8OA+hd/5bQ3VZ6kJut9VYhHliOFt6N27eQ1/HdmnLnNw3tCIFIvXlT9v7v6
6xAn7b3UTlvIKZZvsikvIB4rqOSFCm28jK9zy5RvPERDNK7mVNfFxNwTFAaJL7iGfOTqTYDMTVqx
AXv+dcShELtlrafZCL6SzWfDStplMU40pHIu1Tju6fbeMaWe2pIDmmAEhJfXv0lgmiyT2PUtUcD4
NWO5Y3QizO4nDI2CSomAXroupfeNkhdyFz9ip1ONQ4xtes3xPoe7zo6dVqNGstLM+HSWIUcuVNOF
vzEjVgBlysEivwMIQ1djN+ZDnyYl2NllKAXT8/Y94Tj/vwPUPrcdWxznyfvYZSxUIwufbW6HX23e
rbnrY1X8yQ/bIHdzhKWuFijKD6RDI0xDSIdoNDHwkdRXpx0636zyCpR/ZrK3o3BaRCGzWRqZgNIZ
nDOnARWeXRrZlIlmI0hyD9qteIGN0u7cC9hgg7HILz/QEioLdayBlRZ1x9Ap/FwVKVWrsxngSFLA
xje2OpV4LMP33EgL0kjeHoTI7Vy01MjP3NEqKv9Cgkt6x0lqmlucgaAR0xEKsdk3ZX8PAqfBJWSh
m5KVbefT2erod6oZWhmD0JrQD8sr6zXMx8pBnWeHWNX1KqcQjcXgFrlZG8clfNYD+VW/KxVcQ7mF
RF7r1u/904a1+C8F2mLpqMa9EXdHvgBromBvD6Up0GMpqIOTAEemPznDcwqrNKWz9kjOis7fTkRF
UW7ao+2zdWFn3tYS/S+uLJOC5asNZbts7Bx0e2t6vNF7Gam9Fed8r0s6Dpe7Xpv41so+n129XhDs
i7/Gt0PciSwz1EtVX6gyJ7mSsla8EjH6H71FdZ6CEKNtcf/VUbgqYOFq6IFSCZSzPJX6t/OF2DG2
V9tz/rrOD4wUghhFZDqZ+D4VE1La0ghVfnM/2HFp4EG8gJ6FsjWYDpb1m6R6SQXIhfEg4Yr/syCS
5b/tYEteFd1tX0OIKoTIzslg2Q65a6kpz1/BovrfYqMljUyAAWLovRGPziM/28xMBGS43QuetuGR
OWlgH8UEaPzKTAwNOUX7y+16Wogex8Awm8DYQo4f/BSulHK1GWUqqqfMccMiKcSf6XkTbRlL+DIp
TU87j2gaDY69dG/TW01ZrDfgdkUg32FJu13aww7uvBBGdJf+HEpSx38B99Ud3W+5CAIskmKfKTpL
9BzMvfOTRAM9floaXd+z6XSlvSG3nBE+OpPduIhgHrDzj6NHbAVml/disuxCQ9u+4C2YS2wt3er7
tXk0XaINKLEEVW1JdIKEO6qbovjBr/z9WodZ2Yi79vlWtr9jxz6ll0l+UYOn/UMePR8+UebchcYE
nMK3U6jMAvlAeml2Sq6O4i4mH3MstLFBikNRLg1DrzpmjWnjhlHkC1FGV9jN95bRzwY72JV3UYF0
t3rjc6UHFnjuCLA3IqrWLH63qpMB1nJynuKkWDsQ6gzXYr8G8B+5bJAFvhAu7jrE+LxVMxv5sdwW
2czy/49NHSbn0JTBRHf4bu72X34msPwR15PQWC7FPM06SWeLGFK1LRLkOqJoA9J/OV/vYni94gFn
nbtXRqhRK6JFXLeCvZHHNJ92aJkhOAeTP26r3/MLG8p6zNkdr8D+RTmdXhMcKSmQwc+umxqYvu7f
1MTzY8s6PT+Jt5rk+/+BC8k0NBipUSFD1FcaMEv2k/zIIrHYHteU+Y2JEt9bDkTeNhVyZux+4xoJ
DVPZPBTlUfh36zHiq27fX52PmStrxMMdnBAtb7kD91sQYPphkfh22nMrbFEVq8ds9phc788IFfjQ
FC8bvmuBgN6OUARu+Uq2LGZgLerqbTbV7ahxexVYyKep0FAMgZpJkS/8D2v3/+krItgdsa04LrFI
TWhsGDi1NGvcKXdnrTCzYrBq6pOt2TXVOdfpmnkhpo8CJbd0MFGkYSKJWew5WHyL9xGeOJXAl1uP
NtiqJKj3R5r6DeADCKbZJkA17zS+BMT92qA/lg94h6yxLB43YmpMZtF/lKbjneEFVBisHp190nIK
2ehrTUM43DJLRwT8m3o/CD4/g3Ys7qurBAY+XZXE8tuAgxkHn47LgH3B0ND/jZ6iQWNgm6Hyrl2m
lUyogL8NSUyrZL/5JtBImyjzuPU2EUBi6jvWtUwBfo+hgzm9dZF1kiV1edJdEtXlzqC1lO2p9dJT
4uPSzacPyPo7vHxVe2xaaBJODI911eHbdYIwoqcljdSZ9+cWPzDvmcwkLBf9kvCvP8K4OAKbvLM5
A9jSkIEMUAfXlqL8JIpvX4+s96mPzZhEb63NoNkid+D2Nyribimxg5WppjNHYYgUT7PJzQMl15J9
NIDHPO7+2aTv6Y6s7umFZTjtShR/TtZSuKIEq0J84VE9LTaRAtswScYAXB7WCBq3O2SfuHr8tQzk
sL80ZupX4YDnwIri+NrY+zuqdOHoDvOgh9lwqPS/NS/NCoMsZdju90BoQCfQRuYs3VjtC/aqWz5N
HJE8DtwTc+DKNwgy+YAFV8oYPLdCA6W+EMTvTkpjTnQBf+VIQNAHMLEkwO4wONbDAGj4jEomiZ3i
WGeZW8rcaB9rw6qWMhUZtwN06tUYLt4Nf6i4nZsjC5mUBlJ8yf83X57gQzQfEaNvCAQcTmEZ6G+o
Z5Tt2dj9V8KKHX+IXvRfFjfyey1fDnZOKYTGghZo0QZcVZ83BZCuOFiOwxQnjvUUEkYWNzbvdAld
iX8K/jkpR7rAm97lG3sX8PEclxkqkG28jzdyAoleCsuEzrFx4ccLmPpEnORk0gO4mmMvr0So2GXn
y6xmhNkQjubduQiSQU+FVoc9E4cYcTxyVfzNWB/X2fZsfuoXOPN8wJxMw3/eJyEgP//tYOAuDLKq
McHb5fufxvRz+2Bl8L3KzUufn3bVoXOsyIL+t0qYT0EoacWnAOTPPrf0JWo32K5DoIEtYs2YcHM5
xIdZZjNwb2orrhfsmahyGi1BbGQK+mDS55KV1ajsAx4HxtVKw0AdSUhHgJuIcijUMOMZw8DDm7cu
RlT/ZXErunrdFLWOuL0+5GsoIpRU7p6xIi2Ms5mTrkfaoN8XUlkyEVCZ/R2yvYWh1WoX9QPsnN7n
UFgKO4zTWac7WHFdnohNF5X+4w7DWtr17jQQ6AcYhuOeTHDhCBnvnSefWMXWg3TKf8UqgFKB231V
67lc5VmeYggI6IxBVn6SG1Vii9/vLicD9xB/IsyiyZPmme7M5ZVMC7M3z686fyl5oWWVC6rAtiBT
cIZzt8QDYwae0dG6jCLn3bngJ9dKQEUOe65JE+QmxGCSepUDcLKHUVJtVuLIEE4+xgCCeEXFiWaC
D6f8bSKmIhEv0iAtf58SNqotVGSRGcdzyrdoDAQkNLRKA+5MbDGuC5JnCa+t/OEa0vn5FzOPrOsF
SzdNm8zhV0rOjicRB/UwIaHpfps99dvelJyG0RwzqlSMAXUIDobkhWRARHJZ3f9/4iik87VoekZc
qWGWhBuNLlWzFzpG3FCaSafK/rYy/ChoYyvTzNnjeKaNNx8mnq2dHeqmlk7JZ+fAl0RKDnt/HN9o
R7pw2e/64vs9lfoQ1iVgpo+s4KBaXdm0xnBefH9mZVUhjDaQamxXyfHz1H1Dwsf8YsinkIXsiyep
n9oJYKj39Upg++OmoF+QkfFo9n2qUqhjhXRURUtLoJzxv0pbQNq8HhCppeOQA1qylfhQBQHgGPd5
z/t1IuhbOPjd4mSVl+8hIJpBdwuGNpCLm2DXXvn2INON59wjC1/jl6noz6nFTHiJrc5Sh5jw8FKt
EBwKVwW1aN+yPldt6to+OPJWb5CHTJxNmSiYSTJxt91/nfUY7UdTegR5XgVRzC9LHOHN0d08KnoG
vxKcrkAJFhas4mCB2yot/3jQlp5nAlPmfiPqa+HIHW0rwYOoUmJ/n27oSwOkxodoZZ+xoyuftcs0
5ZsMyhAyip5m44IwPWHOSRXgggu1cHcEjr5Cm8UK4aFh9gSs1qJvyBXlrwBWbdTkNbk4d8Kx34W5
g5mYZL/HRe6TQGoSWxY92QqqFiwdZIaVot36ZEUqZjLsCi1Y1DNDw+Bnw5JfzFwJPYUaIS66wh/V
mZOIfHMOxktNL8gBRwioaORwrBwZxRuHGp0DamrF/Dmh0MA1zQQfwCLvrz15QCrU3SuBDrhWsgu6
u5FmyL2WFMG8UorNgOIgWLLAquGPXdKqS0jpy947XOJT1gbMyrYyjqBgCN73t/ug1jU+svqZrdkd
7ZY+P87lRZ/PsIK2J4XxJeUzDvc9gm/WeerRT73T4CdhHNEteTmmitRUoDtAm+8L2SL228owJ6dZ
0lR+cwIxSFFGRWqXMcY7FzAMVjOuNHmAfnMF9S3OBX41xNi5jJbd85yNu9DEf7HrB4ck1WSoEHb4
YZv5LFbDb04245AVmqJzsXsPYYBx9/QDB9yHq9A/6gj0AC7qMx1/o43kjqi29CHA4vTp92QEADkU
WJuj1mlvUYr0ZMOTSEN/113OWLFzrZBotaTM7IT1UoThBgC1tCC9bxIIY5aaGOmoU79TtKNp+2T2
e8YXg38w53OOr8pV/j45WyYLdSFIKWLxERDISBBKsvuWU1A+tI3dOCWT3G+1kihpsloQODFfMIRQ
z2TjYPiaUdEZgNIIBpTBw6gp3ZKPQwuzLGRBqyeB01LQCflaFQ9MvqsfurpturvIFgz9l/vKuKK6
AUv/juDpfNBYn1lSYWWb4h3yt9Pr4EhJilf7R8eVADXD3IQQRJHWj8IDrCuD/c/GFO9/24NKsNAI
nsnTT7YaU66oZjZhwshTczgFtS7SZkei9mV/jOtelsL2AZrroGhaMrjzQ8gbPiMMIJ/gQGtXyawl
RSqwMyuEmYsTcvY+vZj5JW3241t+GRqmMg+mnFSgszpa0RP4ZQrQfA9IS+V4lBckoJ2Sb96TwP3L
TRSQGCKwdI06F7AOzcq1a1fj6nciNX4KprGZFLKterJyOlN2fjnKqqkbpcZrcDKi8rRJHoGQXLri
5IQFSR5bWGWOJYbCnIhyzDAdVqpGLTaAy3rtGV2ZjzMQiHO3FAg37J6YkpQSYxFy/qqUlN2U1cqp
TjDHZkk3M+oHtTnu5bRmbvdoHpttkpojlGRj7ZEk2VgZ1zb2/BsCze3wzs3xrf3B98RrPaZS+wCH
lV6yPjZlVF/d9aWC0TkupJvK4bOzPJA9yRxVuIlnKtrLk387wWkBVwpBo7VqINz9DxKwIyr03zcn
aWRuhOkzHhgO72b2WW9hLtpe/qmZEGC7uVao+KN7ubmtoHZWSzrOLz2zRrgz6dE5q+zDO/q6Jdan
Quge6prY2BnnaVmwq/vSvP28HOUTKmQSrKNxQTRsU2OecfoLfTGDItLtkQHGmZXbCrw9c8Qv2zk3
73qA1Uc9gXfdEsoozPqIVu1azzihFNyOoFPfWFLLMHY87mqjx835vyh24PoCcx9hnihAu50EyQSy
6+2LDct9Q+9Kl5xUVMpON5Fk6NUDzNUZzB3ShPm0Yghi6gjRUP1TlN6iG5AEP4frL0zLbZXfjITu
K0tNC7Yn2sNH/VS0O/nT+Wk6FEOaj0YExndpnA8ExQU7T5VBCSXzROVPKrHc3UwbloAg3BW4Fqiy
Zr2xb+6ab4spm+FCiH6UJeCR+QB9wjzAzwuT3tEYhgMapdsbqOxlY8EMvyJev844Ih7UEqgUaN9a
F9DpyBf38iZidog+HtWiPhd9mBd7rADX8JEPPFc8n9ICx+ouSTfki2/1/dxhqiGTh59CJuSCMPL4
wsrxj+iisc//d+eiXi/9+0QPyj3aPHi5PAs4BRcCHss+EZ9tDVXnE/yZweeX/sEtSKQhQ2s0FW26
o4+LAkZP79GKnjVKKuAF3BFOWlyy8ewbMRcHgBYuT9Zq5Re2EklWEg4bQ+xnbv5H6MbtP571cfkt
/gOhcauekxKxZGE1PB4PgG+DC8upcJ4P5wxR3qlEz4wldfs+I1i2KI1b25dlyeGa830/qpVS81Ui
BpGTm+J1QYZJpqn99FdMHW1+84IYPBqY/2lDlaNA7KOtQOceIUfQBFCfJEDXbhcHEWro6SCXZqU2
vDZpNXK5XEx6fV7ERRr32HXt8fQTnXNcyyjt5MWlo2iLysCDoDtDs1kuWQhPnjNQO//lJnyojI94
tGtZ9LGv5/T/7/p9FQrb7H0TI9ukxZ5MGOI7cymp/1r1L11WbFjlszaw7cEJMVxXCvqD+u2fRsvF
EkY5UdrXfICk6hDOTeEhp9w1OAr0bQRmURpSl0a87oHb4HjaE7qtSaQ5v7dVh1pIESZ9zeL1iNLF
riSm1DAacVtotjkEw31Nb7VVPzSU2vEjDPT8BgqH1OZiK7aMDR0TsCGzOLohzmaR4/QF8vKPLzCP
TbxtZTgZHSvr2MbFGdY+5235dangAgWhPrjZpt4XA2/joZTzoGrPNtE1TvgPvy89HcT37v4z2B+i
5KvbCGFWBeCvzMmHorwNed7OSXrkeE8RV52ouYT2SpYsgzh0wEjBPQku8AzJQgLIJzr4O5i1NS7O
ElsysXiGCy7URrAupiAiVdOMX2i5P43xspojA+c27g0N99hyexbS4i/FwqOx/iJugHinUkv5uhy9
ozkAeSPKPfQvOQ0d0XADTkrOdkVmpXJHZsJYgEcX8ooT0y5e03t0sEyrMVVQt8u4EFq/7P5aRhM/
VjqCV6CrvPa499fPlcT73lLXm+3ojqUCX8eIScQNG5sTCMRqEhlcDQGn/czYa8vA3s9lQy09MceF
+SZUxXzWP6/q0JFJ3Z8mJBD63HjByrLJEH+9NcxtbcaxAl2pifoQKUuifSG48Yda9eBKa8/VFGWb
azCmvK7Khie+VHS0M1KpSu1c81rOVdjlJZmBzb+l5ytIW7/dTLHmI75nEicUdf5oOO5ZMmyTtUFa
g1Gus6GO0XlLD0WWvRnt6jaBqG+JS7B1cP2w+I3q+658TztFkGuFvrLmkYBNCdRww12SVwi7nKiD
2DXPCEsHFlnNDJ+a24eKxlM08yz1bB0Y4LvWuLaPJjfni0Xx8v8qFqprxS0Q0qxy1wuYYWKZw3B2
mEtRoqlH3YCv3TW6AtZydpro3TJviDNn+UvBO7ohNTHOa6vdW+bz1NEQ0e2U9LTsp3hnk/5lJhm4
Ki5p+G4eKUcpxjae4rG7R0trKLhn0DvMwG5skDdp15dNKXlmcbOnAXE7a8qrJt07E9/NdrDayDIW
C5Q57eGWi+43qxafFe3H7vtxGIlcLUBj0SjvSP/srLlNb3M/JIKhXKzd6XnOlxBa7Bx4ad01UBTF
r73ciWm+uaMCg2lwYZxG1u5byO0sU+nOw2vX3B3wpRuWm0q5zzGKpU8nI+unbL1tddq5Iu+xnRe3
pY1RrDs7mdfuPsh+0m1tZ58nHLXHyQtreYXOKowc5dBqFkBqDxW5FSpM/B6q1wHLXGrfIXVkcBcL
n2bNs+PZ3xbrfwq5hzFEVK/dfCkRBXQJJZnV6k8iEjZG5Ac8uZCLPDMGOBsw5toTFf42TcU09gzI
+1j1Q7UGUl3ZXJAKNxlq11sUdrOEahE9hSaG0f0wrU/nMlqYOIo1GTBO2Fsf44NOoFNp096msH+w
/abxJq2re8Taem8D/Sv1oAltcgo4ATLcZlA/8ViytWvrwTPLbJd18gL68sIAxVFNTeSehSYpZ+tk
/FwKmoT4Cnlvg8E1qRInRFkMh1jjUcb31Zs035wdesTsCq6tcET20wrx/faoAsSsnd4GI5GM58Zg
hUDugrn5BJ0fRyfJycankAL1ePaVD+p2cVqgmRfL3oXvIdF5uPcUmXhxPXVLRXFkU6ssBQrLTcyN
3UZ2m/glLz/E7QdtggZOYjhcCX3lsSYevTvOJhi++HBz+6XmYoKMiMd3+yXp2ITFlRteukBP9w+b
iEA2Xrsu0LMtzZj8tDAhXt9GEZUWJ+Icn/H6myKn3JKZzcUzbgbfwfKgbfIteMMXS912PrV+xUzA
OZInP6OBm7Pux57w2goL4w2EQm9UgkNZbM8cQ9NV7ZOyzxpCaGA23CvnZRspjNOK88SitE190MeS
bAzdIqUxmziNQkzxgEQ80XS1FhcMpTDmytnAnC/CchKfmP8LNyiaVKlVCxNmduYi6fTZ4MwXedCY
6tlpwidfhrLHNqnoA/ugCgxN8P29G2/kKI9wA5Vl/Ntd46YCzvysXBoNCVxNHnIqngqmJ6fTYPxj
JYVjLX+5AU22PswAUfapS+erHFGY3iD19u1LK1agEllIP+svrqBYsCryFOgxIdP1xnsUe563lmr1
TdgA19yzpVA527QK7FLvEPYAExniLWaQ5HKMnBieRpCZacvxXoJZ3/f7nSnjFKIyVLN/yoVcpa1y
LBra1DP7GViTsqJ+b5AfdTl9AMHUPYuDUKcjb5IxkWddW7AoAbdao6jsJp8/HCNqVdFRlN5qQxu2
ln+Xl2uk8GhZh1eLoU3rCS4e2vtICHGTA66GUT5Q9U+eb+Hl7s9dOjK+rn1bKxtwkmbuKIctdYAb
SEheuhHjmtdUafZoyneccSKCGWDG1ucwnTX7s9r5xZN7G13qs/L+5TeuHuFo4lboQc7fQT+fY2ho
qmpnttR9D5EIIAupoc4kwm6uf2FB69QAEdgN9moWqHOMGcMxhYnx2IwllUVmJhAzPWdt/BcmeHD3
x3KCJRSgXxfK8GkN421cBxjxdflgnmdaG3eDiJilk9fsMHUD3TCDse7jLvF2wdNk51uZ2HqOkwJn
RlmxktP/M1ujoKYi4nwtnLzkS4JqGvlmvxOLzvks5A/MulZ32li1hIzu8nFPhhLzr2ZBJH1Ju8pu
AjW1l766ooYvz1wwpriU1cP+iOi+ejHOBUgpR59+CEljbzHl1HBHdG97Xxpc2wGoa6x3K14ktGqd
kKdwRrYbnEvDTcFKSQbZMIBgE2DtklzkM5HIaL2S0os7ljx5nx39y0YP97CvpGFVbAdUXQRnilo4
ch6qFGpsfyzh8ImskjAnBeVIMWwKPqBnZgd7zePgieYHXTPG+35pR5TvVzBr+odMm4nwUeDfbhfa
rh9hyp/FL46VaNsW8peC0BxAYChidd6NWxvx0BOCGV9O4sAbwnzJx6qNl4CVo/Wal7PazLpMBR0z
ceBhbU+cC3vxSmcFcWlom6pJtTlO8T9qxTx4YU1KxVuqzk0TKxO8J4MbRsCsHdI9OnOO5HGuc5HH
z81WLh0+yZcWtc2akEjrr6UHNucCVBCX4Y3jRqfeptRNsocpoyjb1SO8pvxTzKO0gqh1DCn9Z7fP
oCMuHFrKAiBZICTY0vivmVvM53XEPcsgNA2bTsxGb0cJd7LI/CJVVUvw3k3L5/iMM3ByQ3vq/w3N
JJv1LPDl7P6ZNeFwa1/tudgU//mMkdLC/g/6pV4qT7q+Xbqyui3EguIxx+Q03FYwNUnFj+sYKh4l
u5mdCI2eltslRMLQ2u+rnCt2GlUaPyxH8P56qfAKsYKx9aFZTFfV08rlthb5ujVYOyYUA/q7EN4C
w+vT7HpBkgGyBhNUGbs3T8RqzcY6hQ4PkyL/3Wi8rAK/VCy0i4280mbE0EnrXnx+F1QGpVJD+oxK
wOu1yCLNcAX9wU1yNcLyWnQ3Oh7UUxFyHMpO8sffUYWHrakX8hXSymE5PLyfBT4XtaZGZJnAScGG
HKfNi5Cd65aS2UdTdMtkuHqTA6kGVzLj//bwGm/tFC0ntINeSTAAF00YlAkEhY2GSL4xauJ73xtg
glLJoz8TYlcasr+9QKHdd4L+u+nsWN9AZHreV18rkQq8RC2wVSF4hqssoL016jutf/S7jDlfxlcD
s5R7oO1R+aYMXjFvtcK15ygki8DSRjMGUQqTlR1hXdraHdb9A0ixoodUAuDDLKDmlExg4IOoQtrJ
PRgIitsAjPhN9astD2DTcGX9VYGwOK3TG8a8S9WYnQCL3vqpUfLe3+M6hihNh62lBMXlLfciifiP
myDIupPpm3AK9MbYaBThRri26TSwrrzbhdvygHUoalYzl/OMsqfYnryOyMy5WRPmqM6xaA3gucOP
Z/dY9GlHdpshXCheoVkhsi1iZKhjiwMPXgIXcc99wg1bzzONu9lRx6yVLqjTfKVTS1j+yUFdjEU6
dR4c2ZU0SC3HyQ4LgK4lKM8ZiP6ew6HGNSBScb4aQWN4DS5zHpanby4gfY8QagLeiYj0FJ3AwkXI
EzGru/vMVqmkRF23tNF3cvlXqodV/oxZnbyJgf34jk/sBmJxzvzjtkWnkmhUMslDyWmuy6yR7Xlz
YdDTkL3B1lVQkH+d185TURzghltuJhXdYUjtzTYXvWtWr9LqG1dz5QL0wH7xZN486IKu2tbm7HM7
1ErsQd7ZUYShWuDyzqwyWonb5BuDvdl6BIpVMwJuQ7AjJwjcYBITWBUhwpe3qqrJRJ0Ny9/RLWle
J6A2mpyKUOl4SiHUa9IbBgjlZ5O16EC1htNd8u8/8qBs5gTGzWeqTyrjk6n/B1N87pI8Er01PADD
3BngucY2k5fd89Vt5+sVlNIBx+eJxLP8IKNVY9upTAZ7IJgbT7uLu02l/V9JKhqnvVg7RAAXQE6N
YT4B41ZYa4lwPBeNGf41lIxFmL0GMUWA+9ERu08F2ywWmqpD442Oclg3s2klqzDSrf/65xJlNu1z
zneAZbVrA1Zl/Db5ChLZw8Hb22AdMR4UDC/bDTj8JLuiXrOmlnKjLqxBYS+T6Lzhj/XrQ2kelwoG
fEnP58DVMmfIY3H15uqKF5s46S31wHlOzipji+oimqAK8JNCCpI2e8KxCeR9/uUgaOmfHyHpazPZ
5EY2YqBb2oIIl3ty1mCVIEC+V1vlRcGLRYgB9dISXLcyIgrrq03KmXJ4WQluDfjJJlKW/Q7oNpxt
h1Ema28Mj6t+EYjbLgpRNArYbWxXPdIA4rktgxXVt2G5fp9vflwIyTLxlbuZ9GwnE4We7zY224LH
C56FzuycYHFVwn5xmbzcot0Z4hv+CFdh7Ore6/lo2ZC4GFv+qAMAtnOH7hb4VRMCHvl0FbJA90FB
3iYNAWoMBs8XKV4ODW8h1x9pJSUG713Ph/QPHNjxH0UiC62y0dSe9rF8Z/XflU04oxnzcyMC8RHz
HebWP6//wae/XzBlOPqvuIrxIFfXyRE10jdt7PgdEUhrbrGhA3TUxJfylgFaj1Zwl/EjnENDfjG7
2aLwMAVRHzLD2aKBaj660GjZ9UvCrqmWg0gXFEGc4f+pOSUP2bdrvXkyDhYdnMuDmqx6LnnOaVFm
w6FjCy2ot1EOhOg+5TZKUmH1JUkAxgmvzhpk3cR6+h1vaY2B3CmN9gWA8qp0xd3TpsU43my4Aw5K
4jVw1JdpF0d2Mt2ZI/KGt4Bqg7ACgXeVQB5y4gDINNCqN9U+pzWiKHRDd/rFK193aBa1E3JYCnoQ
DBMCFF2q5zsouHS4wnDwle2PNIzd/5wycpISybQfyZK2e0FBrog05ocCfTUBiVdCKexu1vBnUYxS
qKnu7ZMd2rXqgt3BRmEVj5P8TvQQMfZdBZ4SUNm86pb01v82kbU6H74XR4RwzgVCP9FVEpmkE1gq
tiMbArVdpD072I/AtZoqHNqFIft41DA1aKbx6tbcanZ4cASskqQtkHJTLO2AibEMgxMx5JvdvOAn
Ns3bjPmLBGSJnrgbghkgYtRRGGov9UO3d0ssQJ94v52drx1NYuCVYesLaGKbIxgO6RPflV7aNQyZ
Q5kY0mFWCds1DmX0bjwznSNlFHTcNZ6Pq4io9PzzKQddlV+KeJg9xdgKK92TMpy//x7H6Sfd0yFr
Jfh2v8tacXdl0Sq9zB0mb6ecwyIxc3kb43frjfqfACLqplHq3Jg9tQTi8ebC/1CaMHljZDv/dA2T
2Y9GMbwBflDJN79Jt3Ma7vLTMWyAJZM9rlzGKELPUje8mlEkIMG4NlSRmQyedD6jOfwx1PrXUkup
UwNl6UYWJORSngNvJKR/OV3aLm8mAwmgsXtRF+tRups5mNE1RlfPT5wmAKo03i5EWFeiNkyMIYTu
gZKUqnriDcfPZYNmN/GdiOfayXgbtMYSw3y5hwATpf+nfiPUGNBHntRf1fa9BlLT3o9Ja/0bhACU
YDfc4CO1yYdTl0uonAQnm5JbzoxAFPO+HlSoRTXRB/SXxCNIW9UjUREZcZaskHDK57DLT4oMZ4hX
f3sU5JLGLpBuiyZTZhEiQ9ieTfANRKiUxnEIhcWTDDc7JCMWMwrKsazLG4sbP0QuHdqi9rbAVOQj
R7M8L3hdIvwBQufhACMv5bTqKKiVUEZQFtoXKirUYgcAhTPa96n4U1m6w2gO1iCOckXUwAr+YNQ1
lr43y4Qy9cYjfS3Ft3EvmKpvFJk5D3jvGSLXrLF68kApdWZ9Fn2MvQlqDLV2S0k1wmyXukXZ3QnV
thD6A935naAfPUK6nUGDF4UtiGJcOTUcYPL+cQlZK4QvqdlNUXYYBsfsg0SULTHFD9NEAVCgI0iA
zFwhCubuIPQs+nFwsR5WyzDfs1P8AJUIYatSiRY2qzQYU7z2knDbM2xPC4m1CAW7TOdxFLb8a+XA
nVZq9JfMfIiXwwoLckt5T1YeMf+P4NiMll8h/9qUbfPFVRH5JamByUJp9n0/zLhLEyovKhRfpNgb
vKT6nNsi4QmT7InwDckJsyZHhIdI1iTTcx8LD2fWAFwvySqSVV5TST3Zpw5ufQIN/rATjFCY18OC
2RVW1/FgW+vbLk3R8Sx1vhnu1hUUpl/VmCFotElNmudZnOQmZbjSHyhNUITMjkFVLiKZl4NdqInL
hiLbvsuCP17GDYBi+fyDgrh98DBdpBx9+c9GHpGmD60cNmD7kgntnRzmkMnhFLxdqTPRAYumWLI1
84gs+P5byGTHuycKJEshsVA0eLxGAvRXiQKQ7OtV3FSeqQEDpww+Yz7IKjObjxVMwZrVAp0HzniM
OPBpuID6pLxM+FK0IYbp33/FGY5kkPR+BiGepdmKrV7hnSky1OdlwXOjirc5OxNP8k6n/4DwNUOf
gC49UyBdrdAucC4spJkygx8VkMQ5dYqDqpm/N8r4/wPBraYicKT4yuB38eeIJP1Pkw34m6Vf50nS
fnHF5BY+MV0rDyy3iK9v4tY8IzqVKa/JSc+/iqO+RkpNiBsVtsNRlAMzrmoFR4cAUM/8zNR5ErhS
7bLlrgxdfqUmm+8S/psePo7SHkxMe0e9cyqQgMTheW2Zhy9fe2hEUfJv191GZ1QBri4vmqlxGsOB
Ynu7AZ/E5MYL4Q/dKKyrz/Muzf6ukkIINAmL5VC7BbPGegDpdoFnZiCakeuX/Osi5knEo3SPJP/h
GRIvnkIdxRgA0uoiT7Y6JcTCuxvifQrKleCfs9jfzaJd+rsksX3V3z2sXxSIL+hYtNxNXJid/ipF
EJpg8A/vT04RogTaeLQoKwkA+VzJJ517JxOY9I4UqT+RmTGrEKumIJ/+aoxEGAGqBcpEt2Cbn+ZS
8OqHnD9E+AgiVt4msoFuPt2DSe40DUvPhHCde74OATM/Y3OaTCQZQrsDv/A3AOoprCmQYY5p/tCC
uwn7OEuQWeRycPhtqvv5XdZrQlQqH93qmMyxIWCBbfXGzxughPcptxbYNX2NMGBImdwYsH9DiI7x
q1BXZibwwxysJh2UvemVsi18fW09J0VVUGlqquOVKyzE5LqKNYg/AayTIM8rjLkw1K7ks6FChRd+
rdVAOePsLvXVAuUINzV1Jx1MvwHEqQkxSpKrFiVjpuGNCXtJXbDFVDIf+tOJ9Iw6lzRBi155cYOE
YCmGdxwvQSUxE3F9kGafMMgmGHhjvjBkTOsdszWWsWduUv9wlGk4VU8RTsgqSthseUWxMgd5RfsX
JRoBtoB59xMiDMqBUO3RdqppRcVXJiundRa+qf5jaT6z+XvCO6S2+PwrxlFWOEu/zunt1EHnVtUk
XB0fcfpItINnhpHIO+PRw7vbzc4QiuD7G+ooQladx/lTZKqTAj9PbIPEB/LIF9CL9proU7R5+ep5
SNKxq9jOMDV4PqlMBrG/2jBGmgMjdOumvDq6BcxbIoSJGoIr7+RcGOt+XChEeWnWA8ASbhaqBQGr
y4IAwMpYSD4Lt8gk5wy5GYcsj4XL95UuAuCMVDp1IWqpSZ/1hg02lRZDU4RNzGMMwOzeYMQrlIGw
4g+cIxmSI7fjHnUoobxT1OnF3WnvvxJm3TGlYK/Ocwf2wn22s9AfPfL47W145oJQAeIfcU+eTvxp
utJ3SQ8cNh0lbRCBpvKp+GbAWuOKgRZw6Q3f3y8yF+hxH8hiLSHQDsLgS2Pr8Czlibl7P2rWPZBo
rT1uOhGugvFqqt1kxsG7X8NWc6cJ7991oBsRM0SCnsqkM/g0VTbP+fd4K0nBBi1Bamli5uC9UhTL
XgxX7sQ4Xs07osfqciZa+Ei83jcOryPIQm1XbeX9KhaZP+OlvWbOQxNkMfISIRHS1JLTmDBYPux0
OQYZy3EY4mrKrzdQtceKsWQCeFx4EJwiQItXphQqV36pPPc7eFTrpkiJyoR+Ncap++x8saOJr731
qB1akQKSD9QWTdDNGoA93CXwyU5y2EsmTQ3FD/wUjTmeZB7vcmGDGKeiRVWkOndoOqHNox4EZ1H3
gUB910ZuW9Y3NftgvJwpoQbNzwiOvVTyY53mS/b+K9n1z5FKeRwft5Zl12YBxDdbdSr1FpEfVqlM
oI3BZpr0pL2yIhvVwE/+Mw/Ki2zP8VL7LQG639k5NBH7gX+q5rWXGfr0AGav3VsQr5kWr3rEpbF0
69RSnKDqyfWoyv1Ep8yGjzaKwvKSzLQtpom7d6Kd5dGM1hYTIwfuv3PqmxAho/kDuVyO9Tqz7Bd+
pY7bAAltoiLsjif1pq3fRdXxkDxUq95L7NMsUIRH83gle928N7xboawbdH2j88MgM6dluuaipSjY
0onU91KpLjIpMlI2aCu95/Sr207MLBrszLRPKrr7puT2p/lSu+KlXainyPkgdSbriQGzNdJ+2JVL
ToNU7lS3WBIkXA7wFXDIJ5NVah3aA8Pkn9eZyyFoWfbarS/vYq8GCP+Bd3WoDxklBN/LucN29Jl4
KOi8BlxDRuGKYT0wOfgIWLdkEQv0J2turl1LT7apfReSw7UTqPJ3LCxkjJ+B/qLyEIpHSemRBEBt
eOj5RgBpTO0GuShKxkzzo8odxtWubppebqZooDaPGOA70P4kUDZYm5ZBFWf2kokIOIazFDIZeSJC
ZrY20m/uXJDR0POTv4QpeF8R5VDSJH0GPsdGFsVaL9nEp7D1Tom8l2i4mqtjFpxVDcxTxKrNc2tb
d8gLgC+N5sdHydedrbr07s5eMLimVvqso9u1PF2Ckwk0ZsklMS9N8Dr/somPi3CqPjhcSTmqNNIq
V3VythoHHUzkER6PUV9GMRsjKy2LaX6dYwwAfQavyqEaIXEyhasHNKBdWvuV4CKp2WZL0lUGI0An
qWOi6Am/ZAMnvIHsA07uOGcPVmHAQ/NMP/sjmwpCazj7x82C7catPFdk0eTRP+jNcYS88mTz9gkt
TfCivrOtZJW0snmfukMfO0xzrhy9S2mR5ao4JyL+AvyV9B7cM8kKD7V1gCpp39He3Y5Dw83SBxNf
CIwp3W1Gh5U2m0hWvFT31c0Xq9Fcjh7hWxOn55zZGQcMo+8SYsXfIVzt6nnn3IgWJE1av9P4++2j
rVo4fOVPQZpGbOC2UHKpDhKEJq8qljXlAjvouwQQJbO8i5rz42uRRQUaCoip+8OYQ1diPtNjs8A0
v3ZzP0gbU4QyrPcA6td0/p0Y5tJgQ0/LPBgu2Ktp8uNwrmRN05BfHFfYE6RbnlP3rURANqyis+4s
7l9SdL31C5z2nfvL+IG/7C4ueUWs8iUyqAPf+4wqksS12RUjN32d/OoPiR5OVG8PQVj5pjyG0vMm
xqZmeLa7OK6yahOeX5sejl7xFr8EZ6gROa9b41K3SoReSaPOUqGF7E7thIr2utQemy8e8RCcGmfj
1sajLIzoRkkNVvGSXTkajK/0EMpAadT2Y3nfEIhnfNhMnWl8izSqoJGi2aN0G7CvgsamQuKfEeCx
Nj2dMS6WVdWhpaqomgEi3rwV/L7T5PyFcuTjqgDBDX7RPb/O1ToChc8L9hQWI41YnloMEFaueRKt
9MtNjnfwwLmQJkLzi8dVDKmRFUD1WagODGkfLZvrkw/eXScwbvTuzfM2+8CheaWMAVWYTBHq3X1h
GKLLwHMhsDFCiYrgV7YOBDxdxTBzXyHA3Q/6zofw86TPv3sGOpYoCU9hDO98DvO0MGosalhUFfDQ
xWy9gz/OWvR1sx7r1x+bbndpJltc5TrcYTzY8TCOKVkDyBuXJCYQYgIsFbfp6UcT1kXogl84CMyS
FVlbJfEOIRoWF37g65Bcz3OM58aw3TfYldw0bcyXvgDLbH72AQMir/zyW2oCxCmaUMLq8ejPrtg3
r0Oi/yYS8odCIZkimTVZW9cZwr5L2D5GmrLUQjwnXq6ZQPxJpwc/Bxzxwq5Kgcvev/FPEVQcQExl
HHAcdDsw0a/sLZRNSfDk36rPzUeEJgnkg6KpxldJM21dmHS8FJv0kgNaLH6J35Zq380T5szJtv06
+zSVT8I7P/1KkAaHuIgOEEP9RwjKxRdwqYq7r7XdKMt3vvNtQgHTUKh+69/bHi1g9+I2mlSvVJLO
Xy1uSOb8HRmykkfL2L9brWJ3ll5XIjo13l32rYQXGFENZZ5m6EaC7Nhlu7eq8mVewTOXOMdeX3sC
CJs7Pl1u4RcS2OUPoXqSb7dje5BB00j02NnLgWkvWSMbWjseq5AJKQKOQGYpyKbgO6icOLy18AZk
kZzq2qo4oF1833b5+uO104zIjr7H4b+wACsj5x/lWBH7bS8rr/W9T60Koa5tFCzN4B1216wbYHgy
lzLrJxFteaePwFYxjBFcAPpcA46NgdegBJIZi4fIplNmtI5ZAVcZLIJ9vcgTyG4xZJsD0OqehMRX
nwe3pYB3HDv4PC87GHnXc4nfRCUQaWaG35CFpYHR8aq2eqrJhmHWedMPQDobe5jDbZT3b7QC0wMQ
noLeVPFwypiF0biG8MjoeQ8X6qDoLIfYmRnHnmojjXrcz69CSHd/wIeWNvFy9tYp4gu5nSp8bpEq
1aAb3EYQBH5tY8ikk/epNm/clo96tQitz+uqSD2ZKRv7UNQ7T/6EWuqFN8zctM51+JibU5Lj5U9h
r+TL0d7Pff4nJx3siG4w91eT5BkL4S37K3eYk5m1QUssRXSIUMA5eb2S/hWwSFAUiP5e6U9JgCQ9
a1wqfGDfpVZCYVLVJjGaSTiJ7qgCxnIs6u1S0IW4kKDlI5h4l3Y+lQMc0Zjouj1LN4XwgBdEOHR+
zYH5OpOlA3kCK790xcWpcMuzkoAdksT4NQwFnpLUz8MmzcF1WlfgMAKFY9szu0dAX8sLEv/5zI5l
77Vd58tBYCKXdC+T/TBBnXKkE3cZBlE0D08aTTO1UXXfjkpXqAlMikv33/ar8FUbkv9bmuaDZune
BGglRjRJ2ZzVwXCPT1Lg8GhXLRy94HPkGWmnHYWTv0kqnEQib7YGIH9u1h3OAsX9p3JebIwoHpuE
udTC4LudtVhRwuHcvVyOWvKF7j07SAAoZQO0J4Hjr2vGD1iXaijidJsDRTvnihUJQEWwXq53JfAI
GCBympg/PilTAZDjXp33dvOBsF15YqVPgFiTaGGEvuvdJFcIEQGzoHdhD2xk5wmd0z+qvlUAiLVc
5CTPNpQetZRvph1WB0JiGIx86y6VuLfjS2C13QO2g3pJT0F8F/zxdXwCG8S2OBQmEvei7CUlDqmw
llJOJM+71vyDW+Ncf4rZWmV/fUalA3rA0Z+9ceqXggrG5QpxJ0qjORzv9MTyYvKMhrR5haIskTnx
O24/SPbt7JQRYKz9X6wxB+PNvjyu4V5oetZMrvwxrQXeZjFubNrmpi66jPORi42hrxDyMYHfyseV
2+ts7gf/uSNW/Lgq9HXHSn22APkZEymF4cHH+ENKDZ+mjzpQ7Q2eX4VF0OWVGRf92iQkjndOWV1F
cSS0VqtLS+/z+HCKqtn4O9GskHgLeuYHYmNCeG45q/vlCM/eschE/87jOdGMmlbPVZBvSuvTD/3t
/n4gUl5AyAweDno9xGmnhkYNHNI7WPt7Wf7CfbWzqCT8MgQHzC/YwtMTe6Szap/aKX6a/0lkFYNl
ToWPjqJZ82W4pHcbyEEhIBr5pg0pBPOWbZNYjF6q3nIUGzFr68D0P7bjlFc0ahcbhDAukCu3+nlS
yqaH8pyEKkDdlKX908FbwYXZnQwSTEtcopi5sxr5432nMY7RbeuG9DtI7fuK+osk1FUJl8+3w1AV
hYU9B1zZEIw/LWfh0ZXE8MWbafkKNO5zFoH10m2q/yU7CyHZIX1G9YJ5CFCEJumlf67/34v1fdNt
2/NDDQCCWpQYRSLs3dU+khVPq9ZgvDFNok5dLotTrm3I5N5n3vKOqk7GYSgQyeSP/s6iOnjk2vk6
OSqcploYzkJ8uYt+H2V1L0H499KpUz3PmwMpnUvo8ErSN0GdXWYlSNYY1In3teeVQsXxgabzSIIM
9jRvo10wm4yTORihTX3qBESe1P7g490g0RcOeMJjhTQFV7m6VxwnYQwrGJDYxTFNnRlSbVTJIF6N
/WxwYe80oevmLCL5LbLgRPhuZe2ddxOWajsl+0hmXraasH4RMoJ9iY6s0VPwIlXIWAr2fwVPnlzj
UMQHbk/2iLjNxxBrIwALfWzaJ60hxmBovo2g1djjm4rkYl2W0BHAjxdXebIOHN3/v3GKYEc46eZF
pMRLdQqUlx5XFbHtTQoh4WMizWr5FIL+A0fEnHHbrlVIOK9M1kqnHkJ0DGjVvawYKS1eL56wtclv
7r/2998hc7d+U8RrErPqKX7jmh/ABq8TpoK8PnFpEV2CZoUkF/x14i/5fKgC9ejICGwB79RT/R77
dZeOqjbyLv6MgWu3JTeRYfXIJkzNl5SUgR2lIBfGEUI52F23ndr30eVqp0MjdJFVX1ROXIsqK6je
RqpFIaYid+qOMDGmkR5Cc3VeLjRSWBBj1P5X23KvB6shTBLuii4oqFvLnu/rm6NS0rzF67B0B6uP
DOuP3Fd5MPGZJlmSn6FeCqK+qqTuoEvsv9gaoXUWJM+8EodY/QcLJfoJRTaXP8jYDU7DVKcSiJ30
s1SwDZPUNInMenmPnQefjTID5KvTsqHJfIMYEle2N3jGoRAsr8QJcg+ZcrnCt0f6hTOPmG85lJCl
evitmXJ05OtlnY5MLuer+Xs7hSlxD+7o6N+qDvpG5+C9Kj7+CNAc9A9HIhTsWnXDRIV8nRL+sRA2
JKituPSRUtymHpjPHkZkTkB7YDgU7cyUYMLuvgTyFWPftOB3lWPAXFuglSq4qeN5yIZHIVgrTdsR
bp8J++UirRFxmubLkH/91jGd/x9Lfvp6QaGCPlzoO/rTjYtcdGQFYn+oowW7Yr96goU+G7ceRuQE
Z6hOEL3eJ8OGxg8ESLdvtqlN1yit2vjL2yzO+fi6KsWwpRZA5XoTXFLMG+4ia+R1V1jxJtwIYjL/
/PyLaycjkxl1TKZUMa/OZdsyjD5bBWrViY2LaBh3nKP65cTzKwpKhzCGdSvV7FbF2+wwaup0prkZ
HoOGvhSb9GgEGakMY8RKuRg8f1+HkaTYsKPjjyr9WqXrcDIdb6hysb7Eu9i0dYTlqAB7rFpjiZ/I
3gNSOfWeiE5jMqDFKpeXRwd98UP+6fYej9TRdCDYjKWvZz4LsXURs7kWPuZiA/T4QlU71rWzyjcq
23+JB6AAeKQhrIykP61AT3VYH/hNqDmidpXZdomH7VRRoFSs43Ma8vLDHHRHiCZ5YrGwDeY9qxf9
bcOmUm58MkJB0V+uvwT/OOvtyHYqXl4ztDnFdlbWIYLzmK2UpWnDOxX0GkGCHSDhT0yQIFdiDMDg
t7vFJ+3HIFB8U16bPvgTj8v60l1RG31wQzNoqRtPh6PFZlNyTAtpWEQOusSQjCDtvJJIjuzIHZTV
OhbLbdKn6j/M+ZDAl4Gm5BiHElr+j6pdk8yyRblmtQtA93SiGKtY44v1JQTtnvu1L3BVc7yN3j6J
IwXDKG2h9FChwG1rHtsqzGgZot4EtdT6zYnLH5Wh5tRN0icEn1zG5a2e9UxBt5h08hWYNPFczC/3
Y7YKh00wDd7Bmpao+0dZ4lAsCbWaoN7i3SUNQbA4a1eVlJaScR9Au2ClCLI9h3EdGWBIfnj2im8f
AuVrYY4Dnbl0T62Q49C/0ZcDxQM6JzIJoVaf2VPMIV7d9jCOEwjaliqLNVafNczR8IfpPakfbAx/
bxxY2S+8tq+xyPrQL3jt+L2sJAZrRkCwqveYxDzCZcxCJIKhQ9fyLjS5650QaCJHGrnx5rFVWrOd
APzOuqEhTJNMAdPlkbzinSISLTA0zjVrMV9FVKdz6xQ0PnP0WTEA+PWQnmNcSf18AmGkRpEjgVXB
ISqRYWw/j0O4NbRUK2PRyyWUvzfEV+RGXldYCjGuFETzxbTktEyqQ909hozCD1yze0GHb6KhUII8
hGs4Wz6UT4YKfKU7Sqsl6xYwoq3tXr92a/Zq6BpqHt+3k84VcWyGvY44qEPmioICby7SbpDJuZUS
wsPKMCT8CHI8wwtoTut+t4G1BTDzCCJ7RvDgxqjiqe/AgYOTTMIq8iyzWskkPlorx3HvH9qcJL+8
+7CR//TZoMsa+H8m0nSqmGdSrzp6sUAjEkmm8lvzcKVI9QqCaqE0BD8m7/1Gk7wmB18WlJ9R6wt3
YtFoSz7qHdC0ga3s6vTI1qKoZ8IEv6xFa3DWCQdAXhBMG1tQKYQSB75QOnpbTwXh4mhUSfPUW0R3
yaKxlMwd6ZjVHz798u8mjOoePRfjgRlNvE5L4GODG5+CZLR7LFYmInQBVRZlGajpe1YJV9qfGAb6
mYahn63FPJVdguhFILevJRBOWR6Y24OvjNvU9+brs9QbUfMJV/dZJfpWYIh3uiYLCSbp2vzLrSu1
lH6UvaQFKhgyV4LHA8bD3c2RpliXC50B+Krh+37wZteEFXsmzFe3l/p4Gr9Z2cBRDtsYBRrURzuE
pbjA6PZLWNmKBf1bLlvy4fv8iQiUeOXmkdirHHCNxHdR2jz/LRpkKCS89+ay3QoNouor5JWce1At
q/Vw3ySchzpNNQ5OBeu3abTkxs9rYkWJs0xVMNXcP2xW12HBBhDdLlv85wzq+j9PjEd51M6NxQo7
hNfqj2ghsxRskK5GbHJZesOxc8WhEPmYgxReo2ubMdpM2dF5rVEdlzgngHQWCImwsR1ran1wO7MA
OsbJMwGSj6U/DBFlw8XDxMreRxeA8iuUNw675p8kc/voDlh0IlvukmVZryTUO5MqQs8cuPUb1pKV
Vroebb4lbYchtPNK6/Gyq7aI3NKNs3umPZTz6UahXebBiB476h7AxHYoqdG1fEd9/xvPfB9/TBHK
gtENXVkESy9RBZqAFu24ZEZ9qaCSdnbwMafHBRdoim9crJkHjE4bAfS1tg2vAJ+W8asTtMlsy39B
GgfK/e6Mx/xZ0FL2y0yeKy380tsyX2vJaZ/cFXxxcktMV8i6/GxZCJXdcQgv2U4xGoZhzRbdKiiY
9e6O6PLXSuYz0WoCvx1EhTeFev1pkTcc8XVSis4jixhfv8JytVfec7cSDEO7HTgLnztmVouOx9EY
EcMhkzu+4P/iGoze8Ugr3eefofcXYJrEkONeK7zvc34aioCUSh4hdAKmZTzjn0iRlrLu58bBLR0A
F4NvQZcfGfpELZSSl7AmcSAvlLKOzcO5r15NvsRINUB3/EYrTNGNdBSfs6PDrgl7bNWYQulSM2bk
LM5rAPJA7TLNyR6GBdprf63a+6U308xHyaSUhMbg17EJ3Oi8bLdgM2nAv4ZZRMpIbvdbA+Ere0vK
JvSZi92JZARrJgwKll2oZQfdQTINQDLRyvcMl2kAD01F9DKMGhVKS4BZZY2/Hgv8f2MJrzfUMlzb
kjVFS/WctGwZ8OwJBhzXyzuJjLqDFv8SrOMFxPVmv/rUdOTkO7/KCjCDjcgEsgMl5EB1Ul6Ns7vG
h+QMqRhiYqYc78AhUf+K7IRkZUyzfQYQ27Ck0Whcpq5JVjVvbDm5hx7P9DSP7osQqEwNjuQPxaI8
w5kcUWNHREzqCrV+zVIhIxVPMP2uVBeR7XAaZhX5mIn2y8c6pc+vMV3vjbY0uQ2MoYAQZZehFdw9
VQWXof3r2TOdzynpQlUwbb2I2vDiJCOU3BaNryWevsJ0wyvQMM8FHysC0buU+MJ0fivXtccRid4V
XWXiWMu6txiq0qttcvRzSbt7118flBYtD4s7A+bzS/cj/2Vh+zMqn/gFVmaNeI4iy/XHMaHiiFr7
zTAR/A+C/J+nLWz9z+NlbUgkk8BugcdoNQOyhIYxyM5l1neyyu8pQIEkkqATkVrGbsDnWsJweBQ8
PjmHump+qesdG5ldWTD9pI7jmuxJJTZUGx7+N8AMRGMDbvovKU1rxpPFcqhAs9G4wmcBK1oCkIPg
IxQ1DRo0x6Ooov+g3M5o1MTPKDqJU36EwIMEcHa/8A3pOReo17ZYd5nfk+eqAUf+m+KSBy07KKW+
Zsh6FVtCUqkHkceXiT5Oquf0A4p3ccUb577SMDzL/OzkeUPxl+PDf821GsHKs0Dz33mALMCWsQi8
S2rFTosq6d05SyvUxVRaqoTKWwJDjA/R+hTgcxxcN+IxJbafqAd0yochB4uBp1MoN02+BHdwnAcX
+5lQJLLAxjFTrytB+FCf4tv5+GQMjHPfYwfygA1ujrfuLitqtUwyhjpZlhH6UJMpexpYebWsC4tM
GePN60vWdVgxwkGwTbmw+Mbz9DKkLmC+cYHJDQLz+LD6/uzpAuIvseqoAz6NJPJJgBmupqmTJzdm
9n4t/ZA370653BfnVxtNYOuCTKCbLeqsojhERQ63ayw45bJjE3L3f2eXlM542HAk3PU64Nmwv8VX
1HZ8gVKdCym++YdAgwOU635n3qRJlTUB8DAMaeyfU89tEObVT+uSCD/DcAn/B+82VTnOcRy32WDl
oJe8RnB+H9L8H1pnVHC0r8SSY68O49F1nngEU4MzbepYdRr6QUL3hdDDUdrEhpuXYnJZEKuMk0FP
8MRiIlnoEsO2SfcEmzv9zTNSsiWHOBcUpqUenMqUhG4hR7Yxtm8H0kGDC7u54C0ZJHgbQQapa3Rq
APC+oe3gZzP4XQzizvAockvHSGlMUJfGM4jaFwFr4VUnEZB6NWQZNgd69pV6/mwnTAUKHGx+y92J
cnZXva1aEXNKNHhXlhQPEFlnsFzL3iDzre2EaZxkZxxfASZDfvdF72fdua2Rf9Y52007xl4Ox0D4
5SBNnwIAasJiKcNyiC8H0/bhM+byP1oJFhHEAft6l0Yzz19Tf9BjFKhf0dGac1hLnLe2qtvDvJXU
WdgPjk1KX5DagNr8uylrYntGyRyWUhJu6GX21DAGFOkB6hQE/XRzD4gy44rpbhOHRb4ZDk37xAM/
l4xntxZsAJGj5cuXwtjzrayGP2jTXjrjk19llkRLx8v8jIfZfNNPHRx5Pm/H966oo5WfZW7Wa9FS
7uIZQ6I3jTXiB45d7PMZsFlBPZTk7kITO3nx4v41jU9HWnRTMqNtfWiFE1eQBIoxBxPVWehOtydK
pUNepz3zV3jQ3DCqTFzjB+e58Kp+zNY8FJrfrc6nVFOYWg0acWwp99uJxZ1ae7oNMl+a+eWVDnUJ
LL4uTAsd6Pu7W0H5rTTeI4yd8rUsBvv6z3XsFuokKzGqIRBs+oYOZrSG/2R6kPfKa683JJCGmcHc
hb5a1zT4yzV52MRkZDppnVtfrKWuYa6EHdFxUKLEapoL4AAjtTrDewnOLkYyCrOm35oOVfAYmhdS
UIOh30FnyNPXmxjlxdnTI1OegzRlV/V7FANRe89r6dn0Xrc7TiV9puy33WqMY8Z40oYovjZhI78A
RoOrao/hi2BH++GmNPst0/Gg5wk4oARmjccs1APcwh0yrD7r8cTxorV44w8EuZkT+WPs9eSZISWX
zVvAvgDxZ1ng9NFGjNK8eStyQUDFfVuOt0XAjDk9Dl5A73WJrq8C8SG/WFjR2py6nl9h3luo6Mwj
ovBcY461iD+fWR01SZA8VjKILCrGXfdR3PhPTq3ijbTAbFrGS4kMJUdhDsp/S5HS24aRReGSxxdS
NIKHQ1xclLtR5tjrCEG/OenxVa15/frfiibNY2q24ByzGs8RgcebmbPsiSjIoxO0/mc2wMC1Mcg3
XByxYVfWehO1GVn6ndLbJQJusycLfzSpdQBJoLjv8NPoKdf/IBF2S6Z3c2IBtbDROjFpu98qs8WD
sJRdq5X51fqYudCldc8LzrumTrqoLK3DEcvRBHNaWkPnMag7sLYs133vo5ygCEOLB18kxYn07zwe
rc9TEqs+E0ZvwSLp4pY2fSq3bCPdGLBIFvRfhZp96c33Kp976mh4Y8IBBYjOIJryn05O6w0s0qwu
G3Pou/Y/0fcw54LLbfldp4mtnT+PCYI25h9MYWiu5h8wo570QWDeFswMgHuASQq3dE8lrnQUjNkA
ZYbOqzI0EQmjZjGe0E55jRXeYnIy+2OIfQRgdJAbb8Huqa5uW/1j54kqDv4jyO4F21B4BG2EYd+Z
LOUpxDg5DKrbtb7Nzw4r5Zr8xY+vXbvFww8qRlbrwNDR5gHOpTxIaOUg9eoeRi/SE1QoCsi46Mkf
WFh+me+K/3mHNZ5rXC7moj8BDWYJBCO1xGfNpkcC0EXsjo13jqhAOerP3kl2vuAHBaIg+pK7sSpQ
MjbDjcDTSc0f7JQZ2qBeDsbOQgr/t0O9q35JaJI2N4XQBhrOnSgl7uYSbg01i4kSByPKFNItJENw
Ora5eLhXisJhfGaHh5l+qUoJ8Lz5WY/FbLtUkKknK5l2WG85AGG+jxfKGzJTE/ZIiSdJPsZu8L9/
sfr186Fd20ly61IU1n88TeK+YODa23zt/Y6xGWPWNuIbSI/Z0i5DakKSBbXAnU7KXPYXhF4tAHPQ
27gZtu2cM3XouVWhE+bd43lzB1kkmfcuEp3kYB/mfrGvo/PPikreXujPZlEO3yEixXZRgqwwKtgA
RSOtamM8+oVUjeRfcAOl2HUEhztVHNQBxK2O3fj5Wd9hIR2rZ9k1O2vEyvAu9jZkdqdkAQGb9Nbd
Qa68PI142jI1HRLkhmLOph0FuMjvIuftvXGkstj6CJWJwhq4FE6EYRqRwn+938/MMhr1if6Ug+n5
dWRVrEKBCBtomwsa1qHKnTmCeWJEJZHb5/rIuz2JE6QoTx5T8PbPjtPBlLmAOqLEuZpmn3LRe0zB
BFEFSS/KRb1ZimHOVROorJkSG/PG6kxk32CDPeKoOJVpezDUrK5r3RMOX0w0wkSx5+x0UrrPzxvR
nsWPEE1W+U782A4echS+s8/KiTh4QogNyVmsIzkLK24F5D97GIeo1ZggHW4abbOGu5dXJtbLitSU
DHSBsPjD6Ey/5u/sSFPBozFmnH8OC3jZkD2ulLws3MPdajKRxwnnRDSlhzwareRKLhbKN/r5hSY6
WBPfe0+5zCIKJmsMQ9WJeZ0MfhvzThzGaAaS5S2b5aKR56ynqC0quIqPMhDCSgL1Sppmu2KO6rMM
wMT6BfqV45c1ZUje67HayNvJwmVfD+gS0VrpZIlq+BvUQwPxvjc4EKEGuVvAbja1T/D9pCM0kr+m
64NEldKwYzn6u+lDOtl1N3aYEfikicyUfEZAvqQ5bcDSwPWO3r05qc5IByzNQNzLKSAZm+q0QKld
3aiURoWQCihFv/ZdWofvbqK/4PdqoVRz3jrliBjIGcAgseczM5NosUmDkyVWYnzIJs2WGeiCE92u
cX4k4ZPKajbs7kwn/AVkHWMZJM1+vRUQ7T79nxpmdvL6KIxwCno+gn6Js2Hk/1S99PIR/WCNMQks
bBhPuE38H7WQPeiFFTVz3AjusOW1HAoFVQOarUVa1AwxBnPRwz73kRKXkyeIYSuhBH7Z3uSDgGll
rEbC1oaScP+8pOkqIs085YuOTWsKdRde2yrzkH9J9dBBiNs+6RdcCpQxCqbCWp5a43cbH7tGGLhe
0UqE/l1jmrUmKj6uz7LMdj9ONZe29ukEk1WGZ7Hor8i1/TNo57cAaahGChWF2kXSRkDI5FUkhlMR
K31px1Us/D6mo1xRjTQLUIKI5IXUSh0rHH8HHjnB0PllLwerCK5Up34Zih8MMSDeC9gWzfbz9RBs
b0BAC407vKDRZizhKyjN4aW0FaCmkdmjKc0SF8oY8boiS802Mj26RODe6Z3oH7vAnldRzu6w8sc2
NakSC4RRYhEcEQWAO41ke90kKz7Rj3XXJiXq9hDw2R8lD7BkIZRl+LuIXagqIext837jcwfwDIAf
EmeKQxmrszRU16gGVajFLNzvV2Fft1WkMeXeexVc8jsvTPDlZnZGs6NOEWczPtkZ3muN+SRuEo+4
GTidmKW5Qph4jD2u9dbexh1X7qx6iGo9PPv8NGtfhfYK9l17nneqopLtZZjsxDI9Jw4OnTS41o6P
jirSPiUEvDF79abMU8axmq2FaPTec2oWJon0sL9UoI8Bcji7f6uzrI2H0LYOkDkn9BYC0wLNCmbG
XSXU2UTdeY225HPKbwkS7luK/dkHNJeAEEBXknz6ciMvCo40SRNVkGpotlRRn3Ba2r7rl35QKLRK
wAr3xSPSLB9F+Qx7NMwudouPZr3EROaurTtY5XOJfphm3VCj6jziZkYwjrXCjBxUSb/2jDAUD+3O
drCzTbjp9a6CE0oTwl20LDk8Een1iqUJP+pXIr5cjo6qWts66d3LpSj8oR14OpywZCmDFiwoWv2Q
/UNbA5JOxnyawQl4HRMQvVzbMB6YMKxCwx7ZWhSW8eaDtfn47OKhTh1uv44eWvXRVVjw/ETy+YSa
aOd0rpIxMUyN1GjXZnkK5L5ApGX4IR22Kls1FthsmaKTHxPb32KN3q+kZuJ73F7dv6xWjlX6mgjJ
BVyYDqo76Lgf8X0VwPPezIKmgwUJE1NvFPhZhOZQVN/0GHX/uLRDJXts1yyTe3EhbiHX6y4hxVG+
sCey6ZtX6a+2CA69Ux1OzHnlVz+Ur3SdMmiGs1kGywUgQaxwzFLb50hViJDXLGYETyQ5XmPsg6xW
PlgVI1GAgdOWWgFKOtCxfmSpgD4leIWEpelwD0PN7LkdZyt6ZfwhL3b5Yjfx8rM3S1+QGLC25zE8
d9wNnS4BRFlX2MsaRNBh6qX/+KzCWMYa9NbuCuihVwM9A/axeGpybaETuLM4JnVomPpUype7Wf7K
9NHZK4PlVW4fOd+LzoJ19ss/trIfzeZTBoVx5N1XejgrzXs8ub34EwKWNA1PsDcekEgXcStf/cgK
/w3zLGwMJ/ogfkk2KlStRffHCjyTrFrZyTjr5rjhVO1PcoG6zuG+TG2b0uSWZ6n9O56vgCeBW3Pe
UgZvUXQYXzexTKJ3zVRBf1kIu9BIQ1vsMDb5IntWFzfdnaPVagahQUTjkQxcqDAtkl9kST/mfSn8
61vEEwKLind9WTgQVrm6HTberoLtFa3vXBrR0dOs1yBRrkagK7IkxRbZlUGKUOJjVpRtJ3jQpTOg
VGTCSC+mGzS1rOdAQQxotxXi3QKiNiM9y/yvvj8J5DbuefdbrTB3mUZpIxpvT/NgfczgLhEvavA1
x1HC7hi+ChnF4BLSxQnNI0sd4789HFFxKz26AKBsMKtwAOqRN77G2f6HWcDF3Fm/hMuL/6rtg05J
hsZDUBkkwD6mhGkteYlYV4AU3eQugIYXcZGoUBXGDw94kI3ARcXjOZcC+nzluoU0Q91rrf0ArfOy
P1Km9JoFwjo5n4VDmFIjOyilkNXrbH9QG0da40ciURIpOfs565u460ZJJDFK9GBUk2lq1x16k89H
QLh9BJkPnrCC0k8dLh8ANnnzi9ozkKB8LzLxOeTHnaFUd5qwbuEiBFa10rSFcPg7O291g9graNd3
U9Xbls6hJTbhv1VwoQe0NFjZNTdu95CMgDqVIEuLePUcSx5RsDPE4FT6yj2xoGRgkBR8G1SVGBiK
u0pD4UDs3glGFqishChxdWjIvDScdniWBSIzyY9zkWO0X+lrkJVmBTUbdd/xGcI7vzFYPlVGHME3
2okKxC/LQiULm/bLp8a5oWDfQYK2sGQj5gGPWlSkIMd/0McgExejye56dI9Sr2dy5QTIpaOkPavV
Y//4ZF7ulafRMzc8xX90CmVoLmWVNLlMMw2CC3rpsPRZRjrA/lslNMBTb4xFbn178Q4AFW9Xsy8x
Qg/eiP3itiGXCqaUtdi1uU0E8Y+xFTznRchiFSrC8v9TGLINHigTxsQkrDmlmzVCujVP94ZDVHjw
72p6BGhl/6EN0sG4aKJAwvcBP8Q4xxqzTv2ZFZwb3BJuQ2pJwdAVdyPYeQ1tRReh80vc9P+AYfpO
HP5HQYInlBUSnp39PnYutLb/nLeUz/3d4cjlS7Kx3RM4qA4Xm3y0j9zcv2IS84HbvrXEfbjmAyE7
hzkkMoAyKi4d9j4Vj0eE1n2+W1xnSSGnAurH3k8mPSxlcnFEXfPglowvIJpknsBOurQKWDku6PcQ
ssjc39PmT/U1mwufFVLNtwCZrRaVmkFhF8kQvuJ6WgEO5uRLVr+L2W8hCAnZOws3cd8a1pR/5kDI
mB9iiAWLN9edh3X9tDPWzZ+w12FRpOjPEKg59n213Bn0j7JLXso3WOjwqnQJftJVKsbZdGukAT1R
kNJ6NG+GD1nGxBn+Ph3nrbIL6dr6ffFzHgdLt8KtaD/NBG+Ri/xq77v5OX4u1fdZqNXHxOCokSjt
uOHi45lhdn7ge0iEsaqhdimCj3LxYtZB2SR+90oxLuJVIpqxAwUTQZnuK70FWn2136g6bDuGxoAk
BglHheuWYsNm+STutbVjA6aq2YNx6G+RNnhYRqAfNZnqVrO28366nWT+HIgUveQZGvBs7Sg9zqpw
YHgIzH/06LdUuc/GMS/AYJkcW/fcP6rw/ZNaFxQVRQV6jTDgkkzknTY0Ny7JZTLr+kCi93o2cUwh
9pywFo9yxmG1iPB/tRKT5DtudMV4UykfzR90aodtTuFimmbDNnQyHEF0C2m8r3P0FrrQf8J7H0la
Pas326cKjORH+kBKSY9GI/jw5rkTBrmWZ/tBGIjgRhY1KWd0JJaD1oXP2JBcKpcqtSWvxKfmjYoh
xw+xuHrIXF64wc+bpFhy5Q4SaBfACoJRjGpIKKdrT4zYIc3PCl1L2HIdLx2G3Q9WOtgIV5K7ebh3
g4ki8rSQkCouOvffHo4/R3M294qSe++K1/2z7V0mm/8rYTHEqYDA3rhtgLDIhKh4LDgYjXTk09Bt
PXRofS0HtV4dts/hKotWO0QGebdYSBremQKJ1BueBTm7iyWjCHuEfe88RrNE9jXf58/2FdxFnIX3
h9gOvL965Pv+wa3rJpsrrcybmCglIpTFi+EKNSBVgEApam7l9NKr/EmlqLsocKALfct8MYQNw6Z5
P68IPdFiF1oCYIkr1GMrqRKYcHSEASofqn8SQXET0RKG+YwBPLY0fmHOGd69GY5eHJJ1EpVwwBjZ
WKb2bEd9M48fae76hbAo2SBInbMvIwPltDb9a2SSAxnwKD4fJYpSX/W7jTcqPs59z4YL770X5dy6
I2wpbYyZXB7IBiJNIVuz7zZNpGAEE/Rr54MVB50cz4gLlpiAuUrlGdcxb3ReoHEOHV5Y1XbeNqzf
3Vi0v6khvQzuKHOfEhZuRdMveqsdrJ+m9hjISAk2DurEdZy4mHOCNi8mCx3c4yI/uq8FpP0ZfKe2
3pKx8aKd4R3cODMfeNH25R5MFVgMQPI0jMWlR4pQR5rNNZrJzzPFB/dzoabc5xJFTwzyEVgzpRU1
uEcj81t/vjrBu0eseSsCDuAs+AGLAgYQbGZn6d6aFX8VfJMmvylvG3pGRKsRvzwmpm9UIXw/rGy+
FCFknHIuCXIon5KW95P89GimL/GQacaYIDmeLFVSdWLIPnLZ0aggebBIGilG/R8ScIi7hRAx4tZ9
jtgLj9bCAVlz0ccoS68X9moghzhKSqAY7UYcz3heca8N+Y/3nlnZNtfHHo8sYWYHiIi0sx6wZf3y
XjcJJAVJdT+LKZND4vD0zwUzVTlynBJxUxqLdwY1Ou8nSkSKjoh+HT05WTti2vGJx4Z/lXEyKdvB
fSu9mltrdT8icQUOsK8HVsRNSov5rMN8BzaQ6hYatAGrkwlA2aU0SZUdxiqHlRkfIzoXYDUEBnT0
zWvIQ3ZtaLh4TQm5kAfLEgeUdL87kVzx9NTqpqdINMRI4hf1cEhZsk/zWq/YDqRb59WOyHTypMi2
kL/xgwk1X0E8f7M5SkJz16e9S+lka68W21Anm8xuJA1Asr0zvX9iD3UwCQQLleea9haCcsF4QoKF
PKNvXu8qeL7sVnugVXYnTegDe3FxYbxhVunNuuiJmUmQN5f2qz+PWAShl6eWlsDtQMdFt9FVaDZU
oP8VFPvoVFO/MEfaXPyMJE3A6JsFCrQ47TDM+TE1++3AZP8cN93lV2NIh6QQB1upamprCGbTwC3o
RhJJEkEAqOEXK7XXUVY6XrRN5zRZP4h8mQoR80Cq7J8Ap81D92kIYNpuFTcyyLH//Ta2KxR1wAjU
CUmHx8znsW6d4vAiBMvCrvusDAPr4JLMLEUvPdlok/ikGGyPnCWGGy7mxbpDxbMtVje/ueZXIjog
4xXaC4mXhOQjk55FYLuc3wv3ZOIoCCnfTl1knNp6KcZwIEx1bUPF57H4eK+FrvDK1lOe558gxMfp
IOi/dTPbhjU0ZXExk+SpJ/X/LVIxqDRfnN3+gVgJbl89aT1bxu3V871scIWx56bFha+J8UV1W5vL
vTjTDA5BRd9EAmmgV2vH1JSMBCAf9oZUNK32e5VvYZzM/2SbHFhStD6fMWVzOM/OitIc/NnOd2jC
RoNtS5JEFCAT+0AN+PuNFUzurQtS03YJAAi2i4MNekijYhv6c7cRSwmTlE9AUh2vDOYlcyIGhgR2
6oK9WXf5hGTOGyN46OMnQ/f/2cFxunXrLqEUJDRILXZ7OgPW2szkummbSEa856zcI0k51dFfvSw+
yCKVIlBPZcYwLFC70I4ysSjfyj+Cl9bxEISsQGB69svtLPTihnIVv3d+RRNvtBxsTmKhQfMvC/KT
MZB89raYW1dNwyaRmrJpoMoZjZgrDhsabPPEJcSxckAKmZ82xPBTNVvaqEazPomWRtRWxUQr9gmq
owBRby86xr515R/+wPCcb/joNTDD3rJuASzG8oFfi8Rc022jZgnTbpqZI/UWvyjtJyDf+CSoqyPk
NcqtDL8AvH+6eOutVfcp1dGgzs06uPCT7iMSZB3m2csXveJu7n6nFaSS9Q7zag5t3anYUOpBvCz/
yLyruLnLjy9RZxn+xBbOiwJL+wiYB8i77XYwofdQuUEOTpXT873DAAQIBdIqElCp6txOUtEz5bdB
kHJQdOgrFt/Rj2svpkpqB7CgI/Xuecy8MWNN+aiiwl/EDiSo+aEi/QhGTSNJY1QxoN/32u8pP2XW
JyJnoHLLvjiXz1JektlnRwaHr9Ek/8tdwF8BPVM0uteSJO493ba6FKDEYjRQ9C0Mt40IZ/+TQNui
i0jbETy4OiHPuCU7wn5EgWFhyQVAaWROMX+Gz2qLh/x38h3kFqja/YHqaJNWhTjgcswzpVYkFGI9
QVWMEN/o+F+8jSZg2jXrTzNm7v/qoIjzJzUPn2tqXAYXqWylKRDumggwgPx3ltR9N1+ojSUl0ysP
hwHrIR5ObmTFd0ftqmwSlb6cVVzowKBkapPfSlz9b5W1jSLzaIX6DzUrIaSYTCtvOQVdVgVbdh5u
N5XJzGlY6ognyOg2h1bzMO3q+MPfiGBKP4ieZnB5L9Vs8K9SRU85M2t7omof6SsLjSLFjXDDaS2O
ILwJhLhJkYUodnBPqGx71C7TKhTPrWvfXkhu1vFS11V9rPNBaat7lHfLdGiIV8zMxNhLv+aMVRJF
ZgASrNqtWTOblmm6YblZBGDhYK2Y+d92tkLwQJ7DeCxpLp8bz0LsFg9TFarSzW7gz0C+DfR3NR4P
YaeZffAhxXkbbZIa9KsQ87LeS6OUuB83sjmhkeP7z3LIcb9j3UINbKA6I3yJyxNQmuWMbs9VJ8iZ
cwiRCBYPZVy1IBOz72sIRSUNwkk9aYwwLpNU0vgeFJn+GxJXrr2KddZ9Gwxevi3REdEEfLQHSfSe
95BcqCECqTrB11/xV8QmV4z/4ftm26zuPCRE0wU2devUt6gwHjteAmJ34ONVvXvcv5lNKrNVVZMP
R6ISHo0hAtn2ey9YKLaN2NwdlU4HgRoSnBDLEeVhujCgrln7VI/CeJG475MrpZsh8COZLhpWL61F
X5n71GN8MAzF+wvSQdSThFGmIc6OV/W9HKxPOsBBTdDHzJ2uFwMx5T/YxEaABEaHsUQ0CNRZft2X
qu+aaWW5LKLBjLtyYxoKlvZWau5tDobS3ntifu4socp1R/m5umz1g9OD0xya2zaXSzdekEPO08G1
rPwuyHuTHGInEKXHDZ3jSF2K8Xcr6UmbGw9dUemtCh1Ln2POrbKkXXHicJEyu5kkjVlejcV2Wmq6
eQH/Fd2FaMZTEsf1NnbikgP8F/mvBD0m/KwUBlEpJnK4CdE01R5b3FNfW1BML2+cdRsajr6FH4q3
mn7Wdq2LS9GWj8umShH6zKINUJLp47rxB8/pgKtjOG8UwERUF5Ux6IRsYBW4bg0YvHb23lgIpRtO
0iZndW2HDlOY2lLb+K2uF4QABkW8NfefdhhL3tizNSigDBbuYefNTXnZyRY0ouWY+qhNi82DER5N
HxF7FYu1nSvdTDlXMh630nofGHm5Q35wTqVlU9c5NEYLgc4gQHIxJPbuZ2DzyzicMAWu/y79a9rt
KhQXPOFGUjCOrt1zHZU2QgQWBPz1JkYpHELKtog+13UWRZd4B0Tma79GaKHx7XEdMKrQ7Frb6dhK
LvCOZil6nbTuAplK+hefgJgTWD79vEru8uExm+eom0mQbFH9QvCOBTiB6oZZ3UqqpH6/P1fbsl/J
QuO+aYqocSFUeasm+jBqs3hsHkwcd2vBoQKd+o4Z7kYLei6ApQjJ53+WHc7LDlMroe8nb5tl5bWe
W7gNFz7Ji+4tLWNTx3JxI7igRvKNihlZTAlD5Xj92R7NzTP8N41VOhNUZhQ4XbBiCXFvtCeztrO2
cwgFZapZJDOYwpjvq7ILwOEvVNlnYhgf2C5LmE+pvcZ+ayJUM28LQBzdz0oLO9HDAqQbZ0wcL6CM
S5/XTLwn+2lYjyhfpM9Csc3CfxUstK6dube25503pSdPVGW80NK8JGv1l553MebKx2YHN1GSjgdp
O4kTExZym1GWuz5CVI4F+0eNithdkBSaDkXDZW5U4bbLTFqmuR518a/wlDz2yLe1+VP5MvquDRIm
CwTLqZ4MURoubJqKR/8qQl9LDB6FQuDZV/BrX/dQPiOm16w9sIYLojxBtKe7+S/9TiJS+VhhF5T4
lktnylp5S2m5qPgI6/Jgv+4JuSSeeAI9a0+NAORK37vrqqmWo8Wd5iaTx5AsBYd6xEC455lVHwcs
FHak9qbadsxCG7mG5DxvoK4jOB9hDwvvSJhF2+FgPtq3QxVcgykvFpYuO1GlB0d0v6qBh51K1kqr
gc9ANxM2BB4b4jrsLtB35/fa0GLV4u103g3LN12zHSPbMAE5phaghTjMvuJ5u0bN/VJemGp97FfK
LxAL7YGrNmG4mhFb5OAVkCN8W8I+P0f/UDlMGUqx8z/AMIYehGWfqL1NlIVM+s9aCaGRfM9tY8Ws
bMRlGRcw18zWFv5Z/ViqKD2JKQ1rA3mt+IIkLAs9g8UDGSXeY1hhD5eNUdCkK3D3Ap9uAJQ2eomZ
l7dnmhzU1vz+u7ep/+BJLHHMLiPCQ6saU7fiT/4ZvqrT9ZCuUmRX1mWTdutjD0wVlGrO+7p3ThhG
FGfRU1DKdfE8Bmd0smEkWNuFVjRYoL9/f0LtMEEoQGtvDnYTBkMZ+B3udEvVFy1Hqwn6udexok5x
ejasNw6y+NXChjYX0385T3gGe9vpp6ewFQtN3Nu/y9vUCgzJxHwXHnESU6VBOH3LG4LTIYWg/oe9
fCE+qjMOsV3QTNYvU/FIIcrbQWtjHNAO0JsbFDFg3W7Es4iiitmKau4Ts7SRS007h3Asfci7/41R
cVVjfSRAzxbg8YnlWisg0CvExIjuw6ceKVXWlwaVM6VnRbwzLrH7U4RSjPofmIF6le5dsgHSROmM
JwVMGorPPgUo6YzUEse9Fy6SxKpnILxuLGqj4yAYsZgunEI2/4Jtuzk7absk+aUHeFJjdqE1BvJ4
Qzwbv+NUWHwpnT8ldn06yiV0lHeq77P7Oe7QycJ4RfzMpE+CXw4Xn/0mAK3zhaNZyPo524wWIelU
tT+G+jLRJEEhVwjZJ3yIbaBGoZmRCR7AUk0nvmXgQWdYGPoU8Dw2HXF5Yj7yk7VL7qVot9geVw4I
Qzvo+D0xQ+HY/NPadSSPUkI3wQ7mXszYAAC9ImQpKoS+pM83+ECVMJ2Dd56SEK5/znx8zb0Vgj8O
5p2SNc78ikcUputmSZHVdaATyOX+NP4hjXet4M7nng2CQl4dgk2NR4Xcmu4iP7tpN8sWOMtwa5f5
KBj/b9wWEaVogbWzE5Cda+RHbAQfAGhGMdj4zxlnr4RhBUEc4Hyh2nDL6Dqnx8eM/+rocACckyKN
cH69a+P4DVY3jvXYmCyuSH7LYYAV3UeA0m9atE3ZqT9UpbmI49MJi9Sfx6r6RCICg7bozn7HdJTB
4I/jbkEgOAV+66ZBoOhpPqG3cDMQtUPR+KzT2Aoj3nkDFD/hVi6wK4Ip10w2xfngOlE5PGwavpfj
5CbmmVF5YEbLJiwjX+wAZ6GZfdqRghAV1X6uIDmc13ZDF83oraFwl7esXbhUCCxx8r3zFx+Tj0uU
i+UmyjKtv4mi/R0wvzFqwtTVMdeiVyHDxgOIVYAopVsvUP2LCRqyG6R++uflKwBB52pBiYfxxW3t
Tj6hJyTrpYAgBIcnt+Bx2qpKH2JJSZr2t9SOr2YlYGXn4XPVky8HQ3fQ8QNQc/dOAh9TqY9OdmmK
73Di42HQHW5ULQqr2VL+Obf81XRtt0oTD99Q+n/ZprMd5BsoiY/rB9VHFBMceS84hY6mWlTlcDHM
OIb+1OUz91sSsI8YG3KUj+LwkHnr4Gk6nEiM4fbSe3X+CoUHyjc4gRg1m5SlDNa+cEZuko20dYyH
h1aHIadz8JUD/9qztDI1hZytgB9KgipGovV/d/u3ky3caou145JK4kDsVhynxEZ5+zJ8Py2s7amg
vUv6NiMfVCBg8FvdZIDMWxP7KnYg0De1rXtm8/dAZP4ThTnfbgxCICP5dbC5tVJd51Kcm30VNMx8
isrhAcAnZICC6moYRSFa24bKDcZ17GC78foQqqEeWZ/n2wyjINiQ8a8vdCK0Ti4/Stfv414jNgrx
mPyKVPGl74yMJxIPOXhhaElbQXzttXgo4pdIxwlWMGQjaTVf2MG2/iYBEXZE5oSVYtDq/BeaeURJ
iBHFNFH8SgE97Y0WlHMKTr2GpCjsdXSlKz88PrAwhCYlsvDYfJYqM28/kj3kraRRJUasevHv0PxO
h8epVecRUU7llIUGwNUmevEO/1R0f/IgmyrYgNl0C5nOm1d4lGXZZNUI40x0hWs6AbRLqX41jnjY
g4XOBHibpHBb5biivQQ1k5not0xW7Khg32ULJiBE6NoVaNu603wRWVIW7IB28uJPXJKS4OyE0aJq
J6MpA1I6lD+wdNiKlxKrGKTK+UDrXxN1o+JjE7JMm1eW/eQ9V7tdvKp5LgpKrNYkR2wh6B9wv0UO
SjknL6cvoRffbsHzVpufXJEzIFzZ9wKH/VsJ7WR3YxPZyix38LX7FE9JwhHjZNGqxUthb36IKCYP
ZJ2SozscVu0hgJJyx3nciT9mZseTJaLo/+Z1xqUez5dveHXCOqDDHI//v4DLICMu6qUPYQCqS2bF
QRSyCA9aFByYNgx670khY54sxdeqttDQiCOnGcS+VC8fnkcsCCvPo4jbqIUgfvpcg5fYrzmUc3E5
TjLt56m6ewOp1z0T/BHkP+Tp5M+gLBoP8NOF8Mo9wDJNeHztzNwmH6HazLczJ1o9G2VLdcmU7s3y
B8p4BLWlI4oB59JMT1HFtfy6aThIrFQkj09GUoTfinuK4nnV9Uyz7sPWi80EQUM+gFlKFhRho8OE
LwUEOzOLkc5mfey8k0sj3wMlr/C6kQBqQZ/dhij6JwjA2bmaQL7k5AsHHibqFwTHv+WO5Ss3Yrzk
Dvn7QcH59Dvg0I6xCl/YhPQeF1uJ6jYbFDAdWmPADX4KxjDyWFDJkK8WuNOv4BduHf0Osz7gS8/l
aVlbmLdQ4QV8yC87VxIkeBMaPFj1/SS/gIxjM+zKV7/fwdwzixk6hCcof66mLYD4WPp1JV7p3V4v
Wfwc45dhwT07N95V7fCnZuRGErR59u2DOksNbunmCVMuEMf8L+22AQdCVin3lsR8Z6FBcS7WZldj
SQLDrnO2XNLtxePifu+njFTJiy/KMhcUy6pCFICeYZC7IPuZc9v8HXoBXm2CFiQOdIEqHDES1mGv
TTuGyZyFVQBwmLEXCbP9394/ImLzceJkgV1zTeZPfQK7B6QgXEqjEuHjVKCpbKXWtcLOTFrfo8l/
3izOslWPY0FqdLUdPVZh75hb3imKKNx3jZcOXvE/syENXTSa6uqe0k+LFNvcRrpPIrExWPCsY6Tn
RojuM5S945unpoXRtidA3wDE42Us3uZacR8/6f5Wj2/qCDdeYvNQAF8JlBSi/KFT7W8ZGz8oJSCH
nv90TQ/cyCueap8rwlgT1u2b8f1CVII4MDc9pDoW5FDJ2riLjdeTXs+SZ+zSij2Flot8bPzAXnDl
EAyv0PLkr7kwara5mZmBOCOYX07gAT6if532xr/VzklDhG+y//TFcvpSMbQizTEEEI8hnFFQ/D6R
NIIcnX0DAXsOrnvfD1p6abusWZeKG15um7HM+pPQnUZBKmB22bOaxN6oQkuBP1PLv8KkiyqR5wu5
RQloNF8sU8Rz3LgmvccuwH1uMLhBb1B5SJKWfjaiQVkNkNLndqBW+eJfBrVLJiQMh6tB7/hgXttT
2uDNuYfIqHAeibwoogdAcWAxBuTiQpKLrwu46IiDMnJlk2ONjYD7iWO4Gv/Yh4oqn0XMtxmVJ2Jt
vSB2kVeGjOf+4Mm53M/OYwCyAbOD/7C5OBpbaaaJhPBCePRK1w9PUlFfNtUr5bgQ65w8birJNsPX
RqIEhxmFNAspozSinB3gE8qgA9EvP82jerCrss0qGZUqqItn9IIRcjeWyIk2lfXPcIVySS5d8P65
mKfx5Fbz1+U9jjvO4HiDQdyLCmdjjMGfBFfeXwETcqgwuOcp7dCTd8byOC9cfE7HXy5VK079y4no
RB3k9POGKKFD9gX4OQOd63+XiemnRsqsV2ZFIrcWqnBN0eIdOQv/VfdVX/vmzi+LJXxD3viDZ59X
hnRE9zrEv9wtj0vNDPSklwlU7zlXMsFomxoScJIGPs5XEFPEwyjHSxC+suWmcocGLIgFxhy/8Zzl
BW4NUjatK7dNG7THXChM5ifJwWAAKRxEREqEBNnoF87MAuJjtcdjDSBubCrM6sg5bW5YI5S6kVc8
a88JnLBv6Fkcv65f4/diyaHWekWx9WsLWJGRDDqwVZF88UoBColYJUbKkOoRZNdSiHZwbdaBLPRV
JIRm0W+kOsg3+kK9bMoCjp8aEBSRJ2zX2dR5gtI3yh/TjPgEkydYVeX2Tiemn/4kCUzMTDoR42KX
BkiJSOarIDQCZnfh0YiC6r2v0JlF75Dv8NH47J4Jun5Or10Jv9NQPZxZ5xwQigElzDfrvCN2QgE8
L8NDDjbEC7VTr+GY+5U2FibqqsTybZJqOGDuK7+WpUNm4+yIOaAirFTGX9zhaPmAzvTdKh9w0Pku
luZu4I+HxbWMVilUTfG5sP/O5AhEzIEad3mg5fvhG8cS+6AWZyciy1uZibGhgTafYSJsQXjkL1lK
0dXGH3HoFYdQ7ZATM+f9TNXbI+02E+n+wqKa6s6oJNQJWQ6p9nFjIjC0UMj5qYH60XLypRPVUn+g
H4NlfTRf2g4Dm9l67a6YN5hJBYQUGhliTynVX9sY0+FJ4yndV8Nhr1mrf5OVS1hlqep3nSw6Xnvz
NvEdYAPqZpYtzGY6DfqtUhzVJhKUzKKG1BZMR5fGV8v6jwOWFXzuxRq8sWS6Y7cT8vKFBRrfrKl2
Xi0OYib1LODjjFxBKl5xiFjma0ja3shRXQS4bbvfKS8jQ7I4A9tp5NSsk7/7AISno0up4D7AuKhb
pdUjcq94KgCl92ffSumsUh/Mw03KJETiWZ9q0109HYJcEhVw0Pr4vaHjfA+vLJ7dw6kgoo+ahbZj
/c3miCUd3nsuBqW9IxXXqisy3v2IYb2idkQQd67nfqKzGf+fymE79RRgHmTHimUvp1ReBqgK+9mE
O3aO1+HuuN5I2qK2ciEuwdWpCjrFKPFtrOAHn+NuX/iax04EcUROXVA0qwdxniXfBQyz4FscukVx
ni+RAJrneaeq6L6Vi0kbVb5FGI7PT+sv0V6scv6La+sH2deOgO68FD2y66ZLdJMbjy3n5xuctKa/
m8LK5USebD05mzTvQTeyR6+fT/XOzd86REX5z6RX+k9TMqUUgbMz2vRefm9DXgQFt5PxKVkeJ8J3
hLSB671V95d1aeSbP0A+okx146HKLUSG1+H24z+bEjZdd6UzKSEyK8YZchcW4JxfA+P0zJrFBbQ5
6y5oLVu03qHLbGTYs/X0KPO2J3dYwdy/OTu7TJ+VF9cbWQnXulkqx5EmLCP0MTODsOg59XRFW8Vq
5C/S5Oq2Zopk7TyFnSfQcwSetSROERZQNLkHPvAKSB+61XcjU/Jcp6FKkM3X4b5naj8TdHex8CbN
FTGUFXYPia7Dg/3j1d3UtoJblrfupP3sBapE35j/fXT23WV0FFUdpnfBmVQ0h6uhWXqFagQeBezy
3OJEGvPC/tMZn40iyeTSeASFZIh0RhpQNJeSGQ5r/PFIuXzbt6HkqSu96Cr47uoqIFzASRKkLx7m
12y2QyyQSPRpWPHNWLYFdrM/ANdzxTFlFTuJuSdMNspmvxPoraK83CFjY43Qzd/sHDjgFUZv5Wf9
q/PQU8ac/h8RFYlnZZCVlOD+eQiqgyMzuKhkv+ZGv+gNNNxNG8pzVufSh7Gdc1ZVmN4PT5MQ3mH2
c8x+38MhaYphzfqMkpSTFbvf/iMKR+AcS+/49uFDSoSYFzJ13qr+flfA8D/4TF30lGIf8D2xWAWD
vCNtjP9yLlpFL+VgE/iesTFCEcBgtwY5AAUltMEjvVBsSP0BEiQDh2Mq+Y5YZOgEueDJkMPsuhWV
Aq9F3l2BBlYcoLzjcSreuGqGw4A/cZMcMnUEV1g9I8mNznMaSPAKua/TId2A/gZfnpT8A/dib+Rz
q7KnaUNBFuPEL+1ZO7WZjHAK2H5UZW953W5SQbh0ibGP+pzlUPb9Ubt/a7qt4q8FvOY95+XAOwfp
FqI9mBePI0+PI7xaTl0IdX46SQwaVhOqo8H5AviZ9yYJBQLDoYz/qa/Vuh/FLRmHvI3GL3p4aLYe
npV+VV0MA5Hk+to3UAVaJpx05MUkySDakI4OloW7vNu/DHMb5Su949iCJxNDdC4yqkkXvCKFowfD
Xrdtz+Z8roHeetSKajTO7xwHG/iGv/JL2NtnxAaslRyjIECtf0TlGbqdxvQSq7YjQiZyl9JYVkSt
ksz3lKfy6SKyhSEcEkbPkIPNjW7tiOZlqljyMpZWxlEpfTAiDLX9R4UZAqf97IazaqjsZ8E/l5DE
tdg1JMIEcFzNJKsVPsFxpxS530iJgx8EpkoGQMHnOyL6hqRvDugWrSU6vxWjuxeKwdwqMEmitIqe
PMfxQ8HfLsl2TKNN3Ys1GeJCTsdXkMCwTWdE4k1YwqhhpjSu0HmiJG+Rvij49IU5xO+i/zEUR5J0
BwRuQuXNfVWA6M4V+ikq4BkTottXq9IlFRT87dE0pyoxpC05vVP66lTR4AL5lxB8+QdWRmWDG+Xg
iGcegYEofwm8holRSYO8W/L30Ywp/3iSfghBhV7mxEmJeaqun3X53v02EjSO1rE5Y0bAuKIi1NaU
kIyrqv4liOt13BFrKHPxZ/P2nSKVDRZrhIK8Djb+G4x86jFqQInb3t60QvnJcZM4TIe+/HSBNzp9
FrhV25VMSpio0M5DD1dpVRh4m1ZHYLnFuBizGh2bwoHTaC5YDTN12LiGCgJzTW9eHJLXOVdewua8
Oy6pI/UmjmSblz6u0SxL6ghec4e2hi8r3NCVIAoZJsOuhnVpntUdWgIusgWktnghBxZinR0roaQb
E0lV1y/qOrcCYH3wiWQNznL87l53+v8v/Yp27pM/oW6AFlpcxxgLsmX4EoBk78Wk1u8PH41/r3Nb
gPaTEOzeQ8p7mPzLMd5jUUxJrQbUCTpd7tY0ywwH/kyCdFGwTdvTRFRyF/E1Lpd3P8yD6czCv0xo
Csc9bDvulnTviueaKsWd/BOoipJQDzhxawpNUjBDS1RGoHMMwQ5XYeDig4wjWMWpwDDlUk+Yc7b4
DxMHbClclvqnB996XiIjfk73tCSJqgDvdTnyaPf9U/QEH6f7WqIKbaEaQKFU9PPRGWmht+E9Zmrr
WzWJQ9n10cbTu7H39dWruRDiwtqb+3vIT5p92V6sIE/cGnQGCje90PmNtmriTVwPNKXzmFOoIkER
rk/INb7VNxjh4PbEpoK8A+8bClXLs9PYB49xiwvNeHFEK/mWPmpElwW7xXEUdy1HBCa8peZTKtny
sLn742UH8JW+4w6vKhjFSmYKmafkyrXRyRg9jGF9yzaaX7vzy+focaXbmXEAxWNZOrQ40qr3ISjo
o79sUJiNzY9pfWTxyp2VAHPBbnfDTiiUdetdThSNb2CNPWiTrMmohUnGcPdXY1gR8TX7nrTAGLTt
RLrtfGgeXXWMcGcONG/Utm2j8TNGPG6OJEHBwchWZum0ErdDtjoFAnDJBJsW1LiEkBT40NjyMT1p
WcEStlFVPuBmbPdHxEJnbSoyU1BQT9iRQjIvh59CD/ti/RpKXQX7e2+wSaeuu9Q3VTUpEEGH5uzw
Y0N0BBNrxrryplKg4g5iZcpWXnkM331gC+TeyI8YNTjD8JotKVf7UZX6A9jfVY1iLCtSfGa/mHkp
D4G0Utc71N9jGWLoI0hklbuuwDlI311p51Gkr77kvATLzeC3YmsO74isD+iQVv5g3QkpX3WNXiWf
nK1umGIcenjFBPiUJC7Ju49RHTd5Jfwznz5eUoSwccpJfomdemSvpXlMnZBg6nYWA1/mahUVcPDN
t2WL1+lt1jMFbCCksGkXGRMUmFLgweCpmIqjeK8rw8mN62Phn2T6/9nIMXO9TEKELbexf6vKdM4Z
TOfcsuZfw66r/lV53aCBMT1SiSHNfz+1VA50Y5Iue/wCGQZfTCQtuvrrVs7prFwM4j4aHZFbEvDA
DJ+G+B/N18n7iySNMizS6coNwBaN1haVr3jv3NdEymkdDydQIm7D9RHZEhwFtIoLzABbK3e2mxZJ
KwNnbqsKv5504tvclXt/Aw2WBQQaJCszOaOkoJ3SO7g3H0WOXTQn6u4p2F2rVfUqfT0eJvKaIG2G
lf9St7b/lnFWJQfrUB31w5W8ymZjXBZBS7n0OA05EScpa9jYVaLmO8JE3FDLNPw+eUuPg66VULEg
gtjssWdna+QQI4qqWPWFttEjVVYTek3uNdVYXm2SJm0fAYx82cdQPEqjd0O0vJclNNnnpU39Mopo
EcQvVAuHFzFYXQ50wQZ4X9TDfM+U9rei7dCD/BPdZm9YxPU8OzfhBC1gH7PBh1MLyzYycYs8HGC+
4aJ1QVo36VQ2DFHW9NxD21g5afWUy8pLrOt8TD/Rlg/DC5TPbxnnB9gw9lF1vHA12JLyciUh5iCa
Ot2OdBgz8CVteKg51hgUNP9BAqMAsG5+EUYQoq5nAG8PmWUYK8MvWvfHFHogcbxa+CHy6Wanez5z
YAxIov4JqDGRTMM813eOSUxRB/8WxGNk2x7v3xjJB4ii4PtaAY/qdlDA6xOHFpVAIeFxfCeqVDPI
4gnJY7T3vdyjLh+hGF+JCzLeKIsfaiV5otno1tPBjqnx5CRKoJ3/q2pc5fAGRi1BEh21BGi6KObd
Bym08Aw2b5nbKuobzNNfdM8LjHFDV+UAi2C0TBxXceUrQ8fivtw788SrOwu0JpAsTBFvWfBX2DlB
+jA2vVYza6AwgvpehYj6D0zmpPA9iRIBJ9zFuezAfbfa16EpX+id4BgoklZpngtinCqe7WdwCj+9
KHuIFSyjPdae7fWImrz/CL5prLn+RdM1tNFPp+nw/RNQlnAzANpg4fk5+jWw+g4XD2xAmHLdNFBC
6WU4UNdSD80PNlom8YAw3Sb+mlnnKIT/E9DE6a6B7XganD42YNm8tHU+a0jGksCXZ/3Ah31Zw8r0
d0U4ab9bd6EDYQQ8FdTsAkxHMw4r3AUVjGBKShwc6sh5NjjmfjzBWbtuvvTJae3VyhR3f+FeLjcY
w5MrzOn+0a8EVnUeTeYPkronenFikImb5jtn1Z9V/0gKZW3ZiqEuZ83vBHEwow+1XYWVGuh1nJzV
OPsOZH+nc4yLiyBd31FQiLfn4JGIvMiiBgE6J012RzVabwOYaZyMn7VfHT5O5Oj5w5aTUxv/y2SW
WBpAT9ml/3GZp74Zi+7IBbreNVeLhoc7vSVEcDy33r10CvKWiD72mUiwXg+3BkZslh7+4Y0N7umD
RhUqA+JkRFhYqelYOQjLcRkXAQQekoF03lAgrB+9NMqkZrTwzMa02AGsq9glRZ6bjWqW315QaQ6f
XnFf8w80LBPYfPCtsCIiIoM+7uvnvSoZ7Cp5qvNRBfwer46tSwPB4g/AjjTm/YNf7UZz+FxxAFG8
yPTO69LIuPjEGIEGthHZXTEEAP3asUD8DEMhvoNTZJ1oa/+GB8DjLyF3hEyDtAV1YOsVj4x8R21f
WGoBxXmumd4HdmxBETAaFvY1iOCgNbvZ8tIsoh+8hcB5iS9/06oa7HEi1H1wW1IdMiO9UNLQMykp
9myZByP4bZRk4LCKrknTWS5zYP7+h7DAuNwFFkVDGfoXfol3At9scicLbmUGsf0qgQhzdGNs3sBx
NtFPgujwgs286yo9SUvyxY6RlZePzO5AcoJnb5zXmFQ+mHyj3lsXxs7gfiywW3InlgeROesuL1do
C9IvEUBUn1FSiYq6+obh5o/J1MyNvhdVEfLL415FSJvu7SUkZzurRTeYC31b7vKS6seODRUFSq8g
viqpGOlslWlR1/7Nf/6kEhePaMfY5zxbBf1jv6KWCBS+ZRup483Cdaf5fc0315r3MlghJ1Eimyiy
rF84h2eMT8Do8yEXT7DLp7vCzPRVILCyNAa90yWZs6Xt1gUquvasbuRYJzyFHE9VluKhtG4BbLZ9
hO6i2XM4bf7eofuxoLdw6w35ZK+3IEoQtFFSe76jNuCwun3AUvH8hCVlEBkRjEvdSKiSlk1sMebI
XC1Fcu3sAacGKwbKswAxnumJnk0KRqTD4HWJ+R9NMf/6MncVtTf58MQbvBpgRdSjzojHrV2Rc0OI
Mb4bYUZODIi1VOWVvE0/gJwC0wV/vVZ6UYE7FxiaNT7FnZG38Sc+x8VQbN4RtrzBojf/kdO+sNUL
+KJo1qVZJJIWs2NYHuweiDIUDYfRbWjXuIslcX1T0BknX0l8wHka0DrisyGmNYysaAkRTVEQhEiG
p4QGZBvE5dpLFVboKT644eMqOlzFIXjLEQJzgeppHvSfjRz1rwF10IKlnv4F2qwjPi0Wxa3S3P+g
KIX/qpniyuKPDHugexkOqQvYwyG0HXjqfHdE1cUhiMD79Xqj5xM7YIGQvodbLUWej6OySJvOF0EA
P5cBApn/eHQikqVYiW/F3VGpIiOtcbC2XOQFoki0hVDF+Fc32J7UEeKNM0e/LRg4d4kSy4POZcyh
+S8dz7ARABShH1rQzUT5vflcO3dqgaUF5rzrcDxuK0xVSJMgNII+QwxnZr0yENcy+h45gaEauBKm
ktGbA05fl59CT/F9v5HFfpJQekWGUXBNrUhAJKd37Ujj/azMY0FczEnkiM6K7AgQjnGRAXBjxJzR
ChghDlqDtuRjwf+s+GpvQCyCguxjOp3Dy/m7pEVa2XOspfKvzHoh9spFF25SmrGREsVJ/sUIIjbw
N1x5mpEa8F6PG+aTej/HvAa3z+9QJzR+xAKPw4PS8agNp9gIt+RDKdRQhI/5bIkoEh6kPtrI081L
TPuMiF1Kd8cWZM2ZBu1D/SExctuSZRXeXfqJ22h4eFx1KxBGZK22oPCfBAD6ZePju4nbLq8w43v6
ln9Fve+jsfkIPrara0bVMqBRWieVKU6aINu0xxkBLIeqhDcGYy6IvJg/F8PMkTMPWoMMVYm/vcjh
mwapVAPPFGw5fHM5YTzFeiJRhmxeV9VWvHeThQgZstWgiaOwXAwC+5pX6v6zGoqmb6sehMSRk8N/
UGUBLtXv4iqgodXof+ksQaLuhvXjAy46kUXBdz7S0WukJAjF0aWiE9qnof7Ap5vj56PZ4fbNCdBn
AxUhuuepBjTj2Yd+tUSSx/sxs/5UY2Xwj4HUrXmz5jJA+zAG93u+vnbpzDGdx60f/E954pVSduL0
vS5c3xJK7WJ975+uFNJKq8vOvaV15olv94v17DdessL8VrtOFqxwl6vBWOcuccNgIKKldZdou1hW
eDeR8yVrwFf74KN0d/BY5TRxZVNY2q4nFtPn/wYzzQ3PwqRm5ST/COStjLJIt93t8LcCzS2E00d6
aJPcywFelaVJU8ckWn74wir0RZ4z5jRxuJ5lWMcz6CgLwAopWF9JePSbmvRuFtP1TSgMNDeNAK9J
Mz8PEIgSJOlb7H7Y7lQtyDQ3UF2lVXHMA6OLo9MjWyIpXbUQsMoXWRI3GxouVg89AQbuNhB/XTTO
+G3LLjXQItf6jiAKZ84+2rA1XzIDg/b1Blc8nroNvLUyAHY5fw8je2qq7CSWNX33tLgIKPwXIlLE
YmOZdRLRTWaDmsagZSC0ohAzKp7d8r3TJKuywOmlvCVSRvDyb2RAgOnRx1YoX7K8JdsZwCwSBnRS
NdPNKR51vH/k5uXvjNpvNCEEPSY3sO9e52dLeoQROJn9bRRKc4DQBXIigVlF3iVeoSRPD+Ct808E
IlGuiOh1zm7xKLxh8z/MVYkX83Sz/rRtLHmtP9KswlEp+5k/y4AN83RqKy+W5Bm7o7+srzr1f+xW
an3rU7aWw4FGXsbM2SNv0z2cKPaUiEoaTsY7b81Mkcp54ESjjeEeym9SvSMMqa/iW3kjr7x1Sv4o
SLeNdVMO5RksG0gl0h/eMuVkAqdVZi5EJBYNiuQ38Jy6XyvLh9J6OjwqG3+EI21xQ8uuymuTJygL
i/y4nt63nTDua6nf66uYwstnXaxe5Koj+mkr1kWWK1bkQz0R42Mt3/KMeUl8/iaWMnSzYuXONdEl
PqVC1Cf1bNu+ycgnQq0nJ64vez7RskKFqRCe9emrehg9VQVGLsrVJtzf9DoU47ujb7SSE3jAi7TY
ZxjdrNf0uN42sAj1ujElHhBgVCvv1/mHOakbTs/8NjKNIMWQw3Y0iwaWXtSfTWzTjyUlSiUcCcHd
72gMIPxPG2iLIngDgSL0ERUP5aZrst4shEE3eu4eMbTvJHMVELZzSUmKEPJMUVD4AXXjNLI+Msby
ZyPcg4SkfF9ddMdFda0O75sA0OFXAv1wqkVdpuZAZsTYNBKwDIcXpIhcgpi9DZCDPuG4eTc4pDjv
DeqtBr8xCRg4Zp+ArJq5eqdPfF3GxMbyKHmYuwvc4MfxAHtyBaDY0nabyGnLjJ2JnfNyeywnLN8N
0lnHykfLlTOTkiB9OfDtzlWqwgSvh8VMlBvhhj4V3bpPZ5R8LPnsaUDi0y+VHUaAr5swqmJgvCpI
30RRB4CLha9iKokRX+J+b0XLW7vl9ageeyC71qWflVehgkLzGYk7N4q0osf1gemFfXL25Ww76FCy
vw0lpboxgBMj+Mi6g5e25FfEVsNVDy1srJhHXJTvKIn1NhEHL5T9xsEjtlbDXerejhcQnL+SpD8Y
MgGVNJj2FCv+dQTUf9fUCyNPSo5WLShJFwmFhTlMdULpCIlPksMipjN2KnVFB18izoAwuFGhMwVp
q33Bz+w6ECDBOjlga+msiL+GUulfNA5FZOr5FsxAeDuO0p8pZjBfJ2xuyV5p1mC6BU2h9LC8sLco
y+rTGWpIR/Zaf7QsWXwCqhLbLHKE1U9MPBmPSVrFQXGq0tmfeopxh8PnImeqYkltm781zW0eMWvp
V/RjIsc4SYKXnEljy8WB8zjZ1TBiF2dUS5xjsKFPEutvc0IszqOq4kWgJdCNqJdZvegjm4JFZO6C
oZ/7jZ9+xifSXyC5IP7MkVgfKX8b4QHqljYqWcnJbgRHa0H2PHLfXjdcIZmRPQ5d5xUJiyFDEE0U
HMUyN3nak0AtvA/6RP0uhpV1yt0iHKFmv2uu4iehKQ7LlWZO/q6yVD/1bkErFg1uagENuTysl5pR
K1kY5Kf++cPDdlvsrhpnEfLEhf/9RJs1wTzLcO4kJAhwQpg9ak8+rqiYWgox813/Xo1GkwR/mkkZ
x2OB2ScShAR9dwXdxLxKYYZhYXvhX32tN9jEYixkKFa8BtP785BRpwtQpglX+TdvF6SRdFrvR9LS
VMw9Ypvv4mNduv4IrW8ag0R5rQm98qVnJzi3T9Fg7wsioUeYICtkBj+zaNt4Zoq8hSukKRANimPZ
50eoDoMQLpwbgIcCNx70HzSe+9GFhmPPsombDiInnZgrvLsFe67C594sjO6hKEXdrdtDEOL1U9Z+
1uz/f7uJGaksMXTe6l9ClA3KpVWlU2sr7ZmTrkfyF/0mp+uBG+WIZY9Dq3PHK44LvV1KkBqvA0QR
7SWNO50bOWm7UN1FDe+slPvLfce1MaBvMy6aIixW98I2GDSOwnjHcxk/GbTF3tGyfdHsOlzPbW2j
WpZBM5UT9pZeZRHd02xOkBqN0QFkb8XDB/RdJH3G8jDL6YV13OH7oQQ6Me6d+yYsAZ414Xetv8Ok
auZ/HDht3DL2vrF0+92xDVM4NeoAfXKBAn1GdhHHvkJo916RXS2OtDaQwi4e5BFKdrIjKw4qMUlH
qgeoD6ncfQW+2NkWbZXH1WsVuWKDKBiEU/qQSvYAA90AuBBuufrGC5y5XLC2W2wOAaERBMnLRyYp
COEv7SRSQzUUOa56ein2uiSSVXnogPRWxY/Ax2Bv3fQo/tq/jHvjDVoxoU7/2EztGT2ccA5WG8Ff
CY6V5jBg2KLH5jl9ZPaCwJ7iGLv1q8uxD5024n+K/mufhi/PtTWOwKIENkRXHFN55ZLvJ2+nY53p
XWNO7KlaDDCAuCaH+C+PLJ1bhmkCZLTR/gAajwHA4gAXOKioS+J2FXTnZi3cUxzP0iW2momcdzVW
cg7GWiR3EQ0JPWeuHAvh2WjmcWrJ2ZoRBgluIVDsAt7K5JQpcHpdet4WeJrDhTsrbGXl+WNHTXLS
cAVbY4/2Zep0sv9bVeig7qGM2LnJ4PQD0s6/tSgqPeyKm2zHzMFummn5GOUqe9Sq+POncbgP7GbY
SlE3hDvTiTzzdfxwoo5jgqbGqCNeKuuGfyTBqwazrOBtNRuzpcuu8+HCe1tJU/4OEbSNLNkwJH2r
z+Rjz4X/qfDvL97ySWBOAtnPnKca9fCyUyARO5PNcRXaIXK96cFi7gBjAfBk80DeCogtrLG02iud
28g/hCckG93l0YB89QjUPOn9V6J1HRViZfbqgvre6SDMXXNtr3AjwzzGezmoKMfzc+aUVNQzwIxu
yGOZU9aLYJjwTROe6re4NYkH3WGdiOnbuSF/xZ6wJNgmI+Pwgb9q+XVnBLmMANTWrKVOHKCG2Z3U
ZCUPc4DAKC9nI/SFNLWVH0U9TDScH6OhQ2jx+2KJB4P9ftFt8rwEVoIoWclVC/t5M4YvjUetE0B6
naoOEJrqRqBk+LEKgC084wlgcoRQAdDR6Vdgaxm6J5QDALKV+LEAsdr8ZfmDm0lNGaWQES9Y3UNg
afW7C6WvTXSvgkUN4B0CYi6OZd0mmDfCyPBhLokFeUCcVpoTjwmBm3SquApiPmGNX0STCNc3J/S4
Bk3EgcnWk/JLlUHTmPY+wscgqXgPcEIxlkdjIL1pAN8QCgwPHikOpmpmotPEUWeuHfbSiEdAnIGs
zaaFvVAOz6YYgHKf/+fBk36h+n02yslSSRMc3ybXno+Dh6qRLDEgkuIInFhLHMrLXs8hRckvqlel
jsYHhsV5dqIcSAbOLypwKOwOAWw6yCrpAVP8iXNOqoHsTYd4FLZ00Oo2evLpTElV7IRV550VPRnF
Dw+opdjENpCx4DvSfagw9lgHgEJ5ugPp13/nqy29i4l0CE7/G+3GJiLreehrlAN69sWzGCEHXK1m
gAyPhg9PrsuY7JFJsA1pVMC6JusimbqePo5XC/Bc6E+koNLWA+iBzLrq5tx/BcETfPD+aWWHW0wi
XEvcLoygcLfviR7smhZw1o+hFjioU7A9kC3Elln2Vu3zFA3dcs60X7T1gM4xdH4qecIwRsuUkBRR
0jJq9qrOQ22MoE2MGimLrtfRc2Ib4YSWw4ZoKrVyVzi+nvyGOjTbOemeLsaeqx91OaRdl/HbtE/T
puwZLSwaq9hcOc3td/I3iA/9vuLxOGhWrbV6UG/D24wU9ECY0iF7WwKKnMuaL5LZ/9oSLrthUWWa
FzDAaCKxz3MgwiUyzt4v9AOjQvfFZLIPTWQ+9FYb4nqxWTUah5GijfEkAr2RtJ9WOr6sbMXocJmS
dJpvtm3FSReqF7r4zd7QZjLSIPcY2M+EN9hvvdRbhaP0xkrIJ/n1teXUVpM0krZH2wDFkpWRALWc
fOu1SzMaTvM636QMbUN3tI/65M/g6eqN5kIplFw2m4wO0QtIoe/8R4MgjKkuK2ZP/Kp+efRls8WL
dCLH/VEC5yy+6t/Pvzz3sugnxc2Aeb0EYZJ9yIhtqCxKTIdBDMi83IsF40Sms8hhr8ckrnA4MZ6m
XvDEiZ99hskE8LaSHpP8z4I6n1m70clkSBaXlTYlVwyn+xCviY2/vNnfq8Kq5zvlR1Y0Vi9uYBsP
X2j9DgsGw4mCqmwgr2ZHSmHC6ebaBtHlmmjMowcgflDM/kYCInFAyVzUEztHOT6DyGyNZidVfT8e
pl2gfJOxSvcymGukCTc6ovfgI7i2ycfFEyxM7cJQd0SHII+YAPVR5kxHgAISvwp8vcsPNB2XtMWH
5QItzvZfPKahWlMJjJOlS06szeCjkPtKdqh5XiwuquAInzVAvAWH//xoZ+xByzo/v8/6BSRejuPG
C8gyvC2S7+Lncnx3fXIpS6OxIvvFQ66JCpUYqIXU/pkeBz7cfHq9Pe1FP7XO1TItJ9WYUHmSvWY1
/uKExZPGo9zgE4e3BXYXLma+RrY85l9aWZkSCwgOSjtWcYwXlUlZMCrgUf5Hj+1cgavwPeWFAFEI
thEYOT5otN7LgTY=
`protect end_protected
