-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kaCYPH0js1VTZJe4MKyEoKMGmVzw1G1ef7wbvUXT56ThRNbocKqVUkrInbRSFmsM04FH1z7w4aNA
4eejGQLfSRkxWoUn0Ehw2nZ2Fiqcx/DqtEywCv+S7mXmgGBqVOAdjO6TsPbpNnlQ3z+Qmlt1mNY5
Aphi0ICYCsLBZ+nIf11JGjR8B/dqBqyU+lO7lSl4jDmP/iAdkc+v6jheXrgXT2EIDBZRENVIyWFl
7clK8r9JL21OXsGu7H7qDo+ozPgdytTdIM2JhImJcf1YbBTXBNH0oG30pD/YmBpTeY/pvhapY4Yg
zciWrr/vK0j7W7ENGrQbS38UrDbikW7bf/jd9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50576)
`protect data_block
LqYpTreF1B+p1YYDsn7bdWoEimzZvYDDqFuZWkyktU4ZeD94xVL9LWoNt0J+JhevaCY22kNVZ9Rp
Xtw0Lf0Tukbn5+XQq35YUYlo9Y+Wv7YRoS6tP45gkaCsLx1DArSOpC9K73NLlfqpuYsTJJpqiuhB
rINtPEsOzhUOI2LVyzNqZYOzSKuonEwkHMqFr9YayFyAq7Yem9hoa6A4tV0gnWB6N02rPIb6jwPY
/X6V9sN3KMeMWLCIqAHsqOIPz81bV1zoHhmHqtac8pBJr+CsIreru4tM+8cwKDFl1ZJRPDsgX9jz
Qp/74IdJRLgQlTlvFMaAI+33f2rBgVyLqEFEYNtPe3A8txmyCT+XtOzkMcPwPuhi/rBvi2CZAJyg
fY7i+LAFVlpUGHvuT4dGHI5NMOqpuYYyCNpg19Gpc5bx5ypZsYjoDCbe54mnqnbKrH3p7bDXFgvt
4kcR+3mNKAWAlm7A/N8l2chgcGtSG3BcGJUKTBhPVQqfthfKPay2tYMuXb10wfwZpD1i2M1Zq7yq
E1pWw5WjHiWv7BmPoPh32cC61bO3dYpylEPUUlxDeviF4S574fSS+ZJ+h3Oz5PiMSFl4snuoJe94
7Hh3a56hmvTQ720OTfGxX2/vpr+yzRDk/bamIXcarzeeRi8J9rvy5AK6EyZ1Rp1WU+Ith7PoYHkU
Mp9gv9qZB1qcLsasrgh+V5YfXLIpA1IIkHd5Q4fFSeqFwTZ1CtUDsOMxexQArO1mBdP/6KoUBM5K
xS8zWjmiew0mV7i30hFvDPmN4YdQrQ3iSp54jRUceia8YPNNNTT6YmwMLF4BHMsP7dTtvbgysocY
O3uYdO5I5sFo6yXIg4b5cSX3QfOzXdQ7D1eif1c3nr04T3fgazIoA/rkeju3UOHoTsAtm7sT1TlK
ELW0maddkluj4XsjwuXgIV+/l6eMDmIlhT4CzeSno85hUV9r4XMmO2e1GYrqiJgPP7Y9zh08sNNc
M0dt3ixuHjtoQwHERNzNUQ4whN8Opmdh4S4XCn/Yn4BxZQC1hdNQJ6XtLMIlJ9RgnRyyrtQJVCUb
QQJiX0mu5JO9v4Bzia8e6GHtN85wSMioLgw6K6wCLtFFExR134INglU2ldN5guBcNz9zrwzoKF17
9HgrSMCkSMFvyxVYbzLYFb1NQL5EA7/vBSvYZH+SDnodGcaWk+t6pKSJhSfpUyyTTdPT/TNrBZLI
fgwyibNXVBMM+wDqPe8pmLWjhh6DMWuqDZIEEOsu2CwNHW5NrlpVTEXo2Pp/rI0R0W+cdRCCqxkS
KwBAbrcG6ao2+vaVLd2Z9zT5vyZyoWSRimzwlbBiqS3x0CGXo3pewsNlK/vYcF6ScDoTOUQZi5gJ
mX3gIqKfbWzcaLIQoh/X/mu2LRUx+RIa7j72GCceeA8SmbB9dQMTlF3sKvAHrt3fwOP8mhKGkVd+
T/nhu231x5Dym80nQWDh0Klz5HjhKEl1b6wfoAYCTNbMuMIUv0IeI5uDQmzB9NnmV6GbIhFR3Yjz
EzfEfSQBFuAyE4qLylmVgjGF+xmbfSzok8h0nRHsAGO4HN5nFbYSnARh7Z381Vf01BsY7lI3Fr9R
P+2fqAvYstOpLuNR+Qes5F4AUvSkwVwRDleoOm9/+PNbngcuCXnfu+YEw7TMTAljIpz4sQ0764/N
4atVOiFogIcGVRBNv7SEmZBN33dWGUrhXZ6qHL+WO3HfViLsv06iniLKHBDxeprLcdbtMR0f1QFU
A+nL0fDd2+a3BxTWghGhnxLJHQo9YHlqO/BBwIF8YKo7qYx/P7rmxWTlzVJiYcUcqIHPkNPXLD5E
/EjT90YgjaAtEOCCITzUROinJzKAiH8hi6vssYA4bXw2NLSx1Y7k2+tszw/RGZybmiRGK5Ns4ToB
VU8FuospSZg334Zs/GJuA23734L6uYumJsU/QPEnk8JsgpFx31BDzqGo5Ly4UEqP4HgTULDT+wNP
iGZci9aGj+AkFC1gjyVfUDZ/kUEhJxGruMbAh/QBmMWydMC28MModJXXtSQNpPJDKIfwrzRn74IM
lHeBxXjTcuNeUJOBGUnTmwmmk2oKN9vje1bq1AOClmPeUeorpUvGK5kbT8sePGGmU2VtfV3C4r+W
QQYOsgav2Mtf6f2cS3dG1eWD05R9hxtyvDUIYXim5ld0T4AF7p2y+IrEX53Zp6tpZR+iWtjyQixS
dITFID3GKloUI0I6oTXWf48q3zsCcRCfPAIZVqSn5mBcATbPOrO3RVFgZzUDHMGKdUJV6PUGNT4V
rFeiuiuFX2IV4Ayf/jC/8PFAZmjjABZVVYmTHJf58t4eQ5vTRH9Na6V1lnbhxFsp90WUi2qac2xk
wzKz/Ejxotzkyy/cgqKaK0xMGJCQ9cYZMrknvlRWzxGgFbHzjRucCBTOKkwF+fcLCk5AivENTDil
yGyaPqwMRHMUOYtwu5ef4ZSs43/nPAvy7zAuW5AbVehRgAFbjaaSt/cNx74rBgof8ZIB0qVfuw2f
KFEkr9ymVEU+kQBRI85QAPXLvQj8pdltd+85PXODq9DoYcnrp3HZKafWXvOlL55N4NT3ik9lAPUh
pKB+EAdRljEZN18b84p6CDOgP0z1qEgjo/73a+LwajqVtCgM5yD5Bth8HMGZBANU9hEz6nJuukWi
HMDhYtULjce57waRwB3mKtISiggoCN76/hnniZ+uLE5YdqQdnkce687w5zgxs8VBvz61K8rWBrCP
/NgtOtNtGXs24z9DCeDaA2/j+blKmJVNK6UPSiOyuOtUStz/AZznxjmaxxK6jtsTAOyqEJUTOtXa
M6Gx9TQ9AZitgaakvR4w39aBiua1VKWJmhq2+t1DKxT+qCCEp5N3F2tz2H680q2K7du5T+fS/pQq
YL2P1jIeFNvn7T7aMFcA9Il+wFFJ79fQ78ZqT/UzduSnP0/6gksCZzSqnG49cdiNypj9FhmclVQD
fEv29QY4qr20zChKhW9vwRooqYsjrNLen8PUiSBEKDcw5te1sgS9CtvSirh4M/FER/S+Dok2w2Ni
FkwpvNcudKLTKdsb8NiSTFwDc3exDwh4OZco91OMkaUPwf09KvhUItBtBvZjSsXgSLnqqnjETn+7
lYWRVXL/+DG1UXNCPxSzld7ApZrv4AzALhxklOv2Ws7iNpPu+O+lag7DV1bueaTIpMN67jZPjx9O
kF17Vk7/IW2N0xHZYyqg+8X2ZUjUUEI1IRwby2pJYo0JH3hQAoDgy6CfUs89+7fZyMGE6R27MIJW
2n17fp+peWi+7ErEbwJcbF3hfE47pZARPKPboWWTvEq8Kk+1mzRfzaLuLeUuhxkBELhu6uiswbWz
AUYZD0QCt8BZlELRA86MGbgJwNToTRfnN7SAQYxdtml1HluQNUUeHP7voaEjN9MPy9aaUxAqIFVc
/RfaoMyZi8bRukldWr5Ad/KdTrbbHZwRvWyc08b2I3CECERP3oLKQpPFNgToPOWbQvMj+Af+ePp2
dUQhvspqdDJ8GklKq7IHqmMvh2CDc3ocZl9uwzJW25N5rhPosMguTgMyvmE1Nb1V485+DHGm7d7A
gWRbIXxSQZ96RlFTlCQ1lv6TF3lyG8TPfqAzA553Rw2IWJ3JUJpUBn8cFoyUFf6VP93JeTYENuFe
ebhAZgF0kjiPimQEO5BePoB7MS14fKUu3Y5OEgjaVAWmIfwR9JXRwGc1SB9SeEmYVYJlzXcXjgcw
OEEIPbLgJggvLUH+XRdhoBkH2Q+rmZ4XD01eueAc5w2j+K6ntDBzscNp8mCRiJwSg6iuSRvGLgrF
5NOuI3XtVzRndoHvKf25pDNTVjPNeoclZwEMgfkG2ECLsebxaGQoYo7u5CPJSMHPpPkkF0ySGsYn
m/+qgHYayQDqJuXvFvNNj2mrhCNUyR66h76JXDvIzZeZ97inOQiRyCBOEowb4Sgos2As+ap9vmJS
X7TmnT1P3E0BGQ/iWajCsii+YkMU8HRk2aw5vD9Szdg3qe8z7pkrh/C6lpPHW5T7RAwJJ/nWocG/
I7wRNxBmetfmMJFlV8PgsHmLtnSu40LQMCRq078yduaGt2b6ftc3mZyX+SPnq9gfLHfMj873lBQE
jOTO1HVyIyX6RDpGANQ07Hc6eOdz1bIgr4MCmIZAqqwTuvcpwd+pXhM+daoQmW0aVmGITfqMrq+e
1ZzLYnMncU4JGq358xqWdc8Q8SxVQmwhhoe4oaeLdCvSL443hCxIpTHmyR4qqfuaiB9fikpHGdiO
4t7E7/HBsZfPKIeIEk+UTG5kBTHJ9JomH1SkafY1WVQW1ldlKt8P0e2Af6+lwKKGYdzIGovmIut/
zvWwm0ULJwQ4UwUJ8mF1uFI1tdhW7FDZw46Af82nD9G4dck/b79GtCgMOs9BzGPiD2fMB5F26lCx
rdeXZy5+Nr7taMF9sIvDRptoo8QhRA7UJy0xrT6G4zyc5YUd3+qTgB4TZLD0qn93pg6aGEUPJNjf
8YQGZ61GvpeAIJoxGGs6WHzsxSyHXbLNDSxWRwjL8JYaJZI+J0rl6k/IlauHMCeyTUKMhCrSlwVz
mf1sjogHqP2/aGTB5aG1wqDoOKrmIRAg4Njo7298tY2NRcqu/u9XR+mqE2f4n1Fzb7w3dSgGrbYA
hqVtlyxrRZZVwQTRuApM2YKiUpogzQLNAVlT9CGJlu91DqOjgWAAl7Sc9DgWNb5FDNioyeae2/V0
IT4ZeOxyQUOc/hbJ3CeZFhLc2d9McFNLx5p+uNETSr9Tpj/dA65TVOaFSbuQk7R3WlpjGXdMq7bc
2pMSsYil+XcBTQd1FlOiEbFdm1U/Qxzzo6u30sBz5BS1dkIrnb6nBc4nNVybGvWz4PoHtlQyfC4h
ezfB4ULT2o6toRfxZAOPcvaWmSSC6MVG1JIwVbPzdrICLa4N6OL5qcPnkVwgDgPljOIEP2CKXEeO
uu4pHcYknH0KgR4j66AcvKACDo4ShBY5KUJ+i+j0g52fcuD92qzjQswkecZmLOhfkBGAEfKf+0fM
+UhOj3ul6ePur+cCIwhIiVRFlLfU8ZIc/thgpkSYUCnGBUm6jRuKGa0eFcX2JPSf9mmlfR48ftKS
/DCsRyPmsSydXeEu6xm/7QUDqWESmO8bD8b/RTCvJOJAc5UuCXKxOuzcRGBbzYDf9mRHBnkH7o30
mUsZrZ0BBmwrF2A4CCMGkoX4dStye79HOx0rg4uRv7SwEOAohMpsAGU0eBxfEUeHSyd5BKUozvuT
fN5u7mD1g03Fp5vsfGJFRg44I3A8DoIiFm5kBSMCx/f6md/XizjgeBHMt0qr9eTujiHbGUtgGNGD
k8Wh2FcKYfDUmUBsUUiSNj9Y6qJqjs1+rD1a7lPeQXTPyqQ7dU2w9pnp29OetbBEcDhjeCGXrXkz
CNW5s/QULmt/VKCiOrUYdiRL5mKJ2ecWDqfJk/tCiev1f9AfBQLUFgcPz62p9i3CN6SnD88JKcHi
QnARd4mt/5bM6avA/nRv0j7YbjI1/Ja11YRWZPQeKYpS5pZz27xeq3KKniCTpm5gTXPZZGr/BWyu
395OpnA498RpEm/veQxLazRdO5VjyoBzfdLWA9dwa2JWw8vs/BVbbUQHRXaPB/ZD0ZFu2J5wiz4I
SxY7uejlvjCwvx59xKjKm9BG/oI2H7INdeYqfFs65r1iakHymYRBvIzBdrhsk8RFGasvg4LGbsn0
RHvPaZ1LayDQmRDHALT77m4FenOojZuEgFrh31xikTyz5wBCZXrZK/Tsa7ydtwjpw83iLt0hLMwJ
B2HDhucbiX1wEvZeu45m62Ybq2O7yxHvwkugiSvRz0MqNgtai3fK86XFd3HQEiJRc/1BVhVMz2qD
KmD17Ika4QJLcNO42d6nyEranMmuIBg2KIIHAUgZTjqaLub8t9GU/T580wOwJmHtu/64fjTraQo8
4T+6YdRy+aPVWoTrUOlploPHXOCHV7AtMvn+9obT9a6nc9r4KaNbMhD770FV50VSc6fTSVM3Qe0P
dNlJGIutwrQHDwq9SuUROb5/3JGLBKmQDK9HDbTrdHYhsKgomtjeAh2UnBVJq1juTOyD4R5sEP0v
1Xend0RrllaM+avEUsXh/geAqossF+AnIjY0f6NitrR95tA5puAi98kVm0N05S9WCNcvaDAVRhfH
RlB+x9HY9ylKeO5QdI+QxWYXxklpIBbEa+rd23qMAgsdbSAw7Twysc7390Ulpxfoa6+eTqy1zeKb
AHU9LW37hIwxTNV0qEz9BPuc7VG1oIuaK2axxV/EGQjehLLCkw8tPEyX4+VL7Ssciwh/zSIWa4cI
kpqvqNy0IECSERq8DCE5OPm7Dy3+KBU805xy3RFySfgPqPGAbHTEPktT6lCfYRmdADYIpy3s1cNO
wlOof8cLPZA7raBJWmFICVPa0XI+yjDW4N9lk8xclj1dQq99unEPUPBU3aNJrfCIU785wj996/JX
Z7ta0xTcKoSx6brGOeMuRb3tnTDXMZfitch9ALepcaAxrPdw02jQaSLMAapyGly7Q6Jvh3F5ml/s
d5wqMl1Vv1aptFEfir8FtMrSPega0e4XocvJtxLG/6Sx3108ShmZFHx/bnyh5QTXpFp39aIbWjva
pT5yal04ZL2Af56bdXmD6DC9ttGicyefv1irK1Uvyttlc4Eh+OFpzvL0PUMWbmnYCpo5qqRwN/tf
qO+i1i3u3s5ckVlqPgezZ3tBUM81tnrloUlWYd2mITSKDv9OlDwChDgUZjqlnzpVuD8tJgsofKhx
Z3wv/dcuCBKi4CgJNoePpDUn+Ox0fEF0XfE3FOajQvaOLG/jkZIJ/K/pVcrBf86vcHOQT5l/9jSL
XHGDZVMVln860pd5zNYPF8kzp9h5AD/UJVezk6SM4u7HYMaUUqWwidTh3SKzBeRYvrrblILyy58n
szSJLvONQEeS5+i1xzyakyYhPbgvakAMJv7K7+8C42RAL1lnmFBHAjSLoPgBZwxgHrCia/DK8RgE
2dbr3TSkd7g4rDjHBOeVUrueKOQ3ipK0GTYQBukTM7WpjT3aaSWwLwSICm5928mESFiiN5NEzwpz
fc61EsY39J7PdpjQ2FD332b/ZbYmBJJ5Nd0uPpswS8yok8TsQVd/PcKFTv5A17f11519Vm8yJxdU
BvKfRM6AAQanG9DoKaCaRP09Xz5sZpPZYb/K1Vox9qD11+cUv053nPTUXaRrO0ahuYNDlXjsc6jT
suHELv18h0TXUWqZbn4Shgdwd8rcPpYanqsKfNynRjV0qT/hvSk5kKD7wXR17yUPkZBHwrq59WI3
ymyeb7hzGnaql+hK3dyNyXMjEhm2PtJrmunWRdlsdPqXOhotmF80nz38WLhzxhmnY9wiWTfUWGUi
eiyMhngFFqLhYlWShI6EBRq1cOnKBjjE7S8oNxkZNUR/FoqWe1A0p3EK8sQTBK5vmN1PxzLmt83f
Drt+nGCohhRokGL3deosqVe+7AVdpzs/dmSp/S540vdeEeu1DSucbRE4zVI5HTYA0TVrrJHWwmvJ
ZI4gWTOpj25lJnxEgyNob0sw+/0GmyrkEKTiuxzZxXJj8UGSyhNGfGrJ9/VCZUeKwyehCQiY2LRq
J8/fTe7SnM4lPGFqOV+cbN/l7z2N0pouTQHk5KdKIiYx8MVExBfBDjF5gCGt6EsP7qycyoly2DI8
q6K85oryYapA6RGfX3gTOfPhBf2pxfx9Hk85fiw7SmEKqMMFofPkJ7VqvrnMu4p2AcWmM6WYGxFN
kIH7czicD/IhzACPylTxiJdRxwyWFekyrlyfsNjBUndsjpcDOaqSMRf6geGnrYfOzG386Dtr+ZpN
jgn6rQlr3TTNw68OLukLov85p1rt2rm/lDtyGqQxNSUlJ70PX4PWzW4d0ZT3u6BtuXLdgD0CYV/m
6XjbORdRnAaCjiKovZq8g+cNv+TLHAqYi3i/FeC68BpmWWfji4owAcHOYnsbyb8yGC/Ki9voYfYI
eY1kMOk4nlLLc4EfxarNzRNMWCpvvvnaOoj9xVGZWAdaYM9neHJntCeerf1JE6Qw8B+a9bu96ndP
AfszIOvWv6JHaNf4pnvarp+YvHrOuNPWVGmwJwsrBy36joiMf2Tv+fUuA7rDAVLk6AUQKREH7LCD
MMDZkIJgAeoKBL+zye+9v+1mpQ7S1Z2RbihDTaY2ndvlKb5N1pszTm+FjkZexZDNr/q1YUQhp5mk
zlLWzNWHGUOVB6o5rJ2Ma24VcWeB8u6wJ4SZN008SuHI4DOmRz8N6jkVOg9U9whESVoQF7EXVIxd
7VGGERKPNZyQvfm+FAeyrWKoh72oaxlKH7cZmslB0qvuwd8VvdvBfehxmL3pMbZHdF3JRpOWsscz
7cBkSS7bqoRzFaERtxKtYLCsDGADyZAzkGoxzh5w65KroL4vmoi1CI60d7BWg76GqkPYM0YDLnOB
ffK3nZbHt7cOTVYK0vdt8LrVLufQ1ozQCXdQjEcw8YEvoay9vjuvlOrCRy2Vw8ZSMJdFfdPBaP69
HdPWdrTvzNYCsiSSLlj1p1gI3ENokE/5mFjOvt/vvaPS1PssgxFvlnkxtpEofDsyFT8uhcR43Plt
22tet/uYkkv2e6TCQn1vyA9bvcHgKsgwwt/czu59yxy9vovS9wu2pmLyJDA0amyDQIHiNz02cJK3
FqJ1dGG54csxUQ0m3AKWwGBWRXNJUFJWUpcpg5kgDMNYV6OmwwyMYa0MPYQxejU9wqtjxezmvO7O
Fn6hHhRFV33tRwBO8cQ/GXCuxZm1opfHzr6hD0mSBBqiMWFa/XQyCdue5d+JZ+1x19eiU4zeC0RL
4363FF4wcNm5mpXMKxRKzwjtjpQHjuXS864JFqgpf3Z3XNcQLnHauPpg6jgH2VFv7QJ3jkFNptIm
Wi4NRqKfgKmzmJuLBKDBYX7UtrSxCh4WAxBPwKw72mWnqK7a8GmsYGjVglXJ10xlikP2x2NbjdCY
7nKXvsV//750XrIrrYVSCNnhfri3G5NvXSX+uz+DJglh1P1EUNPGxPg0wHmG7JIb8t8QATd1s2/e
ae4Vf72DYdk7yJ8jOdKyl6lMPS5kGHSl6P7upd2DkOSsMPQsh8iMyaykFllub12p9Cj4ehAUBlu/
zo96jMj+6ulcRccWchpw9LBV1dWL+EC6vyq73aV1oz4xp7+os6Vga8IKSKaY2v9ti6ymj1AaQ14U
40HE+tkfcqloJgWzryfg7mPtxuQLLwb3FlfunPWPsreFP3VFeKN/oYAZFMUWKvrKgcs4VPKnL3+d
SRafWVz57OdIT2tGyfYpL2bhHcjaAxejZfs8UbUfX5mZp8kWfTgsDuUANcOQnQJLhVIkEjaNy3jW
iIxaDwMhVfQxAcYs3DUHTNInHm8yapOhMBx3/5CAzsf4kiNFIYJ2zER3Tkh2yrybvHvcWU+SRtLD
lvckdfx0YPQqX602ia59T024fJegedmNI8yNpP6/naeRsSEhzd2MVnv7idL7gvdvv8UywpeEn/yY
+suOq6Ii9w4+Mr1JxOUbjcB+FWtFjctZ+kmT4m7vCXc/+mhlPVs07yDWWeVsxYXT498W7BdrrqMs
GMCF2XR7EqCRa+wDbkMUlsPiglBNXI11W2Yv5xydS0ele8tVuO9tFPkbJmMFkYKApfrsgJGECD4c
5m+B+FYw4dKSSuGg1Fppj/398lh81omjDcxgNCS0ZS8y8BOz5NIpP+867yPOd4QfwCzh7se7JdcH
AVQ3oGUQFX3/zZON2uILpQWtGRDolw3Qs3UXeFk0oGQLjQtm0i8DUFuh76+rii93a/RB6RumP2K9
V5Bt5VDoslRyEKbcCs5KNtnBEwd/HngEXqQdAoA6uInqxiDeuFKuqo6r1rRc/eit0Niypbj5U+ux
2DPqNA8SeCRej0nSHn4MT14apHJQn/F1AlNVtAiR4R8mBgVSh2z9uudyYvOFYmaToc61UaXk/obZ
jgYVen4F4hoXsQmaDcowh/fCKl+C3WoZk9iCwXYXZ/IhgEhpJT3pqyTwMan12Y56OmhLG4w/aFBX
9vtHcfgaHxUIqEX8D044dg9d7EURXya9xwINbWT6r91UNSJQFwJDs7NJGc3XwmAN+/chwlbyuhV0
+D8hazjZLzj0j5l/NFTv9VWdgJhvQg7PqnH24djCFWXaan48T2443rcr2nkvQRYwk4d8tfrvrvd/
8tBU+6Vf42PF1dYZ9mVol0+8mPP5Px63ij7/whv7mn9wLB6JKI1AMm38yk7jnGupnh7673KEJ8Kz
9r2TuUvSXaOhaSm53EWh2b7YA7OQKHLaXKKYfo/eLHcSq6GgxthTdaZVAR16e2BFXC9mZnZJ0RXU
5JcjrKm8ObUrtBR4D9u6d91mYidGSzxf6P8EcwZ+9sedUoteDb+87jHyvBe+6+v9uHdOso3nRyia
nijxnXdf1v8wHSkBNrGkE7GyYtuZE4s3snT//+//NgT0Cq+OEoVhQxPReIkjqloM1Lxlw9OjRJ7Z
3tsKCeWmQogvb3pxedFvJY3sHu2x9qvYsji1k2PNf9+0NJpoxGN5cMuW0TxqEXZXIJ5zaD5zFkqn
d4J1X6Fd+0cOhXVWX2nyT5kHqyL/hhsZenAYlUUlqvlvAuMnuC46Fk8GXk92mZx33MdwMEVsYa41
6YUgxK2cs0eOFlT7jELQDLUEjNlTP6LVjTibm5hlkxfsJcCMQVUgAE2wSMAzI5Dscy/Ty7c45Kgf
XhLdS4PFgaSHlWtbDmz3OaJC3hqFQv6c7ZtoBJx7EGjymm+yhKj8vOUs0KAeO7gZ3Fs189PkEc1k
TOmd76Xy41wSvkxIrQrTCShsSitiuE/i7XaJBtBao5BYCUanKWx/PsT3STIg0hagjKG+vYameAG+
JcX/eAqO95SSJHkSfq5DKFHYFEV5XC35P4wAsF9mL6iDIB0TpWOW0mBzMT+d/uv5kI4alJBQfSZw
vaGtcl+WwNa2Ycq/hhUOSvvEyudgpjQt3I0oMtJwb1GOFg4Sgwy2/wgNKHpJQF4QJFmyf0lEBvV1
wwrdkM7ITXWO75S5qN4OBG9SjlBr4jBForR+sxmcRWjIwY8K1oyfCrzO89w1mScoPBSsZAhJ4Z63
Jevo/hhudwrfAFtELA3+M4nRcZUe8APWrC+5nGtXFAnuP7N2Ev8oYFADQl5w2siyCSVAAYKcewLx
ZEPjBVP1vNKSSg0gCjI7iIn6aBBBZY/oD6207kTw2muwdCDQkXwdEZPTGoVpbdxCBXSXOfiW8NAi
pLXhEKt6zBEs+uKEU4lokD15flO8i6pEk9MEj5MAGs/YWIzhHrcJIt8bb0wF65M1zJsr5orOHI0D
63OeHqnqqWzZhUzcN+RckDgSRXCsiYn5wO9OD2NTK4T3eByrjfbi5krJ0YH9Tb7QwXT3evPF5OV7
vrcmJhLaa9IhR8+CSnff9LamEGk6DXbmsEo7Aztrxue7spf1FPSWdMhcmO8lgzrHKjhoKSkgl4tX
vfdCZu06CnGWJ7FQ5rlvq0A9vsPb/A4RVTUJNBaUYN5fV2WOB4bhfHmhFYwC1GoHGoe8fgTIDN2R
ifdOMzzzrRHvWTZxt2Z0jAkdzXnvNQIQGIgAWBX5ms7yb8HTdxGpooocO1jUAw2upmpYtFQQBQ/8
7SMaGeX59Y0IyZ4ReQgNTr6Ea97hmzqMsm2PqZ10hdhYEFk3pzbXUNk6C+eEdmSlbaC+gtev3K3c
mwizR13kEH3/xkFCLR2vuzfegKbuZIoWcqk264Rz1jXU+slSUj9mi8u/B4O3v7On8NChGG+XV3gm
HfzP6SYDLu+QGRDLTgRLSmBmXJGV2LjGyKpdXo7oh5uEb4gpdJYiisoaPuNuBt9VkEmKk4/HnZ7D
trgXdFc+Kr3nP1wrVkMIEnxw3s2J5UTUicKI2N8urbs1dBYfBh7ZjX20fFcY8EB5Yhh5RCJKdHec
8DlgmUTTVBd5km03RIinhgURYGLXRKE4VyBqdp7jjyiyN25wNHEYw2I2EINqksf9LZ0oJLdYZP08
EmPzgzZFTFF2l5ogEUOAlbzNh4uOYi0YjMvRXAC7JOoGYMaqYU8vHd+nE19RlUa/Gnme7EMZMeb3
3UFuVPs2SaUijV/ABm82J/4ogcT+EClmNLRTBKmV82bDNZ/8+vHSX1eNmI/Zz7gHMfsET9+o34+P
gMfGhsMXSCIDzXPQsnFWPAH8Cl+ebXG3mDc7qaM11p0rcuDojzWQO1WNIKSnUKUOhtOqk8Ck2Dow
aHk/uxvZFeqAHN/BN2O8H6tcJT4bO21CH4AIMQJBAeUHHkFxduYMWFoGucX/n5i0CvouRxiyKcV5
qTuHD5FOyw5pN+yreBQf6KqjELVd/xBoRYqYFfJifVaFhGDTucbnA4zIlynxgw5n/RpOgDQDsCog
MP2aIxjriXQthyXw9w1elVIxCllbLCt6+v/El+4+tFKBiBVSq64q/5dv1yBorCifBeoRGMJvra+W
iWexdSGVsY8tf0/Z7TSH9SlznDeOt1O79klFrV9ZQ9l0BLT+kQgjHTI5jpIRw0ZnjY5rSLTG2fux
wXP5tBOiFZk14ocubleEny2STtLPVSLtbUregs5ziB1U4vZIOIqNDdUMYtgpS7E2HuR90MSZSDdW
Ht+ThGyp4g4R9Xa9Wx+Lc2UkQGA7DIsT6KjqvhtMtciZ6tAxIJH3IGYos7c/K2Tv9FDTcvnmwGjk
OpoKnv1EY/W1kDk6dbt2FGor/1YVaDcrtnu/4QTU5/vV86V2qbzXp5/8lk1T3WmP1K3jQi4rlt/N
zqd3eiw1AL6YNVzzo2LaoQuJC8eWyZJvKWjusXlkNGENvO0hoadSorrG0h8IV6i6c2hMS1yPdlSX
EGs67fTQGV69S8hK/zSrTLRoC6D1Zcr8jhENzPQU6pOj3E4ZUiodWNJHHhWjKPsSixxrEliVt5fl
hO4fbp8R1+O1z+1Tk9lDC3RC1tRnPE/gITpeZurnK7+G1WrWWNYGMDRLGMGQ9MbfaVS90iYsn1e1
otts4BNVuO5CzEhAcy9Yg6IrOdII82NExscQqBeg8IIxkIiFuljU+7TBKM9G+8g3GQZK2LQ3ODNF
EU4b1VkV+RD1E9A7fLZj0xD6ftrpo0JArRyTBNuJI7a5gwI5mkPNEE8d36ebfTjkSRl7MdueucdG
dSHNFwP4EC+7kjjJ/AWgPFU4zIfRiZZt5HTrHfgSFQnifIEeRIm32LFR5/dvobpM2/ewMLrvKrAg
cp/jmvUoBKEy3cNUAxbSw+mEuD8pD3SqPkw+S9KMbswGufRz9wdtzbYz/eqFcJB96MnEX/vCFJCn
YLpGFzSD2S2s9eoVYcL1sWykGXd3QmzK8BFCzU6vP1OBtUUFaanjUGiVS2LPeV7zIv1frDCsiKHi
ctzE+6yifVZ+03Z8v5P9oCBC0dftIMsRyQM1VE3Sjy9dWBWcO+oFqgxS7di7GP93YmnlvOCmUR/1
5yJZT11eSAQenL+doXZf5mwtyqS3ORsMajNHBhAn4P70x2GzVljFp03v8xFOB0hMyPpK4CAfUh08
M8UUBP2tM/P7eiUdFnFYbmPpDiH6j7tzbYdyCH0leOsSO/3OlH6rnv53e1p4pHog+qCb378KU4OZ
d4LCqKa6lMbT3Lleu1OOUm9yCuVOULt00Z5jVQZ7/EWr72UMtZyvUQgY4Va44bllOcnC0CnEHl0z
pbvpluD/cWkOKe6fkT4D85RR+GEE2AwdnR7gZA68wmY7iT9TZ8/DGzluzN1Vy1jWEpkGhVF3g/uu
Yh39xph0NW0EPghTu3snTKdiitDYXAqObgirfSAqtELt7AHt9KO6gGZUYaSjz0IOBlsBvvsm2dKv
/7MUXT4QMrj4pijNnxpHdFISUI+HUL91eSPMmH5qBushAG/YwxURStwZi8nsKXvA57V4J8/3yxY1
IEiQb1Xr1+Q8Wl6LvkN6TVkyP5lIPD7B5CGsNASjbg9T9T11hCA8I7gImQswhD6T3lDBK0UxnmzM
3qq9KPdlCjsfD7x4OPXq7+38cDfqr8UCWuWh8QHTEcfCr/48t7aGzk7KKIafmhBGKTmavD9dx6Bk
1cr3JASOwh1psUKPN0bGTu7dTE9zNIFknkd8ZUN6OF0GLEfTxFW6GNrhMLwjfOC7E4oTmZBww7lm
fv1jyOKC9rwAuUVMSSWThC2RT/cP0hec6nYFAM9Y334t/1+rDiwau+cSX7x5qWcEX8TyMuQESV+G
L6TiYE1+6PuV3M/8fuFVYakRhnifzZWZdX8vh0kOymXaXyiQthN/kOAXjV5oXcQJDKOhC2zxomeg
xuocCUcIdnJiloa3ARD/ylr/nSB9yPCCZPx9SYPlv+561nyUm5gtGhrE9Zj+bf1V85PJIPYP9Dgr
/Lwds+qfbva4pkDw0y/Ky3z1rUfwsAQbRdgoQ83xMcuwTUObHYhiGRQuDThr56VOZHFpN5hVLJL5
/PseILtCHgkOjZ5HZ5pKGVfZaC05Nl3u5jvpH7foN8/KSWq9Uw7qg+Ux6zMWaR20qgXid2HrfXVk
nbPPfQ+VkUuO5TFSomPgzYt0gzpWpQDttSsTjRmv1W4cIY96mTGmEVi8N06BNHSTToSl27SqDUbk
I/OKBKxP43isDUD3QN5ctpKUVnkd5uCEHwsW0tuFnPQNUzZOpMCX4YR8Conjwfv8PDzBJZmwm6b1
d5wQmqFplKsr63ES73rbUm+Di59jq9bmm7Dk1f8JAtYebNGjtWOmtHZp51KCCJeaLQaPJRrSOY4X
DKyE3nCCIePW8CT/2aK12LGhG6HUI2Cmgt7vMtmAdeRILIOgzHUs/es2PAUkAz7QoZ5QIyE5X5HO
40xbvuiW6vkuekWihGd1KXLnNVav5ws0wvuhR5/AMadCQV+uxs467Y6YvAXNdQdiMqfZbRVnX5S7
syQxHG+hciyczgPKDvcpL8DFvcz0r+JhZlWHQXodovMBZfJKSoIqXyUVsu74lxHOWE2G5FRkG/PM
ptjZVy0Vyr4TZrf1imB6Ml5QraLtBq4e7F51Bqrn68hW+oZE39Rh/GoSCVrbB1IThML1oauUk/tA
Z2zflaybX+9kvXGxKLz9dFw3t7fsxk87AfJS1yl0JXOjXc7ZoIVK8ctfWB9m8Ioc+VQqwCm2Rea9
EAOAHy4DOtmsSxA72GfqFZCDQ7bEx0W/wOL/zNr8DqSe/McKIsoVecnANWE7rVYhggvA6c2mTpKm
DA4T9II9E7j/GaL0n0yhFtW0FfZ6X+sxrCWsD345E5G3++V59yzm/8RQ8kZ64AWNafRRs9vbAFzV
e4w9Sa95S5wxfa83vaOntJ+EZLjSgj8JX9pSpuAEuFfUe44mG1tWZe71m21eIQNWJ56G8a4YCXQ/
oJmoyGkG0knK+b0yx3Y1B2G8gqw9MjfFUwBYY+E8mx3mGTHNlLYYIrI03k8i0ELe8Kvb3EgJs2g+
TKQ5uu3xdAwbfV7w25/24kJeXOWw094DnBf4ymyJayr5KEdgng4XGDEeOBZdBj+XfYBEkR+xDspg
E8gHpn04sVISsBhJfNf5MQPQO9/S12/VQjI3zxxRJxZJSkbPMeYXb0EEac0yECAtGZj8mWTGERA8
YnjPRJcCbCXYpyK4srcIAyKOWxUzXTx5Beg+g8e0ikP3rB7BamzsfizS5zaUvkS3c98qZ5yMVAZw
meUpWHuKsyV8znl9jWppMAYCA1W9N3oQnTfROHHe8buYVDvIZLbe9UE33jG4Sx+RafNVUnGA4tjp
HChbA0b8XTCQeRyeyj6BXZOYbUvulVwfUpDmvtGwP8PKWE5IaCC/ElKsIHiZVh+/BQ9xj8kUn9ah
dAcFmb4dixHF6Lusys3G6acRQEMfOdUJNSF3gbekWR90BroLh6mGC8Fh9oKCaXJXv8sQlBTnRYa8
HrtXPhFQ0opo34wJuEZXTa91t5gBc43n4ydRZdfw3RXp5ea4pUQaEfv6OG7SL/KyT435rYkoJMbb
ytvv6ZeKwjJguJcUQ17mEN/ATBygF/2hDlZhxtp6k48bz6CbMIII8kXDnayjeVue/VkN+OHwV2AS
/ZDCBkv5hVKUCHfId9yH5NgUvkHjQnVv1hdJQzp8r8Av7xsFciry46pShDErlWb73zUR8JCkxJx5
6S5uehzO7GKeOxzsudKCWgrxtzXmt6/denlM7JDz3UrByUeneWCMt2yiiFPobzklaE8TK8z5PuIQ
a69cyXrK4stMJwV3RulDs4ttX4g7hGUZIh7FUxt2wXiCYrYSDY0Pv7n9UETbL/3KIlmGgI3QJSuj
xJ1G2sbvBW3eCSlUabFVyMli7fuRReHMDnT4Kd/v6RWfmAUzNh6x/9IsLaOmwK+GkvbMOA4PNkKa
ATBexZOx4PEWbW619Ri2v1cZAsBIDRiNo7Pi7mt9sZlWO5ifF+PfGNcMdt6LljmpV7mx33DC5mVU
eXg0XI8jVdM6pMs3uz31iXWeeM1/qVySEgpVWL21gGXCyzAWAbVXkrF+qTK+cPqp8k/ZtiRu53nS
fHhXVTLy4DDr8bZcF1Mf/Lm4aEib0TP7QdSd/s0qxoEhKmd9rtcTwNmVA9Us/xyRAGkAr/mTtDUF
eHTAzJ3dZEZz4Vp68AAGL2cmdCnOBkQozP+8qTUh7En7qPOVirytIWCGT9fy6GVWpcj9p2g8haWg
uXl549qL9hOcYQaKU3vNi6q847sar4wNl7iafdCixSlZrQeue25zQSx1PaJpTUykeDUt38TSooUw
owOBb1JmoxOYFAdvngyH7c/01AOM/IW2gt7xZc4LDrjMXRGU5BGpJdETUoVukU12zTG4qSegmb8I
ZPBu07ZRIi/vPwsE0SrIPjqJyzViD/n/YTOL2jTC6S6TiFTh9hhjM55/bv/Hdw+M/k+nGvk679rl
3P+426M448whAJ2Y4GZyD9QDR9O9N/jm1wbcSF8iiw6G02eo8HRsSDNMprkhej5KfUIhRVH22LE0
PsZRlhevI7AO0oGyD+YAHB4HRS803RhF5igO2aKgHkHcHhABMtcX2F5cpfabhn/k5UTU2LxJhbRd
t4BZNGTd9LjDnkLJY42LWsi6k6+PVtYpve75F1nwoXJiXWOtjmYDCE0y+rL1oX5qKyDXQPE+C3t1
o8mXQ24tR7MUncqSCPorYhAnBkHmZhyZ4ecFtXqXP320hxCSdOBA42BoqrLZtlZVXJzH7HGxvXaf
fFYW+48I99up0HIMmLe0TWu2otgmhW13CNST/wdDsp314ztu0BTVU0cKhFhgsceCHNe1MMhHs0XM
ae/KsBoOb6jmAGqNz1nO6+slWL+/880jPypOOwkp0koIMd46iwjBZxxUiXTvphTEg09wCncV8vt5
LePO79s1JRACxUgDXA4LToobuPphKtK6z2vZTUWNAcjb3ITfXlqDuaQDXUlc/ZUFO1jjNjZZd/Jk
9zqmb9USKzBZz3MjSOwsK1S63eca/AS1AOgqCde49uZPjtVsyPgK3zsveHtRuCrJ1vjt4mIxmIWw
9dFoanBUyxNN9BOEJVszmB+/ME70U/J3rvlvOEwht1vk19zFC+VCE307WuTWp05MkfSFPSthmMae
xOoVWBcy/8eM56Gf67rc++DlHu7qpprCbGiwTge9yXVapsDi+puOBaGyE29yW6SGMvrNdVpDzeih
xMEWlVHRu9tknq7bgkd4f2jYfGlvne2eusYyhADfTdd0p0lwdtiNTpnKkWeSxjxNneJvUOg2Ce9E
rQmzZCAUbuzcR5ZAG67jflhREIJ2YDrE7BuPsENAwev9tA/qe1fwHNxpyPLyNglPsCI4penSV1Om
iOfj8qQfijhDKI6d+hFhYnSVYTuK5nZ5zrL+DHY0G61+sbvYUR86eMD9JkusZG1F60ezQDmYfkSq
zb9PHtYOp+OWMIAJccUjzFuTWueKehW6TooBar7HbRJ33vQIOsQbnC2U8qd1O5BB6QMUEbPWIMbb
8ssSNy8WFx40mJVj8Wp4McBeK71/eSl2xn6fkaAY8LMJ9Pt3FEB5PN8GOv7DwJNmdltLWkd8x2x8
V+VbBsjuTAxinWvhCkxrCpi9LmsS+h3dEu7yUiBgQ4A4h/1PEKa8tHzxZ1XSjthGXPubfXjCi2We
OeF2btSA7GZkIjoD0sBYTo2C9WJByZltZtsmD6f8k09I0TTLeV96UMt4yrG269aUZLaovRGLqsK2
mUv7Ob8HsS2GgkIj0EoRlMdi61WQWjGFWCb7V5M2wj/2tZ1hkQ5+kJ03HO8aI8Gc/i58HLrL29GY
AhaYDnuddv769fVwt9DC3IznGvQRcXEMBpCl+zcnQHaagg03CT6vg1ZvS1Cy49LYIkmigLx8EXue
s/mwBGjR8IQx/Vx1SLnWlkbyRHDDxpluAyhOa7+lTkoY/mRMNvae3shOV1kUyR6esgtU9NEhk82R
oXYQcz69WrIDVAt18/QBZvaquVDJLAtWvhug5qMW7X7+ly7w4zyQD+dH94tSOVGYh0Pt/gvmXC2M
0VEflA2s19ho0SIhim2bnnOsFyYwfc735HnHg9UqjKccYxD1qp+XRIU1zH3UsYGYulV4T3JFXkiP
wMLlXdM1usPDv3fmpejHSpbF0Wi5DDp+tG2CZk+DH4aNjXJhtrbCPqJZHZoN0xatzLGmvhJyom/L
qB/XzUQ70Sg+bVjSKKDCd6JYu6yMLhONjAhyaHIZri0iYhTUdz0QZvXAqSsU0fFPXrI+56Y0/5qH
31cbz9DQCbIU1HG92OiKL1x3LtBo3ORm/suTRIu1GBopqSJtQbK84iKbw2OAqtdnyzqv7ZNDcUhz
fKCkJTV15jijshdp+lr73GhmL3N8O1F5gZuzCQw85jEMWrMwsCFf3lfo+8QKxgzp3pxw/hKQ5UT1
SRcw/wvBLTGXIJIIpbT9uUEYLKtOPJl7N0ARoVotaq6S/Fnta/ENzXXn7qBFcUIwWkMKWCLTI1Ah
cirSYrTlb4OhInbDk38MkLtFnxNQKZs/9oYja1bvAfnaK09BDPVwEbSnDM3XrG7tVhSjpxb9biXX
ihkCveI4KwkIBngFcn24uVKQlVtHDRUWqBh1J5Ws4daZL9XQLZCd5g68C4rUsU0GSb9K2HeyNL4l
mPjlMadpPpgcwSbNqm+w1qhnUly6xbnCkuPp9RUD+h83m18VvfwhqugqPXzWIgBAD/p3enLMz8ou
JXLEplxgW7sn+zEAo3Jjh5ZNdPweT/dth7497UE0Er8pXJMkuMKxZ9dutHyjHJ5Kn3GobwPhhHFT
FKEVkNhBUW3DG06K5/pAtvkJUNsnit9NDpF0+a8crfmetkO2OkBLQrnB8R8recA/l3ziyrtk1l4Y
GWB3cb37pA2PzyW2oFE5xIg1ewBtp5U0BlaptfRFRTnGhuZVthayEDHmKAP0XHJynKSCx6DMiUXR
gq+H3A7o9WtOe0vNsr1Xkah5yzZgLk4MKs45qAS1XiFCKvNZQ2pytlL9jDevsmnGlZlv+oWW8mZI
kNGVcMJVrXOCdYqp//je9BOmRexbFnR6vX+4bf9Ou0m0twTHpAOE/rV4J0JHQo9lN1IBjX2o+JQA
kSj7rzqy5e0gSxg/Y7KJQgu1Ps0FxTSy/I4PY9UK1uhTSGGmEC+Sg5Vwp4nuEyLyJ3xcVf39+ONQ
Y+GCKP/DzN3gzpmp5xBPa3fEgCzEUofgFv4mo9Oqxw5698lO0bnWYDipGLfFMQI6FfCIdeY8w6yO
8bYW47mCfJXyFeNJKkALS+r+pMb+imtz//2Pw3gZh9fEmOs4ne4upk0cIzvq7FvprQ3O5d37RFDs
Sywwtzoz+E4ByaAtxXDywLzVg6Dh3jmT2qbDe4qUUumKQRb4JJhYgqZi26X1gl+aN9SGQCEe5DZY
3Z8jb/XjOIpkkMNVJhwuh1yTJp8JSzo5LmnT0fzqsCcileoUSNcu8wJUismLIeZrKAhmTrVZlW36
XrtimQQvKoydXc+szxDkggOPiqd0LoIl9+wDfeukVT8XebvKf9SB+L1Bcm6pk4RiEYIFoQW7O2Qy
SiXxo2uoMy9TLOxr/QEI1vIALROD7lXBYPNNALQmlJffD5rROFDkT2qZghnJs5w6vkyK2zubRVRR
+EQb4GBhfTCGJ9havjdpPHtTKn7u5axvYqqPbE56hASrVZTPA9aexg6HWy83FGnyqiPBkRQIJ8qQ
d8Q3tixnohjTJOtI6QhPsOrI3oPxrM6xirknuNdYJjuel41E9bGPf7HK63nZaPKFJLREUbzi34tw
wXEBzW5BXiW7g0IgAly/FAO4MuFwdDKsWBJOn1dB0gHVFTWvGjNKDoCkRyX0COD1ogBwwsdlLB2Q
uIjiuru1IAEqSQqvPudIar0tSwm+kiFAog1TwuyGoImjKRFiaMhTAOMoBImdBtsdtc47lV1KVv+c
QvNKaqY1wmnKFrwxb+xEZ1KVeToLnGRH3nJUG9zbSdTiYBzWCDCUvPqJ46/VoEl0a+pduQGbyEhv
sME1qC+SqXirsajAoVIyk3OpFTiGB6Jvbr7puQJge9NpN1Ol2GgnpNwuF7xtsK4WKAxX9kDX0b1p
afwYoB5OWVcbOv38plfDDstQfVKy3F4jljTbUmvHc8Ll4HnOsZUK9fgw2/x8Em5EcuajCjASt/xr
RwWpHjSiHmZqHDyZ/EwdnFQ7kT0DWObjqeaqcTVl5yjliZpvdHJOIUMXU6KQ5Sf2uNkyAfIkGDjC
fla9YnwDdJRg2Tfa7+RUwL6LTzl5mnxbyeMPivVOdqN/qSQyVGs2PqQTnadSMbUYpxewZVOtfA8t
CueJTmbu8Ergv8oR/Pwyf9FNahk+L/gZw+4zOQDd2suemc2f64yUk22+tJx3gwJOVXOIar3NfC1D
Cis5hfD0HdAIPiZB5X5uHamg/viL9rH/zFy8tmmauhzZHn3WFlESY4VFBGNS0wh/kQQRbJ7NWP44
shNfmIlFsVCid9QfKMe0SluGC6WJI9Z/fG+Elvu0zg7ZO3+rw1+alU53mQ15H8GofgDgo+CgE7lK
10Fk6YN8dm1URFY+eDH1sK81ipOUlvF1emg4Aon7yfHQWu4REYNP1Syag1bWvtWYGtzaiVSgKLMA
w2qXQOvpe5gKrdRcHsZbGWgJ/jicZIFSW189o29il4P6WSrvcdFPtkf6Dnz7UZQNKnkPtg9JRSOT
Qz5sK0h/fvuyT/2oRisIXx5AS8nhK0/YoIEkNDe3gOlzWfjn/c1do2OCIYqzvHKLK2uBCZLxvquH
EggP7thTU6fwSgDYT8mesyNzBx5cjyTHTuuemcelV0SJnmo/OWA91IZ0JiY7y8VWPRT1Y9B5kjUW
AxPTMmgqoSG7hRE5Jf/sugGMHqyQqTm2sPuYJutHAGD4mC7mV0EDo9uEHEHtZPj90KhfGGk1mPZE
Mlr7KUzonhKG0NBVzH9zw95OGe7HMXUKymzB9u8aVKS4y+qpMvPow3TGiOfHVHBPCk0LK7YjIGQX
oZ6fkIKXuEJDZUsZtC6eW93eZPYzn1VFSOcxTqotwrvDj+ggLzk1Lz5Xbk+nl5pBtDIlltIJWxa2
MtSr4lCTRV8CiviBeXcPy153fhlvedqjJ2+7endQI7fK1uOd+ZOr+MEhjwx09DeWqV11zvXfot1f
KkeFkpSDCgR/faObeUOXKIvrekPwYSiW/szmk7tW/GwyH/UEMkoyKjdMIv9O9ZMO1JX8+lujvE2Y
OrTJWzSt0BjzzTtcAsvA6CGqE0/Cd2R+CzlNfPC4fgmHhGsegRSSlrtwnZpxXQ6sWoinb12PsPFG
M6jX2dEBKIhPhuTGvC9c98etbF8ViKyaYPq16SapyDNvkzzYjiM75jOagjqDA4axNNaDhKEdoNMy
CHgNn6JV6fghiIMXWGQmztAcr6qOdkmSV3yPSu5o4vYsPgf/GZQutOtlDBb0cCfoZkWRYqmoip36
sOCL8+o4TVWk4izFrhudVK7myCgrT+0B+O+CBcrGM5HPLEpeV8kdS6AKxDLTsSYOz6nGrQ0cw4tf
RXA2SiycPXrTYLgz/7I0C8VTP8/M4mRt1V5Lsl8xuFxXpQfs6hmUh1RSCiKl1JlQAWgIbQDu/gF0
o8k9VbA9OkIZQ07HwKt/eo6ZNeTMYvupKJ5YPzSC83PokE1eQHxDRSdmGK/t4NZLx7aDX/IfUt9E
QYiku0L0t02RNMhd69qk4UHc3Dy86g1NpV9flg5GbGCGFzqsl/9nFLAb0n4XrtC67EmDiv70tcN1
zCELE8XhW77og/fj0ZB1BlI6Cx7RwSD2S+RJW/sKvQ4PbzXt35NYOQC1Fw+zF563IKic9D7Bc/ni
HDcHvD4G4UXKUg8sBy5uztctc9AHFROxY24mNk4xS4RbmbV2gHeGrphs5Vpfm1ACvgbQEms4CSDk
jcz4lxD9le+AYVWJJ7LRvxnK6WCGv2+Q00447XPNBlWI9yRp8qQEcsc62hf/p3bMpGJv4oPPkXwj
7dX6/a05gjQqQa/+HIw0m7TpcoiuqSD22NWEqY4PjKEkG/VYcoBwRFPH7zRgDtGCkXhLg4kKDRwv
qcr3EmttuIWlJH/HR28dnsNEoNMk5OJRdsK27EVvtS3TRWUkC/w8kg/vOsw8F9aIjnImcUKKDEHL
1vLr+i0Y6ZFkRTwujqpvoFmv5t9aQ+ty/+FGA5ztH40wwRaJyzh+aEd/ja68DtVOrM1i+zhfv4D+
XN7Wvbh5r6DCglIkR3fYJJc90BfgpgN0vqtEYFkeRcM3LAVrVyYD+ePh/gQB4/q6ZRH9+aygpVsG
XazSi1jQ6kgX47cBYcqez6cMYrHB1LFtcRe6X4PaufOQm13IYy5odQjmh1i1a3QmnzPXKy5AcayT
6McEukVTrpmUStWiRz62MOX8Xc+eCyn2O5IKdusrZhbqod56F6A6cHO7ns493vuUT2QTDEIuxqLN
YV6lgL6UWoEDGacrjrOCF6m3Cr8m4D9o9WUMmP/1rg6QK7Lrv2lOsf9uGPpJG7Tsb+lLnanrbD06
BWVSxbosoEsC5iBzTkvcjarwmFgR97srUa/Fxtj2Wq0Grg7fdLpl88Ae8WCdyaQWxpdU1E5bUyDR
yX9RTevUcZ3a/uC98UffTBaKJUWe1DT0CFaDqOGQEjFti+zHU0I9gmcTqZTQI2heww9D0SyMnDeK
pO6EWB6zC5SmfVDsYUc13iTcnA/FEvzN2diKORYw9ChO7QqRWJ2RtGrDLBQysItLydPIv3y8SeqO
IEm16oXbNDwcjFQHzWmBvwxZypM4LTSuvZt0hI42SqMZRf4fuwKrmqFym30KMGhj53OS81/DQcdS
yJbCw6c6KtD0Xv5mVKeae6YEYy+o/hyncPTptA3LKNMy4Z8AzpEcrkr/mVkvvftBmlHLSeC32LUP
yteHC9RvLTwnju45cIh1e8MT0mv/wN/wCUUeP1c9k9mHz9krJAnB3KeYDlcgNynWgbVqOzegAdfN
Fw2wnSwjBiPzt3bQGzGvSFPSqKPNHb2BfzZJSiL1LPCyvjegHiDIlClYBKgVkdOx7KmIcVd3HxPI
c6/AJUbuvu0G9I+7j3XNtKuSuOeUJzVsLuZ7SSyTiCisvFOYxTXgh+uuwAqch+lkvp3yewNBfzlS
bOqLklNCkzOi4JMAMxJF6Li7HcAUNJXukJu4Ql+MHzPgKZUzE7BtosOw3ewA0a1GcstIzG+WVnJ2
K8j/5d3fkmXs+wbzciVyCypIC8I8fJdunhumuAc1AqC8IWiWhSG0uXnVGXUwWl5Sl1lJbrb7yhFJ
Cqqv0nd3tTaPwkitCRkoKvox/3yR8mkDkeUPM4RU8/XAq+DAeU8++dXskmDnkjnoJ0+hY2lRRZof
v9WsYPOgHhfzlzlHfBxnlN+xCdDu1gnrLceeUpg4YurEf4zfRuAfXFITDhWZ4dP0yiap+Jz/ntfQ
TBVmTktQ9ICwBQq29YRGgvh7MGeNmCkdonjrYsMQuyxfU1n36SYeT5RLBc4W7BMTEUkp1vIgYlge
f1biWhZr7w0GLovywlb/7gsBJ57g49Bo3u3pZQKc+64AcrFXj+CVDgNWOzyXCF5x1PuD2+r3kNHw
nkLvT2sV0nje2rvxuwWQ+HHHNgPZ56lFqb83SEARDVJ1plnh/NRHq1TMvNQckUUXtSKkB2UGcRqB
VnVSaU+ODMdhzJX/gv1q7/3zVchV4wBuY+yvoeT2LP7/pdNu/GZCPfhiz61n0zSc9zdaET3OfGDV
ihkStlFrBXLAx0p75/4GGIDMNm/y8v+jHuT2NL/QrPctcDL8SE/IVW8r4Of4h5G2pdnqA2sfzj0A
ojOv/O8YKZiu2QNSmb3Y/Kq+FVF6ai0pUALUT1jdpGBaBknWBMjsgR6i5EK0QeHQYMQs6Gzpk0iP
IH6eJsVpYr6FSKJiwnwauxzjQBut4TxoCQzeVGbzA7TYqf2/SQJ+rrnfz3K2JdCuzCQcgRWi2xEr
K4353ECdDSczaP1MnEyBJA/hAdtg4OphtxH9c/oQcpQ+DbIbufuTWCDxs0d60H+V0D2RcgHhtNai
PN1szDxZ9i6RL6qQDdyaaoPxrFPwzrRewNDkQQgcJYom2fj2HxGqghu+hytxbUvU3QOvV5qNn5El
MWOPRbTPsyBT6b3dXLn/NAnYRYMm8VZW7b1jjFnvI4ABlXVaGHTREdRa2HqEsuPLbn+DDRpzn/63
nHG0nW5xtogWoiNmyhxdRVohu3T2jnXy2AgLcHN9kMkFdc0NjG2Q4iTEkoyIN2q1w5ksH0Ub/Onp
DzaGyZfSP2h7k/mLwPHN2XQS9nwjDvLX5EQ1i4UHdUNWo7ckT/YSv/K1dz7uOhDYBml70dyC8TnK
q2KG4aVOvh0ipAnwtqUy2gQF4mtuRL8q0Hn1Snk1DXPGaBmkd9bQlQY17JTZ5iojMBFz7r8nWOV0
jaD9OtCD6FaHMcvuNXnl7WNLTdaUclzIMaWXAdkZwA04c7tFbNpaJccITxSOMa0wI90o3s0Rlc6r
X4uai3f3qSuvcPaT5hieX3cLUVYe5RG+9JPWGArfxlK+Ij+vwTYNoTBsx1zd8VgGIWYljiv6JLW4
eWQJuxpJZiD54vxSNa6tcjIm61ar8hGH+WCTqTBhDp0uHs8BoxyrJnSfaaliLGaRyoeahytbikfL
3RB1mtjmObMlsQ0K3vG3+Za5IAMnJidTCKMhzvVcsHnDiILzn1p6FODkbLZ3rvftkqRS19xdmumm
pNRW1rHcfaejdbnp/d27dCyleW9rvz+jwIRf83rtirAA7L6IVRaQeMBc54xlsCsIUn9iO1logYRV
bf5VgqbVpjgFkAu90hvBT/YSzuPwgpNP07iXDMcgNgYAcNrkX/OPxC2hKhQ0QENbd6WfAELXz5Eo
clk671Cv2MIp1uOG7fVx5lUtXYPBluCUUedM+syQf1L6W6zAq1Cgw7mvOk9UmQTlNYw3PyvXFk7U
Bqf8l0VIMTFBG4uXzqI51y+ELj3Gb6xcq5wjMsvCm4DLbCu25dJWFMwF/KsdYJD8O9VFq5TYv69P
MuHU6S8tyqQIP5zsBoy4t3eLRPhOTA9NR45rgoFOVeZLmkI8/EwJedyzrxIXcq+k6O61TtVdx+XD
Q/urJIfmoj6lMTCpEpiJpHM/yzCypnpWxzFd4o+HRxAcICcBmeljnfjIGnq3mK2zQA6TIg2hxKZd
JO6cYobqeHMaZ32l9iJ2BaZNy+yBQzgcuEalMZPhvW7z2+e2JKlQyd+295Gfa16YmYYmRyPsHiJt
v5IIMJH+nWnVrTDNMFtHXkOCy3YYtaVosVRrkmmniyJMYaCkiS2chPZYKtsRMGOhv7RH6HYa3Sy8
8STq/aB3GwzldwEe0/7bwi9e932uuTqv1ZyTHyHA6XzsohhvgYWMcKiVnnX7NAbJoxA+ro+OGkqt
Dij6LHt+ks1i9OmxnUA9mH1s+JqTzFQp+AFgJm96QBPyESXJhyZzwa26XmLPZZwouqMNPbGO973t
QPPmWSo/WGfr4LpzBRUSqLzvpqRWK/uburL/4JCHcXLWcyiJylygyQ/TjwBNjnqzka7dHHakSbYZ
35C5G5yVR6iGTebfjN/+C24XNYc5PBbR0nZ4Vl6SEW8walUgI13W+3jVIheRvtjRx9YXkBXaALW4
xIe6BKqEWE/0gNSYASqv0Aq0sjrx2oB08u2b37OU4F/ruwSqcmESFk0AYbZJrFtSL9q3VjzZmx06
UxFJ/mACG8G82oCFEf04zR95bYVVDQZzzPpC93qv2+KUUyj6fjr27EDhdPhRjdqleZSViNOZfaoi
lKFD8/FFlzCaJ0btK2GwO+8LCgrC0vCqdw3zODlHxfXLY3tEnXld/4ny5zwVev7AD7N4KBNWY69U
EcObje39mKAUmEqyKiWZZDHWHECYPxo4xVM4q1He8T+wITQX3CmW44zrj8o0/3DUlnb3LsgvYBnR
4j8dPKlUG+sMT/SM+sRLLJ+AIdN3LBs5SaiYMaFg+oXnbRM/jDgryM54McR3VEe8EgHNGw2+rNx3
DMzTJtolBBmtAHpgPgwzukYa2Q3w/z3aePuWhE/Cp0oB+Zieo/XStDwIutq1ambPpLx105YIY2ib
JwICPjdt193bk0zP+nIMjqrHuf2NpqHovDPq7oUOjWqB5RQvDExo9KdMV/Qkms/DAbC1+WIzP7ow
8Hd8baVC8JXcB7c++n764lioQqyo8BigfKulRIJlQZn6lEXtSMLDxo9Y8konzQd8SCQgKSrPrLqV
0z3TXgFfBVNQsFw7VjWw3LjqkoaPKtB8xFNibO+PoyuyDO9C8oIlSaQCneBpOJPRc8yeKttjLnGf
Dmsyligg/dvbPoCGL2PFPhbACrUoIlelpz+JG4Yfv5VcgB59ymXPKJlyy6yDsQPzLMgPtTOUCRPc
ryyrEUeYFToiu33E5vaTyQmv8JdcOuL5Ist4NCfD958s6giR0fFqrQofny1Br1IMpNpMCxycgHur
AD3mOArMamZmQftKS5Xr6MX8Rb8tr4TwIqylxeqnUy5nI35hd9e/DB65BznL/svG87whJ6NprEih
jWdjMazX2FXu8PyulksOTDdoZD+BWzrWmZ3omScPDsNVJuLBtpQOwj4IQ6AHFMgpUHoJ/CIgmlJ7
AmL3mDsUclNH5pA/pQJaSeXZFuFVOAFDetCgQc+p4MOz7CPrPzupuJFpJ0bkFTKTXmhjv2NOfXUu
mKn+HkXmGytAN60Zad9aUeNjAw6vwWjVE5KGR4iHmEpkix72c6IvU0NJH6n3jUeRj0mrRiRq2XJ2
nDDLL+DEZPg7p+0G/vPaKMU/IvUKJPfV2S86EtB+d+u+Ees8a6tQF0tYfQ4y/u9zi2+tkgChDC2h
knrEgCDS9hTlg7iOmN0szlhSfRmssE2a9ZtPmE2PTU9R8udIIWWrUdEBOw7zG4r+Btm0/yPBom0/
b7WGOo5c6c8L0Zg0AOrDwyUXDihUv32+KRgHtvWGyvTtDkAxtWuWlj1Ec0DPx+HCYNSDak4Fsxf8
tyyXyDNqpOib7TK7g4hI0JR2ZaPRyyguHVj1GXE9MXuOPr/wtRG2RL9djJhRggvsWZkbZI00+Cxk
2P2/jtYl0l3E/0knJkvUlbqDoHy/ccc8WZvvQboXYmHM5lAgFihTUbcrtgevO+etCYqeARq7IP//
0UMTwkqHkcQT3y0J7rCuo36ahsQLXLdhD5awS9YJMBSKeuCT4Dhoho9AR6g7vnuCBtu3IFe6ZUE9
h+lxXmrDAGTet0I8j9URQ5AdnpWD0wS/Y9vFvKriLfImiRVSOkzhtdx10VpKKL6HWcdiucXZPTrq
dbS2oLtblaMLKlkrQQLvTFyCoPM2olBeIv00Zz3zHFKAk6egbfSXNewmfC4ACgd8ZyjgVx120sgq
+08FRLRMURBzZWD9MDKhlc4BPp8MeI6Bx1nPUuOJ7uGsmRAJ7ajAK/Kka/anldNDqdZZNlNA0tMG
ZGDuEtxUzJFn/Y1m7MwBvFNnTZqaI+dLt1qwKr8WrhjDdDYWMf9rETKAVPKcDPYJNAgLBuXWgiKq
vd+Rd9Z2Eh8A6GhJpF7yq6zbGuRpioD37Xcz8TmPya7SV7i4NTtLx1LjtmEjuvauJl337nJJr8sB
Xp89gpcc8hTOt4AHatFNmf0KWJl67imhUWaDssqK/dbk+0h9eoGBIrWucuv1+Mknzc1PxL6oPHM+
xrjLj+7UmojrvQQbTPXRdMNDj2qAIJZzDT3XFPgZZ3YigV3jOm3IzzXbEy3nDVXNzGFLxk8/+7gh
kiDY+Sp3wLC/uDdA8wC5E9aIq3LJZfWdNmR6bpNbXcpRMN3Kwcz3sen1gSiYLyyvjR1zygpAzCe3
l4bS22+KaiE1NKYqr1qsUm7W7JUS/+lrzJ26TZ5oiuXN0RA03ujGm2F+1IIhk3po6ulyUUPXoyhh
2yVWH+ZazlcXHGIwFr7PmupK7hCVWnILXyHcA9xEBoS/7XYlGcEJUIdwzQwZdmNDgakM53rk8Yi2
Bohx/OLLoN6E9W6fdtTPqK/IVek3BAMyiqUS3dR593Ruc49OlLCcLjuxVfD15V6KI/v8tMmgOBgq
uO5Wj9hDym3B1bLYt0DqIUlgQvvzRlA17sERz2c04PPA0XbZ2+5Sjc6//dtqHGZH1QGXmd57QnEe
/CevcxTQWxTtUEfIf0Uzik73LxwK3LUu4zom3niQ+BySdkaZiY+w9aScHdmKdjQxW1c3qQZ257kR
P67acs6qSDFILN8b02apBrcefdMynvlQHQ5/n5XZzr9RMK/+IE1Hg+KhaThCEDzfHivn/Db+MkVZ
7yj8ym/A7Xl1Ry52m02FgVuUZ8wXDu2oBwEDihHdMmZyVH5czT+3FbTdpqg6+MvSxuh7qAeQNx4p
USi2jCVGMoz0JZOy20hK/xcze68bcCRNy3BPcBKI7rrNb24JSA4/fKf6zbLBa3ykiyt8JqQ/NnK5
CBd4biYSdZ+h644D/joDdRht4jUIYzCtqDRCJ1YOTcapIdrArD2Jxw6OBMSxXq5O6C10O8RFkkwX
fBaTA3+K0O9HDoPZ4Ew8vV2Wwuw7DxDLA4JB1WyGZ6tqHG3ZjZcyTN5YAnvuY7J4DZEre3XcGGH0
knHX4hjnn+nm/rt6zy9DkCu9ipYTU+uNeO+1g7I5XOkDEyv0YSzEZjPMC3lZnLGlNQTUW4+xv5Iz
t8OJGPPXFBY7tpbJAEXHkVmEyFZlc4gOO/JaISpJQ9Na00l2p2BWLTueskrfVdSoWyquIS0+1KOh
A1J0myEi7U4UlG5DUJz7GR4nHINiNcCZw008ygl0F/jFNfBFDuVaRz2NQG74j+vMOrWbOk9/f1q3
Rj1h6jVDP82L2lBgaz7tkqjOAt7CqlVund4HJzhD3mgQvutyjmOns1mk26TEzIQTCLY7FRhI8Ki5
sGQUOrMeVMg+h5ybew9dulR0INPCLZ17djKFB+jrpPqnjgeScv6k0tneiIwB8UDXeewNl0KVK1Gp
AH/ztIh/RB+gv9I/lpXDy1/hE3VnRm9Q6J4726CemjbKU6nT1qff+WAn6eC3JYQbYBaL36NrEwYy
H00Sboe3PoDE921Cy0DYhNIPQtkBbTZb1lNtGJ7RaNF1OlgCzq5WHsxd8/YCcvN+EpH5LjsurGIh
LcvECNXA9jzoIoWzfjptGHNT53c4RajcTd635BQOW0wtpQ9peZaoAB4cwIiSJgqfJNm1DCrhW8q8
jy82yA/350MJm/gTl/KUmJ3EmwgCOCqBC6laBMJ2KP3TxlR2NVmOTa9Fv4f8WegCy0pI4n5m82t4
MW78C9M9sl9gpTYCRX70rA9GEEnYRfzSRwir/jzfahg7kyJrnzQ3atpRBA1960oeC8B5KtBBsaXf
VGhJwccF6hkksR3EPSXa8RRqmB8ur1VoJNilKzCQF+jKSw18CBnei55IAUd4vRkFjkSLOFKAAzMy
gFaYQC6wtypaBdwVhAj38B7H5bqBdqdRifc24Z2RJcXSwuxonUZodMgXCupsQvwD/Q+QAuBwQLbB
MtP7DlGQh5msjhlOqykxtK+cMqRbNzwRFROQrKkqAaDnOTWz382ATYKkOfslF59FfgTijDlvrnmF
vdYPyYCE3472UfGdIhthVmHX8SNNDFtK6m1PGaSdatstsFg+avQfXRMBJv2jmU05ccfdZ96q7IPB
GpKc4/j9bZsu1e1meUHbt7gwPsXNI9v7HdhQAbnqGcdanHoXJaQ74NKxGmXrhsdyMcPLaKu2qzsx
YBCKm7PfTI3TKDBL0pU9Zd30A1aGWZ0OsnUoeTievXS7rMQzKH8nZQmKGBLFChRyue6h/5AOOAp0
S3HAh1zwksoYoM1dBfx0uKhAgcjgxcgBGvZk2GOFew0ZjoRHDA4MwKffxxG2c8+poeUVXOlvuddC
uMn3u4nErWFjmKYwnqXiZ4T1ZRcACWdxRshgDxPqw1/a5xfTmrPksHhmlJr6eSqroM74Zzgt/qS0
J2U+nmtRhoYz1tfJg9Drtex0MPmHvY0aSvfNkkRL8FFi+fOr53emfsQyuOPntclZuQg/8Bx0RUnM
3IPozkmSgiHpp0OBAs2MEXypzFTqJgSPNeKCC70zz4u9a6vBAGs9Jd9GVqaJuue0yzejFx/zK+8r
FvM76tKQOXs82ulkDE+vNL8kMOU6YB9dSTXOA8Vp+HF8OtI1TGHhTrdtHgBy5qpmg5BW7bR2ZjCr
owiwiBGHeC/mOMAchoBExcLgOtLkh9aa6IDc8F0QWQ+uu8msM9Tvfu2FQUgQZgAh6wEVrVVHc7br
aS4D6J5ql0a3I2umkxR1oFOqHBBbYvDkrxi3+uqQO0Xc9RkR9bTL/kKB1/9TfasM0mR7dsHkMrP4
SqiQukuHlOcvCspyTK5XaxPovRfJERwBSV0EQcdVbD1DWqEMje27SET3dhLpvJnas4duOaqcU2RX
jt7696fZN0Ejqe9dKMZXx2Ad+TdN0sHFHkTGXjFHZj/5Uv0wPkSUsmsV84afcI//1Dn2lgHf8bzx
Uxd2YqGarcRFl81uOMMLB83b37PS4sa8IZctQZruvQ9xzwkidHPghTUIWMMqvbq856/dkI4MdKjE
TGdaYvY7gQqeln2Q3nyMhc0TvQcdkO7wYGJL/54mX/Ul6VPsOIb5Hi/qXzYIo4/MUTMcICFMl6AQ
I2bQ/x3pKqQ8kBq+qaTXLC8mlt2y0+XX8vig397QLwzr+zwY8gdUJXMmjkS0Mm6nj0kWaDliRbW+
cyLraFGJWuaONtZJCRTDnNEbXuPJc2aOgnghdTKiprO1Yo1yPJU49gBI/o0Iwi+QP67eDMNWrGiA
Swrd55AFllP2gyifAaW8ITxwthShtV5G2ckqzb/xTL8g5whGkv34hI9jPHHbEIQyeCroMYvRCQPi
nfAjb78I0nORZBUM9XZFZ4LDTj44Tyuu9/07g/LYzkTJPnugawbSHChQ3Nb3OhwGnhtI3p1wqvbk
epCRWgIT5txZNNpyNYgiyQ0MYQfmZeX2YpVUoJHQCX2WlYhltZ5VcBABDGLpdpMLQ23UGv6OzLq4
BhAqstLsTRWi9iAbwLgNp3WzIuv+57DtD+K82+dsGfgl4P7iTnSouV7FPI8TLfj0paC5J0dZOUjK
pOxkjx2gW/eXrV7378MNsvQJwBPbx50bs7wY8ybzrhJ/dYvxVi/aMNkMphtEc3585C/2RVcPKBiV
J7h7El/0+xY44tvonTsE9HWXe31iGC8QCpxHF97NB718MPsVR4NuUVvVO9kspCplH29wxpmehOLb
/5rORmUcuhmjIhKnpsWCR/b8J6UkyYnLBptbZcEujROczy68jFfhpcLkLGJIDJPt9FqXMmu898H0
v4Z15yaDtpeAUwxTLyl/7K1zipmCz3jb3l+XI8kDQTghd1M/I9RgYDeg7YdAUAAFcdMm3AQtOQEE
/Cd5/j/BrSCNI1EzTBGRZnPLmW65krFr+tKqf/hcQYwefsu3zlnQx0tJGRIQaQNNEYXHc/ilzL91
LbJWQa17a/VK1CmPRO3rdOII/ereog8kTHG9saIW+01YJzpRkIQZxootkPUJ9ubStapX2u87Tc+N
0zuQWyYlb7m2mRrMcT+ooLLqFVZcyxI57RdWftpTkXYd5IUPouS0qLGHyDhzBIBUKyltqRXDfi2w
9bPm10Nprne/fgs12wLjydLJBakgF4CLOW6To/XHk2bEXE07XIdc3mr7SEB5PFGlGrvoi/99AMd4
s9yzGwG8q6Nfs6NjTHA4yqEcs7pqdl2rcNtAXV7RBrec2x9SYYmDOLbBewvK98C0GxylKCqClekk
+jvVOfZt/6Ae1CwZaRZ39wybHd13YbujPSgkUjARPwDJ7+r080zaBpVSJY5NMmXILRAqMBG0YMGX
s41FUyGWTuKmp7d0XS++BLIB4eQDpJTx8hDz6ly96PuavLGDJe+05848VjSMpi+kG9c/exX2GPit
jp6QB8gFxkAdVP4X9DC6RWgkmeOEQ61Xn1OfiRBtD3J6UlttkSzMaMAoS1UUwV4STpS3clNu2soG
pzhf4qYm32YeTG35tEDIpenTobaz1QikYCDpOSu3vSY9MjpyJsebplgUSc7a6bMYWDIkRhW0Sn6L
9onMWHj46lo6LXuWFzudy6bJCMswF8YVAmDVk5ExLKY7Hwkkhlvorqnn/e8uQInzSsq9L8USbCkz
uF3Cxoc+XeGIrpFWU0yhGcL2IK7nmLX05yhw1p3z8NG/BDxP7amEC6abgOvw7MQwHTGoxfveQ/ZT
zYvbz+mcw1xHvIXCHpkKTr9itAKo5uvuelF0SjC/rGZjK9X1naI6XKfA502lOR2NuMesO2GTFmgI
WpOfmnoDWtL7HIsHUJO1PiX1Nf4vcybFDRF985TqgLRsjdZ28EbUte+9HjZWxF09ta0D/BSos6Po
GnBfyfRnVqdE3TzOrJhufuD59K0UkmMzWTs833EFB5buyM2kjRqXrP3N309IxoDja70cMPK9X59t
BlllXGWTFtB0Cl4mmvITlCinTr513ycE7Ojq+lN1askAbhjEC2LzHdq2XKt3zZUNlB8KMtB2ghcL
FifXDwPTrzfE+EpOLXNcm3jggeeQjQ/ld8Mv7e7l/YlVHXz4x7mje57+sWGiV9gnXj6bNqDpfq/q
7BUg6abhglBmXSo4NtQ7MdSDONmDYRlpbY/SioxK8+7rIJHyXfovZCwmcz0iOPNIbRMD58qWpT9J
9A5PNOTr/EZRsF3IcBfxd0biGu8kUdCz0NP8WpHi8OgD4/xhQyY7lona7HyHjBniutmFuunN6AW2
zWBa080BJghZxcjekjFHz5x5Houmd4tqz1VAuDcxtN/AD/vihijQIiOW8POfA/LHtIOfhPQC680P
IzZSygWZZafHUO7hrNI71KaLO6pS7OOgJhkGgnNKYuYGMNucD30NC3QDiFj0WuhQ0lAuRPo7bfMo
UogP+P6nXY9d1sOBgtm4/HuE4xVngkUDzGoKeH2znBO6N9lq271NN/4uBrizWsgmBV4TniLSZTzq
q6bIjwmERwwsixgz0QZy/5LiafAEuI6YJ2/h437X91sYzBrkL0Tp4Cxr6xEQRoKAs63k89zDsjc5
hE7/bT/OD7+lguEQTePE1ZD0ZK3OGQr6mTgoofPUCbydpTRdiWT2Z8I9rplKY6374UO1urt+k7U/
SMdPEFzk/ho8aoCz/dbs8vvo60GLvMJhqQinKwwcJ2UEKZ4jrgpuvzNYNFpDlljU+34llf1WBrhY
LJVxdRN0nibY94+hwo+mIPNn7Nx4jXnTofigAhLL0T7uw9q4ZYYpWmew2FqxidLNiMtv9Fdhmjdr
wnYv6HoHK+hvNatrMafTfxl9vOosLHTxExdkxSAI1veJGHt5E88mLAVPqAuvM5oMXIJFhd7Mxmxh
qpnBpjyRn3zKdOClWYS1u5+DXDTr5iSAxHmfQFuyqMihFxjCd/MrKpZrsTvn7ot0PV0WvcVFngt0
jxPpKNDR21noyBVfbfpX6CGPJ1s71fai9QoU0ZU4V2YVnOPiZmTWDCWr3i5BDi5qhNzSYMzsdQNQ
L1zolI3QOa/T6ixxwqxjnazcC23cQXt+8878CLv4nbwB2ug9i4x0cM46tmUDi0CIt7xvizFGScmR
Dwp/yMfKoDSB344S5G6jtKkkexOeXDoWXR5raYJgrfBpWu5pvxr/t/n98f9vOZzconJVKsj0P/0c
UKffM8WO0o7bjFxckEZdcijZF8+o0R0b2C9vtOqpH8zr4UrqMlJWD43e5XCjLE5fniiaCJO5Q4Ja
POdPizHGLw+7a7UX07VQ8N5eTYqMoITgcIQt08CSD/KnJmBck5MKxAEP6F4fMZ/sUPB6bSMzfBiE
wqI8jfacwIfJKI75z/tezW2Qsaw1C0Gru0dtqddqDuG2f8v3OgDG7QIBQwnlRXn6hxX8+HhiNZ4a
/T3YtYCtKntc+EuTGWY2YEtXWb4mGKoXjNXjwNPpEOAmzJnmB6GF4il2Vti+9dsTXMe6utMuoqe5
X3mwdtSjSOUDHVlMpf8/Z4XfzeJQyFddtcY7KEwfe8zQ7mdC1B+hLrcRHjquhA1Y8SPYa4LDdzL1
F+HpVALSjNIu5YJVFjLdSNcsWb6WRGSzKAGrgGNYPbr+p33dqEhgzSqttNR/Ytt/iqNIOyRGFL7M
JnhNZiummDXY7vyEzTR5rOpEf6+L6o/jfi++mhyMRqCluSD+KtXYxpD6OycRd+T1E5+2m9YBZpgw
tORliPbXio+ID14aFv4JXPW6knmit3BIcgxtrTCyuI6iqyDgwCWz/ZWshRzaYgSR0ModHWKBmFQ5
8rdCDICTmezcqkxPWdwsr8fbRzc7dYWRDmb685IyZGnSD8mEZcVfc3YWc1aUOM8Bpc9vPbhocy94
1icFVuPxSIpPRAbjLvye5ivYryamifFUtFSYDNy2aIOBtt8qkRjOfBThiNoXIkWpVXjHYDnd/Ted
eDKVlt1kHQMRVdgsEeLtzuNjm1G1w5HnTEeTiPptoIc5URZ3rI23bM1ra2o+d7nEUIdpTa6MvOHm
Mp5TqYYju5/g56zS0k9f3kyWx8KOMVm6w1uexHQyk3pUQRMYKwlkf88FHc7VepB7iV/O0MxK6PFy
I0SWBX9gXQAnLJyuhe9K/Vz/rPbkwUDzFZGIUTrIXpUWwclx2BhWNjbb0wgrbFoOqlvitjMW6Hc2
G4k6PpQJnaM3tRP+hldWfZNpdxcpfIgeTeugqS3A1Zw+vgqOEXlQ8ZUKdr/lbQ4Hfq5iohvVgqXw
SbByvWU31wUf0MNGhkki/N4+9sh2Mh4XeUcob2Ktt+5lw6SrZl8T5CS3AzIzXU1cjtcKY63xZ+Um
Dl03KJitsM4g4ZND1g1MYLlG8ZhZZ3rA4BD7y68f4L9fR3lQteKA6VrcvYawXF5BrkGZtpw15UFo
gYEmOpCacW966luAJxOze5LwT07QuCcKt5iTPXGwwALls+QkD+xjw4eoLeSZ4A/RlxPnH3av5b3p
zoCtmtLFhxgXicEWqr5TDd0oGzIeMrM57kylp6kDorYyfj305tuB54SrgvSdrOZQ+nsugGXR2VjE
jdJr/5ObIKKRgmqiT/++p+gVbHtIKE85eplz+E7ZwmdR2u+0sH49SKTvqUfFEfrDwesDDdBuTm6n
Xo8miAJWnEqpeE5qbrkgv6PjZAA7JcLHtrkBdXvd/iOJY9NAVRBkY3+IAGG8MUPhMfC7OLBaj/Fu
yHH6T+68v5CQavrP9FwliBq4qMSj3l8Vd+mEwcBPMMAFKL3egQJUG7m9fx2IR881ePU2An9NPYR8
caxas42JZHgylNkpDphsuEMtpVfJGKWRBbjN8UJJtV/QJDX/6uxg4ak302vKhEBrnmHcEI1R+Iu9
z9HhgPyfD+ZzapJJqHGi5hRKgr8K1giyWszn2vro958778RcmKTg51+ILqsY0EXsU62n/UVsRnqA
p5M7MOSKEa4n4TZUfQqtDYhTNpAJQ9pkFumWOZdyjhQwFWkLCFioYk8gtazcaI6IfSmcfRumBpPm
4hBJPfE6lZKYhrVgBUHe4oBhwKt8VO0hNO92cWTtX/uGQMBdKLkxlynMgGaRi/igl5NTQ9Ztl9UH
XQ3yCyo4oVH6bn+SmbdYMGGBHfDkxmYvwFHiGTFzJXxe9157yQk1+NEBXdWP6zEmORuJ27LYknSU
qFiH0Sr+W55z47reCj2r3mySxDwC0zNM/OpdYKC0tWlObxnh/haAr/F4MSXdCNhfcInZGD86Kg6t
mWMsiPnYTXYcxCiYmpwXUHgNiLVtH+cqNuuoIXDu+uF7BBTObBF3SoBLCWl2aB1OmBOTlAURQKnH
BvTAj2YgvlAUWgbvF0clOHTySHj/gUhE3AVcL/XM0IOrnMn8S0BOmpyi8kmc+I3OHBHcgiEZprI4
FuMYhYllrj5Gd1yIUEd/4AR/29fkniv3VR0fFVzytvKG5R2QDLH05i/IHVkR1Jb7kG/THeSGl+vR
wNfY+dESkUFPgFEE8Nuit+H3zTx4wp5XTqFz2yTY9xxBEsPe6NbPSA4HjEF/VtZEkMK0kzQVuEdH
n20XDhr7EZpFsdO8IMkgSiY07AAJ/goUz8h84mvVdYKNlPId4FhKK8r6wDRYKBKPCEdMzdBoMPjC
sSJ156f6ngqNpONo/uPIZ9Ko9dcHQt83dUhmY6WzP7b3gUqRc08DUnNzdX4NskOtjRy5lzteDHDy
CttTJlHzewv/H+NqGa2322IHRHzUCQ6PvQAbVCjJXKUFGOI4zP9HeO/X9Y+Iwljdd01m1/gStOLt
QmWWepdF+VXG6J0ZxrdvLBUypgZdNZLe5vnQhsHTH13bmVNnWX7iAVFBErE0h1VGie7YqPTRopgK
QtIVssdM6J2QW6BaTg2m4p8Z4m4Ed8pggJhjy2R7EyuW9ngfyZyb8U5T9cW0FMtrDYyQC7Sm2plQ
VAll7r09pzWKZ595edV8+VyXR37gGP2m974OIgAbz4K7smhDnHCsIiG1h2b7oFkSsv4Rv3p3wCSC
xQGzqEtdzIQXdEvUgfTOZrHJTYUpvvFXG858Px81xO0/j7ssRrAOU2f4gD09KXK/nRE47xzAA+lS
Cj31oD+qJ482dO3BdJwUBYoLYMtxE3xPeWf74GbyEKMC/+PG+2l1auiwMWJDPdhKMJAqxG5Vl21l
eovmNWc3UvyIpbUg3Jjnm9QvscZPhJyDq0L1Ra/LLQ+54CovXJ3uX6xtgmnT38JZsuK29TXghQBD
Rb8uzpjgXT8oRg4KpCcDAE3gesOF0Q4JNGJWsgz+6/HVBckkpUydz8xTzwWTa9A99zTdHxZjqJrG
E/q+w60BeyzOoS2NPMlS6fGUyGCip0S0ZfuRlAjr/7FRwz4+OKc9ry5i/PMMjGiOuETaHWdNAijB
b+hvlOpD4Ogc6fFORQwH16YaiiCGUX+hZyLj67RBtH8nyKA3tD9qRfoJEsBOVUyi03+HIH69Sjmt
LgFsUjlrKYzoOTjOFJbr6NORlk0xziHtJZQfQhIfa83Bund1oIjLppVhk8pUayfL3Dzl3RpAZOtl
SLCeq5sZaGTx8pTUAOSGj9+pv//268N7SZOe5jv8T9AyhniZXwSVXnKFFlHfRAFTFsBK8yIeZSIl
l036U8ebp4XkFJmDxjzXnPugS6/FO9tEXnizJq4SIhFuI81MBMxJeKFJstM1pBxNnZN+h2bUW2JX
KLDUEiHX7zOJcQyu+g/BQcNhO6C8jrIad30eqJpuZzjKEplKYJGMIEkDi1gMUYSysIfr2qWZwVmn
A7eVKn7JxLa7H9yqF1nyDERCG70El9+MmojPrK2TaA11DxLt9japkVccNvMAk+pNfNYWuGiwSGg6
d1TQZWbhtJAn1/AE3kaHGruC9mYir+4eYZaMjghfRPzgsBwq6eBnGa1Vv1A4TJdWwE3sedZ3j/Az
y2S1GfRRFbtAIbcTEnTuweSwYs292RC579dgXd9l/3kyJ7Lct8A341s7knAIWrm1nnT6QBz4OX27
QBydE86yeXRFheE1xrCFmTZDV6ABg+WbAu5YQ3hAX62jqgcD+sQ9MbGT8mrGU2Vd/ZoOCphcMxti
87byPckj+oVAfR2Y2OSnAFG4IMtFWmBNtBA8SE3eMFE3B/qwcBg46HpflPPqa9keINrbtHAtyrmd
YB5X/J4s9ET71nZb+vpKJv3FTsLGy1VLSRwafLoJQOh78WzDCSJEvrxPo/30b3Kipva0UNB958ti
d8zjSj/HBMEyUP+SILGD45G/AM9uRYui8++xnNO8YqyPPPviY/twpIzpBHLqTTbJcx5c6UIau1qN
Z+gxT5t6GIAwsZSpkPENA3Z8p+zjZq+JDnsbhsOaWXx3uQgb0CvPLuInLuzeiBFW9K2V4rgxROCc
mwrhg4emMkZ2dNVXUC0g7gYK6flaqBzgdXk7duHO+GLh/ScxryJTGU6wQhlZFs6eDXq+nuunYS+s
33Iuz3CuAzl5N3Pn3NgS9AzkwwecE9nJfcbe4d8xVAnG5qjM32B4RU94LLSkPnVKjeUcCOf3ohQf
ZbkPi83TSrPHIx7Hh39fhAXWHAYgwHqt7jkQr0/jGPHBS1QKmJ3oEbNt7T07U8d5UNnm7ptE42KB
H/OLaAFiW+XIh13t6rRdnpPD/2ateXkV+S5o7cMfbHaJTeJSyWT0hnCHnLk7hUfeZAZe1mdJhDBz
xegJ+fBLHR7ZijeNzpKYfQlzNwIVYTBOFInQK/wDwJtv1iyYgJBZyShffkKDl5H+zpKQtUjclvYw
cHigjDHDFHeqvPzpOSmTWH62PP5BoJtbBHXB4sW/enG5NdeYdC/bQQOMvrk0uNxqMFsdZP/K+gan
lR/2fl4tEQM4S+0Bfmha2ZGWRct2xjUY1+Pd+H/23ITDMlaCFQATAnGhwjacDwqWOc/G79NaxYjC
hbhb5zla2zSzLB1Kf6TSdZYCKS7kklv/M8/8qzohR1buK5JaDW4/JuNYxB2QmiE92o707edPgkQB
731e5w0tNyZ9/Bs7nnmVr5tIUV0YZfv2FN7Q2KZEHKFDuQMqjPR3/Pun5pp2pn+6FPXrg9n3qZd5
1SSxq4tZLsAKRd/DTQOSZkD7XJq5zt7dNKE/1vhvCretfGxIUNImRS93qPkC/D4DgqF1ziXCSBtE
CrDkRctLuwKOPUO/Q65jOwkf7JndB+jgFKZSrbZdcqjEwyVbPMJqV6YCxb3pkg1alJtTgvzILyyW
zORqwC9nQ/jxIo8vK/VQWQAEhebpM++c5vcyNwqIO4foKL7wpWFv0gj0EA2w6m9w5b2efPtfutGb
okZY2NagUsKpjXYb1yCn2dqKJ5dKIHWcQ3cZvRUsJM0UgbRpOOin8Tqldv/KA53h12W6DnEdJSZF
xb7NDW8RBB/f1S3TE48LpilMObMkUdZp0C8YvvLzjXt/1sFbV04iCiOlKpuHGilzqqrcBE1scp09
BLvEkT+5U4rh4Xp1VvrNZUd1Spb5Y2fa/xiaL0ok7siZdcsInNryoZo0/9zKZD4zhnJTta+eiz6b
PEU/ck/oveTCc+3uUCNbb24xUP9L0bPqodbM/OUyBd9dGh+kpIdDGw2VxoPFWNbhbydaZStzZdqM
0WUbrei3dAeKPO+bTHITlJagV46uyfcW0c6yVqXfHtPDbWVZvI6W7CjU9H+QocORHuBUKBNRIUUB
SpItrzHshPsBQHhBxCzrBcImjNXqu0ppWMbR86UCjPEcqej2MHXK0JXnrNcGc36U5legDL4IKwjH
UY1NvDZ/x/M0PWKo599AVz5zz/bNH28wm5wBtfXLbs2Y3WXJjRZgKoiuU4PO+Ka0zIcC9GidQIu8
n92jBaWA5l5w7J6uYqKgTWv/uUwRQQ+BIiTQaRfDb8vNA/Im6uCmxm5/leAIeRpuuUOGf5P2W4Wi
sztExTk3CUSbUmdhqVbj6k61F0S6AFi1m17it1ifIceaG7etOPdstk0+QUIa3kReWBr/Pfg+3Kas
YCO4bwr9Hhe1r04K1X5OQc5aOa2nHdOTwBvb5oKJ3QiTSPX1OLgBnu2ucle/x40I+XEqf+UsvaYL
XOaGYHK6ZWlYTGhl7I958+nU66cghznpqoPwfZ5qjS9lIa0GC8q4pfozcFhwLcJFmWQ2FLa0Vvj2
hc+/2L7GgJ+T2lyqRuXZY9go0/Q2VzVg8b5i/FTfCzfivgDK54u8p4tDhqWb6Z7gZDd+f4LUAhPm
55oPDvh5V98WZJvGfECILlzIATJgsdIzxSH7HlV8k3Sz98iV8lN8URpf1P1+vIlYhhViK2QjhQON
zyZmEIkm0zuBfqsvUqcAThO3HavBUWkw8gNW4oeriCwXHu+N0uTczksRY8BaS8tqOxIQiJE80Xiw
Ye8Qh5hO4ROba6hFSCMqi8ektBvcY/RxfTw4PRxg5OGjItqEZYEy9IJWTfXTSftpcvFiwvQUZIGl
CNoNHXNGkSnRbii2c+An9Cxmwafr7GlMqVrw3cwbyY8ivj8SvHAmQ2MuNhZAgkZXVa7rhVQzs0Dc
+HEgzQHHUxwHBFCp/q6MtMpWNfbIzkZdx2tgFBffUVk1Q+u3bmlXgoRnoKgCZ5+3s6tfvQnsmtTi
blh188yfRyUNyVQz46VHCNsmScl2aIuQBZWVzVairQZHvCkfp7KbRtr+tBKOtj0SaM34uESZrNo2
hj8aGL5Y+piMpceVsIYqyc8h1/jFRUD6m4yJMrpcnLc+/XNKDTwzagKr69EezXejDH2k9zxCSWZA
t+MTE2/abIAF70BA7ZbQFGcKA2wzvbsiAj/9/VEZEuzoT6DvtzGzQwB8jlwMt/j8OOEOdMLo+M7u
Cy3vuuRnZFhgx6c1H5XRiRrJp3bF/4LY6o6jJUkJPKcqJJyHFcO+C/NFmZYjPL4Ab1GR4KEx+oYO
3rSHy0j8ei1zN3jx0/2hko+f5vULQfbuinYrWj/PYroWOm01r6NNUJnh8H4VVqPI9mMiHL1fypGq
+UPlqlJR6VTT6IhTSk7NPee074ORxrqjsLkW2jdw2XuKMQ5bvUDE04q2Q8fDRce9TQcgqYKdAHt4
7VtXOg8LBAELZAPMIO7cdSGtPej2fJcXtIEBujCDdLWNyOfNhPSRtv/wF+Msi07ofL9e0ihZ2uXw
HwqfzGeD4uGWYVUKplw7yP8zYdIiBfV9EAfuBfipsgT0CyjBeieLq8BbjHt4bw6wiphlOR5dUSJO
Ujhr/KJ2of/DSB96U0sDg+2UsHqwGP2DoxaaDRC7den3jcAIv+mVO8Tb6Xkn7VVSmIvlsEhC6yvN
oqXOfGaY/RfvI8u+lJ2NPeokqpDrR5HHYcXNOXm6p+BJWJAPk+SWdsm2iDPmdiRvXmOshwGokt53
X8FBastrw7MQsv96vU1Cc99lXe/P/idngIZRxfIv8Iem6mZLLCfC0HVkey97885OLVNT4JllTXKJ
bsiHZMpdcUBfQ33ceeiKJJ1spki4JZZ05SFt+TmVU3kQtP0Sq0pXUIsMP2jJXCH2lMy7e7OQyFRp
HaQjQ2gvdkIm8/BnuC32UTctqVmFbWeVcAZ+5beubUsoj6j0NhVy6SvTxRw28MeCF3iv8Tz4L3MI
v/dyTbSf0BGLtTx8O+oLQroxrZgEwLkariGdMe6vwd+D0Lld8aCmdupcLFhfxYL/O2moMqKNSfsq
PpmnuxZegEUpVDFpVQd5BHQ1U3hx6GUfkSZgXnBRdjdPO5QuPckf6rP7G01HHjC/8WhyxF/5D1F7
HfT7vDMaiSK9gYPmAYMZYRSf/n5+ye7mS34DuYS/ZODhrS7nLrIySTxw2J/uTRL4ep5miwG10BUC
RTpEGAPQbyAXHMwm3mVTmrx76UX7zbpixgx3wo5QdDz3qp6xtg1wLZNw7Ze9c97S9QAKhbQzD/Uf
HgCrSOrMKT9hH6o7UllNR11eWYh74+tG50uEUBka6QeVy8+BN3iwOz0c9u2t2K1Yt2IRTEj7IlJj
0MNNQWr4Ai7QRXUtsGlh5w2mgg3W2rVjK4Jsj9fHyitIHXVpwMD22u8/zhcGIxhQ0eZBZsauiWWq
WhE1gyutNz+lFYFDrnMftqKCW9mYPnPptCW0rn9Zkl8Vh/YSvvvflR+YrgOquaO+T3yKQIGC+tzc
SXdxSCW9+Fz4mWY5loXRwuVGGURKOwcM46VsBc7oEoFRCGV3qLe26QXVSoDE2U2pvzxHugjAzm5s
l4YFJFqkatdhW3DlLzLxpuME+oSCJsk1YoI38hbfaSrVaFza5RtQh7nWmnGgZX6t0ZYbT5lYwlnm
4rvaeGcJPHGYbE+yD2R7SWoo30U7lONOk8nDN3vFzlzYp1Q5h1+QWTnzYs6eBHnUaGS1LstJ/8Q6
+oPuSJR2LypmRqrdoHA/mhlKdnmYWgKux3irOzsMfUd4o6HXPhjJ+32mvlc6y+mTEHkI9amfRbD+
R1TiXR5b+ACgw9PNZ2JVYs4AatPO32OtKNx19q0uBP4v5ECejacFOby8+w1Vvc4yI36ev6751/tI
UvyanWcUZ2L1O3UW40P0O75jMOuXlTMjtOrr3T7A5Umlc4+HRJOMfjo1o3eh6FtX8WeCD78yCojG
TvBvQcndfOFHLVIcRBYpWWLQiypkIF1L0RpOr11GdBeTqcGditW9THOpO/1aTpcHUnuf8VCAvAeM
2R8DAEy/aOpA4+m7s5BttPdFs0mn6qJDtnmzZO/lqrptoMZs3ptt/+vIA0hQoAMpKK9DJjooykLD
8I5gWBhIDQpVfeDqK/jnoep3nEsBg4kCxBRokwwhDAp1XdXdxUDAfYs3Wx90PJognjgCoe3q4BnO
30NmucHOX//pOIHILB+Www3wn+27d32Iz+uOo3kFaaDBy6Eu8kNYpPPdmUO/IDVW4/kEwndxbPEB
zxRX2LMRR15PioCnb01DckFBT99kJnYimUJKK2lA2IMCW08d3OZF10G2bui4V90wXDbgArtM1RvM
wy6JGAlNLFyxy/zvcwKOzLxKJvfxqkpIknRQQrjy7z6ETt8U++Cs41MN1Q9Vti6kQ4Es2no+PUfx
wMi22HapVV+6opQyq8pAC06PSmBJ2OD6D2Uc2DB+6KdOIox+IMPsccM1WGF6EichDFpmm8wDNe8T
czgYUfil03nLD07Hg2IZbWu334zSnoruzutHtHXr5FCPlJW5k44lZAPX90/eE2OiQO/Dc21+Kr0b
YGAAm4qdMUoKmNbLTvlW8PQ/tPlXT2MmXPU9v6pF+9/d6fS7bHB6xba1ZXm2fFy3YDUSk/0XwcrP
5Rla+0Nq40MBUXHbDrH8gumI5yFwl1x5Wny1tqhHp+cuIRjKAgRiIT0vejgv9VFPXMPhg3eyER9Z
gGkJSjBHYEIBX1xt1k+XW+zpYJqdi4ifkjKOxR8NBfAXuzWOg+MPadWIKh8ZMt+wDXOb0GP9LYl5
7Z7VPltBefz3ljtNdRGumKNJn1bZs4g5BMge5W7eOaTWmVXg9VfwI/zCi522W2ld3+N+3PPEET0A
8PB+nnLpyj/7w2iGmMc+R7cBODinjUDRHxczoEJMEaAIlsdhHminMKH91uyzrkHX+qpeQAtSc1Es
gdc4Nx2loukXefRjuQSlV5nfbzJ4K84nt/DVqGtaovfYhaZu/sKPvpvzUIbzr+n/RXE6koZ7dVo+
Dq5yCfMTC4JtoluV4dz6t+Az7RmIV26+dJWdoZc8agawChL5jzygOqAQp2iLEWTMS2cK3LxYHgSh
HNSMRybNmVzwjJo/uHKWjzWIejhytxfN9zlcoOHysyyj2SqfQCzAxzpcqcDHf5zmQJRQTaEd0FEd
GWPfDezI5f79DJZxLkQvx4pWHOh8tZ5/4J6AfroVxy3TEBiYGXK+ntGRXyVvAGGLaNBoDtP/Z8in
Ze2eO7QRqtdtRlppYVZW8iyeE3GAPRNV/pjOOq1+rmfVzrDG8m2DO+tCY4aCP7Og0CtEoZqwuOWJ
4QCX9ssFkD9/YYKpV/AcEDJmsXQDyW0DBEP+MAC1r/lVK7ypm/KaRXej+15BtkAcwOfNST1STD7f
eETxUBd8i7cf/1xSSFPuVaSZuEQPEQwWjZ6uGwgQupZcj6t0Q2nN7j/ohEBxRrHVfhUz+oVCGUux
MEmlDIbLhm9WsuyF1+qXVgCDXE9I/Resgj8L/0ldqptUQFmrxBohM962Y8To4tPu6iKWha071VCc
TDDhljQDnovLJ/OYJ+SEbsP6vo2BbFkTezB1URN/9YkJszVokjle6RnK8S6IouRi/jF9IkmPEPTE
83gBszG8wnuQjz5MAJMqGmSc2g9xH6zUN2F7IbOsyQeL1KA3Vi4wM0o6Nh2urOLY2l2VvW8SmGWL
1pNtiO8Lr7tkuIEkdiE9IHf7stGGvIEULK9iQRiLoYLlJpXJRxaa+n40ft1voUV0O79sAzL9kWIE
cb7BM7eyDxROPM5m7zgr1GEKpUelXPY/5LxPNSdJI4BQ/zCam3fWBEKsx/1wu/jizrszaz1gKJUp
0wRw++OcZl2gw1YaGS3YZ7xb91GXEQe6C1x/AN3EB09CqLpYOwPz//ng3DS96VXUcjnd7SnQ2y6O
2d2ix5fcp51KR2FZ/nPl5a+Kl3M3f1KONHNbuPVcLwOzfmUuqqBLJgu3yyAxJ7OmeHa1nsFOIXQx
F0kgLTAX79ia2rko7ntBJC+fi4U+0HFTWgeiibAByI++y2D3IKPt8Obh0/oPrwTlMRToJ32FJiS6
q08dMKKq/wfnc66gWkhasEvXF9dL0OrG7TPEhD6Sen5MNkAWb2yfkGoOoHvoqe3MM7F24vTqRDmn
CZ/FR3c+E2pPreJTHXvLowVi4cepqpMMSymfNnzdVd3D4cpx/q8Gr5AQSsxWC8sUti4qKrDdIz5v
RgqsSNRs7OQ2e9WcOpc/x54NhwlFklW4uqTkYB7tgaKYaL0DgQosA0UOow5kQfZn57/5Rm2pnCFG
j1nwnjwiWr4/0Csjl0ea8a56Nfe+SIey1sL6C3Bz1906SQ1jBgvXmzv/COesTdo8xCnYQQHsTppG
Ic+NcB3T7GtHed1+d3LKKPMkLWo5w7ljiXENDwIqFRk6id7JvuuS3/E9ZjuiEZXPKfaMp+Kj2ayC
JcGS+fLTKaCuSTbMyUHc9YbjxZWTcsznx8cD20GVKiFcG02H5Nunadk+gJWlpjjiwWsijrafyzjp
hLmsQH6t4CnJgfpqDjErp6dbgLA/PAobFu5zXp3wkXs8qlF6r7nIuTk/9DjFWDcO7MysRtFXq/th
WMxQUVpiW0SNLc90u7FjtVApo2nrMAA1VRUVl+X1s95kqwzVnrA9Oe3AuXhmdHz3jhPDPwIZnKEL
36Sxf5gjzJNM7beoWJ8798176gsmte7dNBI/rFJAwA+VGQj39GSX9GeK35H3gj15tlFbI0KGreUn
GYr1RzgNoH6cCOy2VPILKBWPY6QSXz4zpfSqUPsjRWxLaVms624Xird22PWV6B+EWPkEER2cPaTI
MWGRCzhCcTIDrM9oSuSeKuATnQy3BLWuwtQTioPEWm107qXuawtxk+gbuQAaRb14n0dr3D/TjnnL
J1sgOLpGzV9pzhVP+9Xn9cgQlsB5nZJjk8lFxz7n/ha4teIsAGWyB6TGfEaR9OqWRLZ8YWFNAr+Z
6NhoAI+Db6h7GuaHLO1OueB1OmsU3cIdiR7WR0QpZjhzL3Hp6lgrhGRYh3poFkVh/C8GTeMdBjh2
7tiiPxAZWd/H8bAmf7JaO2uwWng4Y9PZjSzt0UshlJ5H+qqGUrC0DBBGTGjFubKm5YMCddfmzrvg
iA2tzMTyaK+MW47D0gk+Ly2r/psSaXIjJEK3e/zC7xprP49Fn/X34vely/DsYTTbKglcPkCRPKdl
I54LpuZslKwuT/14h4aZpsAp8C9yuLSJ87rb6yUQI7Y2ctffJnLAf2X8Mc17T1+Ws8yvvge3pDw2
1MSla3sG8bGH7l9XAPfH0koqCUsrm1bf/cjBKRu1HXvC4hRcUH3oxx3lry2GYHAT9KGklZGjenn9
y0lG98FaTwBO1UY1hlXTTyebs/3BxiRUVcSdIa4vGT0HLTxMTP8rjpR1dQ150dmkyYbgOgstZcmh
x5LNHIE7GgjMUrowPQD0gCjGYOnDbE/PxtgMAPiyfnPmSNTfeiO88i7fBsX6iHCll+VOIztV4lth
g95ir9eTA+bgRoIW8IAk/I8+mpLQjlOoXWxqIdQz5MMr7ZRNtNH53a+WEZaaESQhjSVsG8HW5VnA
l/ZsJ3MeKZsjnAnink9lqGYiSfProo7MrsRA7NkHJON3FDPE03T5aNfX2XUgVWU5ALppRkBD/rDx
6JVSlENgdxNUW6BeOSaljvt9cjnR3BVoc2RUaaXzXWt+QmsK87wzqvueRdYUUU/Embi5tBUk9KZ3
pcBJHlD3gSUrKclWwTV5YMZc/7m0GbYlIidtVXFpsb/tQm+nHPl6Vr7gUNp87owo8JMIemyTXOei
VBqmrmAppDwdnwg4pOiLhQ0pHJkbErVoow5zQ9qbWMDWEBuXd6PenajwgGHLfX1Lr+DG1ei3bjJ9
fGgSj2+NezTHVJbLp/Hu+M9dhRFmEETANoOChAtKfevnlMOKi+1C6BZGc17Tf4J9o0GBdjyzI2iL
7xedSKJYAuApy8CbUc7sMrZ4X6PEaB72F9Rl+wMNjGU057w4P6dKGhOgghMTCLJRVWkthTXcGzbj
VMdM9K7artkHjyPYRWLcJU7cSxOayBBF0ksqrwERT7R5g8FgI7IyMghXc+xqdrZZ3iCT79ZywMDH
BtPfEA0u287V61twTIs+lMkKBfjmogvDausnhFTSos6YtWXntG13RH/GlEObbsYN5iGPowuy91NQ
VIcvxip7M7zDTzlS9Wrok7e9ziLjTkTzBk2Wzjpn2hr9C0QsLA4cjvLyJ5xC8CQOeS9JKULZNd5Z
7B4ujmlIiAMRIWDmjw7r/O9N3h0A5NIl9upnIbwlyY+KkfbX61Kvuo5yzhBV5bNducvx6a4X1vnk
jia88RkvLcq4Fsxr5f1WXxQKJgkyVc/OrLQw/+lY+9GFkM/mwfdBVCDQb2VZUQ2rnsPotyJqcvGy
XWW7hiGZQ+P0tj/Zy22lykFZLkeI1TBgjh/MZpFeuFX3YgtS6EQy7ECIcOtdbH27qg80qU/DjyNK
dVQHiTBUQFL+FsgAOhWDt+h6RvMoUHrknfTSQKyaLWfew+GU7G/UlvGXoUDW8qNv/B8lK/rUYKA/
bC3bLwACWv7aLNixSJfrbYhC70nqDaetlIZTAeDBu8ZLhBl18mJNCotLtHAemfdvMvrQu5Yj81A1
kiB64qwnBItlz6wBQEfWsYPUROOpRc6DMe5f4c+6xEfPOe+PJ4hmYxucVj83Mibl8gPSKkhewP8a
5VcBRJ9aLsWyyiaI6Y4PC8Bg5NYtQ+koSLYBmGd7IU8TTfkrVYPTqr3Xzx/uo7noLN6KWdJ30J7x
O+skLXYvmImMsOtRR0vi04Ivl5TjmRRVZTgDhj2PtW7+Vu0pSOqRRw/tfThddFSdNHVIikeJmOox
VY6ne4h/fdPpTJUNxJjMzNMwNJh2UIArWyo54sLH7CXBvv5PSt8jVqUOnJxJhp4yGc9r3fkMwWNT
7SVYvBA+DiX9jICGz5LI2U0YkJ+lrzV88kAjxMIn9A2P/t+82P6QR3N80k4YVaLXZ5vrt1+kXH4O
hAU5EssJGecUB5O2FGXnlXz7wJVsH0xOfO4ZnPI81nnlFaiEMeWHPKspUZ81xvNSZUMV7dK8HO2K
8k8B8lnBidrYX/CeTS0WiUFH7IG4vwyFNIvq9F7Q7B+YOaZwMZaB/sVyfG0blK4NC5KxOD7EvXuh
m0T2XVRicRtmC/zOQQ7MmQLEl2mddsyFQT12xEn9MJVYZrwj5901jRdxxhtl1Lb+xnMr5ceQmPbj
7hMGoUiSmy5JOPnsACPDD9l7W/ynCDrJqj8QFwjW10Catv/0U3YJbT8+J8dl13uKjEWCbxWv9oxU
a+5zahIsvAvIcasDks1KAqRhlZEXI0I2/fzmrDsRFj0haWIDu86N8sjZUPV6b3OoKwRdLhOPgEoI
YvIKXRDlhwcV73p04Qb95Izjbum/r6txX1KjxMPCdw+9kQsJHR4F6r9nFecErdAJZ4j5tfbJ282s
2/ILaSYDdFMDLccc7HVhonETaEP8IR4xMVwdkkyTKjYZ+k1XnyjTEr+7pOTfh0iusWUU6btXpXpr
VBsY4Rqk4eAJ+dgpNZfyZb1M7u//b3QIuo708lakdAVsOyRU5Qh8IKzyDY2GYn8GtYPX/dqMfG4Q
ZM75MPCICIetcm9w51YqrkL/O1YT0A70zqZqHgknKldVrXdlHqiuxntJNFzlOnn2ILduIDbwL54k
re9P4RJPHHumymQnyXQBfqMKLr5xZvqKUjr2JjRiuBTLrt7Ck8onxT6a5qeR2afmM/yqDEcDWjeY
hpPkedgi660+dfq0PQeD0lZAcRQfZvTxnUZNINIZEbTx8qp2FqxW/x6/WNGC8XvrbWVGGPBO/E57
5+kod/8NVpXLE7TSU4xn8XJAZkF47yRQ3Dkk9jx1VKmonaPUEP26KFN0KL1qtD0BUBS8oq7Ycpk4
u5UTZasb2wcOffQKdIEvkTb5qFTThJdHbSHkptqsohON+SV9qvkv5CvNTBQMJqQi+6OTKPQ7grCr
HyEvA5uWX6pA1McPoRy2fqORgAwHhWu5MQWXyDPmVxT5cT4MH8ZNbsw4V5jgWERKPFn9mfiGRO5h
O3vW3NqWAH2H2l8Fo5Wma7r0/cjIzZSIk1Gjial8yP854IN7NfeIP/hoAeq7/nuq1xPEwk3rlSei
cHn1jvhP3LgSD4BsY0ziU01JLbh1jo+NKwaMdkSunrrApVMUQjM4VRZTNL2j+xgd4gUL5ukfcwCX
1KsW4TSE2WEPqc+0tL3lBVbgXFgRA+o6IKrJQ5TWCIzvEm34V2peLqOgUu2JwXpdASlBd1o0qY1Y
FSaFTIJ6dX4u4Sxgq2weqCbC7N/ruorpvA4Do/En58gNlUmqeAoKaJ/9iElvfu9taoGntDaE4aIQ
dBHKSmr4edwD3rw5fqcYWN4H//eXbAYWzaP8w20Mk+qsDBmCD3RIEWu7IhyKsMga6WxIVSq8wypg
z6aWZY2RjrktKplr3XWDXS4VCfEIGGG54xfh7ynno5JmuvLlkgdwsPkeyNSJ3myOhgsq+kwg/MDX
kmlreraFUp3gYgNQwZA5tYYT0VseuGGxmOCcFy2HBXQD+1d3Xm1cZAuPWBPuJysXEwoCA+s+xUKM
pJN2neWwd0lUN5gbkvNuPDWnfLm7zVU8UVLNkHmsqBm8RxVCeXGkxIfsRtfwzvgOyHaMOh/LFIZ8
JWsGBEwIoeXeNfvP6ffp0H4JsiBARdLVUCctKpuR1keW7eAuILhkcS2CS6psdX0Krf6r/+klYcbK
W64p+pq5hPBr27o8DBxh7t2rBm3Mg/Dw7FR+xiwgXw1/IZRfPI/pSIvbTHG1ThX4jIiJn+VukIg+
OnEOs+92I9p+Z6ar35IaBIdKSm++4sHitF0ZpHSQN1v+eOJC3ohNDr5sjrpK2/BsLccT0azDvq5l
/X3Yrzks8dsQqyyXEvfqaWSkMYv1HKGPaS65ZmN7d/Jtqs7B2h+OgR0vSi3ZOYqJwyX7QICctuUN
FfihxrhHM2tgN+sGnWW/VnpTzFoWS7MaWNzDyLehvukfHrgVFkbNCpIiKEqXUgH1sq2Deqbz9g1w
7qNBhLn06gKSKUhdYkBqAmsyS21bTln76Wvxu7MKvgW/J/6rzG1K9omP7bM0OZs/l87LM3n6ocim
bi3oR8Aiu0hLLkMZm/zURJr4TAP4kz3w1P/rxMQme2BbEJ6H6LUwGDEWuNDf5Aoy8v1PgcDn6dp+
7YGHd57yB5o0JlP+/4wweNcEr+oc1MEsHR52kZ2DeCBHglEJAOf/FkAX2VczQlagWNX/4sUxzLLn
uyPcB7Io/FO1/6bg9HKrnSG31tGxauYPmSI78YcqK90TsFKqd0thJ14aR0IsHaY/SA+aI1+NzPsM
4f9Y5r7nV5Vy3byWS9935SPsBF39WOO8WZxw6oCIrlzOz5MuKH+dT3pv3fP3On9d931ltRxrMeAE
r9BMieIBoDs2ztOPOCUeiQFjLiuL6EGJE8OtE1Re+dXuSDUW7/5zsTxaWVwSzGy91nDTrv7sY0Aj
mA3MPQbvSMi8HKgJumlEIaRemX52AUbjmacxbVbW6qN14XN1uBBegGpcyo3N+Ht0AgUEJFW42V5Z
lKVYHjLkimDtOjCAHPXDBmU/UYidrkAzuTbyKyGBOIm6QXHUv5+SnrncBZAq/9Oss0+sbuKT5GYR
0gtiPJSt2lnlBsYgr9cYC8hJlt8xd7uNPZp4dLcehhyKucidzpGASlQkCG3i7FuduPepLAc/G2Lz
0pZ1no3riEZ/a+UMHInvGYsxZNLqbdPR4KqxNyv5G5omtA9eFP3Y4c/TuMY0DwANTAqzTmeRsLbZ
BetlMnmVdBWmtNJ0BMbPFikyGn3JBZkpPXEbX+uNRBCHHSSDVqwS+/zpnB9jriMhOOPPX90Yo8gq
54AfFtCLbSGaGVRERj77KSU43JOjRc4zWj7tBwLIBgsMsgAHgj/hF3/r+uirbXQIVWU6uLIHFL4k
u/SLe0uKAoqAEimmUC8ImiKbzqc7icDjo9zZTj4/M62YjORQiv28KAOImtLtEyHkJ//36FlCqVsP
d4Ue4AFlghqE/hrEdEF88Tja4CKUwO/aH2McPozS5CMc4SHvq8yzKumdlR20FzIcWxTgrMfnAoKQ
bO7dxTssSMgJ+gLdQvGQvjuXj4dW14GcByuw0SUNrhqdeTe7IBlbMdSOAw0dtGdus1teEVc7uzXk
+gOmKfs2YjGt04sA1U6Nz0NUlhBKxmFdCziHQf7Gd8xj/TVc/TNCYUeDevat/sRKEco4ZYVqusA1
0tlwPBWiRMJ0HqoLvVh+76MuBvUsAHuH6mFO0Fe5yfD2ar8f+lGYK9347KiXFLeMGOR3leDwIkYa
qzex8j8j7EG13nGSYQj8WSZD0osmyuzWywJrf+m0lOifQiHmPSDRPkkhhv1/oweMlza9ZrgcOH33
48DGX8Xw7ZCPDCXWztdK0qO1UvI7glq4XjXx6m2EeZMXXVsZuPpPWv8C6uPb1GKCZYF73LUh424N
Ktwgwzdk8TG/08FXaNW82+MCz2LmEDCxtgr6Kt4LN87kvno4ZHKn9/5cFdahCBlu0dCK/bYgCEQ3
4xcnK6mXrCUM1RMUTm3YK5bwm+LF6ZsUp+5xsLVrXq5r+tpAbghl5j3ZOvFFqXi6BR6iAX18fcr3
BsIrmD2o8inT50o1ufwPgAbII98b3YJGaUuQSlcgPKnCpbuAkbiHhwMF7UM0VNx1IMcFHjYVhqPO
0VNT9HA0BIj29gPCrjs/Ux3c6f9AeOz0oFH9j/uzTa/inNALNMTbZf8HiR9dAc115eBanajCyVu7
h56OneZsN2EBMcn8mPpoN7jM5pc4k38Ds8VRkyaZcBYA6UxX89AZUob6r4fq03GPiu2rHdp58obT
KVZltMXnTOc3YlpZSAOAgP1+f2b8TCxTwXywknOlmxBgHcA7thLIAb+9IaaUE+SFwn4U+6uttTdN
RSr8kqjjKVtBgBMtwc3aEw6raE/ba/bns8y/uDqnreEzb44TobUDxuMP0XVrA4B7+qfnJlvxmOye
JXp8U9vb8Yuq9zw/lk8LhC5E35cCq+95NP714GTY3RjLqu/suEpZbAirwc4NYUye+HQol8GBW+Ts
y29VnercQiB4AD8X9PgOV/+AA6hB+KRJX0U1DuDnHmmeFA+Z6IhwBr8UKjMV6eA09cxnjsEl4jxP
fEEDhP6602FEjU/3oHFyxIYPbC4+jpULNLX/1mqWMwKSPYKk1KEIA+Q2bymGF1ipWf2l4bnUusyA
r4uOgr6C+r7T56N3LDRtu7LFy7Nu4Os0vWxO36O0FkGUQ0FWX+cMMaINmgubH9cUMp2+MyWmgJBO
go2r/6dRWKeFNFKhnf8A8hUOyLh66RXnNvNph3GsqIJbSkg3LPBHxnrfKjkXo1ov1Hg0nkuibZsz
JFu8EvEAvS0/3LwxBBXko9SbvvinX+gEbvseJOydyL79dgvYZc2WsE+zP6euCjdaDqarG+WdWDi6
cWeAFgTLU+43vUB9pE6o6t1VhDLAEONmuiujstyqhXXiC8PACM04Nrt/6JM+KkRfLjDw6Tah5CBn
wj33JuVqtK+WxUddl5LZJOE9c/T3JxVi7G5WVck4FKh7ewzintwJlIQO/hFisM4EFsbZnVPXioL2
NA1taDntTTrxEjUC4TQ1GJ7wqBkgU7XDuY01L+7p2KsaCywKX2LHlvukdsL9jaGJobvPIgXkdLEF
6OAO8yz5gt3OWMmeM0A9Mp9NLlXkFc3JWJyazRg+4LbXAr8PeKwefy3MG8NmfATlLka1RToKD6zu
4mAug1MD9zTfZXj+COQU9XQqCt1xFYZWP3nf+HQpQYqhWgz8wxxmLve9ff7bw6vx4DY73X0ZAELA
1BQRXM28UAO4uwVCj4QEuFrD6tayZHfoVWPLP+VuGIe9QH3swB+kDxoJkpDmydW3dB3+fDspRKyb
ILN58/ppGSMUzSvVzbjdgSAgGnaOy04E8uPJo7IC2gazgnH6aSdn7NYW4N2828zjegxUBR7iFw6G
Q7EQ4cqFJCZalEOopSn8b/+lKCJthV+GSiSHgyZUNx84ks4ZSUtGB+anv5KrC+mphKbtbgRHZ4+N
0LDmSDqe84HQEeVNCR37JhP0kHIv4IM80NwNLlyOCn62YJ3km2H0z/oiFJbLa+1lhB0BolFoKuFJ
Lxp+777BLTJOAchWuIKfi14dCmSqJk88KG5JSHUjzUARoKWVa+XsQEPFurkpwFYg5Io56cGyAkB1
z6mwTkQf05/PQ0VZSlYuaXPGuqW1e0e4xag6KUAMn8JfunEUpabiJ6fDiMrJ9O6VkNJ4j8pcs5Sy
l8gHNOYg5M20LjcI88Vy1LC3EfIWFrRrYtX5p/qvpDnCDJUcUogEBOEXfecirX3aFpl/fYZoN+G3
bpyAFlvvmKy08PuhbL/scViJHic8keR7LdbAYHhYj0pPtho7G4RUjV/q7Uc2AtV2RwEagzTK4uMu
Z5vXaUD5o1dZ5TTO7Z5xC5i532q329PT2hTtj9p5Wiucnj4w1WMmP+CljfsOKJOzRtt+CookNRIz
6I4h8jaVMdu8uzxSTx+4YQADkCkD5a/0DXwpBrn2pyrtx8LvZRLskPxo8SZsPM4ExSxAsLBeRZLk
3dnyUqJlFGwk+jfGOAOqWW8h/DqSCE65OUyIUFpOoItHRx1yNFq6jM3LWq3go8+dLiNiQ4uEvvmU
xJ3TKAIznpa1F9Khc5BmsJ5FG+DO8nbRjJJ6KcsxtUGtBPkxhrXsNmOPKdsdLZHDw0q1QZG+U2fQ
cpBDosncsazkEcd9go9bevMw+0d7Xakypao6nIFLnAWbaIJP/b6uNWdjMt6tYhZJ8PFqBjeXOOut
YDnxvj1Izj6m7Szn8aQ83zaLCSzBjqA0N8lJcm3iJWc8sBWD+kmfAUwhrb5nTIg4hxRtT8nVJv6/
VegbLRkRDieHgt4n5HGN+17HaO9qPjtDuiw14SKJ1BBR+sdj8jHawgNsXSCbt4hlHrwlKtsNo7AQ
jOlHqn2vxPe82lQ/ktnBc9kBMFgUBF1tn22TR5iY+Z2HkNGF8EafqnJJ+TKPOHIfQ2ab6hOxAduW
pFsOAc4pR8bVplZXQ3j6IuX4VwFaEGnlAs6IDKSM21D5D7xa+3+AeJ7+Wkt2ZuO6cUcszfg18ybo
83JuoEaJNky4Kar4VZcqfdOIgo0Qo8tzGp+kb9SSILZR2cfaApfnjKgyIEP/GhR14t5rGG8mmRkz
ZpOS46O1tFsaHuSDw62R0HBJY7+mexhnF+tIDNu5DGMXkZqJl15JDgMohVuqeP9PNK49Ons+j8SN
U/oQgQ/JSxtdTcMYQgBbvIi1q9fI4tHqJHSc35iHK3r1w3+jDLJMjwi3ccCJu7YdrroQ4Xq+U1NW
xx0+rQrXMVrTdnUyE1fALMDXrJF+CcFvUDd6mUpYeMM0XS+RPZEAEixRk8cZMJUTMjgvMT2jwpCW
2UR9PL0lWk7ePtboD6WtIW5z3B4kk1ru2EbEcYzJLOppyviGibzEtL69lQQH93HhgzjqF7Mrjjqs
/n++PdnFxrUmqAUOm2MaTO75s+h+iudZOP8opfml4QrTw2gl9iYEeQT2qddtsI0Gol3sTW/czAIS
45wHSumnfPRd9MTCE+ysVDHPcFFfiMDVcRhZLfi5xSwoOd1BgXCRDgkJSn/5gr5i+/7l3YShMqNF
JTB+QofsaEDCSocCf8QxdHjZfhUrYOXUFXzDzjcRFYFTQPmuLf5gj3G6tPPy1P64UOOLKaOsa2I3
UxL75vGRB2MPq6ch0JcPnjYlR4WNeovk+FrflOenPfEmMYV+HX77VNIjYZka4VmIKBnGTyF77pKJ
UVXqrRATtYQgsFkzV1xyfCifhLWs7Wy1eMS2x/sqjSTfRev83NIdqlkyKYyDJll09CgteuoICMPg
i1S7adq8GGLtac6S5vwGnEVNNeLlPbzGS0Od4QXxnh4ZjWJs4GX2Nc+tgfpNmKUq9dFU9Vh6VFeO
W3JHVRMRTtS5VrSyfn/2XjxgDP///ujjVtCEWt0+IbgwEQurf4m3AR+RhvQ4jE0tDBhfOAgDjGLD
uikDL7jN6jqPgYVqOLE42FzenTrRlkgOakArUSyB32Bf7nRfnhS+3FnjbVGpzpFraMSY+jSj+CRQ
yZ0PIW+efxBhc2DinWxrZqlLPriIb3ISt023w1rCvGcy4C9LdGbOzwmxC7WV+Is75n4R12ea5QTM
pp5cFxszSKZpf/gnbxd6jYYgD0VNs33cfWNLibPcOS+5vh+3B9EN6ZURKz/XrPLiMolI0Qd12OFW
mfHOBN5oYQKrg391JcQre6kaaXpZW7NgrqI70Br6doHw+qPqBGkOYp9NFP7LtThNGkkO07FU2OBo
J3rmIqbMB5ItHJ4Hy9T4ZtyS8JJCvKjrN+ozpMKY5a9V++vPp89vqyRgvU4IEyaKHKXCjtIamjRl
4xFz4zoiqsN1n2fNLJI9KYoMbnuqK3RmImOmIFzm3LTZdnGuZsHrysV0HVP0Dl/yWquier/sWM3o
59/ou3PlWDzzzbKDaTwM4MTgTJbOZp9yyV7k2EDpxxRT1GJAEcDat0bTLIPgonUH/f3po4eK3caR
OL14fz67p/6c2vhRiZTUjvomo+PlIbXP7Jg9Rf4X63LOi0slUzzzWiXlDCEQhJcTebdxd19ymqD+
lzj10f518J4rGxMBRfuOgqzpiAB+Qj60c0vifp7SJrl+GU5DPQRmT6hzLAAf0PdGPPN4GEc1ujEX
hndmZSjyi47FhRUMp9WFr70otRA0R9IF91TPBfvy5jFEfC08qFKbozWP2bMjhfPGrFOWlOFcexU8
wg9m2F0HVeeA2tfc8EYbKEPJQE+TMfeoEJawYQv5Y76AufyIo6FGVOqrH36Iq7j9dBb/wkTmdIoB
Q8id3RCXbgkCw/OsU1fFRSOwmykvqk99RMDR3Jf/5z+7Bjz1GwGks/ZYw6jrFts8oiD4nWTFw9u4
w/XPSXdSdFFXaHdWmzAo7839wBgNcL/YEC78d0vzAHOGk8WY2oO+0ULVsmB1H8yq3EgSBtRR1BQv
DCQ20n3Dx553MuyCzIK3p7QiOgAYOiAgSJV4Ivk5eBzhpA8y9k8dduiXY54bHG7HplBe37d+eLBS
81cuTHHNvWn6io8YOlJXpCEyQj5WzlqOP9Ox+TsD+yA/inmJN3EVPvugff5h44Wv8vHiA0IDu0m6
/oFq1bWJx8aD73GfjGGAYSOgOfT+a9KTeZEKrkWnr1qntEUxZlDesbvZ1vB0DtmU6175jlScaG3y
Pm4tEJ2VP5noVOcIarfNZgG1oj2RIz81ocgzhj685mGMhjhDQMd9lwwSIpZHh0fOeKZcPlWozxms
JllKRfx+uKbGlbq+tjsmmArQ1t4czIblfxAFbJ7QH3dSBs4oYSMonIV7wtiOkDPIRCDghlfnziWe
foEzyURPUOJVHACLeNp5GQUvbJCHYvlqxAP2TVIv6IB75P0M171zoXlnLJLU1ESFRK61OiWNWVK5
4mlGzgnYkja2VNqQx5NN8jDXcdmwyYvlKH2awk35VnWV+MDzO09RAh4SNezprSsHz51q93lq3RXj
isD5L2+IzOTdqcO26pVKxbh79OBZbCERW/B/L2D2+RDNw6+pb+f5RjJMvp8wprm25zUznmVyTYE3
XgqzLRAWYNw75KAGOICsLouwTsamCEClVdk/dirg4t+bC+9SjEvFd4ze2D9Az20wjDu3Ioy2DZrQ
4UBAxt8VLXkpLVGavwhqpTJJQKuDRN0GPxfnJPVYi4hsx08GHME+7HeoHn3tF+RLubeDblquuIYl
dRnXmzG/PZgUg799rh35NNmoz0ozsnmEmTLXS/kdqfnOxy46+5UwwxuDATGNUWmLd+QJR5JOKsYk
tvEwLRhhJRtRD5i8Zl8wWNYS6O9cj8TmWwW3foMkrfvQjWCQxy1t+j/S8jGkUEwh45twGzG//xVZ
xrTleKdcoWVdBdrjDWn1CQYbYU7p5JGhhSe5jmQUxYGreRz9NlebWmM7+aOYNQt7h1BEOZvqXw3J
ecz5+8C1J32Ed1cSp/7FT31fv9VqlPGN94Y5UQmRl45wFc0XV8kKCOhoPUkIHQQxTIVUSdY0bdxu
VoOyvaliLZuYYuhFwJduag8XqiFhp3GV3YjF3Jlnu84zUIFEp+63kH6XlBCF/cGUrA2RYQ9ijN+m
Wsb39fRXKfaDAB3O3xBiBPuHbYMSeE+LhHPPI553VZnmlGuU62wdZGa03osjlQHGf6wkZR3AZgWv
m/IjtlIhC/OSCgTXrgv6kM3RiDSuzTRksjigsIXM2zFr+UqW40DlqcGNnZGUMZV3tPn/TZ7lRy/G
ABJ8HL3OJlcoeinEwK6ODAdL8kl9VGzLLa4GWVrsoF9nQJ7PeEQXfJ7oXwmYYfTHiaS59m0PHNmy
Je+r8eWw/G6stifjPPH8AOnWPDY3e3gHK3Cu8TaQwpfaFH8ggihpvTFVq9VAUePsaTBzUUWANqOn
M/SjhQgAk+59+Z6nMngBKe2CLaEgFf/5XcAppqBvD1aygfZ68DSYbHtvNs71ArtuIAdMcbxkQ2lC
aKeP7D9DmU7VzRbiz5rOeKg7Yql5SAWaM8b3ue9YOoO/SyYPbu/qjfj5hvYcmygND4jGWYzPSPd3
LUHefzqhJeBseWZvxMDpkHQOHEZQr8fcxhGkmseRI5+KVtFLUq2QOb2CDuFkIGMg+TWAUPsz/ibe
34HzrXczaB0n2KpX54HXFLFs+X1KBcsyziZBF9Xwv2kg4TFXaxWIXY9WWulEOkZRnYlcP8litsoL
pRNxgdIrY/NZtWGyQJbGi7KWLHUG/CWkOKKa3BlwSW1lImPaefx/Tsi0AtbsXdTobqJVNEbfqAyD
l4ADPRgb0510jqRmNxG3KRUiIqmqdDZV81Bl3PVqqi1Z+t7yZHTLeeuqzLIBMgw4gtVnzYnf8/vU
9tBKIAgj4Ht4PiKJnIZQs/M9pxnodqL5OBoSK7LS3/ZRjTicM38EYCc+biUpZYZBbnX5GsXVVPeO
HVcZ3EkIAUf0RSopxtyhp8qcyyWUL3Oq8OfjMySz37S4F4b1p/gNgaRuI37KdmDqx0bmjggxEDGO
WacikU6oW4A2qhzyb8fqIg0bZk6jI6Q+Q0u41rISGwmABxTDX9yA1bZ6In3ghKYPpqklXJLdu5/r
nfRA1yGuNNBwmh3Wm/KiGs8q+24qCzBOObIDz31iCmuLAgCN5v7xy+UqQ3h9kL76SaAfGXyfB0Dr
Pcoip9QqDFSJIABNaia6mytTB3MGfOcM0lIraQn4Nu/XIEfVtkoVyUJRVnS6f6hWIRVrpIOG5o0U
CfnZN4vIw7ZqQcbAvcz8XEzAO9F8Ujz8p5pz/bcU4vQpPml8u46K+iU/XEP8uUYR4CpQVmfP2bMg
Sz/E4QH0ofnRdn0gUSXH6XP9AcU7hQ/8i798GL1o8ZSLcZtkm8INyw614x4ELepsGorhonvLt3eh
r+EMiASTVvzFxt4zgZmOmiGOYIUy/ierDTKzhquVOu2qBL5PhMghs4OrMVvs0Da9YAdvAWkg21Pd
Irn36Fq5y4XjhSzQUqnIZR143Y4na2ZvwVEGRDL40L+zjLCqttl5MEgnlgCDAG0fBAf04rVzm1r+
eQHzVrJZ6OD9kdayvIV8ZPFkxtFpdnG5GMzyr4W+AQpmtGfSptwg3DBimbUHyvwTp0tmIa/upMON
ym5OojYvFr1wusJvyky5NjOSX/wcjJOQGsgrWT4zL8/369guqsCGbAMvfZ7kwr3sO21/QH8yfww/
D3sTyPZ/qV8jn+gz5JF8T77qH3aRh6M7TJDgbRm7VSd7Cpcy5b2ka85t7lZrGBSQJKTYMwCQmqlj
OOO3MqxQ80GzqkxxGXg8AAl74lhPGiIQtNs/s+djZVeJNnbuo4/tVLQh288JBB2EnINWcAjweo4H
fxcdopi0hG+Z1UZVwiZ7lG6jaqT1y6rIc3hGy+G/xzdxq9VS5Zif+SCv4m34czyWw/xL0EXlo7wj
DD7CmUo6GUuNDdB+IcSf2Sju2UobakvpuUDXGqhhQ4iw4zEK4LKzMU4y9oC6zKxclvNO2Lo2YYzB
AfR/wba+PlHpR3YJvhii2E3nbAHTEJXijWVsgpIL4j7CHnBAA10alXbSjJAxl/+kZXDu6aua1DeD
db90CYJHMQ2joo0tXQlekkepuojb7RDzVDp6sOEST5Wc1Ss0IARTT8XqCgDENeDDt4qpQ2RaqtR1
tJaFMT/Uwmvs3zzkjkriHt6LiMTkMiVIHXnJApZXDKwAfLVYxxU3o7ty1tW1c4zShnaWBenWSq1r
4icCMSJyUjeHdPIwo7zJoT1sKAFk4wvonMQUREAMs++qDEkSnlPDyeULUhUwzSYE/9AHD3unUxIM
Pm6ozINs9HixfJzacEJM4eVyVGfLg51MsvTG/vEtAJxT4SyQokc1ZlnqTbZ8OCk8X19+fxTaQhwS
05W/Rwi3DhTXXtT6aNNULVbA9hse3B/+XTVjhJL/+oqtpM3yZ9GPhS7Qb67bh4X9kuaJtCgooDdH
GsfWNuDAskMpp5GQpriEQuuyT+ifop1etQFuEuRi6jFdVEqx7YSBYOV1fGWvSMXr/ObEZayvbtee
POIu/oUekCr5YtQLGP0KqkHNzRzgbrw6NwSWrQ2+N45GUa8CSIMKPeeZBfWaHpLYamycVOXNQ6V1
lBSB+KhnMhebDFJSN2tAWii3Vhu3+rio513Oa5t9Mx/S+p5/ZmYpdIGA4nNx2NlOCwtUoT67fZk6
+9a5wW8LoubaFGL07pmQO53LQf8FCtSBBneWs6HD+39IuZrifLwznEfXKueH7Qs1ly1n77tbM0vA
jIcH4WGO2OaDvWYDd9P06uMMXJ0GeD1hjhW04kJrekxyX5oZjnSF8nzUeLO7QOwr4GK7Cxdbir6V
YiD6jCM6tcjNFE3t/pSLimxsHFpTbUFGDEWnICvy4cTYibD40Rnbv0bAFQVOX1qnVsBQybMoulPL
4hDAgq/ynqBCqb4YNGVEbtqH/PPe1vJOikQcGq7lqZLjorHjh5hfJLrtnR3YXJ1x0wLgRDa8Cjop
ObCjC6nw3dGR0OUXlDscUYLK8FvO5Ww6uUDNzMjs9iqzMPWJQNv0k054b9s70ZyUjw10lxipLXho
9/fVeRNeh9iWW0W5tM9jeMCYrYYHt3v9ONahidtZA88VbYL4uudcefxubHCI1UGn6Yfl1sbFQqn0
Cl8nYqyTldxSyFquDThoSWkIZAFdKFOnR/Sf7X9yCukePcxIkufr0iRHYa7sDXwcHc4tX1/WL/Mc
jpEJJ69GxGjs5NqD8r6uezwegSyOB8TgkcgZAJsr9jmDGshIGUo1do1uIpvv9u9M3pOBMir2MCxS
C+gczEFGbqOV85r7aNoe5L7VaUmr1PPS9Z6N+oXATKjzlnwelpoVjSGdhvIgDQ+TylJOHFm9ftAT
mB2jnyklEuxslmZ/MQRSvKMsFEsck/pjmc1950mA2w+iTK16pYsu7AqIsWC3iW/CnFQ+YOpo/qY+
vqtTp2CjLfVdhmjaAgEvfNJLR8eWYR6RTNHEzrwh8yITPUpgCKKTgvWxETlRZ4G9Whu28eVTCrOv
5OCyZxJmVIhAYlwx+2de2m2J4gWvtcOcW2qYkQ1sCRSm0+Gn6Hk7DMZxEug2cQjOgiWasB26c6G7
lg1sH6Svzwfa2hNdfaYc5c04HVpiwXw36IzcwwbBnJdSqoH3boZ1zIpsT2Z3IA5LDujkp6UBkUXx
PvZhaI15rYke/7ft5c5prMqPjZMwSCubm+0iZO7IJWUdSVLmEWVdXoj8meysXXDC/ichEry4OczH
qFlHfaOSKyKM6jMsw23ExAyjNzuEuZoNO8SYv3wTWcQXU22AH7eBdoFaBA1KJFgS0M6blp1H0rzr
H9e9kuwynWZjQvv30NaA/gpH3SS5dqeQos5mJZ0qhnWyOImBoqHt/myCrM1wNY6IC18zHBwxeOgj
gnTV6E5p2eYhM0hXGpCi/1ezgmLToEhF5j3esEt2rR32vKmLGDTXUdeWNS/u337FKZR0TRzKWEIP
mbYcqTJLZ9ttcZ41O3Kd9Ak4M2+oIyEXLCrvjyS5tL9u/kpxSPWgSdIUkswhNVxDbmRFi0hpw9RK
Rz3jagWn0rf5MAUUPvMSi78R+nxVVeSSDNH0VJ1MSu4TgwdW/ujQwWIcazWwWArcRtjIT0X3qmjv
HTRcLQFFdfpp5JgnnmxjXVXqWKHX5mBSmzlUK+jkT/XvokU27vwT5qY0DBmwotD4lynDeq2wvrCr
aVxnB2N+PlJaXBxzVJZ3GT/0y1HvV3BDIMP8FXljz7YHCH3oQRNjMi3iWCwO6mb/RSjBHKuC8EM7
FPX8skHMlSq6h/y/r6cpp+uNKtWw5TzuZ9554flPoB3uLMbtfAPbKjqyYiEisy014S/btZ7ZLwYT
BRisc4KVrs2PGatJWLnNourvsCyvRzeMiFk3bVbyhdPBiXEq4AncAaXxX/HxSRTY1H+3djbiRAsl
LJQ9isdcjaOXCG0ln0owjZ5yquBUL7i25OxS1HqWS18biDk3ElxDo0UGleugP7k8zp8kuUwmv5V5
T/DhBbIxZEZfqOjXnlzMH8bO/lg55QYz9dtnDYfbkoQx/b+wmP/Sq8TlSDJJMTSTPwqlWV5q8gm+
prpWViCyu6mT64UrOzi5l4gy+RBsi1GIAHZ0M1wDDC5ZEMS4P/oGFWaEEsORB34NZIloFEcMHYY4
+MT9cc95Yphd3og2qRgxYU29+NTAhfQ02Tzvi9YyHca6uJQiS8hEDtCzzNY3Yq8uZg9XEVr16U3f
sj/7S8NOoPBGCpXj2jQkMaUEH3ABzYDK8l+dbkRPh/gvH4ULMsJ9E5yNGsStrnYDpSEeMZFvYakX
sGuIvYC3K9LPf39xQ9c4AdK/Umd81Pt2I+2oGpE4m8KvZNV5JekbzziPC/dCFG4UFFq/2HXQYLoR
jC4De1D1bLSvAxs596JPyD3LyAw9+5RZLyHrRaX4tUBGdlMMHZDHNjbsm5PF2q9NXIHLvamOz1sW
pBziXyf1nCfGbP9xFqwcOAWY+V0uGfJTglN6CLNUpm7yPQ055tunnECOOcLCZm8KYiYEOK+Orjl9
gi8B+IMHXxnWUlRjXuKH9eFaLNaZXbXBtCg/GGiVyijOpuQRYFlA4A8oQ6OzaCV6FzduqU8R4Ur7
OsLFvourYT1DnETDNVqLHrhXWdnykU532Nkw6HnXv0KVcqr1ELkw4tkME7tLtNYB3CSLoj24RiGR
VtbwDm4XyF3BAca+yoStLGD4omu+NBntQWIySZQy9CaRBAy6VPAWM6bDX9YZ/gqsTvM4qK+xn80Q
QaH4Gu7BMAlNK283DjebFQx+zXzOn4dnHek0hteocoQCNgUsF93PWXQeJF9gopxmnJSqiOShACKg
j7PeZ/fZSssIv6IoB7lAy3OtQBF8eA7NYXiNtDebReX/tlXzzDA4mGSGdW/4pw+t454g27wmmpYX
5IacPACYEJ2DW5nR+q1ezm7DoA/Qq4YL8dEWaQiCwXY4Sg3FyNb5fsV6jh+P23KZGAE5Inw5jtA7
jLFZLL5ESjjmcg0iF43YYCZ7R3SK6oQjnoXpACo9w4YSp3QMNmYmUTNyubdEKPIl/OhJeIeheXI3
fR2UP4ldL19IRymKlSy+qaYpZGGD5janpoF8f6TTgyGCR8G1+LQjhVEKa1lmllF38jurqz4pCLoO
hATJersYJ2Ex9gulI6zf3mQj33REE6YMwqOBM/EUF9VOnIYS8+H/wpAnYB4HvBAGnWxftPX2lzyF
B+tXMey3yIQOd3ziizHUNAgKsx/WiAYR2eXjhG8pjX8ui1cOj3mtKYtXtc8mX1gvJPa5mTK/bMHX
2QSk7VkoTvyGLxc4KSdH+Q4IT0qIvirNpN/uz+0hV6J9UarulVetUheGxmJiiTZX+8H7D60mx45x
Nb3JuAx4cs/et2wZpMRD4wsZDkXDcrcHqHtm3wtxITaXnteWc1zs4C9l6kMxjOLKHaIkEPTSuvaN
r0ygkE7RSvL9pI8cqkxNBMzH0Y8NMBim4adduKmWd3eY/zw0NXw5hiVAFhiMsWpe/KoYk75e0HFd
YhKJh1CbC6YjaMJpHJuY5ArIduLZy5BkXvs/CzpIu4MNzSy2iSYWf8GzahUGowGNRGZTjn9NzHNE
owuYPo9l/qkcUrTigxcKGgBMVOSmfVjjJjqxUHNPuxxg8FvcYHZvhv3s1RSx6BdlWzsnPSJHB69V
xA7SvR2dMlbVXlNrPk//jgrHmqiGa2ao9XkzBs5khAEOuqlmiulNSRgLDoQPF5Nyo70vKx83JeDl
cbxhqjuSFVMQ01tuD8RYfvDmlkwmZ/W2qxRXKUmIPwrw6WWbQhRom0gTyUQ8C5zhzGc/s+p4YMj2
/wXwdk3mKA78Qr672K4jGUeWOyFT+U5h9MMDQScNXKlaCnvt+O5qX4YG5wf9tXcb7we4m1egIVuy
vQhuSg69GyjHOgrv8OtSwlPlMOfvTh5hmhmlX3zzP01jGsjkyZHV8VkOqCHFgjhhBN6hcPFfoySS
5nc3p1NJ2TeK6AXECEL+Sbf0wARtqhNDCrSXlaWPC48BLvtI3v4m38xQ4wjZXFryrVYI9qD/Y+W5
IN357OIP4FqfovBwulzYK1FwgAJ6Piu0XFx+qDbn9x8M+gpraqxWfY5LMvfrufEzyXcNwe6lDsiC
LIoIwUQiI8ONLr5x8BR1F7wK6V2JcH6iiHBDB6WLT6jAVghF6r+xTZGLv8oU0kqabfzKG88WBN5E
0kbFw4g6jGqHsQamqZOLAr9Tem8krGvvkySVHk3XiRkYegRUUJcGbE5Gk8yiDPmLuoAyI7cqikVP
ANL2GkH57X+kF01YUbY84258qzzgewTaSv3UxTa4Th9zXFZjh2P2kEwy5ldk5yThr5eaMEl5gqZb
Q8nxPPlCoMwSanOZgBZ4DSEEFseW6oV+RswDkR9TYvfQU+gQBTOHt5kDqsPdn/EypbVR8DYPa4sP
LVmVHKKwZjRk6Lirf+Nlwx5MeEWI8XR4AMdVuzB603NqB7lH7tkHg2m+ZKncbAG2K8kDYuDxpGsT
xkOc7qYgF3B1842Kxc2V89CE1ra3/uGR0DSe3pNX/q0+idniSzW/HIzs//NgYDdUYgIzFFaD4aQV
go0XW5a2jxtbN35DpgCtb1HnfJBBE77fE5nMc0R+VP4EZ+xM0RTSq2rqkYqH3lg0rttt8hqNQZCj
eJO9U2zEczavy0aa8cjgmKgtOaP4Y7WRD7v7zpZaulBEm3xKdBEvpURsfFfsbOXrKGOdW5NcfSAb
75kGTQJPXdHABQVgBAipYZe1ZBX41Jr9DYltQNIqOFosk26iYg5j/BCJPeJhffBj8LyHN/J27cnQ
be6Sy2X+tYRsi6HqexK7QzrGxvSy4/8UsaGy5wFlRVJDmrEOEhbpiTZR2C4Tho5c9a8J/41xK4U8
gWGUEq0muGyUgN1iHoNt0GyKEewksZslj8wlA/7IMMis14SzV4/+y5JgNh82iwxwbtJMh50aKcms
NFsDT6S0sqIqTOol+sWST3Foaq5uTcPkjpvg5a1uwOhZg5Fyo7XZEIPSXZxy5ys/02qjUkeci1YL
+UO1tpajpeR2IFgJhpEz/ec4NbdRIBU/Z4o84De6wQ81W/5fYcnbMoDt083nLKu9RLJ7LpirZle1
NdKDBLOjBPzfXqGWZVUDEAWB9lXDxaXVuBjmFXL9UfxH2oeFUuIwcOs4+OAZre13KJg6VfUbZ1+v
fjnwqVgD0k7w8IGti9eb3IF9r2OTW4sxUvtlmLDAnq82vPx1SXvzco+RK+W67biethnbrSONm0vs
JLFssOOBNCKgEMVldNWM8X1CZYNELRlUFUPtN2ls7H+6MCXveijoV/KHMdAM8Q1x494lbECCwwEo
iuUHdWXEt2NEUrPpTThW5wm7iibfF71TJ6c0LY9Ba+13XLCnrMSpCGiVVPuD09rpjmn9kZEd+AE2
V0WPIqiZoaUeGsx4ia3RKKcf4lzKkGcRXbmdgQUJrpkDy5+gduoBZXgTL4NytNzzT+6Fud67PWZl
5cOgYqK103DAz35Tkg/WvQlvLBeP+ZR+rG/2cMWigFBVekl8Q85mitrR4pwW10hYVEGKts9PwfnX
W59u5LGUc4Vqelhdru7LUU6MXdFeSrRNIf/zfUitrrULAAaDYtlYywUZcCygwyIsRhwpYcwGuBDC
pjWN/VOb0bc59ThDbmKMNGnwQBpWl6KIBSt9ONm0A4MAD32zyCKCHU79fuGzBLsIwXH+Nn8MvLn6
Yqa8Xil+EnYQurJVDqtQ6ppJrAtynAy9joGh47s8ZlsKdf9sc0pjp7c/6Gus4tcl3tcgWYQuhZsJ
XS2PEbKHDH7wX6f5HK9vHFgZFcB98AZr6JcD7+PGAaG1shR4KacQDTWVPmTok6xy0TJGEnFi7Dqb
qFnvfVBnkn9Wj2bJrbJuUPtDx9pErGHhIHnxsfKG+PU2/wjmOXnQNYXzACq8to2lDpDpojvjBUJ0
8bKgcCV+OU4hArJAQnTHeBgwhgm4F1FSXNI/O5D1RtHIrfUDcdrESxxhmk3ogmKeCDjxofQo8ycw
J1PpFYsZny9wq168sgWzmNgW9UxymCA90thTc7facuHLt2K1Gj+FVIl6Gl4O/AMuxLbYpCDc8GHQ
NK7SbfpSMqHzkRZYdMmbCRBDB7girAEJIN2qJmcTc4OxYbHEo5coY1UCrxSYGc0bdOs3j6JQJyZh
QzIj7T7FYGICujxfE7tPtRXDiXdnZpr4sUSNUKFrGiy7twu73bLN3YlusgrpknFuwIwW+EDBvN3w
qN01utL/2SlDrwXUBFQO3yV4wJHI46BBO5f9LeCWVzioxGn1i0hD6CHqEzFP57Uii0zfuL2IrXZb
IbSiSA4+4XgCdrk5e6EnaJJeWRRn17QOwSp3JNwoIrQYAX7AKKd6SfdZ87pR+xeSdm0o2FF5V8gd
KOf839k/4iSG/S8pcuYGGQvq/5y9N01LjbgOdkmG3CxAFm2RCphUdml2YqH+p70uQYMvCuxLbXZV
rsKUmHDdOAA0Mm/KY3uHFftLFPkEESzTQSd+7s7Ly9sNYlnQpiNtVU8jvubC9RFtDJCLz1jrf9jY
Cd1o3gMmp2aqR3V9FR8X7Ul4yqe5tPJ6UVB8Yt73FfGiYxeTG9IHZb8n1KV6fzahIdo/M63eWT6D
ZmH9Qh2yuyGcF5FUBw+U2apKp4kHhpAb2hR7Ai0yKiy8Hc5aVxAjy7Ee2sZuH/PeSC55c4rsrXn8
MKt4KXX9jJtEuhKs80+h7DH5O8rdFvaFm5oR8dmOb6wdQcdoXSiCV8Es2Dh/Ie9PxgV8NRYZe6ZR
ppas5OPf1RLGFsH/Rw29sQx43UUsO3leFE0izpTSyxqOfKsBSoKpUL0Z3WuiHVXx87GSslvMOTdz
2zP3JERmwUHdoImz6FpcLdmqD+7x8BdYtn8ocoQBSxSPwEslHpD/2ddpT44cNYabagNRZkAp+niK
DFEp5aHUUQ1WWs/OdIraG48Xfd+yd5TTjpw+f8svfuHA05QvUWK88ky6IESkXjt7hYcmx+MRhhZJ
/DAW0ucoIZuI3h8Ex8hGxZl3wXHcW9AlP2XElsAj6M1ufVsMnAO8RK2i98kGNgdi5BHzFxP47Kgd
QyDMuRT8MdluphqvyEtbHMAg2no5wOMWjQLJaacNXq9CD1gcoBjHWd7sVoYtRa5QPSN2BvyIKofx
lwJh1BH2K0YKi6qPTtvI/yCVjC6iKBvvR/KrsOa1bK1GvvaidM+46C0mV4H6kCuY7ez3iZN7Exiv
xTxl3XTNzqe9QiEdXtSMmPySbWvxnRbJQWm9pvDbze/Y5uF91wfRGLmkdqAk9+se/nYIA+VmxiMj
Ks/BrTJ+4Vt3MYJ7F/zupyExWjCpavES6lbO7QhrzvRVCwGEHpZiEw0aLhKIoREsu58ZOFuSodxj
pOQZxqu1BzR1ezqo/ABSu7JCjwZhXPF2z8F6PsXM+pR1SEJNoK2/dS3Ghe3Rc7mJaD3CKwKVGQ7D
+1HL/1ULAoBEZFch6aoJUM0rP8vX3ZQ654iJaVZp57V4K7UCbTfaoFpDiisYQ+bfYycq69XBI+rz
fRhJf6UlbkOqSJ7817lswrYTnBjMcYfB1mN6g+D9m91FUVgG07JMQCwF8AH5TwMrA9KOwFSw5ZYQ
M1fG75eNuy6IZFoUcegKIDgaNWJYlMH7P6icbsNFsysRJi79LffYF048QTJn8vDcBfL3zQ70t1Kq
oKZ7fMegPUuGrPJplHrNoSDT2MEuuSDJlSamRiwI2pGhogYOwc3Z6ys/Fi6GWDzuduCDYZ8cbwVD
oou6fLDLL9S9ySTQmH/rMuTsgOqsHnyAsBh7sxETgBUAnmeWdK8DMyo8Z1QowKayQeFIc0wQgRxf
KbXSQ+Rldm24ud9lp5cNtHQ9Q+WSdOu/E9YFOVImw6u9uDYI7OU3IdIozg9S2hHhff5wSgxhC/3R
sDoRkTM3Uuw3SOYVAW1mYLhd+R5nsax5tAT3dzggmZgrqEC4SaxennPq+04bwM48BKqoXmUEgzFG
11L74CE1HzGgSKN8SzTFeT2bAVA+VYuNKiFnoC1lx5VzIlEYqEejC3hgG6cFMFA7IZliL6KEsu15
nm6ntN2KUqYxCmbesmpX3yGl8T5C1BH7brIWLlkSLSXFVQMAA/9dShgAY9hbyGfRjU82NTRAnlOT
Tdzb/aSv2/LTHCXexKZ1aPmG3CgaWt1mgySCeOOlw4M2EZJxgr9WgHCDaA86x93CXqAl6zV/k4Bl
J+K5hiTvY/MV/kwTsQsPOxs=
`protect end_protected
