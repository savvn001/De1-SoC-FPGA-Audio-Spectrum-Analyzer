��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	i�A��@e�(�(jڱ#�����)����z�N�ףh'���1��B)����0f�q�B�#��qBh�%;�hj�,^'��g��p�r��7+Rֆ;�Q�e��d�B`m���g��yC{s^������Tx�3[ԅ�����E��}O����pL�|���%������UV,�E�#�+V�qq/o�83vv�P�T�3��@@F�Z�i�֌g�J��鑼��8��X~�`u���z3�b?�ⳁvz��6�57�#|��r�5��ә-����-u}�[K���#i�4W��� �/iI̞u���۠��$��BOMJզ� �g������|~��3���U�خ
]@�`ɱ@�#�	��BB��iy3r[f��.��H��!��{�hyQ��0��l��E��yt~%o�1dC�V|��k�4(�T�@R�N�cF58,�����Yu�5 �� /����kr;����,������9���1��X�85=��6l��H*vnC�u�6�2P�&�I6)�2�8�����{��w/�uz��[��(��̮��hV�SQ?��'��S��I.{ ��U`���~.qOU��7��`�a�.;�k�/<�8����OFov�g���JzF��Τ`6�wR����+4˔tÆ 1�7�\wXXXGx�0��$�M����)�*߇��2ڵ>i7|X,�$�q_4 2) ��&*D��UG���m	���1"�^N��G��ip�-4�d�<�i��{X�*��R��L�H�r���h��{���kG"�l,4S�$����yi=W����*�/c������c5��У��^�X���*��ߢ�5s'�Z.n���� �^J]�o�	�2�i�h�`��������o��%��@~�2�C�*�u���jN�B��т�(^-q: �o���78��(�m�iaC^@
��$�s��-v[j.�1}��4��͌�p� )3����<T����{�6�O���p*"덲V��V&A���*��p���1i2�vd���|�c��J%y磥P)o���M����
��G�GFJdX�z���Kx��~4+�w�?Nw�1sGRE[������-��h�9XH]u�L���gJ���w�%5��6���ؿD��B
�>/l4�ə����7�A�F��آ�Q�}�ð���1�І�-ޱ�����e�6��-���"܄��1�V�֦M���E��k;���9����!�:�P�ɟ]d�ҽ�x����~��*��ۍ�-��G[ux��!���u�g���_��,��*N�8���)�Ph�fh������~�eJ��n�h��{yѽ֊�"0DC*$ʧ����ݧ��(h���f�辒�A~��ܵ�#h����Ct�ug�Gҷ�bc�a�G��i�<��Cתz*��2:��`��ޔh)�e�"���gC1)�~y�+~ GpR����q\�ߌ�����g"��u�z^�R�,��Av˂Џ��N�JJ�?OEQ��v��e)�,��A�싫$���ڵ�7�������@i����ye������<�S���_�u�d����ѥ�a$8�aTγF:2���l���_���ue�o��U�>�p��i��	y��A`�ŉZv��j	�_�U�7����c   �\hPbxJ�����W��Y���c[�X��K1!^7��fK�+������5��(���=�Ɩ~IM�������&�/������E��~��u�X�N�%	T\NO�C�a�}D�'���(��m�����S��MY����87v`U�o�ҁ�6�mD���S�SKB��ٚ���_�F�`]��V���cA%��s�	�^�p����9�w�	p��a���c�:���SMm�Ga녢�#f���K4�N�i��5� t��� :)6�w��n��A�n�X���Lؿ��mWJt�8/���/�\ ��� ��go�,m��X[��Fnlr�K2��`	�v�0���v��'+Ac����╢��<x����8����Lj{ޡ��_r{��1P―W/�qf�x��f�<�{R��z*�Ց�.N�!���|���F�A<�c��l"|O�ֽ��x�6%!T��ڄ��#��M���I��W�8i����lߠ�>#<7�̈́{eһ�F^R�Y2�_����C�S�KD��)���-5�7N����i޹�o񱖢׵Ggޓޭ�m�5��e�*��Bʉٴ��?t��U�o��/�\Y�eA��x`�B��f���7���`m<e�t��n�A����"��7�q�!��]�9�Me/�9�W��T�N���%W>nk��qm���X�A;c�ަ�P�E3m���V�Q��^�mfŢ	���������HR����l����b�9���8
����*�*}�z��*�vX����V��c�W�^"�g�q���|�Y�'|�"u�����z��00pp�$��h�tzނ����Y<�A���? �g���=�K��zB\�XÜJ�f|=7<Oe��B��Z�h,c�%�m���䲏��k�R>�&����p�iiR+��*�����E���d�}x$����Z�7��9Juy���PQ��2�����)��o��=ݲ�I��'�-U�e��R� �s(�a,đo�7�k�&��3�hx�!e<� 
�a�nY��:5LZ��!w��2�b��X��X���%i� ����9�)ؕ���^_��Ϊm��M�<�����B�!&͋mġ5RAp���Ơ��ᰃ�y-oOLD����b�2U�%y��i��K��ims)&�C��X��n�l��О��w��l(N{��1�fS(�c̻��tE1�(�X_>�������g�6ԫ|�+do�QZF&*'��i��)]i��;k/P>�������!�����Ccp@����{J�A����^x�'�-��t����"�}�e߇�z�>�t l�_ίx�7���t�'���bf���:u���~�NMk�%�Ⱦ��jbw�.E #��y�iPg���D�.NS#e$��'!�bN�85�^�MT�����ᒏ*�~K�V�&�̫����`��x�O:t��= 	��S�RYB?�I�?mҺ�������W��16�L��'C��G��f_���3��3���K8O U4�Z��/�����}}�V�b��OC����$�q"�yO�,�p��kl��#�J�ҙi;Q8���͉]�I[��7i����/��Xƥ�^�E�^G�fOlM�FxQ�;7�sm��g�/¹xx �TZ����0r�:@�h�!��`�y�����Ļl���Y���_�(HBnq�8���F��%O���O�1���+�I��9�+�qT���N�,u�=Q���=�_�B{��t�Ȇ�+jN�(�r@�{M�n=� �dV�/ڮ��^l����u4�!r�o9�w�1��p��o�t�g8���bqhϏ J~��*��2�����O�ӣ��H� jO��W)8^x%GZF�L�����zS<z����h�h&�"Bd���ф���x󿆣e�'3(!�=B�y�`��f⨴��<m4�Y�k���l�峽?�����w�ڋ�M���p/�:ڈw1#չ�Å���0kMEz����^�\C��xGf�E������1?�&)9�B�͛���)���m
����`9��!J��M���oW���U"���a�D�[��B�8��~,�v�W��[��4���)22�� ��Ě�O/V49_�����:ͥNu]ߤY=����Nz������I(�n�֓r1lY��B�R��u���]�Ua.m�,+�;u�B�ڈ�;��m�
QY�h�0v�	p����i!�=}=�O��Y*��R���� S�a��=�m.a)�ම���;r��)nt^](��+P�F����(�5�g�Cr���3�T�Q�;?0ő�u�TA��S����
|��x�3�Q� Z�V;��z���U�9��8K�`�Cb2a�*�"�?��ncog]-��þ�멎��\�ނ��������y���8�Zm+Usd��CS�<�ɤ�-)RO����QqR�4bLЊ6@H�c>,��i!ϥ��u��uI(vP�g���>5�ܡ�y���(�=��Y#+l�J� ��Ӭ�SUA�*���N��?(jj�F�3)[�_�|!�r��O�:ށ ��+�\�h�,�"E���1g��Tv|sP��ry�&�89���jS���#[�U��e��E8/�������� �(ZF���,�۷qؼ�!Ps�K�Eq�FMC�##32d �����|	&�Ifg,�|��X������bW,ZEz����C�5{������cB���O����t�w��m艑�������I���L����oa�|l��)m�&qm�+�3~x|�N�Ğ>y?�~�Y�,�փW��"���\,�6:�9��t�/����'g�=R����[�2�	P�o�4J��s�R�V��4N'���Pl��B�sa֠Ţ���`�,���ݔ�/����W�g���׮�s(%�� �U�VI�9�Z���^g5���ф�i���ԁ�45�H,Qˋ�ڀ{l왨���i���l�A�tT�����^4��'RauT%tIF�W+��1&�+Е`8�	R��AX���!��bȀr-�h����Bi1Н���?��Ѧt�~���̭z��@��i�����r����fu���ǳt�){�>0����|2�Ҙ���X�����P�6��s�h���oF�� V��|L��K��~��R��z���8P��+�{�2�yT��d�d�X5��q<#B���7�i֊ܲ�Z�0~���{�B���
htڴLSc��C�#�1+��*�i����P�&#Τ�i2:!��=�FˑS�:��s?����������l�|Z�Q�W>R�2�^�h�a��
й�ɦTvR�P�k��G�`��=�Yw��tH@l��O�BP��vcC,�/�N�`��vh�<6���`�m�X�d�r�'��Y���.tvA�­}�2���YΗ/%{IG�P����&���?�N\ @>$u{(
2��9;h�`�F��O/����T~8E#s+J�tӪgs��ʃwTQ֎Ra�=��=�P�$��?�w����~Ӆ�q�
�ǂ�a��zdT{}L�D�p>K���N����uYY��n5T�ɕ1?��<�&��y˨��Hd�W�U[�'�B��A�<�P���ǹ=�#Jap!4̬FyRT�@X�ǜ���ޘߓ��H��>b@�e&<$�+�!����p��������PЏ������AV�$��X��0��?3xKA�?;8N�'�:�0�W>��y6��U���;1O��˄����"%P1J�(<S��s� ��>��8Ie�����ݰ+�����_1Q,.s�iR��(W�Իz��A�6|��.�s��;���m��}��H����XN�[̩�x�T���[���Q�%Fڣ��+�B�h7Q1e��N�&Y��YM����Q�)ic�i��d���Ձ�
�/�͊�k賙�bGr���ʮ>�[�Q�u@G{�o��AZ'p�cWF��2rT�=�Ë������`6В_Ƙm��̈�����c�\�݇	����/���x���M��7��r7X@	�{e��[DWJr ���RM|K$@~�84d��Z[����9m��Cv�ʉ�����s�k��0*2��Rqk���e�h���2��3T{��p��6Z/�-.3&»�m��o�H,�Ҝ�:XW7N2\l^0���><6�������,�����i=ۜ�dx];�K`S�v@X݁O��)׶�f}��_�`&_f�$$Y�$�M��F�5A#t!�OQ\b���x���m%5�h rGŘ���<�t�i�=c�������;�QS�`_K��W&�lc��i�B{�����0W�:��&-N�;�i �ܘ+p��[��bo���0�w ����c���t�_T�R�@?x{�\��h�{���h��|U[\���ߪ���=��7��{u�@rt��Z �6��r)T-Jѓc���CH�o����i���<����9�qՀ�մ�����Ϣ}@�YLǠG��F�9|���"������mm�d���q��AA�Q���Z��(j��Y��{������.:��+�U����.9�jk�pQ���ˤ�)�� � ��
Gۆ����-	~�!�%�p��*���?��Zx�LZ�+-cx��~o�x��w��U"jS�a"?�&�y�Z�Y�enA��|ʔoȰ�R��d��y�YͰ���ED*����U��[	�	�T��v�N?U��k��G���ڕ�}����� ��0������?{e�ܟW�R�����"�[�A��<2cw�P[�U��aL/T��ȸ�ݾٽ� ]f>��c2�ͳ�mSv���PYj��1Dyێs7�ؗZL�^�OL�Ssh��8!w��aw�z��Q� ��ͻ���kp��H}�����Bf吥x�6y���H��׷��pR#�S��4������oH����!E��v+��x;?ש��*
|�o`�^���Y���� �b�{
���f�x���� r"f�p_ҙ;Ʉ��L�"�'��%�%m�a�A��wȱ^Pd�&)�{��l�]���HJZKu\`�"K#��}��b� �r����F-;,p�.��W��Ŀ���dU!�����/�v9��c�;�А��څ���Dt��{���x|q�=��$��
,6o�}{�+��1�\�?���W
�����0���=� �"`��9!�I��'��k���= w�/;ȫ�0 K��z�F�,�9{	8q��=ք���C�kqD��j⾮ކ�'%��v�1�zf�q`��B�n~zWɿI�d���޺\�uӨ/���	TT]�ڦ�&w�nݲ��X�EE�[�y��(>�O3-���X���_dYcMWLN����f��n|P�ß�^��V��T�����W��n{:3���A�s,z|�8B�=y�\�W(�T��c;X�=������n+T��*��*M��Lg��KEm���v3��&�H�4��C�ڂ�6MX~fvG)����'S��a�`�!���� Xx=	Bw��Ѻ�'טy��d���쌜��	By�,`�R	5�\$��J�Y�1�|$zQ����&Э^Dl�6�<5�w���;xDh�����ܙ��KA�ry��GP�©j~Z���H��5ؿ��b"_c�#i�� ��Ԇ��		�T�C��E��u;��7&ܾ�~z�݆�T��`�=�Y_)+ͤ���vY��ua����^��V��9���fU��&h҉1�P�Y�
	Y�@ �Z�t<q����]ܣ�I͡Wet(ٔ�`z�#"s�ŗ�?�٭��ҏ%� ��S��b��DN��z\ �ר���۝�r-R7."=?`� 諍��-�W��]�DR<���rX9����,r�% ��lu2_�2O6n��R?D4�I�г�e����j}��uJ�)��8'���5�>�>>���*M=,� #}V��t��tG5lF\�k�0�����e�\b�]�:�b�5�U]��[H������DJ$x����ܥ6�������DXc"ܦZ~�蔲��-o�����_V�3���47sH�Ӻ\��^���ү�|!��Ɍ�^�͋�_��T<�9	R�"��bNf3���Y���9nRA�c�w�K���'��L��Z�d�l�Q�
ԂR�3CZ�^��=M��8�(m�����׼�XĠ��;L{��V4���q·�L�8�Y�W�n.5	�#�&p�JS�d�YίB��z,e�Ⱦ�M.���`��͖�aaTC�RQ�Ut#���.���P5h�����\�����T��=���$�HՒ��"e��P�1��"������c)���&yw�u�ԕ��s,h���.Nq�������#T�wW���J�;�!�|S�طye+�0t)F�^j�W�&I�R]�(z%l��G�e������ި�3"Vy����Fr�G,�9n6��`W�H�s�o�7դ�J���/�Sgf��1��~�0�O�}&��ː�@�`1Q��~9T�Dd�Q� �։2?%�ְ�Bo���-��h��d�	�YH��&��[R��l�����wKE�)j���.!kC$���rcV׋ ���=fX5*Ҷ
�(�Q�.	H���E	7-~���N����-��󀮩0m�]'"�]-�5��ϓFdƦ�d���`����^P�<�k �ޏ2�A����C�T�:p����B66�w~,SY���Ya�}�zÉ��>����kP�gT�7��}�D�����ǂ@M��=�a�Y�p/+� ���*�<��Q�+�>i����ky4�6a�o���f#���X:۲��ƛ�\�,H�ǂ��g\J@�Id�[
�G�U��9�-��B�	8O��{��d�+��3!Ǝ��&�9â��VcH`��K�I��N����Ǆ�[���vI����:I���~�G+�ZY�~��t���K�ݰca��1�u��c��,]��2�^���-�;V�m� �,�#4��z�m؛(׋��{�:?=��� ^1� Ǯ�<^���r2/��ŷ�4w/i�)��q��#=)������W��S������ޡy\2WE�M� ���
.���XL�&���A06����!�`����a�]d����qn�@,rJ	�X��S�L��c:X�?��zI��0`�����n1�$6c����ą��T��1_�5`��u��/[���Y�晥���Z�`��ҡ�i����K�6���X��B�J@��ϒ=W�:���#�k��(Yr