-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
p3H+RrYDhJXa+34bWzp+XiRZOmCbrsXEOGnPQrlesOwchBnOL8ITAE1paJUBFQqTJR7VsRykOnxL
FgpcL1nh8JDde4RO0qYoMWGyq/RpgshGzRIW/gR3fzsRtRPFPIjywBkuV6KnQj7HRM33VL7O4RnR
zyVqfQAsojlP3HNunLLxn1tWDOYxKm+7o/xweuA1ROy0FUh1P+DUfE3u/JqK5Ck0/qpbHmq5mCqs
MZwaXI9at/2OdNBG8jnHdL5CMS9zz62yW4GBmB937rkwEvwFJl6Oqu50jl7DcSLoTXY8eTHTL8Kt
LFnddI9eWGRsbkqliXtg+bmtIgVgO8Wab3oJfA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
ZVvr3twzrKoIB2iNcYvx/UoP2CCSHv+HFBRQdVP3jbSwIDFPj5WsH+gCcWnkJh31LbqFtGytGd45
/5z9YQvecGm96trKO62T/VRTL8M7f3ncKe+5Dsu/QAfU3ZVMWrRT56bunKyf1NFNZch1U2GP6w7b
AE6L0PyJSvSRyWqFOy9AeMerwsw0X5evOaEWR7aSlWjEWLT9ubBboZvebFvwicKsnkRU/6zzlzog
AjmcO/mSgKxW93tlD3CsufCvcnhJA9s3yrW/mVr4uSVznOu9buv6A7wprLq1BwVk1Q8oD6Ce/EAA
mGIiGKm6FrsdNBnGZQ5lKOb0sNcKoR3bq+Efkw02HP0v1Bl1+l1iK+x0RHbNjjdRb2aJBy3LSotD
FAhrqO0Jo5SxqxeoQT6vVlopb5XTj8vf3Pb1ejjX+6cTqDB2bcHJSrHaDOMufA/wSkHc0Fx2nsZ+
3EUcQ6goUotB6s3Aq6Kkj4QJsl4ju89juYyNrvVIbv2KrhX96z3f0KSbJ+Hd5hC5caNcE+ta7GGb
exScMX9ctq5tDCTwEwlDm8hsqrQlGdTLm9n4RQ8sqxCgItsNvGjnXJYe4RSHaxidXNkFg9+MVzcx
YgRYxd2QPaWA85+iFR3MpQaSybIDikXJeebxfZj6s+M3GehwbH18x4rDWt6HtlD+Ktv3NGApxb9z
Xl+uIfpUSOqU1W94/ciUftPwkMsnRJhkGHLhIJOhfCgSdZHwBkJTIyGjCrY1NPRJJq5noHI+XuZx
8ztgIA3AJTNRszMarqsd7mJjZvI4Ysz/ECbzJwxb3dqrBrAxI5fcOMXh/f73sBFaSq/eeje/EkfL
E3OX9ipeUizjx/IbHGzNpnsK2gFz/u2xdcATRo1XGC/tbMv7vwXzCx24HfzwmIk5qy8FCjItHClq
Z9x4TW/mJO0nuwVw5EMEEoqfVBtdZtaXqlHkwTL0dTEXDh/6g2CB/pwEx2frU0ae02A2tXCr2sk2
3JFG7A2kdeJozYJvyhE1c4+hg46uE5//7zzYcXM1bflyk6RcFOZJ+Xf80eza7JMQNhHhn572SmSZ
WUym0L1fP1vWBtEoJR2ZTAy6YIPFd6zX+DYv4y+b4H0FK11E0Cmb9pYyY9imxBYBxr25hTqAyo/s
JrFP5hWqZVPt2ImIVAuOb9I3EfskTeEtM3c/0g7bmuemW0CCBlRghMwBpIaT8h+fQDEfGy0fbywv
WBMe7jG/Q3M6wA4g4lAfgl9c2ncNkugZCwQclzLC9bQIEklA/913l4FRAjmrOOZ6+hdASGTG8jBk
Hy9Sh6eGU24q0mPuKIpMz44P9COs3dNvrEAaO9q5Rm4OuvXMTN5I0aqPootHt1vMTUX1bgG1XfBY
qO5oJiqe86XfnUK04OrJZnGtTTzA5QojxQlvosorVp7QHkdFJbN+8WVoE81QUZgdUv07rh9T/H1E
g7HPf6PfDsVvgQkEkdhYUIMxEnA8jMB1zhd/Ex97UIXUxk37Er2Ti7LT14ND5Tg436vNuV5ckUf7
FmDw5J1KCfi362WwGpW/cGIkKPzS1SQR98U27BSnFCmKInIgksgQi5az3EHwIHGlQN/+lC/hd3KM
yFbXTVzJ4QPJh/46yQx1D3fz2QE63nIiO4a2KUMEodEqWZUub4voZPlBsm1XyTM6EhMzRRfdSbOL
JxVQLVncG09TDpNzfweqnmgkXBVjs/IGWDkcEaWUlJZlPPRsVA6NRLLvdFThaDW/afuwy3aIKWSc
1sQQnp2OoqdnQhhdL7jxKHtklB5Ua4Pc+xohoy6g2CatUbzpeM9lbv883BKBZyVkwgvGH+V4H3Rb
uTobs8UAlaGJGDmpmzyFpRRgf5F8Uwq50TSQ/6AFcyiPOTZL95j7Mo2lxp6zoDP/Hz2WD8OUaoJN
tbe+d0zD0mzAZzivwJFJPGeujPqOvCVkKZYM9dEw9E/CU4/jtjNfs0VWFLEwsE6w7xpsQjvly4Nv
qr+y1vKcHfZYhtNtajD1EuuMDQCLnlIFrHgPsc8l0iej63l+9h4Nx7AaZh7QqYC+gHOtGSAvraow
SjlDIhEouZlFhxeI6Mry+RmPaiVJ8Ls24Z0LuBh+wn52/hTTOXxEjejPm461dYhOSEoYfWnJrNFA
L/3Dhvb3KmRL/cyFq3uqxvMF3Jw5hz89n9BBT2/ahB8EERPSulSJHOP9fsrIlmBX8MJ0tHJaXfv0
/nonYi5IWhaEfDOKDkTz82xUQgx4kfYDEQ8s1ZBhbxwZmyKuNtnGeZ9Fx7MsINeBHz7YfxC5joQr
KO8QJqIluvCBbjgrMEFfI0sCLrSlWC/+L2G/D6BUDtlu9LMgHhN/KMgQGXd7NLRCTUJaxXxTQ19c
edpu64TfgFYg5ovexnwIDy9yrPQ8Fpt6g8LwzSnY5cU0TNQNRxoWnDGK6YktDUbCp/71CF58Nbiw
Cu3d0xRb7gRb1OmKtVHxpR/5+AY7cUdL3yRcFLIcrXkOjB39xYIqCHL6fuJ0slWx0Y3roopp+dBF
S/ISai/MibJniw0kqsjKa61NKBmSN9fhZMrfTIY62WLtdWecR9oFkdf5W3xk0dUQxWN4Oax7y2fX
VscC24qpGdiis+c7rC0YOURHd/lZAO6NB1rD42+Ttp+kGutrS09mkpINg8hses46BAy6VeY+eGNe
BKgqJG1+Usn8VQT/1cS+vsBZ5K3JxSCCiNKTtdHpCScpc0HN3m37GdxYbjmPERT89k4jzy1GB+ww
MRN33hg300yzW0MWnRa+bShOJ+HKxiGqGGK3DKcgl1ITqTGC2vsbDq6iDJKd4a4btcqP9Qh2GlAy
stO5WGl6LJY9gRsDV5bdECAQmJeZbbuJa29FmaVeqK8UYDZspnd6KYNrrGD2lfjXxQN1a15TBTSV
NuoWBDHhVz/DTcD81nqwbLmTmu+G+8tVSh2vMVDu7/mmKavjAC8ywrK4t/o8tC8wNKfTQVgBBxVG
VRE6REtFifYg3544EZNcFbU+LPFXnwM6/7/DVVcvbpCaizzc4bX5xsyaIz0epl8+50jltqTrhE4D
tgWgSqTRcdViGmJxuX26tbZV9qVTEhbY7CwasuF/1+N7K12DU/kV/EDXDqXzXajEJtlOeCI1jgh6
XP/G6K9de1tzFXNFrSWXHYah8HKoHopMSNZmbd6HlWJs/JLF0trlJVUfY0YiWm0P0EpMcmIh/eSM
5zkv2IpTC0aNdDkN9gni4vXhSa5Rmc3+BMH8T/c7ExgCdUFhHt6egbRSTWJZp9K7zocELkmh/nF0
E9wFYWzK4i5VgChFFkwN3BmFPmX3GNPFVUQ5/VQ6ejWu3QYpZXJTaYnOecEZ5VCZRu/pmVsQNS0l
3BOXKFftV7FMeYPIF8f3L2jQy+WPDDNOiq5Ezxn7a+VADuUQ/IJBFvn2kr2+oKcdtPekgMYlOa5C
0zGnaIuTNbD9yPf5D2m8l+an2VvIUpPyV38ga2A7RFzSXEVpPm19WqeULhGXCTgsy2rWBOQi09m8
4RKncH+r1sLtz08maz8dTRYfYB2YpxtUibhg0oSuyISs6akBkxcsZH3Xo6vAscMBUpWfiU8LZ9Qh
82zSJOrtiHtTHnGT7Yru0Z94IiP1c/GSOLTIcaOvr/xS+pUeVhwSZwy0nbYToK1vx6DlYLWi/YcP
jIn2+kkpPzFfFOx00mFJRDCHmQ+7J3rVNgEJ0s9dNOCma/pGspSR5WIafyR3wtbXhkEWDwNcTCHW
i0scrYVtJzegbtkyR/g8UL9h6SymQLm0qIwDNP8inghUKx2LGaYePsLmEihsDe6eN3T7L/kdqoZk
i+l2WNJqhlmRUqaVgZIHBNXRLXrgKns6zsb2FaE8XX5ZWuIyeak5yr3XIKaPp5sQflbZS0HpQ4IN
hdQUgnFX+t/spJE/EEtf4h/obyO/Fi46jx89zYrjwn3k0msxVd4Muq3AC/OadvbpdKQcVd54qHOi
HFx7QDYCbz6RcKDs+GRhLvY2AfJLgasiBeWXVERveiYv1FMhmGdg4D7FPb6NXMuDKVvQDfiS/sYH
K9TvoWzBCj/r98kA/09xJ35Sg1h5AbZUmg8NwfW6qNSDy0+8NRMWBtnt4j8NPkDXVPxM1WUlzCst
JE9SqyJaPdObU6ANJ4jULdu/Egd1xmFpHYuqquo3IX/6OX4sFFFKKylumEJHZWZe+Hd478QboAEe
W8cp9oPaRHmx5O5d+xHJmypRBBfP5IJbQaYXAxzla294RcZJEYmYUrioFrGrjGe1zQDBT0o4yQoi
zMbY2hXW9LxT7m9/ZiB3DQnNhL7yO7q5VAr1T3hVzUeeECX+lnM8M4R8954UCo9GIsJeK2gKLhwf
ui/JaPSdtERl/13HSIT2qFLQY/gJiVkBrqZ/Dk8r8dvJNKtJHMDnzbtSQJX/iXqhc1Z9aCG0w2c5
ZK/21rBauY4FoVLGfsFFkYZV24k/bgH9KwPUwAdQrMmIPSIrXOdtaTfOatyyeUvKsliYWwgYsxGw
4p4Yy338cWT2WKbyx/WxMYXTplqARHvi4qFQHRWEf263oGS5YhxLHvQSFc+xRsaw4tUy+ZJXoeKr
eynaLuXtgbomns9I/SmEjj9ZA1aoKMk6dcIcb5Q3f7qPQrQtqTZeH/1zII+jCvoS/RQmi/drqBU2
MiSnD12O1VaGy24900rb2nbGpAxfxw2K2uWFQZZoKxde42q+Xhhtva6ify2KflYPZo5zRoodoSYp
aDXHgAZFWcuDi9rIW2Isl2aw95eHAWz6vTKC9ikaoruFTdhE1I33LW8sy+X9RME3Pjux3nMw0bw5
cv7ZcnzmrIidV30+yOp9nVt6IsNIq0ZvqV/dM6qqFB2fmvQOzjXz9WHklwyLGAI9SmL1Z397Xc0/
DSM0qO5RZPBP/eSk4Ri7Q3wXy+Wz9fJXtllxDn502yJrmvaJDJpwB67NwlYuaysHtSGjb0XKPgAz
wpU2/Rl3czhAvtmMH72f6e7+dG2KSL1WG+6WWasHPSyDfNcEvIgU24FEcilGeX7CKV/tFV9z9k7d
PLGt5KEOecB1rcOhOKBwiO8myegHx4Js7caPhd7ZpLLX/jlfUTUJjQhBPzsrqagRhWVn2tpZFXT+
D9kTiMrH8A6CUJIoP4DFzW6YyiPhme0zrbwCoyagGsBQjhNeDuevB7wRyERiglq1bujOEVtJ+zHd
VtSlT04m1t8hX6GUb+vQRAqDfUJd67qSRoLxo5cMMtC4p0Oh69w4AQMKQuHDmB9/Qz3n/DOOinvM
jARY9kKuQaAPGCNckt4U08dpU6ndDsrdf+bi8qOG1aB6qxhFv5acXfLsa+KRysnMJWJVCA3Cncuj
nD/OJm8Y7dIVq/E39FyAZmV/kKrG7wVmwTxI9mpTNeIRPdYuqSk2+JkORDsMtfyZ+hxYJHhr3fCJ
cks+kNTrUERYRkyfB6MP7RggINWXlpZsnghhfKYcxdpzaXbYXF/xoPl6P2gwe4HR52hse93BYHvb
zcXXMeTwFpSLNO4X7vW+06Tlry745gmgIqFoMHDSYoRURvcCyJy/X4rmesyfctgMqVUvfCbhp4Nn
FcjJRMLMiWq9V3SXRfr7e/MTh01qBtJFTj2tfr/+mLHzTngplvTwqDaoRYjWtFuUrqZJHmrmZ8KY
aKTgsHesF4rIYPRDeOwF8AvonULLDImu/lUZgfebxbZMapxnvJZp3w1VL/Pt2vnUZ7opevBLm4Id
RbbPFY2jHx9wboBTaB1lIj8PWTIohGEzA24sYU/TGxfViod+IuOSeAyCT23bc+W/eD64bLIBe+0w
v4SWSFyhPsL2imnZ7EvjuCIaslpz+u1w33a+ca7qDKflg2+79tpXYETs9PAH076rfzCwpLZmIoN7
V2MBHUDdAVQLwQy8Q0qxk/Jmi8dq6obhYbINaD7mBZ+o3bNrpSo0upBNNQG78EsCIkBoK7wow3mJ
riQgd17Lahq68724HDMWKUyKKpPogKNP7dFkQ8Z4+/4IOosFGHrXc58VPtBFZTBI7bibmEZQSEx/
zjEgkvWCU4hB5uUT9seLvKMNlHBOtbFiU/F066X8t6eqWe2xkOXuVEop3/HTH5AVV4tNBSreGkq3
6ElTPKtMOuA1hATSt5qJ5qaIvlTDogdU9Re6/P8TfBGSThR4xGY3HA0CqAJJ5wiyNOvO1SloPEU9
jSrXkDvC8xlKuUmqJNN9mcMPv2iF3dXk+b7vBsNnF10B4kouT6hBAfraV+3c1RnQpFfwFyTA7n2v
c4qapu7UcjAwI49jFKL7v29aqyjlb9YEcxHugZBLSwrCWwnnedMcuiP3wYIjuXhp1Wqx7pILKs+P
2bis8kSnSZdtB/OAgOBoIkg4BlqwOqqzWs6DNyR9C1tQzd1HvydrY81c5ojc2SHyCGtly9dJZG/w
DcK5LYsp0rHWJv3hRQ3ItcpZOOZ/uEVt3nmm+sS9Y1SPE5luVZeRQXe8mbklj4VGEgDWORELjlDU
O0aQFmPVwNrbvq4Ch2zxccvw6nxmT8ZPq3W/YdyM9D9Tje4CL984LJAzHSTafmBd3bUwM4eh3Fa3
gb1LQ/2DEb7UX/Ugzo2r7H1DxGbogdBOU402w5f5xQGT0MF5ZAeGBjodfhpwMc27qo9cexe30SwB
+qALzbE9qtRE4l3OpKXJULXH+T77rJWSwe8tgWrUVdKBSub7q0QObW1VDueUxwOt/AQTpT/TJHxn
e3bIUjudni9gHmlN3AFt+HcsiroDZbHJELw3BtBQZ+e+TMM3EeLM8G1vNax9+exLP4CzRmUlo8ps
e/Yn7miZxOFcBOc536f8pbstCaEyWsXef7ocBbaipINNsur+LgFgbuZn+b3Mu99GNkO+HPDB9WDT
pOMQlRKoonHrY5siRxHooGxdzz/4FRMOJsU8RD/urMmw59InzDOwyBkvVLe0WlYHJUklWAgUifST
ABd3/BT/xKdiuclNHYGp9L/Pg+EXC/kqjb3rSPFM+PVeSamV6Muc7mjgw9QZmWXXzUgDGDF6kLdR
xbHFQ1YhTJv50kXcN/l3BHaDEcQd/Sbg0MouF0fqA2TTOhMXFFe3GEF1oMMX7r9RDYeXCtkOeFWY
iD1ykepTnLyu/PMRybpL2lGqBnQgo+lmZZDBEk1Ay144p8wBi5PUR+FS8DlE1uCoZTqlzwGVwN1H
sRWx9gHrk1EkPNI4bp2pQTr2M1e6FjI0c0W/rDCOpJAktcWBjKYRrn5GA+4o2juNLGzBIPX7Slt2
+tFum0DdlGbV0g5Ob5aSc2c3uRrFLk+52YJERA02dpIGMqk0A32C9LrB2bjT42gJ5QsfoPS/lIQF
3fN9Uq9fTLNug8n4sedJEiM3G7jJm2bplml/aUKfNkVUFYE8BzgzPuvnls+urX36BfGqKjimWS66
80Zo6CbUUNzT6uvjQHBo3OEqZb7ETINp5uYZPe4UsLZ99yYkCqV5pALQZ39VU5cohjlLw5x6P+e3
Tvw5YXk+ibOB1d18TerxK8zQN80zGDW1Psub9Vmygsa5+LhoYxkmaJ6fMhdEJxeKwHApr/MU4eGn
56DofVfXyQFui8HPglhkSTbpKXjQIaYvt7OyBC2GivS+/UoYEh46sK9UUFcYDu/XMhzumL1tA9Nz
3lMxS3Ys85kYTBM1frhwcHdWYboHXVoYBhUs3dAZtVQ5uBxtfhblOUhVUXfsBkKlIBdjr5qtJyOV
25zaIEFP37VkO5Of+FeHT4H6tJSyf89WkY6rRlqAprJ1YGFU+rkChdMmEH9ZtkJNvZMu2jZbi0uR
6yIdWY0lHfLPxNuoTiIN6P4i/wXfgowRoknCEk3b+pqnynKdkopQwvNGsNvv3Sw+6Nm/KI1I20oX
GebsbjJbpb9oAzTixya4b/ICHWq2m7NGXafV25hWeL3w0aZnO66VmPIJwate/iAZGd/0GtMt/wQ3
+EWE+Gf938xqc0bR1b7s2BksX2fcogcgGIhIYZdms2MqeCGczylTXl/pxqY5pvV/ExOkCyNCQlZI
0NjMkOJB+PYD+o9g62M8umbZkXsdLmI/Kt2YfjrCLXd5J96T8NjFjvQC8duBqOaB1bn5OzT5GAI3
AUpI4W6ouM+W/JtJPFtCnbHN/2EkEKufuEMKAp3ME6c6w+fgF+oWmyhyC2LgPesc9b528gGR3K+c
bdut9puYKQL38nDmQshXlHX2Y4ZjKKOd0Kk/CboDAhszRbqZy5UXmtMiw59UlFf/DX8+w0C+jMdW
0iYriJ2xRb4opZQXUwZbviv+g9wVpPaIkKoJqvRFVuyoYi7nCCmkhRocvl/4TqRx3UZXzHrSAOGn
TYLDOMqiWEupJjv4Xu0bXcAm3zQ5Jx+Lm8r4n3cF/MJ1oueIJKzAjQrOE2Txow2tYEwnYMiN1nu0
Cvkqtsp9iaYwSIfSio2U32lMeZvxoEH+dM/mTUWFUAvt2ioIAz7VeJ7Y5krKj+wZhmHApJW4hs//
II3aN0/4HHC0nQs6/cEGaGlphUCf4IEkj3Bpf2VIQiD9fwQDe63VSCjAfWicV7azZ1a+gHGL4ZBI
mr+lF6zPzEAAUEV/WFutQUvH3BUgTZlwdVFd+dtIawlDBLM0ZqBMYcEPneuGPFGJDEPdX+2XELww
+cDX1RMuDMAw3oQNEKIcrW9MD9ji4JTqMoJjCpdChReYG6bin/x9gfIHt3iKsZJalppo5OH7BcRm
na0yyqFIUv3dUd6C2ojhWR80WSEDxsM3bL8wxYQ/69Kfoxyc64dLGuCQS2CHHBXZp/YuPx57IRWP
Ga0PVn+MBY6ktXjvoc6Ta7T5EPkil7ubFDLJPyhnR9rRqylVKNQT78kzcn32MfYWj2ZHFM0c0x5G
jBNDq9AsWBiF5GUxeNGSNlS+Be34ui8T4ciGmiy0E0WXX3pL8iMgspwFpDyxnLUHiCUmnOU8493e
L92s4iDFnoNrOcK58CAxW1893mbtwcJT86/mNRtSjtXv6/GO1rdBCKwWQ8oKWPpt0hW4LfWpHbKr
h8T4RBiUl93vJK2tVM4RUshmqTE9u3sMw9/RteUDfk33RBlEbzQRlPgCGfNpn8qMnW2zruCb/ZJU
ReZNmFqGiTmVEA0J8LbyG4rZwvfFa5Fs6+W8yaQsyQpV4AYwU4UULvATSc9IgpBEn7BAAHvVQZjf
lS8BekaYVHtDDfqSOoR7hFeNeH5oyEg/qGnaUjT3wFH/e9j7mH2LAufQTPuirNj6n5a4oOoZWM0S
b/CJ8sZ91Rg8zoF3z2c45BbyNq6azCElrS606egGfYjFBeSrxPOedGpeIZP0QmoTiRBHRP2wAjHG
MIeDKwT0u/GYjSenSCMbMj0HgUQuNKINQY+bDuAUDWMvkjbVYtNuUGD7MDc/SzNtHWbQre/LUQHl
UaPkD8IllFlWihnL9emIyzaEr2xe5U/i98+TALhDNX/vVuGtoAfyUW7Qza04/ezriqLZTlwWf1qF
Qza8sFIPJP9t2STkIiCradNzuzHpWMEJURXyft4QVsOavC3FH0AsZFkcoydR1OftaL9CVpgNNXKH
9B6EdU0MfQXn9Ex6kseceHBUW+Szy85z5pCY817aDU5KSInMwCjOmZ43U2YeKV17Ox5wmppml8Y3
XsSxDCITg8s30OKWY9pd4kcByXWdxXJOtH2wT1bOZlsQ/f1RUII+8ut+2lYq7n92vZKpzrYMym9c
UHhpMCA+GWT1rP+xnF2E0eLuIW59N89bsiqez47PrlxlcEUFko5b7nxR/oYcJeGVTkSQbEc9tDL0
4PUE3tVYi/INVr07iZjhxhb4axQ3sTMYKdHUGCMkrWjsGxZ/iQC+pZ6SoPd+aoBK+XhHZxaP8pAi
9Y84Ctigds65QMjSaWpdcX3l0We9bkJcffgWn/aHkUwLIRjx9v3DfuskCOAfU4kJ+k5x5106Iofh
OYPuzTsgC9LfkExt1zAtW3k9YzLEJzzcPiS9n9dghJE79140cb4BsmEzPgf/oigEh/UJL4bGzEFJ
3wma4rrL10gO07no1q5u/l2RKZbkGlLuH7dfnHUIO9zgmXGSkYmzZCbDRnR1xIRvZDHRxWCxuLIm
Wdk2DOTaVXm18aTOkeD1RdD3I+C+9XTsncyqTdr+6rP2KMI6AGAaabJ+D+IV5grpVOUbUcx2PI60
nCf4mWeKhyWymPJR5wJj08+SnsKw4SVrwq9l1pwNbExqFQRdMpV7qI14XdT8bLS1TPW3bAzai1yR
FOqjp1VEWZ5IGQ742HM2YpMvXpwXslhGsMpDfPtwHjBspHS+3nhsjNIjGkUfzoI+n1DuigBsmbNc
zUf3pJSW6oL0XdrIwzWJcrGc4MG1tD5WUitGFGp6CynaMsefwgfTWx835mYiWqs97pLB9SIWDpm3
cxlTRDElHc9dpzIZCXFRA9x6MNVu/+ssUgIDjGO1PyR8aGb4U+U2kcgFZ3f3gKPsPm8a5jro2z/B
fwJ6E8LaAH9H+ZNg3RKoS5ttslOosLUvp4Ed9cyzOmNVF+erpOJeDDvw56vimVMZocdRcxGuygVC
6XzOVRazqNqyutBH0gzG87GpQLR7Pu1HVlLMn061eJA+3K6XMCLNZ4DjDr+VN/lppXgdG2KsGcc0
W7x54q1wtzZR+mgpwAg+oxS7wD1aHvqTC6iV3CIMxmBsceRokf+MoPhIBEMiQSAqEP92saG+K3VA
DZ6p+/60/aWmwS0otyBIXymhL1E8BIP6yp2KjyAYNrR7euApgV2S8Z9erAzBVbMXPQdyQUvaKcGx
bakD5o7H4rEGxsVyuyEh7SPqISQogscf6Dq4mab9nHmXWmkh79AH1qFSC4b35zEr8mAp19Ni3cF5
W8c1eMvXJBDVk66puV9crqdRbwLM1+i6SmT5s9HFu50Su5Gzp3eokBaQ01HDEJkSSoUGMbmsSkk6
zZoG30MnGzayyh8K+yE057yXuvn5rwiKvtyKSJ4iU9X5nx0XsmOTEo8H/WTrDWpyacvZgKFHNhui
aaypHs0IVzGU4kfV36OoIa2V3UKYgnARF0B20/tEnCARR5pDvys80YF8709OVAtijFOFWz0Kprrg
bRqcH6IEYyEmGIQxVRDSjBqaNUOx5Dy5vwDVHlTBQplTF1ZbfOwrCf/9GNJazrhkkuGsNpEVg0+l
zWnfnNS5QxJaNbEZN/LGZmCN2bBNkXJCc8+hjLQWf6vgL3aGDszKfZd5ZDrK09FnTkvZaCVddtOp
y3msUVT6h6xTfXMxGSGJMqm2qSLc3lUYJcc7OHcG5tBHQUHquamVdAXHYVo2y5Wq/FLN5PeawlkP
nK2Mmr7+xt4oE+N8gXbHc+QYKb2SvW3KsjrWsPd0Po+YhjuqxGyEgtJue2sAE9uwGlyaCgMuQTdp
8FXJb4XpESGv06YXEdC+6aN1pCVq6qv+B78k6/ufVJ77aX3QEIjfTDR6wzMgIgWS+WniIl+or+Vk
yiCZU+31gSewtkUtzp7WIeSi3ieskolzXkLUzjNgwLXlHZ+uawNpPAUh09rgP02Dq/hn8+fEp1OJ
1K5FeKjlewOvMCA0DCmVAElJfkXIgjR99ur0L4snUNcN2v+U282Gl8I1pyBGoI0XP/sJzY9ZL+FI
E5VTUd8EFo1Kccl5c+lRGm5JDPINdkdX9rVO+j++514Hi1Od9NFCAWawYlEHBWlsbv5ybfgUyxXy
M47Czlw8e67yzjgjf1Fu7EFyuAKxkvKci4YgNd9n4dTLhpKoSweu9CI5hdFBPVES7yjgGE/GNdul
nN06e3opOCVgmWMZtXt+8LL4PyWqc9EIYvnjXq1kh4fkKHOgmLFuLFl1PSshTAB/iRup9ctxi9jU
J6JdwPv0+1i8063dXZxt0wVbvcr/GDuOcZSh2qQM/Mq2qy7jFb/VAVATHxlCn21CKT95W0oqaMwy
pRq942IhIY/rVl8y+u94X2D8T3jmilNd0TCGmsVosNbujf4gDh1Igu9DtziEaoeMV8YUaDA7F624
G312Im2yHSoNkO3TnF8CoCUDzU385OwOIfsvqeU4c+2pgbMaBIb8bwDKott0CgonQgKzhqL2MbBr
CZtEBshMJTUupBaz5UH0BGejxwIRiXrBffXMcXATRr0UVApsz7dQXJHRAAHTqfKngfYhryf3GyP9
zg6FIlvSi4CfVxvTBmVh02MaJNNt3MvLvGBjx1B83mo6/fCsVaXIZyYlogX0uH/aOQagRMH/zXfH
lJGRLGNxB61q0hsZ3oVlI+fjiM5yyPExfGPEokpCI7QuLh7Qjw5WY78u4xgy/IlrQBjlm6/ONceM
jwr+vbqGdB9/uoZWOW8ZbNx6pNXzO3IGvizZ+gSw7xRqQ6i4i8sXPvti0wBaWxKQY97CEzljHSTj
cmMRnEFlHY4nEY5BE/zo9+qObltO+v6a/Xxiqh/xMmIG9FSTjJBjBHaKXqSO7htShH4OW9O9ONB0
pcUTUrc0blLOvhz5Daq1dx/TfjSKOxEksNh3r0h+sgg6pjZNxdZJD1Ra9+9nB/fahtnC9acZP2JH
vTlfnCFe5FZgtwA9G35hyhskziDByFoUDn8zFFgOS+oOz7+OTz87HnxluMRiJkT5fmEnBTToWe5J
AYVb1SU/yJ/KNO6wReQZiQWzsO7tJm7OYEqLm1j6rlp5ZKHIDLbOJ0xjztV6eFifPt77S3uTIW7O
pC7C9LJ9sgz9qZsFYQQMpk86DSoOqo9bxx2UODUOxxAYOUIKlaC9105IsUMqTRjo4QJ+wroY2/+C
g4WO5nr80ud6IHYxDJsWKNj3zT1WlR8PrRUAekuBtrRHZ1ThJQPC9jZewI1wrvRT1n5jki7Bajg+
bcpWu95ppc9sKCXLhlP3C5g44uS1R0Iv+6nfp7CRU8hvDdh8c6emjOsb/yDEOM7EFDIZ4qszxWJn
F5K+a+1OxdszFXt9f0E6vPrxeWKw4nDdESOHH99DqT3GO2YI8fDDIOQuII1m/cJA7yUapgNQPzg0
giSXaH8QTSdSVbPL8Am1zMWeP0Be7E2xBwSKDLBceoBUmcK7GLPqiC2mT5SL6woqFUALlm8fD9pO
ZnvgzF7m7AC4D4dHAoXbC/bcaxYmOa4rXAM3mmNxCL2ztJjZ7j9x7weIitP9ED0SOcMi/s2gFWYE
iXJOyGX1uIwmS3nYELzlLF2a94hiFWlHbrPaxvyLijppUg1/HvhVhDM77j/Xj9UELeF+NXgeELWN
+Yh21jElOUSdFCJDp2o1FrS3xBNZh4Ist9fGAq48GgkOqRpsXaERN8xlUpbs9dlpX71ldcElXZP9
vFcAop0RrhL1WzpQS18UtOj8g/ht6hKDOcEsgoIeThqgjtEjE1s3z6VgazH1IJdF+hCiHqQC2dGw
iJGPviUYMBWMjk6p+f/pkyig/3Yau1makFhqjy1TJuptV6An7O9DN6/BEpBccZOWiWuZWZVQoRe5
F9td1TSy+V6b+2ZPoCJlhd62iF+UZ7FXtYou+rjL5c9B8/3D1YLbluZldnG8jryGiFkpRPO73o9X
ZO2zepldUbzUQoBnj1Un6m/N9vp1wDAXpw5pfu/cxSQ5oQNppRD/FzvzKarQFvHXhaah0dhi3fw5
KqWBt76rV8shg+TYWvp+zzz/sB6VeaqVAWB3xzvarmS9nRo4Oa8lCBDaDMejxV7hk29dFK11uclN
ddad1FiDKL52dk/VwUSxXHTQaF2LWbAL0Zlrvv5sgVn1D76VF3rT8hqVdWN2SGRuxEFfNDqU+/r2
dd3QYrS65aDvj60/R/yF2qyJC8Ll2fYs9UbRsG7rjiaULrPXqu8YpE9TVBXLcom6gMUmvnqHTQeD
8Tse/O8Ob7F0sGhVJakOGV2gKB7jvzOKtWyEVPQoW9qIhUZm0Yq3KJ38gnKVlt8TR6zjcN4Nhbxc
EdsYoXogGkAGEeN7GFroVO/k2qEvbeSCpFE5/qjRSYOk7jgj+gk1YzV63oB0dAx4a4W1GO6urDW7
jOE1hIdvTjoQn623wfqDUsYBgb2DqFOzHR1jYz0zeVlJtAAKydaiQJPFGTx7EP8SnkOgs+1SPAlj
GH69CedrB0+Xaomz3vlv600Ssm/XykZVMJ89gjGjrKtgTiwQf3f6qfd6gDxUJa7dXvfg3t+4mMv8
yWQ0Iqv1BT4TIN+4ocPNEZJIPPKx+lXTleMTMuFDNeeAzQRDQ632CJAWqhj/wGltVdX8WT5HTh3F
yMU5ZENOdR2oyEXpqRivduAfT2BxlSUODEqfAq5Q9bG3F0p66BMtUTNqJknk6ZfeMqHuXWcXi0og
B18kNS6BVfgX9eDTazUuTn5icVkFJXer8owML7SkaRjDeCk+SVgqhFzJrxWRGQkY/cFpqxkygbSv
aZtI/FDxl9NIrGDJVublv1/ws+2YPnEIVXpNSq03J5jBz/sp1RTjAH5LoYOU+5cydkoo1/uo4ytS
WaMbM+yKJFfjpe6E1E1ujr6jXSegBylO/SR3e7LZLryVdNAWGyNI5IZEii9dZ1LodFBX041jMbpc
64I6RploxaU7yFhYOyMbkHLJcFkYZh8AAwTgvtZGKRshMZQITOEYjQuDreYklk1emHMmNaUoQdQY
QCn5/wN7n5TgDI2PrWUcjpgkhVNxlN7kr5x94aEj2Bm1HPE139/H9D5inhY60egxK3D5vv/5Ingg
1le5RnIR/SvOV2EVMPTgdmXZvkYwitlJmOeEyN/TJoerAB/8HAIGyxKVWyivN8oVaNTDLfByvsIk
FQIaTL6PQxnp89yxGImjmXohjQoBiPO2XHi/K9AjjbMDKj6LGdy1lj6SyVZB6jNT+duHy44PVmEx
XPmVCwmuhl6YVWdtvkNHczcmSGb3+nhh+YI4k/M8aa4YGz6pfifRca1STIT4mWhXYANUnm9+pHj9
N0FAYs9u0sEn/s5dzXEfE80079yrkydWriM+7JcCi4B8fj4NER3PEx+7LOSaMePMLSS9xmFCnoMc
XES9G+ROt2lR9cpZxG77sLjoc5IJUjSuxb62tiN1UyJZdBcQ0krf7yluTXKrapo/ss3aLzDS9Z/Q
Y4eByfb8It3cuOsACGPQZsO1qrLgBLgMxzijV/dA1/l1+zXaoX0hDv6jATgx5XQawkvAvV0SZBuQ
0i2GBQ8M2OirJyuS3kf9JPWTIFeEsfEMIaa9KjlBbGkF0rQ7galSDw8//oaaa42rabGc9vojOEOs
sAW4gNNwM7e9tBAwnM1DD7DdsCWo0pB22vPTCZj4FD02JuZp9NpPUmGGSutQBCbuZ4CbqMqGQomZ
r5eoqX13miJC2Pim9FngNQIyOrvUvQ2IdoxSrpVwG2s8P24hRdC9RsBrJUriqKtCJqnIeVDb4o/S
Gv7RahVe910prftgTe6g4q6BFh7MAOQPJyllV1WNIQr2Cf1qyXFrs/ihpkVvSJLCFhHzOwwse/e9
Bw5rOdDKoTpPMXiZQ4lGSGPd6JDQqDC0xLomTOYwhnzLV7IkEQE3aRnhf9ZW1gfsElzwjVu0uoKd
TCwpUiVIYnCi7qr8QgJWmvFRu1G9PAhQyAq2u+eaU/SD4GUgHTTRyFZV2fsvMDt5GjqEh4nIuVG6
g2ErALO+stfpfIV/IFl742TbGAJhXs/RK0kbEM1z6UQiMIrOBgtfcHU/+e10oq3zgYX66EY9Njnp
T795jGyxscQvsTH8dIVLmTxdzbknW1zOhmh+FsnoEfE2Lwl16fZoP+s98oCm+S6eaRwvUYPg6BS1
HO3kWvTqNWitWX2bXV9kWNXPDmcDquLePQMyLiH16eiPaUWuBahWWBxs6+hjjMokDWahmrt6R5l6
c89HT16KFMO6OLJRYCb+WjswGC3AGGGBQHcp4Y90C199aD13nUN0F27VWv+IeCk6diRdGE5NORyn
BM0skt3y+V4i8hVriMtvZ6BaaQQJQJgiY/xMIXLbjneiSTnP6WL/QYCuQ9ENR4ZLDYqXhIbVpisn
Iw+PjsYstTCVuiwNQDCQRiAyQ7+jyraalZ1wK2ZNzcf/0LFTO1YNTapzPRp16ZFTK6YnGsceXOwL
xSzgyivwCb5P6FfxGUD9ExlQZxt3/nn62jW6Vp/fJZRYd0Mg3AqEH6T489yMRkEUepT4XO729+V9
r+qWF8XEsnkn0DgA1YLsdwADU7WDR8Ru12cxhialOJF3ixBIyGTo7HDBZy0fezPtWucWh0xomIgH
JlXY6YZDBbnZ6afmUv0Aq2V+CQXHyEoQNzLK8HnuE8zkC9TcEnl75UA97O6ZKSwy2PLLKj4Svbvg
FCg44O66/pjORKrYzzSnEg3l1Xb53Ps6xmo0SK3rRWupzpJqUQ1vNibB2JOqJ7nlvyUzJy+NbXZ+
tdm1wUhzymCGLqn0eKbNsrOJHysF0y4LiiLTKN5bPF/6SYKBldFzf244owJ1fF/ExNJlHl0wCfXr
6CXz/W2xbeeOLt00t4BeayOojUsKFYUgVaeRsgGQ5WRlfMsgj27t4RIiyHWR5vizN9PSRQcwfUdi
RFmQ+hrvPcvpfG2594sGgItMdI2tE3jyaxQP69VM+iA/1sjuvwyb4Y6cFkqpt/47z5CRdUcxKyNk
5BxG5+qi3Sx20cakalsjRToHpRi0EAUxvY2Y/qHQtVG6g033lmhckhtCg+tFdoLekqVdQVDwZxXf
U/wceLkafWjKtPUX//8GKWI+M41n8MjGmdvEhoIFDpruZHyJgCypyVg83NQi0KkKTa7oWZQAvllP
MbP7IEgM4h03Xvb2FfUTATC1IViD3CUg9vfAEZXnzaHapoxvF6T2k6pH83ga1lBgoWhY9h3H6Pco
t0Z3ZhEw2RL78E0jNp/IbjOXWVM3YBJNx4hWqHe2WTAoiYOg4AA1GQYU53Cjq48TQBmBwsXqtJuT
vTBZAtdlAxfZtDePiSeHWLEMoloM5Sf2kz5uR1W2nRK3HmeFPzK8boB7do1vVqfQb/PqOxx1TewU
1j0vQT8IQfTrTS6WJ/7hq/42y1Z1T7FuxPGiu3ZmPBpUEBwvJ5sSLmvsKPNg/OGZgrvvOA7A/TD5
yn4TBBx14nHgwcnHe65NP8/1kbpks/CXSyhJMlbEUJArSflWgBJJQdPZgZteQmHXHd83SHJNsev0
eQ/NF9r7Nfs2EvP76afCue3/QQ1j3iFauLltzx/VRM9cq2pqV6FLAcYvg2N4a0On1t0ejiiGG2Co
YFetCed0FgBf+SwLDr0kiFyLZB27RQLPBzxKG6jMdh1xykiLt2IgjbnS0JNyxiWdJ1WkvTUMSVIt
XvUO1C359mbxRD6a6vcBQdgo6xBgnOufgaC8ccTa1a1y1f24LTLwEpha+wGfCiI7WpSIfTiB73bk
Lz5goKBRTM/bYiBD8y/gbl7CIVeoaUfC9xq8U8rtUPPPDKLDKzugIfjzzd6iJJaHQZKP2uDYKRZp
/oarDPXyOkIvcLgMvnatG/bn+5gkMr9KlYAXExd/RRiy+T8L2KsRFzoVa917t5agHNerQt2sTnDd
LUzAHp4B4u83q0tSw513+k2imJmxAuoQmraaWQbi3Pry2qzcH/dWpzAsPOy2DCJCIkQqS3lEWYR4
0wRYystYDMcfWoA5LGT34MUaTVAG0gIOnM3dFCxXmT3I9KwmdjVyhm52pdBv9WaqYQ9HMbfqAzoe
rAgYymN1CIpI3/K0l2TDtDcWM/l+KahXEwXNEcmnKoiBJgbzEhCE04puVLnkCMFKdVDOMugrOBRY
sYP8Xh6wMOL9DhUDslRxzFwoEbTEegvxV907Nasv4uH4SQ+wBnxahIuS5KqNYKW8Nml1ZIV4tLcD
wmjbS0cjbClbpu56/kaU0S1BVpu5MRjoOp0OcHsJJXo7ioSxT8VJR/kLSe9pnpPN0o5QXQ1GIEu4
m5So+oUJw0S3vkQUeIkAyl8iSBEI7xGMtSdjkhkmt+Hy1DzOl/IrXf2h50DMik0TUfqlFGGfQ9Qv
3pSMSanJPH+873br9twOwH2MSSO+4W5RCUkBK8vTi18+EJs9sSPaN+lyrZjvMyBalgWvnugOJnbK
WuBqgK21rXYfvy0JVKSQAge0mIURlRF98m0iByjKbARczHOVaFX8v2NaNOYU8reiHTy1Vg0aA2RO
SYKGcLgXnz+JOn3gArH/mBc0yHZna7w4DXiOMRUnMTegNl8hT9U+513mua1J5TWPR29AvhgqnhVQ
9QAXGxCDLqfJi3Xrm+GRG84uaA1linPB8VOsRysJZ276QYPtbw48kUBVN9X3z5d4oVPO7GG9hylB
OI+fvqeZ32D/S+NAOia9SEYp1MaZyhRhpZBCpUfAC3WQUItWbcxtXtgqwFQtb6HOdC+uWx36QpTl
6Gi8nS8x9fWpar4qe7ga5C6tgtahyQif7HCghyrChgUcLk1e8KEWZ3y3bSCBh08a+GwZrG5HShnn
E42rSYpmJ7ho6WHU9Ub6Hm7PfdAHrIXr20ljw3IY8/axYtUG99kh4nibHH+YTgnEiltWtG+mLXB6
Z1/PaC3PtaAM/N6cf4QAKOBNQuVQXrsVJJJVkvHHF2DRxiLhuufR24q59IxKgMS5G18gD+lNeWH8
ebCg6suHhmeTV9a+fLDBzyHt0zjj9FWRRCHTRAhNEL4+WgJg4bdldrPICOD7/UedX2ECAfccY7Vv
J5h2KBVvDUa0+37sqIduKFTcd1qfBoN2aSuSUofngKcMJmOwh43UcVMIKDTdegH1ql2RH6G26GjI
Ahm+BtMUaqQM1mYOUm0rgmv5XxJAwyBmK6B49b73cB/qGP9rtURpWr6thWOvndxlugosUbxZVnpa
fm3FRN5RunKwIBvi1UXwEmbEtFsEtBzFSxbFBYwa8jqESZgjXs8L9INYQOHb4fYwFD1RHDVb1o4O
1RvsktnLL1lAL1u157tE67eefFLtqw9n9vIt1zl7LNthNMkzjMqXoLOt+TVkYrPNXyPi1VPS4S75
UlZC+icknyWqHrwjzOLSbC+uP9iSDB3y1S5Vdvr9LWrRlbpcalwW2pnO8GrCgfAgmbpI8SVjTtO1
4/AtoNDytdL0e1icxUwfnMqpOBNy9RbAHARJtedumZHe8ZEP/MYRXTS3Jm9Ts2fiXh6ZjyfxgEkC
j67Luw+5E9bqMUP+nOaSYlyPVrerKbtRKKpR1+uXUq+aMwvSJu+LK7xvlM3z0sEre+z+Qmmao6Vm
agwZfWp96m311+oFC9AwX9tvCthVOl0OFjTTU7rkAvTpidLOYjTI3slwsXh1DDbtNYEMzsX0kst7
bN3y+iJVbtHDgiYsK0Ndb3v/DlFT8LkJnqVNXxbDol4NMt4f5vEqeR/bAqQHqPnL/szi0ygHX4n3
K1UdrBcrcgOgbxyu2xY+EtfyYcsSmTF+QtJr5zTJucoZEvm9s3johe1lYVkETjjI14Dwlb9setlS
ZqZfZMGBboEH7gTCBdH/BR2WszjVuQYSZziW+nY/6IeBwMzC/f6a4H5CYVcdOkKcouRpCFzlcK0k
e17r64A3RFcOzUvqZjCcs4U/DwRkO49yzqf9n5tnNjWiRXv8OpffQeMR/sVWRzD7rESCVkoOkrD3
NmqcLFUD0Ro8CIOo2sCOSpI7V77q8FkkZjAEbMJfzPEtFEnYr39tCX1IkIPD1jw4twHolRBhdSld
09VDtnunsBy9nOc4RONSnVVFxHCoYHur/0foH8Uez4R1ZPHbfkTXvLyDaSP5qGBoaDeWIvsBxO+a
KCOyGx6yiU5+v6zsVTxdeIpyj3ItQWFXxh4xUmjbIMRxouVqnOoqP7p+1AomZ/Mp5zMp2sAbbPar
glSPjUnmb7Nyg81uRHH35TXAFHirQirLrwRZ734cKjoZMD+cc7TBQN6wz4w8MyCZcg9+fc7Nmk/z
UbOCgR+plBEIKUirI3ecaZt/CgfO/gYFTy5Dn/29+3t13rxGHH2Ln0akxViRm843A5Fbmmtz+HqD
acKL/y65Euq/VXyJhFkwwszCaAUg+GGZy6d23qiCgCWGkiqAPEd/x9LDEirR/cSyAqpu6mnUdKox
xdMcu3yHwxvr3y29bwyJvJjmSVOY5yOZlcsf465PUAHZeR/B5o3FSnCntlkQvZ5oYI5ueBlLk4uD
DX9XmK5U73foUWgzpBqoSwPMz3LE0pdpaWCVAkFlion1l98eI8JDWtH7Au/XhmspURFyRULgcfbH
OAM0v/9vzy68qpjGRKJ0FxJFnUWrdnHH87PgGJZPcta3i2fwwHilsbXtHboZmZmQYk3sslO3g8I2
NsJZ/dJcm4vbt8ododBpgNIAgHmp/LRczvMgME6FB6WW88PqGLfHUf5MjHtTcFgBGzgiFxCGJ+An
+sUN1KiYMPgYrwrQk+9rBiopH8mfZwtirXmQ63yjKRi7Mnkmr5HMChpntG1oeZ8iyDHIQPvixbU/
s48G5b/f9LGtjqAc3BiFt6fccSP/+EgX2OhIrSl37bB2ZRzTkrd4Desf78a6Ef4Jk27okFM20BK2
cZGylv86h6NNzubIWa1jNhqhi52rcb49CAWsSLaNJ3Jwd9dKwXQAFP/ryWmBw83ejKOACWe9FNJC
SQHgfT3BHr+KxC5lQD7F3hjegdlfqs/BaDo89/UGWkMiU+JlpR6enWlbcTJVuaoeh4+i4JrYjwEB
3qyS1+E3qmjm9YyR5cSWKIsxsnj6WTMTfGkJkGqLA/05JaMqRK9ZNrAcQDY9FBLfnEj3gnNjs9sR
aR8FfkV1MObY6tsBe+cSd8pFVDgzxRrIp+MDOvLV+oLfJmjZ8p+1JYM1s+bB4fpzs9jQnUxNxMVb
eXSamX+dEF8FRDKkePlpaTcxJUuK7dZ1cT+KqEAwOoXcvUB1+5+SlOYcx7uhzJTRnTXehuRoW/Gu
znr5OXZJEcT2MtfLSvqJV47SQax0UTjBQ4cA/nOu9XoonzwL/L9GUmyJyhI5MIhiJDXvuzSd+Bh2
GIfaVVQSpt5zQrTa346gIjgGP6RkgdU+riuHMRlHgTwIZbIU2VI/PrMAUaWpPi4Jqx5mMgB59gZ1
7OBojB5qx8KppoDEcUIvysj7Uhl6STWOWk3f2IsTIDbAzXyGXO2yPgvakfg212/f9X1S+komZOkB
SkV96PtD8jvQPPCcFjqHW7X3GMci2voChKHg1otDJHF6FAJ5AJE46IPoRgt+9HX+Wmx7sYH5yN5R
ZSgixB+xVjpIuw5agbCbniHiEOiTBFDqkUxTHuuKU7pZkpC3QeIgLFxW5b5RyiTw14yw4bVcmtBx
EkPMtaPh43mcnnleQmXoxlX3gsgVuxkjpAwFB0fFOKBm+c0auQhlxmvaGePo+8fqhV+VAQL5vj0u
rtOEBWwdXbiAnREQtrxlOUKysaz0CPzF4TmpT+ubcK8RhMCzVhETssp2GPvrdT+AVbEK0JuC9Hb4
/lhSiORImeEh01nxVlggemAfRwszj7MK8Narz2oT2Y1Y1xGbk37xloELpEe/BJaADXgTPk4Vt/pM
duya1RM/eWsMNEr1mTVrVRNrVTwE87aNWMYIfS8REMpTK8D0jjpsFWemnu5xRRWfdSMsOEtLlk90
Wcod/GpjMAnw1lDgf/PyvYu47BLbmtpu1M75infa1AIjAMr8wCnH19E1EHQn2JahmZpIvCZR9mOv
wnQ91QPvzBJ7nUi/SwnQVFrlTlrrqL0tSqQdJMbr6azyeOLme3Z5aujVz6LBBiOK9aSDx90iQ8YG
szqQ40DSunw6DQbCbZeVCdRpHG0gqlRBriHcAqxR7cC86EW0SKziAf9IUH50X+cH/jN4nkGO5J3T
uKEVFcA/GxXcqZ6U9pwelj2n4BGTzIrsVE/8DfEKMOa8wXI9KMdKMSyTIgq2bDoCGn+T+UIAnndS
At+AnHX6HVwqdaWKlIcgqBy1AQ3Uj6cow2w3dUNiWTxJELrFLaMn/30O5zn1TyIdEGwfK3yo+9Gr
u+VXkXJepwjQet6hDOtr5+G0RkkcTafcfi7BgM53ayLZxlETTeMsGqadWLwYFHKGKqLOSMNReyp9
LSZ75EbF1k2PKy/H13BY12dy1EJhMTAVRJysYtZedlnqOjHTRAABxIoNChCBqEC1TSdTzOeQXh1G
/q4WfCLbnNZUTCPC2oDlBKrI/bTMeWvaRqhj2CV7ycpMY7BaDUlj6ZNY/gsCZjq1CqTgmiQyEYF0
BKlZG10AxtKn7X+FvsbSSisEi3WiEYVhYupmhPhEMfK+CsrwP/O8ZPliQQ517nQ24HG+drE6Ud5N
wcuw/9e6UfY1CNrF8/V2tH2zwDDKtgS8adiTSAF6Wlc6P7elxIpEVWFQyzOK/g7iNimF7GRls9Cm
Wnzlia901bfCLsE7NenSpl1xtSFbEVLVU5ZS6mJbifPus4pInBCf7Kqo1x4Adcsu3gsHf2AzSBoB
ttpGI1l1ze6pv/R/DngLIkb2y+ndU2KAUG1IA0Fe9hUu5U+a0HnFRrUWLc0eda0/mneaz0a6cpyN
hchE8LtV/2BcJxX8QBEPao8JJoQZDahCDUKsdUbDPDz99DNjSRSuONQgr5d+7VheFXswe7cnUnFG
M+glPPot7km7Afpiwd47BsRMZf8ygHkFTb1Au3nHh2yh02HwL4uR666Fn2Y37sLAwx8Tx3aHD4lq
IH4r3wh/nBHqREYVbCyVDaHkipmcXFPNfGxF7OZofOZMUDa3nqnixX9W+zY/eiSurgicH3fbwEMo
rmieTKCqyGvAlf3HBWHWwEESpJ1MmpokuqOflQRYDmyhG1ylNtPPyZKCAPa1qoicW7Al68Ic8ttk
ZigfSUhNoWD/z++EJ2HGSYLnMSj6ZhfVTV7BGkpZGHw/4R+irJrQvRjRhKh0VgckNFQFShZbVJ99
iyuRahj2hT4Fl+L/vRpNp+0ySmuynWHc7CROpPKNJU4fgLcQE94cBgjIUX4m6xShxxB5sgJR+Gzi
2TqxT5ufD0bI4uSWcfqApA48FRONuQ4Msz55eKxQSoh0Z3NFTlug2WZ9ZYMhM3ifZ6YcnTdFWbq3
peJ48llUF/NEpzZElNRotJxjwrpRUBK6I0slGRRSGHfCYSgrZtGjwu+fHEOqvoWh63P53dS4/VMJ
nfKm7YIwQpctwwfBNz55xU4HyRx8bV0PRJp+TI8TJwLuIXalZgdQT6e0vh6c5L5DJVvRL1Typwbp
AKqzyslXR7ixl4m531180tu1MRO31olmVtmE3bclmjysYiSI/cUcpM4kljyABug3ltWKth8s579u
BsY0pvwQeiUcVBUr3UEzWFulBKBURieniPo8EOowcAun1+SOmcB7yi+CR5LZM0CnUiQ60VwM1E5L
xuco2f9PYBA6vMNBjvbIIzANd5AQ4Jz8zM/0q9dUQA88JdYQh2XR47DUSHIO62/Ee4QxReuvjtgE
NM5yz+fTkIVoaye34pl3UTw1mSFt7sZgag6t6C5MRSy9ZQwI1TpSUpe+UyxW6hQl3CNsgO3vw5kj
gRYkfPzvuZX6wonRL7acXQCFaz0uAkr4kqWQJtKKM91tjQJjbBaVB66bfA0RpH0/MjvACqf85Ly8
JH+tQoRErFLaMdankntgaxgrEcIlG/lsLgkNNl85oqLQIqtw0IJffWAdve8+wmeP3q0q6Eq/YJxx
9QO1a5EVw4NV3XucOHfJ71bl2JoltCs4Wr98bCnLrfI9jiYjwgsCRdk6sLSDc8UrnDyVBp7Lqw4F
qwxkm9SvZbizPsqtsHiJCOY8J/09mH+MlXf20mRAPVwOorcfUMuhH7nH5ylrIveLdoeRuNf4u0K+
uRn4Kb4Fn8T+XRDcr+7BXbTpOp18WlS7k5dfagFLKJT5mo6aut6oKf7eVXWg188+q5S2UbiXi4gM
qyIxBQtX5ZWA5iPcCgtGZ3Grhhv7yYFBLddZkTrcYl1LRM8w98FK0ZhgXSyxLqTqj/j+11AtY543
mM+V1iyomLxoRiAGCzclb38IiHSbU//RW31u4npeAkjxz+hH5nXT1a7NCgmEspzR/0iG3Oyo9uSk
DTtDqAQzIRmT6CxGHOJxwWThzX0OKPy2AQTvhsM//ArgvIRu1f2xH4kaS2Ktpvt+RspQiO6K+46u
sZRwmErl0jZXlb5Ko9ZwgjCh1GWcXUWprg6PvSMF5oO44iJpiHVJw7PjK4JIrlvcgrh6mvVnzJvx
8ZvSrvI4JhrzKkqq681F8OQuBcHpHxeraeSaqoJOsRYU4qi1Q6jN20Lv/y342punSoDAcgzz2PhJ
b4O4/gP58OnJxMbs4AZqNjMAUdqjQWCrRL6IxYzo3fRMCD3QtNlKNWSHZTMWlEYm35QsADmMiD02
1J/AFEaAljd/HvVD25J7hFg5HeZa7qgnSwFfMwhx/aKuxowfPhWvQThBvwrPhOecyo5MhWPH7qTw
SKJ78V/N0GTM9j7vaTrHAbh9YmXQw5bZ2S1QHtOD2UmvCdSmS2lIDIFPR2lBs5XUaPEeMpzzZat9
TH1ws51oeMYu0DJn5d3iJkapi/Rm33xS77tw0zWw8FyszuiJU5SvlRTlmF8Drdr3cKkNB/f2McvD
lKeXzMy4R4o+Ales+z54MgZmTmVyEihS43qCNRtsrJJGrPbvhxrC0xt7n6utFCqGGVc6zEvRVZtf
OqClQpLTWyeEGOuwUn0l/a6AMHZNPGRnbD5unZ5VMTD8Rrx1hUDtH3Yy+dbfesgQ9/MOAXlvI/5e
ZPBC8mOcAGLq2kFAf1mHuKUsSFtSvXeClq/xWOFWibR2bofcTfcW/E/qfrX8dBbiq/IbwFAARL/z
Oz8r6vSfeFhDrblbDEUU9XmzcaR6Wo19ZFtOIYj2Q2RenBVe0kDJaOb6DdNOm3rvdgY2koOfCa0O
pPGDDI06j29A71iIZwtHN2hyia1IkCl3jw/Eb2C20Ys1oivQ8Zu+bcJ0ge6CySoStNViEBOS7qhP
FHg/5f7xcEDHi+4HLI5c+4nOj1CkRRzjl6ySDS6S63aArJHxh7bGHjj9fWvVkcXojzHVAsmMhzU2
dUUzaTrE85Jp0mkRHKMIgEv5a/ByM7QmJAgzC6wlBkwmwToetVdrt5T7xsMWb49IFiTnT3HQvYK1
y8vyTd9BQ5ug7orrN5sCxKkYWLHpGvasJpUNMG8xVsYFG+wLfNHpMhkBGMKMNsKlY8SuTPteR19Z
W9P4mVdUMZ48eMoMfgTpXg87Obz8U2Skp8iRI6XXPlLOQsQmy+c2cFMAONsu00tXuvJbkOqH3s79
aNnWFjl90VX3OyEpISpH4dJHFvUFn0t2WoFLFVE4EjWyWqsifRIiAGQ2kwYDd2/ybuFHrCnqLLy7
jANKijKiKfELYVA+fd1VNrIUXhMqSQ6x92MNSOSt+7W0Wy5+KKR1npNxPZRdILhmFIwOXMx3J4EG
zctW3LE1jfcQdbgTlYnT93Abr6zEISXiUMNrFvJVM80CRH/Z8LHTuJaE/IztgMCkvycMSJjDusqb
paAED2qyZNJusBWrJ41CBI4tm5E9SYRP0p3sKUCXKCbI40TfAxRH6mNBfIsm/6vCc4O/ZMWMRe29
8Td1YYkfcuch3TrGS0NdrNLFK57blJzu4boNNskTnOH+sP0U2bYYb8Sx4nTcBdDBMqFM5GuC5m2F
7zFTd+PfkOCy67uIaS1WCsNcmVvSV7khVhQ7zMuIL7Hhti9cTahnu+6qQzopLufHc2XHx5oPLt0f
jJQ+kqMA/KA/y4JYAOPJfX5i3vpEDunkCFRSCFGtAd7/0rZCLV/ECXwg3NblrXUWXWHx5/FbtjtD
ojhUtNs4NYNR5892l+WIWlqc3qjhcM7gAVxsKu5n47m7HpwcNJWKx0ibvJUp3eg6/4sMJnHY+XxR
RJxZtPzLqBkCG8CZNXHE8ZO2T7xh4QCgABCBa4AVugdRg5URQNvuGg+0KPFzqJI/p1P7fb9GteeP
WIVvaXlL/RXXUwn4ExmR9hRsxOr8238D3YlV1obWpTtZ0enCvEu6AQlhnc3XhB91Bi8bKd4wRIdQ
CbH2+az8hncyMTopct078/Zp7sJav+TPum6Mnm/rt+DK0liaIFKfWyh9Ua3ylWBcjLx3o+NmXUF4
QlkquSUtvHnD17kquvku9E1qKtP9pyBn6LO5U2QLjk9BHBYTKvxXRzJ4Y89J2/j6aXTt/vNq9XAA
pw7bk07NiPJNkOhcFxcTdtavIlDs79Uhu3nGgaVIPqpBnBfI0G5p+mXEkQHrlL1B50aNjG3maVM0
nLFjC8U5CczIyF/1llaqOhSb0tdPqS5WxtdNA40OFeeMg3Tpwhx3lQQpONuXa+I4ffFH5PfjJeo+
JXvikB2nLpnnPHonA3R6/9lzidfjtpTZlJR57U1tpUCkYalXig0k6PnukIMHBFkauw7NnIMaSqXK
MyBiO4mcYTVyfO0fDza7gFmwEjySgsMFKNWO0SF3rWFZzWNOJUj/4SSH+yJRV00XwtvqkOSguzuB
5v7UiQjN+oMIdydPUkXQ8JU+kCHG6S1f4GPWmEOp7gAlgmWho+RBNziFktbPHH5qo4TndlNKDvbN
ipeIy4Ul7OL+Hjp/IDcpQ5z0PUzPhXsjlYuxeDPazvml4lERUGDd1HgP/m9H8xXWFCtLnGVjBun2
vjGqHonVj6UbW6/XSnnjlhscK8QKTugyCU2lT+gBz0zQnuWb+r8BQs4axgR832WLJJJXlOlFtiOZ
hl91VSnVCxsnmM7c4xt5UZ9ARgPHlFz4OgALHJfdjjKIfTqMuCXZSF35Tb3OPB6zWwkD2j5+L5QI
7vaTXXHfXdu/FZxmS0uzgpLpcH5sn/QHT9ziUA9guUVT7PrkY7aeh+O2gIN9WeYRZJoKSWTcjYRB
bZbd0n1BSoW9bn0nwjhZugq4v8Fy/GR14NNBkpuHZ123nTSKd7l/5riSTdNrc5yTaHvEQV3Lt83T
k6SEqAbOivyOnuu76JV7klWGAySo1+hwQSYiuewJzeawzXDC4MRXUr+TKINqiEU7B54l3gL0hsGF
nT2+bETpY7uQCwiI7o5uXo1I5cBuUsRl1DlMo9qyB+7nc7b33YRKAvWjrL+FKupDuSd9MHOfuLpR
rIEuj05bC17x/FKOyQv1prrf9GkPRJ8pRP7w/uqxdtZ5xCn3+ObLssS6NKYCNYvjoIvg+DVMh4md
TabUMVrIKvKNfQb/Dklf77PVhlzTW0ZSNGDNVmAfZ+rnnZPej+uV9jHpAfuVOykG0inFhMnECoZW
mfxAnkNn6IIu1NNpm5HYqlGME7xwl4K0if5o0L1ZEbTLHc95eeh8tATP0OzNVA0dsslCnI9KU6Pe
ZvHTOYydXxWY/xh9kMMxScIknNpHXcNiyVA4kO64Mnp+VP7EdkAHQivBEr5bMEIB2VubXQQEzoZH
/h7eMTpnn+GttEPCt3yShMWvPHEpHxGKsyqAP51WsdCQm0lv1q+5sx6ydRzB7SSw39+LR2+zSx0T
oHhRvcNmyYzoOKWiUkPd9AJHRcfGwv7KCBQ99wBu5NxTE4SiF9N8KTvyKCQNnhf/JHZjJap1LmoP
k4ODGKFhpZ3b5JJ/lV5u0xh3wlf1QPbycPhUu9ubuUFWhJkmo81AbZWWnenlFVpFnG/2SW6nyS38
uQFUjTD/1ZjP4vyzhU02OiZE/zD5zmGM3rQBjT14ro8GlK1mQ+8Rp/YhNovcX8m14Jr8h4BLcvic
so3f0LvP5DkTP0kgsLsSGYT8/xUIGdBTryAg9SwnzuVOaEO74roM5ZP/1RqEn1+GCcnxliAUtm1j
JR3gvZwL/k7VLu96VW6oc0QTw2j9gE9eweBV8JIhY2yh99AI3W/Tm21szBCRzDRweO1ldB01k+5X
rqX8FbL8Dp7sh+Hm59rlxd2lNBXjwk/PUcj81Po3WZHXx3OMdElk2rU+uCOe3VoWGa0k1FEqf/Ij
Qf22oiJH44Y/8UjZjTjnoWSdEaqRKBr0ZaOZhFrVzLBTPKkRd77d8eyVZ1wQtE6uG15Gmx5gPx90
2ZrrupN2jNOexCcDkvnhYv8zDxGNQhqqbD7yy29uGsyryAF88a31bdGkTHdfNCX8SONA12lqhIEq
PsLEizvqReyZBzenRPZyTVsQSjeWo8IKXMifmIy9I6htjBabwRMslYG/hGrKXdovGwqJiRH+K/JM
Kv5blDT7CsPdIwwzStyDa2AIPMCmrymsmAeL6KgKXEnJHfguRfLowWmVwGt+d1qG8DR8YWgk2VMB
I7u+UjRVO1NTw90b58PFziJte7tR/SfCnXJRIdnSrOLtKjVpK8x5ksdPehGg5Y6GGj32eOe6jlpt
0cevSQbkMs7B/LPFqL+caCqf5PHIm8meePR8YlShHqVfAOaD+VCldD9O8HOPafdjpBGwwzwBVQ0p
Xf9YC8o6QLZoERVFWDXqAOjFVilzBmIM7UDDpKmHRVtbrax9SWHFP35mYtoQ6G4ZVc3DDB7dx/Et
wYQABoTVCA3VfUf3f3BhAgPTlFjWx0IIEILSE5xAZY89GsfE3FAnhFRnQzLe4UbFR4UW0pdrCkEN
A8LVaSGI8puGhdgL+hcnfOEVqbPZsq/vct05KM0X0vWgPfSOYuRH/chzTmf59VFhJrdTHWEdbymh
seSncDG99EkWrdQg7akOmGqSRj//IGxcSAMbCnnq+jbMv5gZLHAxUqYTlrjJ8pBWfMd0lwFDO/Aq
YYuXyxcZQoFaFwDIQUHmu3Ffk8CucrlFHdXeT90Dmri7EOLALhtu/Hfs6pqHe9c8/Z3xBrMRj72p
XY2lk6SUGEnokDDK3B56B8W13Ach0VmqvDtwxB2D8Rj/hN9HBz8Szt4v8HIWM2RQJm2pdBKm0loW
anzJnsnZiqsm18MI2yynjNGQ2b6qwx6PV7wFHjX1MyJKGyKDztab36zOb56/Esb4jgpL2xbevAI9
sp6j4HD28RYi1w6FjcWFtPA5ffIvVPcIKWr91JmSQNREPGXR0r9GrxrMCvxNb6LWqBVIG8AdTNU2
TvlPDo6e3xoeYwatTfOYXn53y4k9m9OynNiiQMB1v9VHplJPZtmdmgvyLtEZMPBP15GAK5ZVcIW1
y51715o5GRYiGCD1pRwcOLOwvGeFdmOzg5O4GblU+q2NzUVbjnHK0S4XdvWB24mxpUq54SBHR1jh
IMdATP90bl+0buJ1MH/Z9WP2xadgrcP6AJ6Qk9vDao9hX49BfibrnGuj3rNK7j/x6AEcReA9+yIS
IR3dRURkc2w5UyBmHsmowZsFX88721CBXfwv0RxrK9l0PpOfGsfbxwQrF7kiJtUugZY9q7/q/fDm
8jaolN8E1atDaAcTyK+R5Lt8p+Prc+fVnEQFhif6Z0QIEspsexmxbxP79zSU0bBeeRe2CJZCFgX9
uYaisD5HPi9fGpxd2DLw2pJsnFeUCnkczWPltewg15jjYazCDzpxcNFAe8kw67821zky+Y6CZ8/H
7y1RDFIYTJSaIzP2So5P+wmkxnLtNSORi+eRgDl8aTzDZglF+rErqSfGRq5/rpzSqmcaVGf0Ub9E
MQxIfdKhnrh0juPyGLs9TGLmkk8YEV2iIcSvkAegcjYht5hwXkuOK29bqV1VrBnesa7Xy2bYjTyP
WYBPFPwa91CaE+zfzYO0jIdeuCGw4O0RGwO6V8Qj155+JKxVN7N/SoAc2ysbTlWH+I+4NxeZ5u2D
QRpKrqil/ij4NVHCMTkmZRlcnEjyy/MUmNWDkZ5ZhHbZ4FTKAs1Ox2j9t18QrCUvlI4BjoRUuNZ0
haDcQ3rMzgA4C3+YlYLHRY1a7wiBGwoFfDBImJuy9vKIw5sBX0o5kv0RQBQj3o0BXeT9mRFa22Vu
rK4/sLrBJO53rZLRc+LAY5E4/Uxj7XNPIpxcKwbs18lgNYLzWUy2cPa/9ogmtigqqa4djBx5sthu
L13eG95SjoqWVbcN9p7dBR51rmrj4uerNfw9oDh7pD6PhgYyoN8EqQaCbdjR9A5fTT+HgTkGx4Qa
PsxwXaBINPVO9jdNOBB7Auj1kwB2OGQSn0ZLB/nNx2YhKom8GY11Fc0CawHoP85WjPISbskFvuvV
gQhQWdxupWRZ4SiakUZas1MZYcpwe4yv+xX/Zno0BTNqyKDASh1+YEsI0LHVl9supjFD2S5ydX3x
dmwyL0l9FfUIJkInnKlLryrREz7VxJlGWEME983WvRsPZTm793CWVvX2Q1NQ50QUqoxO16PNRImI
avumUn7M3mxel82oP92fpqQnQ11oEZwo6VcbQ1Yh/v2BzNlferBlvxCeO5S6kIhnzlHLyd2zjXJT
oX5rz9NAUSsd6AqfQDNECjeu2wFz4HF5S2mQPglSW8BSHJ+vYrLO840n7Am8c8RTKtwH4GS7Lx0+
M+oxQ58TcPYik7BgK/p6FklS/odH6sN+UHN8Zqi3mdZXEZb6DoAgNrxGc2XmOYgciHOOCfV45Nb4
WvLwuBueGhTfLMMPMGiMYX4qfK6iEfKCN4PtA1YwNdfZ9wbLiVSia/PLrvaXBQgbTw9N8mfL8caU
+HIMAYOPLfvnu0YZtz8WmvHpPpigd8YeQC9cn2WGPbP89SdWmRnww5QeUwqni7SzZ8fh3RRHdjKE
x6yTAT7NJPPupVQYpS1CCtozoyDa7AlK90kesraimkwyb8i/1r1p5IXUG+wop7y+lBwLdyVgGiwM
TRfKvL8vtWO9T1TcgVRqBQXgylEJhIUaIGGyPpeHF9EUt7mGRJ/QeeGSoAK/9nkhilwVH1C1T4Ps
WM/41F7F4pmb9AyhFvOHHOkfGowCT2gHszo4GKNiAF75SQ0iQMSJ1oBF2aw2pVOtOwKm2HxuJXbY
0dMdoUUjm0QFivNROhTUz2t8F1sbzmkY4mHjEnuDOBoJmFeRIylJYhPu3+bkw+s3CpQVLNXAdwZV
gvSjEU7sP16SxECiwb074Lv1BfB5eGB/0t6jM9GD2I+WzNLVZ0i2fAhtK2w0+JOp5sT6rWWJI+lS
NyMLJL6d4ss1S51Radkci4KCx6OQss1NOZRO3aZPHRuQo0NJH3QhNbDi8LYioPf2lbgO7zRc/TJq
dVOlr5RNh6ZTHdWqnaLhcEVLDH+Rg1yuRn+gHoolj+0RLM1Kfk3HXIaIF4xMtxFCQoBXjL/MoH80
wRPH3sJon+fBhVYwmnHZ/ioQwUFwIbldUk4BIDYNd9UzgiWN8MaSPlgxd/K3yWlG0M09KqqkXcFo
g8yB3XIrLGa4u0+5RrBr1EKLhV+mZ6SkFpNJMwpgw91IrVaQSx6XMvuE6jSPHl5E+CKRed521h6i
RndWK/JpkMLkvwhfwFTsC0h6yy7Ws9tt40XnBj4Z+ZKdeSbKMbao+agbDEQB/HFI3pKxQJPwg70H
QoYlcdVRoxpviZZfAsm0ZlgRvV4ynVgx+jRZCbOodxsLHoMQoJf2DJdSRu6or7tJG2p1i/qsMPlD
LAG0Qd7t5v4ousLQ0GtO7Y0MH9jXOjwjK31tVR6G+iaxWxVDiJKwP2gFdEV7pwC1kykcWdgpijkm
MMzoxgs9G/ODGm9OmfBXHroUayy8uEDW2XA88PbOUoQSEBK9Qcj8IveSvUKoIw3q0KfufzkyNeio
rOlnJBym652ti4kRl33c+oTzacLYSBqBOrUAA1ZvO8A/7jJ6MoI3MzG5unr9nPLga5JGpbuIuh5A
I4Sw/RguqQzqDKHQzOTaghaCX7bquyD6GgdwTGGMXf3pKVFBCAaPflNixaOuIFINU7EEnIZ9Mb4Z
3dk4hLdZc6bbbQlA1/cpoA5cmG3KIf6Nk/i/XkdsjKiOTXxLsS7dxbhGjRtf5FTqUpNYcAi0kQZt
5l2XcuX2QcgIMk9deNq/UAbX2oAZSyas7CKDQAY5R+rYaBBKzEAQhzv1tkQHcyAPfDbViFXgHQwX
hZJWd68YcNZ6yFMCgG8Mdm+EVoupOnGeb5PsoRTp98LXPNUSJc1gyurcNX4b3mMwwR4gA1IZ3HlM
iwOQLL2PRGwrpQ9PgQZ2Pnap19jvZBSzW/8yW1C+cef3HYS8+nVq4OnS2J6q4GxhOhdTH2pMsapK
p+L1PnZsdpKIOsDF5MPcdL4njg8mKf2+32T7oY1go14fLml32e3RE8hNYpqi8I0eZ7dD/IoHIyJY
OMbyean75HvttQSIdSZSCR7OrsfW+8nwHSNrvKrUsc9UlOik6LqgeYBHjEB9VGFvETTg2osyBsZs
3rLS96zGBaCZeHXPORCzXh3QS/DGSZKBhS9+qCqBl0c18tf2fwcPyDV1+pAyGfXKCCC+H4DSa0P4
SGQE1zdZ2MGlYpWJslDm8QOyUaU6eu/8gVSi/KOc7OEyn5QIlkyK5DkZPCMicn0zeDQV7mt0zQsm
oZFU4Dr+6x88XdfwjT+Uk4cu+B53Efu6AOboRwyhDlF24Jb1Cmb+8H9ViOsWlfTK0Qc+TDYZfYvE
sTsheEGNi+RSM9YAcUZbQz8bTp886/dOTo3li0Hd8YCbuOr9pHePwgOOAb6fmbOb9+TcFDY+sQ3x
DE9LDTLxZVjh/2q1BfXbwPHa7I6CvJ9PM4yo9ijqgqoaXj/AM1ykm3zeiaBsRTPkpT9DXK8nvuPl
8uK3VXBHrI3J97QZs1AIg115PsDk73nM3PzlxrmH1dIwobBYdF9d5gDoAL3wYHrlXPpeY1XDw7rP
zXjuUBRqOt8bTUqE3FZuiuOYLyzeWDmP7nWWE22piq9203+bxu5+My2UKa7G/CZQuJjP7IB3LIDC
AOMsNND/yIxuh9tebrC0QgL4gzg8CDnDksTU55oKkP7FZetb5ygtnSgM/XX7Dbuj6ScrF617Ssp6
VcdC/A43r+32gjA8KoLPwvUrH/X5ze6XptIuNZFfzIA0sk5ddZkqGi8aqiLaDrqq3/wEEJOw2Y+7
cIiEgxw2TycBR8T/krYDr6+TWIVlqmqpypEZd72nPYzFy4cdrZfCXApNerk2PJYN3sSqLqHzpiaA
t0ywrLcoGIRjnUm6a6Nzr6tKeQ5gFENewW6pfUxIT4WwD8sxPEh7POvXDRdmKEuSCTpafqU5ApdC
7WnZWJdEBPAlOiZBud/bu+8FafbSe98sRkOwWSzwKzbGHxHxcTuSX3i8d9G8SSYgtcl6gu3tfhMV
49jdWzrPnkB+dMKUJ3OjW2zeVTlCevKZyivE2O0oW3lvhM4MVJHH1vMfswbOHQv8QRcZA/Kkb5Pl
/Cpfw3s9YvMFxTRudXxcO204ih8gnLTZXmitP8qOiVig74302QyDbZ7GJjBH5WZ4/VwY71HWz+0v
UaiquzSsBMj1s6rvg1yEvVhmPveO8QguEHPqt5aBT/CUBQ7D2eErZP2DPVRXCt6NzyI9KEFLV6is
l52Ge6us9xyqB8lqqm56Hb4aoNHFgpGPKa/19RiPI4mSWGyMQxqYLno10Aeb451KjyHcOYGXbEWC
PnxvfMHIGY+nZ3a7Kfao03k55XHTUQ7fsv9LhDJpFDfeLzWfGGCN2RqA9Ax+Xw1qQ5SaFfBH+lP8
G9zyjQXTL8rYipjp1ngqvxvlFiJt5E6WbPnqknaTJzCsOm0RiSnHvDafMa8QWHbtk8uED4qmcNmZ
9ug3XQQQrTG58eEFQjem8tPp+j7k35j1BPPXvX7z0SpiCSrg0AZU0wxmNhf1OxTNKWtYsJVcW5VQ
WvLxiPDXx5NwKNFGvkm7qDLHvNtLQowhQAEkHGy18kkyk4VUiNocKxriZ/fHMUKGgGs7kWPTPTEz
IE5lkMvsXxyWbg6zChiwBXywNllb7RM821v/mx3LJieXaEPJrsRMf55+n7LKhSe5SaEToTp4o7EH
6DWPowlhzYUudeVseqKr9ii1Mre8YwHGcRCZtSKb63sLoTg4dYuNeU8LU7sgkP9HTfn/0PAdhpuN
jKKy7gyBXXamU5pkerUre2j/IYi/D2jBDfzjseyqS4nbdJ9KdjkDvsf6g9XyAhJxtkIb32iMSO2r
kfgU0kFHXRxk29wu7nI6Xf+1k5ZiLmAgiVGoVq+C7BqU6HP07e8+e7zFQVFBuaz1Q0Av99Zpubke
6fGrLjDB68fYvgii8cq45GMMhuZJfiEBtqFi9Di0NPbQjKCTFm4K0gHeunkYPa9mVG2vGyxz1LTA
zJu73/LQqduaVQoXp/0waBldzBbVtC6DvLFw5Fk8BGaw6hliEpR5NLxV8FkP8MM0Qud4AR1aALZQ
ujLG4qMk2KgH++iMX0DoPN0fIBzGKFQRxHmslWgl7lzsygIRH7EmLmhn4kGErJnrX/2lNsjswx6c
3ZhWLDZi3Kq5knjGKL3H9opFcjspYIFAIunltSaXVsN2ioCJnHlEXFzDjXZULuabvp1GB40ZxvUt
Hia6ff7JM+qdP5Cqaa/cqW2ODs0uDO9Kba50csGQ9D9F+b8NbXlFx31CJ45NcvmjP9Km1CdLcxSf
GyHtvNiAgSxu8SvM9A7aSvu26sEC4zMWZdoRhfXGCk66EkUmLJser+rctoVdWg2hZuAJKvxl2gZj
v8p7M1CztisiqwxdaUBkuja4vfcJT1ggrzIanI3LQ1DBhJgA9uBsRObMkpDn47G4thp53d0ixvW+
wAlFeOJPn0iX9SCRXTQR2fkYujfohCgeDf8bNFKQN4e9zfsBOvkSLxrxmlbQ3tLfHqz3Kg7WzQ3Q
53anbfimECrYk2qjVU6HdYB0LJ4OiuEmQyCgMgVdoIreBYst7ALOKwuQY010vPkRWwXeMIL6edSl
a40DMJ7yV5qc81sSRENDsGPRecMvqrrakwdA3IXLsIDHmLNiwe2d5AO9fjh9gkcX1J7L+3slqOGw
aH9Oxolh0AgGbcQDEaLxheHVRUQXZkLzBhYNq6NsGWhQ16Yh12s+7KMD12CKTPCrr12pgkPvfn2d
ahNxwwOUgO8onx6GF8IvPiIQSFGvR5BawvjAsJyaAsPYqNQOjNTbt+B9/GBPKMuet4Pu55kcDPhj
Lql85O2voQ3Y5O5S/DkFppDMZ/S0pKKwqruexHYba62exT01akQDDEJ2NMkHY247cwApNOMNupCH
mqNeawQNCHI4GXh1KqGVqCcHeJgqWO0ctZ+NCSB1DwPHPq9g48TuHnxtASjYSEGF7e8rSSF1tpRL
uqPP+03r62bj9vEbCMzRUZlbc2fw9jSr8A6tlg64lXqo9MrPjfKUCOtJNo0+H60prbDUJnr9I2Aw
D71XHbs4vtDqpKaNaEG58wklw25l1ago3RAjhHQm6DwSvJZAYrl0ymCm4MFXmV5kKoZIDSVt+CV4
KdXluph+L8KHnqJa/IWtadn8+f2B+A1ifsodDkUm56XhIFRdMDWpZAi4wp7GuW9IqCJQYN8IgLrW
XgN3kCbNM3jXzKj+e9wPZ58UbqU7EOxT0C4YoRTm1DnZ6m7CzBaBrpIct1GYVzflg2Cd/cGKJcNm
qVaaPknePvBH6Pm1/wCwxOlv+IDFX/5OtgjOq8yW/gC9oiLwew+eDlcYTk75wDQlq0Bdvs5jaylF
0c7eclnCyhARyp4ca3r4NtqfR1anCqRtfH7LnKU+q9YHrZMZjC8wJuejXmPl/xhGvCNV15N7M0Lm
SDfozpoRaY+NZbVW8kxwdOx7/IFWqinQnaL2vji+9t/FfMN3/fKLLxairr+9L4+25FB8iQWhQA7R
bjXLhePKBTDhZ6NM7s9+tZuAjzSFNUw4xCxngawW8mHeNoj3+/dbt6/fFlSxVuOgjKCu3W/cYmtL
nguVMOtXqjK2CTBlRidZzpI788Iw6hV695FCp/u0PKSymefjr++6yxLhefIr3YqCDU478R7U2ag5
mpqMf0TnGnWRrIViSijoPnjBxwWq1bLzGldZWXT/vLp9ym/V3/hMVmL92I2WC+i8S/yOcSBgn2dP
buWRBEjizy7drxjjlOEM3pkwKkIsi8TU0UmBrXteGeIDcuHvdL9oAPz0aNRXuG4W72eduipRmAb2
b/offjqYqH+VhOOxoQ5x+gOnhHDjb/A9KkuvvWKakdstVaW+nZFgYx7BepjXhhe/90mNtiPqqn3x
iwv8yRWQI+lwfta0CJe963POP9608yBgCKA/jyOSALMoRux6IHnF17jd7P9BfvfCdyTVMATFcEBW
sbFyaJUuCTwBwcyrK7TxJxnQxVviVBQELCGTqXZyjC76vTHATszi85898n3z0tt0eL8WnkbGhVtv
FC3OW/95rNgMBEgVVTAyBSQYMPXZL3DwyIohkV5t/uvwKai3x/dtFDVJEhk9jWpgOU8bvuxEtxwk
UsblMplKULApBXzF6Z1xvRgkoT3KqthV9rt9uv5NRR8Ds7WobmNG0+ZE/dmYBdFWXRXEWH9rwU8H
OfsP4PxRiOK/rlcla5aN9Yll+SQcn7Et9hAFU19QYxy2OV9OVrMMaHvOJ4zYuKQwLH6m5UGY5lSJ
FhYR6PaKzgw88wCvUkYF2zBPdGAZx3WQdsY7Vz71JvFQBo4Jxla5A6xnUbfDZ02y0qspySThJbDo
dJtV5XHWEYj9blRplbgjCkRnMHaI9tMMuz1Qu1EERLKKPChOKX9bAPi22lcxZsBMSvoz5spWc7/x
HfDjz/KXUsM7MnwIjkz4JsKIlBnn7m/sf1Dz1DEcLAXceu5O7OJeNp4WfqI+PfpHnFfQU4VSCdLw
G8KjLf01QxYTClJs4YldQmkHHwtDpHZ7Gl5r5Wo1NkpsKgG2rByd1qRtcFFcc3xKyCvcFfnQjdGx
mTNaqlSpm+K4HgZ+ngkoLqjqbhy+kk5by8gFMaw8XNRpCbSDWSgqQRxswB8YlheCBbDJ1xhOyEWI
hsikNVjE7SYBC7onvVNUAklkS+877J7p/zX2cYRg+hshSR8jL3q8WQwy62kMyvyEB46nmRBharm8
+HKxFlsEwS2mHh0dokNIwWCpqFoA9aXUKMIoXnKwmqZ6z534Re2onq7BqoEcAKBKCWdsP32ygVb5
xgtM2Vem9l2VN4RF90m0k5i/Z0eubu6EtTQ2/WkDXA84StfyO8vHuVD+R7a4Hs2RftcEs1krnJYI
d+X2pMdKO45w/BZHnxVvtpRNoTpDUfhqV6AqHNmu1Yw2yQDtDNDRWtLkOiFTsSn0QwFEjdi4h3XT
ZQBMUhBgqb2sNj9Nx9uXp2NVgGBpLvRpUz8qlyVE7P7gkwyCyX6WVHXiMTUDpHbX3VmsTjJodKTR
MnJFS6zM9L4nGmXOk8ZgsRyEKVsMa7+m6dS5wGmy2MGHbEcPH2fKdqEyRq63NqPn2jKBc/jl6RhI
Mwp9TB69N2QdnsVuIGRtdxNHt5mwaURkOavoaP8Zz8fTWIMYUZCZbwokEnTZj3CiW9lddaJLtlyC
mYWKgL9A5FX33wl5pPPAk3/B7PKe2llWrk9xeQP8LYo+gsjCvFS3xAOBe7MSrluuQ/GMLGuoDrMe
maufKZvhHdBlHxVhIwo1TePxyGWyN9GORR21W2QWJkpci20EdoTdfbchVL3ju+HYW4b+deFwSzr7
LtrngMNL6TNWVaWSMnqOMDkgytrNFjLc10k7pgB+unp4jKUzMNEw0lKXZ7qrSNSJByVPjitN49og
D4/5j9gb2CL/RWKoGl4waL3nWOU/g4+TmpL6FBipkd8fZXc5rxr+K7RHmM/nAGdrowunJdEVB8fI
2rcI6NG9eUcdzBiLTV7/V3jDpWgHRU9CPjVAkFDTmnTVDVX2D6kl6FPRo/WImgOLRoikbsgcmVXL
St6XRC4juG5s+W7yweuxuFJ+kmrE30y7XPeS8wrv/1Ry4+HrV6bqlFs4CyDT64L9xy0/PEZWB+Yu
yt2FxUWV0Pe1nw3+1NKyncZwBrWHXymnY8zgpMzqpmxW30UXstqS1vkIW3vwqRGDIJIxxPYErUUw
eHnd4DY6IHeZCcRLbItqnzMduVIajE3PAS49/0FRwh7ZNAIECj80xodNJ9QDX8som5OFfkGIATpX
+UduW7LJYk9FE7jpF8nEvoUVnlcgcgGQ0DyMIOOigKQlBzfhUr+HCsUVnvJqqczi5mAKx2NCJDEz
gwpV3827yEwerFZLQyD3ls3odPEWOHQDnqz38OxxFAjP1/ayX5LTRWkK+H2E/ePyImk/8bRF8Bh9
UwS3ZeIASrefnOLHl5qeGfs9hmJazsVHVkWqiP0WIbfIvVeR/0DH0dyycB5pbAOLrUv4LRsqXmOs
E8szy45wnNH2g/uaVts+mMbr4vsNvVvYD1p5TRR1G4i8QkPNnpjuvF9JrwFUAtBiVrj0TEjLQstV
QJ91g4jFZ0NOiJZyAoPm5s3NjGHu4Vg6+ci42RwYHq/XDQ31q2bIKsJPF3uhpnwoLi0wRMy6WRem
3YrLjkHajncxl61cFEe3vE3MW0fWt5pPNBSXZKLidL/vkDHaum9f9x9hWbo87dxrbuqnUfqN2/+/
mCycLm8a/33mXsQPopNSU6lf5fNNNhSYQKd07oE5e6CdfsgaBlMpqpn81P9aTOeamkaXNfHEOQWM
FW5w2qJjWJ9gMhhX+2xt5k2qrHD4Wr3vpJs0AGCxKIPqgkYB2K2w3dWdDTBYIUvZKOXrZnj6cTH7
dEig9MCBSF/aVmD1jNV3hUVuV3SeEfmRIg5RWr61DIcOdOlT2bunB/Qd5yyELr7/Ro+4yIKWiW+i
ADbcMr0BqzhW9CAykAJLPKN7sFD0KqnyYu52WAhQblRVepPEwo7lIqbbah4ikBQMCk25yaD3pidB
cEup3C9xieKoxkAoq+xaDg4sBoq5X/lAg53WPi4mxD3qaPAKrno3pTBeH9y9QqEJJWMU02g3QSkt
jRa6j2aHxd9dKq3YkRtfLho+h1w6nl2skIWut5SzIA5ea7PmJLHYqvUEfZMhErjHttXYy9V+jcsM
WnFNXfrphQLZ5hB/ffVI8LB9TTWJTblM64A8LdHHGypDBSHDypKLUDNKO3rDlgDVG1+xYklWOL7I
ye8XYk1ngJB95f4Xev7B+Phh8sUpzH3g7THr2cWG2vpjZquCqOCtcMJMKOVCPfOvaW3V6qQxePNh
EgtECEiOKEmoDBOMJfsp2cL5OwI63G+pbWLkV082NrxGVjJJDmhC3uGlLDOtpCbYVcu5LtZZZAy4
8u/Tw27D4TSZETj5752XJe3KnhAw/3a4esFvnk38WJFIqENZ8LhJKSIjwm/HB5+WaHzL21nYoBeo
6e5IcM11Ny2XEWG3kVJADy3nfg5bqltHUrbE3ssnApEIhCy/s1YHn74sYsiVr0nJP74eO0b7CeR4
9e3rs4j+P8yIjQq5+yU/Wv6+ZakLeGAb6Xh9sAq+Smim/nZOIo7KMcV9zhU4KsVgBmtMgj42gjUc
tqEHg2HbEO0UX02yrRdXrO43K0O4v2oDPjkI72VuSj0Yz5yQF9N8kqP/cjJN7T4wLQwTkjp9ViOV
TA62eKZIavsaQ/DmddCLcJ8rx/BzxN21QT5TIO4jKhagGW1r8Q4Dd2nLDl9g63dgvl6WEn0H87ib
8x17vMg0VEIYN+MsAW9a7/45kEyQbGuyyb40he8YucDIKRUOOHRzLaUNnqUVbjQKal2pO/yrfLNd
PFquH3iEgIdhusGm3cuk1jpmHoefti8olBuSDoO4Ffbn1jOf6/CnJri/MWxR7yuosUUd69EB6+RW
rtKpirUPkpc6ryiQJasSdw3DjcpfNfYL/jkbwuHnoqBBA4ioowU2eJnhgytj2uOqCaByGCUB2DUn
jKrGii8de6rrkVHiJqxggfU+T6QMcJ8Qszt+onz8tPKnl1c3bPLAAkTq2gKdnSljGsX6bZOpxWgs
FJkXt/+feassFaI62wdjMckfqpqkPO8Nzu111TRSidCuJXAhMZFTJfKkYTZos9FR46WedrXBu8CL
5ntHpPWk5qZL1kzQPZujPoHChgNs4RUSCqd1AJS3hVB8utcmf7cwCUFE7tZXDmoSPwB1aqWJ4rjH
icCtv3w8KcfXvdyc5m68pD1skkT/BAeuSCji1gTySgzVjN0HYWtjXXOrP+Z/XHEClTkf7BIe9qvN
44Ffhg+k1YSGD7Dwi+J34QK59kl4bDywtFu7nh8PpdBIFCEmHjmxmR+ZzQ/8eOKPIZhLxsIfE7vz
fK/L6FlFHL2xPYSkvBhOYYU9XYdSOs0MMBus6rQcKbz9qlXUEJK6zgUUu9RJ/wx0e3gAJg9u9VfE
w0ygVlzADNA/28ACA4Vb4UA+A1T9c5inJC8n941xxW+FDVQJui2KdRrgcxP/ulzpxAcOmoguGF11
RDNEKagaQ0v+QOIOc9SrIvbmJ4QVHZ3IhZi/3efeYyzbf9tTmoayUXibf621w2MrRZumipxWa4RQ
9InhyVTOPJ/sjLe/FlByPWtp+Y7Imbdxt/3cHk59cPPYKPCaZKIS/YiYtPW5gwGIP0XJJJYDCpPC
jCp9Ogl4HVSY+fV0aJwVaZbYekTQmJpSNVtHNh0TW6m4hFZNClmBGBk5rI9/Du/Xq/4eeMA/89z/
VM8LjrluxQBT+CR6lI7/msiUccUbF/fztUidW7juPAihil3OIzZCxQQveBg/sRpGly/eh1cOQal4
yBA1NeUXd9pLwwJwMXdZstXXT6/lWgVVQMgQFXFJiAI6kK/6pSmfLHyfQbX289IHUi6T7sy4/2dR
PcOOHqEqgA3+dVzbRFbYMXQwn+8cGiq5I2rKubw1F70LTktJL4//b4NjnBqGHvBkxZCSLF7vKVPO
AyatWOe43p4tyEj3EKiLI5Ieb9iQkpTbZIXoEWW3iG3hdACQEqxYW+JQTGlr/gu0okFO5xOFo7tX
TnQhNAnDT++f8R03PxpqSsjAlQM9XmCflD1hUUvM60rpuSxLWKqidlyOjwYAmsNw3a80ky5GTuiG
bUXu1hddn4MdoEnH/Yvp12W1OsabPwfmhlmlWtgKOnrqwXXo9tprF8c38y9MEL/wX0UHefHF9MuG
QDBbThIYd+SmPDz5SR6M9DuXveDuLaqUipbB6XQ45L7o6lqFoQPAl35SBmypDV6YY2d6otT8Hg1s
BcU/3j41UiPABc2n8u3VRIOlVuQ/ejgmUOaR8ZRYw/9Dvz6bR+KBvDwvAdC5GGFaH3ui8XJq8rbc
hIBoFMN0auQri9SFMF037wgPe6FbcDU/+Rjtohd43v5dMO0FmU1DIC1W61TklAeDUnR6pesq49uS
+kD0YPTk1PBPZQ+Yb638Qid66yangv5bZgYq4+xYxV1t1riNF2zTa5ewR9GJYPI9o60EsnIzvBZz
nuj9wPtvolWnMGss+g7+9HXk0ZAkkB+bw7ZAVOfQ/yPpDiGBBu0DfwLy/rpotDwujsvDYXENLMTj
RRoFE5i03AtjNrztK6+H6MmDEFym6Kfrn7dndsROVeOqiEpaBzuaviO3vO+/ZhYzqJmwgTA/K5hY
2rya+r6owkeVtJ+KI/3/CKA2PA+Iki+r4eSfYRx8EOXuAak/N+Xv+kGAo1EO3XacA0rTWOccV9Kj
Qbyfh4KhgKJR2iPD9WcmO7CQvMGM6drR9BXb0dTw+I1Z+nwLo7QtIFMRRyexSrBq035+/OIL2Tmv
nHs4L8vBvdXEaJisHG37xGNKJy0FpzaiFPh/vsqYX3YuD1vF/VidvO5Kdh3kiY4SP+fIzc1EWaeY
CF/DODGVcl2IEIUvLsg4umjprzGj3F+ThO8jYaaL1W4/3RiUxWNHMgzLOTN6if+o+gOgIVvPvmao
v0uhUMu0MM0/O5Tsxfo2EXMKVZIly39S2M3qQQLHoF48ked/3rBvvTpesMVvguT9TfjVk2XCrmWS
KsNYvpjucO2kwVXgdv/+7JUyKClL5Dia6hLA87e71uthhSwY75W9+8OCY7MugrQoKRej6jAGyvdK
ErCxQZ/bMAJilirwbSJGY5X+FwHJczBlcvZxMlBViS7gyMYtvhhiGOEfIJiuheIqtDpo+/AV1AvO
xa2LAIPcwxHWsuhzqTMkgVh6T5kz/8DIChcYepGXPCn4fvJf5VA+bRHbDATt6ABtgqMAfd2DgQVv
wiN/ldxOdY39FghsQy8mPo/LgOCGOL4cNrAQ+smmJ7rTq8AkSSg9LATlZhGVc5p8bacuQP0NGxrV
Yp6R6fIIphrjaPwAMmotvxeY5f1VJH1bz/JYIefbmdnRfwA4/qpKlO1qz45uX6UVVimwiwP14e8K
iBZTn9Aeu/HuTZJ7ag/P7i3MWlWiDqBqwH0yyyIJkoJ21CHPaKw8mcb9in5mrwsShviWLZXj7hGI
fBA6RCEP3+5JPZd9sLHilU38qXxe+e6KuoFv7n4vR2VteIcmRXGx1sZh8EnPQANwitzgoFycZC71
FS6ZdAfxYQDSBR6ewHUwA3jRQVRqVEkym3rS9T7pTbhgqlkqI693TF/JA7zSqcO8V9uxHVBAL1d8
b7KyXD9Yv4ztHjBc3it/acVmQo27YLcbVdixxmsJ+ziujYhCWPJoFwtV+Ct+8KaAAiHSALrnzh9I
+rU4SIGpMEgynll93xs87ek0VbDFrTT/wVcv9Vd/lL4Wl2owPmasQMFHWAPtrpYUIfktm+umv/i8
1lP6ga+0+Wp8ZJQk8fOaGXAQv+oHj7jKghzU8orWAVvLJW2HUhPflwgRGK9BCteLa/fFT3bsifk8
2vZQm5vLFCvrXkFx8q2/CV8F1Q0S1Ws6iCLorTm8/lyMtaDFLPViW3cfM2YSUse8QBfbNcbi3ank
3lhcgblQJWB7G412ipSvampSN5Dw+iHNtIDxWmYAVmZaN319rsbfiMAhH/VdwRpYx5nPZEoObtwS
uEiGDJpO9stO9ff6HJUBA19NlFSkGXT0bNNNqcCEnedKsYUVfAZgHwLEqA9PdGTaOslNqlzZ08IE
MeKcyde6simmzBXujCt9gCz17o4tHKPOUBB4v3W3bB9g+ejVHoA9euG7yBoH25SA7bXp6uWUU/g4
UKTWysJjjCfvcSWwnWrZoj2gOf5t6Q8nawr+QBxBYOZhxhUpXZ5hcHq3+NtsB4hfPJd4tfnP1Ro+
IRFbkptaQbv5cA3BfHBXnI3+EbQbyiI8wBe+9GkvTdnGSUBnI3qdgxiAnWETLi8ouYkv3BxpF+YF
mCTQGO73iSX/VGVwAXeSV9xoiE+JOhKv4Ke+YGyy/MoNFSD3ZhQwCvN56UIQUtxtpAtN84YLNbF7
ZpUk1XMCylWHE26VcSu905J6wMJ0kh5MTheO5GVYrobXDZUwY9nTtIZjgTnoygTXYZHV7wyXnyVD
HOu5TC3wY8jLGQYRgrklQqC569Yg16/GanX/9QVSA+5LpYhbUfDNbp4ZuGA2TcQyFyKzGrRpzc3I
piLoxkYUqCQvIxQgTeiGc8gOnw93TkiPmhYJaNpll+B6AXs4VxpsoXOl6Kb5Gf7UFW/jfRXNa8Yf
d5b9Qy1b5XJoqRIK3wk0f6HZ0Uc1Krdm8MuLYpNpjaQlzscXdECe8YLC39iy0rrqnn/GOrFQGXi6
5qHhBGv3YVQsH1aGQnP9oCW/GcI8xgT0Yv/e7IPhvVYdunKnUYABvZKclRq2xlH6fNQcuAysQviT
A4y5QBd7X3n6LjBVJL1NaPhTR9XdgiD8n/1rxKn2I4s57bFw18u1VjIHotLh4AVTfMZJSwyHrzCF
BMUPiio+XdEkd2O+lx4OTr4OPnVRIFtrOtIMvy6BsWm/M61X+bHVbGNJ2klWU8SFLUc3BFC8+2Sn
FJVpsDsUenWKcw4lkIEkjEkTqKwnezd5wdd/lLJiV8Ppfo38ipTfigr3dxlNVFifNEUrNfHW21fB
NsgLart2U1lv1mb7t8eIUK2w5VbQ9iV2ld84C6aVh+2Fn+4ISXczjYUZwotJgVh9w03dH9PWBos3
FR3emn8N4nd1hQUesEmCSdmhvNvLHDIDczrRyJeku2vqqODyWRv7q+p2gYufF7HpRA4W9+KzATaC
FH1ExTjg124dIErOiTBUUU3ti8lxa4ScYqSPaXnHnA4AyUD0GjKVLbOZMSVRO/ufQIZwMVipNz/d
b+jAf3XbbXDJq+gcK9hOoBHM2nRDk1aGoBWfCr9jnWTEt77Ojhhzhwofan/PUz/PSxaxJSzBQTl5
5TvsYxGbZQlGIzzCkChLVUR5kqqfsBvEdvsYUmBPz/rOjPTZXEcdVkutz5Alb4wWm6VY8wIUid+7
7flcgMNeG9xdbk0MI1BQjP+1KX5FYtICIM6n6PIQScF5lL4+nsb2auJM4Pw3xgwZNgzr7beXK6la
NEmjU9Vip1Bt9gt/9x08Yzl9KngdpnNYPCckr1qjyuyaEWihS5CEAKS3Ty/5t8iiAMJtE9Jkj8/w
wntxn0k6kLbm7RB3zUmTKoAxdaZv27Gxl/uNwCU7Uhn1JNzS7XLBGHgtskf6iA4jjMYAXaLnqlF6
QELqI8RjPan1Pvk/nztoW+UirFeS5POHGpjFFl4dB0A1otacRlhfgfpOxLPL73FUYR7MQ7Dy7pEu
THHQ3wTFaUIC4sA2ptE2priyOBHbkQz+fTPxzZ3xKBvVNAD1ur1uWCDOwfBkZ7pe6KjPNQGXTocV
e5oMJzPWBoTvdoDgmTFAjs0cNVFejGi7jHELqGMs43kQDwRxOBcXJ/qNpecLgmcWTX7q8o49fylM
nzT9xfBYem6w/qwlXIlQnIYVE723XldyHwGtKNnpk8h7OKYHSkjhHASBkYbffP+MlBRQvxedICgi
wInslEZvA/5adCjqpzfNCdM+YYik+7ZpOnZexLvaedht5Jjfs+rX7lPbzC3E0JpTlDv9VeEpCGtZ
nLqgEdiQhxnHux3QFsoCG0HaRXvf5BV8IDsxBcEh5nFkUaKEm79bOLLB/8tpYqgxg0dd62K5shsh
bA9Ucyldze+sSz0Wm7/yyH8H/YgIAtppQN1PJP7490xGz1lfYA+prl5IeJ4lcvMNt9N1mmwwv9mh
AvyZukIle9bItaYeHdUg+fQlSpeBRzT35wWrMrn/NUsWZcTyfhQsjfnynDWBQw0kw8GtlEV9OUm6
dFN/exbInkSuL5buO4Ov7mW/wVcHs5g1qhE+Y7xHoYB6hNBDMr+TKhPdUfQfb0gH3OYCkLwIP/Vw
o28eJ+fxhTZ5f9aO8PCHQRm5AJaWD/wOsX3BTTWvulERJLzK9pLdhw1l49JVaCZH1BcNLltDjXGN
taDfFjkbm402d04OPr3frUpYge3EmOjCMKMSEbBCvGQsarDmILPP/5oiZmE8Asey6ohpFAOaw9Br
Atdd/tZqcdJxZX6Ny1dp0Dh27gbJRRZIVa9Gsy5XfpjIZtgd9lzWfnhr4+GUuDwzEcIWKTFVuPAZ
Bcxu6Cu8SJaI1Sw/Zzn2MX0FwTXBN3FxjcWpxLPnJq4Yj9+DsDQkfkfmaz2wyBdL6ZmSJ2I2Dv28
+L/KHDmrukZlwdQV+X2Z1bF2GsgT69dOQ2r7BdwaFY6TEByMQy8qHYgHsIO8ItoU2vZ3CXfH6OYp
TjVI1xR84u24RM1mWyIdoquAq5YVw4Qifr6/DiCIx66FodXSss3bBWCBGZuJoFyuQgg0WYA3oKWG
yvljBU+2XnOIXM4YZfpqQewJeHzezEMdFD26kXEjbt07tZe/DzAie4qPiPEkBtAoY2R60O3p43gS
k/dTIhZW1gtz0vNQtmDckosklgxHaP5oYEIYp3DKB5rWJbO5sRNH1cSOfPlY0DHybtOp8RDqDhnr
mp/ijY/+dTyPVKMUAagYh82WCaFURonzdB0ATa2pWdVPfremo5mCfciAzdIM5Lfo2EezNvW70GMy
2ez+snhqd5NVUV7DqCBSLOkD6hbAWx8e6XErM9dp/YL5BGFvJiq2HM3AievMUI9EgmYqoa20/2RN
eVdZLJzhKyv6u/n78A5zUTdqN+aGgHKsl+jVgXhWMmTBQkmZ2yAogSE49sq3ANX6wX6AzB7Fm79+
yAlrPuQf+eXh7pR4CWEy+QcAxSwvYpcTPvnqythxWMx1WZdxzZdkc61b5PnP9uu+w24hwWkXs0lE
DAmwzXWxSjY4sX+uqL5dME6Anw0JhfbFZ1q4o1sUKNu2Hjbo+rZ3WxukYAV5p9VTfZDJBta2+nUS
ERvy5J0tz5vrsAvfXJlllkFfupk6Tqd3bx+8RUUN+9Di7jj8ZcNZaNODXFS5f3dB7tm8YsEBidqu
/cIEl4AQFQfHz81RQIjFvnSogX80+5ZOMsF43r9Lds2RaxtAL+BU5j9nPznd84olVMm38e2ndoNg
MVJ6weFj3q571shf2J3CVLCX4ehfRIENFWtDWXR1CrbUR4bwrmnOC5pGcEdQYSg5Vke6YPsVFsFZ
lOjJVurVotkKupzI7ZKkta6RrhZEWj1TRFWDbsHTFn8uY574niVT7FMm24iQoekZYN58s7BfguRF
/Lbez3z/y1zSx1Rv/TPSE4Mruce/xGSGq26BjIK0AkHYqZ5CrlWnyz0e2ZF/qzV+aZ/WrwVRkelV
bFOCr0YACmQHQwYLGsc+nee7IBTWHDRjcaBtN2BTFVnrCgthui193wYClOcQMYIi/aup6/HNq4hi
jeQsbd+uzN8N6yengNCxjfVmE6sELMt1Il6S1tmIQVwE8+s4o0xPkHP4xd2qXJ66eTzhcK89v16n
b8itQq0ChICmd3Q9J9iNGTkaqQcTkwK+ghQhRgNs3NE+bUn9+jkYKXu2+qO9bDccacjPnMkNbJL0
j3T3vRytF44SZ/rqYAeXnPcXPB22R58/+nkCJ3/XCQdKw+bzvHVnKvTSdhzWUOaFQ+p4HUyIu8QE
MmiRxm/EVk35y5cB1vhKqSR23hT6LXfopCadMAlg9R2QPlm357WclSFrrbjz4rzQeFae4pdY7iYl
MP0N2WQX/LicX/f8d6PgyDV9Dqf/xIzymSjc6BLrcdGOaxziqWUulyDFPZHwtxiCz0WJTVPR64mi
gE5Dta3NjvT8q2CaZQCxYTRITcLfn4mZcUtF8Afh2DHxotfsnQfc3Rjby2ZmNR3Z6h2hXBZPvNgN
HbRu0xGIsN4Jn2+a4a3O4XFfwjGp+wNXpbDNCkVplwSkYg1xaCQipPVglHH/t0E7JNnAbdmaL5uk
6YP74QwvRVvs944wXkEcLMUTxRyO0vsr2xL69PWzTJedEPjcBfX9LpRaONV1QlTHwXhFTFtwuk1p
qyVL23/ru4fH5WIu+mZZAg1uuUcHoCeK+kweaNO6CL8l0hJo73qke5D5BD2ucFc0J0cG+N4eJ36L
kTqoH9UuR5LoWpaQ7ZI9JNUCPim9dlZJdhIyfc7SFqCwV2Z/VXVQ75uDPpufVTWCbkATxti9Nrol
3Gw1yP0itlY9AEae0AC2zhsZa4OMJ28THbMBagP5baEiC9hjI9sLyUcJH8lr/3qSaqF0C2yauqnR
7YCEgVF42qzvuDavKt+Z+9YaovyNKSQ+NQeeq66bmG4ulPQ/P6lq1BVkcm3Zm/n4xftiBdaCIYE9
VHbsNqDS7kDdCPklOt4qtleNyFuARPAnb2dc27VJRjFCSXccYYMuJGoraLHrEeE8ey2jqgtIhPf1
m1UV27hNwBx4iY0hj8UXcJkAV4BySLYp5aIbDZSrb0vG8yipo+/8FA6Qzln0noxZ1dQdKowEi01e
WsuKSLgXChrtX9+TbWpaZJtGRf9dBGaKok6KzfU9ecKgYYpFSRTOXrLkMhr9jh9zOeqZTlIHxrBJ
R8vt/BHKStQvR5q+cdAtrbzIEZBAHOuI262XBBay3UPgk27MqLFhmYHLYP/ExKTzNcMafuLvF3VM
auQBOaIzA73ADSeN8f/KDRiZDqo5nsv8H0nGF8KVJqyg22yqAhJ6tzxBskzwhTpTy2WaAm/N4Vo1
lgL/RMaDAgGFBlDQ12TMaghZWj+6gcMwkTVnr2mriSBKFTl3XUCJqDz8nZHqxDPzY778mpD9IAPZ
CgomGrmi0kaYlW1LNrsxxI+HzPFeiE50j51bfA6rALmgVF8Jg/Z6PBj7gZfipS+s/fORwBfqzX5h
rryKGc+UBFDQBpD8W4+TMAptwwopS2ZNNEfb0eL2eGjfXaZxIDKtjY0OG6P9lsRmOUaKYwXtvFXV
LI6PhWMXe9GdDXAi37FNoOj+8njP6gq0Y0KKeFvcIsrqDI2n8qjKWAVAzS03pZhlPSkC9tKu/RZa
GSU+BQ2781Zea+x5kQv6Go/1VShGusA0FAql6WeEPcK+R2sFTAFyA6ytDHO9P1K5raB+2VyrTIE2
mZ6U7V7y3URQK5hLlXk/m/AvLhjRyaVwNrnZcSEUWiu0wWMCOVgshkX7EhW51IIi9cWt0R7J9zTE
AmuAHIDvhVNSksuKP9SZPmw1nhEZaYrDleKRvPVJFyZE3wiKoi9ufvyLt10RY6FgWUQK3JywRLV9
AKHnsAPAlKQqWc2eE6cIMP6008LFRywhBNBnRqYsNlDHfWkf1B7Rc12l3MSpEhdlgdJ8mbiAxd1g
TY6RGVJoQeJfuu7bKun7rGpZ/RX1fqT8E4N+m9bmVBm4KWvC14AmsmvxvQFYZCxM5vcYXgJDZAX0
X7H7cGJtbTJclV2MG/kKbsDWVmE7juQSbwMLPMrDmZNNLyVkiJfpMLTY7iCoS3+T6iyqj94fhC5q
Bw7YiUbxa+OggBCGaCZdGc5A+p/UPZxtTev2FnQuVjp7vlQZJ17hox+dYw9qv4iS6lyQqg/GPOEU
ZLpLhplZDMuZtKB8bDQmo0DyG8ENZXqFBM99cHdLvvG9cweeDeTXLau8VuFye5freKd/uVAM/8n+
2v8P3Tv1HuDGAKnJc89nNZTE43HVIWU4KWFlAmZu++hBbVQ8neo8duYGZTklog3jT5zHiT13IZBQ
gHxb4Er1Dwrcl7dqvYiQg3NjgkqC9BfVCy3GewxxvWlY1eG0wt3mzWQhBxTBO2XYrV3XzeTfg8iT
U0/+Mo13mBadgkqF/grzyPWTwaGgfMjddMn9qM7zMCmXgG34sar08mfwVNBqcUgRg0VLt9Or4vP6
QzwTkSioKSHcBttCqnjJKabt9a3sdYBqyvVDS/tuwbMYmCSdU5Ok6hHS4UMrX18j+wnFBek54JsZ
Kdmh/oUFebNsUsK6RSITnxhUKIsI8fz1qeDZGGlThgYUjaVOPx7Lz3NAubDMYgZAcOlNgkBJqb0s
5cmrG9C5E9JY2scVfZAy9C/npo2VjSfLnK3p6UBa86f4ZH6i85YJKOYdg36Ctb/7iyMEKYrIS8C/
iU+C4BDaqdQIlPRvo+3XygP6yw6MF6CVHsvoj7dEZzVMW/VJIiFH2aYyxOg6A39FgElX9ezidh8O
0/06LGDuomv3r2EOyO8GNq7epAZyXaHXlmiTzdFjKT4vk/zPAN7ONwD3KpG6rBWPvQA5xhNDXWT8
4HAYDMITokp3JARgN79tqJ2/TyIDkA+b80FmbzYhRs5iLzR6V47X3T1zISfWCaOS0jBSEOxvKhXH
i3EZe1XDUuytULij1QkQTbREq7RkrrfeN9Odbqpg9U1JFHKXwzKuYwq9PaxLmOK38QUhXH/wz/x1
4EDuroN+/8pVPbV1gDhQQKZqIkR8nL1KiYDDPX/cy1wvs51zEJqlHUSi9H8VwEE4ZUBjjiO0kDZs
twXGRcuTROxFn1g0eWb08lr09yAdO6Zh6wmKcATZOD1nnVacIOVXJtLsau1ilPg0YneWYp7bSj7h
gS5mI1pgx8IByrfdEDwfddNhK1VnsnPB10T8y3dIZ15zY38Tt1d0OYvWCvw3HJA8j356Ss5S/VOr
09QTd5SQ5VdOqi8HzZmgZTBEXbLsPEy9eSGA66JmJLyiqkBaG1Fn27lkrSDi7zB6wwFpWKeDWFSh
zjS5iMIUzxLNw4PlZsMOVeDthF0TNJRLvyg/c6NP9mcx1CfqT7yZvflWUwVq1g66e/H8G/vejYaq
Bjlek1E7p3swA2Rwjb9QWm/sWobYJkRMFvdlLvC+28VyVn3u2gnyiwec0AWs+8AQ7uHqJufqBMsr
z94EwLrnAa+92nnry6L0YYkWY+tjI+XZJ+WEwrqbAZSvKNTfVJArp30C/iiFahKU1IE894rTxgiB
KPWywi1KPoLf/oMxdt2cdtQvUYX+H5yQootRDCCnhSC2rbCRD6JZZHiBW2MpNCD8OCLpbf5i4cuU
yfbn8B+cgt4lCMS8Mkd98YWb5j0mTEKw0sYHso8g1DUuO4GRtwObYD3oIBmUKNVoNJ5Bbz3HeEaF
sXEgUOKEKLVfSbt3DnqLUWvYifT2OkoFo0QCefjjyqNkJGGxT5iEXj7b/rM0YXH7W6Y+R7tLCaQx
ldc/GoSfVlMGjZibbtSkXQi+XKN4C44rf8DuDZaz8wyQAt7YAljB8rq/pFzVTd8qxf8gd+xIJ0ce
/j8ySQfOmhofzvS54f3gKGwFmfyUjW1yJELFdjSDs7p1avUr0bysZzytXAn7iXi0KAl0UqhKLVfQ
ZEfAg+PU451uIoI0KDDOL1rhlHIiYWMmYmrm7nuYT7IJE6eOi/udsk0Gwskb4td/xkPE6eUgrtuY
jPnhJ22/si2SgdnHXenClqnfH3m4KIw2QriYhM4JeoxtiiBuTOzDTiJdCha0XYcWHzcomTTeRUjJ
Yd2sFp/hVNlAkj8WkNJm5aQ0Domn3sV94MMMn+t4I7si4idI8kOPw8aBT8OZCS/TMNNF6di52otA
lZ77ixWs2ayXsFBER+dtCWI0cp2fOSY9imotGnVMSESGdx9FA1ppewxleRG+BJGvIxGOpMwwaYZ8
IS7I0BOVN64L3OSC4gzRTw/zSszy98QwLuTC0FwBzj45rZTpGqYRD+QBnMwzTXRU+MSLAsePMgfz
/3PI2NWrYUXKqeaw9j9VkX0cw57pcd2ouzWmQdPbe0u/8NMkkmf+qpKbcV+fmswfbgNB4mST/3t/
sdezcXYugBshfZkLE0FVrUfsS+Dq8oE4SIieQdssX29M9U+yAaT8M1v1gh5UNWYxx/EB0/RjUodv
v5EJFB3GZlGhquMTfw5Obd/U++HOkdRHEpJFHNMPzNAKxFrVDuNrwqvtCvYzMcmZemxYjVJEU7V1
9FdnaM5IN9j0V8eQXmhI4ycAbEk7JmgXpNczzZrURf3F1/vwuKRPCYtWWVAi0TUBFKiSBg5IcBuI
TFug5CGFobkTGyfwrNYV5CmDuIORozCnAB/vvnKqiLQON2KJgudRDa/pUimtrN0vFQkx/VfyXDm9
9xGSnBhbie/HfWFcS7EZk4P8pnzW1T3ZeQhMnUPJs60EgjabZRT7uRuKvJHR2ys5GRyqPn+gj4IZ
mHfeUeGsBBNiz1hMm26RnYcS9RdiEO7P2kbrke0zIopsSkszQeYQt7nfWaxA79r20UEpKFQc5s/q
75N6u7ZPx0sLgr5RkCTnIQQOde2bisLn3G607VDMjUZkdpKoDsMlhAhQAtsunQ86j4W1p7sxxOp3
qV3T6AtLz6TF2ks94SCtQ3sbbfXzhh7Sg2mnFtJsSzS1wRp2rrDleGexu9KKiv4a1wnhVd7JXFsA
SdhGOihIZq9ZUTpCK+0Klbg5mouAuCb+/lus7tX1KQNDbkwhGm6WMU54YSv0Qxfe/CAP2XqrldlC
KJw2CmU9BrlhU3d00ppIy+fbvO1S2/fa4d2AVCoCMn9t1CUq7DWgj0CVf+dqfu0iJdOb/TwziMwL
1lOpKQl+YiGzIT8HTNVevSbAVh6PH868vl6WmzKSOYqzC5nyC3zDXOE9m/JpO5quTWgXGlH1hk+9
DAc6OBc9/K/oXa+rfoenGM9m5q9O41QZxx8DPwjubWE9PhjMkxmSSWlQuPUdayRQ8U6wZLgdEosA
aDvJqeRIjXxPoc6J69xjS4BCO/z15OGD6hH+VPlD7gimHSCZRk8N8i/ksip3Fto/oLygrPVPW6Ei
Z+Yxzv0/3D3GQUKoZv44SDdIvwq+x2tt+JzFMW7/CPzzO6i1m+4kqsJ2Sc/mLUp8v+VX3+Vf2ubW
GP92hOqXWzE4CiIffwT+UPxdnkJXJyNsrw4N6CmXAdqIWf2Y21iQt/HlnKR/YjrY/1xfotdqc49l
NWYKkrsn2hVs5XX8ckEFYTTXe+lSYjvFbIpRATPoe7iBUXegEx3vn8skFn2tuMeIhYyxQQvaTGgL
kaFNA2ceHyt61uujyBNqwB9H/pk42nGeR29aYueDlnJpuuVldaYnUCCLFR2TmKDUCMeSTjVBd9Sj
MeOaIyaJZNCgd4Km367rKTz3WtSkbmGi80CjVYFLrCFa1mUGs+Yh1TbbzVvPs7HaVEYFHT7dzjF4
H8z+nLVJ3DD6SnQJMlJKdk5UWdihvK0zAzdd8bppG1FE7sT4qWk+rPl+R8/dVBhYOWb/eITtmAnZ
l4FvcDEzvxyUYP2SqqINGzDPDzBb6TE4N7ODMu6zkYR7M6lNVBPoqfgxMciqNHqmuChpaey7nsSZ
AAZqQnmu8mTwT9y/2dwI6HN6jxz82aETy6NNZgAD6IrikPOv4FNxlrlAgCvjT6Lsd2liR5GPJ4aD
XMcOAsEgNHL8lheA1u9rPGdzttPCvh5hkHGwB0zhxd+duz2sLJWa+UIkAAF/KQCotHA4LljetHtq
m8otPQVN+XySoq6bZqC9lPFVeefVZeE6QzzP1eYZIIfB129OVVtazvN1yF9mEywCByva7CQGKjE+
shJNCITyxSqeH4NMeiLwbIOCINNHfcA+hV+ABt2qhNJJd+Tfu7R8LMb0T1xraugDRtdek5oN+IfY
Umma0k4MDnD51jHtqCAvX9WzMdcwlyNqUBv/zTpvc/3EXgmTd8nnxsISnlFaH2ve1cWidkrfl/zd
xJvZTNNbSK0HTiAggOl6fwwb0MVxezs4EOCvSGLVnKvDtbHQWJBqqXtrZZXzz07VORwBJiwVen+r
viM6MCcV8Np63A20pU5B9o2imF00OaTXZTcd8R6KLHjsPQZu6TRrT3fC02frTU2uLuH7Hy4WybeZ
BIc/KnJEjGMJqZV34/UMeE5eqPEQPpFS2O/SwV/HquJX8CdBNyYsM7MxvwRf4W9uwLSVT8rKYHNH
TFIuO85vChp/+w+oqeEeorTjB8MAOXZqkMy0XUcG9/kWAv+davr6nxWHVKUWHTN1PQ8/aL7XYVwM
ATynMbo2NshI1BF1tr59dYawkzNxyd94WYMAR9iLUl09KlExYzip64FlOgZasVaDSd2liFAJo1he
wBDh843Ks5YCIf6h6b9XhbewGizs576a15qQfYfj+Tyin89sBHu5YNXhE89+xtcbsGq0FvQGZqya
Us22tnhcSazsgB2MJxIPuRtwNBdlz9fnQHHuqBiHDagzjOQexM5a0nwk5NOT+4irnIZWViDRFx6I
7L2puBAeI3s/n/X9cql74wW+udRI82zbr8xJ1V0hTd9eDfQ4i8h9TZnAd8F2QE6+zqzS1K8q3Et8
QZ7C0i4Ky/9UpQwsGpMHLIyMu7HNaYLoM7Ft6YzuOn18SCceA/SqaPEFc9Rqcl/P+KyLU4/MeFUX
0aebFiqy+XtFaFA1ENqj6xz07A8e5pWUoRDaEc6paYLB/PBro14yRa4NbgwORBnHrcLkLUbNSxW7
IMyJ1eEQN+u+HQOJPP/xNswzuEHXUTz26uoj/vx5XuLaZyA6yoMUZLW9KPOtsRKzj8SE6FTqCZPi
U2ESo6OzZzlerVZ8FgD0nj2p6B0PZykn9Louma1I0uctNyfZH+TWrVmv6rp8+EzsZ1dfMjv8eAsR
Igyx5QM6WHbP4gDHH1bP7OypvCL0pMGG/Fg1iOyrxI1UVEzDVrTAIjOaFeGhGd8Cdaw2OKPjFm1J
v61qFLJHv3p1k0aKOSuMIwOS9Ml0VW/5GueZsQoZWn49y/skPOKrTSDzpUAu5OeKVSreNyx8w8lk
XAVUxgrUv9AtVztxhgBIqwnMJIjW8n+Kql34ubUOpTnJa92GjxpOzfvuFb0zKKAP+qohc6DEhAd0
y6k0imjnbMKe16CqRrVN9adYGfdQMdimZ6/JuNI6BVlLZ0msKQ3uLuERjETobwR0zmoAn5uzY2Jc
jPl4SpIXTX21LJ4dfpt4G+0/sA7NGq+xsDx0kMji1cywV8A4TbWXx6J1kKc+8z5LpFdiDc3GVwvm
bfsfriHJAZpfd7EiAqP6JCx1HwnH8D6V7fIpCkjtnA2sdfGCEdUejlSguL4XyukGL2IYPXkSwQry
0jgwUwmMUqvQvUX/4Gw3CZjBayprLVHsDynjFxT/PBCd6Eiv2LugJqarB4aWtFwrGuisqhtAqeA5
1tDX7In5J0UpBz6wmXqO0UwvZABg39ufDWuydeb6uM8a6feTJEKE7kJS+V2jPtAzfr/p9CfIkwR5
zfUcHxhX1x9az5yWxF9rM/pevKMp6USfMM+3ueVssE4P02NTSbp2LhVT1WEa1CsL72QJkIYbd7Lr
c3fcSW1QL5ph5DMTyGCHIrPuUuej4rbZZbmVFZ64l4OlSEJ4mxoWYe4IZEDbc7kIhHSuodSCKDMh
/fg8gcGg6fss4UtGfc8z4ePNW33F1ONhVztW74uNYsLZP74yqDbiPE+x81/QWqo/m4aa2/fAwRGD
r7HWfHA6jATW6tW0vt3DaHpcbz2D/f1YyRhjDPbKKMCyIrFwEKkO9RRUbLosEZAmptaOtzIffBmM
EkemOwtwsv/2lWiu17JhM70B4EG3Kq1CKEd6Cv3Vc5NXhzEQMm4fa/0j7pd3sZ1ck7IW3gvClHvH
/tLkdxlrn6efAcz0IhC+EEoJBJPr50aMMJwMb501rc0WbJP9GKJIrgo1c4TcLZRIcoj2W8OXtycx
ZWvguKZhx+s9R9xgcp8HshNHm4ngQmITCkdXlTpckhH90XE0uCq4XNiOocsqvNUzELvVUcH7SKTI
ctstNnCz+g9c6eFz5H2g45Sf7N606Oww2SmarAJ6kw6uh+4EkoUR0W/8rYGCWsBsWGo6XAx2FsVF
R1363nPGpH/J0gBNzI08a8WM3DaZ2AYURwLxqTOExTDN1EwVnQzQyvcLeXJ2E1ngwh+rFV6bGbX2
sz2CLefWHloWplcHcFHz6xaAuwoJo4WqCU2ertDQHSM6NbWeqhawWxNeOrkyPyAcia85kg7phaUU
ZEaGKsETJ6oaeyHGginikKkIR5SCXVhtrk62BySA88h9FxpB/0AVDuk0FA5dbD0e8Pizw0VeZoY9
IYGJE5qB7W5hUosPdZETYuDsohXehwMrUkJ+f9lbUSA/1ALCluajgMkWTdycC9WKD+JOVFd6N5TB
/roh3PersLvjQgJ97agBfxNkgr4fP6xRru7TcnrbBkcNOozQaBIOaQx4fxAe/qxBv13mXKhNtxk7
VXQTD3wJsj8mVB8CONG2AbW8E75t0GZbh5tkW7n1L8zkcnJ2TO/OY51F/Nor/FJaANq6Fj2xCHkW
sA/lO6Vhkv84TujgvtSlQcppOvBxxysi1rTMnKuKKSymatSxHjd3sVd4PtvtQofgqE7vXvVfvAKk
3olVw7KZP0rthWUyitLGU4Lmm5Q/Zf6ZtCA+pqaQVJAZCWYtCsfL9/bdWOodIxQY3xrsstx6TMqQ
Z4q+J0sTgyH/ZCj6hoKXLUkKeAORVoaJ0jEGkLQ2DRrD2sx5SPdX68vAJy5hXnolBbXhZQx+2ZXI
P+ruJT1wnAKH8pw3wLJx+rwcFfILqZBH9NjVXNeEM8fczwihDKcFWdeEtnrURzYa6QeRY2CMzqIl
gVy3LzKPlC4ITsLEKBkzJuSy2VzAYA6W6Q9EA9/CQo5P2IglyhUJHAaU18Jdi14u9PkecFethxts
u1bt3Orn0CGpGQ9+Fv5WPNn9/NDWIuPsQq6eceQT71i6zmvWUbOoSVxFAn+ScU1Y0K4ncZdMEBMH
RzMwWcY8k18esgQD+w+n8tq2FqFKVZl0cDjR+j4x5Mi6jKjTV574yr4wWxtvCxEUc5E2KpCcnGgE
W1TtowTZ2GnxvfEjfQUMHmD0EVzKNDX60qXUm1Ptvf55r+e9X9VlXCrDR7y6AIq30l8WPjkTbiAW
Tc24Z2vuuIwzPvjN0IGxnCkDmr08XdnVBrqlHK8L7vwF6Zxmoi2h4BykxIWguIe1KnRC7hagvTOe
gkDQH6gBKEIRZBEngfX7SbmR3Q3ubQauIAQHKIVFsX0OJNuMrWRE/56pxs2I4e/Cid5l8qRiMNeF
FiAsfzDY0F43mTl/TJ/SLNThPq5luCGT5W/NoxhNLBKr1h34uhSLYPMVBmhoFkR4LTElqlAuu1Y7
zbcR2bDFa/ql0iu6HdAeXW4FRRBz0zNl4HdH5H6/32K2AHjzJUZRMDtfbR/fQ/5gGnAgO9iz5W6o
XN8t294PL/mZCudXB8GnhYRPXx2gyG1L/Gyqm+47xCuGMtNm8HY0/pEZYIkr2GdyPeLYX606H7TO
hXKa8mlcGEtSgycV4zz2Xa6sVEg1t/gIKhtk8YGcZGPMewUKoVmtgnd96l+DWNHwamU1UX5ZU56S
tAEPnzufxFG8Bz9jkciDYLWmMi7KObTuffaqSLsGp2rY4SlUDjevdt3KHNTYw9O46ADAdGWvkqZE
b6bfNMWlwAAKpaJ1m/cQN7E9H4Ok++geRnSI1jL5+eLdophQssQZO1jXUqYFxlAYGPwt5GXYw5MJ
gB5fg75inZzmxOs0HgdEh6TvIsMz3wPJds5qZFTAcEzrogRClSeXN/s68NuKCjja6QiPUbSuU9tE
TEVYQ8DouIPqtWIERg+sx8Wb71w+2tznU2wDVJ6pT9QryTHpTftEehrdK28feqkhlzmjIl4gmH/y
A19JGvwuMj8iTHxbFAY3ZmHnz6VM/nqn5DVMzShmTeFodNMv5LXVCjtp6h3KA3wy/PuduyY5ZgLL
W/PHN5rq57326Wgc0hODeQDrYkYnMRvq5zGu9NYCDlbTRZUM/ViFYGACLCrtVKX+XnBzvzV2+ndU
RSt05ezYzyCQfUP3y0X6WTLxJXFPiOSqW3V7zoiJ3YutRmQExB6Sz5vAiu7QA+UoukP/aqlsgdkH
j8PTA3NqDeW6dmQ0sncSZffrJpDrt7aaGklTcW1i0Eh1ds73XtMhTYp3EGC+RcLTj7u5jZbUlHUF
G4ZAsPB3nBF+a9DBnlvpkI2EMewLOxk6abNZAXpMzTbBDNg3TX7bxReexKGc8RUxA6GrxclJeKpy
KRGlyjbmcsQFyvKL3quDvjfviWGEFtIx9IMhty/qRiiFn/YJ+URXjcbw9vdzN/yJxcUlLUFuM59C
A/llTex02r4g/uKfzo9RfuAplO71HgoKdyZVbEmNGdNYotVDTsFedpaAskOZUR9wZcvkbJXeXNql
ykquq18f0BFrAu8K+TN1Wfo3OFliNARaFipy75+havmVUvDR+dhpPYQGIMKxlNBBcvhqFej+6R+8
FCKmkjh+RJh4Oy9t0nlpoiEId/r3Vw3Bck+OK8FtBuiXFG+hkroIbPC0Hgt3mgSHQ7hhKIFECvtG
47AR5HQQN/2gtKuk+5Vp57YK7aPQFvoqjNAmwEC8DK7Qf+pNLpyjQ/FJMoOReWbbKHOm4B0w1sHP
BRKMFEqRU3Hig3mxWYnB+0K6qkEUbBOn0aBzRTGRKqIUcHyLVKuFKwv5tGRl+b2OblgmzJO+GinP
CENBONyOIovUvqktT9eKlju53X6h22kaAgI542Jgn2HOKvtZl+XFzGHJHWeP7rnG1PWgG74kyoR4
UTNk3NKlwF+YnwNC7T0Tnjn4gufsxpk/71Ik6QTFHzVUKeYR/0ak9Q6hptpV90eIhsEb90FNjUvh
7q6Ib0pYWE6oKvSs37K50kq92HV3WkqzsveDvNC+oeF3GRBWfZCmDzJoztmTx4RIH4/oOG8mYWjl
AufLgGIhXsIPYVMzlFN8f19SM5lH7GeQjUPT0vUcs2GsM1xDkQORe/7bbX6GWEsgS31XAvCFtktz
nnt1LZeFoF+tFhuyy6jWKwS9AA7D8jEaEsULZbvQgQp0YoVxDprzoFpHq0BSkeCqvRWeGIybGYyx
uqrRvk382zToQiINN7/w3J0tzLy84ASLpS0JCe/cS9KZu85KWiWYgOb83A+5Mzlm+YKwd/2dsVUl
AAaMKRxEdm+ARYaI5qn1PZbwOQloGzt8iOBfR7i8i4DkeGE8wFNkgVCaGacbvN32/sIU9lIG7UjN
1165Eu29tL4IWBfv6BQ0kI0FK5QkqbNbNXw7OQt90D0IqT46bwQW4DIB9TOvXKL/DM7xvzS483Ga
hhyvAODU8Z4EE0RAPYiVElYeA+XFj3IWgapY4bVi1BQUJjbN5IpQ9kihR5FCB70oQ+TJAOm1Efh6
FmRdn8QiWsnv4JR5XxpStyphYckl3Poik4Y5En9jIsRkzM7obFKNFRpned0hd7n5oolLyWJgmBhp
TmGU7hOElgtQs6zUG/VXdokRUd2Y+yROhFZWrOo11/dwDzC5yx+yLrIL3XDQNTzF3bBlQkrfz9Jt
GFMbb9ZJ4FXbQCGXc+AdDGrTaI5bx+EdpgBlgDqWQoTal1SMKN6ys78iI2ADNFMLtyZPemZyM3E/
PPbnGGHaZFh8fTuE39uwY4IzwpOhPdl1Rbg4Dxjsnh6jeE7xpyyRnvPHgSaZ1ocew9aO23NmsEpz
mLPVVDxbrwMM+VsVoWhbrjuoxvtB30yBBPXBAVFyN2CmfodUnxHXXkbv/UDH3RHKIje35Ct16RMm
KuSdXnT77fhEVIAXurbt9MpIhMVhpSaBx0diXuzPGm+lVnqx+J2uJj12QFAkxksfXbVFEbmg3HXj
0H1yL8xMuxQp/ttnWGl2DCdIYk1PHcDWbd7UllmTTwRYCjiOUkm1esVA0WJBmq65ae7U76BgRe2X
Po7DWwd1cO9fWkyHYsw2B1Bcw/s4/rhcHiewLrNg43JOY4Fo4I7R52JmBNjD7tCci0Aw7kyjOQ/W
FHvzD8ksxUuQjU+6M8SggOeUqpOg7ILtzzpUbvTXXnQoqud2XuFiR5y1F047XrxXa1nBRy8uvHe/
Pdi/cA8vESihq49cD7CP1o6xo0WrZcwMwC/CSNUQOdNaqgWilZ5KxPc8X9ztCc5kzQsn9QL9q20f
GNyg2qvog97S+Mmo9U2pm3vbEPMj4RpsnpYiU1x2Uy4NYUmQNj/HmCBI71BhRO2DkRAzMKTGn1a1
Cd7JxCRbLl+zKf6TJO3DZdiql3A3PhEJVEqEudxNdnalJp4blRnFIVXRcBJ1NOx7SJKOesGtx+lh
IucJANtgA5IaGhJbtNIklRQgNaRmLP2Y7VeMRPYGMNd/bwe/hUAcHSq6X0duIap/xzlRjNz2yv1z
9oEJ+7nTBGPKGR7YoE+RQVkWwYzh/wzSxbnlBWM17+ONt6RtHo/06qu0swRo4ro3JkxbmxYjuwBd
fJVBPSwylzCl9ndjzEBL18YxesxejVCqjKkQog//X7rxEdSRxTtiyJI3Qk7h0oGgJULalxwRXzYA
TbBl2qImIDP/Fawbv81C/Z+q3CivaCZQhZwea5WMcrMgXWAY4HA0q5blIIepmZMhB2G78u32y66D
jEZWmfV4CB811beBUk62u1vuVwi7XaGI5yhDDbQTg8V49VLoUtgebAuMOHAlSYxUhRIbRKKSQZaZ
B2A5LRN12tUl8lIGZwWt+CUsQYIyRlkkjwyNzbh9LT5WyuMvnHhpdHS7WWC3+1tLrNtoxT9d08DC
dP+NDU06IbQ78ikNWcHthJlKLFYc3UFjOdhTqIQdprqup1238/+sZs5+R1Jav8p/M+G4gvgWVSIB
Xuk+g6mZLj8gsUYZ8Xuit0Z1rQHQWNHlZZBRwEcDkeAccaNsXJOHvVSjBx2lWTCogpQ/2SY7iD4L
rdt5tF75NTkIP/m6SUB1OUTZzF1PjkBy3Mz5y4QrwGSyvISoaB4PPIvtz7gWUMtZ+AoMrP+WoOQE
/+vo5379dQKcFMvCqmgcMGBZVdCDaVrH2om7TwGRWMzHxDtQOHAIt9KSehXCPjKpw1G/SvvdYDbE
o30KQNVUvAzXEMvMFtmIXwS8mKgXu5Qv7MqYXAuEXC/kA8mrMaZUifRsR5GOnIM4VLuGRYOxWoJu
SRArRHPhrEsdpGsuOr7jOfm+3tAka5zptBmj7N6DtXXhqD3aOTBttpsBmBUV+M5pTtQEtVWFfYTv
yNt1Oj0imj7IW54FXyCPhRs8Gtu6/jSkmQzPpThPeWK00qXS7RLlcAPvba25kibbZ519YzYrKJDF
I1EXU/burXhJ6OCPBG/v6RahDoeP32HMT2k9X66WSFG03t+R7nU6gq0mrS6t6chqoBVkVlDj42BO
uyU+CSFzxOIAzboXDNX0vbzHCVQXdBeF+DvarsmvN5zdgM8W/HddE0izDIzmgBgWOVpwn4udemQw
R2N+QFKvQDBYBQnenZWhWII38GSMxyWi/vDOpyQidx3omJ04TnTWHcm6uVE2Qgq1HhegA+I4cu6m
44eTTBMrv5kBYIAA8oYoOx7/v7mCpDSCjII92jEEqxLmUAKCrHX70xt1P4rRN6LQzJyl+0GSTTPn
xBascWPqJO/3fjzEqlnqWdfkLeMQY95rXMoF0XNiGxU8KM7cf80z4v4W0Jz50Q9rkQ7T1zcO7PqK
oRfIzF/ZUqg2dLvCbQQ3/32tmblSkmsqb0Sjms3ysUuvxQBsZ6lE7obWWltb10iSs/zTIoOXHA7t
V0rH7vJPp/APT9TnJN+9tlI49rgFbYtHkZDOBUP9L7n8e3Z0i8xLhkFsBTnH5W6M8ILeZmHd1zoo
ZXZCjHyeR2H1tV2Y4L8DoVhOk5VCefA/ve1La/q2DxM704FJ/Nf2RNjM0qTyCsr+htpYUW/p00gc
e/7HBr6Lb1a97W7l0LyDZ2xLk/TCblevm6/PO6VGCgbxlJj2b0n5aZDbxPHH7qtaJzqkyjmrDLw5
QUxRwYLB0mbuWW+90p2l2oIYrCSJ3i7qZDDlf3o2AzW23daHLoUOsCgM4ArWfwgukz9zNiXLWt3v
vgNqeh3OYFu1GYeWYn9moO+prv37S/FNHTS1YX154g+QbUhiGGzkNZf3EooHD+bwNwpcluqDW1U7
8PYQb+sX7o+U98wnqvdxlYA2OcJGWnfgxLRRRELbHZNgxTVqCKgoNFgqf8eOxj4LncsbH7K2gKaL
0bS+U1fEb6iR9hKQUpebt4ZhECRMo0gyhGjY+cDSsEnhjmjUYQbJoiH4hM84RNcYDRrdLQcaZkWr
xiIu84s/c0Mt7xQ2uXjyCXLgGdarIIM3OzfJVT7ycC5pzaqcl8gywUXQAhkG2gfAiiUkcPHzygOT
lRD0yq4e2qYEqkipU/7OER69tWpXSSgbJju6ulIeVNPo8lbws70HYrfwYp1u1aOrFkiTt2EQ0VQA
2l/nCRJsoLhNkAX8JK3BbVedbB9lrl4qIb6JPOgk3oHgmJgJ5RT79oQEXiRgJSuwVSpHfGKqlJP1
PDeYGuCNPdvOrv1m7vLOnJLJoL6HL4AGgtjSkW30aGRcZinKL6PZ/JQwwymb1VVwatE/pg6nElvH
rpJ3DIhcS4R98RxOw5VWjUV/xS6VmiT6lKtDZO7dPIjPl3QhhwL/DrYp688beoxudN2fGxg7j3Wy
A3anlEaltePICZANztjd2TGfQhuaI7ic/Tg8uER/lGvNcXWb+/9D7H5Y3QHHIOkr9i0fFhGXmunA
tAkByCCp1430hEROn2UlA99d85WA7Ty+HIQGiczy6sJOCJLv8b+0LoW7peHREZjmWL7EPQ0PJQq0
bFs7yY/Kf0zQ79UfAx20YnlycuPA+lxwIwa6S292QTiThy2RKGu+uyGbsK6v3m2m9Qg9T7I21Osd
iixpklvw6j0BEV/HUfT5AjL8LRMKwtiolsuoC2W0oGNJV/4bGSTJidjkqPxDLS07h5DKkWaM4Iph
TMb3JjHgbqNa5hOWIqRRD8jMv7dE5R9SEGgICt+LM/1bIeKLyqOWb9uw6DAyyb8maESAWqV+2rfW
ZWdZHybrsnAhdw6AFfdWjB9v0hWveXYRuT7Ub+P88PgO/kKsAP9A9A0XeJjNcdWaWUTFK8RsbEpB
pV5mEEBIECnNX6QA0xByBFn4FwIQQdxD5TfLSQhp6hxtKQwkn4K7mcY9RfPOK/ylhQ3s3SmJEN9c
DpUKp/2Y5vBVqVkclq4OPV/l7ZncB2PZBFzD9/Qr2jXZAnCT9v8L5HG2M+IPNHqtW9pzP0cUZTFA
NQSi+PVUr81BnTkYAkDAZjZXC07uwHm0RM9hA0RlySzS53eLfS/+XgdLtBlScQKqhhNcsZpSaWgy
kFrso/n3ZvbyaGeOvwwgHxpD/SWW+09nikaFLSYgddTU21lw6k/rymzypvmTD+D/3QM8tl08DYGg
d0IlmxFMQDk3BNDQSih3LeAYA8+4IQa/omSsqaB+NlqQikb0uBp1JfW5DSJuC0zp/kPB4cjswUER
7GfA2JPmxHEy7vEw1HkDkoNY6SYlLK+jrrRrxKpBnF9Ey7BaqWCSwLGfleGeEsWdXKbGS/zxgGGw
27qAftJphAqFXusyT8PGd6/Vdlt/dqbFtYtkmtxRKVS8+2lpdivYkFfqbgiJ4rblNS2EMETbhmCu
tLB9RCmyiAuU+OWe9dbxFpiRLflzQlKAu+KMlrhPI8NcfkzEDXIcTWxoMNgyCQzIpeWemKFPCK8E
B9Bv52iCxvD8SxRUhEKq6/Z+HTPSa/bJX4BEo/ieS0BLvGfwx5yiuiKvsBQ3Fz6B8UVti01FksxE
udPh+PaRGsBYFUGYlS+fZm7aXsgUaXovjE4d/SHyUF2w6k8epW4evIzFL94krhM/cAoAGTWRSyjV
8Fp3pAWoQ2P3vigaYl9JBb+Rha/kDJYG7SYi5SP6yolrWkok7OTXFOPrnRl0/M8ckYVN3TfGVzwl
6hb5+rct9ihfZVjxKR3PcXZDqDO14b4MFUfzDcVvw5PtNliRJKlxhc+ZvM1/CJB+vPqxRRX6U6It
a1H4MSk/53jxOjVWHrRClGSxzssbOt4tOnVftpvNgekcnG062Uhc00nCJ/dkRk6QA/tNwovuSP9A
Ct+sEqIiXIs6UgdWV1Pf2trKmKAaWL4FukfhYtenE8BdBe4X6IObfBlKg4QcEYExg46NoUXQrLjn
H3AjC7fo34qgMmpjAiorKxo3jgqkGAYnBfmOW6fxNVRDxNWLwDrytqOaOJcxZ8GMWGfPImYOYwBA
oNObOEaruuLlYtDHVoQB/mALla6FfWR1fQj18LQrG0xLVzjy/Kd7X3jWf/cUQFIo0SR3JPWM0PT0
ufXrrHbjVrCNZHVgT6TdBV+/iDXZ79rcaSEcfF1lwa9EeqFoImHRvY9vwDKn1qwp++emJcmE5YJs
lETJrTF1aurs8fTZgsny07Vg+nUil6Uy3KYJa3RplNfoS6ghmBSh/Mmn6KZMW78S3NRHAmWLW3oI
6PCzFYHs7lPqcJkTkudRulyxLy7H6zStVbNCZnR5mcShMo6tOe8MXQPS/zEHpn7FloxuK38kj5io
Jwjo8F8LGNoQPAE3OfZb4YqxTlTX6RxjUYWBxDMJEpvxO6GXUQfmHODfhi6FTnelh7+nxxlty+7s
/g+nvGxz44lPHDMG+fTorJAHyWbyTZhy6E3XeHHXBvHP1Z2/0ryP8dx5K2HoQGc1diw6yvA24llW
PM61V7oyErOz24pL+SEGKRsOOgRiF4/HZHHmijSWR05GWX0lJgSWuIgcO/dKX9wwKYaGlG5XoCf7
R7FoWNf9m56IIjZaOgU9IxR/T8XRubJgRr2IyKCJuEF2QBPd26lR1/LUcA8M21hxwp7dg2sijGyh
UfKAxq5nT2zuULCcCDpccVyJTYH9vDMP9tNhG6ma2zrIBdl9etOx1pubJp7W+MO1L0G6kDMpQOhG
npd0J1Gw1KTe49TKauGiwatZ7MY3uDfbt9JKIcMILzP+nybDPSRPMffUAfixwr7+/JSeGXxYgdL9
WBPnlioKVVXcUHytMo1P6AKbo7kctcRnriHzQiRzMBxUct8L22x9nhrN25Sr/7gnCgZw6SulwX5X
fQAs4yjqVsQY82gQ14N6jEFrzVFbnrFP+MVATEROx3rq0IVKgdLG1i8l4xhtgFjC/OcIwN9jLEXj
62bL+ssMJbfHNyQaP18mdxqulvL474iiEq4TpKLk0g7UT3sX1ybzAMqMxHcLAEJdiETsXdbnKLbT
ASFz7QXUN+jFzIq1MpO6QWl0ZstwNXkEkaToftHil6j7NfQCF0/mGXGD+cggls3mMbJ4+T0bYtjb
aq3ouhsXHNewncUULm/xhLHCeyT3LGWnnn/W+CRcGCNz2rEoayPk0ZFhj2GdSAxRb955hh5VQf5P
y0ZFb9jF5UoSq9dV4YADwyGpmNASP9iGlz0LPthINZHgAdvM+13sGdBFnYYqBTHKD+sdVdZFxN4Z
wp6QS7zQihuhshqKt9n3OmJ4JXjsOhfKXHB9GgYkHSwZcMVtjxp11sLaaz96b2qwReerMAGCjrkL
rg6NSYe8vkagUYdWMhGeeUDgYIX+yvGbsq88iez1cjvgwdWCfpQTiwy/59tkYAE0GbrkXAaF40hj
A074Jo8ZYjGblVJlH3NvDrrX83ZVNMRctXoZV4iYCXSIwoW7K4fCct7OxhLVLEFTyLB2Is9ArpbO
340AbPuVmYPKNxxYpumjTCPWmqDc2WeiGptNh6br8zEOOOily7Vns17xVBhXORYzKpeBQgihcuh3
vcx1bjzcB9rUwyov1P5nHKeRnyYApBtss+TcsGgL53wTnjoIW5DIJeuRecVTawwq6B5J43gGgWng
+jmUvbo2tRyA9usMVRxTAEaYfpbbqHGM67alqHaPyj6Hyy3A646Thi84yhfHupxBwBSWArZY3uxy
0nsI0VhrJxNr5K4w2og/D82EqGoHWu7W8N/Wrszd0p2FQERHAlkFkauKxW39S+iK3e7U1aRC69Lx
0ZKhzMkc0W16gQfZ4ZPVhfZbqkC14jg1jaeT3k95n2F6ky5QeivEKWpr9cRF0njNwesk49pPhgTi
wiji8aaNPoYJ/ZkbJu7QT0sWsD0OgbR41QzqwTPi4fWhx+kMfbVjKHrKo6WgIrRUUqFfAZ5rB2Km
tp1wUU4Jh6j2x/Xjrd3zoaK6UqKu+6C+hW+LSM9xhPmCTRZgc/pI09fVGBpCennAqawxzLhW0K0n
BJtH9FMOIrAyZnmfccmZmf0cNAbCg1vUPuc/asU9fca5aeHUwSDSaDz57VMw+FJsHkhf8TSM5+It
IhtC9oERYo4NSFzGroYt9zcGIln1KGarJpDyo9y/0Z1SNI5MTfMf1dCY4gITxPZNgnG6pvUW1clK
2MBNn3LKHNNjVlHSdoOsyIjCEIPt2dmpudPmikIE2j9dk90+TOi1VysD9gLJKus+vAIiFzahofWJ
AcgbMGGdWvjhZcsnc85Y8aqG3p7XyIoQ0AmSJbeGFbalHHoy6qf+tgovjL38cgd0rcVGHsI7p4ip
gh1c4YJfHys8JY4clU6y+2uwpnTnBW9D8LCb7SdnQCscMHfYjIsDKsd1svv6Sn3u+UCWOkNR2D5V
KOmKHHEKAaMwg8eHDrbn8kRnuPu+/r7RclKpz7zAMaLuTDLCjqY+YGNxzUP1A5APjwz2jw4WxCPs
vvrxkipX6Iu6W9rzxlavAnnQgyaNdpA9xzAS918dc5tAWtWXZDnuVzl1G7A8S7rNQUmIjz5jvNfU
OQStEITsX5Ul5GGZmdmOtqCf+qYxTM1KZ7ucJBq7afZ+Fh1mpa7Gan5uKyY8wkwW4h6AMZtlLzRE
UC7WCWJoS/QVLaH106azPQGPIaOALUoH3UHOkTgTy7xonFgbGZVRXDccnY/21E4Iu//YZfmR8+KE
IRTiH0hIbeqB+jj9c7sU40RpiTfq19299oWEgoSl6R7Q1fu9hJfjegrxLnJQxL5s1EuZIyNX6aQG
Jx6yKPdMeNIZoAWrA/Ojo6ZprdfJt54T+YnSrJUSn1aiqtLlEExGyZ6nYQcgAx8Tmzst6uZbliOK
jTgjyrCnEQET/VnvNT+WwsSk3dyk/ppiUwNIjcC3ztSNqIwZiVfZuvxRovcKwLVGBH1r1ahpJzAO
GdccVjcps6qiOvIvLQTO7umOinjqUWKgM4nmHBTl2Jg12mfP2+h8Fz8b2YebtnR1htgJimhFu1Ro
XQSozODTui0VFXX+zYMrSX/Lo6r52cRmQmItIe/NC8oO5z3fZG3mS5NDd0Lp7zMvEkSgTSJuYTOE
Aa1MGbs0ymBTJHLBYBqytixT4hI6WZ61QoCR6pvAv8Yu5UNb4/YMVdThesya9+lzxWkSuRR+VHts
cqF82UGpDMkjVsU4kAaQJxU8UPJx3enRY8wFvg2ZEPLOxWyn6uLbmQ9o7fDjHVkontF3b642QW2T
GhcpPCLZIv/Mf3+KJUsjRvRx039YC97zXccOUult43pYkevdXPvuKThj3ISUjpHMX+P4egREEUkb
3tmFYrDAxrSlr5Ur6a/3rbC9SeXU8tRt5RatKQ2Xyy2ektubQQdllhgOCPaE0SX2LqTcat1XA72C
nQhFHFEXc7vPkcSVMLz6iC1qHc4dBKZxx7jSHuWLpuzpkXSIFskFRpgzo+slhZ9Dhp0M7e4OjX5u
CDWwHIH+afOH55icKdn0B8Qvg6Jh3yGZoNgAnmjepwrixZxM5vgB/lNAGSmxj+1a+YG/uFtgB2AV
cFZH74IXFyQ1YxCWZHqOi8MYu0OnzhUVD5gkRNf7wIlf4ATGRiPs98Yq84WDOGNOJMRqg5U1y2Qn
E9ybtHDFu2AG546n/0m8VSZCu1v0Q4xLHmn9G9DVRmJsBSNfgi4IXiEbWrqXdnFKC35ICZ2cHPNj
3DhK0YpEHLXP3WoOfMOZ8MymoX09MZj3rImUh8LC/e8eQO32AAxuqnxIRTzgqytVjqv2WxcLm5I0
uQSsCbpxG3Sqr94AG0f5bR6KyGEMVyqXDtTIslKR3fFEHvaFCYp8pnoT49RAXAS9O7AHaVIDmKrC
Dt4X0tJ6nKwonXGPmRyMamiCqX1Gadu/MlHQfnVf7v4UcEfKHuOj6N/iUYpOWB5dDfLeUh8eH5Cx
AupVXnwfNu4q2bjcKEenWRrmd7FQLj5bx4qnvuHEWnADUB+9AvqS4H8Vgh9EOYHZHtFCcOe8fqML
q15BgIBi2CoOj09dtNoWAMF85kyKwQvko64Hrvci4gvw6Gci6qMG8B4sQSA3xvb47l0AewmN4nmS
Eymxh3JuTo7ZF8tq606J/hyaffJUQYiTZwvbEPcth4deW3OnlNVxxXJ38aVc8QZXbf0ymqFRZm2v
igqE2mt/+Q8uSCxpOXe5Nhm40+xhqrIV/iidopocR9kKuUVF9wRYZhyweRCQZnODDRIqlr6UHAxV
ib7/d4w5S7R66XbV4N39ja63VwPoljcaLPanRD0h89IrntlffB6KVWNsrhp7ROaCFlPu7W+D+fSe
SUizHzhapLEDhfqFWjgretwl4eYJvKYdmw5P8hYj5d29otHT3w0o+ihuYC4/71vk1+68mjNn9/Ng
Lhy+/9Y1J/wrARs6VOxsxN9GHyOOXTQVDA3PAHsEV5ZTG4KAscuZ4M2fZcF4qqfFOnRjQn7IB5ah
XkSkVynKcst75CM7sGMqA0wSFArDI003UeWSkpuSb+F2vGSzhGiFIlcfCcJQxw/NZe7u/8r6Uq4u
1ns2grt6s8rp7isqYfNOlRGAlTu++rOeu1uIwan5crqRksnC+cZo+4K0Y47R2JmYkYFscteLQsGN
pdyt4MIqOR4VHhp0uMrAoH8gS6W7sucoJv+Ccae8NMgU8HA38sswuld+DmUdWaNkdt4VDd3WIQ90
cQCGw7GNZQQGXutHowXzlaYydQi2Us433j971w/uL4PFzlj+GOC5lOdiZG2HcUCQsAvzXDNmVaSv
mZCJuDWjjF6CU9rKYkR3MKDu0F4VLd24EeqdJr3aiA2ihkwVGDdu4nSJCSiFYm6UMGlOXG8RUzHa
CUh7NceMRX2oM3afadYXR6mBptiAyQKs6L3YKe/Oi1HmCyTI+7G9btyrPXO6MMIBsaL/HMWlZTr0
V5u27/0n1Kbr3TmxM+d4LsjwpsG00+vwCtG57MRx9KMCg1KhbdGktXrGeZyPfn/9mrXiKgHpgwBU
N1CIvsGW5mPtrFOVMTnKoDi3XC9oPXe6YRzaIoRDRPbboqWJXxZsSVu6IwpX+SnKU83BUkHJxhJU
MDypAuf5L9UQNhYF/1ltL1Ed3kSUG0hINfgSBuYTAarckCvMXpbEYUj7Zq5h3Jio7MZMeLPKEJOQ
8fVPl71hj/QdXOsdLvA3nTiAx3nSQAoOQ+6s6w5BY2nEAmicsO48zIZivs7LNxPRJ18mjcn+iCiM
KwwT8oF5DgyOz/tORUqRNjtpz9o4/tiUqpmW2VL1s9p1h3k8FVpXu7QAX+LyMvLoNPmHhiB6bCte
0fokuVrGhr5mhFq1D2gF9iP7/FvFZQMq/AoyQ66EJD7eQkISJKGC1PSesGAV2KPCtiW68MkvkKJd
6HeFVLs9uf54cA9nnEZDMIsacBM99aTXYeuvQuOaLHGV6qVX1MCRhkYdg23nYhrCvQpmGQSei29t
73XBeFH0TmeLVw9aiQrO4TZ1b5k6A1dFdEWWGqP369HfJgNApQsXSO7YkufG0fL/0HejLthCcnMZ
NcQvoZxaQhWBVDO7UYH6DMENcVkTeQa3uO9M9YtxBv7V9iNBfP0G4GoS9jEvcuHENXZiUmU0lbyd
+NKfq1j4KuN5m1UczC/bIgHijDPLSYLx7d2bvwZ5b8AnFSJ5BvnRq963zZMYtd+pIi1RMNn9DFfD
L79SuI/644/p7xHjinQNE+UbJVzdZd/J2W4rjQTuBld+7ASxbtDrIwxdrBvA7dcg4+K87mWs7JXf
M+sMsljcVUcFDzGoEUN4u2RCucMFI2hWVHDujsycvgURK6YTncV0AvC1/4xgu9IRp/bdRFCGKPnj
E6BempoHxPhVwDX1SSfXA6AwnT5OJhbY0yZwsRoKuoYUI7YMoxsF8HXMV08onke9EzyV4Hf9M7aM
05tu6HUf8NGmkUiC3hxbtHKyV1TTfAjeuafVR80nvxSlzWvSXPnkLFpN6/ylmXG1id88ObEaqzVs
gUYBeCaasgHAKtCco+7VhWQz7D7WKV46l13jJiFN32pqaul/hkcRirzKJ79vKKqrcg658Wo4O3a1
IcCwMbN87SjSVIjU/1yO4d4JalGlJN0goHcXBRJzj07XtwrPdnCKz6fF1HMc/Vr3sgnUIQwZb1IU
Hq/+FYNIYcPf/ZYo0aI2Vfq4gUQ54oGhKDnKA7yEro/icG+yLyngZW+0tAa6HqI2bCH0cf2/rJv0
oftKkqHZOCe83DRrFk0xfX8xcSnDT47PxsCegW4ISHMJFGb+/KjtNSNnh/yx9F8xQOJDRjeVDCG0
FMI4Op8QX8n+5RoCfk7fEt4+0TJgWLmLV+VDFxotTkJlQOOlZelAlvbuJQ8DEToga1qwvYbmSoR3
q5wYoaJtw9SdtYRWuB4fBGiL54JLdDTZ/4VejIeh9ja89tOsLgY/Rj+KHr9IDEWu+bBIJxhtJMgu
4wWOrPqNdFxQtbcRilmpPSVSk0xuvq/IaMXd7XTau8eEJRXPZMI6fmwxImCdpMo1rjjY/9c1wckI
Uu6iCGV6sDC0cWlrT7Lvc3mxTg4Cla3qOOiBUtMeyKlHvpUUXOjkn3QrBaR6rwU9lZG5BBTzKdTP
UGnSUjdBGbK4QeOEKm94fynIUefM+N5nEbSelEfXlIaxUQp6rNhvZiKQR9RbCItgJELJda2Q2Tk4
Xf6En5qRCsy+rPpZXAzSSY5gXWovp6hBTgIdIrlw3m/Jfx9NppkWnIUi8c6T9q5PswqmZlwbd/KV
TisQgq1mYPHqzVozC30thgX/cg6RmeEx6GpT0XEB0AGntPVFKlV7Hw5Y53AXuwE8H/UUYwOk24Ec
etbMVFaTthxpzztc6NNVYMNwge9Jf/tk6Lq8bxrciwzQZ5IFUIYyPYbtIBOZDMiOhZDlgpbv6bYJ
1i4+nvCgXpkPQf7omJwu9MV5NUW94sjJYWZ4SITuWyfbkwGgC4YaVjCUiVbRTPttdvqiYlHgCwBM
IKTELjLYnbAi2hjQ3b/7X0Da3c/RjO9UnwGiy4bl9rSnDpWb+lNP3Ue1QoGQaTnxAjFcB2ffIQoT
CIOxUlr6z/MZN8hnVX9j0bCY9q+2iPgHRwtaoL3DSYqQ5bQCWWaMLyl70cb43KEHHD9SfGKmpKTM
1UYFGqA8vDi5cs7TvK76fEi27vj9F2KURKDDebw8BHE0DpXhafcc+mcQlqvxrN6Cv7W6zooRj6DI
dNeohPMHsGOHrMAIJ+rymi+FfFThAfvuE+EGuawU+aMCRUt++wpZ2DWNSxFnlA/KsrvmGvPW14yz
s//L6q7c1pzXyGdO2cj60p8RRCwAzJDLQWoL0vwshoYocNXizZcVm5euG3IKEZj1tvT5tlnLlgnJ
Z6VCggZclw0+WxN7B5MI7GeROFqazkRbhSvAlm/oPGJkjIEByN0KwsczIHAtIwLia2ft6Y5zVloz
lB7jTRh4nhHF1d6j15+eEt8OgxuayRRUn/nXkipl+rdcpNLIh+gKkjsn64tjhm8I2PtzxyrUhf3b
WyUCYdrXZxOyOFG5o2cA61yCt9hi1V38+W9Ml73pqymQO9WZcYvAEjaqqmF6U2fQrAdGsr1Qovu9
xSPFAqi8caMT/YaOlNR/HsO2ZH5vOZke0VhJeR30cQCVecx1rN2YhaGDXMv3y7Blx/VyQgMcg+Gx
M5BYzHufPgww/Ru7DHdrHI/vDXSdYIkfW34IoOXTooIMdVcek20f3IHiqLW/hZ/C2vGxtVtfTufI
0VKWGXl075d9Qjpll+4WYSt6EcJ5uqOPtDnhFUM/xYtbv5FG2f+6Zb6VfNJOJRgmDAdW3HGRqJrq
Y/MnyYFIlCh93qOBGcOIV2EnkX2ixuKRbCarZ5Y9cON2LaPTF1EI+PFuPjlytfUC5JznlFosGjVc
/J+I7kwntf41jFC+7Ou+OUBPsh70vdw5y9w/nApU67fGkQAFOPTdKXrESJ8df3mdXidOH27+ywYE
TO/O93emleRaEAQ5LsGFXRueJptNXcY2BkIEkbuGqc7ryBdFLdt61j+uDgu2vNqCqFe1BMQ4AJFF
iAV1k9/YAtqUyFb7TRb7mUwubLILwcDNRhaMDthGq5eLBk1N/0Sf997Ieqg4V7y9lzhYbqYWkxhS
m0m7i1b3Q463MzNAqSYcis0hO8rrKeq62hoR0GnyFESekGZUHSTPjJmszZBMV60OsEFNztxL08QR
h/Czq/o1qL1cZSDtK8qiWV6AXfkc1M6lXWFPfrxgtRJm+cfJbx2/39oLWHLc84Kt5VOieBm/xlWu
GPd/cJQs7eTuUpH51uw2XoDtjLa+dGMr0ZmVur3D4/cwossrghdApuK9wwI7Up5o+q59PU/v6HCB
gL3z+imXTHOFnRu9/h1sPkOJ5jvVcPFgzWJvo6tzautttCHJt8VS2tWSY3OmewgazTMyvdpENVwK
D/wtXqczHHz40UZ9sGs49LnSiVjtuooNydNTM9jO1rrobAvg9wOrCP6iPHfsFMzn+x0tJP+8cfeb
+A+bdjV2NkwL2QMKLcKsvEd3p8NwjwR3woFnqXboBRS8O+5uVtKfmSJrxUcSwhvZJbZhb/JyS32W
HzHobystEUyyZ35UD9z6AjM10oGery3Dja3R22wRqGWk+M6eDhdl/D4nNYyDBFbY9vM2Z7N9jZxW
Zcfj2KbKPRv9IHE2jkv8Dl/w2H8a+k/kD+Q+9f0byv+0bx/TjPFOLu6DxbApRki6G1pwUpYB0Odx
MMEYH7G3mJVK8eROYnVgYznLk3QJMAXSB55XxQdagwdEWDOU8if6etMAnE17pMQ7f20jtmL2tbFM
TfIR2dTEpA3gkV0bNRfak5xdA1BH/l61pT66OPmXZGt9U8rKRMUGdFLPSDjYI69UaUQgs8n8WZMN
S78JW+F6cvMNeYorZV2H8in/EhVMErKlABg0N2zVbL/THwVPVTPXgmYAvhKs6b6JT32+z83AAbQ/
ogtwhzt8CoRlTkBBMrl8DTfKkMp6g0Hwj4sQiYmp724jD7zWIzT350ePA/bQNkcC0cSeq/TuDJMQ
bjIMwiMuRgnMsDfcX9gxNQh6hPflmtkzcwsgUyje8/y6hELPHmv/pt4A/efDRva1e5NwTfho3GrV
Kkq7Gph/4zF4WgIsWdov0HHXXxZT41bzCSDAqFty+zHhqB8C0zCeakV34gw83OumAd77Mo/P3GxM
hv51GRqmnvi15QQZi3VeD5JPhY2vFotuz4sEjjzZpKYgwDYsDLE8RqTsIfmdlZVAZYBFECr8x9yG
Wpo6I+PzIQ7qyRZ5iQOSouO7rSHA/9OL4ycQDFfh/XMnhT7IE+pvYVdWU7/bhGLysWn8GhUgi+Xi
Ex5tm1Hw1EbJdnhWzhOqnqPa1GO4qrYmi2wGwuCILYN2EGMx2pvS2euHTgwp/tYYXREYYrzNompi
GiRraae+CkvnDfw54qgwnFq9Kmk3mE6j+NWuPnBHA08z6NDETXIq2eDK12Yu6LPNDFlwggVNGuQ/
67TEsmTevaBT4XLJxPZxPDME2SqmPEZ+91qhf5ddU9coMeMDU/Y54ximQPpX7ZuNhObHPC+246Uz
OWobebEIkafUVOKdsV+SbJ6Lw+sWI3iOoeDTeEJ4CK0N1DGHl8hUppIVYrcMoAu2aVo+LOG3t5V7
Efl3ab9o6ZROKpCGHNavQEc1Q3tXFkfcfw9ySnC9uSr0TwddLFeju5PaKvyD7KbmigP1u3zPFf8J
lEvIU9cUN3hcVmpscLKrmRz73YSQFpeUvF2I7K6sN95U6ouBrWpBO48G6yrMkPFuQ9Rc1sC4+VHf
gLuyUkpKavhX4L4bgZCr5QaKsizuyLTj7UFIUyX3qbdiwCuzKOENvtzCsw38dxY5/T8AUq4/aqI/
mAZv5xuW+5yQ8TFrJG6w87srHDZ6uDr/CrADysXNztmKX9pHtM1sDcVeO0P0130ELtcYkwC9/mpD
8jsj67BI5uswOhK151uq5jtUsbnbBJuBSibEwrKUtiEXAuW8VY5MQpdAf/AHFJ5zOInJhlNOksGq
8KLuwacc5HWLI88nfwdIzJkeIYdJmUttgzjW0VEk1PYUWipE4V0iyXJ1c20aW6a/9piyuvZ9jMjH
tzdNAXBY2RCxYzD8Uj0R9VaV9kLCRlAdRv1prGOOQSWzJHPnUQec+lXNsQ6nl2zcUb7UjQg3U2TE
uCO/UDspddoFBsg5Tkjc+ohrtdqLZX7WY15uUOvczsLUBu7oExrVHJ/DHS04lzwZM6F4yODiOLsu
mrWEh5hCkwEzQPaBJFDrltXU56V4sU2g5IFnG7XtkEgbH7bYW5WMbmhKFJJSHY2dscIBHavXKrpz
rbvaYut84EZoxJIjeZHJCoz4ynMt19v8HrFiADPivepi5DJ7VUVw5Il3Q7QPUcy9OtpiwuNiaDc2
hbkI20wbbGFw1eeY6h7u7OM4kauyEGApGNsq04DO4NAWXlVHGSWI4ykD3gbDvKE3Vo2M3Dy21IRD
gXdWdeoDnhCKO3Euaf00Vnzt5ky8UnaxXVBe+0MQHPdynNKMS7LsqSu9jNF+lxLGDhSoMh63X30H
sQUPzqzzvNqqdTEFC37Z+wgA+CFPerexNHQjUbulSOFZK6cqCIOLaxBvumg+8EHkcjEP9rOVPKv7
Rdxl5HxroEDd8zm4pI1egDTXkaUfYDVpVGA6httOC6wOJK2FxdmduoWiqvOgq75TVmBbprFBL5Yl
s2GGddboyFTIFL47R1c9iLYbSeiy9wCwnGO+a4BJhSwBbC9R0O7NvkPziuLnPrKJODmUawNsrOzL
+FLarJ7iBe7prshgyCJ4T8jF9zRdU8utMBEHyRM6rERxz6fGwUCyMPwb4jq4uxb54qA+wzHICkuA
TIsHkWe7jijPS+ezfMFLJIn7sOUMTo3w5UZVXYAQqdMpiHboRabz2vhOEXDB3pMu0a02GjE3C1Uw
zin9EhmJwscA2+9cK3OU4rgHrHv9GvAlQRs9wSm2aG2ElF7YcIDbJOhGSkuqE6FmGov+5DF1nnrg
caCr9xn4Yv6RS2ECzeKmvxJwHFsiJ/Epmz8ItrZ9c13IxhNlG7kVFA5kGWl1px13szjrfE1H6yKx
o1XFVNfJ3dHFqEL5Fw/LsXLdLEsI0KOqO2Tq2N9ynCG6MfHXWD/QTN3S4nDbB5CNJrRziWaC9njp
R5Gi/wH7vD2IapeRi4A4+FJ0GW8xT2ZG6dQQBerAFFoSn5dP65WYFwkSiMir4VfyMcFCIJDoHp+o
2LAkrEkDVWSsbCGWD68P2K6+IMeV2/zglmg/e/chn2LkmFBZjylgo+GGoDG8IecU3BBe1lsC73Ut
x2MG7XH745gjIGRbmqe7ooILp9PPueg3xBn4k87akF1c1y6X4mm50HZroPFlppiyv5mTYVvaZVUA
YwJWxPDD+FgYvmC4wtQI6zBFbHqONS5GWx0l3Ce5+4CzFg0+1AXqTsbUqZBvKG5W2j8zyFCOZpjb
oSce4EFzZeU2+n7/Lo8GDsfxxN8ap3LWqw3QnOox8S9q/JtRhkPt/V/JcnkXgLSFCaHA4H43zAjH
JZnoGk/kA3A1gHim0bNYLDJRYUCB33UuiWD9BYG3rbQtesutl8F8la6gT8mNfxxQaCUl3Za/gWLE
RUhqhDRBTPWCgHpvUc8bJ9MeCQn9G48Xoia23X/NqvTmcjkn4cNjZT144Vdh592QwJCwAtYQg/w6
xfGEesKA1M3h5UvTXBs1BAs5WNBw+N/kMAbjVq63VGCruDvjqiCPLikf7pPX+8d/YXggPJlXl4ut
8/45tuZsKNKGoJN4v5HWdZ9h5LnhHKgG/putzyPxwG9luPamg15cm9AsLrd/iMMqX5SB8gBFg3eI
zTlI0BqDFvbDmD5yGX/9HcRwfKRZjRMaFbwWJMIQ+LpE491BxMxwlwtc9SCvzz8dnnylQBxwUvZI
BbOuy/LYBunL7hz6AzyfRJihuiD0zM0bVi3/Ma+HV1AjLnOs51pzm9Fjx2YjrqhEnGE6TX7tlbQC
UBb3QuyBJrkUGh9YZyN2EHcbIwqwlWUe/7QvbqlzcuAjcGkGNeFA7GIbJ8h/9yzHK6ySa9Nucrml
Zxqaq0k3lsBeS9CvBpoJb0e1Uq4jL7ko6dxjV+4p+JJThfQ03hVoB0GTacm0fFK2TAP7NAI+fCSK
kWU9mjFa5Ir2U/s5eyvguSZCX2xDGFRpVmErH373ERsJpPma9cFDSfLPdJf9GjHz8+KY+58vi9J6
9RxH7D8tPEosnaRRylc9RMo3rqnzaSDxyXiY7S0c2dZOfg6VSmyQFOkN31X4wUtCiBh3iGQl4K9/
RWfduR71hN9jrT+fLg==
`protect end_protected
