-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BsanghYY/Uzw6kMCpvvaSYoIeC+HW3kHpIUyx5fZiCydFIMBdtbP2qoCjrn9923XRfOGfXXDyjig
F5rcYBTdZYdWvVWklTH7HA4sQ/AoXKQB5Hm8D0urbV18VkTwaaQFFhpGvZOxbvWszSRJ4wlGixPk
vAJ3w+TiFegZ2zqo4najcPvV4eXL/Y5mXZO740i151gTJPSc+vOLzb0O6SOHqjUgINh9xO+CFkrL
6mS3O0sPD5nkZxDGP4sPYenkq8o/xxpsjg6vr8g8LAJmvyHtKp47LCow+qmh9V32gsIcNyfIgqLj
+UhNpFX47hbW8jEXBxItDZwynBsQoXGCeHHffg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
cgDL7vmonTxlIkIdRJp6F+QXHVwRnmjelkFSuKaAAc58QOBsNS07132gZTE2FshTw0aRv+NCah/4
XUyiZyvh0E5NXytasG3ureyzI+qZKreHbxqmd6sj3vx/O272QKGEsU0xEJME/SyXOW74ctNkZfO4
YgLs5u5SJYLGqedMa9P2TRij326yrbh8PP12NZ3dgXWESwG06Q8ri5TklPBxhYSpQ1xtadXjGEw2
wGZ1hrgo9J9ObRnDgD6YWSk+uTgtWRcebJKxmF5n2BPIoUsT+EV8hCouz5F8dtrxxFtZK4DT+Z9r
tSnd78WO/9Uqcl5uUwq/TXRaYEqdHgpd7sLnftUwAb1EawxxpHN5AFBa4Dv5n9voHIVxeQTfs+Xc
X2g+P/utTviDk9lhspxbFaNsxIbbydjaoZmTvg/9W9hXtjCBgLkz42efI89p20yG0LDpsGbLGJQw
U8wgjDqmzGdecalgLbc4XGEx53MX2gF8/FIXvNYbSL+b4vDFfhIX5iFpYJpzHq6VedwZfBed6r1W
G3A+TzbUL4WQBFt7Z596VRt00XBbvju9r8Cp3wyhOyA8z5GWDcP3nw57mR6MYPSXx35ZCekVT4BM
U+vcovE4T2ph79DV1TRU4DIJ88rjlOvVCZQTsYDlkxiFhF1WZOkkVHqsL2dL7Sy8aPx5R6DcO1dm
5d+8c0D2sX17L71qXEW6V+8YhFDqS0FWxShOBL3p+REdtc4Y9zlsOsmK81cCBPnhf0m4wJm2n4v6
sX7EBcG5T9XGF1tkYvvU6QWQt/w1E2Qe1qNOQlHFQi9YFuIamrbkzvzSdcs2ttiRP9EjoPgcq9L1
GXj4gIk4AkCFczUGLwLt2dki7I/eb4ncWuRGPUiMCuyu+BavY0KGUmTq8nmPUwNDJ070bfMXuuXk
sfi6XtLMIxXxmDb2XCC29tKI5LPxXPzAVB0/XqIKUCbiljVo5/tYDKKLOc2RXv/I2tK4OwDPT/N0
OXa2rBGQ3CWbjjbrCCA4NwnCrHRxV6nx8bhq4+DrrH6/Ei6S8xky+IrsLFvpdz9d5IficsyvofBd
/+xg15q0tm+e9nBQo+PVuBfBhP3+nQITSM/1HW8t08jBFO0Plll5CnYodiED6LMUbjjdbEW9dxGY
awtwnQj2YQIG40rljo+WzV6Sb2lia0lHvN1QEikbj0BKtg40zlZSJVsdYsJULlY0+KWYhJD6iYHj
+QllGmM0VXjBzjYjoE7ARnkZ312QVMBaQ6zL/gk9+GJTE24bhWywaf2Qy8LS6YND+rKPrAO7rFVc
MBFiPIbvXJzUhkp8gg06A/iQ2U0sRhMqj3HrXSgTttMh6mZS/FkOpRtG5ahm0DcV5lVucb/mPPAq
3jeCe7THJjuop+vg6l//CevitwiQDy+YFhm6eeaBW7/YUt7WLUi6fi2/Ljd7jnH2ZHS20tc99HQ0
hHNlMM4WbsaD4Xw3dHF2DELxqujEOhdMvP9Gr9XhPgb3hI6VOFL0IZKfEL6XCdwkWmVXLIdQacEz
c4Um4UfxVoe3bAEIL6g/DwB8wAXI0PS1BJYcItluWS9lU1dhLCDA1xN9Kos2zLCm5EyvNyftcIXG
nwdRETmDaGIusXW7j6BxwpTrsFDzMBjm28pvwGcKkvtfnQlqCtGW+4a2ldg4KTNYMHDHPeOaHzHn
RlRpLjRNNZtq34xxRYE2wWW3E2CeUq7Q4TuEzJ/tBPx5lUHHPVHvW2pXZ1abFjympukhy4ARc2yY
su/lAnBFdEJZkm48ElfcHiqg7bar7y0RrKxVhzPlIR48GYDYCBeH6NXIDOpq0RfP8Jg6AoYuVU7l
+uM3Ih5TENm/NoO7mnXPa0HfbjYWz6D9nyf7OHw37hrEkRQuLvTpqmmQVE9PY5mIMddadyrMay5u
ZsgKewlcJhlm+/AgdxbE8cwQ3mvNOQD3uBwdz8n4h5O+e8bWKksmCWDqdbOnSrKnHfWb9137hKzt
0jSeaLk8Jt8xzA0SAOEQegyWYnCYV/+fELFdw0fppfCpkxqtYlyV77kKoSOwnI+d+2ADTcsDvxHp
bqIAe1SM2FXGLmOZH/+1JJ79x8sCJsdHHT2uD7dNhqhGahqhwHU5DFZRJBG/iDcPZpoMNw5ijG97
L4jD2dKbm+qtroNemconR+Ez8Fo1419tRnztD4VY6UTT/iGv428u/9hLU2mtAxnDzjcldO72HHzY
92CL9mye7pBNSwIoX7G1wJ3LpQnilNUO2pvLRPg2ZTF7b7WacAsGbVKxbNekJaMerJsgSrqCWGhP
bdHeF4aoo2RUQiuTJQqHxS5vdGjK8wOsHn0LehjDpdlbVvdboEoNZjBdoc82gX1U90Lt/ePUMfFJ
kMDY1fJja3vneWiC4MYdDS+L13zSkiWmH1NqkTINTBkQgEjwlzVF3/TZ8SbbwLbdlKSoYHcTj+EH
cmjJzWPMcCF/sMwIhxpyfMnu0FE0GPhGB/ahtY/wjX1eJdXzx4GkELmBXtPJ933F5AKgjqDtl30T
37q8nJ9pnUQRGCfs1hel8BVZCDQ6aNLAkJBuA0uBFDix7zDJRzbAu1m2Phw3328S7VZi/Nr3U34T
PMuKNQ0Cj3KfxHR/UZsNKYPaH4vPAbRVfwtYBp/3Cjbg0Wd7O2Ftl0kQ5QzNxr8kWfycg4MMwqwM
YgpXIipskW+xo66u6jwgWXPjRG0S21n7e5afCiaeG76Dp1KZZp3K6JnP85ZFvomPMxegSsGiu9s9
zivDNjG/qKeeH5PXZNii2HeF1bt0nC28DWn55Z+IHOxy43u6/ntXuCfK8JyDhuoES+5s52V7q9Y5
/uGVCJillqlmCzqJXMWDsCVvO81i9r+nlB2Z9R5TfhtAeNX4CfnQTs+eT8IxktPANy67nslkaWWC
F2tP9mACgqYhZVl9Wg9DHFoj0XlHDc5nZyfUZj3vk9WEbuLVOBPPaRFgz4dApxoEXANQeeTPaEjn
PvTmREFTDk0K4QxamYpVeOmHKvUMoFLfKcEsbemz8QCnu+jnINZnY+Roml3WcjcLbGahnEdnOJ/x
EijfD9cVSedfZWZpjLeuRKk/L3XuuGXtINx4qYp5MGgVzTlZ+f3oY5rv5XsUHAX5FmQF2+fBdyuU
/SYeayaqTmX5d5y084Xu4DE93+CI97pHyM0Tsg0RKtERCj/jOrcTHzUa3jmHsCC6RDY7YwKFqqxo
2kOyxhhiPlx+KOmPqXiFTCUqHf33WskaGl64bi2zenQOn4jdh4kn9QMrwFyJGifKQOLDv2iYjLLm
ii55XAK0kUB125fxjBPbkiPibtW5szNkmWq8roPbwK4uStcdpfcgftCe5/vniuYCOW/NFKy8fs8M
AvG+4JsxDwJtuyp/LdDl7aMwccLgZpPIkCrS1OvIYCDWxYKKQTYSYiO155PnuDbXrIq0yUG2sSsc
wMVa+9LAadZmqmIoCl+zGe/Qid7JHMXeO+2jwRgqM3NKrlZkpWXzb0cMEZpkWMauag5ddGg7C62L
ZLC3uEYDV6ElyPuxnu6JYW7B4iFThYs1iaVSjERrkR/V8995f7UOI6f8Mqr469Dyrl6sJnAgC6PQ
FwKK7FhFVqXzhclja8oPyl2th20HWm0Iq/QWbAJCVlOJkCVqlnRFJaBjP5uPAGmjpXwpnjFJZKws
294UXFN/QGmL2ro0kDTkbrvfIi0cXTTXHiMN+WgL7TqNSg2Zb//pt0c2XDG1QhfZs3pUbqC0gxJ+
JmO329mkU0SBd8vlcRFXCj4i5k+jU30Ckslo9C0+kJ/L75pou18jkExQSkeqCV15sQ+pyCjBAs3r
cYzUXXAAQR3FMF3IIrpN71T/W6StMh4LNC4mVVaoFianAdMre8SWVlkBp3uLViUd+PFcbRc7y1Va
qngDCTSb9nIu/CQaQloDHb1AWzJ5FFXi+eYWtBoKzmfrk5vPvRs83aknA/GX1Pzwa589WKXz+gvN
93wP2G/2Mu9Vx40kLYaS4vxoFrTCmRJHxy6Vue7bQgm28lNdmc9CQavrmilwkBdv7P3JAOBe/7DM
D7Bjm69CzTcqMM3KsVL9iCCs0qpQQ6+r4/+Vmw7tU5OHub29ABKWCG7xMhX/6sPQNvGVod2n84z7
DR5hoPo0PsNi5CGXPv5ARflDVb3pk3zXt0rs2jTwyxHMnoEfnTaSSSbRZIG3irQ4jAdTDDjr2na/
3COIT/eXNnB1Pc9DH8lnEJP/Ux1BDsA6uLJPkWPdQVD8MZmByo9Cjp932dBFQCzPbalu3CwWyc5o
SV4bljxFO0pKyPzLGglYcy0zR3CQtp75PkX33jy1wq8T/9LKORlptU4rN9Nx1T1YCGBQHjrBbHar
4I1+tx4fTdEegsdpvBbk2mLrzqlXJdSrMV0QVFJKE56YlRIJiLVxNWVPCxx++I+9z1MExem2h565
USC9ja7hKH0KMXj8wtVHNzFiEcvxQcmVOhjC8tA17+zdPFx4zCnDTufGpcuJy1SC0Scp2q05iXfN
sExJRyL8HgjWpJy3zg85J+R7bw3aNPayAvT7OpD24gp24K3XWudexHcdcCfhWFU4c0MOgQrw4UVm
eJYD/tHVfyLzG/zsP9pSP/XVjm4vIdNcnm3D7//OI3HCEGQjGQUrgB+x0mP0qDJTERhiJ0yhqqU5
3TmCI6rxA4GeRRk4VL+FOwG6LVAr+d/nlrxd9qmUeUhjtiQmhCh7gMzsjuRVkvKvpDFBwJ9TjQRN
+8JqdFGr+94qrj4ezNAx+1k/JuPuYzbqVrbNrmOmTydsbb6UZxfAa84KoYEBa6KnshGfPjpMWdfH
7kw08Ro7NOv9NZsz6cuqWagj4ja5olCN/9xlJdFkj2fdHFhkKlpK48VQR86K/e5lfnZDW40prcyj
mtuaqiQ/E0vkirTfnqqUPRUD37u/tKn+Hn2miNH0Mu7kAd0fS38GomghVieCD+wPWn+droL+aS3z
V7wbu3AP/1FZ/vFG0PRlkCq4huihfjkjnjxLkc79x/UJpisWSKYqD1Kf+JqkqwIl0nD/W6JO6xUH
GmPygxrEPA/jMVPH5tOZp81od92c0x/1UxnzTywtKGf3GkfLWslArQOeFDS2qftlqPyhpGCuK0j/
scbwH1xY3Aqy3E0gzG75TFdxDV4baL+Em9ypFbG5+rIEG3mqqTq6ADhMmJQgtB606MWsgpOCPrS0
eBp1/aYICGVokxLhSp+Xf7n4j5lU0RkAb5fDjmDKHkDzOQ9l7ihUZXx7l6NHLAATIAhDErOhHiFk
1/+HFKeshhMicM/iH58c6ZRlgQze9FVDN7AoG1WL+04skRuywTynQNHN++Ceq/ZsN4C1+wMfFlBg
YBp4zNotiHn7QZG3KuV381Qhfy1tlYV/MqLwvIaYSxIHaxxVKoQXlk9MJuS5K4A2e9lCH7wTuLla
qaa+sOv212gEYDpxfxC31ei/sZMYp2lUAgf+5LTtbjDO3DFpFeTNJFMeYVV1O6aDKwA5iYXTC0mL
Pfljgx2EEJVD9lp5Cqn2PgfF4DzluA34tgAXgQSp99gp8TPNku8qkit7zmm1rRx2MF80u6Q09l5P
t0vhsNGUcnaAdtQ7iL1X9ZGEPFKShJynHJvG2rib7/5wefTupHlUDEHIpPentI8lN8RY9EEslBH/
/eJX6LKE5mc65iGVyjUVRLaNTLGsjngV/F9taNtEK4xj7f0sQ9zjaKoaUXiLUGdFe5SAHzUmKtHg
r3S77zson9dNAqmEF6AZBoR1NUhsm1LrTc0m4pgeiI95EtpdKZHnqB9IxYcB5uhjYmykfE0ziN3A
X4PRrGsRKOBlisHmDamvBoMrm+I1RWeR0GsbrXppfVDKvQB8sp9XEJjpv1Ge6JmaFSyuW1xKJ3E5
mVgZYy18gu9hxyNHvEGmr2yPKPVhoquQUhB+ztqT/r+O6mrMF07wYMqv7KZTyOwe1cHEKiSaU1xc
nC0wh2lcsSgmnvyj/2OUrGwgcJ2Lwuex1v4VBQoIiBoqB7E1Rcffw5ZNotYLzc7JWgn+c9vL/zC0
Jz8Vy8K3Y+EDcc4qIkt0H5wcgvDhnPqeFN64UbGzyMc1SRwJK4e3ZWzgUSCPFB+kv6PBGb0+qiBy
gerIN5rrJ89AlbdGLbU3Y1ImzxTaEjITaUcIABEifpm3g2SJZq9olmME0CZRk8b+cKOz61to+DFG
D/X/yGqXzcfsqcaPMJ3ANmx0lT8/HziQsC7FyvPbEcUzi41q0WLno22I31lLh7amgEj6exTyq3Gg
7CGi7TnYRQVRVN9gyZQSB6YD4OuIdb4p1BhPCRX9jNOFGVR4fVMlN4ncmuVw6lVPmELUe5FZt2Xl
Wkh5P/YFY6CEgn59/2n5Wll1qgBwyfC2PlWkTQORoW5ejmIAos3vLpTsR9Ub3vgjDciIWWciwJVk
Tox+J2cCvUjK3H5x05pXBL3YpWwdyCMsVNhRUk2UtxHeBFAOmIfGv8TcJWK7nblty9RXuTodPL93
w2MyG1ycWeb36t4e5/LvlE1tk4v4GKP7/QeS27Rwt0s/DiZg3ULY0r1xyK8kN7UHYAM1EzBqDgKd
IbRiGpFapeVXHxe3qIM7/JdqdXXsNCpAh5GOQDkW2wY8ZCsgwpf3dy6MnqO+uIDOa6bFx/7q5VOD
ztmrTYFng8317tLr1BpNVZsuZwRuYClRZApq7TMQAObykAO5y+qwzulWLzU0jC3Bau6Ik/OHULdX
6M37sKISivXTYW2ulLLxjvBc9vnbkWvi29L5tdUDQHjnh9lctGR4i+cDR+7lbm8bqEKfKVlYyhy+
oRj3ZHy9AmwZSKgLOoRQ0g80VazOPQdOrBp59uWL8VWMSBkS7to0DwU2IS6b1otKmpZMP8HqKCtS
e6/kCUbRRFM5W/RrsZRYGQ5+i5b/nNsoFf/bJ2VrG3XzzWSkJlZX4rzbOpcEWCu7S+SD2WG4gOOV
mBw7er3MuZ8zUtMZJLnh7Fy/vnCk8+M/g6c7AgcD06ORo0ekg74hu342xyQr3sQq8DihtoUWOV2o
BPJey0bPFKv7nklyYSyzbrJ5dd7LuQmRzLbAvl9kTotL/jydmP3GTFMof/az0RR5WTyBB+FjSOsu
oZklcpL7EWOU6lXWM2F3H9kzNv7cxUQZ2HGSe5ei8O2t2q3CiNI5PzXgtBF3OWQaYFpsgrnmJXMZ
F31Ids6wN++zk9CqfUD5TuAUfHG2KAHub214ivzSgD3Wg1T6Uzg4o3nduT+CjBtDc0oUIKTtjhgb
UvP5sgBxUw6tnB90M/A42OaAiOeXWBFIIKV6h+Zb+4KvrGVrHQhMDALrzwxFXdHaDH5Mk8BRj4B/
YaagxUASk+nraSNIApipBdg9cfSDB8wI/VBnVKy+1l5/D5kLxbXR0oMK/nqPw02xNyOw4YPgb2gP
ti+mEx3Lw8bqZBKN/3Qe5dSLqyI3Asu0eEj54RMLT4bVTHaYCyEsW3mBnZxg30H7C6W8uoE5QVR4
NvW8A7RaRWqwQQknbh43x53N6Gij4bxC2MWDf6BRqnR964w40AXLSsghn41B0i145UForZP7KYmL
Ep0tf/SGcxdecqf23ARcJlhQ7UManpr5/KOa4wzK8QpEXJlZZ975DnQSbjtRu93dhldv4uJJfG71
WqtLSIIwGC0tN7D8AE/iqV8eabKJW+AjAuQfU1Qj6X2xR5GPX7kRnVLdHtbL0D6xGifwk8Z2oWdl
LRPc+SzGXdP9ImD9dkHf1C8XbaDrEN0gUDqKSlE3lmVcj2rdPWKHfKpUZxQL5VbyP9ntxxOWn0Jl
2RGOiap3ab21FnEYo23gOME5u05KcywzqJCQ1qUPPEB1upFnx00MRWGXX6C8bjliCGpZ2qNlm7Lp
rswcRPyoF17XKHqxedLOV9J30oTsJep1qrrpijt/JqtA1n3il5ybXC0a472WMF1ME4edWqRzhosu
pPClrvZoWKnKLqkGsDeHkUo/XdCmrkwyXq0ELJ0eAFC/GD+gy+3qUSXiV/btkTA9A5RXTE1Jfe0Z
FgNxko+8VddqDAyDMb1a4Nu6/Uyxmr76RrcRNTQLUSRCVD6/AjsjHwObJAH2S0IHJ56aw36PdQ0v
bwsnJGZxxsSuY52lL0jmbRz2im2EAsNopKa88in99eTxc2syeYzStIVRRaw15oQ3o4NYFq4sSsNf
DFjpmFCBDBKRmJ9YrT2yQFpqz+55TvKYEHzyOZvnsDa7+UDnC5lTDRsSaurrN8z/eWeEVq++X7+F
QFQcyNbge1Gr0sK7tQ/M42q6jzme+jbtQ3W284XtWQhmzzlsXYMSluRdqyImqg+UNeDrJqhwYr9D
Ypes7+GKkKGZFBKy7ljA6zdWuw8XXa2vVvZANV0crF23EL/JgWCoVNVtJd0XAs1sZdS1I+bnAmmM
qh/xLqWvjmsMJEhcNEtsBrg7U7AlyfQeIp8Xi065A1CAKG9mxd1ormOY5jdhI5krF/AlgiJlNnP7
LB3erLAPseo59vygyFHOiA+8jpyAObqiNpojpj3aS19BR5KBohr4oRJQtNCteKId6PkqNNsLBNsi
XvaQvKjpnMQxGnx/LkdUZGwQgcNBZ7P0/km9OSxKargyGe1yxJ7a1zi9YPIX/mvHOfDCCiNMSlGm
gLVTgtC0kT9bMLhCVBxpJ6nQcGSV7UUPcBWeMR+Qm31rgeeJSYPnywJR5jNW7YGeYyegCMds2GIJ
PhBRmrmiYvjBnewbezDnoRqgwM6uDv/GHAvJgagRBV2k6ctS6OtNkc1hym+FBum+x+fNifvs8JQG
NjKL8oo3Ld/NMR7CNRZJv0PXt5VvOshMxAV9z+gP2hLHcGHVJmXFIWHiL3fVqrK+I4pvsmpR7NoH
5yNbDlcoGoQAIdCjSLGw803V65lhs6+NxCaRFtkrppMmuW/EpTOz7V3suR+Xd2MaSR4xMa72VcM9
VU1SYmZrBsL/96f3nUZuZAs2q4IVrIFnDNmYRfDl4Be0lfuGDR9Pzn01zHYaQ9jgeUkeil0w/Qet
7AB+AE1X4ZIgjVIB3N5sFvtv6LopTS8Jz2kLGxvsxCRu9Rwv4Wxv+hdKzXcNWYUcWNRw3UIeco3y
s7RNo0oql9oQoWBBWPPu9J2XSX5DPb2UvsSz8QSBamjw/2VZnpIIC3aBAtIo7hoJnRKOhxu59TMm
N6hhyBLeHDuisQMquyaR7sYW8TxTAT2LYru0rj4oRve895z0fIJiBOCwryfuoZSvDVTv+wM8qDwe
nPPVTWL2P/776ReIuJn4JyZsIOzoIAijrwDnV0JzUCrfri7sg8pRVPAAjKOD7u5/7Jh70KeXeLIr
ob5ppvwMGdcuw7KuwLd3eYbD4Haxz0R1UMEuVhLZ4n+dpmfU9kQ3xrfDQT0g6HjvWX3E+tMreOel
tdNWl7aNPL5fHMLy5EEgOvL53IzDe1KUbiuZynS1x8Orgy/p0CgHTjFFBqFI6R9jMErzSXLeQ4Lm
5dRb/YhSpQ3ULux35tC7rr0TIJHd4dN7n0hGpqkC5VblvqyCxJXHYKvRCwCjeqkhakiaLS0554mN
Lj7WldeC9xi4OJ7xPtLfoD96TcNmXacnXXs6ZZKZJ5kyRY0Ee9k8oGuIuYECGoyxVEyx/PRi8ogv
EJKJ+R3DA1O8uDho74FU0JGszed2oZ0U3+1F4Vp1ZNhDM81VI4yk6q1KpLx1YWqj4l8YOtnljfGC
elm6A3j6YCCNyDE+JBwCQf7x/gyGngjxyjkWhtI1Bap9eQThg84E3sqMLqmy+XhtOD3X68drIHVu
tm6Vri/q8ZMqYCXeZjQncD2kjsGpvwj3JwJlM5kTo180KiGO2OTJUqs0sen05DQ/K4/H6gWjme4m
gWg8N7t/9uDsUWh166FYw5QkOQHC0bQOxSHHqjJxXr4PjVXKXoqlsDXimqwUmBcw944LIPnlQ0uN
sZhF3xD50PlkcYdt+D5ZNb9MfSbxQ5QwL2O9H986VRl809lymNR9uGrC/cqOhAzusX+ZHRlCxwmg
7e9r5Ma4oL3WVNBy5/OpIMDwS2wCttjLn/fgB+EzamqRQVTZq2mB+byG3craQlrpXV1C7zWXxPbV
X9pdH+8An4RBAL2LLjTs9ppVcQM572ZlGqJ3QJgMbNutMEShjGyrF5yRcKi1pDVDa8Kk/HrYCnVv
rSWAlrBgRqvjuUj/AAJF5UasLEfhwT/0Afjw7dju79uw4emdhZvpsUyw9SjgIXdU2oeAdZCK1XDY
kpa9CyASAJgPwW3LyaVWt+h2OSG4hZkHCTTSZ4vlPIOIXLMcVJIhNC6Bja2DDxMboT+DXU4FNhzJ
8zw1ue3OtjflffUeXwmwUlA8YYc3n8T8MHlJ5celGEJVtKUNYH3tBF1kdmYAQtt1Hcaw3Ut1qD6K
eT+RBcZusgyEtMZDsbplSNRshzT13NGOcC3Oh6PXcqDEuzuSSwcfp3vaE/VB6s7hxTrQ1hbYHXpJ
9JNmxy016K7d0BgHfr1+UIoN03SWsunbIUTw8cYsAjEluj7xFnMvmSs2BSwH0/SpgcFNUpA0/4B1
gAxXpE14MA40UYeHAFDZdZv+3G3P75WrjLsFoTGXGPtn+lWvnGlnYJm826VhBuvZeNX/z2TQE+sh
jnThFyoNbb3m9oMPXQ6CqeR/4S9pfoJzKOO2aonUCf01oWb/+fdcPNP2sw+1blmdo7/udKNcNxPB
vyxAHW1NUtxzmFiBAW3eaalivG7/vh9J/2MfVuCPWZkpDPrVmAmHzZ/Iqrtx/lP9MweP6q9DdV6g
/kdcEYpnUN3RQmLFh3hiW2uUiEsjc+9TaJW4l3kGQnEPMaKTfaYcD11oTtvyZPQR8SRGj9nKL+eJ
0KEVvAGiceUu5+ktOMviBBBP1EF73WPN/OM/ta8PqsM3aB9bqgAWBkffyq15s66Sht+hbi7kynRz
rYxiolHzJyE48WJyawYBoDOmWmVKyugjiFS1500CUBJtS4ER0rxyl+LreoD+/jalTK4NCciM4jJl
19+Hesku1rtV91nGpg2qxIxi2Empc0ZlDjdrJVmeCtFLYOHNtgLKbrcYB2doyOlvQH6oDrbhWBpS
mSKrDkM25bAYvkivWucd+N1ExYDV6mOLyTKqATWdatCsmoJJSilGC2+lq11Iay0L6EKlP8FJFjyw
L3MjiWoQbmKpGm5ncp3hxO6BuVo0KUYv/n3ziuShnT/8Ji0E+Tq3EeruOYzp9Q8iavI1qGxJNvop
26KQmF/UEuxKaQnFHbFoYmAqla32erKH617MCQhQ6EB2E+XlKTVfWoNNYJvlzGf58S1tW1pbE2Om
4gLmk4R4xnr1w4n22oW4ptroieycqJWr99k2qQe82MCL9EmaGF9swfKuz0rCSfNI4+WylvEMwP5X
EUEEnJ+DFvUljcAiOdRGz02ckrphjQNm0kOo+q4d0Cm+j3VQtvZPziKaWp6Vh9iMF9m4
`protect end_protected
