-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ptHFO+z1yIr4/kRUwQctj3vaU99YSDKhsYT0AEeEWb+v2rVKbhmCIbHPqxDtUjvQi2NTheb3+Mt1
p9yY9x/uZLf2niqXZfQshI8t7nWdc089PsHNglau4YWSY7CRxCKdAVMdwIixP6R1+t6W5k47I6S0
nJhL+ghAKgGhD4SAvcHcLkydcnBIZDkggZaKisysdsOTamIyzMZ+ZmhofVgNucUOBNh4RXte+0nn
0zlLZLWo3jBkHWXgc2F4Fgd7AvrMP6noyCV5eXyvgE+xyj85OMs35fZaPg2YuJgRatssGD1tVaSL
dwoVgHkTmO714H+9XGNhPVIMDcTj3wb4JzSQHg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
XHssrrDworGLLUYA7FuPP2Da34/6uWFON0URrBnpIXjKVWw6vg82J6Zd4/0+HoYyIGfqc4EFCtKY
PkKK8SM+bIUAwku8rVy9ZHmJmKXjC2ZjaeD6IoSV+Aify/EZ3Rf8F4OW6jj/WYirJqkhRJ70Eam2
4GBwpCnNgY1zkpf3NEAQ4Q4bguHxUHGbYQC5CG+Ws9Za+/h0Tx7GOhvBG5wqq8U+1ieJv5xrt5NI
6dZeEU0o6Its+gmm7Yg2MKgZDti0PRWx/rssezsRTLzW+ntiqGkePeKWbGC1YqhqivVc9P7mGZP1
/v6YBNJJpN46A1uOGOW6AgelbAwYFTi1sRIxiyNilpSndc0nSIITnTB0dmpysFRIaXwYkYP6F0ta
+DImXgRzsrVV30jG0UOAbsDIdPRSHxKNg1CPoJCVmWrz+a6MGv8Les4IbfxsOBngkgij/fDB1drq
d0EpLtS2Bjr24JNpDNVWZr3MKotPwOdE6GkOVPTJa4NymMl+ruoloOTO6ZW0Qbt/wWtnkO/MD9hh
0MeEkYMtY9CQlXBTjC98qyb0t5sUL+l6s4jiWcEA7BxPwFm0KUiKL85AnIu8hjjH+nTUxl9yZ8VA
7yi/1cCIGHewD/RWb+dJfY0xttGGojtkrHbLKsdK19FUn9J+mpseX+Y+7r6bIG3j3AshCt3yAX4g
zsgqoCJLYRzW/3R3DfK5ozS17Ua8zpwsMvoraDi4/rtiooR10odoahzI/YnzXtdkci1PEBrFkA8r
rqDbs1BdzvaJPIlOMb9yzRtZrrXfGlmmUn/BjCOLeVKGE6HyVSdLzg9hzpUuXYXLeSIcvF0TSh05
BB5LztUQq6tL14kahvgD4fZBZ4FJCLtLlXu99fmF6hxL9IXmmBpdpvmz1uesS+hZ4FCsEkb/APp0
9Jzf4HRM9p248tPGI9J9Q0dbuf1JbjiMYjpTMjaF2SD3PLAtmEiliS8fCZGynGHyIulFEu1OH04r
Y4NwCOvdN36V6widKdNbh0TLreQZ47dr6cYMoF777eWw+hZq05USsHX3i+jxW9waZ0mAE4eX/bwS
Mt7IOZKN0f9SJJIjJnQRge3wbQUw+lbsWY/X0gMry8PqNqMci484LouKao+jsP1VzjoopfMxJumG
uSBMJr2BrYHIJd3bo+qZMeqZD/H8QJsx7bpoVWoEkapLoxR/FG6mTtyXo7zcAVZtdXIYufwvoaCV
h7InqHv2xxsuy8BHu7rHor6kKeMZzL0ELvjwfV1PAeg/UJ54eia/5p7AYo64fq4xcoOyn2m8Mu1W
QjpbW/YI9PadzSyqfqa5SuQyelsl/PCQbmIzfxyl9quC8YmvNw8+eoOc5pcycCxq6Srmd72GAINa
t/FyWZ6KH8kDmYjT0G0WvjnEfEERw/WBOwH3M6yUhJpOIpxj/VUxU0CwQ4Z3G8A4J48Bv18apmek
+PsW2p0KwnolRiOpSsbCcfNfZT8Pudc7+r8WQg7vLuPo/vLU0b6K7r6x3yW3tfBpcqe3NmY5mEhL
o4dPNKA2hcRxIwIyPDAci5X4s0ddjwoO5iqYN+ezJojiMzYwmV1pgeG+F4PFoPFNoU+YM0vWBalk
RnmMVJOAsXnsjT5UBIoBRSCiTiHdWEiw3u/VN7d7L8i0JPIzOlYaa8p00lVwDVtIaZZw+P9MCp3I
6AQuOHFvfO4WAn2waNnySmy0WoHaKnoF/kBxQnfd3wrHZI+1XcGXxy4q2eWHAOPRpkmwmhpfyBX3
w5iCNqZfYJfvgTCaCl244KsgJI8FT+Uw4x9lGsf5ynEHBhQSs2hXkNFZdMtk/TkPLSV5H9PJBSCA
fkY1aMtyE/ViiI61I/yMN9SoITtrBm2ckUvmwlEM8vPMqUXOptiQANTuMakxuY2gK3xlvYRl1q2G
+ln0DpPfgfhaLlYzvuZMERSXMNYRLcoGG8v4aj8ql3x5hdw+INh4s0ER0gK84ZLFyB93KDfUE7iX
4E85raYttO5bdmgJoso0Dxlylan2qmCFQjn/87ygRKBCmGpbVGC+o31utnlkmEYEgPzHSslwnc/X
RFPOAfpJuvEzp+U9W6eynApeyVI4qemNbyljnGmvEthmlZbCZnk9doyIT9U1r1Y9XdgF7/ZR6V5/
sPesxgOlETvEkXCEW6pz2aYg47Dt/xW5iy94S2jMh1o8epPCs6w2T8KA7XdHlx0HHWnnuO+dsGug
sGwj05nrjVahYFyQw6honoQe8/rNEM9efRFT4XsxTYaujNpbaNE3JPrOYzQuSXbXtJQtm19h+cFi
kc8OZC+0a5G3qmISMkpV19vrRYnPpGWM20qYlb5Rx+ZmqAlMNQYvtPLidoZGr0wVvO4INOKQ/bhq
hluwU0RjWq5rPRRzNInaQ/Xgh8S3nW2BrOObFbAGC/hzANJvuNzxy8yCTIB8imqLvdEstVN18dHE
IrJK+xsdIRzacXhWg84721LWXhEd7/CRlqF9GCjzCyNn3a7lwvSBRzHAzOyWuk79koKU67jNWiVi
aRu6jYujwK3zpkj58S0Db3QE4f3TlN1Bio6eGUB08An9MHuRSH3OhjdVeXQh0u8hA4d0VCMUoNS3
hu7MjhxcmM38JT7NqKRFYpNjk8N8EoRwFxX6W5wb1jh3FxAhm4fz0Mo8cm/kz5zsPMd5ClN/Gh2j
iwZ2IXWmxUCb25cr5cQXVrWv/UcnNKUnEtm6/1wwdGmW1TUnSqkjaHBIJ0wd6U1u3wUsCsRMyx8M
xaTm+rS8PJrTPR31mGa3pW+lpYPmbx72iOS6fajiWVYrMkPnhTT1jiMSTbW9GxXbqy5dbiFQfbje
F8JD3xsLWR9dogsgNKOvcBRgokXwAjgr3VqpvRzXDeP3iEtI8oKWCZn6OvvWCwdDe3jeWsMSLksC
vptL5ivg7aqZ1AqUO6SZO0/3+VR75/tcTnWvOnPyQQbCqAB+m7DJ/2WulsxAzkXArUsk+keh+6ku
BTOgNDJUS6bp3En3mZIo0n2WA32kO6icMQtdqv+lTF46Gw6HDj7u5kXeohLXWDy/LtcWYJ2V5anT
ov+VO1kQd2tRatSwtLjVyzUzV5Oi2i8QQZ7kJHB9Z8u7PxyAmpsE+RFPVxgJnvq3xnohw/0Z8UNU
W1ir58/DULVNk2oEgZW9kGy11cfQ8qO55vK04AikvbCBiiQKjvcJvxQ9tRnmVt7dJixWqKoKHZuq
AWTShk9yikphV0fZGh+kCpnEL6KXj7rmC46REHQehPFoqGFDHS5i+FdnzqQ31AIvBNQxonQHaa7j
mqW2BDHWUcrro9pt97JPvpsddQP8dsftF8mNbw5czdNdPOAaPqvKEVJP1yOyE9PlQci0/vAslxas
eq0R0+1bsP+4oH0wrLobDCV+XObSXsoudlYoa8LKb8dy4bceHzACF4IWKFgiQJvnG2Tf18FI8ZWg
9uUgih3ArNNm2/Ji/+JiwNIt40EAzh6L/2QgFRepf//TlRVo3iYWamaaJGpAHaryMn9H+qSNLuu+
Hc9mH6Qigd53M3HiyIMZS5fJszkAeFcFrEALNcq4xkDf7YZcVlyYNw/vvr9ZmqzZwJhcN5U7bK/3
Vpc8I2LHEk16PoWVqRfcyiGmQSkQZHtEgQ6LDkH+lN8G23y1cDsk6tv/aIZZN0lu1kchWqPaeF9y
m1AMI8wESSTIvTXOhlLPmb6UCDFWayn7OIUb5tC+wX7SCbQSTl0LC78aJctzYYdzpRDJe6NUhF5t
1yg+0NEkNU2O/+gBH7QVy717NeI+XKiVEJlwNRdt6l/FhhhMudgwsezOL2qCJ76PYXNUx02iXUMb
LNCIPaKLhiPooWGwQX31GcZI9UOBs/VvrmBKfB3WewWxq0fvzsPqRx8zw0y3EOHTzGJ6BWWlfYwf
hBGFaaIvJx5mvaWUWFDPxZ/8ruymyfxhIIOjcp2JzlRragxh3+xUb5VP8Ld/foB5LnmmFO/XVQxu
kErKm+NhQSI2JfXdd46dQ6s2neBZxoaVyB1UIxh9eGBQU14EhuIIk7sK1L250RVT3/l9eFC4g8lK
ZIcMJR4nrpZ2xFtRHxLsQeUsVUya4FJh0FpY2oBKuPxQ8yyesyZOTTMaD2L8gHg1DKeL/1gxrVVI
tp/8dUS2sTPg+T0eeGfZGMOacBZCH0KhfZazQkio/R+zz6oN5vLqquCa5g8Xy9y18mAK0tBL2kK2
TAlKEbH/5AGdlq8ydlATqRtdGXCll6muFGjsW4vXIE2Y7PIL4Ed6nlQRv13IETYmKd2C2k+sVPSd
2+gnmEVYTqC6bgAo2R6VkhUu91kPjV6hjpsQEjQqB5hBqYBtb5TiqY0L4AldAN15iigfjxp6QIh7
caKCxVVM7l3AAZMOplNJG4tp6oph1FjD1jOoI26+DeaeaXFqmAw+b/TcpePx8XAc/x3XmJVELkTl
2KWCwHn5hhDRmXPCBN1rK4yuKlPxjzauptAsz3IF1C3H4DADxZlFHDZJ7AepdBwTtoxwZoDpXV96
OoHzIeVT0GtcZCoGFTrFEjI/++CZ1xoCbJPvXm8IgcpX8W9tAbki5rXbrLtcdSLyoAhrXyl1+wXs
H95Ar3NNH4msCTMkka1at0ihvxphcJcDu0+Ad4RrsAc2MrZ9DwNa/mWywRaANImwAHl19BHPSnPq
tdsLOA1rIdkeQW7z+J3dGHo4CDOTiCpwvwGkfcYY42L6wq/x/IqBlucRZ9YZHjMQIEbZKoA3ZIZR
XpsAsVD8usBl7ewZ8LPXcU5ZFkJdNecYtu7CvkOnrd9Qozps/XbtDEkaytthodp29f0aJya+ChyC
nLtkhRY+N2yPz5RuCgGVmce6IcF01lm6SHbM4t9ytHGU7Hd11vzQFqmqV0+fzLUcjVnQMyy+LCy8
hm3zfNhlZDSKQZQj9LB+oo+Tc4OFtDaxeHSbaTIWj1zxosa4CXBePI8Y6BIrmxC+EIKoiao4jW1B
gLFdD18CKCjI3x6H1ULglq5Ytb5LfCweLVS38We/fhJTbTMtgeFfh827vS+EdUznAF3qczcMJtFr
YA3VkgcFSHZ4kBEDexcB+A9C6JG09Uy3+wmL4MdZNWllOG8vHyy8vX50oR3mWxlK8G9qTdKJo8su
HqdSNuh6c3YgN2//ZiTzJ/8K8WpFlByXPu+Z+M26xCL/0QgAjVHcytOH2KE9FHeB6SbjCYu6hDzq
NFsyKoYNi500nlEAHhmQDpcnmuuDm4I2arzG0NjszQmnuvGh83hRfBWF2ZRFtLkgyUCAbZAilCDe
mteyn3iKvpvaKgkmJEyfAW1IGaShdw0rr81i0SbsVDLk72y1H/x2Hscc+sfATRGsixl5Z+8MTmYa
mes5LPnhyOnIS4N7+2hJSwNjSZAQGp2w37uZLyAZ4cO32VQphGmyhbjVnwah3nlM4kTuGf77KCNh
mJY4a3+JCJ0iNPrp2jMxzXPZ5Tfplb/68QiIMuTSsE0J+3ZAx/I57gF+6SbVH6LKpWwrM3hQtaOg
sraBAx03NA9twqd85ornp4RvG3BbiTJHXOA+Y6sToTbCVGKEH4auvybavORZS1F/b1ztsAAYng/z
94UUrSySjHDxNtesSQ2NuLRNUXxYOAHiePXlll0K444vqU0otUtNjG6ei0FZm7FHooIpxe4n8QQC
Sc8v8Kkn+SV3oJkXhxzlMYkRMmXtSJEsrMrX5fGfD2KxzRFwvpp+RR7cHWt82Wi5uGK2wFCK6F7c
RxevYUadYMle7VJjvvjRQeiQ0EH1D6cI8RuHlelQavEPODwxtZ7TDSYlq+/Wk6B8+shccE9Ipgdn
pE+5acnQ9clGXj/Gs+anM3GF2FXdcVbc8EAOAONE2rEZL5L5Wjp8evxEmj8hItJFjJJr/4HfZ3+K
wqF1KgBWiNF3cj0MymU5jaRbvoPYVuYSaP/GEjf5wOjY2H607BxEINIIlV58QwAYD8IWPo6x7b4d
nzSFNYrt+ldAIgppqGd6cUy7NPx3Mre7aHouuTXIrvsXDCCqF1NOHfwipJr0qUgLNOPjPAHNmang
7PMoaC01rdnRa98VGRFZ2ihXuc9Ubq+ixH1CsHIHVEDivpNdujWCquQ7nY5obXed0Gb036azuZJe
OUs83UbdpzB9bKQfmU/jsbio2anhWMsNGDKLd+u/hPMkAX9A+bK7ACP6/l6ZfYpW9f9FXwzuVWmZ
7KIdNsycrbNR5SgWG2cMTFRyToRiqXMz8eWLAg+ls3kwxtKmn6XUYWFdz8MMciLvHl/QebOwNPy7
NdizBvGbops2SBrHCN9N3CfIy42dnYzG2rK5jFcAvCqIJI2M1/wD+88ByRWr1hJ0K8EtSS/1S5aw
L8E+3vOO2ISYPmTMeOXsAjJopl6B2k5BJPrt6hJS8nbEgbUSFmyGC6JhaKZO0RMc83X05J+1KWqm
pvU1Hyz7YBFabRBOr9MSTu3UOgFiyw6VPkeKsyUNev4oohn1+6XH/dJtr9LAzuB3k4rNPbs90XKC
yE3UG+assK/+LFD4CnEK0GD8eECw95NAIwDcv723X+gUFRebuLX9B5RlET7cTr2bRoymjsBNM9O9
60MVx3vpak4cD/i7HmJm6Bmg1T+5bRPlNGUgYU+UpeoUUScRPcnrC7IiPDTx8RY0dG+W9/xeicS7
UGGp1PdlbNEzkN7aZWGyrPgIL+4MaHAHCG/Y9Do2l5sF8zciknDBrHFjMQ5cbDlB+41yZvTtEvgm
9rxgfkwKUVxJbBOjzFhYDNtDsPbVXibJd7CfJfCZSZGR0J3PJoSYMOCyhzHYIm8CKtlyHXRCYzwg
wlmiQ6pWQTwqDzplgYNT7+L4ogR55D+5hytpNj5jrdctn7vr2QOn4uC8oW1VB2XXdqAoYC5Vsvyu
N56Ah4JWP53+cKfxEQvnmrRUEUluRTBI/BPmRSXUgeDKCTGZ8TeqrhFvVqGX3/jnBJzSwFyNB96R
TSoVSIdiNIsxBibPqNJBXy2IkKbJvFxYqPWsAVJ4katb0eOfCTaXvTFGgxBAuAkT5c1hQLcQx8OR
J//A0ZoWQEugF61IeCiL1wV7VJd4jsI51E25qcvyd6WfAuyoX1xOg5z1Clpdht55iR9bAxD6fnIq
WjAJQhsYm6LJVIT7VpO8LDgm59jXGRG+t/d5pSm1N6+oa0aWEwai8E2gW94c4EWMCxpcIJtdMG9i
m6TpGuAdLmswu2uYL7mYZU2hbgc8P6pwuJ+wNzWFrIB7TgwousXy3BawLy88iTcsDRv38yo5UcMR
rR/dNlRp9cgnJu5C23nMjDnIYyDdbjoW6AaYsP5PXKXFtPdmIxyE24cmHYyvnLsDaL1ThbSfGH2q
tA/RP1mgk6GGV2dZgwq2iCf4VKwIp3weLlGUkeP+G3T3JvyH9BIyAYeuzg88SBpwsBQl4Rkb/lVl
/n8gFIg8GARl6nFAHKiMVgXp2BC63MxDfXRl78lAvsW18jzRGCuDYaIQB5Wo1c7mrHihhaun010m
aWcJsr9Y3ApV7oB6ZfMTnJIsafHS3EcZMdXIYX5SnEXZqvW3y3zOBnAaMdLqccWXBXoAvkEiWOnH
+kHqFms2Xya4g6BrXgoMFA52OxNu7pCgrb/uKjL4XT5oF4o2w2BE3yqz2IyN3hz3a+KlaFJDjEjd
Trx4VkbM1XzJuZsfcvGqK3NpWx14aGGb5LIGlt1kCjYFPYyXpFOOuUdTM9tQxa2HERXYKvLJEFYw
BfqZpKpx+rJsY1IE0ELRs2sLZTbO99H+YuWw1vmIHlaUT3mTgNeC6rlM3OCaVh+41iPmH6ZP4ncl
ZTXZz+XBpzpm6zAhuWGSIjWcqEfQNC7+B2TQsLSzGz1MC8Aoc/6hrj7Ff56/2bKw/bh+HMtUhAE9
loRocYJOxwpF5pDFz0Sk2zOwetfsPbV90OOksKthBCvdIqwHMenj0xcFMZpHwG0z7eZcX8uIVhML
3g4eCWtqmKciolrFolMaLjayrPtoTAzyIzfdd/0AiueHX5UC3yNbO5GbVes0PCae0A1ZdjwVrybj
uzK8uEtQVZeyA9vkWk8fKLzQNwOTs1Ov4WvzffSHAU44jFHD0QaJ1RFOpTTa0tXGR7aw1QYOY7pT
Ojfh5P5WWnrlsDp7GT6R+kbIDGQtEk9LCTIvU+QjNAkaJnzNqxVnPTui7KVcl0a3aap6MHymC+Ka
ZGBMJ/bI/ahP69BJL2RHFjjc7yXyl3ik7hgyE8pvAfyDT9zbJ1ZNWXR4bjO1WU3vfbhKRe7eLIcL
c9p79OOmlDAMtCUmsMk22+6/vn0NX8Om6jWBBdxUr7f6AOYnYH0cyNGGGnmQIm6AiSToEe9/BwJX
3KOE95cxDD6aXeFQAHEHufVcwZcd0NRRpRPsBTVRTZJxl+apcsBmSSuFkP0PXiXO7sAEBtyGgguG
HveF91n728J38CtTSVb8ZmieDu5Mv0bq7xAalb+xw3Hot2OwCoVNQ9u7XG8pjwBfuKa57JZJMgZY
Ujj96rb/iacRBPxXsJZCyfX1lwJkigJRKMR6m2y7diZzeFPOp836yhx7lNIiJGG88dhZioWLenU8
HlbqJES3MIqQOXKfBepYL8fVVZPzeFnyUAm7S3i9BfGrBTAtJC+w273tZUqziyYCrgzMVpADTrSg
ijpeDGcGK3YM6WRkJwNP29DibV6b5vmJhhAJpsWsspowPtHk5aBlf+hnSZFXVU6h6JEjo/uOMV6a
3DQtD2zk8Rxfaz/KkspVhSzSi3zooT1JRzmfSmHVOsYu1xIfnTXsozk9JwBZ/ZUvMT3MBWXxENoJ
MPYVm8EOx73la7cC1YT0lkqWcAqxAJlUeoLT1QG3uvvDbZdweSfP7BjZMi38goehxxIDhgbGah8/
VTQqb6I+iJF+c0a5HHMnozDgkl8j4xzSdzWuqSjmoIbe/qdMsZVjnjGrl2Ip4Cu0mM30V0d/cFys
8oH4gsWAAqDKzc0mCTiYaf0b3NELdbo5HMLDx2sS/LGeW/9c8RY4BOCa/A/hqCWnqNKXntw89mzy
wySXHCMvOyVKHJ0QftK5vPLc3FDr3CkIS1Vx0EtJVfLEY2x0dtdpmbXmGZNowS2N9Z8rpoLgg0st
073CBQYTu5ujnE1hhY4DhhgLhVKhhPqXGBJdZ0uo3pwjQotiuE1J1wQX4IyMnzRvyygwZ2khi1Bx
R7f1IFTaqJ5JvqxDNpJCN/uItLxG/JAn2sUOZYuuSvBLgkPV30UAiDfLejuRa145aHqaytRI5KFV
ElqNFKosq9vLaU6s8WYkdxQdZSsewxRcpk/gbMfOxwx6V2G/rcdTEZGY/xJGlEp0VKJlrKgY0GFL
32VgcPW5WFtjrBz3aI8AZDCmPje26a9suppKLc2+ExO0emTD9TybMeHC2ArvPslRynXP6ZTkOnYl
m/btfNKBe3Y5B1QvMnwrVxUI4la02PCchPRk+z9w4eFPaGl6WoisPOs6hRdCkOrElARYd1j8Y/TM
5Pe+/dw/3jSBGRZv3Fx7TKyiserWBekbzFIgwdFjNWEowtiFAzDVlt3DwstGczR2XZ7lJF6ckPcG
GQQoP8WLwxae3YzLMYjdXv6ebLju6Dh1gzDowsSyVDUg5zlE+ZqCh7opZa8L3yZKHJOZxApOP+nQ
a8iWPdCyRruukeAb4/ZxkitK7xpVZRAVrkxks2oo+sg3U8+UTeXNdEHEAsOUJ2bJTDfAFu1Nf7fw
bMTFVhkQf3wdjy0GZrPlDIRDcc9hZi+UUWgkfAMutISXtbY5hfA7rvfbqAtAvZlOVhm2e/Hxm9Uy
X37QznE5Z/KFNIeA2VDwcj9tFSAJjdPG+iYFSZh2OXcuFIhnkhx4WihnGL4YwAKVJVMf1Sm22pjU
tE6K+oM0qn6a672uqNyc0PUMNxmOCxhF4Y3au/SGMVD/UxKrRpAfRfwzaxsWwjYiFJDYazfeqkpz
tBv1OdbnjSjeHlS2K3rX48sYx2OEYJIo+DA6aX/ruRFTCn61hvLuy+d2n2djAEO84/JiUhU4ynUK
be7RaNEk/57UpEJFobdWdY/uw44WkJK5et82of14KpSy8adqQZciz+aIYQyIDJ3woI4ClM3FJlZa
YS+kJZ+Z1i6ci3mJymP29kx7yB4dE0aucCpLPb6h0dUUx5gSY4jTooYya0iF2dNPyQMb9pKg5boa
BgRZDF7m+aaOKmRaJbtqwLKqSIPQlFZ9Hig2gedQB0Brw8JBACtunAhK0x7DDp1cRxD+t4MIYcb/
1v+Vd4lhI11DiLCdl+ePL/fZ+GPHMD/Q2/gw1VWISXPFg3U8bMVWt8cKkjBzxwZqIcOeQ3D0wLL3
UFjEkEWCw34IA1ieQ0gnQCzE2Ek8dSR0Xl6NDQYE7qRYQg8ICof586DmA7kWJLAfHNnp3uhuatjS
IlcqmSJBaNm1VWHqcFm8CIFOs2XnhfQhx0+Atceo43UX/glKTjNOGYNu56t7eXG7iCNG7X1Tgfk9
Vu622Npvtez3YqMvmWF9eVwMI0JbgjPLF8g/XqKeYGo1R/RbHucPoTz3fACDFDx7j81m3TrgIc8I
Bv7eMn0hV7CHeoSgA2TzFCLdqcdDWX/C/4k3RF7UfUvF1u9ASDXhlY24FK4l/Zc65wyYTQWJU6+u
efauETqYNj2fttKILJ0jDre3hKz9fLgG/9ptduC7Wp10+w4EVyKi/YFixevoGG8WR2zkZ2D0ivt3
GYDFm38Kh6DLpWl3HT84tGfrmgmdN5TEdPITTxdspHnzzdyAkZbl3Ma8Zbvcw14PR0kNfYxF3JbN
55HvKp1BI1OuUGmW6hARCkb4tQQJ4GPxMQViIOUBod8pYNqJBxySQUjSzbFw7yXQU/6BDRoXSXAq
yysMHGqFZsgNTPo8QkQiFlFqDpCKa5sMRujFsyPYWvXIHzxXdp6fRKdq7TDpoA3VIDUaNFAOyNaL
B/t78hnp+N8u+7slYygrqyau1Xf9Mh6bAE1fMZB/54y+e9ZL4bbGDA1vQm9+KbatwmSKMXmRoq/7
SFQRPov4teftfQq3qaN2GSjxwaGtSRCNUqhosgRrpdRHjz/AWd7jCxKurUQcEoWx8F3+h5BNgNr6
r0qxYUjoCuDOSiFHp91CG5E4Plevx3BV/gApVgUuogvVEyDLgdkVYm/Ahk0MhdqTDfkX7i85HYuI
4CgfQPlCZ83NNzZsMdHAEAz2g9lsmhAvSCEov5UcUxHLkCPJizCSTQlEiCcc9Pu9Ud0MIVZm8ZTh
eV5qtZ0PVx6tuu76GFoJ9Ccm1+VyncDmqHFpaaPreLFqP/f5BjcabeLOrBgyMVI02QLF9cCKWTBu
yCmBPFgfKAxSrZcAMYPru9oWsFHDdQCA1HZkyMxO50n5Pi53yEbdu7egtXQ7hnFCHwvhhRtOHot2
4xUfl6he3PjlVRpKE6RNXLGBnIP229gqIbpAw+keGw5OQmIrpMBvD+1jZKvq0iNbUggt7HL3cQU8
KhN94mrFz9zAdZrjwMJfdVbO02O1b4ZO9XneqWC7Ceaxf4CnnbDJJOTqams14sPgwT+VDDmN2kCT
p6Bwn01M3Gy/PtXjkPXWh+EY1l/S3V3YDuuJ9uWcXs4UF8pDvt9T8L7kQujaXtvgjsww+8wHl4oB
erYrMINoiIK9wB92SSWOuAGHI3cizqpkkKbvtGLYnSXBGQhABq+cAX61LYaLEwvrcCAdkNNCbSqm
EZfmdjwOpFvZTEsNA2JBOkQc1n/1b/Brs0dlKEmezjwRR5jMUL6CEFCHI/kde7ljdFmejokJdS1z
E7WoF2mx0GADGAEveL+OCp2wC4IWGH6Y5CqYQ4fvl3pnGuc/oE7FQrBWcNbbJ8OpNqUE/RsgJttQ
6X02CvYTRjo8BfhpG2CZYfOnBcrOopv0N2Uj0EvvI5V368+UgNLSJGR4rjQpbBfvsWMQYYcz/5UR
81LJFzyov6KkL1aTAiav6Lk2ft0eZK2kbroCET+mXxeUytkPfZpVTIMR8hwQAgLfC5OXuvZ3VfQu
FrJJDy1bYF2TlIQnbyCFbKs7x1L4Z4YsLSjLZULgDjr6swWXmghbB4fVJb8ACdHFZ1AmCgzc0HiW
zvxUHtkQb9IgriPRzFBKgPGav3ISDf31p2R6Xsb8EBivrGQAqb1+7/aovjcQe2PA+IXP7F4CEteG
GXm9w1iyJYzEXFPAy8TSj4jueFV3v1DzpWbReN7bxQUzM7j6xn1EyZR7nNcZgH5x4f2MnyZZOnS1
ub++TDWXOd1E7tjRGjOiF58x7wucNPX7quHwE9i/eI2NU8fKk7GlayKI6RWft5mgcCvOff6Qqiaj
m7WVkKOFHkZ30UWSn43XKPxkxhiRuqDPBw7MBC90F72XND3mcHlm5h00IQ8GbXvj8+3swpZmUCPF
k5cNA3TZMxVaU306rQJd2drDRgMPRoBNiofwGOWaQUfh4tQlgy0Hac79PMzFCrbIjkqyP8Do9PiR
erqpWPFA8wTtmBMB3LT+tKMqEsuYRfFAes2eyu9al0QrtCxpJRoBNWkI3dvoqtGqVYJaIr8GmqFO
+W6XT9ukhfMyKi7jelECYgVxMS4UEy4ZxSJz5AlHUhFfPtpqGIkNItuWHBpwMhLzT6v/FJZ4egTh
LwYOAQRB5/HgcW8EPgjy6NEzyrwmNcr02ZjHwvfpdd7sK44POjzmx2ipeqZ3VkWdCj3cZwfjhQ1A
bBhjV0L64lMt0U0va++ftBL+wOtllLiXE9ixZBiQWi79mo+Z4JPF0Imj9PRm9S7sV/RM7R1nMb2H
g4Ek1K0UHmaA6IeVebV10wLZWXK4WzODXFj5QNIyMeP5SxK2GfoQKfe73Y80HP4Yez69l+01R8SQ
x5lv/4QR21BTiyVPlufHIrqsiY2TxkHyNPwHkB5l0DgDt0UNhse5ObBsCsALrP4ptqfv31FMKx91
6z58p7qwzs5f842UPbS1PWxKrUmLuZHKk2mOJLqLhEHD9PB2kz9fFfAS/4BHRf8KmjZKYlHQF8br
wOCWFSfUjlJvCiZaPmuq4zUKtnp5YbzCiNJfyvOLDV5Gg3deguKTyklvuMbfqUNgeRyynV4pOIXU
+NpNRWfSSRB0sJNaFY/fBSpgmVu/2sJKBWJjcARXO0DpgJt1r+Eo0RlFB6rYnEkP3J+a31TVRCb2
oSdZNFDrq1Tw9vojKq/Tny3aoOyK9JrgyUuokuAH6XiPTamgBtIt+/abSUy6ZRWzS6/fAe7qMZZ1
xCZfAJY5VCFE8TA0eq5TU0I57uJJqjdSaVs0zLJs2oH+jwXyToVmGcoMQXgfCDYR/M11dWytheVl
dwfWmhMNRNhBo/JDb+BqVh7Q2CYjpDyE14EXm1NOvfEfm89R0IKc6jJoMRxQk9a9VttidrHxCt2l
BI/ShFMSiGd4y6TUHzoRNgX/X9GHRg0Bf7f9c9pEbGg1peznkcDMLNziLkXI9PSR+mIaF1tkInK3
kB+fwdZ+FEQD1TRfz59J6d4tJCAZlzof2sRvxB2tH8MaBkCH+u5WFbSsdKjRgOVHQ0jmGiQtGYgu
D75lhPK5m+E1kuG5ZA6iLoRVtYMFcuro1hiwvH/lGluUXVDnu2Ct2o0izr+aOKZj0pw2PdOGwsZJ
Ms7uqKJuXYSld1AFBfrLM29bhxqLrt6LXvWcz0ATA7yHhhlwil8rQ0nNWfMSpnVvsw0zsXMTBRX9
iSVfKOUWPXz+LcOmaosS7WvOO0h/kBJrC9jJAEbJIEQkygEI6oOh66gMwWqVmYDAYFsFnQYcGgQo
BJj3KODkzEqer/JXUjipl5m5yrcRYK2LKWGVsjQGpk24Bl0FqARUjIm3AetLiKzEkRwSJR3jbp9z
gYfe56KaQlvtNGnXATVdQkQzm20N2eUbcaaJcomtsc1Rl0kKvjqLfDtkFeSIkHIvp7Uq8lZlyCyt
xW88sY1M52PkbFrDU5vf3i0tYDKY4NulzDmvwVNmywKsOjtl3rLpiThzMKJexJv8aPQ4TfLAQQoU
ExjG5ZjWDdOH0XsUlE0HWE+XG9pR5aAIh9XOYrautRNjY0WFiejVHcNJMfm0NkbVkURVfvMpf2T4
Xw5jbkZmz7FePKA7sKlfOFRRDEIlLxMpkqlh5RMX8RPBPg7JoUcT72bmdTe+h4WbbTK+BAnKJGRV
RKfCrxVtk0MHkm78DWCgoT6rVG/WOwGegDyX4lCReh1VVkXAWex0QicN0ZIZI+dX3/GxRAb4nkZk
hQVskvnrKPXtor5qDQxxsRwyTwxoY66TNHA3ga28thkfDUus9uA0HviZMWQ2Y7svE9Kpf6iyHSrU
bopewROO1HQacp1jpd9CAaSfJL89m4iXjBl0R/GovyRUW8JPC/ncGyQcZJ/tqcAsOtovUjELZgU3
mJ1mYYWKzXJgL+/wHefCDvli5wTT9Hc07LsDVqDxOwJxxsOguoDqRbo/qz5ajqTGvSuqqsz5/J5R
NsuO5yasviHkJ2AM72X2Cx4HAuO8s72d1BzdiTEMiTnV7mJP+bECXlqp6c/nmwtJXq/ayylLj4ig
hSj5T+9hGI3JSzym3rG1RWgKd41US8A5edsiTn2GbdkqHW/AYfYUWu3F4rv3I5zT/VZC2O8QRx2T
sLIb2OdQC2uJrucbJU/Bwvbbz+fuDv1qExh0F9biWf+0IThFytDIV36l8+bxLB74n4DnTPguPoDX
QB6Pr9AWssLAFsspe6+se0YQZL3CrGTYJRSkH/pO2HgTwIoBHebVi+ZttekARAISm+NrKSbBvvjY
LI1HGkugxbFrYW6oZFeJIhnky0Tlc62oVsDyvPxtGABjwKCl569WXeSzpxoJVjNJrwlcj2tiR0ya
8ariRjYii9mfcwEtqOWSqS+Zh2m+hGerzAyNJveeOwjPu2860P21IHYao9i3DI1sIZRqX3Cx+guT
5dRKJFYVOUo1gJZz0ScVYuQmY0Zef+H4LBJYU5J4b8/uy4KWv3uf1WOnPqw1cPxykXsqmQuGuhxc
O7csIVudUlmlVWPkytFSxYtwC6EKcPB8wJ2tShKhSxHU3T1n1AMEDbhkWTlZIGwDfazroMarAA+y
opkYCh2W4rApcAaz7SMUDU06XQXuIDPUVsmdVJpExygQgnzAdfX/llfn2VctC+2K4T+X+2oag/Bs
mRHgYf0M7bHVkFkao4TqyNtA5bg7wRz1NjlKEYe686dZzNdymr9eF+Bg8yxMmp2xebEMKMvpUvFg
UZHR5hE5Datov/sneHpwomND4JuSEznceXHDr75CVRipyynbjDLlkaxLiu0SbYiVild5aMLZE9yG
pVSFzyDJ9oLAWARgW+GmiXKU1tv10jUHzHpDeYh4BG38goOGnnk++O468v+xEoqdb8QQiljRq8eq
vs7IX/+h3O30wutVGHeY9Y5DLVg8qD9BLYs1OQD+hXF+BtCO04E7rV8mQQDSln8DDUz0c0XI6CYr
gC2X58iZJJMds0uO2fUgWzs612sCg2wjHAUtHkyiFl3vzBsJiC9JDt+bYJcgryM+WlZW328+NFHL
/Q6YSGIkXdd73QUPi0MQkNCyzE/Mwkx7kmDMKWnX7bpz8Tf2rrFchSAQ01r1hIHNj30aj4C/elwJ
DUah6NGT8WsUXB11abeFB8tJHzp2u6tWmDLODAVhhi2ayTGsj1GcyqT4gYKn8LUG86dg2eHPvD9t
h5tHwuFmqRQXudSPddqmi3/0O/qXGjOcsUeObwgA8+RDQo7sJGW3IAsiVHJz3Z2v14P+bAlgYyDF
XARnx3hSbwo6VZJtFZOiovy+9Oyve7+niDR7ocft1kgaQk4dogd/+mrWbRA85iTfHXTbEXGQbsg1
P9wie+miHus/pD4dEg8qcK4p0P9m1EfYRiOHagr+d/EUsvy8tFf0ojIpUSLXiHhknDQfIUSwNEUG
O7KVjtrSWRBmlE2iYV9/MUlLYgDcTDPniC7nLkA7+/fCCGsQibB/a1LmQ8Uh3ohEv0wHvb9L+IBw
O+aaQz2FU0n2kW0UVC1XpwFfQV6y9Mhd4SO8S7uDCG3JMHRyUEXT816q51NF9gCbV976x/n/eRGj
0ASCI4/NuMRF78/6SKR+0EtIb4q7NV8TsCAE1geRJqoHkRv8ncA4pcFwlsj1j2Mi5g6qr24i0dhF
Cjei/Fs5xrxi2gXSIcYmQQZKCWAleJa3Q04VNH8CMuUKLiUfmXFrMgKVSkmXpuB+3QokwLJKFu2i
OG+JVxui50Om1TtrQedMwNKr04HVZFIRKJ+hEwdmiz1BNmZo8RwW4bvG6rLevBA1IOYUOsU3mq6p
LQk4BcZaT2LaVlQCDcIkbjQ+NNhpUkeWMK29UjXLsI7pc0483oNoJvkUoZMY2kKhph/3eN8OdOjH
oX16M7gARYzTaoB6ntpov8gyjfOLmxIL2QpvL/2qF8XGc0CtN9SfRRzOvPzzi7+qKxWtH+dg9bP0
SVochjm7c5PVtr3Fj/3vZQqpo2nsWekBCKfcPskRpV0We/Jsw54tobrtQ3Z74Go1+1rAaT362YI2
E/ezQAPIQpbqKebGFfwjS6TvGa0/755w8x/OzROYlCyTbtRmx6kiIO6Ir1haTP45e/y2FEL9twTP
kSdqSiPrj0BZfICS3RST/IH0BK3+VYm5OchahjbRbN9MnR4auhiuOP+yWNsPoWWEgXGNfj/0Il02
ji/23qZUt7cEbMZTfHsCb0ur1bD+Cth2CWfrOyGnolEvNGXML2vVpD3tFcOzleXAaVyRQ8ifJcLo
x+5Ac/hnKeAfB4nrhmP0uNjl5sbHLLy7SfmTqGDIuhp8GGiMc10VhJz8/CglkGSCv8pgT13usB9u
0ZqX+scXC2XZIl4Pthtoz2d9XbQVjelG4av0+H0shMkzQj3d23IrsFjPzP3BLhHzwwV5h06JAfGl
BCaNH2Tav2558Xl+pxUb9wiJHMfh4ZAQywLCG+K/vyBpqGfWQa4v3pmvhp1SZRCvRiVcSmvKbc42
QTm9+BPGu1odnE4CVx8PvrJ9uqEmtdoJ+gWZCUzMEx3Vu0hjAaLDGdPKdU9YHOlO40gD6PskuJAl
fPP99uWyNYG8LXgYEBsNKuqS6kWdpdQOkdFEiZdLYb/HDPvb7lpQ9W3B6B98N5ia0kMQSSM9WYEg
IEsQYMhTVRhf9mRhOC8Sjiyprgu5j2yR+PlXMyFyKxdC6EPIHj7mRagPxDhPRLQ5rm6vqGffpckW
TkBmT82GuqjY4mjFyOuDcIVTuabI19Rs8dBBifHv96vkiFTCFULjyB+O1r9xndugZys9hmOKPoS4
ayvJR2j19ik5w9CVUDW3lwF8xe4ISV9RTSB5+vm71sPq65IYz4nYwkeu1dNPFGK/O7F+AZrDhJ3S
7HVhsT127C9nM6dYoKTVrzXsJC75K8T8HW2jXDddD6zu4jpf77+ydWlFKcRNwrnOk5reB4UzHmee
LPqgT8gxxOeZrKfmIDdsIl5n1VFhbGCotdUhx5XlWbbtJkILlWCzsqDgni4ZDidjlpffl9QMCWm+
OiMQJWHXUNAYb9vtM4Il2CcmwDhhDSoZU6cp5HHrL/mJeLCemRkPxFnkLt1cjL1wiDIvuR7EVF9n
48ecFezpqUMuhRuGsOTMGfWgPw6TLilsh5hM9ThrUHOAr/NiRW4zFiMcGD4dUCoX1Cs81AOABCQQ
GMhkNzz6dujswcwiMiLGPZtsiuf3S+iATLEqUfKpbtmOALLaHjuM5kT1kHq9HfhktIDjhlYM9Wzz
28iEC3UkuhBJSeAJB0LQaEQ/ekL78M62vRbvawe9YlR8kbdvUfB4ZDnyvWIbIT/x4065rQiVNueM
4r2hns8kcDU1mNJtkEepTfPpdcpeStoEyLlSCx6ohe8xmIrLkLgF5/s1Ie2zrk1e29vKoHIl9AjV
Aa2y5qF87O5Pz+cAiTJUKBCuFkBAN5ABevaLEGa6H2e8pU1zy9TTQsJ3VDKc8qjbooJXGtRywyId
48zigNC88Ho2SSVLFwYl/kykTFXwaTSojgphqfz39EtHh+kQ2sGhvarEDS/IvOLPuLPMNgBbplO9
iT9V/kgpMDQAX4TFvdEBm/LsG556A0HC0Xr+vi28rcd8W/WKq5Eww5ocHv6yLqbu7Gdat0deOlVp
KE4bPjUhE+THWekpWKYeZ4tu4h1qURGNdMKeJWOE1vaKYjtS6Mv9RjmRN/Nl0fPtNaq2QAau3QMe
veY14CKL6QCE0eoO4XfzH//VmhyX8J6QmeSFiAAPo8698DUdYxMA186v2YMsUSxsFauTStqUX7UU
XSwTf58Sn3tj+4aP+UM4E3BEbrTRuoi//7kEU7ixPT7U/Swm2AhGwWYhznxxxYV8d4HTb1ZRZScf
VTURDmpCba3S6T16KNMPdDWQfocfBzu0OISzmthUAUMxho3qQBmyGBjQWpYJ2L3EdWU8QeFG8sxM
QeH8nCNgCTRqQAA1sZGsQmqeWs84I7TAIl4Ji+5FapiSVxp21s+mhaEHGqeSt/Xx/8PinS9mAYMF
8moAWbNPchoYqR3dBmh2MqMAYncdB8pxeGx9qxlZjFzQMCtzO5wz6Re8sSggXyOS9LoYnz5V1Yrp
3V4MY1okLY70AwGe0RrB5jVkieUktpiXYYK4UcxwaR4Jj5fKP56GTw/gLGQBmlHJTIjTav79EM/6
6nkHmXYE927rXmGwGmt6fRFQ72jjQ0u4j9QlRTNSsXrQotK00GYOGyK3V1gtskofEA1Yur/cPern
OhvM7WQ0rKwk6ZpVROHXusO4mqNZALsM148WOIOlIpeFjfrZqrm109JNYt/56g8ecWrwmJko0jXU
wdaNhEgmNZhJ12C1/OPnEyqYr/6foQbN8qHkba0HoFV3rX1V0NrpkiHXnS/nvwIwr4w9LukW2me0
Enwd/6pRvncW+8KU/G9Y6Ka5/SwMTV1cBghTP9bvqbuDR0eY35j3hujz8A3LUpzJI6Fq71jWD8pr
p5SKCq1DCfU20R7X3MwkFJfg36YqlR5hxgtWw/nxGJycQvB4ahwDYDOvHpQFtOFWfv3MicPSOfZA
QwCx2usIWF+EbFRpGU0zGARaCBHCB3sl+w9FIG6K6jyu9PnELLk0KSN8VUVRo15gjcPNe85AoJKk
X0LLdM3lj/HhWieeTHypHaYvYe9KK9MrNN+FRl2NTJjzqgnna/9c7j6O0y/WHxpFoKSPEY4APeMl
RefQKNveg/rT6fL0LmMqv5fQEAhU+Pc9PagiZ3tBeu1HxbGwKa0paxAE00wFIMdwD7DTzatM4cVt
OQ1JvFoEPKT3n46l6zwfeeoIPsIa+QEyd4VcNj4Sxvp+zp0Ro0wjdaAxZFcwHPoekC2vDhP0LhuF
5bHhNRX231oA9u40WWQ0oZ/Ma1eqOC0Iy0VRtECU7fdPJ2IqVoQarp1ObCorecHHwqFMfA1R+y0/
R4UnHvIm7QtdJkVPgwbYGsVXu57v+I+Jk5m5NunCDK+tndsyuPcWfNCfz0SOv8mzun9d35COiSBI
Fh7cdde37d6znVYlu0Xq0OxWPGWbPxQVcIgKpj21akpxJe3KYoqhX9/fqmvBSpecywxAdpAW/BnQ
EtaiIkYkH7MLBD7KDjU/Gh0Vkf+80yBgyFFxYxEKTZLZBaB5t6sfjfEOfmiZONFurcpjtn30B54X
y+rEzEbyef09OOXCUqwznEaEzMvANw33Py59Iyz3GQwV5SR0jciXo6Ny7ZLvREeg7k+HJYAj0S7w
8jSJ/dHzeaLB1+yEKj6L5S9qUYdQq5UtNNKCcTEnnFEJCFuWHjBEdO3KzPhbu8NbJYJDk9hZUw3Q
LJCe+HjIHSoOeQUdQviGxnyJdbXtjubYF4PlPi3iRbyOu9ucksMoGRyOvb4htGDKNQ470KLIREE0
mL0sJfGnLosH3wA6TVynzb0DProNpM/cUMre2sjMh+cK53V5T8W2fv12srBcypURZ3gho4bnGHJ1
4wuQs8ZDXUVzXUb160z++eWiJxgKdxAQghMh0vvhbDqB7f4xJ2WCxFO2CAW3tIdbdxiSNYYba+qa
RXqqPg75gDfBC56ZT06bS9jJiIdm9mTT95IOiLZdB7TIcGCC3S8jNjaQgQSiJGsgP4/vSrEbMWYe
rP6ijreg15nvZleH2dcmBEEsk+C616UiY4J/66hOE4cr4IffVKPFKbLaQz1KO+5xxf9Nwltg8Z/R
XqhAWUIJWo6sjMo9qiPHmUClzTH2D4OjbJOxt732wlTrXyAWk4UmozT43IBwZexUy5BPDikC9vNv
JcrNiz9giGFo/XljRqILZQ8+We0TRVEDnjDd9hE5Tjd9FCvzwhcR75Kj+Wi4OxIQdlRi806DVGqO
CEhHCgl0yDlruXT2Vh21nFZk1ETOjZUnW6JyQk+OsavwMwb3lGA09KHyUOZFavMQTxR2Z5uoT0+D
pDpdbvAPi4hzWB6mxVTWs/yz2xKjdf8ekY59CDJa8AKlatQFhs5umVVAjZk3IsT+/ImP7KtEgFyr
0bLQmf48pyRV8Wwp+COUE5zMJFmcZIbLHfdjSumi0fKgWTapJAEX8ESvg4AJrO6gU2JPr9htqZFG
Bs1Fr0F6StlBjC+JrRIkQYgbWSa3UC4jVEW/NR1g5Pj11j6tzfnLj+qV+NPDTaj7oc0biHWdE0gr
XVCTWtLcC1yweevKUuXxmTruG1GhDOMxiNi4sbe5jhR5suwfRgtntnMtNng5p3Ngb6MKByRcGenP
o/85IuYOtkmQSQABfnC1xSnOgS+G68xS12cEhne/YikNF0Rpcy4avh0ngvR9ftL6xJhyrRSkd62f
cEGn2KC+L2NYJ//pSP5FE90vBRr9Li1Khku2ExnX3E1dmxoKTKRTr4vogJn66+Hp9FIoiJqFlEg9
wSwcn1QA8Dp4zz6iRTJZZBMCCoF4CsMjXe2BbhoVsqyxEk1cbkHAA/XJvhBglaPsrInw5Ghp9pkL
ps42H0H8NNyTqEgpuYW6K0iFigKx4HTjqR9ThHL+Cbot2dWMhbv8BvQrbQCqkUI3pDy2So1+U5+6
HnuOsC2MyuZXBnC60+kzuBMQ3CDvxdx+AZnlF9WOWxroRd7FplaOpb4KGu6xybE4ZL83UbN4n+gA
Hun+fjyCkDcGtiFZEYCw42KN772TXSGdWdRb3Kq8phrGI8OnX1BBEL5V7fN0D8/yOVgdK5L/y1s2
KiJ16SrE/6/MlUzEQaM0n8va5mMclgnicQ3NOJD3hsBR9sK+5atUefQxarnSTxiluivVOSMERrF4
fDV0Zvz03gkkI/lVSuKo+KaOwLR7/TJSSLBgrEy2aFzC6htQxVv30I2FZbnd2PRxU3fA7f66YW1i
ahAIwnKr0JUve5FLkY105tbcNmSRZMfp4fID2GyNcq1Lg400k/r73Cjxsb0UYRADckhGuZvzM7NX
2b+XpBTJpruL98vtXPzWpAgTpDejgqGGiTrT2kkti3a7QjwDMM3lR/faXL159UAi9mS2+ifkZfdh
bHDyYYKoMC6JTW9xB4Inkfc6zslY/s3GrfUxZwMZxz/uwnjyLqyJEhr/4yDSfeF72nsI8avJ/BLU
MBlS8EWLgXmCrIMNaddgc4u+b2fQDFpj+tIrTCcfZaDlUFmcKoNlQeKVRrN0BzGy5nMHAFr3cM1X
AZdtWkx6VRfg7OViZYi9Q/SStuIy24g5cyQaBeUcw9Tc9pGxhv4GIpzZ3ao/y/JUXwg8no4OW5cD
CymoYVQJ/1iLs+sSdfFYGsA471H0Rdip9dSaCKD+mWdSezC3x/86d+SQ/SC9iPwEA0wxA97S4m5+
vnoL5eTnqsVVM+CHugWxBsV1wSrULqv0Ya/dNp5bN5O79i9ouoLilVdVW9kBE88N3pp98Y+p3p9e
ey9+0yunwJw2OWjhEoCaB1o5W/mczkHmYTY2mUQBiBjo6pGa/RcdyVtg/0ZGrZqjNZt4tzVdXPk2
aM5DT8McTHP2lJ2m8wTjtdH6XQIL+MBpWoxn/MfEkVZ8ypNFh4Q1XxzuitzG7/03rZQLK+CNlFGq
12JaaoBkaQVEJaz9B3Jfd1eopxy/fxIc2J8zUCnH90xvGlxCj9F0Hw/UFFloARAnSUSn/TK3cUdp
1ge66u4ZQByhSdcOpdWlYiT2MmRekc+80qd2gR7UWHgBD+oQdBcZeCWXFsUXY0MqyrcTPFmvr8G5
hhlQlsbqOmy2o96oE8OJGDWeBoennJYABH0AZtHAkTgJiehS2kHFLjz6EOg/zWp3o7qaqfyvzVLm
UtaTrf0mbXvvyc4FHr0d78RAp5FPspJDorp+gJskQiBhnOZtdqyxj/VK6k3OSCl3hYOSAGi/6NVZ
NvLsU8JBf6bIe/meEGaS5RNy+s+LkrU7NUiqGvxAoVQ1tQm2+MQEXvUVgL7o7ogJi4hXltqAE2ht
G4DOBcGnfFRFpDQ9ltKRY41hvLvgTlhSfbPf7dkMUFVpD3Km0cctAHnCIzDh/f6VTjslbXHRxPIa
gkbjgnMKEl/z46Jfe4AMkDYKqnJym+7whgne0808h26bFT+WocUmLJKWOMoVMTncHRtGcN6rkMFH
0aUleB6+geC8UZAJiJP8wGysaAHlAskOvWV+GB3nNktG9T1T/lLhJo9HAWqnMzHh+optU7gL7t49
d8HYCCFA0rX7P8Dnh4WbM6UusmlvNcCrEXMWNkAnocm6izZcEJdiSkdnV9wYSu+ZIY1XfmAcUz6s
qlbtLY0NcFp38zkzp+tNnPSeAW5hsL4G3L0ZjxHQKbcuV9SPBTZ7T9RxIdYQyOZo2UED7EMSQsiK
HupFQnSRg5YnbYjfOwsajZa7G0bdk+TDmFu+M4ZIAYwP8+c03iD5nN7ie7ObgIhj6DxaHlity8jh
MJtxvGfTe/BgpzEk+GSA9oJOPrqixgGcv89iRyhBMDGPeqO1ZCugwg6hcapZ9RMREOsUm7OcBoUL
wyhvzvvJwDt4D0yv10lcwTQige4YucA8b4+8n96J2brBQSUoEEMGySxj5pTAMlmXv2RyAf+xboLK
Ri3ntQJQUjPp2dtTj/ZQcejHJAXrsMvmK8VeFUya8tj0WESwHvPae58/XF9oxYPvGbi6oSayF+k3
Jp3Z/MixgkiivPY5RW9WOMaXrz/HDyvMPqW8ACA17bFtwe20JT6HOiOijDj3gVE4DB3wGa3hKfRd
mzC87nACQyL7tTob/dAXQKAKTkbhJhczaF13kSVSwdrJMTGaVevZwREE6Q0MoEdvqnf11CjWKFat
xKYKOrYlpRrU3X2vWDfOEHRdGgG2u6iKrJLsi1/pipb1Rwy6cy9UYQk56M7CfdHrVrnlt8OmtMrG
4wsKVi90n12jJfGWU4adRQQlGPR2Aa0oU8Ghl5lOilMAj+Hzd12wAd/1+9sM8RAmZJGCj7G5izqS
/3meX6n8L33cayQ0slesMSwOnKgJvYpXiGbGQ+CJ2rm+TI9icVuT+ke7wSK/75m5dzwZNjhyVTGO
LuBpE92d8MxsYU7e8nJ8HgCScyU/rnMUUBqDb2MU7n3jFZ4U6zni3gUoc7xoI8SzwemO4rmEYXWf
arTyi1GthY8H5jRqX4ysZ8B/sSkUw5TRTDGD92hyoZK/A44Lw32rSmFm9/IWbSyBPoATtN1GtWsd
JFLTIf+B6pVhGIQHT8YW74fFk8XAOqTf/tIaG0nx/m4/wwIcQWYBAGnd8SCzd722cNxCHcRhZ3hn
1oYdUuM2FbEleRR+EV45ewDHRdN8LhswG/V9s75dKHzH7YJkiBj0Ul81cZk7qKL/ZT6C1MVVPgP0
kC09xZU1hJfqB5tTJQJExqT3VU0xBhYIUJ4LLbv2b1k7gaAxPqw4DlUsNGiU9/BBZXkl6TZ/SGxf
jc7TnFaJT1mHZxyKP0a+gzyuG3q7K8NWmT1qSZgtcRciZYEyFT/W5e5zzUmVoSAIdHGVdYaGc3aX
RGddJapBOlZ4AZfPf2NRrf0eTUJbjWaBrdey0lcZb5+68BFmmQeD3EDFHgKteV9roh5NuF0JSpKL
oFBu7XXYTOqBuU+G64K05QXSpk4ANMEG3NyVUctWsrBhPY3pC0KXmBDlCLQ9UBaC3XL+EaKMJ7JJ
aqRCmafuBfydp5WtN3GfBc0Y1ll8VPiXSRTurpqUokoAxydHe9quDBkPyjS0WItSUskKVYIjGkbv
fYJIv+W38UozRtcYiGoGcg1gZ5qtIP1Na4rd16E+2TZi2JP+ewXPELOxmt0OEt0TynrhMHIepbP9
P9kBzSl13FuWwx0MeOM2hgZfsBdeMcZoLE3UFeu96mcsILyY+uY40tp5Zz4DJsGpJkGVcUfGFUx8
ov9chJ9108P1PQKCc8bjNM1MaJSfOnx7kjPQRIzeKOgLtGX3BPZB6iJU7GKDIXFrTIFf5U+FOTPq
WyyXkUjFBZ4dEiKYJxvTLahHHR/0xGl/dUcLhnJGVUzhi3oIeo7BwOXeUnqMq6CXtrNvzGQwgJPX
vSHBLH/5TWF76Anlc/0iShCWOcGtzhVzu/3Al9R9KNkoO0jIwLZnn7ve5UeDJwAjriZ4IuLQvWRv
0Vl1HEuXMVhNTZgJleOGiTZ2sfMbjRMbblob/XyeP8r+xl10+lCB96a9ahpWKA01CxFzSczkNM7j
LHGzFn0BerEFpPedN9FTWk1FOqEorxvITLaAinKdskVnyOYaaWEikkCtdk7//c6FRlGrVqKbuIl2
6XqQdIWXms7vQbyXycgHh0k2ao6VKjYqNadoRR9erOIuvqJDZeEPyEwFHSim2iuyQ2KpMKMmnql1
JRFq5Mhe9jF6AvOZpT+Nhn01fYKKQKAAu7qdrlUwN4MEu+Dm4XAVtI48j5KIH0DXo8C57cX82C/1
e4jscom1BaDL7JAzu3c9sMX6rBi/HgnjEGDQMGLIwuGEycoLfA8zQ9QIj+5oLEJQXMPC51RtpKsD
6A8qnlRFOG57icQW67tLxwmucrp6kafVjwKneD4aDuNiNHU/oP8uhUOpnPmA37JNQ0mSNmXP3sKn
vWma6kONET7EjChcG3zNbgsDnd7ydrmbhT8o78AJdqMIVr9hmg2XnwLiXW5cwSIpKgwjVHIUZiMV
PoUukZWnmRPN9wWZl4jivzcogO1owPIFXTV+zI/XCPX98FvMHt/ANFXSGz1tlr/sFSU7NYTYw91H
yIyu86HPywyoqZgm8RX8WpQhfFobs44mwHyGTK48QpcbsbRIt9jZ8+XVH3qe08bXUMMcbvGLujfG
AokOcxrCCJRqsbQBCuzswYhS75xEB5uZqJEcZBRCsPLAx4r2hcmNt9nWtj1j+rRM1jChdMcPrxlQ
vzvN+hi5fAWZK0sArPYEd/k24+gKMemniQ0igr4wE+hyMJteLMa34mnHNQ1Gjk6tU67+D/JIljr7
NYttJmZVur+YqnfF5iY5WdHkVvmX+Kr5Zdmv/S+KaMM9EsQ7HBSkcdYu51KJYV/mL7Vn1HbcJVqj
6tjNFvMhGk5lFg7S5NMqNFQYaWRhBmT4TrUG56U3zTVMH0e8eUyLl9keRQXfHteYFlswX3C5f77W
6GgnUbaQX9ECauYnin93k01jPLrHGDM3nnHMdCW2mOR1ZQrNn4xfhEf8pOnR+F42aNwHBKO0NKef
W3yjETbUkWo/Xc4Gq53q7yIw9ZbVk/jnNZNcLpL8ootf1uWN/SHzvsDVW9MQjqruiUdrhWaF4PhD
NHE1MZIl1el230ISj5W7oc+KwOS3Tb0bq9N9bb1CUiVJmuMomcrGVCa/yOwauFo9gbh0veCseFII
VW1h10usu2MIYPrN6jnnnByV6aQsUhK1gwDjzOmYcljHlALdn3TzE1QNk2JgAo6oCUtTqNgHNPSx
azOCRFymIrWIlS7xZBVETjOohpnB9V4Sx/dm4EIFUkJg8KgEmsEN5i8ixyagK1ZypnagLd1r/7dD
jVRyvq8avMUHB2BPl9teZbdI2XshJgvnRIqS5gVR4PMoKZBJMNn2jUiuK33TjYFaPwrlf+xV5Wk0
3glnDxgjzt606AL9xZsxIQGlPmscUKJ4/fd9RODBqyHLwnrdpq/xB4OeINtZg52FQaHbA5sXkicm
k98FW8KiCF7jGdpZmpYFCR1hfKd7pdrdj/uX9twpnrFcFxXgRJQl8fmUoMKD5kJxyZgAF1QkppHo
lLYYV73x4Lr6F50H775oXiJ1G5cYm92INBkUkg5+f+/N2eNPn7x0TWPOFAR4bFEpYpKWrU5ksnAn
84xD6ALDLbx1ffAN7l8WX2ildvx9RranqCdmvH+L04HgSqInkAx43dWpk0Ta5mvWZMcV6wtHCSw/
hhAjEdG3A2Zb6K4q98VZQwiyLTFeqtVj0QSM0+RiCfLdRV44jecE4ITZhijlzmj9WhvXi4Hgq5bc
W522LdZyOSYJ/l7lvFAuLcGrYt/wV7HAwR5hJrPEwNeaod7s0pqDvX9iD4b8pck90dBfvct5XDnh
tBBwcGyeqj7f0bwuHIUU4Mrh4IXswuZzsHJcZObIwO0vNMWf+roB8Ys+tNv38wt0+/G0p/0VdvFr
gJ4dj6LJvqeXAxTE9l6BKCBhCNx6KBGu1ikPhjbNSliJRrz/M06Hht4idnkTN/vfmqhNCGmAfGPr
lgysbeLo4jHV5OXuMWJRs3g/BNS24ESvxw9GdlTlRgb1AUBy/HEwPPgHUKhHLm3Wt1sXLYH8sthM
1stc7fUmtO4LQfUK/rbzxEsVKXYcmcdvTxPvUj6bAZnKSRgSvlwv661a/GQQcMByVUp7WA+MEozN
cEUMIL+H1sBwnbAEgdPt6+B1aINh7JLE82o08LLZ1SOEMmXIhJUT0fCyAKzHOICybbYCpf6WbI3q
kzEdVA4rx1sWYxPsyqPF+ocBFxPFdRH7W2Br9t7EArH7wr/mq9KRZMHuQdgsK7x5s/DSRu2O51lN
Wf2GYoueks767D4QT0qcDRGnt14x3IRZgp/MQ0b51lbzpYmasuzK861o84R0hLX7XfbMPFdb9Fy4
I4pkQcbEUeIOzswAaTH4T47iY28zWK/k3PqTv8ZXDl4ImCdY6scdAt/WHB4UalOhinS5Utmzx+2E
8Y0YscrfAcjW2n6irMieaokkUCRoLgDOA/IHy2diZ8/eXy7tC7wNLwU9rRACyENhbTlQfAQqX6I8
MSA9nZmbhsguGxmhbU6f6Qgw6z7ICSFxrZl45AD7bYbJTyPKyvJjh8hQBzx5EqobZpPQS/rCZnFm
z6S1VbBIziosb2FplHHU7TvaxvIKWjB3bMcaV5J9nGCeU/P3FkGSwhD/Jl8/iSVX6xGVOceuuWbN
LRSqsU0MHbLUBz+bxUS/VxKDDBtlM2VDP4DpWIHwS3qbFHo9rRN5ft3P7RfqqengQtLpx+I8kKz4
T03/rHnNd562DGVE6nPW1EfLfnu5iTKiGAIbP/81p/UP2iDQBAMMl3UEyMYfbyDz3l6VV55m65Nm
81WkhxR2zKt2hVOoZRMot2GwYg03fjkWjLra976mkySHjrjXD6kHHZMvsfB97297s53oMXAN8J0F
iPyvlYHWLjwj7AV/Wlhuhban6aC/E+TKY3KWMhQTzBSH10x54NpSu02U9fO/VSfb0iNYgvbOnf/X
mkYMQCM1ogqFwgIGIGhYLFXo7I/L+yM5kWZ2LMUyAzMehyKVoXKVrGc1Y3o57IkpmuHZyTdlIgB9
L5/QA9+3VlkBfy6rsx+UES8YYVNV0liI9j1b21coi4fxXZqBotjb9tS474hBpcHUG9OfDsK/vcH4
efZBQRqT6bzWxHOQahigu58gnRquo0YOqOWwWB9tSQaYLKbMp2DhpQNDMtonOV45AwRpwtDQdLZa
hf53e8oEDVZfpBRrsFOr7S1Ozh3mDUcO+HmlLRv+GDBHtyMpMfSJqSKcGaTjP6gpAsXQq42YxO2h
wvlaKJYeU86tNfLQH+W/uzqqeRjdvo6MnlTTy0USASm/FsDx+0kCfnJtNbKojRnDKKZD2/Bz7fxG
nVL3qgFJm9G3jmVee5BHH1LNSY7wApFV4fGiDcr+Ej+cd1F9kqRMli89DtVTHpo0Uq4SWbgg384R
aQjJJwNB15nVjY5Rq+EyegtmKq0Sfr3G2II/K6VlT3V3XqTlpG2U7x9DlslP6ZizFgbSGfNqTyMa
aWAufADars31wy/xhIwk+erdCYuoGM8+e7QF0NAKQu38EeoH94+njtn63ERGKx+GePN2wDJ41GnO
xiOm57oZ2WndnPYYmBvPyjQRHFpc+kLxFvzU6GY/WGHk6O4eNDF2dB23J8XI02FEYPa8vyc1KGKh
Q+HMmZbX2m343AUxAR3B1ArEwDqt3eYp38CYXi55Ftc2jQjcx0N+097dFs9cxNe5jTmqCFXN77kt
ySnvO6+kkM4xu2Zkx+FY7ALcxNr/
`protect end_protected
