��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	���}A�0l�D��9�s��Ž+�K���{��%�s�-J�k��_�	M�X����6�ѽv�eT/M��=�t��3 /���7xӊ�1��أB�c܎�F�Es�i����h���-�ۂ��i5c�7��ӣs,�H4Bu�ޘ|b_c����BFE���!�w[A+�r�b.�)VG܎Z��x�4 4��͟�i���MY�4gϮ�H��RpR������5�M��R�1oJ�(��u���
���I윭ɬ��	��G�?��E�bG��n����/?Z��l_��5�HR��bz.g�txS�V
uh"$�ƒ��u�j�@�\I�Ǚ��'�g���B�M�� �w�+M��9�:䪻I0�)Ơ��Y6H#dnKTS��vڭ<�啌��\�!���q�+|�.*��[ǪaR��{�Ùo~rCpюۖmc&q�O� ��d�Vb�5om��m-c�,�D�'���B����
���X]C��-&�= �Ց>�j	�����5����ſ{���)�޺�n�ͽP�P��(Y��í�34q��%�j���D���i��qx�4$�!"G��V�&���w<��,��$M)�3s�0g����xS�}�m1��`�=����:a_����;�^�OH|��\�Sr�����EYN�nଏ���of�"$�j[���d"��R�%^�02!����Z���G�Ł���d��Zz�~s'x�{/dR�d��ty��ܫ�Ԯ�i^2�ce��h� �
VݾE���̖D� �b���U#���Zn�nH:�	���Aʮ�-[Ε��U.��?_]V��{�~�O�,_'H�o˿�sH�:%�P���ąj�N�����ۀ��1�)=��&6N-�C�h�B0�0VY�[�6w�sZ ����Ԇ��Ɨы��P����sh5�s�j|��=�����RH��׺��"f�:�9��V�g���j�lt��utQ�n���r* _��q��sN�=��vc��c��+M�%\O��s�7ged�������-�����ꃌ�����p�r�,*�@'sW?RM�P��+Fn�9����-�};�Frz�hQ���g���;��N96��7u"��S�]"���)�n+�}�3;}}�9���ڞ�S����&�x��t����j~��'k[W
�(���z\؂ok���-��vN%$���b��\�3C�=<����Z�~�_j�O�,P|����F0e����Z'Lh�f��n��@Cco����:�
�2j"�[���:&��� ��R|���cR�GFT�,\%q���v���8/p@4	ߑ�������m��E���x#�R!N�-#���j�<'�t���z��Gi�ǯ�RǻP~��9/&J)4Bvp
�ڷ�c��6Y��>7�c7�FRz�O�FD���JP�qv�5�D2X���^�f(�V�սU.:��T]�okڬ�W�d)g�?!����>7k�nrF�V�S�����Z�Hʦr��m7����<,V��LY@j_�2�'b���33���vQ�_W�=�&j���>2w�Nw���k��$d���3���R�:����kn�W�)�fEkP��u���y���'������T�|�$?��_��sR)�}�R�Y���c*���<@l�}��՚��.ÿ����d�#���p�P?�0x�D<���DcY�&׶�i_p&|I���s��Mx<�o���^8>�ǁK�!B��rN�4��*�~� ��[��?�����;��4�i���]�wg;�J<8l�i�j��R�/b���]��m̀|9������>"����~z�X��:�Y�����MboL������{Gصt�iJP�,����������i� ����x�F}`󸘣W��H͞���O�:"$�Y|�٧8ŢI2\+�Z��>�2a�;w2�2�)��/�꼈cL	M1(��q�&3!�� �Ħ�IWk�~M��a��>{U�fJe@:��mm��)G<I%y�O��+8��I>�+���i�@�惿5��j���֮(0��u���2�}5``$�P4���f3�љ�\�:��R8R�[4��|�;!�ɬ�p�����]��I{��f�J���_���4��_"�HJ��z��N��M�G����&�0՞8�F�m[>e����⛫d�0���4~馵5���M�9qQm���a���Y��/����~ŻУ�C�<�ţD��2q�Va��:��c��o���rd_�/{��F���7��"��FH��k=����E��u!��7|�S������4��*nc�@�O��A�C�kq�����1ٹI��T���E(�a���9�f>�E�).͏ITպ܏��,�m�F�_|i���C�߄tx�q���'e�?��,�,��v�����^����a��',k��g5a�v Y��Z�s�LqWs7AruS�M��16Xr˝�1��-�&��j������V������pk��NPR���?<����D_����|�[dt���`�+$��lb��-d�v=�̈X�S#�^F��\�xr��7\��b y?�0#X8���]���zH�G�S��{jͤ���1k��$�(�r��5^JC�(B�t�l�vwQ�ȅZV{&v����'�mT?��)7hď<[o,�����H�D��;��#x�S}��*���u�;d:�1���_�hIp� gmP/u�.
����;aHw�`lc��ۖ����7��:�d�'��-��7o��q��M�C)�Ӻ>���6�{�����_�ٳ�3r����,� %���3�tv1��y��6	DgQ�=����K�:�[���§v @i�8A�y&�R���WρJj���6D4��?�f]�bP�'^hM��ۜСыD��B̥���R]I6t�sd{�jçg���6u/.�*��ŠfUh�����<}��\w�� ��|��8w�G�*jK���H��F>� �Xʈ?�nN�,P�l��\�Je���5|�O��,�B<�~��Hh]t�8lH�d�М:��l����e�s/@>F��(P�@�^�>��ض���7�4LR�K
�@ŰlRy7��e�+�C���qf(�~�II�p$���VX�rc ʂ������#6�tޕ�W|�.�a�Y��}�M��3`��@F���?���w�}�䌍����1�����~Ew�������D&���}S<��,!�9��y* $ PX�M���.�������!#�{����b;�8C�we�aΩ�$׾ފ(0"��D���*C�����ٿ?q��!��d���%^/(�����!�t�	� d=���&�P��0��N�b�t;�����(y��*�;�{,�N
j|����aco�Ay�Y�q>]ͳ;��ζe[d�e9Q�K�S���$��5����QG�2�Id��g����91na�����✑'�P)�=Sa��+c[��TyU&G��z/ojlu��	�҄����M��#KS�9�1�w�r=��
z"��t
jǋ�df&n�j��>���D�C���s��w\|O&�T�oCY^�~��+�(ԃ;��B��G
B�|�	Qc F�	n�mug�vY!]�F�_M�ʝ����38D�cs|�x|�	>�U�"����S���.y'�	�t���K��`P�Ϙ-������ܕ^�U���&���;_��;���7=�����9Z%��\q��԰�KK����	*�A~Q�{5;T0���<�lH^r8�Gl>ڏE ��ץNYiy+D�Dy.�/�<�C@<�1���uv\m	�_QUg�z6�������s�Ꙙ��V�œ��XQ�E�C�s2��.*��r��7�B7R��6�|x��Q��<��I,n�'�]r�OS�`�*�O��Y�Z\�)�ͨ�����(.��wBKD����=��F>�A�ξ�~ҋ7:�v ���/k�R����T+G_�@�jpe7O��.<ABW�8���(a÷�e�0A�鏻� ��p��ē���$�W�1���iA�?8$�ȇ�iP��|���)�V��W�LT�"�iZ=`�a���^���A(�W_0)���$<�\�?�?��[zB6�7*�ƮG#;��46� 5sA��C�1��ϯ[�R�YVභ<A/�뎡�ϊ!�q�w/o�p���Jsթ�}�낸N%u8�wJ��%���>	��
�-�vmHٕNL�RfX�oY��,������/�K��/9S#f�Cc�g2!�Q)]G#6�"j��J��6S����^�yɍ�ON����`��V���t+�[L'̘r�C-N���E/\���*�BЈ����|��MEG��hX�t�7ǖc�=[+�o��,����(s��5�����d���(�a�}nОj�T9��K��l���yJ�{}�YƼ@���,�raC:�:�1!.v-TFCc��Q����_#�8�?� ��Ȧ�QB@i;I#�8�LQ�>�s�8O�G�<\�w	d�W�/9RN�WpC�V�3Uzɬ;/ȴ;�	����0`Bn��*�v"��^�r��n�}m�_fԇ�>���d�bȫ����<Q�T�ǳ0)މd�$:!�Σ�uDE���Wwk���F��mu�bھ"��[�5���.;����*�Ɲ��+(������&~9
]���:?��ܠ���W�u�߀�����?P�h����p�MB�M�>��-�i�(���^��=<������)�}��F?T࠶�r�5lj�~�s�+��q
�0�]\Wﲟ2�L��x��S�U{�l·P�QM"�t<z�d�������
-�<7�vV�Z�NԷ�c�զ��6�.�`������iXK�fb9��e�L�7k3��*گǨ2;����(���5��Q����!�`����jn)��Kry�R�Sv�j&�ľ��Kj���
�i9����ꪭ�z�R��|T�O_p���r���B��o�s�G"k��o�mZ#۷�D����w�͠T�'�Y�B���Z�7����Օ¶݅�����,�;>:T�iΞmy��X%6�V{UG����j�߁E�m��Rõ=GS#n
&��#y��3̥�����A� ��� �_���LG?<����y{�e���3��ig_Z�j�2Q/��˿�����4]i&��4�+��m���J�r�%��Řx���T����e���e�i?�F2qCW쉭�s�K��!>�L�1K=������T1tۜ_��&�P���w�5\������0�P��]T��y@�լq$U�ѐ,z�0�E�Т��\�|�ϡ�xǹ����?�w�@x�vq|^�}r���+ܾ�ֵ]��"I\_��mB��I�<��N���쁴~��Ƥ�RpTYN#Ə�
�����D$(�����͸�[8�)�����eR�/6#.�'�iM�u���wR�8�@��5�'����*�VЄ���'�W6b��\)7�e��t�ƋE<��p=��1��%+��HC��}�
3��P�%��������%Ӭ܄�.z�p�Qß�d+��#9���i)���4�<V)����ktB���{������qI�T��+Vs����[�xt�G�la�/�?�j��6g_l�uŏ�f2J�Z��O9{��#���r-2U�[������J$�g �O�D<���F�����h�-�c�Yp���J��GV��
v�[��g�2"���{��bx>�����3\k��/C[c�>�q�b������vR��n�s�Vw� ��m���D,@�8|RA��es�B�R� �I�F,�Ξ�Wjd����夐(l��W�o�A��m��L�x��uҏ d#��)ȉ��8=_w�#Nh��
��~��*���:P@���O�"�[�x;)�Hh�u",x	#�5�+�H�r�!�Gk�=��������g(z���c;_�U�pQ�@���:��5s�YJi~�
�lw��w���8'H�����~�@E������M��G��LZWP�Al��a�P0PJ@y��0	>��Z8�.#[����.��t��3nT�^JS�Β��)�w��^�0�-�9�H�q5;?+�:\���5��U��_{<Ǡ�E��y#dc��8h����p�c�p�)Q =����]����0�~�Ȝ 0RP�����n�{1e ���|i���!�/��f�}Z�qDo�U�!x��İ�B�p�=Z<���/����$�^�+��pD������R���Yo%�o�{n��� �\���H��Ň�װ�F��0���;Tx�LsE. H/�A�z!��gD��ql�:c�oeh���R�k���Km/��F�ϚM��U (=�@�*�]��G����C�(����M��|�׀C�:\�-��왧�^J
�a�ݙKinz�l�YX�^OJ F0Y�OYxM��#DOm��{��m¿E��{S�ʑ}�A���9��1Ms�6=��$P��=��/�쬂�b�K��Ut̄������)C�');!��fcB�����&���>9p�׍~�Ր�-��i�R�I[�eO��] ۼ�#lϥ�,����.���څ�,-�W:?P�\D||�U�dVYV�L�q��li�v���2�I���@LJ�׭����wl��Iُ�����%(�+m���s����!o,�t��D*���Oe��L�o�R�YN����?��Ĺ��}�%��L��Jq�x��v��R��i#^p��)����j�$A��ŸU�3D*��N�9�+x�3�"B�:�6��Θ��k�:�7'��p��g���l�G��J�ӫ�s��CdZƕ���5=���j�v���/L�F�wvն���a:�8P��(C�:�a.�������fR���ˇq����Ev� �3���|~F����Q�\��}�H�G���7\��������0��#�њ�9��>=��$����Ž~).���&ה$~�|�	H���w��TEN��OO9T�ӄe���<3.�~U���v��6u��"�����u���m���L1�3]��:]�K�g�lM
���˫�&s.gj@�Z���
{J"/����PN��І*�=<&������:��S�3/UC������p�DQX�N�/a��R�l\2:�q��ޫ�����>��i��-���Ċ��=R<mӪ/n���D��*+��Y�a�]����<�G�~�~���7�"�����&Le͘�=L_�u�S�GqAQ�Ĝ%��
Op��U9���RH��B�d�o)��>�ukP�AD���h"kknл���!�G@��fXR`҄����<k����jF��<�cщ�ڪʹ���@�����;%����I��<O3���W�}���N0`���I��(R��n�O&����-̢H�����k�پ�z�gb��[���o��i����Y��lN巵#�{us54�WMy~����E{����4U^�������
H)�%k8���w1�ˌ{_97Za)��o�1T5���80FU	u�=m����MM��9��8�;�o���R'́
oTh8]&���Z��-p���/����)�L�P�B�,��Z3
��䊚��6���)��vDo��l�`�"+� ֮�t� ����;D`�q� ���=�f��L��R���o��yi�s�`�q������[�ß�9V�.�W���,,G4Q0��U�*[�:^��H��}�t��<�"��wab��TQK����߾ꢑ=��Y��q��M����ZM�2N#��#�葫;Oo=�F/��������1Wy)����|���Yp��&��S��r���^{L֙d�L�+3q��ղ ������-��@A�N^�Hݻz���
Թ���(��T�ƭ�f���n�mw>Yi�Ɏ ]qZ�Y�+���U�2�yj�(S.� ��A9:�V�?Wӳ n�������B��~n���ɄW��LFﭥ4�14{���l�&���tz]�@�h��q����3�)�N���o,����$3��im0��?��ǎ��U^K���־�TR�~�i�p�^���[4��U�+��r+�>�&�u�hҎB��M�K����4$&��W'��1FwY�hA�P����������}dˣ\���u
H�+-=�Q��7����r)K@�T[�j��N����C�@q��3-ԉ՝��BE[f�)=�Se\Ek�a����k�/�-��a�+�^��B�\�2ٶ����5��>��p4�an1N�>�]�����|O�Fk�}�2�8��ޱ@`B�0�>�b�lr��&x��R�a�A��;���}P���g��\[U��%�|=���M�㰙Hvp��ռJ\����IL���w���K�N�A\�A��v'n�C)I�t��H��G��S!x�v�\JP^KՍ�m<�Y H�.?4T�G}�3�tr:�P��� t���4l?�	=g�����3N+����<i
b����I�#B|�#��ĥW��٠���>�@��̧V	��������V.��Aۂwz�Թ��wE�Ds�l�;g�ڦ� fw��,���V���o�O3�s3,��Ƶ�˰��K%U�D�"K��	����3�-Gd����z���E���cߩ�!i���%ug��o���C� ���q��H�
��h���js��z 7:A#s���SMu�9��{$�6�*���������/|X��ϓ����$��[��5��E�c,��n��LА*2V��NQr:�B�I%��}Ýl�����n{���(��D��;��c�sniv^�w����k�d�
��c����7S11м�Q��K� " sa^Y���l��.��l��\,�?��?�0�5+o�B�G��� c��^7a�O.%S��y�T���Mh��M�Z5�r�zS����0�a�:�Oe�A���F�c���|�<��-{��+�!K-`v���I3�2�$�G��[��pI�4H�ҌXV�=�7�}1��v��p<��Qn�か�^����+�[��Whщku��ͽ�E�A�xm��MF�U�<�M��.�]p��c�ŀ)�1B���1�hp0��|��jxtx�ٚ��R;N�t��o���A�B�P����E�z��뿑	}}=�N�"?o���{.~�I����&k�bƊ'|�y J��D�tlG9e���I��҈�c�ݝ^�ؘ�0��ɝp��Hh�ƙ8���Ǧs��Yx�+5"�0���A%�B���Ng�\}ܲ����}y�iN�P�"��73~��F�dqu"�_դgjZk��Y�2����9��pM�{?����������O�{>��qȠ�ό���S��mΚ�y_����oo6ǣ�$IMA��F��
/#5�hW�
9���M�Hy�S=$\�V�b����Vk�I.�"	��;D�U�� �sU��h���u$�(�0eFr�A�@��6���;C3���;hq8y�R�-���/�4���M�/>*�K}�XY�n�tR`n�'�F�'p����у��e���G���I�Ǌ�P_Bg�&WT)T�︗�H�ڍ+<���L��R���]�at����pd*#􋆁�����{_k��ئ��Tƪ:�o�!����F㐴�z�䥴���-�Tg�?ɖ/A/�׽���J%�)+ �X�[d}��lj�����+�?�����\;�v;!A��z^������*.�Ԃ���4�����P�G"_�q;|ixx���j��1$y`e1��r^c4�а�e���zv�hL�b#�<�I"8�u���̢��gﻬ*����i}�����`��]!�eK��q�6���%�_J�f��UK�� �����o��q����( ����o3��6��-m�΄\<P"e��b9a�p&��K~��';ۏ8;c.x-y+��}�ƨ�O]v7�O��&�Ⱦ���:��"0_��+S�� �e&X�$��h���=�}������{��b[���X]A�<+\��Rj����I��E�n����Q�O��څl/��t.���iTҗ�{��S�W�N#A�j������F�޿���5�������Q)�6���i$�.=�Ү44��7F�6�R�Q���Z� [���$M��yj�+0���ݯ ����7!��|�Z`/�w��7/,�=�>�*R��S�S%���5*^u���B��I�"�����6�O�*ї�[��!�k������t저�� x����8IPp_����3��D�fꛐ��2�3GB�F�7A}n�ߟ"�����Y�>�S��g9l�&��a��	��$�7s�G���Z�.n�&�b;��5	
eT��Ea�A&;��K�7�=�q1����˓�Ж2P-�����Ĩ�HxP�v�L�@�@�:#�[y��6��A,�ۅHb>��R��48*t��-�gԥYc��bG�ol[o�!:�dHk��Z==n�
J���2K^^R���