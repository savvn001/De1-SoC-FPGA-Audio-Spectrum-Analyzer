��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s6�\uz� ����ۻ�TΤ��p��G%*9O'X#pJP�n==�=�B��=F1�?X�+�1�d'�6灨�Wg��Z�/�k��(�Ѐ6I���� �=<��&_FL6�[��q��O:
�<�k�]�ή0�D���ɂ&j*���C���?)@���+���K:��/dBNz��/��Z��-L�.�Ux'�6o����3p��-�w���M��`WN��'��0� .w�
����ʄ}�\�����ROR�ņr����ǚ:$����l���O��w�_x��fC,D� ;��ͬ���6ΰ���8<�0�-_mGB���:�M
���+?	�PZ���x�Ε�)c��R�+ꊩ D����u�jTg�
��p�Fc���dK���e% ��C%��<�V�+=���@�єF�.�>�i��=s��G�R���%���i�N	���@�"�}p��d9�i��:H���:���#q⒦؟ �Թ�+f�����\t��e��|2/�k�
���}	���a�����c��qN�(����wWV&�ጋ��N;���/�3��v�@��"�y&�*�H�S&�a��=�Ưs���2=_>�]���џ�._{�4b�w)808�A[�)E�DF��r�xwY�* �df�2�	�Jq�VCyQ�67�P����^�g����}�Z��AT:�k����qҾ��� h����BP����[��������T��hXj�Ry$%_3F��V%9�\��h��As��u�#� F��@�l��}�|�Z����Ï5�Ri��(�/ּM�~������3�"�׬����c���X}������<劑�@]T��z[���˚Mt�P����<��l?}�V t�?z\���Y�!�#�|��F)� ����Uy8��&�B�o
�ɜ�Y�,�� �"�.�U�In����{�����Q~�+Q�Bl���A��}7�.�?�
��џt�a>S���b���Q9'>jL�O\3��w�a,*Ru�v�г!�,]f$T�s[�A	��92H[�.Q�T4և$���X<���kY�bP�w@yS�w�dk�>2��+�=���ސZ���c�������`۪������4/W�|H�cE�=V5�]��>��b%�Ά�M��}��ʰi����Z�(z��~�E�"�\��S��/	WPKuÆ�1[�/�T*=>Ժ��a��U�W�@�.�	{�!�����?����W�z�� ֕1�C���0�{	D���j;�(*Y��L�k��$�Y���\W�8�F#�׸m?5��P��]TJ�7N�
�K�"�p���'=r�n���,܋�4�h�'""�C�Y�j�f����}N�c<ۛ�ܧ����!�u���b����Kud�D\�2\�ۇ$-���||��� !���h��n�%���O��s��	L��`&ٜw�)���M0vw�4��"�.�(L��^d�q��з���Kq�����_�w�)�_�'ď<Pҍ���U���L Юˣ�c42eG�n>��Px��]�pt	��9����"�9EXZ6���d�Me�Ҁ�v��?k��Qn�Wﺬa;Q8%3�?�W�@;�k� ;?� �2�=�n���]-���˯������ک	�&8��Y$�.p8������Z@^X"�s��W��%���,�]�.���b]��Ҫ���a�NW���w��d��7�=h>P�zb5ش�*��L����c�݆.��?4d׭���������-Ug �28P����M�o9��V:�B�=���CES�x�x�N�_I��]]�3�A��|?Eb͈E(��$�A�3��G��a�%��}S?k��gY�?cPe��Q����9������y�9~E��c�O��V��/:|�߼VR��F�P��6b�����z'��g0b�����Y}��Z`�8L]��{{�p� 1���8O��[T�m܈sQ���w��*|�� v~��������j���)��H}>�'�l|���]�%ˬ�5�Y�l��d����Q/��+Ȍ北R����㺺7��ć��� D)i�����`~�BtFwB�ηu9]�_�T��n���X�����R�Pj��m�� ʿ����}u%��k0��u�?"�.3*]į��ǓC��Q��uY����hE< �ѩ�1��>"�r�5���&G�������@<��r����X�����g�F�����G�����Fq<�����=�Y~
�"эR�������[)n��km�_��o�ב�X���(-;��>�`��k�O���wi�0��D)��`b�a��� B�� �&O"~����=* �?B�ލ����o"0�w�(K'i��7T���	y:�5H�;|���;1�1��0����q�V�d�����=#xT�2X\����U;:y�Vj��p1��_�pF�=N�<���g���|a�R~�B��~۽B�?����˻0�-�67�v�[G�u���:�����8��b��8*\f�2����$h��vx|�x�w��3|�e�9u=�бX<-+Tpۙ �[X5�/�'1d��X��S)����StS]�)���ݫ�Y��:�����Ј�Cd�l�}2@�gRQ�U?4�����eZ���D&3j�RrLW��g侫�t���0zC�pQ��	�z8�V����W��d? ?��)������\�8�	��H%V0a@P�q��|���'2�Y?�C���e춭�?1O_T�f�@ul$%g2'��ο�/k眵	7��(�j�%^>'��Ou^�30D>��q�Q���%)e��-b�Z{�Nێ���y]c�F�R��Kx�!c�Zg9�#��m�ى$���.�â^m�����P�L�Á7Y�K�s<�B����zz�d/ԘX~���{(����i%�Q���p�2P�[	�ihBp4�s��*�sKZl% �@���%�e%&ʘ5q8
��81����׏�E
��E�rnޣ�_�d����O�
�tx.�[)Ni�K��Y�co�+\�7�sTʻ>�`���v��;���l�ҹ�e���y���� �*i=< ��1����c��R�k�WY R��@���WU��X����aK�����U��	)ph��iiɤ��P�Q�Ō@ˆؚK"��#<�ۄ]�%�"5��M�z�)S7�DH%U���a]	���H�E��w?��*�mA �i�>�yV�v�i�s��m����F�ed���N%���U�f[�5s��W��ᙘyWYc�qr������yg�ٮ�R8-���zh���<��2|"Ѣ^��?dZ����W��,Z�Y�D`�ʓ0��7�f�'������m�1ѱ!���࿍��3��=pV�����T f�zN���cif�`s&�o�vB[����) VG*���)�x�{ɫ@�VS&�tX%Pb���H�3�|U3� ��M��k�&S��Y�cj���n\��W��L%庱�+ �Z5�;�
p���hn�qE�ӥ	���M�q�H���=���`� U�D'�c��Co�G�:MTU����p��@��=lh �$���w��O��k&��:f3���B-�XPU��P�5��Z=s��e,��iHv;T�-M��[�Ⱥ;R̯���[�(�`��,zFA���z-�ML�	)+�,C;Ie�pO��"���=��[2}3�u�J�R�A�e;�LA��rU�8��l�1o�c�-]��L�]+o��Y����y�Vi������uÊpJ�B=0�A�䝻�x]O����|��	���^9����8=��J��5�BA�uIIKh�c��J�R��e�O�W31 7�2�-�P?�}m�Cadб�Y�! }|�C��ty�XAw�V;WZ�M�H�T�0h�ւ��\�S~��-`b��
"�P�+��ۆ$�5@D��,��;��ڍ$�����˝r-Op� @�k��tw��1�Q�8�I�`OtЀPտV��Vŷ�*f�]��-c5��f序��߂ȡ(�6���"`P5��R�te�Jz�rC���?��7�g<���_.��Ո�{F�>v��?��A��sSQ�f�h6.GU���pe�]�w�)R[������m���"'���0������j
���,\O@ߣ�j�2[����Ch�М2:0�ƴ-�%�::��3k�� �+9\�=���+p����
ԇ�+0Oq@�����Z^90�"+ɓ&�:��}����d��$W�g4�h�D2n�n(J��8�!	\�iy;J~N]r��h�Ry��将�d��1V��&>��f�Zr��(�@3��#ψ�+����	J(�d�3�z-p�0=,���R�66���Fǽ[P����1t4x�<����ա��Y�h������S=��eX��?s��H�K��R��zw䨑]˦@�t��fs��VӒKV.Fw��[�χ�tpT�R��yo��Q�/m[Z(���U��d(�w�^!S��EħYn�}J{x�K*d�H���w[�b�(=��~:��܌X����`����� eh�S�5���M�{�Z�Ǔ�["$.�8Sn"Z_�{q��i�n����g
%��H�V�x���R�V��Ո�IT��g�\|;E�p�)S�q�8�@���4�s�lo0�>�#S�4���;F>�g:0� ��G�9�O0��8Z�p	�l�	++�~��
�Xꅈ��	x-��*K�K��rxX@gv����Z)��ۗ�u�j5�8�ųJS��!)�����3�ο�HK�>�-P)-��t!�wk��)�V��ȴZ<��q�q����*ݝ9��u�!�MM��Ӧ�f���?A�/A�� bk	��R��bߠ����N���h�gd�K���	��-f��uq;|�I��O���&H�ĩUZ�7Hw��mdY(���}J�IG�ᾶ>�̒���B4�(^C]B'_ޒ�|��׍��+�M��YB�w�MBy�?*�&\
�W7C,u�`y����[�|���4��Q��_�b��7���U�\��y$�,�>�H;Yi2�5du�"����E����lժ���P��兖|�C���%,�k���囮������h����cSA5��=�2���MB��o�2U	̕����37M�5k藫��ZΨ}ϻ(�(�k�r<RD���,�2�����\�9d�(�\���_�FN���!�<� �,�����#>�b�BJ�13f�n=�\D��}�gɟ�Bh���1O�own��y��(�;y��O[1ɕ�����o��������T֮�ф}Y5l5�/X�����.VKI��L�{�ɂ;]�uw�%i}x)>���t�'�= ��i�f����>?rL�}�46"L%��i◀H�Bd��z\�F%oaS�E��L���L��{.�,l�1�|�`nnW��`cB��m!��Q��߯� ܘ�_|<�3�HL#��o�EA��"?=��XW�6����c�Dc�M��օ�J|&��''@�t��V���lyoL_��5�n�KZ�`.8v؅�F�7��<ى[T�a&
~�S�)O�-.��� !gX�XZw�}��
���@��;�˽��Ԇ^#٧qw�>v���ˀg��_�����Lo�й7�P9�R���>Qd@ʺ�f���U�i�ֺ����L �35�md�<z���	,�];��%[��0�N~������ɻ"ï%�׭1ڠ�қo���sF�e�o�� ��������H��R�	uS��b*�hPY�т�[#�ԆL��s��n*Uh$�B/V�'�P��Iq-轉��fP�dF�؆U�p� ���r�Tx>��#2� ��"n*�w��!2�6b�`��e�&^��'�m��,���Ł����q��b߸������;z�ew.��*a}侬��
,w+�Й��Yr�dM3�m-^�_���cQ����6�>N����$�A��Ι)Hgcڌ#=Nim��QK�N�:���m�У�U�ٹ�&���O��V]��ʇm�Uپ����I�N�ֽ_:X���p�S���vD�������Ǳ���ր�W�ۤ*��F��Q���"�s<��]+��~0�"1�2��)[ɀ�Y�3AػAp+(l�����^�<�Z����1�� �d�W��
cs`��er��n�7!tYtl��vw�aK߉�,ϭd΍-�5��ԅ�u�eI�sM H�9����	���@�Ѷu^�~�֍:K�8-Jர]&����2��n{�eV��㍈�G��kG�(��p/�K��ǌ��{��R�r^�㠾�}��ϟ�h�]�%C2���.��%g$;|B�־��2>����'���\J�`��cl�Et�2D����!��(@} ]:m=�=v#rB�fXo��G�Ry���:m�4����.�����7�<p\�|���ϔTv����-��b� ��-ٙ9�^�����N% �]�����g�XM��=��S�b*�(� I���:ǀ���zX�s���`���?7��*�Y%����L������y�6�{l�o8LV��L� Q4Wob���䩯�\?�E��P�u�Fo@L��l��	\{�W��vҍ|����֖�h��{�D�W��a �thR��rW�:�BD���c��mr�A�t��4����^�H�2�9.��!��2������e���寄}4x����뱎?c���6���dv�wPf�D�ޚ���̬u}h���:,�)�I��z�ґsmk��g�:7l�/<w�4e:90��'G��4��
����;\wב|�/1����j��9�BD��L� (L��T�����kY��������T`;��ʃqDa���9w'4�E��G��7�>�wb��1o�b�B�`ݕٜs�,���'k�[v��i!��6��5���P�c�׉I$���E4�������%��f�W$�~GFѼ�%p�	i̒/J���9� �~jC�N3�ef��K���C��R�C��z�m:���9�FDwp����V�)���d+�d3�R'�^�AT�����&ī����Px�hW��C����찿,����?÷~��u4��&�{GxSFLՃr���U� 3�680ߨ�|�P6v
`A|4�^Xqܝ���b��-RO�+�MR�D�8疆��=�̓��g#Ʃ����R�� ���˥��9t�E�X}KM�}�6R~�k���Sɫ"�{ ��Ă�7[�n�9�O)�Z�����g��G_<$��aֱ�:X;aQK����Ü��7�V�\��[͸f����/%�nb�Z)�v�c��?&Z'P����ȓ�KM��l��swc�~��@�bxF�Br`֛Ǵ�����N����ETϻ��kI�o�\b�5C!�j�|H:KĩU������=t��uν|�c����$'k�7�&���hֱ]:s�BD�^��Y
H�\�Q��w��� ��
�H�v��ݤ8 %��S��`ås3��:u�u1"O�<�R-� E�%Q��:c0�x��S>w�Zm�N|���&0��ύ�s�> �Y�t+ �J�-�5N򼏨��_