��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	5
����a�`���~X���!�>=���(M�+�#�	QQ�-Cϸ�����Wl��L���3�)�^�pI�2��x�Ĕ�[	���<�f�7�uM*7���Y��{�h�_UP(k������<����$�ɭ��|3C+U�#��r��>2UH�-6�^��W���^����S�����T"���k��X���L૥�����C,�J�y�c׏�J(?�:@��w��ΐ�U�!��9�Pz��|�4=���R1C�ܽ!3Y��&�.~P�L��[G*t�ؑ�-Z8�bmП-_$a�Gֵ�c 5Yݚ�Y{C��+%�f��2ĦaP�)W�P%pxa'>T�jp~��m���󋥬L­l�~-�;�8`)%�Ŭ�/MT����iX9��I����� �e��9�p��I�VG"��!ʱ���PTm� I
IɽCbF:�Ș٣���Dhp��3�x" 黯�3zV�ȢoO��Ԡ��U�
G#FRDC��]��:��՜�y����(F����L	:�a�|if�J�>�Šˤ�F�~��B��Q́���W�}6
�uUSD��ߜ,��ף%��y|]g��j���~g� ����aM����۶ ���[�t@�4{�(�2s��,f�C����ދ��u<�D��u����Gu���ю�e�2"q+NyY�b���?���N��?P��0p7�#wѮ�kθe�SőS��18�Ӵt_���=sh�VVlP�������[|݁C�}EB�&��O0Q����:����+�N@��EB��<�xVC����C�"Л,�M�@�ՔQ�\
P���~T���0Ӻ����Iy�Ϡ]NE~~����%_�=&���ܒfGoҶ7P��ZR���
���9t����v�I|
�8��09(..`T���$�>�k�2C	Կ:AV��`h�P�ײ�[n-���/�6Y�ɧ��M�GIU��A�D;��#HkL;�A���S.��`Vr���4N��<ppJ��������J���jG�EN�e�T��d�v��"��5�E
EY�v�vA�eo�T�o�>�Z-E�2D��#AL��D��B�@}��!����)�{�2��ݶ�0��j^;���q�Ƨ�o��/������BR�4:�cD{M.fEhy������d�I?���lN|��׶v�&��8k�.����`�r)��f=p.B��JX~jَ3:�O_1"tN�/�/y(p��:ĺ��:��mɍt�aA�ݥ�b�}�f����	�V,WlVÑ	x�D���JCE&Rjx.G Na�`	�c��<W��삖
g
h����x��/��*�D*���b<��~/�O�.Դ�a��l������4������k���޵ם�J�k�;(B??��L�V�� u�bd����o^	.1�	|�ݾ�����ᒖr/�:�1_�����Id�F�	1�`����=u�l�Շl�M�nh}����5�;����n#<�}�u]�h HT���t��`&�q"�.*U��vж�o���v��]un���%s�f^Uy��*�C6
��W/�?�>[�Gb���`|)V�R@�_Я��\�^�䪪�UD�0��zR/�)�Cw��]�d^�M�f*�i[�qW��l)u��y7M9*�����*�}Y �c���4k�kyh���Օ~
��w��Ń���Cs��b��̴,�\o��td��Z7]�͊XEq^2�P �R�/h;�]?!|��_Xzrb�>����1H٦2��j�Br�EHW�/�#�&��M^J౨�Z_�@��O1�&'&NטC��G��~�k�6�)�T������F@��m�t'�~Ŷ^y,��%1wX]�f��&�8��Zt���[Q��|S:�&s���[d�&��%�\�A��w�^�@Τ+o�\���X�p�J@!�oq���˽����'�o�i�>�W��C�Ej01&Q:h����l/����A��]:��mL�ׅ37���p�}�y�0�X`�`i4,/`���4Z.����#���7�9k����'YS����>��\�STI���ޣ�\+���������L��}l5�,�� �e�T���Kl�k����� j]�&�f�t���\�CxhUb�w
@d9�D��T���� rs^������u�u�i�������`�;�e^�1i�MD�h�})$�Y	�g:aK�^"W}_�RL�˲�&�Q�)�u-�=���'�T�h�l������l�KI��w�p�\z�����n��%��`4�Sgg�ʹG�+G�}Ӆ<'�n��T2;ʌu_�O��y������_O����X̭�4|�MÇ%Li��\�(���+�Q�7[��u'd��$o}}}�A��[)w���\��k24=��q��d��#�]�sGk*=l������U���U�lA9\JeIk7W����9�A�d%:�n��6j���0�x���UF��9|g�Ч��(떇��w�͉9D��v��%��w�թ$٩���Uy5�q˫2Yiea�+.�'#��j�J�l"Tc�A8u�2n��OU�8P|����6����Y=�Y�Ē�����`�i�۳�]�]�<�#B����,��vx�]��+m_7�4����
����$��KChoFfE��ޏ�]��ə����J:з��l"@��$ٕӫ�"bd��������&q�g�F�kJ�!3ti�BW�qK.1��QcM��szRR$����IVI��6��>Ȃ�f\��14W��c�a��5�T����Q��t���_�C ���j����7(�jFh����F�ak�3_��'f�븞�kJ0�H�
���E�Zj@9�0g�-:y�������3�s�v�c�V� =��y���M~��&����p����A���P��3����c�sl�ǻaQ�EXW9��.c�E�MU�1�{��X�	/�w���N��&�B���4|�z�w�y��� U��^���0׍���k|I�'�nȾ,�d{1�<�PwL�+�'���8li������m�����o�V�M�{DW;�;�V�"��k	09 L�#�u߈�g���p�4�D�$�_��l�[Cܥ7�̥l�i,~ѷ���!M$��#s�}f���olY��	� �I������'X����kޤ��.�B�G��(Wg Դ"�M�u��������@�LL�q"'F�{ �ic��Na���| `��U�v�![�z��p!�����Uș3����*�Gg�@�L�Ki��]tv�8�\�^�����rX*��f�.��[W��Y�!�u���"(IBd�/|hk�\�`�&���b<�������3��s����pW}���>��9�|,�Sؿx�{j��1�J8��m�1�vB��WkD����4,�-��q�G�B�ܑ�B�9�����XM��ͭ�/�l�D����������2kJ�P��X�5��b|�4i��	}W�6��ɽ�k�����M�"�ì��)כ"(�� Ƈ�1H�4��>�+
~�3���Ě�������RS,3���5w�����Rˍh~�A�
~���@*~@�y7�EV@���0�t����0Bȳ��?��$~!i��6�]>`4D���)���ߐĄZB8�ߌk�(��[����03�+�s�m-T���[!������A.{����Zk�����}��J�gv&�t�^[����5q����XP�'?���)5��ޓ	G���|F�rZס*�9nӷ�	�vm��ٷNW[R�(>֏���MF�[���������l�u���c���|
�x6�� o(���\9���Gφ�O�T��)E%�6����%�xπ�Nbݽ�S?��&��O��A�b�INi3���}�k�O.�5;pz�wwK&X���� �Hؐ�^/(��i��yHN�o���K�_ѓl��|H\�H2^de"�C��`��ϭ/�=��)�<?�M��A���F�}��sZ@y���$"��b�K޸�Xk$��i�J[qO�'��;? ���-�:� �_�i�S0�*6��2��}��fҔ��_�%9�r��H�Ֆ��Q�e�L�e��}��7���V���j��i�x�g-��Y(�Ϋ�^��k:�}�P&g3��^x�2�ge�\�5��M7�4S �按g
��I�e�{�!5����e�d�7w�(N��/�n
}�1O��v�:�^6�V;��h�a1�j������v��d´r{?�\�v�T�z�og�T��HsFMm��~���������q�����7�q�h%�.9J��Һ����P/#/
�ӽ:��٧3��C�m�V��t,'��8���~����
�@A��Kx�s;�Qidǵd��	�!b�|#�.�G.ˈl�佣>�=�:�g�i�8�n~���� �5
��US60,���ĻU��܂p���)u^�yS���bT��yE#�ا�FL���w>E�s�w���{8�KK`T��-� �7�a{?����b� ?��&Y^5Ԟl~��Bg��%Rz���m��m�Z�'����f���s�K��O�T2��-�7/b�-{� Rbl�I��m��a�7�琇)����cp��+����^E�܇���e��1�k<~g��e��9c"2qsޮ}�����?�� ��2���tE'�v��="�Ȇ�!=H�-o���C�(�e�.3�H������q�m�*�>���GF6%/��u��t_�zjV����9�W�ǆ�h6�L�G�n-[��7-vu�1V���l1��L8.!�ȇ�4����2ƗEv�m�ʮ����E�К�@7�(I�p��j����.D��M�Ԭ��܂�s���w�c�Λ)�� 	���H[�[<���Zή��ޜ����O��Q��|O��Q B'��(Y/��8��um@���C7W�?�kr��Ai]��q�ʦ�%f  ��\'�K��:��t�sE=���X`�1�0��E��g���pP��\;):��d���wHY���&#�D���r�����EC�׹��5M�����9L���m���s9�I�E�4��Ѳ�InY��񄧀��X�`"��A�ix�����^��'��;t[�-���,�����P��b��wu#�5W�CC�}?���JϽ�m��҉�)1�K�#;������K������
Q��R.�"PSqhA��xD������rjBt���Cck>������!���s���N2��C�op�ʃ��[�4���V��]��̱R� o�^��[����������F�zą�]i��ﰈ އ�����֩T�T��� �u�	|�W8����$����q;'���oUO>�Mn:n��Q5�!�\���bP�"��U8�7�Gر�*,�Y�0�G�V�8�H����앀c�F<h��+�.�_o �qM��]x� Jm��k7e��U���y�D#�a���02�����G� ��Ez�4�`�����%�e��|���(�4v*r�p�7"�OWq����8��s�=�T%e���+�Ǻ2#9%]�m��/^8�|�12�V7����M���Xî�ªv�����D����O�8Zv�����D_7@��51����5��ݼ���6^iۆPI ��I쟧YX��=���\MT���3�ۦ�jfˤЬ� �� �C���_�=�I��e;��;pm���M{9�`���v�]'V.@u�jLor���V#g:�Ո �?�.���v�o?T��V��6��I�,�u����ۍ3�>��	�kG��_��l�Ύ���죊,���b��	�k;��u�]tϵ����B�n��9���EP`w�3��x*���>����=z�y`%dWPX �_����-����-D	��}??��H����g�ڵ�)�]Ak��@�X��%�4�G����KR7U�z��)�g�`i�6�@ƕԵ��ۧX�(�I�zO"�B$�u���yBy{��/ҧT�$k�ȇ������!���������e��L�\��̦�����\�"���S�j���ӿlsL!L�Har�toiu����h.
�^�])���n5hcY�H��}"f0���Y�2�߽U<�=�Վ<1#Z0���9��l�e�C���C�!n߲��ي�v��.�M:f�~�'�
Â_w��n�q��Deo oC�G?�� �t*��>��W��ekp~'�ɱO�tR��	A7��8e9�e�i9%~��ΰ��`��L�o�B;l��s��c/I��L�?��|ԉ�5u��Yt�~��,�!5Jv�pU!+�'+����rSF��j=檟���K�qP08X�S�וf�e�(p��pȐ�_}�A#�iX���[�3eQʋ�j�F|ϵ�quF·�����AW����Wb�f�0�j)(�C�w��)��d��}��Yw����%vo��ޚ���)��ù�Ā�r<��=fo�qh-:�����Y�S0}�����)���y���Z3�ϰ���h�:���������͜B37ֹ�֒#@�}ǭ�y�.1�p�]�$���Ip���ӄ��~ �˕ʜ�t���.�
(+��W	
�����ȁ�m�p��>B�N�3a��Gʦ����վ	�fI�'��X�Z�oD��������gb7��y��كe��.= %�8���k?�<��!����J����]X�N���ҹ�٠<�i~���A�f!'ʰ��ᜏ�h�#p�vNd#7��m�#����&o��ݻ֕g0��>��i��~���Q���y3�D�V�!�z�X��2��?�I:n5l@��FȠA �>x���Ö:=H�)Av����#XBࣁd��l"��TMQ��S'�ВF��v�ۤ�E)@V�E��Y�� ��gZ�Su�h��G+�1m5��63��ٖ��2C`�ܲ}�IE�4�vT���p�i[m�#�Z�־i�li�)?]���EoW�Zګܮщ΃��eR���y3�	�3���E�͸QX]������@GUkߨUIʊ��X1
i��[DU�'M�t��!2 ö��Ϲ䰈�
d&�$�qpz��n�Z�����(��V��K�v������[�@%�Q��J)0l�#�WOP�y�#��&d�M�o��p�$�"�K��`�0*;�9j����d�*�y����C)��ѧ<aX�p����ܟ�w���xD��Qs���V��y�Vs�Rj���'����1o�U��+4���Z/�8_�!hق7�n�G��Ł�c��#H��U6�|�]X4v�o�!o�)���Q�^rxh���e>�]��2��C ��C����y�*^��3�W!��8磴�B���.�2��oC�}ߤ�
]�潺�	zJ�$I�6�m��V��+�Eh?���g_���jy�-�6+Q��N�i�Mf�7�fUYh �A�섶�F�6�U2������D�8_����f��y���ԩ��9�1��}�������,RL;����l�YHD!��k�9���F�`�	�V�eC|!�os[�cݹ�O��WqM��s��~lq��Z�X�-?|� ��7 �aPa���MS�U�bN��!��鍴<�N���i�|;��&�'�4u�<KO�X=��pS�S64X �$`�#�q�����\թzf��Pj[�(è��[@�ҡU�"���U���c���vvn��*4)=�p��s������aR3��c��f�P6�mS��Q��{:>D; �;Hx��j�(�E���`�h k �mƊ��{<^�~�GA�e
�u�\�KN�cf�����}l���b8�pQ^�	_}�^�;}�Q
����vH�O���X
 $&A�S�(�`^�y=���8�q(G~ꢕ��'qj��v,Q+���r�␖z�;d��VC��?i�'D�a*�^�&�����}���~��k |M@��>X]��Ԫ6�� �/���+��ҁRL!��B,21�z�&SU�p��#�ɣoīfbk����(�V�r��0��ϯ���rq!)~4�-�n�^�ߪ�v��j�������n���o;ɿ5�L���a1T�6�k��n@���������}��Z��6�1�\�����<�GG[L�	,LD�d�{�;���:Q��ߧv�����;��JT=�4�����.Z�R���oE�#���|� )mo~{�:���2M��hA�".�W{�;%��K�y��?t� �T5W���^��((y/*�c�r(�ر��� _��q%�B������")�����	<I���$��z��m�Q)>:�ʵE�DTg��I1�tf\���ma��b_š�5�0ly�H7��Q/щ��@�7��(B�)��7��.��!X���zqd!�.�;v�W������x;��W/\�Z,�2��˵�|l�q9�y~�@�[	��}�@��5
���e�\Z�������Rwca!�B�u�B.�On1��'8h�ǨOޒ(=?�Z-5��^�$}L�Cp縍�e6?IOo�´Jct d��_�e�T�FJ	g����V�EpB���LqS��)%�cA��x7ϝ�dW�uq��=u
��*ܤ�D� �{U�I�5��Rb�T�q�G��4���j+�ܓ(�����q���)_21�?/���U0E�:�#�R�WdBD�8�qY���u�t)��`�`�Z %���!���f$�s>1��^<��a֌{�5_ā��g���C4pH�a�Yf
j�9�>"��44�L!P3
�+�mjq�%����OOrzx�)�_oPUtp� �AY��A��Cz���xG;���Ҋ�p��Z�up�^���[q�e̊
(���:�S�ۂz����z��
������k�o��P��s��gX����(�}|�24O��z�s����ϸڅ���UW�V �~�W7~��ʳPy?-X�Y�u�[�Gw/�	�Fd�u����#:���ޖ�բ�4��C��w�xo0��n5Vƅ��������6�+gJ^m�f ���g=P���}�Vd���**C� �:�5ۯ����[	�h�m_�V��h�$m��a��w��g��ԝ�6�wN�܄�-ZY,F���=��2��&�0���:��2�pg����\j_���5����=$%�L���j��K�'.m��jٿlX����@oo輒v��w�H:�B�篪�I̯���|z����ұ��@�3�� ���n��MPJ��=ܥ�Q�D�>�ė�%S���7��J@����Wd0�����"��}Z'��	4��eޛ�) ���K ����r�'Ӫ��eV��n_�Ŵ��֘R��<_?��g�-JO��7�<�kF��7��y�NVL��὎�M1��\����������c8׻`4�LP��Z�����#�U8u�ɼ Y$C�%c	�~�;� �~���f���	���`V���B0�h���R~b�4�S�!7�E%��C����O�{�߮�Ա�y?P�8����M־7a��քU�X�@F�ߋi;:͜�m���J�ȓ���o��F��*�Σ�i��}1�y�� �'�L�RJ��cW����jo�0�)�vQ���Ĝ_{�EH#7�Y;+���M��*D�ȲBa>Yt�����=A����@yV���Q�fi���C
�A�v���"��b�Y�0}1��������y��9<�T	�B[,������!Aƴ-�bC�蠠u5�:����x�=���9�W��k�����vY��Z!�����CP�GN&6@R��u��W��с��,�|-4̢�Ǔ��F�S���?fJ6�2�=�@H�{�py��Vv������؄'�#���Y ��ݛ�j�k���=���e%�/�99cܴ�q��ԯ��䛟u����؎Ԕ��}*0���P���*$<���Ci�5Kʮje�qs�)�^a�-}� ���E"�2��^K�r���16�r�\���9��jO`��L�-�^2���݆˹�?�
zk�#����Wr���#�~�1�m��!���ϽTc��$.��i��]�q� �mic-㚔]u�=,��@S��?G�{5���D4R�C�L���B+�����p4K4�Ή�$y/�r�/�޺��)��܉J�5<1����%P[h�I3���]��\���ͩOfU�1Q�ڠ7�{Eͷ��( �������q�\�d�Q���
�xb%�Br��Z�8$�~}
\2\W}ω��i��f{@s!�'�T�,d��,�K�O�g��Ҹ�{���(��HXұ��m`�_i�ĝ��#������K/_�-P������=)Ug�����g̈́Rc��4�HF&Z����5��:��"�9�C�v�u�Â��n�w9��t�2���ר�^e��#����u��,�,�ǖ����T��i@yo�ȓ��\��,c�ࡠ#�/�Wct��j۔.��G����EU����z�ǻ ��~���s�w)@��_0� �Pg�(Ph�%X��$�w%/��	N�o�`�]9\��΃� ����AW�Ş�24�z��PS��&:
�A!�PbPUf��\��e;����\˖e&��d|��5P3*��s�@�Z�9�)=���WqN�J��K�?{�Y
��q�Q��>���"��.����R�h�^Z�G��K�W�Ѓ��'�E�o��y����0cv�<4�(#�;�	�;��%Y\�Hy�;��-�ydœ�bXP{Z_h�R�����Q���B�7�%p�U�u�t�x���o�S��1�2�U@W�,���G=�������']�l�&�Z����:n,��|>vf�dd`+~,mwwG�	m�V!_?.��1�U�ى�>~�d�K	�{��f�!-� ��ViĦ��ݩݾK@�jϿ�P6�ғ�ޅ�!���2��h�N��b���� ��5����qxY��Z	��H��^\�/Ӽ�^�ƿ��ٹ�@�����������4�K��Ȭ�TA��j<�W��2|B�9�dx���!Bj��ނ�!4�oQ�\.(f�@1�`���f�1f[���zW~�ex�Qe��BIM8]xmHX)2�8X|�~A�9�1����D��L��-�e���Ǎ�,��\�� >��Zu�j�h�V�O����N�(�L���4;�u�T�q����_��"`(^i$�P��QJ��VͳF#����h$���H!�,�\�PMȒ_�O>PlgX��p#5�|X��D��߲�Be>Ȼ�2�s87�w��իp/� �~e8�(~�\5˒�ef��0I�q�ژ�RD�(/Xu��5@6�S��������	MG���u_m��.f=��^F ��z�`��m���a�s/�w Eڮ\�}t+�i��AY��ң}�_i��d���~4T�jh���u���� �)#k�[�$W��E�>�K��/h�
��Y�_nR=$_-�m5W�'�~��E����+gQ��X3/t�= 8{;�mGyzx��m�}�q��,��T�tښ|}�@��J7h���P�v��V���`�,�4+ܨn5�$��s7D�2�1��Jjû��Gĳ�v_�Ex�C7V%ڑL�I��jw��N�"�rnԿg�#]��p��΢�
u�H}�
C���*E�{�Bx��W/�c�M���5�Т�w$�tl%� �h�'�is�N`�h��y�=b�h[����1$�px��A+<�Q�iCbˆ��ul$���Q�BK;�࿘��^Q��gݼ�y�)H��7pU��R1�a� �VpԮ˧馷j��L�H����?��s��M�ߒ�k{D0i�u0�Ŀ�^�H�O����2(r��Rrv�~w*G�,���h}ǚ�R�	�`��Cj>�ݣ=�4C8��N�K������ "�s�6�� Ņ�H�U����#��S"6�׶������1��MW���	4J�p5ّ�J�UΒ@C9��}�'����ӢtH��@ʵװY;��~�XF@"v2u#��CQ����*�z�-k���b#�:F�8׳����9H(2x7	1�:�H�7�\�辟F/̆{���0����j�i�(�[��yl��(Lr}E�����4�d�ͤ�%L��Ol"Z�"�B�r�?�ݏ(i����i���tOڍ�u���)���|4�(�U2����r	{��M��4/���H%K�hd������30/����;G r���Qnwf���5��8����Op�7'��*�������#SS�/!=T��=Kt/�o�#>U"j�4�h��H��yw����\�Χ�����L��^�X�4��E�����#LIu<�~���&3�-�:;��Lr(�u)��Y"?|��K	-L�X��س_s?d)�'P1b���>�t1�- �����1f�O�`�2�L6' �Z�W`D��(ڒ�4}�{./��yvv�͸�Q/�!&�[����Qs֖�p�5+}!\�>��`����-���ʎP�t[��"OH���)��+-iȶ���6
�|�\�]{V$I"����]Nh+h���2-bӍh`t�n��R��!#�-�qeQi���K�+`�GD�l��L�v���U����N��e��&*r/g�¤�C�H(�<��r:��Nx)�� k���ҙ�%x�Ŕ�DuL�����o .�$�膤���C�����FG�zj��{P�����{m���x፺��xU/]��w��IJ�^��7�aX�>{?�Nb��I�==�]t�`F�#?��ۏ�9m�d!l���D���&1����,���sw�9�\&S�yМ�a.���B��o$�#��~��'�W��=�ߨH|XI���oG��J�/)	
^'�e�h	�?��[��ai'Sj���E�\��	�7J�h4w��ѫ�K<��ʮ�#�JfV��F~�xe�ْ���a��-��Ox
y�%	㶜�P+L/�� E�d|�Z�>��q����a�-���K�Q�͔{�������՞��'���o�
>�ߗ$���ũ���:�<׻hT��!��|��Z!U
�����Sq�۝"
���Պ�x|0蛘��ϸyުʧ.�UJ�����u�ؘ�ӵj`h���z�2�����qޛdJ�sn| ����M�<����\�5���h�	�d�~V0�Y7�B�Qؠe}�
��1#F�'���ݩ�D���M.��5߷�o�Av��>\p9�7�'"��>I}�����.>�6X;Cr��O��WG��4����@g\-�R2Tmn��>�öNi�F��8;4Sp�_l4y��%��D��=���dE!�&Ϝ�w/4��C�����G�	��_�97�icK9��w�l]�23��9�K��D_��9��ҿ&Q�蔎㧂d��C��-�[�G@���GV��k��VS@�����`K�	�cb�w'z
�bHzL�{�uKYn��=����ԒkY���%B\3c��ͬ�>0��%S������lVQr�^�ST�^P��j�Ǚ�'^����+H��)傧J�o������$0E9/��#�c�x�*��kI!Z�kH��o�0��>$�r�̏H~�~O�����$��v�>$�,jC��w��r��H���ϙ���wy�9u��C��USdUM��bDe���p����a�NȾ�@y�vk=3��Bq�	� G�VhP���텭e7��|��i���[��YX���b���
�_�_��Q���/kX#q����rMV�c�7hUF�����]���8zv8"���[+X۬gv�P��ׇ^/M<$ȒO6�TU��A����
��I�)�tk�q ["�U�p��N�*�P�}��*b�Ȇ͈c�u�D�S/#�9J��n�Ȱzզ��d������3���f����v�A�jb��接[�!��,<2�+���|.�^��vl�;�NG2�4Ҿ���؀]�@$��E�Ӎ���߫V�u^�1y��ý�sńH��ĀE�;��N�0R�r�}E������l�6A�Ϭ�nd��s�����;xs"�#��Z=UJ�������E;���=0f.(G	j��K�&�	����tC%��v�D\s�>���)T�4v<��k@���O�$����|��B fd,��@7���þ�?X���C0^���`���z���@,����������D�Z=C�ni�JG��'`��QZ%�R�*xM��l�$%'K� �@=��.���}G��dcgy�E�0��i��>V�Ni����Xu��|�w�i���R���*�043vj�(K��°�a����Z�n�щ�]XM�T�C��'E���.d�t�՗ђoh7�c��Är�V:&�j�Y4�������H��:���K�\_6W���.��SFک�������?�j�XdЎH��p2�F�&�Qx@Kٟ^2f��i�d朡�sFD���%֎�g#h�A�k�p��~?מvQ[vvoۿ�-�����c�_��!�ϿS�9�]�{�̼��E�o/'*�I�'��:A~�#�9�S�Wc�ob�'du�e��U,�z� ���Az��{
J����~�ٙ��Œ|ުS��_�����Aи�b}�O�����t��u��nOA��>�Mx'w}���^�4F ����*����+4�l��5?>t�L\+��^;l�X�����,�&,7S��
�ܵkꂍ�R�ܳ���=E�-��ܩu�@���p��<%vg��q�k�F�2�d�{�,X��-����<��l�ԓ��k'�ܠ�7��uU67.=[�"�?�@H&��:w�g j,8��z���������F��s�=2��Ĉ}�g����x²_�	���D!](�P��"��ȼ��<F}��if� !h��"f�~A�'E��$jm�=h2�W�s��$L�C���R��Tp�0�tc���8�ֵ�=������Tᝁ\�Շ ,�"��l4 �}&F"M$�7�OlvN�~X <ǠQ�޻��:Lb��l��^m8v�?���Uy���`A�����$< �����o���3>3�w�V+���u��l��İwm�yP;s���E�������qf̩r6ǯ��חU����� �z@#��cLf�͒ؿ��_~K�=L���#�]&��a����C(�nF���N�=E S�UE�	����;b��o�MK��v"�)!mK��c))]7���nu�i�K��8T!l�H�V@�`����u?qՉ�\�?�b��r�/\��8|�I�W��#݃�U�,�(<�3D�8�K��b��!o}4Ft�m/K��.�?�������k�bP�'r������hƃ�Y˧$��A�MD��٘5�ͣ�w�(�$h��Qt�
���7��=k/� \M��-�|�_n:�+B�U��r��/"�|me����ob�Ěq���;;��f&� �>�s��t����r�S(����l��_"0,�#��$-,*<��n�LF�%|���$�1C�-F"B2Ȱ�A�uǮ��U)BQ�e�d0�DT>%�Bd��\�� ��i]h���]�¶��>HP�d>���`�{��w,� E�K?y�`�$�i��9J}ޜ�-�V���͛he�g�׋/��hK��?��~`��{��5+��gK6V`��U��4�.[:+��]t�wv7��vgf��3/�xc����P2�R�4}l���6��)	̻ 3���3���U��Ԡ;/-� �f�""���"1�RO
��9��f�Ǘ�C��9wڜ�i�����͸z����J�6e���G�ݍ��п�)�Dw�T�����KA@���������0}��m����4�I����X�B��2�%���2�r�һ픊�Fz�W��tN���xC.�Uu)�f���x���,�yr�J�7�AW�(7�`˦�򝟫��܃g�N��>�D��I������#�%�)j�N��v�