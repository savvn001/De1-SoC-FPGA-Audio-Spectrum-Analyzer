-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qCkCgx1gp0TegwYR40CoyxK+reeTZ0J7ikepv2Nx9VfqWEPoMk15ukrSXL7h+prvrcp7RMPjH+Cu
D51lDyqJVD+6Mf8QO96Ui+qjFq6wL41xKVZsuSrPOvLLENYeM3SKltIqT/zZ+nhLDAtcrE5eWH+D
qJaZe+BfeR+lGVHQGV+wR+nTxuN/vsUk7HoJDUZ92O7hYlqDdaVtIiqK8Vaj1sv9jPMoE49sbqGT
nZj84zHgNkBH4Yxl4dUacJ+fJP5beFVsqz8Ip3T2jy7/zBnk5QgCMiborZ7+ibzP+lKXdmFpJgBG
4WvvpO22enQXzhfHK84xvV+Svogn9M8pPoY+GA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
CHqyQmgGp52k4YYRZzrAavm7YxjIXN77B4yjVTVERBnWWFytZ3M+jmjxl6DdcEbrmrrFsHNcL+UR
LTx8hLA19rfzWa8XUINvCLN8vsA9DwDTVJVWg1urppTNTbvzqVBdp43fKQEte0ltMFHMuLYshsGW
AaM9aWSDfL+T0cplC9WRnKlF6lBEkNyoKjj+bxp86oNmvUp5MOPseJD15O0A4aspcjpwU99M3mGJ
EKAg0CFtkNBtrdmNXSn9dGXe4UasCyYuAUvkaxk3K68b5yitqL94S7qzS+3TmphAn5pC8xzQdy60
HDqrrvC3t5omlAKEPXZ7iNAe5g2yaxHcfy7YQydRPPNc6tnmhMnds+VVqzvVWo3zcx+U9WYPZJS3
LiPxaHkyYIcQpBL2lnQiL4QQ7N7XAOkIeIU1xUztcTjCe5aWy7ZuyjQm/2m/+Gwxwx59ZlmRiksK
4IgXtqF23xtNFro/LZVupMyi6xXcGlprhI1KZ9bPzWRdUPB7wTOVIl1J4WSmCn5+5jm6hR5NiSto
2W568s51z8fMem/SOHoDdVlogIwPMVk3RWZgTDKltnOFGiSFcueVZCubKYlIb0ch32GhNQP2SLnm
WQBOx+YID6bsk5R3X88d2mKPpGpBAr1Rj82SbNtcGS3tFSIZOhqEtSUjQ2+7wgjKCBIG7hkJIMji
HHw5z07fDiGc08JYdJvQSmZWiMjcggxchV4p8f81Zy4zv6dgZg0c+cILrFlbf5sI6EdNTXfrC1t+
xnkeOpWAWAMUYDxB4APlipNk2jwGOkJiuiwLkxO0fDeDCToMxt51S2SIxLNxxaKxhVG5Pw4+L5ge
8yK6wtqmM5NokdcqobYkwjFEx1kr8AuLFcUIZSi8fSgJUcYUBEicvvXpNIGtOf4UDdvFPfqi/RPE
1T9bSrQuCHttdu5rXHFL7/DRS/NI44/hBtRV/OJFthdNjtwEIEkFndSOr05YjH0sTkBuuU6F3NlQ
t3omHSMRfouo2NiMa27vrYsJ16I+l9BavWtedjf2GqwMAxN1ZdzbFMIbtAZEBW/Roo3HU57d3HQx
HpaHfXpYi0lzA1seKuHaK2gQ+KVBjEfYDSRnVgZj14SMoL9oyr20ktAhE756boQ2pmDEti8rt33V
8rSJvXHXo6LuWcSa+OGnxmICCSr3SbXr8E28qSkFWq8tYCTQ8l2mQmlg3co5HPyoJG5YLofbGlcX
Fz04yT8oTLn4reGMYqpIShDXQ5Ka/ItRbW4YcDyuCsGCypntZWlpm6ze8uD2JPwxyywn9weiN/rh
INGLg1w0NKNMQCkBF4rz6s4MhEAsKsAf9Hr/LpXNtrhYbCTpN2P14yOphw428mt66fEHtV8B7JE3
Y9Sjur90BehYuAsujb9l+Isy086LfhVO6OuPUS0L4fFdqDry2U4dBw36QTyCYF6rf18ZkYOu8JXb
8ZiFQ46vKnAveAMaIrMtZEu83wFJ6pmDICzde7ZcfIq77CXm/6AP18N2QeK6mCI1VFCYQGMoSKZy
gx0Yr4pCluhtavEHE1NXK5Fwfq2y/cwu8UCZSa7W/mtrVo2p2UiWLffR4Nbdx1HWwA3h+Ci3BRkJ
4yIFaAAKh0PVdX7xClOCS9dz4VQ+SWv1WSa2auvyQs/Kz3YCmEq9JZikGrvpuk0AzG8sIdAlagzI
x2vatpN2bDanKwDjaPdKN3oVBLObdiCvENuq6LsWlZLtA5sAB5878vc2oN1Aakk+xDg+SeU4/wPl
BywO6rryqG+gC7w6JUwG3PBClc3s9T/RRjrrswaqp1tJLZlSwrebXZ8N/4jJl0mQDQvUWgxq9RyM
275W3LLW/GLI3gdmcbL6XotkMBWsdPAa/3kC0VrdqHM/c1hppar5Ltnt3YnOvt8oo9Y1FlLJ3Mrd
/+O0fXG3aLpNQEmrUI3U6OrB0i3yT/VSpW0jtVZPTsXOIdcOC/SAWYAST16LQ5SsUYxGI170bmQM
gJd989mlgFNj2OSU223692tUcEubkKXVg1URoNqG1HXOIt/4pGyuMzpMmQLYrM9X+TtPW5+agji8
nr5/951NERdnsBXOCIQIY9OLBdnqZ6nQ7tdFZVRZvoQlZ+SZ7wpNJ67gaZTIDxp+Eandb3v2GoeY
XR3npQepeA/Isgc8WOkD+JcRoyCqzYYb+zFWItmZhkhyYzXbGHUqkJbTpHziyw01fCiJYjFLvT49
mY8JlmO8BCYJEhsWOC+zIFH18TqRpB0ZComOVwoVkWscMDkARW4XAJXU0lGY76642CBquPHHyu8U
gjFJNtgQaV60vxnarIo1WZjsFSh7ZwB3yV834mjvhsOYYvjVY3jGDvNOb5TWnquYqx6+Suvagmok
oSapOF4rnsnouUnz5CY6c52a1gX/7g4HM/5HKTcBfniT+kWAVb3NBUPwNDnoMb0Wf3fmMgWhJM+m
tLn1koXhBA6s0qi1ALQ2Adb3Wo1BCwzlEtu76S1JjyaF0XGc2ua9U9qN6K+b74w5e/YQ30kjjW+c
2a7c2LktQzLcRmQ6IKZPRCYjJpIrrcLSE+2xMtbPHzKdgilGdRUVlKFrje3bhMT+RKdWAwdDGGa0
UnRF6sgGc4UJZSWih545yNQEond3QybwJvUFwjPTpWkRlf1tZaYL9KAOEV598EuRi86vDVksnRdB
F/4OhivCL35lqXeNEvGu75GzNtkPqsQgVCkSo6pMMCFz6O1Ut/t7GTp2iNwSdnMRgjsRhohL/AlG
IgFuhh64kXWKMS3sRQCtIxAdwlR2hReMgMsk94dz3QC+HjTRu4XP2JFg+Zn0D71rFaCVo+xdQYKO
K3sOnj3qb+XRd1WsIDbps05/FTQrCBfVdbULH38wA0mxUFyMszXSQ6NG1LIeAQszxg+oybZcOoG6
Oa8rr7RtgSM1ROKB73MEAwcMBV/WjOMOYesYMX/ge9gLIlMjz6jCUItC7TusmxcYKlf3w76/7YMk
5AgLH3uslACRaDnFlKU+ym8NIZzyH1wyM2bW8zQAfZWlvuTSmI0Lgp6EQaLmYfwUezjamiAwxjRl
Ds6aPKoxkAjikHf2G3miq7SkK2wtFCucfSAbOPzZ557rLXnKx+FGp+GyOfG/uVvHC7rYxwMZD4Q9
Thsb2aNEQ6e9WIqsDS0fwdYLD+7rK4A5A/KZJJ2E/7sx7mHR+8JABFPbLCSr48y29bq0+lov7PF1
Tf262PgF95lXzdKl1Qmrd3TCoLPeuLJ9qeQjclCB+rhaD08cJM81GZVE2Xg/BhCcl77wpu/XMzce
b9gNNYrbfi4w23DsvpPXyVw67lEgBV+qAnSVwi0DKpxB3oECTk4KmDnJxnPeIyWFuJKrtXF0R4Cf
HjxZCV6esM2euzfy5G8MGyzN9+bpOORNKbh0x1kFaILuoD7glg/Qk0OCTK+os8HCdYKs1ziYW+8C
AI2IkDoFewEyo2625lHsXj7NuQyjgxfJLDpsMA6QgjQyfWvf9W0doYhDOQ/vutEQ8RvgFCPKEftI
HUDDy7t2vXH4za4XGiKghFd+yTHZJxECk+WNYPcAGDNcIGmZbwUyuhsyNt4Y4x92n2gfYwqx/phG
IZovXSrNHzCCmANqo/M7m5KEIXiruGzqunZyzVNfAlE7Jn0YfSL4lfnfcsD2AxvTi75tk6Aw/3OO
N0oqWqsYGPjwyXB+SM22iHW96N9T8+9OcvTs/9ZYiPbytxmbfV6LKqO5Hu5C1UaVeaLVaFNNGqaY
W/H6L2RuoyZiL/+OutFbX6k0Z51ziYcg195XkKWvhmXDFzMMVsqiM25D7tKXsCcq228Hz+fIXFLk
k4lQJfgGAqqP6y26KPI0DkBh/ZVN6JRo5FgvqIR4wLWc4iu1ne7DF24mGt/ndSq72rB2oQCcQ6NY
k7MxUSp2uvwAArYycgTAXPnUgqCJR+qnECRu/8oT+LHgG/DThDyQ5bq4Knc3xcs7d70d5SjGxyMI
jH/YnFyKpFL0XwEblKVmc/b+j8Ni7PMkpSQAXAeg/3VMEQbITRRXmeagJ0R2djD9ZqhfG0VV/F6x
KBw2jJx9x2F8cVeFUHHSYAtmn5/8WBm76RCxl1cjhkROtVGA6LLro0hBHRO5Gp24Y3eiCKPzF85h
sUOYc3Jk0/MLbHSMja/tNv+aHlwmtGS8wVgNtAAGva0rfLGqY1oLso+5sonEKpomdSmJrIt5eUOY
ubiX+rHqnrp2AxEEKsT9G/BcwfYeHA6SrESCw6nlEPKb7D3qU7zW4Tsv64Y19pDPWe4rYdwBZ0L5
9AkFETKNh7De1t8k8wk9onsA7d9SGCvoVQJ3YHS6VWkTFnQNbiwkKfrOV10ptbwjFzSJcXhnDQsC
y9ssuKJAqgIHETlY1vxPM12T120ESbiI7VCX+LqM7GPqYnRDhgZ4kDRnqXQAcbaV6CfuhqtOrp8P
IXjCiPnhD2JEywRqgHxLgvzFL0gqHQ+i/mDxU5bld+2gq0j8miqWDmFls8vEk+72wK9b5K45UyXc
gcrkqKux6utZpp/FOwW75YJNzqmEH7NCyJXcBEmkoo4vXon3u9Xby/3yi1nAyHdeUBhthXX5QJB3
AfGmUfFPouOnt3SmLe51nfda5pUHdEU3Q974mklzWdfxkvY14FaSmMXYEqJ2o1PDl/6CSvhWnlA/
LWY/hTSfHKBMHAF9pnIJ8nBGW+8dQ86jdzP+Qn9DwLRU7jg2ft2oPaGyyzornnp38NDSQY7vW0VT
LcH+mQgydZ7leCmEHpVUCW5joc9+N2IFgnOSN4lbeayjT49M23UtSJawaTtelm3aYZR5q6wb7yWk
4b3OMC8Wv2zNGG26wZImvCMMYWDLS2HMoO2pRKzWv8jTU5o7GtLv90JIT40HsLnFd8j921Gc06JR
a5fkvG+rmyn/QgGM23dH5crVEVCIfadiLlLiz9SfAs6vBeB7ODu+pwCermPaoz+VrqjJqhk+CaJX
7iNY/MKMkJcDzKuBRn+1r2/CTTaR1VWZmuYPFB0R5MGid6+HhALMAfe+Emu6DlC+p/vdx1ctvSVr
ZOCgPUSr6FAtghU3HelaePPkTvN8gkUmLiwRX2kQdpcSWB3+X25PHp+1fLLAtP2RCPn008ddwWD1
2j7o6bvog5JR+bBOhQ0cmofpQfcs++0qs5p0mrXRnQO9sLJyFmPd+2GU8qRz/9vFJ7DmZefm8TQr
1UISF89AcSY7KMIOILiMll30kir5daop0PfBQa94tIszZPzxA+DFJ/KydNcNyax8LveXrCisEeuk
K+av6ts1p2TPQuLkhyuCl5pThZ2qaFtfQ7+ExMYbVZZbJQKDuU+cN7X1ngrPxX9ebxgf0czf8Ylk
yy3tb/GE5cCDGwUWNUWdP7oa8PoDgBkrI1OwxO8XUJKV4oevLUvCeqpFygF8mE8EtAJlbwr9/3k0
8pxaI8M/5hAVb+MsPju9RdGRLTRMCdHNrbH6GtV25pBKJsrEN3qAcIfDemb5PpG1506E5hqcyTeo
RiM0T6T5U4vZ/Frmq08ujDzRYYRt5t/qwrudQrAdBn0193JiaLX/whOhmqIYk/bMyiumUbak+Q/k
auYNjroDszrv4lWJucxCpw1Yac/HtNHeEE6KvLXiYqIrGF8XjvzjANyQVYueAvMwS2qymaw7jH2E
59J+fZ32prgpoHBrHoEGy3d/dNE/p7E01x6r2yst1bGG5z/eBjtgguq3MlxNBVwy/vJuCyWVwnMn
tLDgVrNHUtpsOHdKFYZu4Mc+dEdFimTkT4a8pqfPE41lB5IgNMifQP0/xuWmMI5JfT4+8Z/c/Sx3
Op6Teo+n0qJzfoRYt+sxbApHf19IK9B+bRA9kR3AaF7bjt87uwYiI9pAZjrQgU9i/HdS0TATIzOO
OnlkW2zfZ12ltoW4n61GwEbsXsUpfWvQtbslOTbgMrC+zMiIjLDVAqu5N6lwG9Xct5wO3zv5oLyr
3oY9Nj5z68/yxTcE7t2DClvK1qU2TGcUppJ947uy+xmGJ7vDDE028XH6mukpnOijXEL96bFJChIO
rGM69IRVr5QoDwpSBGx8aIKPk458TZvGdsgYyc6YofBH9Vv54hwvItWqzdZQLydxiXoIw3zOYoIC
/6sy4Epv5ePbI8mDpBU8RKrWscJJDTnVGsKCUbG1ieBDZJQbQVHqMFuIGJA0RHYBMtkihgrmiSdQ
Sab0KJTh5JHToQPA63S1JX+QT2SooA/8jE2xt6uZBHUP4EjDbgu+esnMzdHZ/ucf0P9ns0ypWiNz
8aOKuYIHt3LYh335mrdw/tStJ9sO4LPPfaLSd5fsDBb9dUfu8mlIug+a+EDHqN2RLXOagJTRaPFL
JqtxaWWo5HsgPIcUeRyGPpG/4p3JS6VVfcUJt9xIemsqhurt71WaNq6F1AWt+1gMEWTWSKwJoVvn
PxtWYQnYJSGhxENQ4LDpVHKbgnYE+QhFaag4yd00Slo7pZ/XADpsBGEywSbVKL3TD7z70gPuyvDA
5N+d99SwvwGpTAsNWlKga7J1wtFX4JkUbV1NophDLm4A4JPkS3YbxCh1ejPZ9ckG0bd66pMd/CJm
oive1vlxRwjLJtD3Kuhl5fipvLY9hxIhLezzWI2tbKPYYsoMoeFhQ/laC5Q6ayJIkt+JxdBWglXW
RbyOomjuAU/DApaRQ8kRLR4CsupjkSbKIibT0WK/jT/d6XnlwN6X/MZxJU0WkWE1cvPJLZPiVBBT
5PJy1/0+ocbfXErAyPQc2EnwUQ+oM+Egcmb06CgeQILZwlo06s36UweT46xiUpZ8Q3MG2biSbL7t
xjUsWp/YpC/mNB5nLkmlnDg+u7YZDQ235NQnIhOI7a/I6fTYOKKj+dEFXSdwS9O2zh4WE4HwX0FW
MUgf+t5RC28F6OXU0Y0RHMDmqM7Kz8uedJph8q+e+TgitDBA2Q4vrJBj/treljDwSuJ1njP7GXzI
UWMRLVTyT5wu8N/NqNoZ9iImT/ar13KcUu4XJt/Y5kUy3NW0iq59Sid7maAN2ealRKB1nqGCx7sM
Q3bkHCAPXcwSbnyTJRmHV31H8ZecUFX5fegXypJU+ikQ9G5srPOuA0jSDyqfbEg4CTZ0x2jryZXt
4Q/+jExq9Ea4Vormy0HwfmiMa++YBWtTS6U5pH31FqPzWwdFht8KbZ9Ds9qTTB9iTL0I9v853wAQ
Zr240kcJidtWqhW0STSI/cBgbnvPtIwfolt2aPcQYVzvNyxDpjfDWD1v3TTm8GClJpugV/NGzuIN
iS+ze7ZPF/TTtY6JsQaCEiEkAif8EpkbZuH4zPnBQICad+039kRfcL5d/ph1TvJNejQ91ofDUyJz
PPVCW8VvzM6R9ohQZc/4mOvzzM/CwUMw21B7Am3Jw+1fTa2c5T8WzKyz64eVMpbUf7ahkJ4+KYiS
kv9y/Sgbm5/0MxhlMfhv6BaRuTSUu8urN4tmCHJ8Ppx+WdIZ5BOnLrMPpXRAyPa6DDsjRWjS1SUe
VIOljHYB427NvwSaNgBaGCxpKuohJQM58rYkQdyAQQ4dwQzi800F0MMtE8+XeBfgSiXd0FAYx6SM
ec+i1DAXg+6xMdU70kXjKp4W4aGH9ALJX/dSlHbqAHk4tx+QGFSkd1R+MRqrxz0/4pI8sKsIbLOy
NUq6FF7Dws20z7yBgbgzwnhF6TR2n94n2Z2oW7xBzPdnZwASIy1cVODueVN3gT859aCHdeJF75Z4
PTN/dlBniMKNyj6wH64Id9TBE0IJ3n0C9HEjNF8lr9ipyX7KnwaisSKg/DN6vTJAXBeX4E6R++Cj
N4hs6vpwZlP6Y0rmxhFMXbB+diINkJV/W8w4c3Whi9k5FPvmJGvqeJiC/xit6Q/mV6lF2CTo32Br
fpx/MmCYW/hhgWzCQN4FTRQsOp8SIGVedKBQK1hNx+Fc3CECKw0GuNosOpjaqf+Lxp3tqdA+S9Rd
gzGh2pzbg2XjEMAys0fR7qANMm0P7uOK9wTagaIPHx2luRNpglLWu5yn3RUOGwReUenSX4EL+AS7
Nz+gH0pC6oUFuFM9+V8YlAdh+F4LmiCaBDpVmt0TeeEnKiOD666PzMC854uh3hDeabXHZ9JgNigf
lZmGQHgny0pDiZ2toVTBii75Xbo4lToaWzrl2wPniWYkecoJ0Dl8kYniiRZNy7gWN3whfMof0Eud
IMDMB/q3QhgIGQgn1q+vJZaYR1yn7dmt3J7ilDNnBgGaJbn8wFYi1hydK+FbpesEd9tjVfX5smlU
sWwgGlPEkxdJ6lpvXCnDjEioTpwJPZKamjPlhltwUx/bTZWfXofo6IkcP+4UMoykByPDl/HS+5YE
+i6mbNzwbYKHnqqeZU85ofHuM0tqaufiF+yiQWMNYAkFdUeZTZaLvL64IhzbK0Upuk5ZExMa13Dt
wKWdT5tfz+r9azZzy6qyeqPG2I24jcCIC6xtUFI/RYbPElXJizr+cKnq5YoWYRuK1eJFyC4Xh0ky
tlIKJRb6rK36HeMnn1oTDJcvwP49tMYbkFA/GsE8uSMItPbjRwyP6IPKX8zAK7bx8oMwK239O3pi
clLKKCXnifXc56Ne3prLad5lHPfn9myDVhZ5EamY8c0xLR7Nmc+KBxXydWC5FEYOcZhOQvLYMlRq
lpKOcHHxtcVoEG8z6/zVB8RUQv3b4tZV8LURaLzxa34uLtbjJsJ5oDBoFBV7ZOQL7CnNJG3WhYTL
RIgo0Gw9cQ5C8cFVum6uOiEtC+f25zFkAtNddBMxY8pCiwhEs37irS/PMdIbi1RxLT0Brm/uKe9e
EPPNr765/C4YU50+FDRgwahez4GpYrEvEcaHn9AROSkS2skQ3bYiBYFhgTtYjbz1XWcT2/Khvjt8
HXfAvy2n2FLRq+ev1I0wbmy4zY70dLAAezbI1RDGXa/Gy+gtDp+IzGHx/IQg7FR1Dy2MbhRvZEx/
z2qKljnIrbQxxuUPLoKQ3BwTKWQKXbf854H8ezH8BiqZHpMWi8gxPVGXt59o6B4N2qL3//qYlNo1
v6BBwU2XoMTvJwIDA6u0mMw8/im0EkZfcgkBbPQSPP+AAvGwsw9B6WUgR0GY+PbcTQZw/nsCjUDv
ReKpiIlJZbr5FzMduN4sTMBnFLS2O3WkYCzGFozMLTIKIm6t9ugIZK5M5RN6JYu+UNDsgKimvhKx
35yNBmnbMMfAuoRXsVom5f/O8w5a22o7b5jwebxOt7ymdn5kSQmNlWjaBJMUYdQ6hGG6+lgIvFV5
LmjlnPMUaK6RZ7WZxw5XN5JSXjRHJiCKGTxWEJ1mycd6IYtSyaqI+2oGnc68Lhl7xZmNKMrXvv9/
mgw7vx9g33XpyA/rdHOyeRlXuHwlnjZVR13EvtKolCNw/M9XvIO3po6l1Yb1MBUyV8p/8/+4K73U
9nKHGAUfqtp/BxyfJiLA7q/mfqLGkhOl8wGEvFHa70lgZo1XnA70gOS3OpK0CgSXyxSBV+4LMueG
hrJgOQIniuCSch30NkdPtXWOnD1HOcQiEn5+11jmru1vMk4iLDbVElBOUVYXtLnSlRJ2HSyRPDdt
zK2nthXMtDNjMic5SP1Gf6MVapLUzjFd9oWmg8R4daCnjHR5NXJqd7s9TkcaKgZ+m4NIj0TPQxCT
li+i687nCpc54LJMEoHHz1kFRfn0LzN81xNvxVDI1hCI1bluun/g+glrUeSKvszcWzQfXk33UW/3
nv0Y0DOKjPaPtaVT1TfnWWJkCibo7K/gPUzloxt/IMAeSb9oJd74xkzzkkbwSrdVj1TbjQiyxM1g
MbG+kN16Ht//kGSZ5jgZprUcG+kL78PB4Ktw9rIu2Lsz0kWhd4df9pkLa3XUl00sKTPs70e95Qco
RgcaCPNdRNygNsWMpXT/NDY8tRk7ZGn2rwU54C6nUsnHBIOMrwMcX4nyQO9fhYmvBXeh9qzfT4rq
+blgjNigEsIN+Gq4PWVmC/Mh6AfnLY87VYJnIDX5OhCWoiuHJ0m/WiZWHen1PiBSqQW/h3QdZUrR
hkFCtk4XMGxjLKewao3Cy55R2DYo/3dEcBmm4RkX3O0ha9UUM5zGJ77B1H+88BY05Kl8r51Gjd15
q/WtXBNBr9XQdgk9VzY7VtOVfVJY82gh0r0vKnsK/HBJpsSAou/DW4xI/x92XDmbzenpDGXRaNXK
k+OQzM9VYGIBv4+hJxOE/PFMtENyvfUIy4bL7Y3T6Kig04qJjcnvuCz7ElNUc2jnvJOlmZmr4AwI
Xudetmwk03kioD0JR1zIZvycHeEPhidhXPH3pqPogVipZOIeOJTHPrQfMS0mLoDpdfEu2UQcxI4I
ncjpDG/TLOpIY1Au91//IvnqgBjGAX6I8mo4nmi77EfguskGoV+nMeZwQzqu8QR07EWxfJ6gHDYv
HaJdlmQ+iIpCb9FPRulc8hoARHClhf5n3Pm3AZ9NSJC8rXXBV3lTxxr+j2DscSAoETqfiesbYQ2c
ToCdISdpI8gfz+inmhXCHylg3hG7RK1m/4TjfzOUOLP0WeQmarG4SpzjENB5rWzPKXRfrAS3bbz6
8Z5zqGIIiAkkKK9Sq0INJHII6d1yvZo04iib4spN9Ra4sdv5r8Btsc1L7sGSdiH1cMxFBI1nSG9u
M5l0tPVcY36ZWgL44xqucvaj0PAjcsCINW8tBn6DmWNGRLUndm+DrbNDDgT2r8Y/ZT9iH5hQBdGL
d/R/H47S7LnB4kJ5LuJ2G7VYhS1kLY58po4csvv3p/JjNhvCQ8JrU7yyWRHVbQ01UCSraOiYXVgj
1sLB6RCfe8MjcC6PT3q7UKKgAAJAMpneDikfseT1vnvmAcXHfL9Jv3RGToVycELUy0adVQ9MIvdq
9M+wjzMlVhgmvtBAmfBK5dKxh8mng5DBbpeV60V4r+MU7MJNrXpW4KRjfvUVaYRFnJJy8Dr2Qd6Z
Dyj/6ixHe+dsQpmrPTtNX8A281VKmsL9wDB+ltK4TaZ38cETN1y9cWCxXtqgw6r0895BFcCJMzEm
420rT42YWkLHMZQQT+q46sXnQ119L1BLE0GU8eZkoqHI5fXp42jzdYtDwspC9+YS/kiGoUag6/mj
NCmIpIRm+9WSt7TPjgT56DEWL0oJQ4xMGQgWI2GmsO/lRm3c8AxNQZY49zANoV0prW2fyoaeG/pX
ZKyOn5vxkF7Btnv1kNqYbd0wHbfT2HwEEs0kQhFkjL7/HPLATQYT5Trux9YDsadlYyVtbHqBy2hO
wxKjncaebo8HYjfe+s4TLP/TqlE0QGH0KmsJc366qPvlSHXYVSOLv6DFzLoEBVr82stBsQByY19X
JF0vVijIg1hARRwYSOAKcYHQCbmvvZ9ivytipLcsJH3agCqDixDA1KN5Jbm3JkYnJxAP3s/ELuQe
k/9tBg1EJYTOFzpueV44zTijAI+hQUUuLH+uB//R54Lf/CpVNot9y7Q2mDoKrNXqpW/Didi/u96v
1f+7t7AD6u8qGbH/Id6zooGLQeh+BkSe6NShW+WhRs8OoBdW17Sdcsrly4J+hUCMuwRp7fRcXlWH
yZKRpkjE3javt9oBoEkBTet48uwlgeSY9lrHh5fnc8tCT8kQh6JGvwCq8nnRYuNNv9cIAkZ4zaXv
s4YxHIhwIb1pk/LDXF49SubWndIPxo84Bz6klQ49ertHz5WEkfhKtTG6tbJVH68VUmnf0wt0ZSAi
gTb1QVoKs7AFMjjarcmfutHkTppsxd6KXgnNeWpnC3sZg7nFN7FNTJq6qh8Vm076I2gFGVTQn5mb
XX8AZ6aTiJqNLVdqgjKn+BBUguz7KrvEfDFg46rYC1/NERhMLGx1gHW5qsTunsKTUTX7X3wkzqqe
jpWJYtC2+/12EO2nVIVLuKq7jFLaINTQ7h7lICriHxmzO7UoYzLz4hEZ0pwlHnfOBQvnjihNpDuo
dK9BQ3fuCyFNMGPXpSHonreAMp23TfjHT6W3AVq6O3DXQEtf9VZ09sQhjkhOmhId4E7tuSpU3m3W
OErl0c4dZTdfSuTtCVzUwWffj3OJGii6pIVmCe3CnPOVrgT5Ytbn02MrfSpmw0d8CZXu/nb3Zr4R
tM8H0/GKkCv0diFUe5/hffP4RDLTuNJDTjckHCpGCy1VTyAgLh65HjUVVV2hvFJdEZhUHHI3PUby
seLO01WxrBaxDorFhVqrj0hFFCPj6nfPW8VBtAmxoYyrTOAlDU0NlFv/6aruPVp05bHgUeUm81co
CPl+yI2prnwHdpJeDcDZd8TvKa3ygIxTYT9+Ilioph1vv069D7EZjLAbQTL3klygRhoNiQCAxfQG
zgofliYGYtIGrIKW12JhxQoTPHUTg+586PMijHABPAaQeA6j4tZziT38UAviYWe6loAAVGwHXXxh
uvxCAAFH+lBh7feuCwdSSoRl3Md0T9V06+RTBRBMmTehYtVZuFrXuCyLHocWzHhSz7eTefvXr5Yw
kikqKzO0StNE3T7ITyhI9jgt5uC8hWI4j4hdEM7t+kT3jmbcAmGQNUB7ASN0aE0KHOn0iCQJ2psF
IXFi1CIr/peUmVEKajj4K+ffw/LfPw6EavBPhMVlyT/B6lEJtRFnYregWwbSuY663aRtv8B9zqV3
bsBw6OcY2O/QQ9DBIirYFSrbkal/ZNFuuoWTaKRR6u2OLXN5VYIUsI51/c2Xx0LShPZqQQZW6ICY
EF5Hw3ycP67Z1dqNLTA8TiF6X2uuYGUoIKePbv3SuY1F0pamAxMqSfn53B+dLGNQUt8ncVea576E
NXuXdI3O1GLSAVugnh8KUNYqVTp7jW9TwbSO9FGq/YqKSiqbFFTpriVDW+KWmELIQ2QkV1MqM+tY
4Le6R84SFGBmnVAo+655AFv3C9TWzrLHZry0XcOtyISxjq5rPni2qJU0lnMxH5p0XNDcgmXnrAVK
x798A11E5o66bpcTmtOj1xKTa/uo/I3NdDK2Ocm5SbR0L2cjlMUzpM6YDg4k31jevVxNR2wg7E/h
XbpOrtGY7dIzOHvyW9HMf+s+9dCfmhFGky9RXUo2aihiJvBBMmVEos+ZrW0uoEJ7rvh+kipWZb9N
DfuaK0+uA8YxuQ8WOw6UWQX/FCtXG+qaWkMsK+OJXOrC9lVm3qnxvZXADsy31yBj/Iskx5DEY3AB
IP9qqtnCIx02ElFXfkEFk+pZq3LRyPJqdl9/KwjpNpkk/Gs398e2GzShBDwPk/QFXkNSpjChj0hP
BgW0RK02u6lHOfUsH69gqwNe3F2qODJwCfkfqPVp1tLF9VeIp2XwGxRVyHW16cIvVQK/6Lv92IwS
IC0ajOdixIQ24H6weNiYYErwlV+dK8qYR2sSdEuswTowVdkxIr1k07kqrv/O4d2PIbQF+HWHHQK1
KETEXmK+Z1ve9TiqoquK7FiAt/9ArnCTNo0+XcAYcApdGk5NKlzFqIAewbdgUt0Od6lHX1AYv2XM
jHamk4YRYAKr6tKteckdnyfMqGMnPXl/zq034Ql5kXKdfcAV6XXYW8o0DJndi6MlYUavSj2EFtMq
8vh4jst5r9JzvdjM0TxOn13Z0MxGxA+/azy76yBUhs/pPbTAPdTtJl7ywXq8vhjt0AM97DutoAvy
v4pjgAsibSJNQhzL3wQH0soz7F1AvbYgCUvEjA9nin01sccG2oD0b6nKNCYqL+drFs+XeIQ5i6sB
K0BFNTOzYfHR0dQ98Y28oD47O/CZuFdXVVR4aE8DyRSTEKBsvu2LYtjLJSwtvzp8x8pr13k=
`protect end_protected
