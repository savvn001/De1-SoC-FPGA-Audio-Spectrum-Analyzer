-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
saNqHk+I4jKFzkh29R6nexEyPNXJsaYAj6gDFgQxyn9ypxweCQYd4mMeouETNAG8j+arGVRdZkYR
xGXu0v1DqWbyWA71ZNoiqBPBSRlKxmsTeFC8dToyXpcrEi+s0u2jggVCzzpQoqKp7nb+fv13wnNy
WNA09ZDzWX91d9mlZ0RqwvIdp1BsAjjLWW5YhmlR6qeVG8Ci/ZEX53j0bS+zZdixWOH4NT1DZ90E
qCHIy9vyI3ZMYc54JmjoW3dL0H2j7303g/XOxDuZTTOB8jaMg5vhzneIT4unlA158eEz5K6rSd9m
8KQVr4ImGOLLIlOR+x3ilU1WCoKCXrjVYnjpGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
BRRf28lMpwuDAcKo5oDWP/vzISKWCzmc7bx5s6942kC+tHUeW+cHOjPjKnncJ+rXJxXeACxg2Aix
eUfK4Q2urukvSPlHb7PZTKtZrTy2J7ZX3yGowyXH6vyrxx2RMIkHW1kf2Xv25tMXvEdBL6WJy/aY
bX/kDyLzI9dW9pizKY6EmCjBJxLJX4r9/3K3ChlqFkSiXqww35Bm/hQejNcpC3Gs6JobOz3kisgO
i57MuGpeaWT39e0Wm6L0c3csY3CjYnlnV+Fc9RRM8SLcxoTHylnUqibXF7G/uCbZckm+RprFG/zS
MmTiCOPFrMnSvUdrLyFMjQdxtdyoonh7OaGPehZh0XCDAhthbSoy4+GwdSYBsJ4pC2gccpYFMtKP
HlOy6vBvYM/LjPlxmQB60IAu+NJcqLDwx6iSqSmPDRCtMM1QWMXvWnWrpHEtP+2onu6pvBaoly5k
8SkaMU2YHIjyS/oovNBtVRTnUAR1mScLXyfkXhfRvd8+ZsIPZD1bsHzNV5Mo139OBR1wxqO1/iCp
z1fCgwySpot9iIDkZkGKbFax7cY7Io7qq7MRecjioqiuUdO3U/iThbGHRHNw3qe5sHNVjnNH/8VL
OPb/esyUb7QsauTWaiGZOVZn+Wa46n3obN+icyfpaVHmBT31DJuG8waZiE73AWcXd7SF04XmXlAt
rYWyzVYWRGJqBWtN7jQDZTd+/lsev6DQ9jo6itE93NDBJ0MFOU68S5dZSSuhlLPeagPgvHWM9TJz
EVr5G9QQ+0INyI/8TL1sscVsAXYNPwIsmmx1RPtGrqXsmRqFs8KPEFmEvPJzYp3fFJ43qwibvt9H
Aj15aImGFyQewnyWVnCv2D78JENOcjLswwSA1qDCP0l/EgD8KFty2eld9qWM2sjXyBt2kI6BbL15
/qmyT5MkW82czsWA5LeFM/XGlK7GuwlMpEgqsPicCra5rYDvdERi4FLvWhh5GqFMcE0idw9XLDNR
U34RSiEt8hZEWZ09h7OVnKGHfBxgahmCj4ugfFbuW6fAvXwQKE0wOGI5VTrPUihihtNhuHD9Goyg
F4QwrqgJyq/m6ohRn7ggXg89gXXXdsBTCLvfmAd2+s9XSja8IMlDsUkEx8LRZ12omUAfoHqthj2V
TSTlnkFN3bJpCwLDWWcMq+ZLqWhxRcDmpiHnlX+2kZfAr/Du0jAqJQRre2kTtEm1lbprHVSU47IK
x4jIMptxdybXRAbx9AbiIJCgiChYr0/N4rCB347iRjTa+gS6wtRPdduwy5QSlir+Tko0Xi+aKXqs
aOeY6OBGnPDOcjTcMe2YYFeWoqBuTVHtmvXVf4XKl1Nty0H114i15os3SQsi/7fiHQSYDmFE9lXZ
pYi+jApwshS8/vrAunLngwc44WFDbIR4oZ1opLylPAcsXwPDxI7WUsSJzpYsbIwD75vtRGBrMKB2
7ijg+3BLZCLdCx2AwB4YCpvc5rBsq5Ex8fnclmIPQ2VPiUGfAFol3vTwMW3loOK52dcCGjaM/XHM
9PbeV8uasQGy67G+G076zv6NHrJ8BoMLPYJFS7ZKPnAgFskEqiMV/0nwPMJ54eeQEJK9K5gOhd7/
eURmZ3T1dZqK/FEgyL/k5dtaKXZAOzHq0WPUclzAmr/DtSZA/gojxRAMtXXMCpPqpP0R1+ugClBG
cWj8fz2cc5qXpFH7qGNS6dBIACeICSnHkmf6SF2USyLowKhdE7lm4LQaau4fW432xjkmlmtdAHtc
njH4EmUb2J9/OYetF0AQjcNJwEQRlzhsVrbSYiPchIqUjW7yxRA1Z75fDavZMpf6p/vBs2Ps3msR
LgTojKgCMrkYRkmOL6Ms2VgdAe5mUMhZznxOCnOv1Z03daQ/TP1BWOeB58dUgKiWMfBA8MMVJr0W
Jvch0XZKXAUqg3N1dQ44UUYl6bDEY208w1HrRft/sFGnuAenZLIj3frFhqIOmaR/RgoXzuYkichD
nC2AlIRW3kDnC8nfPRBgHdzlpVNO4H8uwIPMekGzAyd7RlrSXh2VOSlT0QtWPVHJo0o+Szrth6Sn
EruoFj0urORKVqdQWnqYS+6wL65CWq12YIufhSc3qpWV4s7t6ojtK9gp4uz7aNvbJg7o2Nb91p7c
GT+lxNvMpnz//ApeBmNh7nnRH/sPaEwLRapX0OzMAulparf/BzDitn0Vm5BA3pluxKhsgaObgt4a
FhOCFJMn2Qb+hC8phhqMxlZkyUw1aEp8ZRyos9c+Noai0DDA/xF/YAuKE3RXaKB1e0zbobQ3vVjQ
N2fUljHmhb0sIKjOdN1ynvrXAx6SRP9pAdJYtTYPPAeJeQ+46j4iMV/Ky/lfhx+EEIqciIedtVsR
T+BCToM6wkZ/RjVDIDRh5so71i+GeYPCQ+4Tw/Ovpsl4QwQO9hLr0IWwhTuRaKHx9hRBmQ0M/27P
t5jFZWgwG6C8qXc+hmkG/RMaRmgNEQrxRAHzr+sNNcp1MncwW9R7l4g8u7UaPYkfGolnqIQL6zFo
kP3UBDT3FwFZZhiEHtJhNvSu8I1R0Hi5zvwOzObS9zsXlZhaQAlYLwa8ZebXsS3snrYAa2Szhm8i
yxAG4yzGnkAV8fKKj4eQ4LLoTYteK2xfBTJMhOzUVW7vMh44bYxzYc4k20/HxsRNX/GYJcfSYksm
typR80k5E4TPTElT9cu/839S9v8xagG3K+Bj0b9WzKYnyEphknm6ufrDC8DU5HdSPfTPSuIbG7Xg
+nVTwg1Pev76nGiINjbEkZZlMu8K5tv/NFmOQsUXixluR1i8Zeu1KnBj4l7L/qNoJMkcxf7JxgBG
+N6vARH5x17FbQcxpR9uN33cYmWckUjIRhvA33XB3tywkpNm39NYj0+IRJWdkvvHJG75KJq6txY8
JbD4gVU6+EeOykQ2/zkulvrVlHxgYiRc64FY0qVt3xRXsPrGTED2Z5Vw38cQEJyStIwooKDMEGBT
D+f4WWTbc83BsM+cIPQWTdQgD43kfsnKvVa5wj7Gb+9EWpmj7Zl8AWC+bG7aqeN8UK4DdhNl3JC6
mwc16o63Ap4zcTqebYIhAbqx2wjs4BcJ8NE6eTVEnShXCQYL6K7QdtNYuEIq7g7LE577PuBmaBD2
4/hZtITTPFstqfPRRrJ0R2npcjHJrlIHo/FBzK6NrgwKY9HrfUoaK1VfavxM1A1jpJNO6gQGu4IM
Uw9AnOBaAe6FRkrTOst/aFzT/T3bE7WfGTFHs8uVSuSQW6WlxPgDIMqfItcIQSPlQQNgtnk3ssoG
jxYB4PIXL1QJsHYmVgyQhLtGev86YHHYmrq0+JNIX9j7KGrxpN+Z9hhEQ96TcR/hxhoR4Byv82XK
Opw0Udj3MjRixMT+x1JA+Efovv/X7+1i+cX8GbJKzuWm2amfqj5OkBjATnryLEQDpzwd5pRXCS+a
Gv3bydmChjNyNVXJrQav8VMveioc3mv1HbMQogMWkNDnqM8moNHgnmep9+av6f6F1jIgVtyi7s34
hEWJ/+A45eD+Z+cMTsCH6lKS6nJVT4+116rVmqtxHx8RQWLx/v6HUt4/eODtHp23xc3+uBF4rKtn
9kz5Zf5K6AudCi2kMoBTr+K3HbktuKsO3mpqkSGkV9deHteT32/O3L0O5JCZD+N4mGE+bEbnr9ON
P9vi+A7tIUk7fuBTefuyl2X316SQDcKv+pSCn+IL+jkmyBvVtMQUyj4DZ5lEtag+J6Hu5dUEWVGY
VnyfE9OOIexwBBOeubse8oZrI0Tq9FQKrm4l2CjPV1z/AI6al3liFDrKRzn0oPhObqUcOB7/v27k
uoEvk68PMI9pKzc4hki0qaFL13c2D4XesVIzIkIcWEY2iMdhq/o+V+liU2MAy9aufwp6UzdIwhOP
MwTLIHxlaufHhEVQauxfomF8G7cWMpW1vYjfsUqtCjYoyjFttii3UFtRObehA4u8xpzZ4sfsjPV4
l56N6wrNFNWpZeP2Pw5mYSpm75e9qYhuH/9Ez+YWvUINyb2mBXkL2bg84331vxvjVSuWXsZL2paZ
vwTES0UQ49mHOV5/4NqPkF4/pblOZlX9ZkEbIgbMq7UWie+egsuL1olWFmh5q6kAgUb7bFkGQYgp
3nIZ/Vh+GsA84L+BhaZiIvNNQiDHjSjg5zqrex/rhKScRjBx5gXqhnHNAEZhjYQKxClha1rWA9QF
gif6cM9EbfPgxvLizhGcwShsI4CRN1Z1yWgRWbE0WwSXZcSJCvLAiRYUURUBFfydjjj3cpuUqWIf
R89KqGM/ZOi9ZlED6SKnq5HhFIOsTUlk8/uX5B2znVJ4xlpZX48ION0EdMeSrv/aYZLgmsop8aGt
EOMDEINKGd0PLmuAAwEm9pkA3/+gw7Rf19EGBvkbykrk0sIShhbZfjgZwfrVPjxLIHi0holwjyTS
bm0r7eBec5SvKYAygoq+aIs6HQgemg/8hwn1DR6Wg2iVQyTKYAHAN3DV9paMj9tN4fZ41raU8nhH
JqBdy5UovNy+A9SiwHRA7JOA34VLwM3Yv5aFLJej+2j5+tlUjRJgyLqJ/9dPBjEMPkg9ljiSc6ek
Wv3SxCopSL+S0muobhzJs61UT+scxL4qaDBC4iHivXEpF2SuDM1nTAsdls0gJryMStl4Av3TGaPj
XTFNSltnsMSfryiSF8/Ji4v7KQxsckKSgGvYdxX2T8v8Bvtfxp4gPCFA5Oa7zG37ECzNVHM0hiD1
PFuJeCgDiMcAxT7cE23+mXKBphjJkOeJi7Hz3AjnB5YdUQylM9uSSaBR5sqf+9i+chmy8tPeZq7Q
bblV+k09mBdw0TiUHYtpnaLcO7eMG1x1IBQ6jWWK9Ed4h+s25HtbJMqAarzgIipiewgIM3FBLIus
cLxB8jvFYsP+xcPdqGL9geqlDB1+zkXoktgsQI+siJdhCBAKQtS4fRgCAwkofVodPQFOp/W5h+5C
gTVHxDfORnc2RE/OYroANx/2BLEeMjRjp8TQ7Fth0j7q5NXcdI7WZ9s0tmBEzZqfzUMQMLHRcBNs
fINdRC/AOVeFX4D0nrmFSDoomW7nAWhAeZVbYTFSAHK4NyDHjiucgkdDTjy/mSqqYoRLOFaDyWAs
meDBLXR/SW+3Gj4VJ1byid8l6WxDPa0uMdhMoDnUTQHIduTpo5zmzNTtVKGfS2wTjqKTIazsGIYM
9T096Ezzzb3y6+lr8Q+YnqXWxnLZARzD20a4UFel/NAlv7nB8Bv/WuOAXUPYS+u6mov1prUs0m88
mFxqIS2hdz3EQf/s1lbA6Nmieq32KX8GG2/cuQ/7w3zvz1qzrctvQRLPrl7Xyg9KVqkShNppxJFn
JFfcTaKly/J0JTctoGBs1E27XpgKUmoaA7xMGYrlu3nBcGOBV7GftPv2rmCU6UfaWqEGsKsktE2a
boD1v3H++2nOM2E8o+jt23OiZ1MFIrw37cr4I6CvkwEd6AgbwabpQ2WwjnvWbkJ7muyKhI6QJBcX
mo+ydkQEdh2NHgz5d60dC0I2pAxVfQDCGrcJ7ve9tyongjZPcENyyEGxS1Twm+sA+KrAurv0RFbX
fRQItiyYmBszczVuy7XuN1WTvP2ePxIm1+8dhSAd0VQtzsT92W9mDwFLwFIbmfko9TnKEoBapE6A
mLxK/eaCGBj9ZGDsZMqGrw6skEN2X0uf3n2K8VChvW9cMfcBuZjzOSo+ym/xVcTOR6GsanGZTb+m
dYdej4KJ5daG6VttIE4ceWFRMlwZv5D0uBFdA6D8kJlNakhTZyvxAlbkoFduY6NH6iTnPMR+Hrl4
kFXAz1VtQ3bnpWVIRmmqjWlMpWnTvMR28h5KPmyWRMs/1ZepzlcGnojRs2OibwDKXEi20tvW817k
8zYxX3j3MonQCcRC+W6bwhmYJdQZEIKKmg9P3muEEV/zh37OBq181GwnjxlziZOwnyKAZhu4YCeQ
E0CkJYIxpKYe6rS0zhc1nA+aIVBmLelMFzyyf0EDfnWZZEQ5QLyqX816mJFlUPjaFPR3RigRKD/M
lY0BgkGCAb7yAw19+j6FZRhtFfqQEh80PIt4EGx/yAeOlUT+q4WcGT6fKS4In6NcKp/AgbY5J3Fv
itFQcOWtTcJPrDizZiJd0CGdaSfyXdGIvtjzRDsvIgh8eE/o3tfkzqzyfolJvphZvcmDFgz1rG2t
Rfko5Kf+zywlfc84DZkSPM3bJtvYBvU0ftdTq3e5wqiQMIMTsXQ1SbNTqKcvn4gBPEE+1lrn6BXK
tS8jnp3UdB3OfLeys+VAImiX7wEMegQFXcuTDo2U5ypXWFOYTJKNMP5gEGolaZcoAqWv+EhASsyZ
Xm0FDKh61hnF+JCy1zhrO7RUH86+8GdqUrQBdNSqEFNwrdzLT1B0happvwkToPoRCugyQowKnC4q
3fpDXj1TGDRtnhQtYTF9ZAReh7F7gUayf5nfs9J1u5gjpIEoDYfYdm1lPMs2+vTgHDg3dOcW8a7D
UqA2N8Ox2ubi7Ryqv8v/UG8gXsTozo9o+Q5mGeBt59XofkEiFMirlCQX+uFSLUPBcMmmpBX//AnB
MjL6QijQADIg5xvTBYqDsqUnzvQFoj345xtb0R11ZZb9ZfkSK4sqWhOE9GOLYXGam261+a1ssiPO
TvbZgxzCJrk9SewRnZrKrbGQzZRdC25umed3LMZKmTwVyEWIn70wOAc4SiOueQgvhPYImMtYdWm2
oKllkJfgkUXBpKgvNXPKXMCB1p/G6wm5xkBaWbqq1btfC7vyWLmjUiAxhHVIMKzRBcg3fB77JmQ9
atnV9o2m4KMvMR/HRRdARtFUQs1kNqQahexwnd2q5BbesZr2PJYlmP3dHxhx0HYoIziTFxnxoNrU
JJkI+ES0jjI2lh0ayuv/8kyltkKjG5VWMWrrF905WFGD+E6UooI34T1qTXrktHkgd4jr9+A2sFyV
MBB/HqxBlSP+q9uNfrAEPb1tSfOkpeSRyM6V0FzzlBmdFf5uK+4N9RXudKxDopBFuWe3ri6WmRoS
BZMc61GVvaxAC9O2eb+uWWTwZWjXdjQoeRO0NQ3mMszUHM+oMegGvCE/K1kroYsQwbi9JIAmE9//
ff5TBFEUq/rByzWdv0WrFgVajk6GJCm0TYu4E4ERkKYLvt+/+tGwffpzIAWrH3Xr9M35wQh2Fpnp
buvBq4ST4D4gw0IPxoeaA1mdniOnvaBK+0HTZCAIW24qGD7bHFw3c002iu1tWKuGxeMON92IH1Pf
ip+XFAqCTZ37DREeVxQoBM8DarzDR/ELpFMko84MR/hN/nyuhPsohx/L9nS8tvPLMv9Oo1UKbBp4
TFx5PBli3j3t3o4ZaQPaHSQWNxy2LqQJTX4LfSnA/JpLl7U4jDvQo+BeRIWtrfpxj+8B6pm8kFr8
wq5GFq6Iv/i7GRV020ghEM7BpB8Vzm1+tTrLig3vQwi5u+EqMUDApIIAYOegxIjtGH7C+CYyFbYX
8Q/MYwvP9GGJ+fGHr58fZjFP2xw+uiYcybHOcnbFnrb0h+VhzyVQRGj+xCU7hEuZY4mHEGSXg4Bk
QcD/2BlRjW66tN6Y8JhDlrwZMbn90TouopWc10pQkDOW9jmLHyXpoDVkj7z3kRtdQ2F/1nSsrMG2
0h6BOXDModt9frv5K6gSHHEal0sQld79/Gzbq9bgTBN8B9ny2my1RBkLV/fhoeRVWPK2f81CKl0Z
HB75kZ+F42KYlRCsUFN+TZQCHC6Zw5zsf0arMFCidmOB7jG6gHxRKx21ejVQYzNzioJckcXFLGF1
EhUwR4p7pyuOs/0La/27gSpLnG/iQ3N/WQsX6h8eiTbyCmsuVqjq6bc5Hzgs80jlzvgVLisV7h8y
a7HftJ5aU5jXPjN/NEdJ8jh326BEIRfSLi8fsP38QQiMu/q55UaMNsCgrCxNIAMSBjovxu4Rbxyb
KoEA5vewV7cqZIpnNvU5ZPi6xSeX/+sEkwN9Vt1BWiXO3GLyYaSnMldLozXFIgca20sjRdcOX0XX
wCv/hi/AlISF3qRU390VHb8hzTA8/x255CFOxwF5IVJoTB6CcnnJJofFvKBzJaK3uMXnCA+BQMcF
qKvYEFgRNGpdlxA+0vacVrTiYN/VXcnaF/G6Zf/vjg8DNXv8TBU0Q7wMJhOQ14Sxze7QeTf+OKWN
IeUE1Dt3Qz4CROtRQG5uGiXbK1jol4b3D04cRVdC0NmsVe4qH7/IEVYwsxip3yGmZOLfzZ1GGp5T
lGt+U0/o+uNXDp9X9PyM21lebDObl16kbJ6d8ld1i116UCgPa9VGUaBevlxb38JbbZ06voxLbAfB
D7rKNHCgogHxBIfpbmMS19kyntXLUbOQhhFO7qDU4NXbbDQqwykm90L3spaRcGSNxVZcEG7KACLG
yUTuuuEAp1oiS96bYK9vFPfx2wILg+9PQvSJVmINPIjxzWVWGxc7fFdi7Xe50BL5KxAU1d6myLvu
suo5HPE5Iq2AUKkFvKl9QtOaID0LkHDYHaUk+YOIQhXFxWj7hl0X76vvTV2brKoR8e4jl+2nnbC2
/lleUlkBIGjiM9o/m+qCh/k4hV99WwNbGcnQGKlpspfwirIafNRbiFgk4myW7BxBqmaVfbIeFfWd
1tsvhOvXAwfbkBRZ2KvUsX3OITSzvrf+w7hYoWuG5H5UGZUagxjM2rkY1GZxwQdw30SAUfqIsOYY
Xe903uO6VkwXIvDg5H4UoFLOwsxU54Za/hhvC1/P5UAoUm0OjtEMofhlE0R/5bYiQYIIqVGq1GeS
E15SwELPuxsP8RaEV3f/okLs3KmY4BJ3rpNhlRg9Sr061CayyDL90A7+cXwJeHT8QjKVqTV4awn0
F0krk8hCelpbSeo4+rrtYjSqaAqShA+cKhDnVyRCIQxYlyKii/SXJ9mXHqSODE1oIHeIz0+DTx+P
yboFFEiHaEkLN5qjZvqXzky+mMg33kctFjcobxXPNhaD1rlCxZnJe4pTR/uZ9B37P6EbOR51/Kdv
ZAoDzoR7Wg/dMDP+Du70X3g7GaEUjfnsfZBqwyTYn/gZEOVSF80SnTidjCo6+zhx1jnvnbAIfykv
4goehDnzshI1cz5YE8IS40CfIKgPv5B7Iw5K9P51FC3uyMYROfVdGFxB+WhXPgOr7H+Aywe0cJLN
hv79DrBjmHsyXG9JmnapedEGUpggLZiu7d6bEeKteehlUOiYTnqHueTIfd1YyM9UbPWkPd4LdR5f
46ezblyFd2kqLvKLZVlYlAAxIc5FRb4ZyWxz48mcTFVnzAUGolAUH7QH4Q6R+s0LPA8L/lOkJXA+
+m99VjsLR/yGot0a6AXYBQb8CuCityg9G6r/37q/E8pOvW+RwqEXK4XJfK9vXKSWdxLAiTFy7j/Y
9p8pgcNgHb66HfneHe0Pqwq10SnM28o3idpXT728C5udKXtbbBjjXt3WzrAXPS9B1Pdn1HXn9Bg5
IVbrO1aaewZzqKLrQXfMUUUeBGZHDbpVHyhIRXt4iFyPWSLcW5l4WKyxk4VuVHoCzzl68yFzUOYr
MTAxpjn53lmDnlx4v+dBZafuJEn+750LIgQwO6wDwkI+ZXEdVKTu9+8RUr70+ziUZldg9tcHpbyD
MNZMlgIrhH9dtmukzRfjzBH86+wjro6qusTdGACdFFdtGj7o8ckXBrc0aNsw5LA0zmnz1qWC1Fd1
WsxzmMfOljr/ctdFuX00RzwwMIaRIXJWWw9Gvu0Ph9pbS4AdPakSfUzogyTDaoa5KHB4nwwxMKp1
CKUdlHOF0HTFcuUXf5JdlYbL7UoHSQLg1f1Z3blH3MOydhROdaMNiVeqdorNLmx56yXH3E6ckd+V
NwdKXdaLDltA/Ae1NglijXBiWjFL5MlHjLuEqcLcPW4F7T7Hm8xmLDLYyOXtC1Bgxow79O9zJbct
bU6qdeTSJMgGlP6IH3eWbcKEq5LJwzJwMP0Xr6mTfJ8rHzDKYCLUrd4KEl3/9aue165Gg+73pDRC
C7PFXZI4lWCBDpugHL79B9L2FkBJsulX9/1tI5N+qMso9NBzxemBiCO+SO53tziKpQsGXfPrGoAC
6tl42K5JaoTeEyU4TudlR3GxQaFDD01rYZlVD8q7VpF2NmtDX2vOWUAscpVz7ZmxUNk2by3g1dmy
DYGxD5T4+xy1eHrDL9o8tKTVdIcSnZyT/ZCt2Z8V2oBkupaRRYaaJcdjHK7IonzPSlK+IgsictCI
OxjpJmqePG4RuR6wv72EhqBnZ+VsS0NwFxLm3jDF/n99OrrrET+8A9nndHR1eJxKLOW3jirr0iTn
E9rVlF1jeYINaUyIS7vdsAedvUt4Bi1pw8ZBJoYI8Cd2FvGtGr1T6Hi5r3XFEdn99MAW1c1OzLxn
4hSHrS0AN3nnxD1b5QJlZzE9Ee35LF4qGBVAoAlr7djzVfJWALiqkMHLldzQWh/hruPxDP4UiR7K
3/Q4zg/2QzdOzdHZQGbe+TwHHO4Vd+8WM6EVRdE4KsmHyGrnTMm4kP3UQb+/Fyrkd7ObRY9frD3N
+3iWjSJ826mWBXfw10OqCOSal9mNgLuOHAv8wLfOntE7ZR3OW1c7ZfjNBdXfDUPq7Z2Pd1OlKh8O
fQg8rClfYoGzWXbo1SiIZken0a35VOrI7OZqYGcp2bO6a2opU2hMr2WPNsNVwcxzbaeKWAf7c26l
NKmAms5LtXQRdgLd/5G9YbJX2nn76cszFZk6S3/9bTX6fQEdlML0VvBlsXP0yzqohY2A+a24J5oZ
mk0ATzwTZ6nIm12ccx2uqSXiJ4iA+p/eQoekBuWzB9hWvg68jiOt+1DXD/VgeDU2CLDbtMmejFVk
0KvLaFiIt0hkhTO72ntlArZ1PsiJnSybT57tRWUj0pti83M0mcWN0qV5RCzHYQJ09VAj5iPeMrPE
Ltxg3DArEwOTLj/ee+tMI7mOr97hs0uD4FZG1C1iFyZQ0BB0fSyO5zfREhjdyslxrTDtn5UTtiIe
lSKotRH47lb+ZcORl9ItuvDCNyPFQqy6Zb+pYjf1AUZGSrG/5M/bNbr0HCr81FhFbeRZhAHmcD8b
HabkMHuMniN/t0RfWOAmqp0mmhesTqONajtDy1/MSHcLhG2P8l9T9bBlFS+o5EBvMviBFqHyp9Ux
a6vM7ZfeTUKvCDaJlILBsrAAeqMTW/Niyr3jdpL5Golsjg62ZsbHVii32HMITZEM3S1fb4Fz+Bny
ptZUdE94YgRBXSAjAjU2bJDafdDK1wrZM+zH9TDvdYds88XCV+0/ugI3LnEb7L9BFDcqekBBC2Fu
eQNEAskj0PtRKG31LPHN115DqX+IQEB6KixaK1t1uBSo5a1rmIUubUg7jPdGJ069iXJBfk1YlSVg
KROzkrJbZqlXrIa4g2au0i6/BHHyKJjnKRx3wNn0j1geJubXMU4l3izFQ9/3tyW07tozhxTbfZ6L
76va6unB6gU8tm0PYiENUr4ffqXPRY3gQ+7lr64httX+NzIQMt+9hAKPCdCR/p+CTESunCSpu3kY
OI9DNjgvxNS/pOGGBXymQYLeB15k1uyAj54N7OUbMoGx96ACzDbmtQigWfwDu3ATaAD+ptZnq5us
eayYSs4b/iS+cDLManX5vle4rQK1U4q6K560SpZeXaEpn0WxMQiLkFXVNKP8NqD7EI8rJcmrWaSZ
Yh9wMwJniqPCYPesa7RkGVleEKrXX6fKk1bOgl35PbzY/9V4gedJL7UtZTobEbKsJf5ArYK2sbRQ
0dfw4BPWl7+CHz3vm8px0bbKXLiReuUD50LrY5nwE+tZByofKhmpq6QCmSLU1p7aTCvei5hgPl0f
HyRlQXCin6s53h8MOekOJPvHAjfCdx+r2MBlNgDQdY1r6M1cuiHieW1iKNLNFnJx5z27KUAyVx3q
yFph78GHUwYYK/Ocd9BUTE2nCNkgr0McwQGRz5/Pgs3i2YVzsS2E9dj3Wp+SBf7C9oyyk14es+ck
F9vZsEOt/XIH+DnAaMh3psy7+y3XnGJZMsnfo64F2dlu98ksUf07+dPszCf4e3D/cTSA5y8+5WAi
DuJpTuw2m1gvLIS+lQZzMXypjxnA42+oV49DCCsl+IY3y8ojeVl5HSj0NDwQ7XcAI28FtYMfRr4s
MTjVdxvhqwgFAkHUFxxU57hrjXlkEEoG9U/9bSLyQ+tS+fWrO4sNjz/S02vm+mEzxJ99dHFGxAEY
rtYxscWqHphxYA+JPCK2wP5ykpulTv6H/dxepFK470gjDExN9DRkfEcFh8StEEIyJw3fzh0jjnWH
RlXKe+IM9GTwA2wERhPQ+HBIJrcfnlCuOPhGweNm9DVeAXZbk0HWBHAE/8Wza6jrgd6e9VllEDVu
59/SWjWSVR9UmsmNU6O/Z4r3OAuzgY6NjgoNRJx+TqJai+6dtU9pWQva4ixMucFwrj99lTdm/FuV
uA69+y8PmEZC/OToWTzs+TrJ1uiLYXVlcYETsap68Q9ipCRa88ZkiV1tLR9WqYX0+Ygn2OrFz3Ph
78ayEROYm0YbHSSRFUAr7pZy20CJFsn79D3j+hKxPu4BRgsRLCGfaiN0BY32LyDs9ZrJhcKBI0Lu
ccp4fEcyMKz15n+FYNZMID9XGhRKy2VIetno6ZOnzj6nds/TSJPU1kzCVhlkvWtTpXH+KNmI2Ad6
8C89seh1sVjtnDF9v8KcFUZPQeKeg1UGiuIzCx53HINp87a66B9Rasf8FCMe6glAR4lUJHnSgPYx
chL7WvhQcXYmaq/fDI2FNkkIymmmB2kji2nn8zwDstF3ay9XNC+NVoCB4qAFqWr7bllbIxIhYORW
2PmMuDvnxSshE+TyB1RhhrJaEbWvCz+9S990v+9v12y/VkQI84LlEIidXuSNOn0D6Fd5rEespdDk
k7Qq9Mz/vkeBqPXjlKT0QsAvmMfEkm/V88WLjcmZoYcsavAo48ykGCXkgwe9i5gToUsCcaCeaDiA
X+AlGE0Nul2VHFo30wMM0ngay62KJY2ogIfu4riZA2DNar1vrz649pIoMOb/SfwAhce5IOnRtqsZ
aqFPGkNASL+wgYU6YDAwra+f0JqBJapcBo1uds5yzbL68+DzQPoNit2rAKQHbRY1rzKlB4W4McDk
/A5xWsJ8MwGIqd/wfELQAGJTfFze/hQPXDIQezl7XDl+S1DQCJAqq7xJJ/XgUC1wGNk95/m3j5z9
lmX2dkRkwu1eMGSW79lfVZRv5PxHHqK2F1aa+iNika5sjN4mBRv7fjpIH1bskEm6HGcUAy3yWIw3
bpYNwdpHUZkcwUANWwjbE/4WNqLMucHiv20pvzSTEFg80uOqAEl+td+qbqTKxXxWgFOSqTzK7fEq
odMnmA4RIWG0zvTJ6YxCe0edEUsR87yBEyyygaD02f6WBYKtgfh5s1SiYLndDqaxEb+tseQNIx+M
fGKMM63jqFM01D0szF1wWng63I6cGim7EFyueJsFwwci47DbCTO2fGlX/SLhrv6lUrDEmtuSxajI
OQFEElopooTqAbKki1bmU20F8ZEqhYkSgj5tssz2Rm6IfTElnin5Stwl0JGNTd0kQFBYDWO3+a+q
ZzlEGfPApgD12mNg7frR88ZomUvuracpOD7EaGM1EbM/CbEAr26WGjFRlPWFtcHFsXi7f1Gtlf7k
8ifvwqgFfX/b0TPcdQBIcJBfPQxfcucaWwTzlxcQlRsyd7Fi/s7fG6xOFsXrFneuTgcs4NhDfPA+
y5aNGbavMZXCWYtrdt+d1qcYj0BPlTeaq0z/K+xEUNwjimjJQmlNuiO2K3tmRZO5EXbcNqtoxj0n
nVHEB5LRddcZf9LPTM7ehiKM9ObLuC35QY59ENiRjsn1L0Watz9wBOoKsSz32ozBtjzoId6uffRx
cQLO1mUHNOGNRi1PJ2jKmSlvJ1hED62p9r6+KjymuZFg4aHUAGSIBD9wenkXY5PIRbblPfbIsOmd
+eZk/hPnXhAKqhP/sCpdIAnU18Q6kAYKYwkKRN/A5yo/W0Ttz3mm3MmSU06C8GJ+QsC9AMpMNA54
f3p7yvoeUQf01jYVJ0kQS00B3PmoDgQq+TOe7DCb5t4qbS6Uj1udgJDSqb7NMp7nri3aSssmZIEY
txHz2U8je7BE8jQcJQHPH+Mz4GH4mfc+6Mgy7WQ9cFDpFRPd4DjeWw7INFhY/UsfrmLAQvAE5AoQ
5gWBOOouXIuVpHY7nGwWmzTN9dh2NUc43yUyXzp+6mf/905ioe8xhURc6HEgXwZYC44Rwa4Mle85
f1OxVbPSy2QmhS1hjFvoYstRJ2BQle9eGF6bKhC1isU2X9C1EZZsFE2XTqFB6Mw3AjDQ4DRwytJm
VFWXUODM8a9BdfyvatbAUE7GGfbwmkrKFUNJsAXV6lrC2XsUSoK/KYRKBHSuhiygtClRj5s68uKh
8o/d4ZdNFvKwzQ1QiVbl+bU+G1cIwKkKIg+WovkSaLCFvbVKmsxMntNESrN/5k4YfXAjUMEpu9tI
z76IO31wkdMnv0yCZL3ueclxHQcBQUcBS3XPmvb16HFC1RidBW7GDRL5jjxEqQ58D5/eZxlk48aP
+P9sWZGpvJR1AA10lBCddt2Ap5cu2dPpJhMKo7gx/6HtqukivbGeDx+yHR5lFF2wMbG9skrJiaxb
t0CK4KBtxYmjtI78V/W5lgaGROLwvaYGnw6hKAhFI+R2VGi3SxRXNre1rkw61ShnNxPmyPF5guq3
yxWBHopSqF3sXnBAv9ptbAe1Kp10GOrQPcCGD6lxKor9ymC8pPPMBnTtP79soAaG1U+w+jB9O00q
EU0cc1OlSgeQmrEZZecqKrQfzdpNF/FHMZMr+2p380JbhAt9hgsfGvaa25mMkGNA5PUBX9vnuxCC
1xPu0C+F7QxIl8QW/YKiT5ic44/tyvcQwquKNJD91BVWFfOTAvC1AgkZe8DLOSZ5+yHlr/pJOfUj
t4nQcqCbSwUwxLZ+bRyXOMUHsIb+x3AgWi7gzvGb/XhlxM8TUpwPZ29qoq7JL0odsnwwiwKfhSsT
GkffVDahLtUXYs9LbsJeMNFAmRws7cMlIgRxsNoqEUPt/fR9DBljTHgtS/9YtsIqYLlt4fFflp9g
sZauWxZYKLwMh8hYtq+1th44GyWHRTp6zrYkMQnd4OY8sMkmquV+/Mn7a6T2NhoIV8dTqNo+DdmE
aa26xZ5T+HF72G+tBE1w5JYJ7h2Ksny7AiOrS67hCfSN0j+Vh45CvnynMJsYv00D6pWg5T0Mm2AP
6W/A3VazP7GQIeaKD96bg15rbCItAztEQmLyCMvmMRwhsxG/GlwDLaDEHE/5w62+fjnMLymp5zoa
09kx4scSIKP3C3OHWsk77eGNtEspd0mPjYliTaWihbmaFgSYbIjgskMrfyD6Mw2Psvum7LoLG2wk
zyelQMR7JzMwxUA+6Nyrj6OHF8qUtdaomoQKTGEMPiMrm4Rv73Fg1i8LhdHzYdUaOUdQKY+QZbSa
SVyqaUYp6IVUR9Yf2PUw6mMgp/BHsiUS8aWTcUk4HE1mK6+ciWTgAFs3hFjrKKfjN6K+ke8UgI0S
uKOvnJpaZMseLf9FfSvcOchsxEWE0sGxxF7Q8YKN5msOHmRz/hYcXJEYgavgw/VAHsiaD+zT1p+j
MIH34OCvZ6sd0kK+2THAz5c9rNKc321PVC/y0ghNXFJWmsh9p2X0Zo8bigm5lQP3AQWZc9M4Guao
Q6i1Q/vxab8con68qfni6sPv2gMiffgDnLKGtz0HuVlbGQaPs1ih6G0hAh+oRbPxuDnLJwWZxmcZ
HY8VbTQ7IIGIbdGIGz5tZ4aI7EAnS93l+018kmcBGgLWsXVSoGwztKiN/llEh7/IHOAIJlNucBjO
wYHaNS0svZOr/l2VqusoWIyTofSJylAhvJThXjBJduIRFbTNbMtE1/wocaweOwnVFqllpIFPL+2n
zs6TXYV3SJhV2QbM2tb/3LCmGdLeJX7xr64upJU2UkPrMRhfMgoFbUCw9jzdWPWGHSQl/xUCbMM3
dMuFrhHrsvWuMAPd6IjUVb6EmdZYS1cKmBFUxxKI2enCL6T4KSesaVWPUYtDURWyXz0ROn5FEO1p
MkKXvDI4z5QFfu/BLjJ3a5rEA3fCXXMjLwHiX6z/PP8UZfL7CUAM/37q5cXTwExtxcvLdbAP+t8W
WBMPdgw1rD21DdR1IWUGtoDD9QRt7Dgbj45VGYa1HdW+/9cbKK74xF8KEFyn5DGNCJyORCkg9YXy
lrv4MtBk8oz3SkWmyw8w3Hw4A6HbPuOWYKafrTPGb9Q+VqUkXNEECGlovqPAapkzoBSMni0B7jHB
WR4Z/P3ZsZHKA3a5cZA8EsSJYpBD0tbmdZSpH83COrFpRXyxVKMWiqG6VVkSQsZ93sqnWIz7QNRH
wGZ+w2OfagqbJIbRf04/PVrXgdwFnYZkvVszd36gK2v+on3wfBNs0fVX7zsh2rKVcPAnMjwExOlt
JrxcFo2/Nm9grH3yK89N1XPj7GAyZQfX1NVNLq3gS2UtX7SvQ1WrfYfc4VrWpqD7FrtsV1JtDsHc
TZ9NthQ23OBMfnyqHpsvEchsZz6FzBl9QTq96Y3iULYO35vSYl/C/nV/rybLgeVyzVgt/DjunIqR
sMWIMdCL790C7LhPevUuos9G0z/RAiD+W9ZvHZo+kOZLw1dnpo3ZWbX97Pv7cJiwfwU3XkfHyr2s
UD7NL4kSV2h4mSVAN+hY0Zo+vSjKNxqbdoZEyvdOHM1MgSV1qT8p25+kR1uLuFsnmcPx5PK4mAdx
K0XijjrkGu++e3lysCSueTJkecwmsiGmFjo9fdwSyBnAZjL2vupJztAyHo4pQL4l93Zj8Zh9WVh9
YPN+zObGfjiNZSU3SO46yz/E3dW+VJlpXqnBrhGHnUOhwcOPicb2tcjjr/gQAtpm8fReMW0iJYa1
as4rnkUq7vVuD5Rn8bAYDBQnEWX/0NpMwBI05TTHEOCdxJK5mJiZGX5SmAtyuRcCZof+6MllpkS3
UIGW46DI4cyRL3vJ4n6eWMDnfAT4I3vxN64rIDhVazb3i2IXZbsb73LAM4bW3tTOQZPqf7aNSytU
yCrL+pSkwDZCbs1UXUyE2rvevw6m2gRGjFFAa9RYFjhgVQEssqA7rPseafFEhHfDuox1/GrOBV8r
MxprBaIKLGdseDU5g0cZA62yM2UxKS4=
`protect end_protected
