��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�vl�5�X=Fľi�aX��3j�*�uj�G��;MH�x�{?U�i����,B��a�s�(�1˪��@*I�[�M �#��ɪQ�${�:<:�����k+"��B����-�������#n�n
��հ8ҝFD�Q����Nr����"��*vUٴA$�/�u��mH��
NlJ�M�:�Fi��1PGdסg���/�Q�uV �a���䝚�0^$���<�uNzb�+j85a���5}����ӼN*
��CPd�� �L	+�S t�<�Z�Y�̎�=��K���6�[?fg	{_�ĝD���J��A�q��d3�3=]F\�U>� ��(���oҨ`Im�e0�!�X��;�K�W�u�_�/�憬����t '/i��h��P��?��G�L�Mmw�p����H��E���o��u-��}͍�v&zxbj{
\�L�	[��>*�̬`��f�r3SI�,D�u�q,Ϭ$�,�����!�F�ca+�P�o�H���ȶ��zˤ7 8*EC�!�)q��v٨�D��[ ��G�*�3�C��+�3'�vw��:�(���kfQR�dUZ�9Y,��r��u�"EZ2\kV�%[rM)NH�lI;�d��8i�ĸ"��洱u��xc�n$�2�/�GV$��y*�TT=}�aJ%��)�<1A�b2���Vb�O�M�f�)��ҹ��2���)D�%�ݢ(���ȄT���l4�v�⹛�Ǵ��o��[( &��
8�^���Y�
�c�����>t�%�M0CL�&�K����^�_����� !:`�-g17<c�K�a���2k��F�D�!*�����
�m����`�T��X<?@Ϳđd���&^zp���έ��Z'������aZp�k�|�ݘW�y�U��\:%_y�q�ҠU6f5y�y7�S��n���2?1_�y��� �8Ϯ|Q:|�o��h[k�_���'�(c�wx <H�����i���pF��H*(�'zP'�h�����I��fSRǤR6P�=M-B<R�@ӟ�������a�/^؄�Xd(3�rx#�5�a�=�jG�����!�	����;��b{�-
��~Gx����Ə��ɝrS�)������O�f���3���Wж���o�'��uh�#ޭ�`�;)�7KJ=�w�zo�E�����x�Z�|�A}3�g�ûS��:��PY^®l�1ܘ�.�����?^Z#�H�5X�2ݔ�3T�%W�
��q�	�z'E������<
�{�Kn���4��ݮ=�f���yb+0�]g"|��G�Ŧ@�<4�h�����
#\>�q�Aq	!+�,�S�����!1����k��W����{C!��$:����a`�=�Qh��]_M��P�`B��6������7Q�SuT+!�&6���V�eJa�(�<�(o_�qV<�8ƹ4�ZZ�M����_ܗ�iX�tP�neǙ06p{U3Oz���oS&b��d�]x:ֿkZ�+2�߶��t�9k�vxÛ��(1���_G�3KOeҖ�ǼANdZ��_��?��X k\�'^����E�>A�I��/�〚��w�r�ߘô�u��3��i�ퟀ�������,��}*�� ��=�S��ֆ�b`c��(ׁ��Wu�e-w�y����X��e��X(d��`�Y���3t��r��*܆u���n֘�6c�0�	�4ԗ��-��u�����e�V��'�4s�	�Od:��'�K�� ��?�Y~ϛ��噔��éœ:�����[�t"bx�{]�ȝj�ɼ4�#�U J[1a�����|��nZҨ_����l�$�'ؗf`<�{w�T��Tx(���B0/A��^��h�����
Q�*!�Zhx��k�
0�g,8�����~`���^J
ր�Ɣ�� SP4�N>�,*:F%�t�'��D�a<�f,a=�������|
b-��M��Y��mLU��8����d���n3��m�M][������ȡ[$W��L� ���Ɂ��L�Ii�^LE�S)�kp7�m�"��k<�����%�8V=�f'p�����m%Y��ǽ��Z=:��%=!m��I�0kr��h/�Xâ���&��6����}�:��X��1��Q��`�ol���1���0Tq}9���������T��|}u�zo�a$�c�]|������7~v��׀�[	�h�����W[�X���TW|��|�c�@� �1#��3?�)�1����Cᨃ�%��C�3A��(�S�����X~��?�����D;[&ӡ=Zx򞌫t��π�l��<P��pK<��eԆ��A([P���Ũ;gV���\n��>���!�ɚ{��'���>��C�B��1'�1��#�L��x�bޑi킶Z��:'�dW~�4��ed�Bdτ�,;�hw�����]�V�&���L-��R��@��e�iR�6�p���^q�ƇF�n�nsˠ�zY���M�@Z[^]P
W��(�z�=3�0b3?��CBߋ�1��䩕�A	<�z�Ԧa���/2���!�C�8ý���y�x�8���lxW���*{�����ɨ|u���E�J%��;������w�beB��`�_rb�j�l��c�ݠ�\�e�}�����9�e����p��	�k��e�}�>d	�z?�`ϋ)�]�%�ӧ΋g�B��t�<hsO��͆���;����#�?Dܬ�ԁ���csZ�>	FQ;'�/Z6tl������U(�ݪU�t�Z�/Q����#����~��:%��3�&�zt֤�v���&��8i�x��M�@WҚ�^؍���wy�^"K[5�}�)�a�T�-OY�U�vR��
�}�@㝄C�h��	K���dP�X2a�fhj��(�ϟ{R��歠r04;�2f�PE��{�9���hK��5|0|�˦��0=Q����5��7'^#14m��+�E���"b+g�P��WPyZ��D\C����B.z=��3�.I�%��b�2յ�k��z�GC\e�(*�.x:O@1�"���ϸ�$��4C��D��lb$$�-ȝʜ1y_�-<�*�8(��X'�1)SDR�P�(�a����0��X�Kߧ�3���<�}�:c��X�7r{i��>��iޔA�$/�:�T6��&��K�O��C���]?��{F�HV/@�]��$� �k�BqW��̃���~E9,b#��woS*��R�ׂY��Тi����i3l��J��D�@�j��
׷�	愖*j������92(�Z
�E[@g����s���U�Q�R��u�1	�s�ᚮ�v�9��S{�!hZ�N��56��z[�E�Kj���%�\
Cۮ���������/�p����~�
��0�CU`��UaG~�;2M1�1�������9u�l��Sb�=�	����`sr�3E��Mk��Ɖ�q� w5;�8�4�hk����s7hJB���� 󐶷��LÐ�mQ^�x<���G\��ޞ�S�<?1���i��%�e
"mB��nC$r�F��F�%����ܙ��p�Q<���oy�{�h� J�l����W�@:�ifx�6�y��4$Q����U�eWRn��!�27Q��PD� O�e�  �Z//֋sn�y��tf���iiJ��Z���/r'�DM����(J6�oU��D0�h(���������蚓2-���+'�+Ҟ�'4�g)�X�F����k�4�S���u����m�BX(t;��.���N}B��느�G���B��Y.����}�|�����rfp�zʀ�hz�j}��,2s�o��F͈�ڇ��^�Fjs�U:2��BAs�u�˥��І#Ԕ&J�w�U��И��ݬ֫ZvpP%�V+�)a0(Y	��oJ�@�ٯ�g����o欟�3e�,���_�xϳ\c�������c�~�2��9�\@%�O��l>�/����U��0{1۝7�ppN�����w�Q�~�1�>�Zn�͖C�39�V�v������=���@t�m��
Ub��g��$�=�-�?�ȍV&��]�|D��	7 �"F����[��dw��C��WԹ�G����o~殌��~�v�T����P��}.���v��t4�^~�;� ��]\�jq���wa��U�|_��I�-:B =�k9y�,B�zYо1��;��6\�Yc�=��0`'�g�����R�k/�m���,o�`�Y;�ć�,<c��j�3�C�B�p�W2<����Gμ� X����aZ�+ς������[�im�DcS����i��UL�l~e1;��Aj$:��b5Blu��N}s�?���}�n�x��"m��C!�=��i�Zl���]�$�c�v��z+.E�I]��!$t�.t��5��B2�=��~^7_]k܍-ل.�_[�����{3��]�5��uL�"9Ȏ}27������&d�Z���,��0��/�ky<ǀ(?�A)��ٱ��-��^�V��~T�:��ԓ�>w,�7���o��6�u91T�Hֳ�F���?K��P�L����0����sP����Q�"�4��6�D���4N'.V�F$��L�N�x�@s�uP�̭0��fG˜�4��񋬐Y4ї,��7/B/��B�m��)h�'=;��5E����LU�t85PD�0��V���� ��'�߼t#�\^��lf��v���s�7,Q��wro������WO�*g?-������V����1�q��Ia��s��vm�ȉ8JN����~3��~� ��)~�L�TƵ{{��d޲�)o*e���:�'3��0���+gnq��p��?9��Gh>���a�2B;fx�%�p��m"vӜX�]i��
���T��W��@�O.�9o&+^�t#a����p�v(&ق��zq$q�¯���Z1���SN=ϼ�8ɩњ���E �邼|�1��@�S��i�����ga~7�����q_o�w!�\_�?t�� ��im38�������S�V`v��<,,�]f�'����pʕ�u�N59�.��N��G� 5��ψ̔�!%Z�B@�bhB�Sz�*��)�͸�~pr�.� 4�C��$�0)��4�����A���i��?Bh���a�!o���]�-�|��:x)�F��{w�O���y�j�ω��c�Aætc���XY>��bS�l�`�x�w�ȵ�}��%Z��������/�
ZE�	PM����an�p�g��cDM��Qy�Ė!��U�6u�m�RV^.��
O�g��H����D��s������.�t��O^�T�= �&RpZ
�1��#�B �����:���2˺(��v�8!jt��!���p�G�O���{�Ɉ�*�'A���#Pt�D��Բ���b�d�]Y �������1:�&,�i�����-^�Dǈ	���Ӱv`�Jz�;5,۩�
d7�_��J�}mw�@[��pɿ������h-4�Y��gl��;��S,aq'S#2��r�� ���l��!�+B��{��O��K��|��NKCK0�80> �E������f.��Ü̙	��4�ru#<m�y�\ĸi�˝#Zj��B]�q�e�I0Ů�O�e	)�QT�I� ��0�Mzt�+@V$Θ�`�"~ro�z6�x]G����&r$����k(�6V���u{�>�f&y+��p^c�e��B���XakDY�٣���2J�ۧ��O�ľ�s�֧������"7�>N%�p�%��-�>����r.{=3�F�x��T{�������8��i_w��.�N��e.�l��=U�!�0.x�}Gh�*��c�E�I��K�6��1��s��e�y[W_:ƀ~�3Y§a�:��t����fR�Q��wE�:��=���.E��I�'��'	F�y���c:�M�Xj�����c�3Á��g]n`��h�ٺ\��ig�R"���
�|���2-��4ln�;$SV�� ���
��Um����G��E�e{\����C�v��d;�/^�#��V�Gň�n��'�w����fg1�p�[��Mȿ�J�d���z)N��R����h�OU���k@h%��ƅ��.�.�oHpٷI���~�Z�eW�%�3��DԷ헉<��J�b�8�`!�_y|�����h��`����m��i����f�ݢ�t��=~�8�Kr��ր$��9���,3Q�`�V���mp4i{��|�騉�e�X���vL�>Tk�DcM�b)wh��G����]C]��w�N�u@��fv�*3-��}u�WNY3�ϤB�����ܝ�_b�#�'��@�/��,��1���J�{>��?5K��7{�P�Vhz<�<����1��f��|��<�:3��~_ٿN�Ź��')�> إ��A�`�Bm{(ƕ!��ܹ5q ��u�M�(�b��˝�#2��rz=�6���(Q�S^Qz���H�n�n'^s�͔���9���=��Iq:B/غ�I �!ǫ`,z���S�q�^���_�VOY�.0�>��7�%��di1�NC�J�M�B��!�ޜd܈�r���$�&֓�ƪ����2b������΢�R�ngn>7k3�, �&�䘽Ԑ�X���в�e����NY�v����K�]�9�G6�ͷ��j���}�b�`��f�r��Br��'(�T^��{u��[d��	
3�4�L:���H�:�Ͱ���W��_���"B+F�p�K��nA��I`Q�%g�[�x	�.ۼ� &]�;��*^X��1D��E$�|/\�s��[I��!�^Կ�0��b�'����h��Q�9�:�[ыGԃE�}�x@��U��9�1����<��l�*a�+K�Ҿb��aee�ˮ� W�~�B�	����Єo���^�'�'ou4k�t����kv34��w}�(���\+�c��9���nuFpa����}7v�`�J#W�e���Q�z�/;��v�]��'����yPn"�n�	W���������-K��~I
 �� 6/n��'��=��녩@ڇ|-�Z��(��
M�=��%���5),a��'�=���!�G�9�I�[+�)ᢌSWb��xp�^K����n��q�.���Og�[T>�m�,01B�j��Sv��� k�
��R�m����#SĀ0�eܑ�bc�ל���F@����|!��S$�5]:e�k����g6u@gZ�樉�֪�ĺ�]�kH���[O24û��M����P۞��N�1���C�,Ά���*�a���Qn�~�B�_��٣���0L}��;a���J��A��"VL,U:a(��=�{5y'��[cq�%��T�����$s)yl���Y�i�
�4�4V8=�A�O�Y�<]w�͎�%�\x�XK㱵N�T��F�:\5�J��7��|��d�Y�b�w��8e��h�,3I,���IXp�8Zh�X5܈��Ma��G{��^o&�M�W�vl��2�g��@�����N�hZz��<��i�#�$�'� ��<�?RH�1�4#���? ��F�(j�i���ZN���l�:#zFu�p���:����0z�%�E,�4����&�Lqp ��ܒ����)��YM1eW�<���S��G�g��[dS��@��}D�ϖ����0JnnOL������S(���fD�dbP���:�K5���:z�v��o���R���t3�6xxD�6X�� �� M�*|��t�+�x�S���o
���}j��:�<�Z�2��&��({��r�«��I��P�dj�".�U����T���(Lu#���BR��x�/��&)K݀D��}o��=�lժ�g���c��4��B{̍T>U���;S�7<lu����e`��*s��&�Q%P+��SK�6;s��}�RU$K�q�=����wO>"4��tB~pd�
�?2�%���Sד�/Ŭ�sY���j���=��d�Hf��Ψ<�K���h�f"�X]-��`��@����ؑ�����e�mE�Q�2.�-���v�Ɛ�'�q�~g�N"w�]�ܤz)8^�6ē�E�1���_��$ڭ���EG�̖�.#D�j�}� ����A·�(vh�+ӯWW@'��XH�U6-� �7��.eP�MQ[FV�H��f�-'�;�}�S/�*�ףg�ޯ�v��6��T�lu�KkW�n�	��'B��nf٦
f��%�hdZ����ɿ�(7�cWؐ� }7	��髃v�����[�T�}]��/ۣ�V8�V��0Ľ�,�T��.1�*Sg�V�YJ���X���k����ui\T�����t�$U3�A�V]j�fg�\uۄ�l��5L����6���%>�>���C�|���Pi�V^)����.��-�7�]�+������X܏"��rG ��Db˽FIX|�2������j�iݜa��Y�W�.(��Ԁ�-���ph�Pųh6�H\�15��Tx�L����5�����˳È4�����]���a��4f�;��[@���*sPH/��qo�`'rH���yf7�9�����y�>	 g�|*Ɨߦ����`?H8�?ىK�8g[��~zb�d��)�?^Ȭ���A�\lM��W`=o��pK�����W��m;�pX%�_����q�v�0ë����^&�gg��ʆ�*�Έ�0Z��i��1<KA�@r����)��At��gvg���Z�I�<��|a�2g`]��W����O��K�/�vn�B���Џ�2�,4��"?YMC>�lD�t�佺ຆ4"
zpv��ի���i�>���c���=��z��P�9h��(�8��OT9��riX^L34s�����đ�<y��B�a�9a�A�U��\��ő
���!�;rzkI<w��Axˠ_�G����ls�iH�pv����[�T�z_]zz(roKC���@o���;~jɷ
��p��]'�$׺-�N.s�8�3j�bz���B��e#���h�G��[�'�C�A ��NCz��X!��	���W�A���I�8O�˂�b�2UMB�������{��$ĩ�DV/��ɨ���'�X�[wJPd�[=sܧ[OD�]H�_^�}� �I�4g����]^Ί��δk�KyК���[��ĵ��߿���� RsŋH"
��'fƭW��B"��y�� �?����#W�~��c�]RAҕc�q���)LZY��P�p������	�ZQ|�=-#:O�V��is<��?!��#�ɈA�0���`U��gm��4����Z.4bf��Ț']��QA$A�s@1��ӭE^��A	"�i������A��Z+[�������f�F{W<�6��~��˕w�K�����8��ٿ�!�N�Wu�Z��y�u0��Y�l�����1���L��O�h*�nݥG[QNt,To�;��E_b�i �U��7��Fc\a$G�Po�P��:�4\r���h�̙grAX�=�5�N�z�n��P�,��{���w]Q��կO�pi���wz���.�e:�%m�'����R�Og�I-ّ�������q�f�lB�t�ˬ��!ךD?��!� ayy�կ;2�S��,�[޲'�EڇF`�?�w�I
����t�Ν�Eu���Q�(�S��p���N����P��R����(4i�B4?��K��<��� ��)�^�4 Z�b�E�����"r�"y#��{j����9�i�c�6���Bo7��J�^,"ݪe�}'_�[���Jk���d�Ӆ{�˳�O�#�>�p�M23�[Ai����cV5����v��:I�+3CD=�K�:,6��U�j���U�S�_�Ū��Ն�&=˰t��}t����A"�<VC�5J�n�:��f34�;9��T����E_������h�Q�Q��WԤ��) �t����+���Jk��uR��ǣ��Q4ܺ�s�dl�v�_��e�\P#!J�i7,Ӕ�-�@�4fw�B+υ��r������-|�Cd�}0.�l�9�����0�:{iC2�� :k1�<{��P�V�Է\ �/E��}oR�B������(X��b��f��������{7�昵�]�_��~��1+h���첇��������h��^�阶-�P1��Ъ��[	P���Vvx�4�����i-k�Vjh��`�YR���tB�]X�W9��'!]ßІ<'�2�oF�Ͱɤ��v����k��t�æ���JՅ��am��ܞ[��I	�0�v�]�C{�x\2��m�d�fK[�����ò؅��Oe����ɳ�jn�'p�6H��O�Ø~\��3K�uc�5�p����5Q��pY���r���;b�-19t�3����n)��fW�.��u��#�z�S���8ڡ�����2>6Y��U��./>DnH�x����obq@ZI��c��lH��\Jy�{5�|vq�P���LK�*}W*��DN�l�Z��3,��*��ص�/`�`>��K���a�G-y�������7�������I�u���) %�e���t쮚Duj��c_� >�mӑ)�1��Z�>z��,H�C^Dy5M�F���?0���h�)_��2a�:\_G�'�|2@t�`�~h���W��s�˞݇�����zc����	/�U�$��6R2���!�<"������]��e'm|��%G^���ZS����_�^�D���P�p��H��@1�ƿx�Eb���k�jqЇ�'���ʪ���^�ñ�mL����Y�g9�����9���z?x�����3X妅b]�/�v�v�҄�zߤ��@�P��B�_C_�}U�������2ϐ������l6����elX��6�+{mܮ�
p�����j�7���o�'��lb?��Z���ni��v|����{�}.,����) lR��-�ￚ��T43l��`�/�J���r�"�:q�S��E��9|�2A�u$�\��Z�������ScE�	�