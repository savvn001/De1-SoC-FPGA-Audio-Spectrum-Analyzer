-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
foaCLhn1ZfTIxp1ky7JtfHsoWixjIWNWjroayEoCoOn/HFqbF8nEN9ja7a93DNzdsGCIv/p9HuUj
OwXBjmE6AEFf5JMiF1sYev4a1R7fFTyXk4OYKPGsHdKF+iDhAa4s8mlvahtQ35dFZk2rdfeTo5uL
Pmz7eLn56akQBRGPAeN7dVuGhnHIjxZKGsSQ+davDjwErrxDVu+39YzSlwTgER3v8JcEk/9c9Cu4
2Y4WfO9+Re8U3Ad+Vh31Q2U19TA646AyJUmr07OW1Z5qLg7wSL5mxB5c6A/RY2TSE8EQlKa/a0Mt
mPr+EHNPciG7EIFnuQf3Z/D0JDF7k6dhxV3NRw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
Tck0YZyQgx3ZvmhO3TM3dhp/U0IoLJgnxbBvdyqPCRqZICE0SmGSe7LGb0aaVmC138bh/0nLalrx
oTEn/VSAs9sRdiwB0YIKGPEf7dSSC2I+9LQeOtAb8lEZvh6dh0bA8/t/48myY9cgh3iyG87ZQGvn
e5U+uvOsi4WJ94Qn1w4Ou1a2VdqsSzPBXbbZpAHYLftFVjunwI9ojG2qpeXSXOWgdLsy15LUdZu/
3OQDZR6YA3aXdpQqr/8xeETZMOGeOCSELfTykqxstzHZw7luW2hQx5dvOi/E9DqIhGT3gTksxcTm
RhgEM6SIeULfL/HGKHyV3hhrzuBoECa/a9dFn4tIYeX8dzCQAT88SEj/GwH3JfFquc2gy1+4O+FA
SEbSbS4EqtHp0kSg7Y1AXpiInI3LwAZJJNFEwjLgSJyuf4x2ZsPr5Evy9S6w0GF5Tyc6jg/xM+wl
gRRslWmtc6MB3CwE1XfhPqtQ5uVnbWgHAbSNrUmD7dv55Ew8/v6AlnFC+z7iaz4Lm13Hk1ucB+Cl
pxl/X4cdUHOVz2SuQs3g3Zkbg2zuYYElTdLvxpyDf0gXllJwXa7cF1TuCczA2WTKeGc1tDxOA+m6
e5whhpTfxFIUXHLxX21e1tTU06+nS0zQaekqs5+hmfdxUQMj3MghmrEWgsGrEZtNINl6S7WfRybz
eWQ4VojuWYQ8EjsP1wIt0Xya5JVh6oDGYxgcy/3bHpn/OgRAIj6CaNF3JTXgjUGLa4RQmtYytCWn
ydjHi8UvTGvABQsbYv/bf2EVx+dmp+DQDNnZ9ptrKfBFfOLcUWQQehw2uMD5lgufz6mzk2cvtZTR
FDuIbC1OddZ+Wi7xYxGPI5/CPtlwp8JtqtEgDEo48Mg2Ne6t56ZhsqosLMVU2dGQnYBRj1aSg+e1
v6HJJxJ252cujC09qUbw+pFOuapLpf/LAXbGMq5MPOGkFxmm/k68Zq8oANrmfO9RtZCDlbhY4PTI
KfCTKFlkUwEYZAHMTNWkaeGh0a3K9JSWiFgAg22226YmZH7eWNINk6YBPppEBGlgv4hxoiYUQE8N
XHwy7LPj2EchtrVELt6jYWuYPuSYpYlIYVHNVZBacu8RwU4rTw/Ovyn2xOIMaqq6F4+GhG9WyOKk
6+f0KQ54XxvI27Asbr0e/l/KdJ6Q7P3b02+ekCizg4RaT1M5GP/I4MWk4JJoCvJDweQpIqeFy16w
UZOKF0NqMD0eHwsGBMAA+fwLO0rzyXZa+EMwzbPRKJHXVB1g8PTzUAU4pd3EyyelArZnIoCCns0A
eTPZmFCYwy4FwmLmXCGZEChQ91i1f5/kpUqVgFbYCyoCZe1/TETixjSfgFLs0g2KoINlILZX2AJG
h2yabh7FeRpilYtJ2W/2TNOF/0YYq9yQR9d0YhAlReFzQQuo45/JejBZuiI1exVNDTymE6U7wbrr
4YyOB48aK3W6038yhQjG32f4cidxQsE33sW5eb3hsh/VdYNcNm+Z8H97aF+YmVhwfwJxShy9F5xq
sBNH6ns+IjyVad+N/ojy597AFwqIymfXNQQCgzrfutkBzcVeSnonJRtlQqM0VICgq/hoOD+cuQBY
7HaIoA2BXgp4MfcAeqTvBSxNDTxeQhUj7VPsgkkS5gdiq2QnZ7aUtmIBCk4CppO4c3JI/cGCl2sh
kWrJWBGhBOH1PB2qsOo9amuo+TNmwq7quJIG7lggMdiI1Y2Gf+Ml+Ro5Rpxzu/CjCAOAgK4vMzWw
dwBZgJe9ufJo7TSWeEgZKZA1l+9etPk1cxhNIYChCazRWOlH9oyBpQsPEkS+1cYGuwEf9jZoxc4p
7YFMd6fL/KV2idEt0JR3vKW7Z9TGmZo86Nz+2OFOVUXZ8OJpjDBzwztPlIKx0A460SI0B/hl3bAR
WB/5kWhkoIvY5UuISGgTbGgUuBO3nQmULw5Z4PP+JC55BBiBWBtWhJlevvTkHK86mt7H5o4LSgBP
6PaHofFz9XnLWoFOXiGtSTePxD84pYZSSJKNiNLHMIEBaOUK97E1cjJWc1f3AJxvEAhBDKjETdCO
YR3q0pDWvf3fS6ocbc3PrufWKO+LLFwaMtTRMzw/NWUEqnwKxEzIj+R5TRPmQ8D0YnB/26XE1OUZ
nawcLZuD2dRHPreTMGA4fkOWHGabIRX8bpOjB/wMNnxKl6bf9rzYE628pU0EgrnDRzYnShoIRhFs
4d+2EU9PDimmdxkkdaRwp0iu1R3nFGsC4w5m4AWW+HtF86g6GilcYQMjCE6Fz8aMOmIrPYRfxfY3
5aOD7gT4oxSZGPAo/SPRiH7SuEj6xPPRnpbGXbnE768ISzt1lDtuvv+6JE/ImpkQdTXHkbSQ3apO
Do7r3es2F6eUc78Zb6/B7N37YXUupoGs6kJs8aolz9H+dycntwA7v8PvuaG523lQOLg0HoUW5moK
d4OD3nOkW5FBk+LyA+zdbIAV6dixvyvfYB4N6CfQlZ6OnG8pvy4E9XSjXuXDRUb0L6bVRem1x6ny
Zp188pWQ2JJuE4darITPVfk6QuLXCww9rbGrYPVe9pfjCDyPhmVBPBDhq04npqeLVtb/gVPNq4pG
NEeQVvbm6FTDhpd6j+47k6fJ36eJEvWkzSluyRLbwVTGC9US97ABOYqbiuCF5MyUpxwlV08aYmDw
HAC9vH8qHUmXRzU5DZt8GVj/Ui0GjCTZYfPMuVnF4BORi3wF91FDzmDcoZl3s0xcyXEaVudkQ1Mi
KPv7CM2dbb4LriUElyfLXXEe1iAu9UnbMYmNfgtwxHnqKl4rdaGAlHwZzCxrnIdHlsj0Hc5474c3
XfbJO206Zyw/35RGs3Saq3pB3m7eujxFoPIrguCYanUMiOckO7uk3ZpAg82k6rucTScmYnEehZNw
T+ZmwHIY7PKULYfTuUYaSG4QKhu2u2cUFA+vVsQYUPvWwZ24amC+BmY42JJzBxvrLcYgUNBr7F/N
wXddLDcvSIqOqo/JBUy+BBko8QOKm0QoZqi4qq6//nX+0jKuQcYtOkfNTkef3gKwfJxU6Jz5PpWM
WOt87VcuuSHoiTGuGoRUO6KYkpE2Gotl7aTCK6D3bsb+NPglvrySsdBVJZadYGgYq0uks+OcYN4R
AAGZGA4l/JM2IYErNoGXaCqNqzeJE0pmig0hnJccgGGaoT4HbMjIwm3r3oxz2YYV3WImNy0lmuk7
jq+xRu/Cn7T4RMqPox5v6HCNjFX7L544NYWqenfiYYX0o1UWLskrvt9RArmZ9/II63eG48Lb48rW
FbldO/R/cxOBt7xh3gqb9hXM7LV7hoGIsd97SFY570EJaTzGKRr1foQaRqfKVNBazouiKyOJqZ1v
MmPSjvVu3bb9hP2j5Z0af4MJU1NiBbJp6zlvAH01GTTMXixTILKbdVFnd64WqaGXQh7osKPIyKYW
x/J57Sf/T1Yff3LoJVbE7o1vuk5Uv7+ZwBR9mOlHo6HgaAEABowFg6+DwpheMbaW1qxSQKw2FPCO
vnYuTdz4LiCYPBEWWI840Au2I7i+g0hbMJWyNRWxUzHZLLAw7UGYOuwdoHXvraK5ecBOkV1yxn+M
s4Ap7OEN4C6/NI5j/pGiYjR+Pag9t18VqKHm34GlRgdwFjQv2W7nWn6Vc2zmo15/tu3FUzfXSRvf
ucJkGp1BbUTA4g0cS/onCl/QHOKy+18ZGQo3PMphxQS2/Sv4HwuP9sKH1yEPHy9cTygb8H1WU+Ry
ch9ol71q8z/uDSxBcKTkyOb2N6yYwIEoGYZZaBT2hkSKfbuXIjKNjLE0aZHWORWfD0VP/b39MIWq
vGnv2f581KbvCvI+y6OyaFxfA0F/1nlDsYOHb+5mfMAjYp+pEUWbdkGjkgNHYiESHfUFSdLBHXKZ
osSWs/ocMJRlRAmhG/rkKIpHsQy/igeALjtCnO6Gt7k4ELTfIT9NVOwzqGW9AKHp0RdjI1jQ41Jy
omeoiO2YjiWioRGGdv2Gmrr4KrIfbRd95i40dBaXzFNo4CF1DtCwyRcH1tazT9hE6HKf7vuD6fXj
UX8mW6ff/8Q2OFlJDyyx1n77jBh8r5XSGNLamNwuP/DVzUdHROFzs7sWnvWYkdlQV8fhMafmIf4P
xADSl09eKfMAlirDu6whU5ZHiUxKWwQCZrN4CguCrQoaM0KLW2BVs8NsxwNL2b4xOqbt2R6STjmy
uqffpEsM3eCrpsj7k0+KxxPlOGLApMcbqGnJxjGjINyhVJqtWQmkmpeXTyXOzinudguX8RslJysf
ho0Bhcf3dLG/QRaT1qFZTeNou789wFvze9vG/ZfJHtm9beZYR+HR2VSXX39zQZrFaZ3XkWIz66wF
YGmV66Gbg4XEAxwNUp9WOisfcg/5js3W0sSYd3VMPtIMtjZbH4vkPltk+5DdKVSrbFSpVmrKcF/C
fy7fc9KV8sBlN5P1MCA0RHye99Zervma544t1PHXncGWq8+lamX6g8GrJHi38YLoUMiU0+ivEbOw
CfE1nbDdG6NHh6U/JoITDaLPZy8XXQcKMwUMa06FUxXXojNxKWwHtlK68l+UjAlkLGopvBQw8+Dj
XVSnFrU4nR5F5FY4MkQfzOkD/HeC1fMWBHouHn/kmKCgdbMYZ9nnp/BjNtegs0IJoS80hdZSKby8
FQkGWSFcPimMuelSFCNuoKunYNjJbCVrasYMoCI4V2S6IYAg6fonCoZWp9Xy02h8Qy/8GZaQIhdk
WLnOfbjREX5QeyKcVKo24L7vPRoypGtS3G85YCipxXn07EBRFUrS8EB0NLxeuoFSxatWViU+47MN
IlzTEWJizkbNNikfaSFwZ+gQyrYQs+lAr7TrB9X1e/kKotqpBz0f6Lu8+3Y1OrhXPhBQcZlfjP6Z
dIDBMt7rMg1JtarSSBrHjpbZPrGbE8dhIMCxu0fof1QaOIARcP8URPwOldWm5rzbT57GcERL6A/3
J/ZwRCyjcYGo3sBm47+xAaZKMOOdkb5wKLJKc6mR/PFvJUCkpBul4iIq7fqbgBlrzATx0fIfzfjX
pj5qhXxpl71jBEVead92Kb3xasSJf0PpOWUS4pk2SqAmPfal9PWKeXHkofTDc5MdtQEDU7CRvIAu
yvBPhlGgNU1w5PlPxd8wUWHUzjhZvPwRSX8vEihW3chfX8WPx74gXoK8P53ocAO9wpV/4LneBXjS
8ytkvu923ZYXU+8StXZgENxmpQhRbRteURFFbE5GGA/pxWADOTU5dwn854/deoRrU8pUdmxKRpM2
0XAvWGenrV2TU6vmH0yqHRnylRlVMP75qsnZ4Jh2cfNZD+NcOkhV2Z49eCmU5iS6M9nf+nNQlA/L
Axrg/SymYzWBVWoh7oQTqJT0ywkbogvI7kUqQLU373scr7Y+k7gE9CSis3tCJvgvceDXz5kHOv9T
Dq18HsOEBQSKWF+GK3MCyzM86kDTgZfCIxD3JqZQ0zV/+bmehrIdXlLbLtgychWzQ3zI1qdSjWKg
jeRCtPXQblLDv6E3XrKsZWqQ/Qo/wjQ03fDQ9f570qcCQm+erp8g4uCeT9K0uPdKo4cyIY+MygAp
G33ih3BWbiaP2QpB+mozajfPpsu+khB+V+2V5JCBWvFSWoc5SLI5OmRXbb/EHHsDdIn6Qlcb0lFZ
XAesIm/j6IleAAj9jGDEdD3TLJblWK8w1WvGKxXyPUnZCgDfnmQ4aaT0sFe7iivfGLyI9AoNphS9
geH2/RkmTr2sibvTc9niY1qPtbQd4Ddra/TtC/jytu05PhBA684WzJ/6SXNdEjwpcfcFkEDhSBFC
OMFEp+Ak2/iAKBWujDtUOsLcLsk9bpYRQNjNTpIAR5nWpJGEGzNYxHyETCWInsqmnI/HirvNNjMS
Hu2k/377D8ZkcF9eF4j6czoBObRz621I4JpacR9iO0PT2KFxmcNhcngIgrI3/mrc77VzF1u8ep7E
NEaLIqnLFzJRq1WUBljTDrXK3i1mcZK8YL+zehYD/A8t2TTwRnQ1APZjt3YPsc0EUM7ViyVsHyUP
3hqg4ujOyvHOU3xNXJ/9VeRIukWY3kf6PnuybjXhtfmY9m4RpCNZAw9sttuv4Yy6aT4JNXP3OKvZ
85HIANFRj1YhKiUMURsixAivMw/cmVvrIMaTvYl6QNhWmDV4ZEW1+RxkdxmDcgCAx1bMuYFoX5aR
WrzBIvz4sFE+vDQqEAj2f79zeSN6Ov857R0J5HhjG838f9iDaz8efkHDvE0qTriKh0vioyjU+6+1
+0bhtE8t6vE8T551jv+bWcqok2joyCwmowhUVy3kr+VZpc6o/CJnrV/JE++zhlto8J0gWSDGv6MK
XgP39n/9ch+W/W46FExgkEf7a7yhv5OeYPaL9/EDhW7W7g1ZkybgKC0RocxoiI15mbPYiHgVaBBL
xe5rh1JuM6OBHt48C0FhQ92IeYhuXQbiA5zHF5s3vMpBpm6MU5+T7vH2FW70W/NcbOPc5ucan7YE
V6alY5Ho2crBvRaHfCAyL9rBJifmlmOP4pTa/THpo1oGs/pUU4MHfXel1gKusMsNAkFFXJDbzj4y
QfAOZm3Rj0BUQw5aNGNhm41F/0qSJyj7XFVm7KHf0hQAYXMowBI5NCC/C5bHzZYJmY9Zr0qWKggb
lhVTrHKsh93YrjQzxCLda1TokIpGuls52u+bEuv7OGbCt4LFS9YC/snl0knWOdiI/8Mo1ZHqlAxh
yCQeKgoYDiE4Rso/Zfe889eQNntoydBxCHTZyvj7K27vSZIktfVCoDIZfBwfJgMhvRMjdof3E2HS
23cbqvp6qJ0nUZPkz6UE1lixxFPBB+A+Tzp1lUWf6UW+8UgAt9huVJFWxIoHCcy0UG5Xo5tlEES6
1zKyMlVqLk34Bc54hcbL+sLEduDhZMNa9CIbUC5ZTIhEq8UoLtoAax+ZlzpVRydGzjXghAObjYVG
mw8RwCKddjw8/qja/PMX+yJ+pA9fAgqSbieYd3JWy+GrZ5ro99+AEzoV/IjAAS5IjZVDvMl5MHlx
6dbE30h7PAhKp5rM1uHxRroFaUP+ThTN3hbY59txrgj2+lTNCqVM5oQcpxxaCQovFG/HEI0sxoQF
Nvot13ryMFOLnwgeVwMBdJI1h39nfI3dMt3E5YGdSM2OkIcfa5AEljhHre9ViZTE+Yp6ijE6uElT
wPfwOwdAZiW7sNS2KaegMaNhfhrqxTqa+knWCpmuIa90T6MwNXgRqlWywvm3Ss5PxmgFEpBkDmOz
AptHqghX8oIMvADlz0C5DyatzKMhPaz1n3Z51zpD0uYRz9jtTFav1I9c1W+s1unVN+Uiuh3aMb00
IswmOcROkLr8Y43sBbTnfgAQUj72uAH19huDApnkKhBpHyg0UUqIN9et05+ZwR0xZLYrYzcwEJ2i
gp8/qkuJyunoI5UTqCXno3Q/ejoJcUfaaAbUtfvPn1tZr3ebkVxu9A6b+cDdJEPSr7BygDrsQ8nH
E1e9HIcjniwJVSBMxfEK8STq2V1/GmnUfMbu4LKf9yZ8P7y5gE3Pdnxc59cY8hhbdjFdSlZbw74R
/pxoL0DiH8oxHzCguHzCnPhn4iAFlWrHhyYXNRolXzDxyVD496l1OZ3rhUvXnYhY7l3tzT+fNpEU
ftYuoGfrmnJdm1P6ZrIF9MNgxWDT2MGRsAji5WuUUNl4jUS9AEKDwpZoN00Kr+8kuxp2f8QEvQRj
KsCn3Hh3GRxYv2hryH6vhLBaQKE8oabYZDax5PsK9oWaH4yTNyZxgrCE6M38xNJ7cL6MilZAPeLC
O0kdFTSbME7pijJacKQHBiZpk7N+hoZw045m1lNgZhF45+9iv7tOAgLfcdlmXZG7jGtcmd0amNbb
9nUaa0U/r6XnGakvOBHHo24lQCv88g7ioB9iZXxDrLSLP5UjdEPmJdV4h6ckQKrj5++s4XxpT6ut
nE4ZRUvYBsU9ALg3yh7LcCSKOc+7m3YndDMnYNUKw2J0YFeHTmE9lNQj9a/HVc2tKW7c0D37n6Ri
HjrKKMtWW6f1E0L1lSYgeAhprKWcQ39+qA59xqba3vuNTSpZKPKkQTcLijV+kJIay06DoYkZTfeZ
cZJmS/A21UbzxJfOWQ9cdxR0/SGG9pgxPlWdNjNN7ZYp74NHqAaKY8lFriD8PrjhenhdwkxhjaJz
cOI7ggnzKEELYNWhjiLXFTlEvc5YOXyRitno72ZKiWvhtzE1fdB9KbIDzw1FVm5yil3ke/NAnrbA
YQ6MUETgfPbe6D2IKy3ZU90Q2oFOlbiUzN7P77oL/64Wa2Qf7B/ZO8yWSmLYAqE55i5edtEBIwlG
U1yiYfnbaSS9JKVvdAVIq0c8O4v7NgVPrIoUiXYxQjSh3vftAICXymA4F3jFQmRJ1JfPH7x613Ox
bQunWyZqo2OYkbdBm4AOyHnqutXGxtIqFkENxXv5s5KvOPJC0v4M6nk0Rbg59xC8bh6M6URsB53R
Ht+2G+sOKEv2GaDzjfJGNhOKMyjTuiSPKvui+fD97xLVwR3WRJCVF//F6XSNgmgyssNDANDo5RUf
17C9PPSdh5lUJ+32DBx2TbO/0oQq6lajie0gXzCP4MX5a+CW6uDCWkqKwWo5TNSMMV6yb4MPoQpR
llBeaDI5+xU8sNiAJv6jt0KlFAHf1mR39juWJ7Ejm5l2Yg9sp+uwrO2wq2nbWxWv8J9fQaGq2wer
iSDuXcYQUKyr9VNPfNQKMfU1r1qA4g0f5+zON/bj2kN86Hae4KZYxer1sXURLZNWO0SWLCLdQK4m
/AZO07EGDJbvA84eoDW+U5gH62jcvuzF66IJw3HVDs27SwRIA+xXHmDLKsTSRRJCJN6pcIk0Yy0j
L0eIymKGH+iu1YzFHQbkxiXIoOao082ihSTSA63x0Anu5xS5jRFjYTZKjLB8KbAqwNJvujn0HDjs
t5xWM+0EvE5X7gfpIQZ72tVLh/7EaBGcU0kSI83tHMnqz/otf1bhvPwTF67Ro3nrxcMrWySTrrpi
twREqRoZdpuzU1O8Lf0aCjAGFhSohHucgs+1xnkUC5AmxNm2AE8XBsA1VcL4tz1UbtVOHpUVkvWe
lAQbJ7jUv3JSMlTglkuFlHv31EAf1uZRNzdb6vCPF5xhF6tbkVUQQsBWuRXA3syoEWODanmvz6Ex
kZrnYjko53we4Hlx6ROOPlkVDljvhk6KdUBiFTC8xkimGq10exyYslJya7M1icQT3FJNFMPZ+4Np
hw28RlKVl0i9iJrVn+OVi+jYxJ2qBN3Ty9bTBedXyViG5cqtzD1xwIt48oro/vyey/nks+caMeSY
jgeFaX6MR/whgEl7ZnePjjAtQwiCU7qEsrWd4YMovj0vODBr9x1XlVevN89eqLiAPDtA7+eJcUlY
D4JiTZnBLLKDYcepL3Mc8I7Da7qslKiksgsz4PWa+Dq30CfqunKd26wWv7PSa495wIdsKrUaFQ2W
TyGWlcbgObtY7Y1GisF1kfcUTQruhjeAJiNwVQPxCeIPtxl21AXgBvFOohsMVEOh2tBmlvk5ezV8
kB+nPp0ipxOJOL6Hj/lTQywqJyM9DyUiZDkVwJZ8ypDJgM1Zmy3oive/xq5jKITUjpWASCDQAqD5
UPVwiw7kLkvt9I3Zxxxa9LxAcb/RLqiITRwrE7KIM0jf6Q5pgCJtpbnkj3GSDzPethoPR/A1zfjR
7hgdOqiMB4jIraI+0hZ8Kzig0NDx/i8/23DocvOBcnDSHKPeCrp6BUqHsm/FTblQR+nYjlbPDewU
hxOjoyklMtv/+oe63kvCW6O8rkFuV2mpgwXTXIdQiWg9ifR9WjvtbWuDEnQ7FpOCcQlkMlB3hXHc
4f3HArm6WECHcn5wjxzM3R+pckGkAWDhHD7cPu134mea9QCOd9I1hcZ+jnoE5MI0EMbAXBrOxu/3
ThY2zKxqfnapVBTS9zFMOmGPUWmpnyX6cepQ93pvbv4xmcm6wgZyF7EYMbEWCgReTqRDxI8CDwG5
41//5xTQg91MkiVVehuPyZcjoGO8Jcd0XEShiH/+F+gdRZITCoUulZ+GJBuwpyR0jQylY/sHFXj4
ZD/gE8ZnNgbNnliDdllD8mZzDtoGTqRzOuKyUvYSNTAb5xDWC+bb3aGB1cMb7hXGk7vaSkDGklcN
QI9vjHOZtbDczjE22FyH0cqcwmC9Zuq9jPq2pVZxeXjJT99R4n31rzFtsyV3RGTRs/aoHfYHCkZj
aIdwOzvoMY1kabLZ1Q4BpXHY7JrpoxNWzjBh54IiolQAdQWKTQQgcJO63O7Jhht56gPZ/qkbBu+P
9F92+tUvY8ybNQdaZgbxf8EKxqMKWXWOsAaMAg1cXFhQvXzyCa1fA5nqK94dHcc5k9uyDRz5/9MB
owb/dbvnITZMc/KZaOHOsa0FgpyFaKdYl5njNR7mdJ2LcyMvf3XxFt8kc/UMRfA3TAcAmBQnIJfQ
zE9qpCKasSe/zd520iEQ7wgUI554hWAEq4ugZL60RW71WeQBBL6bHjMp04OHjlf9SQumNZsjylG7
MEFJhPCmsfWXATbsvbc52VagZnDeJonXZtm5cAT3AxmDrIrn/LwJY635+ozfRLFxb0klZ3EqWrrG
6ca7DVJngD/18TjxicOQrZ4QvL/cVJx9r6wUsMX3RqMAEPe/bmJbT6ubJwgznh8QFRQLer6xaavq
NJ3gtPQNAzuUVuvwv/L5U45rcShM0Qp7nkLJ1fCu/HMdbhcQl0jTCIkqSggW0pa4wQgPq/s4Gxpe
wQ6LIbWsWmrxKD1RHXWy243lSbNbYvhPtWTiMbi5hfyfzz/zfn8YU4jXcooZEQR0ObA/KnNGPHYm
2TTWd90+NW6lXEUVHgfQrQvPPK7Ot5scw6Cfy/cpM3pHrOT4xxxcahuz5Fw4rG6I6CxBJifcMNYc
7+WSHEKYNcpMlX6rsBVMpeflghw8dDjHn9ZHbL2g4u5NDlRlNg+Aom/rCHp46XfOs5tv7O4D9o+e
5TA+CKQJhu0aaUy+hAOEv1YuCsbxkq47VlAjFTjAAmWEBfuL3bf9R4RNwiFfu9zxoJn3mj5TT3ok
a7K/AXH6+qpX8SyWLWsHv+MovI8EqSyKpe1TPw03L4H0LIH+v1h5a15S+YwoGAX6OoBG3jNMjDqv
bzSsY2f9xUGDUaxUQupxWFFvp9Z1b9uo+oJUKxIOj5d6PAJa2KbwUei9TDHnv6TRv/NDz+Oq1fHl
llDABxyN6n9PLAX0kWG4LT5Qpt/E6h8vBm+BY8loWbUUGzEVqDNupygIJY2XD0F6Ql9pGtuQzimO
tPQqsA2cR/lgyhe7BQuhAPDgSdSNKKIqiuZk4QLhCWspEU0EQjYF7zWzIOggI6aqBsgrhPdKn/HW
ire9+E8P0H2iE57ggwXbL87OzAeyFH+i1rIpP12v6Iiyu6fQ91UCRBy7jbN3eYKcDFTvEWbuaEwz
Ea+smVVi9EBqhcHg74bApUZbSXc7gZioU0P3DyUh2+3It9IuYm/dck5lIPot1BgxvlmnHkQpREen
bFmWDL5iZB7l2fdFoCbxMGL0EAhOmsk6mBX473qz6RqWXAY8G/CXo3om/hiZPD6zlzvQ8meYi04l
xHRxsXnyb43yKu6Wr9s5thIeUZfHcq0JYuo3+W0slEQlI+blAhgZAc9Wm8NjJzX+V8bLgt9j2PX2
h8X0a0Qw2SuogwQxel6SRfvTfc6OsHF5FuZ9koFKLu7CAcEUdcluRX1633BqP25mlfvA/NpiZyZg
tGB8A0pGtuQeTqiyd+53M+I7cPLLRBVHkGhgPJZ8vlUyoBFp5SyBCdKdHoCEnziPPP5wmmNs2coT
wqQMP/gdl+w+O56btom20aB8+RbysCZjbZvZDZ1xm8FyhK4KD1rbkRDQntfhN34CRwnLlNz37CN+
OodmmGsvlt1Cp4FTFdchi6g5UVTsbszYGuO2SkGERlIbnsKuLHwILG9e4xSvJBRF9ngkOEYHG7Yu
DsGxSU/NNACTEUBQQJ7jK82xodUHRhYzsYn6/1KQIK7e1p0WINzGQf0/HU5qee3VUMaqS2UBzmMB
YWhJfbbMdDn7wvYs1MZHE2SmKOECkVlZ817+z0A6wtzvr82S3XhL/BGgC4UosQ/iyZN5DRAN5L5u
oiQEnJIPWiqBaPlWEdyOfPUcq2iH6M7buI3wPl3yeFDTpomms164gSAovZfSuJ4KmIxPOzxTXIEJ
pf9a+bdoWFcXoBU4kaRxs4FHDBbrudaVrvIgVpWmcF179z4GrKxveuuqtHTuUmS4zIy2bDD/By8w
KPvNXFGFSfZWaZQGJb8T5HoQxNL4Mr7SVVoRJ/1sbgDX5kkZpOiNQF69UR6s8DG3wG5JY0m8sE/x
d2ES52ZFOI56TKHKAZA/4LfXo0Ktj+GM40oAY1b9M8DNCGChkirXZ9wbrmZ+9pXNU5kP6MGVvUqX
sfzPrZKRdMTiW1a1SLOivTqskoQjrI1u2hQ1BAs/jQWeAFMl2bKfEjV+gr/G36QOwe/GyY4wctoE
chel10ikYNAM1Au1I3gEbV0BraJ8f4S6N8cw7gY6vXwCu6d3LKflbjTPypNaTX91pOY0ZovIFGbV
msOa1mUkYCv6yCxBUcI1A04iE+zGWJ/Rr+pFDTQnSQQOcgbZr3Annh+/hj1KjBvlPtd7gK00ZJGi
wRbAUyxNCSE8d13+2Ttxbn4SjIw8NOx+F1KN5WqB0tr4htqawgEZmWIBip+VEkr22v59qCt99K0u
QUKG9g0zQE7e2TowIXhOWDGddH6Y/aFnUmKNDBz22jkw6sVs+iUYgNds2ZEvmKIBpXw8d8fql2eJ
cXcLuUS/cuzSN1BEh2f68fFZ0vaBG5f5PZsh9zcDC6awAHRHsZ9jWCNhF28D0zUA8MTzV/i5kfjg
DLQtufGyl53aUmUsxsn0dmdJQ0bEywMnvZB1hXONn4NuOPXpEEYcU1uD1nrJQhBz3gFIL1Ie/DfL
Jz4VNNsJXAyMs1y1JtRdq/NC5o5a+YuxDbOISpchG/rDuWhgQV2ktk4XC9AX1NVCKY6riD5yr9+h
MuAq67uGimQXXI2+lUPS96Cztc2mgXN07TAuU0dKqC8OlR3VOD/JrnDXVlHgLlZ/8ORSmrkNQ6SG
JKBHKh62ka6q87K2kxvssMW0oF36nZmNfVyCako0pIXQNo7Z+ou/gS65fayhzQooCUbptn8Flhd2
PVS0JjwSjhMiNw7yO2CEKI8MrXi/tAZTKDCk1FWkiAay75Z2WxbZPIrKz3SCgEClF6fQjO6Y87YK
1m5LGwZTHNYRsNQ441UWaFsPGQ6ibA4jPsDsqZJTHDYPwMXVQ+rFXeaL2sD9vl8jOPuwVvFl9v6Q
BCVLA+wQaZDpZBK/RuEQGQtyOSmt+yL4n0aGHWb8wpr07td9dTAnbq40+owx0uvDFRWSwzCWsArs
tbu4ugUBL3lsMiyV3rWLXUkWbGYxo5MfGTRH96ULTuVTU8LBsEtrUTcKJxHmgyKwgOO5DKSxRzEo
WSBcc4pCuoj/fy2E4b6ca8siLzJMTfv/bLg405P0nmHrDyf7R5Vx/tw79eHfZvM2KeNGmI/Dm+0W
wgxoQsTIzGDMEM7ra9TrhjTaBrLaauZhOa1SmfvRQl3PC0ELJGCwRNoTin/ii39KwauRCaY6ERhX
XEFneb98QxZWu7KaaTFdGv8Z8o55dfIIjn1GTOuFjmrycsvfTGsbtMXkSl4MtKRJzF97Zemf0+EH
Bf3G/Q4+2wkjhiL0oA9YZJi0K6o0AahkIGdWcgzeRf004gbkrhu94rk4wOe69m3yVYcL+WzHfAa9
yqtAWaaSXZ247YMRFXmD7XO6IC5y7sVY9fN/1hNJRvnpLk6TCulSYg1N9r48ni06Pom+2bCFqMnn
NaJYeRJZaK/dqAFeCp/x2almG5OBaDizWcquSiao4001Jg/ZGh01l36Oj+B1SUFo1pibK2yUE7oY
u2zFBdWUGR2/8AZYXlKT7N3QRFNmGxMClTR6I/Lf5negKHPDnCssRtujLLLskuCsimsnQKb5GfIo
maP3Ei4tVjgWjtYwl6Y8wZtAzd63e+Z7Ipfxi1K8T1Q5t9QtWgHGNFVW4gapZ9GNwrv9AgLbOVib
nacaoza4CxFwYrZrtXO2VJUnUIJOCZzCU+C7NJc6uIXlpQq5fYK9sSI+1NJstrvJODd/wpZJ5ou0
ujAtnyON
`protect end_protected
