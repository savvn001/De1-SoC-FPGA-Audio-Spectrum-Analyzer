��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	6���C��8_�xc% ۢs(�B��m%����)����5Ý��{��W����qU�s5{�R�@��l���w:�B�%k/��Na��FҋQ^'�&m�;�S�s�fx��س�Ȏ����?A�XBn�uj���KBδ�W��q^\Xܥ񰝽��;i�k�N�@�Dd�L�ɢT�m.���4��W�X��;�Z['�d(�ů��5�25�j!�71g�S�r��$/vD�T��Q�n�Nx-�����u�ɊA�0 p�(5�`k�?	sU8՗F5.�>4Q���Ť�HX�0h��C�;c�
�ʷ��q3���@�h�f�"�]�0o,��x޲���%>G��f��M
�q����G;�͐�KA���q�g�p��F�MkG)�3(}�Cz�9ZE�	BRcY��+����Q�E�����<��j��$��O����t9�1�,�ǏދR'm������$EK�!�<F^/��P��-9k<�&z��ʆ�j�0��0e��3�Lc�e��@#|ϖ3�n�Kr�yޔB5�v�a�ٲ��m�8#v���ە�'|��Zxa*z-�#�`9��F��aح�i�׭ ��2�Hf���^��b/��K�/�������^�)c_劖F�W�-�g�.�ӆ�%�+���P7_+�x@�W�H��\�f:�# ;l�1����^�B��g­R�ݜ�{�ٸ�<1��>Ek�"�\3��uw�o�LU�Fs�hN
��qB��\<6+Qe9���N��QVu�x�������z�|���4�IM��������p�������!d���~�����._�V�&��vm����X�������Yo�*P�����6�U����_k�Wp+�O�hl�R�#��֖��
i����g�2F:+e_Xg������U�[e=��G�+���P��t����@�$��S:�(�l8B�����ʣ��[lS^qLho�]��?&.�Ќe� �����#6}Ԋu����P�|�	� k[_n_�#"��E��殻�A�6T�]�lkw&�f�%�\`B3�1�rM+����3WW�e�����1{�<�
�,��^���\�Nt+uD�iK����9~8-����v���[��E�Wh��Ұo�4���s'�〻�6A.M�5kn��%H`7�!���v	�ʍ��i����03���h���q�#zxq��nX����Q��P|�ѳ��"3��,��}��(�x2�'a�Ի;�a��n0����H@�\�jd�<v���"��zAm�o��d�h�YLG��N���x���0�|+;H�4خX: ��o����:�Q�%`RyR\Jh��P���F�8%E��wS��z�1�q�ˀ��٬�G�ZO�2��a6=yߪ����V�:��IIh��Mj�!��co~D� ��Baz/��8���
[Q�;a4Gp�bZ���+!1�.��N����|���&��.��dN ^8k%��r:�P��F��a���}n[uxj�@f8%@���`4��&��u�����>�^�8���E]!�xOx那i��O���}^�I~�<�Z%�ӕ�D�t��%�8뤈Cg��eb�\�s��t��V(nc�8[e�vvg8�T!��+�� �>%��	�z����oE���$�\�i:^��|*���<��p6������%���Ak⏭d�	ş���rB%a>��o%��A��7�z�u�?Y#�q:�e�}s?6<M<Xv�#�Le�l1�GM��B����Ʝ����C-�ֶ7m?�I��=ۡ��0���8�-��H���_�s����/�@`a�0�r\����_�۴!��/���֜��e�"�_,�$A����K|t8,z�X��
��	�%��*�XC��TU�2�E?�ß�g,������-3 ?!��z�[��ʼ�E�8�"x,�4/��\����-W�|��{����_�4o�_��5��u�XXPQ�'��:�[���۹����<qJl-�%tЭ�����U���.�-Z���W�ޏ��*Nr�N8#�֬���
��M�����k�]�u��\3��W~||sS�PѳC��ӭ�z��'��Y*'3�mJY&l����DI/�)�8nf���k��d��&B�:ы��\e$��稸�#�{n~NP�8�͚D�eA�����`��(���0� �sQ��s��+�W�q�ʵ��'��qe8��?�iը�
����I�gK0����e_�o.�C�!�EBc��Ch��I���U;I�j����Ѣ:��Ѣޤ��3���07��2E�z-���(���Xׅ�S�_&Y��'���?���`i�L�㓷���!X��]�gt,��$����%�UЁAk�M[L�]���I�h�%���4֩U
��\��C��1��QI�N^2�,:�,�N���͟��a{<�}��T���tT�.�,�!������v�?����V3�5���I?�0�LS�뜅���t���{�7���J|HQ��/���������>��8І��R0F!�O����P-L18�G��4�`}�.Ho����!m�4� A�xI}���!�h�K#���_�{��r��C�g�NA=|vCG���W���R���&����Ҳ5�_9���LĎ&��'�ar�x��W2�D�����P�<W�%srJ����E��bO߄��L�s�~ٵ�k.��oMT
 JC#����Z�o<�\���v�i�k����!��cE���mtHd�Ҁ(�0T7��r�u�ި�f��#�Ѝ�Ě�?M�*<�)��]B5u ��gO����%`.G������~v'W��B�lje�a�Ϭ�{�T���k)��ǟ�w��k:�k��Υ����6*������r]O��$\��6��A��9s����+h���®4�)oۂ�{b���Y��F���L�b:���49h�\u�RA�C�
��E�# 6�/��:Er�)��V������`��������hF��M�� P}��;������M5��l�B���?�H7<��ۄ11�`c�"JN�<��	�6˷�5�8Q�΋�k[O��-ē�c�J��V�"���Jg�m�{[N˻�b�Q*��-7�