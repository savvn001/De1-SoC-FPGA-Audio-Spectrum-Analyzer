��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�vl�5�X���N~v��N���g;�����&�B5o���
R��X��)�>����)d5ň eg@.-N��X8�Md>�H���dY�I��'�l(�a��A��������Z�h�x'=vl�[v�Lea�Λ���&�/�X��.RQo���g��������Ĉ��`�؋�#K||�������S�9�3�y�D����{jw�̎um<��jY�F�G-\�n�U^���}[��m	����t�c�:�FZ5�a�?)~ q;j�HY�F��3x�׸��ޟ��tJe�8!�(l����G��H� d,Iݺ��[ϔ�0o����w{DBZ�n��l.HzA]���N\jF7�.����m�u�u1����9n��*r80�V^L�,͘�&��~�`t4Q��V/Y#i��jK̒b�}U�b����wj�V��v9v;�1���W[�������m��]��z�b�2���\ƿ�e!��{(�������Ƿ������X���Eߐ6ܶ�^�K�TE�8��չu��Kg,>1|n�r7����B��x��B5.9˗9�5S2T�)R�lYn+캡&4�%jP2�Y�>��[n�X�zS�]+>�~�.�7S���y'o_�����3��jT_�R�m��-�̱#{�[��h�ڭk>�ݮ��~���� `3d$d����CGH�����bg�я}�����W���ڇJ"hŭ�;�Yt�Y�Wք���2S��|}fۺ�������9Sv&2Q$��-ZL�՗U�Bck|F���£5ݏ���2�Qp� ����{��(R��,��,�	�C'^���7��k��ߋС�NH:uA@T�^� ;~;���2��v�>/�݆R2�L�lX�򡴘�U�e�^��43�V"�M\%Za���� 4Sl�%ܥ�����חe�*����,��*��Z����H��n.��:��+G�WG'��W�V3�����k-��y��h���P�N����M����ծ���pk��C�>/�hsu�{'��#�U�e|/h�CJ�[Y�3�_�J�A�;vR_}1& żT�bo��jFm�I�H�-2;�b�Iy��ږ�XUWQ?��v��K�*#0Ie�x��a{v�ż*�F�Ÿp~�Z
�=V������ރ�u�D�3��n�F4���`^������19�%M_�`��f�o�nyA��MA[�}�p5�b>>�D3����qeU �u��Uk��-		g'������&M.�G�!.�����d��"QP���c����"��G#k� ���!�*~*W���U/J�����<�|��o��O�҅+�KY*}*��U��\|f���/�6k���C�%D�ϳ��;+����T��0|�=�*I��O��½飴�%�/�ASP"���?�&�{b0xdԹ��������<k9������¶�����d��,�1w&׊ �M��9A�({;�n~Z�����#��NQYT��Od-�>�V�R�]�Ey���tzE�w3�H?�e�&��RG��6X~`I�c¼h�����Κ����se8:� }.���ٸiy�XZ��D��ᅢ��k��o�h�C������0���ݱ�E+�8�C�ԗ�[��2�M%:�'D�a������ْKH[ē�"��^���g�%�1*�1������-�T�8��38N�eXH��qV�e�� ���.#ӧ�?�B�g�x�����_=v����DI`����C%MX��xVU ���$v�;Nh�v&��p@�����
O���5�.�b�I�v�5��P�l6��!AOO�� ��"�p�2x;t$ڀY���^�w��x����X��~���P~8g٥�Ug�l�%�R}<ɾ
�R��zѐ,J�V���lM/b�6��_J#�,,b'X���!��"y9��#>څ�U�cB�s{7���P0^� ���5��� =�/T0�-��_&o
�G]��������>�b;�U��V`D�Ա����T���t國���d���\��l�����+&�e(�'�Bc�#�;��Y8����@�[����!���p�w�T]�"���4F����Fֿ3z�H��&����I�4n������ͪ���>xg�$d�����0%�_2���~Js#�#���M&]�*	ﺻ�0�؇�S������a�A�����6���8^n�L\��!Bx�me�c���h� T�&���,�΁�H�y#Tq����L[M&7x�tHX���+���O#�R��8J����,}l|ogfh@b@{ҕX�y�ϼ'�/�m,�Z&��G�}�Zm��N�nn^�%�;�k��rgӗ�0W�䣚��s�vq��M��|p-��xd.�����n0(�/��M֝�~me�?�N�f�4����ݭ�2�eapН��f�TC��*9o}�m/?����M T��2X�$`�>w�p�g+P��g�o]'��1��4KQ��1k��Wډ���N�;i�<�}8E|��5��:�����n�L^}��蜿[�fR ^��;�r���m,Ya� �LD(��0�d�(���E��#HK�_���7c�Һ�Z�Ҷ���y4,I�����z�,1�(�fA1d��Ġ���&~�ɰ�f�$cxƽ�/)���I�x����.�:��n�m��$~j�9jP�
�����c����OѸ>���W�,�ü
lQ�Fo�
��@�Θ�o&'r�K3����_0�3�ˑ~�qb@��f'���X�j�*V��p�D��4�H*�u{������t=��9�4��lYɜlg����J�[���	��{JwH&�����)lEu�9��OFj���u�-ʅ$@�4O��^	i {�r8�e�}�v9�;��Y2�c���}l��A�_r��%���p��kIR��X�X*��a��w�+��aUH����7����R���F�j#%�xy*�;YŦ�v��.9	�&pG#������x+^��fZ(
$�����+PRb�\��Ba���$���QL5��͵��������7A�������Il}A�n�t�{���V�]�*�����0��]�_���?v�)�:�����4�;���q
9/��;x��2f�]J�xE�,[o��6�qy%p��}�]��xN�2?禔��d$@�0�F&N�#�W���e�6�LZ5zx�4=�f�Bu2��ZJ�4En�)�k��Z4���7n���7_���,M����]���-(����B��Kl�{ǁw����[ؖ���^7@35���<��H4�7ށ6n*(�a�1ui�樅�	���)��F�݇�L���ȸ��,�s*��;�@��G��L}��W[�tU÷��*��������+;�%�Q�����z>f�ˊ� �h�;.�2=oy���a�YuL[��2�� R<n��ү�7�c�7ӛ6����`�U Va@��"�|rԚxu\��o��ꨟ��E|0v��(YAE.�Bgb:���lym��E����}7���3�P�;|�$��q�t����E]�	;ö�!~GA�!�K|��-X*<�����L�shbƋb}���	e:���c�^+)gx�Wȸڳ�Be�{ [����2��7��^�ʛD����O]��-�pK��?��94s�����=puoE���{�߿n����	�A�-bn�a}
��2�=�C+��ⴑ#�a.R��ޅB��թ^���i��8���H�$�G�? ���`��&s�����W{Dl?6�l0J��^hQC�e|�}�8ӦA���6\����fb���u���#G���=]�,f��/\I�{�iF`��*�nfBw��Hu&�x�~`��]#�B]Y(R ��Fe1�O�y�G������ξ�}!B8ȉ���ƩZp�哙�S�ȼ���ۣEA�=4� ���ü:�_jf��,��@��?}~b02!:l��!�)��B�0��s�M�3���p>����q�*{3���0����wk���x%p�E��@*��l��l�M%���$ߑ�vjp��|��Z�h���e�㱳(l�K<�8�q���'�k�'a��h/�(�G� cW��������N�-���NC�vk�u[tG�)�����l�݋�KqN�F��%t�t�"��=�!�b-/x{Jc��mSڿK�>,��_���î���~J�S����<��\K�Ⱥib֭�Rr�7�
w�y���ų_%|,�dX^ǧ�! tW��Τ籕Hڝ��;%B�$�5��\<���1��Ru9����$�),T�+*bs<��.�ʸ́ǇC�)�ؿ��zD��<�t2bdka��eF�N��Q�����$Mɰ��f���I|���?�k��3�{�	�]R#�\?�Oa8���ʫ�$ԭ�®K<�yq�|�9QV�u��,��?��Z y�����S
.�\F�+���g��s�H���5�́�13{=>?����>�[�N�<��ɫK����������wuZ�¬���2W
0���I�ʊmb����*�,��}M){�8��)������Aԓ��"�H��D.��9c��-��O�G��;v�u��+�/�d��U��Q��V�1e��ݟ���[b�@��eւH� �*^s�.�7�͑�,�${�j�+�k�T��Wg,���o�ZO��|&fx���@���d�Ɠ���m�%G�[߁ɶ�/�����&���AJ��� �e��y����[n�|�س��oz����%�.�l˽�aT��v�1qL[�_����,'�,���r�v:׼��=��h��&M���?0j$��'y6������'S�����tڣ��Ҙ�lہ�ƿ�I��q�����o�PVq������[D��o�@?����7PVU���"$�V�j�/6�D�˗@� �3L�8P�AYH�̟o�W�ÞTw��YYZ>,!޶����^�?X�u�� �ܞ����:�P����^�vi����i�
��Y��^��K��� �(VJ�	�U������(��:�xa��D����[�wD��I��m�ȿm�������##��{��e��ɨ)T����J�x��srL㒻OT��֧z #��5�!��D��s��ZSv�V?�e�uBt�b>���t�W���_f���3��G�q#nr>�_ٜ��%hN1Osk{���U��A��$�9g< �쑔u�;�]$��\!x� ,�]��}5���G\�(C��e<�>6���������V�5}0�>��(�@���x
�C�ɗ4+�.���Ő{����Kهk�y:MQ�{�S��~N���YX꜐��yd���JS��x��� xw��"�y\F^q�w��>��?�lP�["T߾%�y��u�	�����.�y�}���kHD&Vh^S�R*�Q �\R#��N�*)kO&7��WP1�VK�����*�i�k͵��Bʨ?6fp|�	�c�C��&x.�N�E��rw��zR�_�Rl�(����h�1�in�=��c�?'�s;��Ӣr��e����\վ7�o�O��rE�y��ZW��,a	�)2F��!��� ��<�,K���4�X�̙N!8O'Ja;`Z��$��͕@5@���m}�;�/c߱G���X�4 ,
���TZ>�ێ�b��_y;r�[����_R�>nh�u�����H��P �2����N��?��U��7��e�3�$%o��� ������҅��ġL�[�$����Y�m,��m9Ë�!�797�^����ń�,ػ�_��R�A'��rꔭ�~�����q��XG�*	Z@�;��GHU��JL�_��r)�9â��)Iw�&�aX�s�=��d�z��F�����GEћ���v}����e]O�z�!N��̺�Nے�@�݂{��0h�.���j�K	7ƃB�^>{�|x�B�<)�řQ�_� ��<�5A:�$]_�Vݙu��
�G�C�2h�Us[=�{��F