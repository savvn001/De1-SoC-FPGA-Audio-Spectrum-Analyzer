��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�	��g��R�6����c�l-3wD�L$���E4S@�m��M���צ����T�]9� �R���ތ�����ц�fZ��N��ׅ���M�w�JX���bӡ�t���ksm�Wtp) ܆����\�q1~%E�~�	y����B�^����z���(����Yvȓˍ�B@���l/�]u*1���8�TYץ�#�z�+1�:8�k���z�� 
��7wԏ��e�RuGWq]���Y���O!٤��獈��GsCAz�.�h�-��!������X|O��-@�Ru0,P0�յ]�ąnᣭGM�/!kX�!{��G��'��&�:|DC��b��'#VDɢ�l�o^��&�b>�'��è��Ճ��as#
j�҃iH��)��m��n�S,L�2�x�W�.����כC�TZT��¨g�	&�f�v٬�}�9T�]�+�F2�ca�a�����5B<��V�9a�#pv���KY�y'C�l��M�x:WNٕ@��D?�F�l�"��Ve��h� Cl#gM!�t�Ӛ�����B�c��G��P5|���T���d�����OZ�X�c{E�=�I�/�y������1��w9"(1�����j�YT�n������bI�t��;#0���g_(���{�<�wB:|�{'4��[<�	���n�V�H����+$B�M۞��U9t�qOߏ��1Yr�)	�����z45��� C�M�u<��*�������<���0����>S��G�'&s���'��U���7�q��� �D�����F+�5��s�	ZA�	�#o`g��zd��_�W����yN9J�~]���7�Z޲k���5\U������������N;�P'�im���b������Su_�Q~)_!gFe�tO���ix���8�$T�y%4ɐ�V�"�����ꅾ��A�����L
v��m�m?S9.����}�M��Ѡ_��kbˆF;o���=2Q�����r�Y�Y�QS�"��h����W��#~��A!����U��x��>�T�V��M����1�o�0l��H����ojLݵ���T����}��b؅�wP���� ����X��Ư�"��#ܸa暲������j٬Z69�X��FVHIZ	Y�L�;]�b;>�B1��>G�b��X�2p̯��� T"�ż�Q�1��H���V��yb�=%�ڦ����U+G�K��u �lksp��=�0�<��ً��׌�˚jU����H�+x��A���S��H0G����L�̞Dڃ���ڑ�ß�����?�w8)��7����ӵ��׷��%U��}-b��x��Z������ZM�w�T�}7U��f�;��g�_�&X9K���솠{"1�U�vs$��ob!���mԥ	��{�/.�Z��o�ڠM��������=ٿw�,���E�}dADA�ܣ��K�WN�=���OB�����K�Y�q ~�nw���N��Z>Nԁ,*�O7s�燨�4r��-p/W�J{�M���C�2]��b�>+d�>��ϛpK7�	�*�~,�-�VE���������Ef�EB��W���ȏ'g-I�o�T�[8�����5
�ߨ?(�&5eyQ�t�Ȉ�t�d�;P����d�xxe=8�&�W���v�&l=\5�<�u��Mk�+�iG��S�;�g����
�� ���!D��[-��	�������hf��u[ٽ6�U"�%x�Ay���.0G��� �>����>�R5� �|f��f���B4{j�I�-Z�A\�V{`%�K;k}���dc��b�F��%�����Kz�x'8}�q�0G2�ۡX�h�K�H�րg�������؀vJ��`�1�� e7:ͳ��[�L����o.7d�v�R��L�j��GOu(�+�	@�;�S_ouM� ����c�	(�J'�[B��Q:�Vi��U�
�� �S!V����q*4�TG��!�@��%�dv�w�%��5���eQ��+�jDA�8���(�*�F�M_o�������7ThR�vF^�IC���U@�.a'q
���� ��0�5`9��d�,�D�%BB%���$��N��H��5�e�6���u��c���])��p^�=q�Sy&�S՝�g�B|��"���0	�C�"��I@Cӈ�Ht�ۛYg�$�s��8v;��UeK�	A�T��.��~}�stLT*B���:�����|@шjACj�5��"Q�%��׋��4��QE٣t�|��O�QF�(S�+ZǇ,��փ	�s�U��5���烟���g!����=ʫ�@��ߣ���;"�5�_NZ?�	[pD������"�4�/Bzp&أhs�nt��c]G����m1��j\P��&>��o���F��q8��}�1Dr�1{��� xq�����a�Q����L�H�2y:�R3����A�q�=3�r�*������HTK!9�v�8�*w�@(<�BL �\!FG�8��%^��]�������!B��A3=7i���8"t�Pd�R����DH	Bח�!ނ&�!�UE����� Q�woF��,���m�.M^=p�~����\n�ܙ(ر�Ϗ"���\| �a~c�n��;����d�
��_�g_\'rv
��Ͱ�d�����C���5٭$ԕ&U��+�8�H�x�k(��4��n7]�u�y��Q�Z����Y�!ԕbcC��}�늹����cօ�e1�p�i��l>��(�̇�@�6�؂���{�iH�=����!�'��F����~�-iF�s�aQ�l�6�3��MY��FIA,�Nz��0LH��#~�i˽v������H�}]p/+��&XT��\�Wou�a���)�Q2����Ҫ�:��~}) sYq���dȵ_���p돝pyl���l{��֧֨��PO+��ޢn�/�%=�q��KW�J�0�$c�FգJ'���H� ���tI�`�j��
d8G�<�r[��/���߶o����-���kzd�-��s	N��]����t�a���U�]}tS1����96Id�VÅӇzU���W�#�8�?%PP�搜5t�Yr�i�J�"�Ko=v��d�oh@�
ySD����d-�;��))?���5��T��� �[���v��,z��IKo��p�T����Q2t�b�����l���\ �
��Ɗw�N�.\R�Uu�K����竣|��_'s���>؛�ܯ^ю�ȇ�ѓ�4Qi��gs��|��10�Z�a}Z��IhD�'2�m���qw�vζ�����ﯪq���)y�IŹfs�!%p�����Ae���<r'�;���+����*\�"��`��^vW��e�Z�%�P�0Ŷ��������������eGj�LC�Y�3Ji�w��g��5Ҿ�
��]�ӳ�i��d�<��js�;��K@�X�'��8}-���A�!�p2����ɋ�����h��4�.~���=>��Q=�6`0��#R�a@����Uߛ�s�b��.�8��}�0 �;>�2��S/��$�j4ZWC�2(|�ԫ�ڣH{�~Յ�5Pi�=�[XӉ�V� ��#��O��z���S��o��gf�fG�>���	S݃��n�]k����.a��@,���UNp]Ǭ��ϫ���`��,A��-}rz �m��9aFsC�����	�����h��E�u�\�$b��v��͂;��{�s�8;�����D���y���Y�#r��?�Mс/vb�����H����.A�Y��^����V��hEw�+��$ c��oo|��o"������t��5Z�JH�D��P#H�LW*+i������2�,��Q�A�8x�����r��>�	�ks݁0Y���=����sV⼯I[+P��%��z�x?��h�=P��1�{uR�RI���a��#�zp�I/�7rgR�t��/ĵ]6�Wơ��g��Q�A�rOi�;�����_=,�b��1��[�y�u|�T�ݓ]��m�q�������V*��%��v�ѧ�N�2P@7�2%��H��)^!p�T�	��\�+��G�s�}�E�\C�M��-p�vTxl �b�>���/)�Sjp�<m�9n�Jh��9m+sӚ����vG��H����"��O-���q
ih�:�.HH�r�V���[:A´T.�{3�ZF�v/�{��� "����BX�N���X9���c�hw�hO�����p���A�X�e���h�NY@(k����j�oO����z�h�9����P������6�}^m���kŌ�%��vo���*���s<NRE��9�(�+v��j=oI"~�3hW�҃?3�� ���s�>T?)�na�����`"-{���-��j�C���Qok��\���y��Ȕ��;
Ә��\�<0ϕ�
n�`����+|�jh[��z�NM�I�,�Q�yz�K�g7{�^��-'5�$�~�?ڂ	�?��_:'��ѳ��k�b� ?��ݣꋦFgpNj�iF������\3k��6/�WPC����9y:>r؎��_��*�Э0����/
u�h�A���/�G09tgѓ�:;����9VK�X�`���={� lV�#����it��g �d�6��Yk�(&rö��l�mZ:f��=_�Ե5�����`�Z����O�������۸��������H���K����&��ŧK�CH�r��I�Q}[;!L{ca�������|O��|q2�Q��v�4-9����L��!�;���wȰ� �P�&�V#�M&���W�
�	݄s��0��^��V��F����D��e�C���Qk�1�SAZ����-�.� ׎}��7&U�$�"���%\�.�N���TP�Ἲ� @���C�@T�һ�X��n$��F�C?n�iV���Pc����n�����y�I�n��4���Ww��Q���g뜷EC��H�_T]qm�)�q?�9u��P$g����q�CP�и��H��T�Pˢ�q�YKXb�?����(4P����ᓇ�ڇ!���?B������-�\Ǉ�1��鴜�7�7�b^������R݄>��PQ�@�2�$x�w>�g���0���O-)�/�(�kJ!ܲ��R�~�̲~�����v��%� ���+j��3�(���ڰ�ҺZ;_��	��>�J�Cm. ���e�	BUFo�u�\�o*eJ;�P5�*�~~;n���h������W�e��P��"�¦xٔd��t����<P��դ�݂�B�z��X��
;��ٺ$?��V�BK �Vږ�cqK�#���M�_�
�����
�T���F�_Ωxs\0�c�2�M����lVHK�3���O��r���x�t�B"_�0�:Yߞ�P�6��U�~�r/?f�Y�ܿ���&�˻j��<O�p_�����p@i��L�>Yz�[�NS�
G�-����l������nI10�xi�f�g���5�o�q;0�M�L�vB>%Ff�V�%mp/�s8ʾ#q�%�gz���P.:�5��@�1C�X�4|��%�������Ä�Ai�^0��-L���h�غ�DT��2oh�S9I/Ь�:���
�Qc��<׹��B�z�8�s%�uU%�l8AH]	pl�˘g4��>69
QR����A�c���=�۸[y_����NUp\��-�i�ed����=���^����������N.-�p|1~�ڝ�RP�i�bF{4J�95w�Ta��n��͔!�ׁ��Ζ�;�n�W&�J3���n�]��@����e�m�$�V/�?�� 18�%_Ѷ�� ;=7�����%~g�a�-�⨺���}�`��8Fw�Ppi�#���������8��l|7/n� ���ω	�[T7�꽈{����� p'�����7S�ώ�b��Ip-qܾ}s%$��xM#��-����d%�GW���T�e�Cǽ�Mu�D�ծ��%ɕ3�%���N,�oU�����H�w-6�VR��tN҇uK[��)�T	h�4OE6���6�9tѳ�|�g�!��n)k�8k�J_��W���
�mv��*��o?8ς�iU�\��T:^h��`�ڢ{�]��p�̑�n�
�?�/N� &�dj7�W�q fJ��1����'�V�bj>�9d��e._l�Mo�x���uGu� �\a}*�}���Q���eǖ�+o��Rv�G�����8xlD~Sۓk����cT5�����n�?���z�/js,�:�B�����US���� 1��E`a��B\)��h�����WI����Et��(��_i�T��<��n�;6kd|!��~:eDz����A(㩧�n%;A8�1��JWB��t	�$�b��TD�=�e��]�F}�n��U���T�^
�QxH��1[9c�o�w�q$��=�,�f���@A�0KA,V�<���P�.�H?�>���D�b��b��G�����_,5JD<�ҚVM��Г�.���5{Ƚ��u ��p[A��!:�� �����[TKJC߸*�6��������-u�%y��Y
�
�+������8=d�	�v0��[��2�y�gl�3uf���|����--P�)פ[O��;�������(�)f}J8��aҹ'� w�%}(���:�K�;"GF�����`$��K��)�4?��+)Wʯɂ���S{�A�fp-��g��&:�;9�U<Tmч�U>X�&Q?��B�J�����I��Z�m|��H�Cs8QK������������?�\�lU�
�p�#�9oq��?�s�#���uJ��9/?e��F�6�3tL�!�w_C��;�еN���l�J���h�'��[��@�D���[����ĖO���=V�b��ju�L4��e@�o�!}�Y�[5t���O�Z�r�Zv'�M�w����!
���]��d�)>
��ZZ���)z0!�ln_َ6ϰ-/��2y�8����+�`i�@|q�bʮ�L5�vv�]�r/7*X�h1�p�'8G�E���hp��X�I�?�0�OOv�ԩ��t���w��ċ���S@���gT�z��^��7Gjն���A�B���z��v�Ғ�~!���i��f �K�}�z��')d����N6�ƛ���*�����\�Y��S"��y��	��d?���]�a�Q�L�$�T����pW��l��G�oWO7���Qh#G��,JbG?�����?�͍�[0�)���M,����?���s/C�Ű��i{Ѝh$Z��[=�J@1+t��5�� 2��E%?����0.]�,�g<)LQc���c�[D��
볠���P?�ǌn��.�W
W�$�ӡv�r�@Eo���[X�@r[��FQ` �O��F[�7�x�[z;�Gw8v߻���Ó;^�PQ��4���QX!�G�<0��a{ n�
wtQ��ޭ9�,����r�P{tfRW�s�q�2����~��7�U($T��``�)Mz��(@��qZQ�S��{���V���n����c�_�-w��la�D}X\���_'��~�8ۂ �� �)�?�|�?m�/�:��&M��?i��f��#�ߵ�
�lZ�K��q��-�ҸN�B��I�'��}�� �]H�`Ms��������U������h�?�W�����,��yfUx��S;�����M�����}'��@~>y��j�`�Z	�$TS��{��J�&~^�ľ��B��=��bxM�;˶�� �T��OH�R	Ù!d�'��*r�h9�/�g�㟴�8�|��X���%����l������O��ҙ�c��	Z�ʖ6��b����Bd�~8X�����5ܘ|�+.��tK^K�	�l��ϛ���W��"ߠ�)(�b�v���xk"JMŷ�+^9�귀y�p�ٖ��L��ߜj"��;���.��.��f���\�	� M���:	�]I���K�&��	���^c�<S'��V�zG�cX_.�R�*��+m��r쉨��������Z����V�]�CI����� 7\�n��Ft��:�"��t��3]�a8M�U���ȉR7��/I�*-萌s'�1�D�cgTz���ީ@��t�P�Q8!D߫C�Q��T��|_YٱF*Q���NW�� ���ݍC�5��L�����G
�	Cѵ�b��5}�PR!!������)}��� ���������+�S��^��`dbZ>o��[� @�kic��Dj4�������7'��zf�((+3.��Ӽ���O��\}�PQ�T��ua#�'XZ�̜�����ɲ����A�#M���BS0�̶'�n�Bn��a˄I�����U���-����waоd���q�O`�/aW�HV
��U#����ri�Ln��A��D�~\�[o���;����K_�TF5cǼ�Zo^Y-��La�p�>�<���7Kv��r�u�:ߝ]���V��y��t��ӗ���@;�<g)RBȪ��T�Ⱥ�q��d��cY�S)�V��4=I�_��J0tII�T%RBɌ��K�F=�2��f��W�\	Y��D�6��Ԁ�H�L_0�҅��H\	T��O���,e 7]��EꤓT�A+FM�O�ę���1.��%Fȱ�!�������(�+VpŴ; U�  @~����A�"I]k�T�t��
g���`G��Co�D��>ߟ�����Ļ�V#X0v�w�Yg�A��3�3K �a痫tW�a�W�>��0�R��}$^?�T;2�r��d�# �'H7����_\��m�w���⾨�؄���U i͎�qg�m�%��w��3xɾɗ&��p2q@�p��k�Tpnb��#�c���]�L��U��a��.�U���f�[�
יr.���P��F�gZȁ��\S��JMX��t�R&�LZ\GQ7����I�ɶ�t醈h&4��� ����?�G�>~��� � �A=Rʟ\�[�1y�xLv��23��㊘�FYy�(P-���Jp_ϋ��}go�u�lF����)Y�[(5��8߿�	Re�c=f|B�Y[ɺ�T���!��.����̲����F��\9�9��bwՄ��=ε�)2V(T��2���j�� Þ̖�pT΂ �|4�"��8(�� ey,X�k��e����߀��k$2s���q o�V{1o1��wC'k�:���-�Z���q8�����q�z����m&�B#~t�o�}}��IV��%c��@�*�h�gI�H�"�ğ��n���	�Q��a�|�~a"��.³�䏽#�t;i�=s.�@?��!����e�p4Hy��Έ�`ޘ���W���[�$��8]~�ll�~�Z?����Ԙ��u��BH�5�Bb�T���O/,Q�M"��V�.Fe�#ϊ����.��5�b�kk��~y�V\�l��|�������:|������yb_͎��P�~5�����w+�)���XԷ��?�"P��Q]&��*��'#�]����������2��XQ��}�.-�]���+z��7�#��Kc ��g�š��P���Vi���Y��r�q��Ҳϝʘ�,��Q �����B;�0ʵ�F�fo�"ųa}�a�e(�`7��N�6�=���g�4OS�X@ ��s�e:Y��A�I���!�Er�.����A9���a�0��ߚ����n���\TC�^�����5$,_���(De�F;�b���@�������:����P���>�2��t��ޫ�"=@P�Yż�D�o�TU��R�v��(��AǤ�_���$��40 UH4�Vp�s!�	�������x@|�A�ط�4U�����z�Ip�%4a�%*���t�� A�G�x=�<BY�*O��Æ���FW~o�l�����b�P}Ħ������\�ӯ%W�O)�s�ť�k���k�i����ƛ^kЁW�+XՂ�dJ��I|z�ոP�N�a`���e#o��?�`�y�~��LO�(��_�{�٣��_>U���>?-ۀ���W������ϟǙS��*��9?w��O^̤'�F`� l�`fV�kb�IF���x|iPr�͒�O3�f�O YA�O<Y�$�b���3S$;�'6ڠ�>��i�x�Z�U˰�-���D�␨�X�S��(�nSP�EE!�@.h�p!'�Sx��x.P�:��N7$���I��vj!Y��D�rjZ�,Ter�f`g�!l
OL��V�4��g��EE�q\ge~`��*���yYez=�)\a4�b+JՊF����u\�g5cx��X5��x3.�A�;}f>�a�xj�k�:�N��C�_RƲ1Pܓ#�n��k� �bի�6	~!�,`<j5Oc�����qC��z�ʞ�j���E�7O;�D�l��t5Jbǉ�T�A�K�hn��yo���:���y*��<M��/;�m}U I�(>����Ҟ��T_�QG�z]�(���
�w�A/gW�d�lO��n����*�fl�R�Ca��aMq�(��/cHiXn�����=	7�9���N<��u��E#B
_M���}FY���-�L
4����h��'L�'�Ǝ�f�[�ք֬��g���@�c�O0@Y����l���_�ZI&�_�u)�P�`npDHS52�֔6�R}�5O�|��&�NT�N������L+�����|�Vy�I@�M��C8^ �Әvή���DD�0������A|8�m��-Lc�(W�Aj�������Ys�p�q:��߬�I,��iD�-Q��\b}���4"$)a��쨀7���ǡ��2w�.) ®��WU.�3lly�e�8nq��P��T����T�N�����ɤ��oxG��8n0��w��@pڎ%�97�̧�H_f@m�ˎ�R�� ����8�e��n[��6H�Νa޳�LW/"����J-@R+���
�ucمXjh`I¯���m�\}�`�5���x�O�v�ȸG����8)�Ų:�����
��Da}ծ��t�"����kww~�n�>�]�E�k?&b��Z��
$��~��`�T�"-���JNIp�Ӊ��v�r�;����E���2��F�/�{c.2��S���1Se�s�0o�u�-����<�D��׮Y��*؀W�ɥ���N��Χ]��\Ty$�fs�I�nx�oϾ<DL��c<'�A}�b�湘���8�:����L��/�P�a,�;v����h��s���e�����$M���JgU���̟M<7+���֘i��Cs����ۯ"�y�v�uӚ����g�~��G,fL���ch�A`�S���t�FT䰔\8ݤ�0?�A��?�95A���;�y�p�Q���/�=��������b0Əq�Gj���9-�����!l1��������8d�	��8�Ũ����"�~Tk�E7�w+������d74;m(��ZH�6ij���"���'#��ei�l�G�֥,���{*!hġ#.BS%0X�+w�ހYih�;T��O�+�U$�zn����[Zk��^��b�`������QX���~,D%�p���D�u�ƴY��\�.r�a_���i�]���}M������}p�*g�<q}��!A(��4�
'W˱�-�!����`�u����$���PǅO0�w;�*Ӊ���)�� �0]�i�N��������ny���56
�����a4��9�q~p��L� �vT�ea�w�W�Х�>;���"����cs���' ���-W+FՉ�L�f�s���{�e�qd�~�%<��(�jgc�6F�F�����x$nK��Ɨ	(ʪ�T�X~$c�$�/�����_��P�"ۀ	��d��NAj4�$��2�~wQ]1�r�H��ξuk��m!�dM�R������+���|m�w�������|	/!]�apN �پ �t|!�1��S���ܶ_{��'_/(���5�c��Y6��^,��GJ�سJ�sA��^�vB��m����hC�j�,��ֿ��+���\����KJO��]T�Xנ�o�$�E` y�3��GT_�JTd&��i�l`6+�<)}���%H~�wͺþ%oM��uΦ��u���i��u�a�<?��av�a��[��L�rI���*7а$aQO��4mJo��Ғ�ʎ�qD�s�8?a2B�=�=[�PQP(]-��xJ���
�7����ޥ��r�鄜��n�L�p��M}Bi��Q �"ީ���Ͱ �i��3�HkZ�!��i��������5�82�wz�Ye��u&��F8P&j�(Ms�scI�ˢ�H
wA cx!2����T�F����(�ck۰%�)�1���n�)m���KN�t1\ʽh� 	h(,hR|t��
�o�"F�˖����5���
Rk�>`N��e+��[�|���w��2����(O³�0�`ˀg�Iws\?�D���μP�H�l��*�7��D �� ����Mv3 "��lЌK)4P�����9&�6g<�:��9m�{�>�����c�c��D�f�i�{�V8�?��Bw�|"N��㗬Z�#��QA$�E\g�$��'����(d
�2y�@(4���Ǳ��sm���� �X�{��b6��wx��}��isdTr�}=�U�o~�۹]�quL�]DL&���?�������0>Z���\�P�z��S�Sݿ���԰>?$�r���ϾVDb7��J>̾�d�4�����39�r� ���;��v��D�}�-�C2�X�q ��������lat,�k�=ZSu�����[}�y�@��4�or%����,�6_���!G��
rLgy�7X&]"\d���lI�>,�����c��/�u��Ѕ��Mn*fcܑ���}/_�i@��T|�}{��o.���U��'8��ބ��+�"@�EC"�O{E�V��R���x�Hޭ{=�]�w��!��jgR[�f��(l�b����qA��o�^�\K5�}�n�.�j��n������W���_���I�<g�F3F�C�3��*�0����(�3�G�c���k���jJ,U���@�a��n�����9��3��������@t�7L�pj<�>U�dͫ�i����ѱ@0R���|�����C������Cf�4K<1�����bVP�?�?�����^	�& G�KKcB1	����a������r!i�zI���h?���w�Аe���\�a1_��v¼zרK����t+�����������C���������A�bG���[	��p�c��8=�]�.���@��˒\O!��r ���@բ�OnT.rFǞP�����z��v� $\]f�ƹ������z�v�*lͻ�-T3`�_��+ez�<�q�wh�8~j�rCȵ	���.�C0X��kiY������BUt���Mו���<�ݍ7e�Äc��aq�9�Nj�cﾧ�(>y��h�\b�L���o�ɇ"�]a�'"�����`���X+{x�>�*��QV�u�
��;�9�#�5#�A]C����c�&����e������@��43�ܯ����s-7p�2�N��z�lL�"�6�?�똣`�8ȾֱrV7m/H�x"c�8�����\�m�|k���d�j� �CXi-������q` ����X���T��^ƫ���1@y��~�mZ��=ͭrA�_ǿ�E�v�k�L���E�2���q{�7�ŷK�3F�D����an�H�?���E!�қ��%Z��04�k�M�& ;����d����E�����\p�L�O�?n-.Vī�_y}x���E�ć��f�oK�.�|Yh�������O(�n�C���*^�
]bY�gb�p���$'f���&��`�*�D�%H"���z�6�F���(U��{M7L�I�S��j�f���ev�8(p���a�~-ڛ��-���#t�<%c>A�܋�]�آ���[�d���>�@�o5q�?��S).��!�����A�吴�Nυ�&��U�m��r�:KAV���� ���>��nЂ���if%)ᦧ�]l ����9e�~)�@,L�C��m�[9o�Z������&��q�>ƙS��GB)�l�����Z��1e}��u�0c�x��>
c�5i��1VG�r���lg� KZL:衸�!Y�9�<C�s�'��R�^i�]��Ʌ�l��U\���S�v�l�k~.�c��/�,F/4������"P�����Wc@����j{�,�3Yx���L��.0�-�����}-g���]5��\ن������Ӕ�jNd_��HN:z��?�jr6Y2��;X�gF�,��*�T�W ΒZC�C����o�<4�}T�t�&
/Mea�3q���r�����/�bD�`Nx��n�1Ay�<�R:~��%����� 6��S?U$9o�������|�0<�h��a��V2I�
+��$�);M�6۫y��s$<8��tx79��C����҄�I���meT�y	���:BY��%I�vl.�<�( :L�W�6�*�U�F)Y�ń,�#p�r�t1�H~�(0`�-{#�VW������1:����+^+2�kvn���>�kߗ�*TΛ�ԟ�<:y	��.(�)������_��w#��ΰg����߉��ynIW.4o/T�!�i�_Ւv	n@���� ׃����4��)���P�V������ʃ�+�L��R�xǎ��ci2E�D����W�w��G��>� ��Cn��������<�ʇ5`i���a�50H���Hʨu��ۄz'����m{n�_��wm��_Om��r�����f��Q�1�Ä����V>��*7�b���j�X�H��u�t�Ss��v6Һ�{��a�+_�@���9����2kY����S1 ��W(���7��� T�>���ֈ*�0��Ov�>�����h�q�e£r�.�Ā�v�zd78/Xq���]Oȍ|k�Z�ٳ���1��M
���_� bv9J�޷����r=+��"���lY�����0� F1�R�kŗԚ���t�����ĂPBx�=.j䣧.�xl��K�E�=��i_�a{������LX�E�Б�>vN��"��U?�7^��㏷L�47���j��H�ҭ����3����蚮 �P=���V�`V�+ę�o �[�����GhJb〕��H�)�z�.���)�[��>a���ݳ�6b���ؘdh�o$������L_F��/����-?f�y�zuyr>��ۣ���R�y��NmM��.R}q�I�2E���夊�$�R���kH3�H����7����M��V,�;Y���� ���RßZ�ؙ:dA!R��,<&>�+璉�s0M��C���\D����1��,�P�U�|������S@�=<|ڙ��u@�=�;�K�Q�����_ ��i���.�i�J��p�e��b'�u�4H��E�����6�E�"]��ۼ2\44��X�(��{�N�鵋	0 D ��7������H����왶��:����o/��c��m��x2L:1P��82;����U+�����R��	��Pܶ%<]�-�!���r�̍�V������ٙCJ���_#�H	��=��H��"��k.e��� �Cy����{��.����Q�
��щ"��cM&$.�q�����upn�y�Y���u{uKe�CZy��9!(jQalc9��.2�f�}E��鄭���`@p�m串��(� g�S(�ayM�}:�Cb�)rp2�@���2�|D�Bg�IF��7�r~��+ς��ɾˊ�xڎb��Gi�6�S������̊/�%6[�#�Xh�������X���ɧ"�-.k>EyY���=t��KeOq��tc�j�XUC�A�2���ɱ�L�v�[��u��ED�<�~�1N�Nw�e���s!@�`P2���J��`BX�ůt������%Vҫ�`?��=�������y�����c&h�X���by�x+(xtZ�;��W*�I\%��0n.�d�v�AMWK!e�G�;!g���ƌ��7��Vd���#u���3B��"���lhy�D4�%�GE{�r{�1��muds#ЬcA��8v�V`�\�����dY��7OltU�T�@G�zv.�0��rx�0�`�O\�'��-Y(�<>��k>��x情L���7қ~Z&�І����PmsUg��"'B{���°�G�dD�I�f���WfP������D*���=G����5f�#�	���B�]�[��c�0��� ^���5��&N[�K% ����uH(9�A4��z�c����l�0&��Tr(�βm�U�[�M�ōN�(���@ݹV3B ����׈Q'�L����*�4�Ю?Fu<s�\y�Ϲ��s<��Q���}�tm�uŹ��)�,'�K킮I�/t�����I�� u��us��zKm6�p�2���x�M �?E-,�:V�<LV�9Ԛy0��~f2wU-�T+�|	%�d$;!��	���	�Zm����v�)_QA����
	��u���(�]��2r�RHu��C�ٜ��c8��m�b���k@+P�TTd,AJ���������SD���@-���V����7���fK.h�� �`#9�̿����Y��M�M�������uOQ8���ƍ7��=UPȩ� �'N�ÝM�Ӟh�C��fr�<��So���V��ހ���=(�r1d���L�@�l�bgk����v6mt��Q����;��/��-�K^y�'��dS�Cz�_6H��y'ďl��,$�ޯ|E�;�z�=���r-�AӔ���H���co��|w��µK���d)�S�xۇ����K���[Ҽ׾�tD?�z�V�e������i&�A2s7=��n�lro��:��=z�9h��3~Bߺ�(k�h�έ���y�)R~B�S5f���G#�煀��q�b��!
�Z!*�L����:�z�BWd�͗��c�3��RP���l�I〥PX��V��l�k_�:Hn*4�ѳ|5����P�9��)��]���a]�֮6��?XS����S����z-�[?ۂ���a����=�P�4�Q-;Lg�9V�����U8��a^�{���3����O�W��ߠ��y!S��7��9��� ��,ɖ�n`�^�ۣī�Zd�nn	�� �� �їh'o�]x���~)�Y�Z���4;�!�ځ��%�t�]�'|:���2u�|�&����P������.Rr����G�_�>Ԇ�/vn�+��O��i�[��Kk�ԗ�@-+���"��l����5���`'ƾbf/���]�C ;�W���[弝 3�."�W�yy'�w����L�x�u ��1I��9�F|�^��D;C?7��x�y�[ ϢJ`�so��o;����Ꙍ�ݪ.�w]��s�$oz��\�����:$~��n��S��xs*��㋰�}���7`�8*��Oy#;�΅'R�Y|_g��G�~5Q ���y�o�)%�ջL��ٰ����Z�r���?Zg������EP�iˇ��j�ѻ����6�����N��33��&�s��?�[Y��u%<��ԟ� U���i�X��O���ҸOx���\�mjC�Fpի��za
�9$���g�S�*8�0�]ӧuEw��YBO��-�o �WA#�#�)i����$*��Yw��Bŭ���JJ����(8�`�/�~��KZ��"��L\��z���h�T*p�!N��o�6��+��u��aO�ld�<����F
"��6�p���cg1�F�Z�<���8�wY\���5�j?+�fS0�IV��ޯ�$�d)�������4�yM���nH��Fi�x-BZ��sw[�k�[C�`�G����>5m}�?�3�dq�*����_=��h���wH�B��b^�y��kx�LJ�_YQ�[Oc���wZ{�-�v�!��5I�oۋ�1=C�݃2O���)΋|��f�;D	d~	ӚG: �F��\?�Kw��,�S �k�$�T�u��ͫ����e��U�����O?�$�ȴ*8��]!�$Y�M��l��u��+@�W�N]��N9����$㧯�u��B������
ȳ��X�P���RSǰT��������.ԝovc�tf�C���sr����Q����&���vss���N�{�a��u�z��bru��2 t�v72�d3�FD�����6��o�fd�䟝_��qp�;(�m�� �D�n^���� Nqu]D���Ń��R���#��z��}��ŗ���y�KǓ!���h�ɳ;]��դ���G�z튝j�U&v�z��D{^��&]z���j��� )�^�V�ǳ��!�P�U�2&���%���S���s�>Ǧ�B��4v��b)�Z��
8e�+�L]~O��K�!,���2��V�cʋg�y�WAL�p���������
p���Ӳ�ڟm ��D������y�)2R��@���I�`�&'�yBB����pe(a�y_����<aU϶9AB�7MN r��p�I{2�j�ls��W��oԷ�<�n�r�ƀ}
Hh^�t�;}����mO�g�d��'�*qA��O��%��)��p�~���EI���N����/��s Vp�1�̚����0-C@�W�$�M� ��q��ن 4��s��^6�����wV�UR$���e����������˘����6]�No �����ʻ�Mp�e������e���=@�jbP{�0�V2�5���j�-�W؈Bx��5��ȖpBqmu8!b�F�����㔰��9RT�g3=<>y�J��a��ߓ������_� )�y�G;�����]~V�us��������&�(�Y�m�C?���������"� iThY�&��bf���@@�YK��	��d�
�Ũ��?��N���K� ���H�00����2Wm{�Q~�x*3�_+��������d�"��rrV̕1�ΊPJ�_AD6�N�/u�M�}�2�~ 
%Pmj���p?�A��x��GF���O|W�[֦b�GȤn(�XáK^o	���5��>L8]p�(�{�Lס�(�I^g��+�a4�{�P�l%;����:~��a%�=$�Kտ	�$sp�X�'C��jf��!i�qD<��#�NŮ���~�Һ�����@M�~�͝h��3��Śz,u&~ז�t��)<싊�L�nuS��?}uD�?l=�%@T�CiRc&��2�*"��2�
� /Ȟ�0�kb�E�/��awm��g���s���yW��o����)_(4M����
�C���ީJ�2?uݫ�To�^� *�K�0܅�@u������Za�.}y���|�j)�,���w�p�Oh-�O�h�b�~e2��v��Z��("ki+��P�E;���qrt3���bt�)�o��)61!�� �O��d&-Q]TS��<�1x ,�z�4V�����y��뙨_m3��ġ��j����Ic੒K.�i�ä�S�H�G)�h�{�ǇF�S�gd<o��iM�S�%>����9U���/y��� J�r������6�ؠ���6��#O��M���ݿ@���ԃ�{���ٖ;c��?VP���!¿`B�Vș!����������&���� .�l�13m>7h{H���6�8����cu��L���ɝ��օf��so˛q�h��dܩbŖ��v��;(�x���*S�r�!��� 3��]�b�h�w��ss�Y�-ڞ(X8��*�팟g�� ۊ�����:����SR������1Hӿ(��x�������?�$���h��qD �(
��R��S�/�6��K//�4��-CLk�	+j�XR�"�#[�$�p��[2Q���~_(�Ds>�K������>P2y���昹�A�l}��UT����,��ĦF�MG�P��	�[�����zllbA{2Lj�Jbh��#�V� WKp`�m��"FT �gO	��ӹ�.��T�������k�gȢNVYa�m���`PfuNn���Ka���a�xd1U�H�]p�bhS���x=?����p��exJ��M�8�v��+� ah.V�ld�8�D�f8\�N�)�x]E:r�[3`�����3��5���´�1r�T^�6G������p��ڥ��o�����Lq9�G�8��PToO�_����X<Z��#l ;�#���M<L��t7N���w�dH�=�F%����?�y�ZN��OZ�3���)fa(4�N=��Br�_�_j.yHN�O����8�Zͺ�\jk��v���I�%��NLc�PA��w&����*�?W/�����A�^�	=�ŕ�a�} A�qf=!5��5�$��W��!2�n/�[F��>�.-��&��I�8�G�3CJ옽�ˈ9�����ݍ$�Qy|��U�#��ܓB��!.�s��q`���'d�ȵ��Վ��aW�&���#�S?�6܍���N)�/\�+��~�����0V{�͑����[)�tI��宻[i�N���Q�["���QoB�g#���fh��Z�{Mx	�vG���L���yަ�4)^ ��ԣڝ�`����W��}�' '5���X�l�+\!��2�}5p���~����\,jb�
���(,Q�rF6<�]z��N�=> ��s�r�CHIid3�z�Q��Y"�F�Ϫ'\t��h�Cu�k�����1�0�+@>w^�gS�?S��'>�ۯ;�IhԘQ|`�$0�A��da]h"/k�^xCZ�UF��8�r�m�lx�X�/���:TT^.�兒k�[���2u �7S�S��_�}����x`��)T�s��-E�����V�>0U�]L�؅����qÕ����Y����j�0�M�l�� V�MZ�@	@�y�g�+����Ptz�׷��t���Ǉb� {���d4�����uK[\xBݯPÜ���`�<���葫�%�|E]I��r��7�K���N	(y�Цz+�V�}�
Gղ� �3e	�
@I��.Rc��3���T�����j����~l���Xj[sd�F*�Z�@�������ֶߐ�>�ǎ�ד:�,��v�i8����65Z�w8���Uv�7[�A�⮮VLBD�,��
�F4��U*�Cú�e�a�%��ɳ�P͑�v��/HpLw���ĭU?�͖�Xr+b��6����F��4:�,�?��
+����%.
�!�?3b^!Yu�g)�DsQ	�) ��?�t-(ß�d[}��T�E���6 �/r$�RS��Z�d���_�V\|�7�4LJ'a{Q�9Q���GM�q�z�l�/K�4O�k:�P��׾����r˻�j�Ԅ��b���@ l�"�i�Jc��$�ޔc ���ȼ�U�ڼ��'��4�ƻ>~�e_�� M���Ah��s(��D���Q�i�(�� ei�n��tU>���m�:T��	����tz\H�� c���cP��JowB|2
p |�k<˼DL�@?�A�$�Zo0�6���.�q����2�(8#�G0�ɐ_vѾZ�Z�,z��KߘE�"�[��"'߱����_VF(�?�9q��c9��Amލ~@���vCu3�^<3���)
�����|�uC("��G��{֖c����n�x%�I�@�agQ��8�h���L
��aX/B�i��|2h^}r^�b�_��' �7h*�w0r�3�H)��2�@�:[Uz'���+�G�w} ��#��l�U����b��ELL.k�#��(����ǿ�ZQ��:���['���$۷�u�jMx@��kPl)[��1����m�WP��#���:�D��y�8=5�JB�e6T��FG��{�V_�<�kJ;׊2�0ۈ�#���u��i��y9[�tb��W��od������_�u����M��yĬ��皟̖ܻV�ZvV���,K�K�`-��90��c���;H��l�w��#�,����P��ۚ-����"P&ru��x��P�g݉�~���{�E�M�ԩj��jUL$�����u��5b������+(zOa���K�/<��Qୢ���;�����<ĳ)�xnW��AX�1����󙶊�n*�ʿe	�R��i���c�~�l,YG&��U+U�݌X8�5n�zY����;8�²=Lb���]���h�	���Jq:�{"��7�����y������`��vF�������%�<B�,�]S�����+m��T�!���O��>�,�f�D΢�b�BD_���iD� ���æ���
�ϰE�?�Ph������:c����5ăv�����I'J=�pX�|C�VNҞ�P>��,�q��^i�3-�q;ѡ�˳���'w_�:��(���|΅z�o��I��c()p���;�<�t��	�g9St��&Uvـ�N�2���;�J�=$�|y�_0��cF�4�*jeק7˪�8���y�����5pR^����	�`�Pʏ)�(��g�ᇔ�S@��ާ�(0�`-8�,*/u]�i%�r��0`�8��|ԇH��lH�A��Ki�׿��R�i��1����܉���[�;7T�ӿ���P���3��(/��Z�y���ʯr�,A�F�P���`~)0���FZ9��a/��.�2��¼������1��5C���s�i��-�Db�j��'�$$�r)�5�&���N�H��e�V�V�@H��	��^�&�_���ϭ����*X�	��'���yƔ��<(U����j�,h>Y�h*�q�7t��U�����EΓ�i|Odr�R��Ţ�a�ja�R��Z|�B7��W�&����G+Fz��������C"�th�����yX��o�O	�=a|�h�x�hlW<4x�[�qo`8�6����P���S�S��7�d��i��w�1@W䅒?���f���6�� VTU�sPep�@����i+8;�k?`��M�_��@K�sV����Ⴅ������i6$�<q��)Yd��I[f[��{��7E���ߌ4��.�%K����MU�0Y��.f�KQ�]Ѧ!�D��r���p��cr���1ҳE�Glr5`��qb������ W�*����� $�� ��kb	N��Lƽ���3T�_�	�KR�&�N��Ոn�ؘA�%�z+��ot�_�A�]�������\��6���B,SO~�7��� '�6?�А9����Q1�Ob8s��l�cm}���yL�+��㷩J�
4{���%�l�'�A���V������+ӆ��[�.g����k��||���vQȼ��Kz��=�0p��l㪎�mpYw�U��<�v�WnB�y�X����_'�_�L�+���X28�ӂ=2įt��e�}K`R���Z�G}>�.+x� &S�Эb�9Ij8-�RxE��h�'�L���N&K���k`mE��З19s� �)c_[�M\N�	Q��� �v>�<}Z!_Ӽ��C��7�UɸR�B��>6�j����.1�C6�������6�Lҫ�(��TeU����R�bd�L��oA[�DR�J����f#�u-(������S�ca@�m�n��h}:�b��f4[�);�w�����K�>X�Q0t�R	�����Fݮ�8]��^10q<�3	��+u�da\�Oy3?���D�T~SS޻'�3��oQ������7�S�d�x� JRD}Vr8��������~�5��ݽf��o�M�*r
rˡ/|p�܁�&Nwbp�������T��b�6l��|q+�΄�z�*��^nm˫��H�M��N3Lɋ����Q�[++���spC2�VQ͂�|\��*��q��4Ô��d��_�S�{��h����J�:Ec~�ݕ x&�2B�u��W�f.I,�r�D�,Y���&���2��,�<4�����z���KU����-����<S \S��[n��a�Pe��Zk����:�@�Xln�e�������Tv�՗dWz���҆��#%��ˆi8S s�����V:��7b����$���;�?�Ȏ�a=�st�$W 9�
������oh�x3ZlNȏ�0|�~��� �{��f>��	[�f�r
p��l��������[4�(�Q���\�5p�q���B��k*�x���ژ�F:��KaY9�j�/s�2>ˤ�ԋ����}��?�J����N
����I��/�Z��J�x��4��)������#p���;d55a��8�@ѹ� npa�y�=i�\�\R0?�Ô���O��k\�Ȼ�{|A�A˹_���}��9��f^/=%��x.X���� ^�c�HH������:>]i�Y�	�7M5�鐅�p&S]b�0֙<��������'��<}���\[���N��Zd~��?��$��W��_�����qv~���������;�{|e��%�P�5){7�m4K����ǰ�)�%��Y�&�%�E�<ݒ+x��K�dil{�>5xʶ�b��[Ʉ��B��2�v�=�p�*�������(嬥��LKq���LV���������)QΤ���e���;���F2���>:�̍ƝF/�yp��	a����&/2�O/��孺z�]5��BM����8e� 庯�б��Y:��3�ɲ'���~��!_zh��/7���^�<3�O5t�j��1�9넧��rݭ����(�9�z�Ynl�G!�M���/*A) �v�;dI�c@��\ ����Q&��X$˴�)\�͂�A	��/�d±��Z�J�7��;�;���"o�M��#�H���NўB��z���S;E#_�"��]��*�ܝp�y��b��A��+��b�)���6DLOp�^j��܄M:4��DL��
wl	0�v�s̲zf�:��ިu�2'�'��G���f��}����r`�9�u�D��|�/!�?Ӯ�X)�eӃm��w����W��9��XR񫖉Ԉ���J�,����ٸ+���T]*M�/K�W��sQ�G�zq��Y�9|���l� "tĂn�9��,ʯ�V9�zHY�2���/��b�����8����읐֞��i!C8DN,��E�#4��wY�Zd�b��N=��!��c���$��1���,-�$�])�&m�	�*��\��9���#�f�����?��,�t�ƇޯWȬ��Z~��U�}ӧ.���V\j�y��2W�
�%WB�R�#�g�?��!��2�����8 %��G�v��q0�?N�[yZ�De9	�V�Ѵ�@D^{;�ƈ����T#�g�����Q��˾1Ic��."OD%2���B�ҍag�M�F^�U��<#�!K�[`��O���+0����Ro~�/�E��3C��o�`77'k�9/������a�����>�4>k�N)&8��+g�B*��/v���h���J��xklWjil�ҍ�W��;�z�� 2B�|c�/xfg0L>���lM"i]�㹼Nw��Y����)Хo�m��*�?5D�s�&9.���I��մ���m��;�!R*�yz��JNqb��7߲K �$q#Uq�LY�Sw�)�8igtl{ �t�:�n�����X���)�Y���I��t���E̩�r*j��NFd��1�ߍi���Òn���v���k�Q�����I
�yV��5�O��|ýr9쭒������+����¹"����t��fd&t��A�W�!���U�KU�A�����G^��B�9S��ua�4ֻ��F��R�3,�5�l0LVU���ĳ��C~��U�'q�[�+����`�1�rK��Q��Z��ˣWX�	�	�k\>_�T�|���ԛP�s�O�0�n�g3"6o�lg��vc���X[Ȇ����E�?�������˿��w����L����T(�åg��#_8������nϚt�0����3	.:��8�|�����;C�>�yb1%:�ѧ���ǭ�a1��P㨬�OA�}z���⁧a"w-�XT�1߬�AP�	t5��Ȉ���D�Y�Ta�̮sR���}�p<+��x�CK�+7��ML�3:�?.h�i�3%�Qn͒�=��R�_�^������63D�6����G1��R��i�Mp����=0�Wg�'���6�#�)���{����y�������f�&��^3s?6�}��:b��զ�0�sKGI�'d2�~f� 5/��%�;��蛍fdө�B�b�YMc���F �W[�1w�!A��^���[��{쭹�Q�$�0�N����y�K9�@l{�~�<�n�{}�")b�kQ��<�'rT&�(/����Rm��6��S�C?���C�[������gzV�H4}�ӗ�CKW=�`,$�+��"w�O&W�!E�X��"����ޱ�dea��M�,s�O�}�M'��פ3���J��3!�Aݑ@����~�ݭ��Cb�u��TJ:(f�Y���@?�bց���큦Z��|'���{�k�_��zY����Cs��E�R)��$�O��nظ?,m9�:=�.���I wV�}Rj��]��E@�b����5���R����ΛU�g�0TgI?�sj$t�P��Fʖ�l��^S4��h^f�A�Wk�\8���'�f��K��mO�w�ͨ��xK�2�6�5h�.��tt��,Yx'��+TW;�U�W�N��h�tߒ0�����Ckz�^�0�:�ȷȊ�G	�/%��#�jԅw���%��Lv�v�+�b1�� ��-w�cXE�n"��jìzw�w
,~�m���G1Mw��B{�G�T��� ;��z�d�(�=�ji�r˯�����<�s�8�Mn����_y�Hd5�}����q�X>��˷��Se��_��ާ�C�)��>!��kx��;CT����ӵ���[3-#�\8�JD�2���]�l���
���ͭ�$:a�gy�:��O�EE�"�>���a�n#w�QR����m���_�|��#��:pRf��C�����4aM>����D�;EG���2�{[�~t�A�n۩x��Eߔ�}�s��y��b7�'�p#ެ�r����=�Ȧ]C����Ւ�.K3u�W
p�6��P��W7���݃� 2G��"�K ��ppLU4U�˦��Z�٣'<�^�#o��dV�	$�D����nu�}��AxץC�@�?���(+���r����&ɞ�th���W?���u��-�<�[ �n�n�qw1R�2���?Z��S-`:��Œ��"{����lv���g�2^ݩľ�=?��_��#��l��ce�dv0�L�(̥[W�6#��aM���/�#8��u+������_齭l ׂ$��N�hSAˁ��2�$�A)#�s��P��L�W�ə����Xnrs�XO0z!uͼ/��*�8�Z�_JcfU<����n�1�+�V�Wם0�M��X sĝuN&�f��W�:%^�=�xy����׹�z���fd�^��D���3