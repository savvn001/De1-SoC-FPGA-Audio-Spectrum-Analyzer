��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	i�A�����B�h��f��	;���D��^�*{ܓ�I=I[x.>T�������������R�!i�p�%�s�����YJ���{�B�q�+ҹʵ>u�?n'��pp��)N~����t[%��v~�tN8��ؽ���fT���Ut���\������1�H�~b�􅶑ՙ/���s1K[��{r����W��=��,�b�Bʖ˗��帻�޺�	�:�9E���.���hR�o��W+ ש��A+*�2&`��_J	lxG�z�3'�k�,���{/\W��!��Ŗ9�	��u�ʀ1�r��Y��fN͓#�:���#HJ�AX����f�X�l����6@�;У��6������	R�/W�3k��!=1��"a�'WHz����9T��nkp�~��C�]��t����o	�&���h�}��3�1~V������R��%�^=�<N�c+{����1-C�|b>8 �ɬ �);�l�k��9�zӐ�\ا��[=z����ۼ���r�G{?����tBP�,�2��&%��tQ3	�
'�i*S�wJ�ֈ�s�0�3M: ��A��� ���wDg
�5��<��KҍZpS���u��TǢ
���~v����3�ޝM%^���I&?��mK�������%���|��P]��.â;9��&c���w�2[�a̫���0�ьD�~�$��|�8�35y"|^�Ξ ħ�Wf
a2^��Z"U�]��8hV���������w�&�z|bb;�<���aKG�B�v�Ja�cR��<�eV�kEo,ɓ�˴��&�`�"|���Ҟ���Z��p��
D!��ρ�oBΥ�ǙO��JϮ�V�{1>�@myUA�4#��!�n��� L�m�y�7��� �Ge&��%�L�� �ў��E/�h���ʆ�������B+�П�����54�8Ȱ��/�y��h��X��OVX�Ľ^���)�Fjj�I:�5k���n��MG��u�VP����1��̇�b�	�}D�D�r�T�K[W5?���D�� 3�� �t��Dx|I�C	�`�:zg߈o��k�(�nǵ�'f�T��f��W�29�[uq����Y��y�]�?�q��d|!X=�)CG�ȫ��.
�ŭ{_FNf�F����:h��g�1@�M׌9E�ʞw�u�,r�^�F!�^H��Q��n/�Â�G%��׍T����W�70�L*�G��(h���j��7젨�Dh�q��*{Pw`:2�n	?2��.0���9� .$��;3i
�������x�= �/DQ
�/r�{^�n�<7��F�LF�E���3��2�w��kB)��3WS�p��ظv���t�C�6j~EC�1|}4�_����,�ٲ��B�au�:�����<��1K��5�^97`d�͌�^ɸo	���._�,������ѿm�p����n���߼i��ajz]�?A��Zi��c�Z'֔AfN��!�+���D��9�рv-i) �&(�X9+�>;�B�K�O�/p�L	i0�F��}�K\�P���$Z6���o}�l�Å����2�R&|��ݠ��4mc�a�P�v��������U2�������v(7�q�^��n@-{�>~���q@���غ�!�TC��+�!��L��}����(��h ���m��4��+$}G!����V>:%�|�ca�&S��Bs��㝿���3��:��=N�sbr`<��e�j�����z���(Z��~�x�2 ���N�kIVʀ*��rǵ҉�3��愂�P��gӃ|���B/�a@��Y��&}JjIbHe�6��:A��|SDD��K����}*�+k�`T:y��Vz�lļZ�\���Ԣ��@�}�E}�g^s�︎kM�{ތ�:}�.�#ه���>ש�נ�|vs�~G�y�:�7cJI�O�;�MH��.�ݧ����x���J�v�74_L�$����dK�%spt�����*���>�����r6�]��\I~XB��ʗRq�2�Ҽ���4��.�{������;�'�W�%=QuYF��?П42.����7�֧�Gtw��f�qױ��]����RE+�V{�D��џ�+1]zuy��ѐ��Y3"��?�Й{}��Kk�[I��O������TZ���ۿb�?�ACv�=���*�<���]����`��vȐ�6欇ۘ5�kB��3��J��u1�����4o���
A���+��8�n�ֹ|�Mlz���k���W���9V#pR���O�Уj'�}q�������T��P�P]]�>0�O�bT
�֘h���������xսn�����O@���*D�/�����R)Y���L6P@H18}I+ꫪim\�Ƕ�$
)^�H��_?O���'��:������u��ٛ���Ӈ��f_��ˍ�'@3��f�w�FS�0�A0��җ��l��@D�+��S	�(�p�%�}޿Y�i���(jP��xW��&�P���~���m�]
����N��CV���C\ 0ְ�>]��ӎ1[�� w�
e�])�E۴t+шS��+��>�Y�zՆ<-D8��1�JUJ��D�Y�<`<5���s���P8����#��<%}�%!xxN@�'�^Axl����2d�"�/�cml�hI�.{^�D��Ɍ�ǀA�f9~����^��k��{(�I��r(��j|��e#h|�W�Lo�R�}�HJj9������CՊvp�H��k�
g�c%��'ڸA��-LD�����1�$�%*'�#�-�����,�ۍ����A��B�f����+!��7����Vp�vUH�vt�\�=��\��*�*u�W�Ӟ��
�C�i�ߦRF��0 '���r���l�Һ<�܃s��ι���!7�6�k���5�nVHszoIB�����щ�FL,0�><�����U�4G�m��Kr�n^ e{�e��#�����#�iYHE�������m" Wd�U�|8�����+�����m_ �\~��LHa��QL�4ǥQ�Y��	�{M�he*���Р��g"�;�2[0���˱�C�e�%-��J�;<ן���g�L�n���J�~[\��p`�g���E��5B�j�Ty	C[Ғ��e��B : ���pw�g��2:�K��8�I'}lm��8�w~�ɭ.H0��ͻ��N[ޡy\�f����0kK�5xj/�3m�#���<���8|�Z���u�=]����8��Y�m��_�؛JE�'�����һ2���:0]ސS%�/��-9`���`����p�p���]/-��z�N�����~b��b�-�6�a��{�������C��P���7�Y��Ͱ�n{`9��Z���	��dg(=F�f�pS@�q��"ԂI����}�����I?3�Glu;[�o���k�i?�<�,+�1�6z%!NB�b�^"Թ~�~�I�F�?�Q/�Xwa�ؽN*����3��-As��n2�?c��.�ē��c���-t������K��8��=<W*>�>Is���Jbo���_b�/Dq�F~��o��l�������u$�35���P��2Ք���[�Gٍؖ��4�׍� �Ԋ��5#�� oaB���Ν�J0M��<��AE�O����ގ�����c��(�?1-�M3���̷�!7�Q��h����@��Z�댙w�����,$�h����3Q̀��Ǻ
�mÞ��]�u��S��yM���`C`i@�"(z�6<-=r�/H�c�=Ĳ�?e�^&�聣*�Ȗ�ֿq���6��=#��	�n�!e�%�`q��c3:�c��l��;�y��g-y�����%s��C3���ø�LРd�G� c���ˠ_ym1���ܜ|^��d��r��i�#+�b3� 1�@`a�3܌{�Zfo��_$%���_�/�R��N��W�f9g_�������^���Nt�I�+j�`�����c.`nݫ��jʟX�4�Q����
����e8�DC���h�oh�!g��.�S.�Ü�y������W���,>�<"i~����}��<I����_�+��-���7:�^N�4��&��C�3�|�JE$e�?A�I�{c�S���c{0ZC�x���Z������/�2�#}���X�b�p��<Ah�TBA��<���6<ƊDb�2n�w��Y��wM�ŋ�"ȴ��&:��xaA�?��˭qA9
�q[��B��7�.6bV�vmn�Z�\ո�s���}�h�]J�y�F�u}����;t������f�e��3i;8m�UcYXJ�F~�ˣ�i�����q�39c�艧d���p�Ҿ[�X�Ȟm�bC�������e����"�(�z�,lM�5�\;�aX�]�\�J��m��7��j�4T�Hq�=)M�}������P,���F��^d�8����*�śD��W�k���jf��u�/���TȜ
��M�$h56��"��YhkD�V���{��3y�f?�QA���Z�����k���� �+ۿT��CF#�P>-��Aҏ���A�N.���Ŀ)�Mּ��b>�Y�h#�]�l����D�~����U�M�����yje*y�@��B����=�'f��pǇ"�"��zGG ���$��3�)���LX���Rܔ���D�l0��d]όu��ek����Ֆw0ՙ���nM��:kO���16`d�g|#�����M�,����l���kå�5�j����vzԴR�dQUoL��o\Y������G����yY-��m��0�qԴ](nmO�<��2G��Ѡ�b�m��L���<���Z�d�j�<��鋚CXI�"����.Ȏ��� ����C�����"���E�[1�rb�d�b�]Z5/�"�DLM�bbL��N��]��W���θ�et�e�Q�P�	���r�x}g(�m����RCb�@�Y��m�&���@?,V.	"�k5�ϭ�{wžh�����Y����n�m+���Z���9��J���~��$��HBI¶:�b��A��M9����̓J�2�v���<����3rg�u)z�6�S�Ӕ�*?6�������ߪR��ؔ6�jU�x�k�����Fw��RR��qޖc�)�"P��Np�"�r>��X2�֗��1�4Jyn
v+����k���G�:�ə灩
TC3���RILc��z�Ɓ�	�5�0x��}��{�w:�5�dL1&Fo�6�o�!]<�!���C�8�G՝�O�;'��Н�a�|>m	D��=9�hݴR޹t¾s�g�8�rz0�b���d�XX�b�E��2 iNa#���&��	}�p�2��n��\���nM�'��tHA����8H7�Oa������wS���X����7Y�=!���ۃ���*�Ǿ����q�_u#u�.�qgǕ��%�'���� ���i<�Y{A$�C*��Rs�N�d�`CS�*��}��|�<�_>$�C���\f��dk��'���=LP$�*��)���6מ;o ���	eo�U�{�QL���>�2�1RoVǴ�'3��Uމ�g�-i�P��O!&QG����N���8���z~�]����֧��N�x�>�9i e��L��^b�H4����CO3PL���B$n�����odg��D���e�F"3�"g�NS�v��\�>8�iDK�xHY��,O��]�Ms�{��2�«M��1�ps2�s����ɶ[鉠��z��uaQR�B�Zzj{���pyX����U�h��Eu�J������l��������v����jp�o$#����P���ʪ���v@
,*0�߳�S�,��S/��P�	_��ڔf#��;}���6@k{�T�^F �,}O?+rT�n_%��];èߎob9������
���/:d��I��A(V�� V�ʑܞ����\o��	r
X��R o�U#uR#	?`��]�٢XH�q�zM
�ֺx�B��!=�V���?df�~M=\�J�_W�6�N'��}�~n^�G����n�V��X�ͦ���W����*m�6�F���O��Y���*l_cΏ,?=/��LLå�
�1��)�o��l�w_�2+��9��GꭅR�q|��9��I�R���a�`@� ^2�b>�( ���U&=����f0�V�Ps��<A�rԵu��  '�QD��d�� N�Mw 8��js�!����"Ny�*�[��? �F��r�ސ2Xk��!y6ˠo�V���T�HÎ1�F�{Yܸ{_ �� ]�H! ���:�"�����g�o�j!��n����K�J���3�i�d�/|�5�*(�=¨��L:��͢cԽiA�!�sJTA��,�ђ�E��M�ڑ�rh�}E�;�g'���'��ĕ��3�mf4��E�~Uk��eSԚGϤ09�=��o��:�'��Je�c�c�!�6������PV���y�5����u#-���?_S /�QMs'd÷O�y�|�G�7tB�.��y���΂�6�r�cSz�n�����Qgt9�C{J�'KOI#2X� �]�af#���Fs��@D�2ҫ��+�T�,	g?�G�c�)���bČޅ*xӂV������H�l�.X�@��3��}r�wL.�ô)�(�m��A��6M��)\���)n�����>琓f���^xD�������-��Bhm�h���"j��O������+�������0(���c�}k�{"����,	���O���|���*<�@��T�
Y�%�iX��1��/;�I8d>�0oC�\م����gKΘT������.�C�H�W�Z-Ϛ�+��1,��>�^�σr�9aK^�Y�Ir��W���~Ե��,g(�SK�y(*<�u.�����Aݎ�j��lb�J�5�YJ�
���5ϣ�uah�����N�i9��@���K���9�P��m�!~A�[+��W��+��N�R%�+@U�h�?��N�r��qJcfo����ǜL|�F�_�2M�G�7�t�V!�V�� >����"Eä/�+)Ȯ��ݔ��,��\Q����WT}�.K�"�[H��=&$[`�p�i�~���^
��P�i�92�����[U#����yL4�����[�����<��a�lB����b�V��<�{hdE��d3͉+
�'��B� ���7������+UB�`AUP¤u��i:�� j��D���->N_)��>Z��=/�6Z�3���e�����5(!�'6bZ�X�4	Яű�:2�'u���]��
d�"�|��SR���荤��ɕ��ӱ� M��-{���$8I�$��!A<CQ�a��,6��t���Iu���\8�?UWֱ!VJ��=n�ӛ�J�ǁ�ty��/�����|�5y�\l�0P�bk`���k�������9;}� ����S��o.��W���&(��%F�������!_%�kt�R�
���CG��?�(h	S\��v���)�]�2�M��C:a�������a�b�')��8I����`�b\meqR)F�'��.�6W���HH�n�@���{?օt���6��7�b|)j=s�X������~,H�;H()��WsR�~�F�8(o�Y[ޫ����vV�s'ۗ�.%��=����`����}/3��_y:^G*&z:FQm�	�NҺu�r�+�Q���(&v�Y~{`��y���WK%�Įev8*���M�D�