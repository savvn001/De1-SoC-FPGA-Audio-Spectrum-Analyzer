-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Jb52CWbKyzmyZcCEkLszZ8lWumfvvB5LE4Q3Y3hLAJyWM0qtFU9hc5woxIzUsGr5DZY2wNlRX6x6
JOTd3w52EL18X8dipvRTlfDhzLQbFqIeftHbVCj9rqaGR53PElAGoRpwnNF06Lxbhjevuws7uJ2Q
j9VY4WK1tveiC9/kOFa+/IyXFKWBxmt8MF8DkyNHjpj25a+JoigHeVLKWCC8nVZVaTJYKbVfJNVc
XZgpVvqe4klBlhF/57seWi0NSd1pqZWSAEBibpf6f9Vb1qduqjDakCXOAlyC+5dMDWHLejzQgXDK
zlGA9ghbHtn8O+eJ9Zu57ie9SSRIj3UYVnQr+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35728)
`protect data_block
Nzu8Fb7GGl/eZ4vp4HKQKQymfMCdp/ZD66aiAEZw/kdrlwjrlCGHWE+JhNck5mApU9hpyYDafsKo
OT/Vb6o1NsyP/jZ7iYEi1mIZfa1wB5FaQMqLJl+GbI7AL5JlR3F+sBm0oBRkPWUHhVhhU5YF/bRT
e4yDyOut8chnP4FUlC5sF48itMS4ODK6Bl2vsrkh7k0JkW9hy5qRHVB/VAPxp2ypXkKJUcAQMrud
eJV079mWY7oGiH2I/tXTx+19jW7Pb022BDNb+DAbjk1C6xYjJgU+5FkZBj9xtGvVku9MURWdYkM0
5/8iiizqCszKAWx8d1Hh356F9C6fqDKe3k78fS9Ca2/Qh2s6LnMZlka0mgV//jxIb0IvF7LZFyax
CVmpBW38LV24vSTfXQ0DOTHmOGH1HDRlZs0Nx2DCbqn0GQBmyK66BfIOMCck8V1QbgdQ8Bm1uXYx
XMaA6wgBNThT+KWUhXy5fqLnhC031VsVGJdSdyRe/aDDO7lPJDx+vQfz7dZe+iqn6g3JIqsGsaJs
8I/55n2PHEY544zxlrlzbTnl6gSoCwZ0xhn3ZkpUB4QiJgkPU+5YaPA2XAozL/JwmKCJLhB7fekm
Bo97kyfSPRAPvW5u7nR4X4nr58s2AE/RsMLNMkUAdSf+uL4aBTyXLtVtXuOG9qVOirRV1R/wvQcp
VPi1ItM/j87C7jaj4qdIJfp0b58DqqTcSuXB1pqOXTy4djK4apP7NK7YywS8EAXucDJdgbeBvoBb
076v7ZVRntbVQpQv+lVFqQ76xR7PzZutNgfWocEC5Hh5MIPVYDG7KPrhipua5R/0Y1qL/m6Q21hw
gDgqE9legT0yLEBXy+pNNp+KFnGT0hregywZdglNE5TaWNN4bb5syrd49HUjt9jqUhhiaTUqIxcc
a3eF0fWzZCho30s/xMa/BYrfCu9Qs4q04O6iH0JU99xRiGqQcuZaNgcA3z2KLq9rRAJgIQPgpWDT
i1RgGrPWg5d7v3SvN4M/rmmiSCFvqPRJF3AWS6v9J+bcMGoWptWe3wJwEcN1NjN4dRQTuK8q8MaS
v6dammw+LCvBVcjpLHq6oaOLGEHnaV8sP/Fjv+dTanBFktOTmm/8DxvXG3Nyxnekm6CyC4aiCv1L
+X4ruh0BqYAyuhIfKJ3dSJaSm+XjzIHiLf26ZDotJg45x/iKy7YiwnoBfxl/pIhcrX9h1QgEACzt
4eP1A5wxw87MwbX48rEUX62I2YiJgjVNabxl0chF1trQBjZe01cY2eBGLH0aIh9wVhrJjFu0fe20
DepHTW5n5p05ZOh6U/U/LAusBNInbLLrGcybPB58bz1EvfplMQWZxO+Mynyx8gTc2H8oNRH2/+F5
KJ3e2SEdUNoASNB0Il8dHhS+4Be/84IyS1N+2sBI/9oqZQ4GAM2EPTeRUwYC2CjQJzG4dsuEjQbW
4t1bFq618xtTu1H8nV3pQv3t9hR49+vBuaH25erBm0DScZgZdih+JsYqM6Hb/ACi+0LfgLGIVuut
m0I7pq5gFnWn7MnEBDPeCgSaoCZ7YgSH3OfyE5Ucw/m28MW62FB5PugLao7e7I9FqNX4XEtRkyaz
7/jqX5Eogo1z+0kF7Cki6F0qsyH2t27XvdtkgJQtODLTPKHNh71IjIQ3lMGB0QftJR0YPQjmYkY9
mH++1SYWhmgOFRaxSF+w8xhXwvZWggHX+eKNB3jvfVHhoPbbdcRHanJR/RYvHQadaZwXmhqaYEYt
w9v/wrz3lixY+ftmIPW8ByK/5g/aa7ypdAEn7e8YiVf/yes7TNwBqdqIE572S5NZchRt9W3QeaIr
0zxEj+oFoZMWDESxjWRSVPu5AZwT4EW9qNMQu9MGiV8XUic9S8SFfDgb6BWcjtqKJ4S0XxneAzty
QK+VDep0iR7iKZk13hzCE+pjUG7bYJzxB7IkVvOFtQ//LpRrPlxCP6uweIwnm7p7iXUxHj+H70tO
FbIPF0QGbYfe7Ksge2eREs+ukOs1xFZt0NviBrHJEgC07ZtAOtrlcEdvE2d6unFPkK6Khq/lPamS
lk0VuWH99U1bCQqvFF23wxm8oWYChJ+z1D8oMGdZUZnqqdMBqyHwje/YJDChNPc6GkULPuDZ6TR4
YYXIWrRsTY98UTy2odL/8d2AlDwAS5sKXaIYWkDGH2CVpXppReac1CNTcl7RntshC2xcEjA6cvsr
uyHUG/LGi3R1/PQYmTT2YX0dkg99H8PfAHNtcXXKaV4FcyW8vYYR2OxlMWrK8HsWzGN7TVtSqFRn
WnNznOuUFTxvuCI5lfFzSytHZEbs1cpqBowSRy/RBa5o+ZcRlaFOdotpQAYwf/ex3qvrQBOvCbEq
/hCYvJ6pfBJ6Zc57n/jNOR/dKezWNTOeYxAE/M/s1Zr572cNTXEgvGUZUR9bbKJGn2b1g8MYJpds
XnQwwNzwSNiiqVTJsB31yoBrUHUydMYhXHW2gCdu6uwbjrz1pXRHyq9cBih7ulES43YA6yWLqins
bPN5XrQY5KWefl+v0NdIljSXQ/tNjeEBamubtb20im+tIe8PfpiSVP9wv5ZRnO1eRVXq2RpmgOz6
fNy1Bx8zhqzSM9/Jnl1Pto7vCf/IPlmCmmyg0V1GG8jPJ07IJbZd8hLDf96u2s5+DYxb3Tpzo8UT
w0X/SC3uOMWbY3bY6M4CxWprYSGwfUenkoEWhByp6I+U5K230p1nhayuX+lBOzG6CfTi/2ouNcFk
vnc0fk6v7hVUe0dxUhPbgQOpB8Dd10590vWvFzY9I0vZnyQHk/QOGyUQ6m2hWQmu4Chc0naQnYgH
2u2UXIySAm9Z/B2rhj6aVTHxZBrTB+GDLlpsii2yRLvJw+1yIt2L6TIjBrQ3d761o9En+jSOIsU9
iYSYuwsRANCkZXqF6HhIq2ExaPGUu9SCnSXUfyfTNnKaHiMKXezOxQKg5tCwSTIhRE/7F199HGro
Xj8tHSKpEXkyzNFbAGvFOlXxgonaeZWqASPA/NyVL1/O9Ax2IiLm+ImxFJ9JkvYnHIC+fErUgc1s
KFbTftYVOb9xcZBAUJ9UeRVLuxa7d61v6c9vwCuh6PNTdOY5OKUoms/A75g1ZyUpyLuUFOqfOfwR
MZ85hDjYeEKWGuqzcDDNI3RWweNm+9GU0s3iideBS9d/I97PXk6bSHACXA6em5DHy31INLI4lUiB
JRcHW+jbvHc827TJzwymiQF/MFfg/5HP4lnLi02RlIjKBDi+eZlk00wcdguAFwbUIV2Dt5ojrShL
+c/rI2fognoDS3SQ+WNCsmTEkpWdgi/0LJ3iY2XyByIRSMZu4+6Zd/YponmhQzxVFCDHcpaU/AHu
vDdfS0W1eRAhdlwgNe4CHLGzd9je+pt6shAUHgEb1EEvmqRhNi1chsuDtVpIh75sHIqvXjXmo4Pp
rfeJk1V82qP+myVJjfHwD6NGEwY9oKwv/rZCAfwK+XgwHhDLlanuDUYMq1i+x0ohwgUNwhGElkeJ
jQolryuYUmTgexi7XSPSdsNasD6XhqZy2nbhKzoDhKrhbgtLBX1pSH8l/TRx18dbHBmgQ6VEzGBk
rw5nd0RR4ClIrcE5TTgLB/XtyaIuH4zxnTR9Ei9BwwyniKkk+IaVQ392wxaw660RmQj8XS3IY+/9
FYgqwWFe5HJKTaOHZzvOQD/qcS+SfsKzz/ROO9o/7ra2T1TdOWIDM7S40LmwIa4OjQRPyjwaognF
8/SQrTjQ/r4tOGqd0dCiiA74451vPBZroAFR0oJBJKxbSlPiLahS4pmyBEnRXJMRtePXLRXUso0x
4nuAFpjbCM5cUY3oPNYlgz4QBs2iVFFoP87btwlgaq5vyV04bS2t+CvBL4yuXcg7OQpK1gb0ssNp
F4vrOTyolSKNeANsh37qxCwpNfZJ4UYlbhpR+n4EulBiW3YA7dBzzZ0WZnDuw/ifLNJOrcvEZUlp
mOOUX+Heag/yryiHSYtRq+JLPxF9jB6zMMOhF7krs7yr3OjT4j9LP9l68eA03wRgJY64yokpekRX
VoqB5CKk2rIo2UPu7e78AsA3C0CHUFmQr6Nq2jWRTF/NBf0KjfZTV0pb3/qbZ67KsTr0aQkrx4dB
Sfq/axOrTBvFtqm46lEI1HdBf0uyGafIJ/BnCAdKSHcjTVQFZkvBYkK8SCyDDAvkRjC9FX9zMRlE
JABOoW7j87L+uXAmkoqCjJCZ2hj3x5hJfpfLN+IVS5gLisSbxakzqGj8Vig5hkyR8047wnSxNpqU
H3H0W82hEZUkxHHJ/2LtgJ4L/R11nJiJkV7sAR6s9wyxJbl7pkT5Pp/Q0eRtYIxtVaSRLmwOuBiN
akPCDOMk6V+pVelZQIq/Q0QzSD3U2788qBCGDKPcDq5/4Fl671qD8E0iYnHba/8zF1r4GUrRZJaS
r9rK4qFGp4Lp8JRJEGUUoFJXisFLhWD8cEY+AykvpU6yyhTfKgfsTwSP7gSxAuvMJ5vtIwFLqBvP
qQ3PkVldTeHnct/rK4QWp1pGa446cKLhjhejFwJoPR4CfP+ctW1z4faGRDY1YhRvmHNnykj/TTVi
6UiTUEz0OIoO70k2w283qsgD2l2VuvhIHSq/lX06+RL8y0jjctMwahv/oRXd0PXnQu9NsytVFbyO
EovmM9wMRCAy2DJLk2kj9vHztiKE+zzC6o8X1Bk5lRULA+eo6mwazPwmAkpQFq3zxLnGXjVz4Wtl
Yxk+GrBiBrBGuWwuDEURJrPuiaa5SrsESsYsLUYzyMOnXKHd+DtSRrBhz82iGZ6XPEZvY58vyw2n
xitnhW6KuH+S9PUDUIdBNVRWgeqAEtGS4lpdkgWa++F4o0WkWFEG9QSTmGtLjQXlJSXtXAO49dqx
/LFu3ZatCIqbAMjrffNx94NlExXWR7K544AGp8v+R9BFFwVAQB/PhX8niB6jtF96N0vbPKf/6yAS
v9GrZimZPfq6AT0PIKds+PQRkswTmXoF8AimSfk1ytxlD231ULP6otZ9UAJGTVbuZl0Ni84wZZ1M
QU5oF2t9sf36COz9vU4LtMHCCin8pSgLLs/wvxS1cGlXZACLQVZnZyjq3nrkKGheiIYC4XrMcgc0
wCsZ54igSAtSkB1XC2rqfpyvGJwSKqKDEGQHwNlgUVTe/pEvhmh31+yUqMWknd0Wsn6QSOHLKLvJ
IF3spo1E8L2DVWCP86wFIihh5Gc+cCSD/OYed2u821Z+8jp6Nk5R01lw+CZuaJki3fbq8UzgFDyT
A9Du6cnRDSSJHW9EZqYFStR5uX4NHIzJ1fEbG3MlL8emafUjMassJMur1NqrnC2nDU47sFNF8N1A
yTlu2etK+cEDkanMpo+iF7KGAuhsXypbrHUPZmljD42NcKLyBB2qqNuH+7KGXRhRqIrK1ZSq6VM1
wcUg4eyWsOdmsIZSC+hHobKFJDpTvHSIk3Y+KGszJv3Fzjd5QVR+X/aZWIV2CnOLufSMptNTTeIo
Bf1USmUEydCJvY4TEEU+W+H79XJ7srSVsZxWjQQjYl5+Q8PyXC/MrukBHGBF3BSj1WcrdTbfM03s
9ixRmAYTF1L+YAs8k7wV0c3OzmHB984PGzf8IY5ffQGOyC+3Ee1soU5/oTTri2CInBt5WvDrI6kK
QnZqpKnjoF1XIvzAV9F63i6FjKFncuduZFn7bRntqOgQkFnMbi/GEKgtMzxLAm0IERJcGiI9QI4f
EN/7xOpFWNnUmSnLhneBj+jqM4BcrZxlxsNpWOJ+8iWXnWF/ImiYjyCxSrbilDypzIMnp4GsOxDr
+9j2cN0P5V3QqNlJUQUWZWKzxOwzc/fPp3bYGnT4KK8Z2aMZuiMjVAnO3XgB9JnrKVVVjOS1YQWu
iEkWvtG6XN/rzOn7mDIDe1aLD/bwLqiNTqwWRu4Gi7ObMyQuzhMZyRiu17u5poI5Vq0jRUw1XmBC
3FJ4DnWYX9M27UkTQxQECdPqLzOM0nOjBeHSQCFeIVxF1anwnTKqYe+I06WSpOV/aN69/fvxb2AZ
zwl5nfXG74HFK0Mne1QxCytkU1Nt3js0wJOLACIsvrGa/jz220Jva1VzaAWC6yG6+JBt0PUm8JNQ
XqegvQC0fOpMC7J4zVQwtHIQf8KE2U3YFxU4CQVIv9kTc4H//c3bQqGjB7FRpNg8uqeyazeNcmzL
k/wFXgaqlt7BW07zh6ImSlXp7EtgiBcXyon9qXpq3EJ7edu0fpgrfvV3o65AV9l7UcyyEwoBgo1M
d/RCa4CSL8rRpxTwMFPwJ3eNZxcePzwp92aDnaxSeUI+JHYWSYtV2o9eieEHTPwLx6/ecMLh2Glt
MKBhzmS3ICrhJ+Kw9ebmZZJBj+ZPhB7O7jAjIYJWJZ8YK7BW9ZSeADXIy+6BgJ3QcmtUFf6jGMXu
scbFoTTnqbUERKLv4uMXiarhvNRKLfV4AXdclqnQ0PiP1PrBB1yVr/ClMFfvk5BkPhunW42jv7kN
fq5DEjPh0QchEUZ01x/o0aa0jawUsHlhkgtuYsQkqtLaN89sZPHsqiQ7lJxBKb+WJXartN/kZKjJ
MYBwZ6w8IaUUNzXCZp+h2yh5Pdl30vzaPxQKKMFoIR4rCWdrs3uFgb1BLfVpFgpfbbgk5px2VvDK
omF8m0QlpTYeh3lEfYLJ0bWWLIZGf6JV3ycpgacuzSj5g0PscvS9xUvUKPVJ9L6gWeDCcjr57U1Q
bCSWduv5kyw10Na/OhIHLMhWN6pNP6KQhNrW8iLtvx5BcFPnScD2UNKzqgk23wL9dLMu41CTa/Tl
T/hJochXzB2FVa5cGm0QzMn3cyr6s6t/Nb24+dS0M0v32MyklvCVEGdFuF7TyKOkSelH+miXCAWM
uozK3T0fqwUasOQuYFWEnTBN39ssmA3WwRinMcDX8g8hp6tV/ccdfHWCwToTwa/FBkrnajf5p7AY
RIWz6nwkG+Okc1q38ovt+NaKNfaGC0rFXMwnvZbl40JTFEhM0iADVWjlg9sk5LBO5APOD2VuwR73
vvkoQuSumQAY7UmWgdcd3MLN23QVGt9EZ122B5M1dx8hpXRGl4QwwlS6HzrWVe1kPP3jcFJMK3wI
BKVK4U5w3IA9HiAHN9yG1T3w17GH3JP2xFh8mbkOCIqsGc2YpWlBSfo3c2HL9saYEVwwgfVqTa3u
8c9ZmoVXsaFSTWsR68TXhGmgfvRVX+6glBUqPeCGp0M/bb8wNR4m5XFK6S9TiV30RWworMrTQNzK
Wtq4c/X/73I0kAZUMoIQvd6oxtFy4xAy45Bktu7VMMGNBMI4nAeg2bkxrtsFHFLFBB2KIo9FE39S
loStMqmB+oiOAcYlHHdMmPS/Nv7Wc8Sm2VUXTayzqEKQGw/3lUQksQns9N6WGr6+CHQlJ3xF0dT1
3SSNIMzauA3ZEYhW5/75wfe3lAePMXKvBWkMx5EPGgylO270BVVMX8nJF+9vr53iBHVJMBrePsqM
WXWMBKHnT6KF7MZWO3cFuosQQn1PIJsqj6OSe8r2DT03Kn6vyHRafnRTpT3lcxPNdmu+YUcMLYdA
LGvwrolGVKhS6lzrmIAVTkQ7e5N2/ShXTJpiyR/LN1MVTYOwrQ0qhjqAxz3J9v4zD4iecLA85Ukc
gV4G6fPRplqy8G3qj+Dn9QgUu90r+yYAQw9M8g7u4LHvj9NtAX/NQctPhWJOqrv0DMPWGn1BJxrV
GTmcMpXcjEfxoWBxeeaZ9d3x+u3ZHWUY4FTFjFx3J2GalHzAUU+RUAwMEdLP0+nmxBltQ1VgABK1
J0YWJkge52/BCBGlDAl/9JBkbysWHz1Y3x8jyB4A8ARQhMeXgZetJABHKM0gafyBC4x8JaTghosK
EcCdp01yZsmsJkFdWCE5mDx1sTKz7hlEAXVFXWV6bw7oHemNzlf5bbWrJ25FxQ0c4S3EVH3HB/Lb
NsnNcBzxUVpybIQVxQMsk5NuM7fMI9vjtpuFKW+doVoOHdb/eT89q5y/42i6j1HNiH32OaeWYS8q
McZiZX+5WxlbRpiksbx8mfa802tmto1us3TXp9ZGEyRSpL5LlhOvy9cfHH3clNBSFZi9a3/GHtKf
2viKVgiSoJXWU0huOl61Vc7zGVK4Ne0sqquN9HLtWkRRP10iS5SvU2t6w32mIeHkQAW/T7mRB3iN
kylb+HT6wR9AIF1cRKmfqgCSd5ndqeMn9P84rPpwGZyfFyXhUleupZwJGIaewm5vS3Yh/bZr/wGG
LBOYL3wrc7W0Odl6PpKVtOf8rhH1yDCCBPBCGseI4yYfcZPxK/M9YefcIi8vEzS6S1FiGz47veH5
Qy3P6V/ELGJY1XqQoQY5hMDt/jx3s8m+He6st6eOYve2xgLRddC3XtPBLVxevVAh4JKUDn8zmb0C
lkplaNVzGjyzwk8p63KJmhEPLtQGN8CGPipUnsoBZ5/iSTzak690r6oLnOQ/KhsEZUQ9YgIs7vrC
E0hj6gaFDJmSv0NwbyVE1XabsMMg254Agz6hAruG/BHJ5zXFhAEn/0JOWVqKVJTO8zITNb3q0kkO
zGcKWihnNUuuqTLcS4uX3spFczeV2UhptklUw+xIN6XucME14+Ak8ul3PTbc6BAyrJBFgODSRwo9
BHsjLWiTfTg8J3HkRQ7UAAXpE8pcFHXvxkc0eG+LlnUI4rKKvmlpj3Z/5LSALkESUO8TlbGbhqF0
SKipsgKmnvoHoMUCrvCwnVQeajDOSLqMh/LnlDJd7I2zXZ3Pfs2WPlOFLEth7iRr21npJTa1m72X
Q9Q+fnmSF64Qa77V+kztUMSkUR3MmNEAJNtv5M6GVYPwMly6nCWy9EaNLfg+Que4LakKo7I9WDTX
CAxrTSHn851Xw8ASTRDfxX6mUsd1ma8da8Vw1pl3F77uJLHpZLF384d5P2fJsifTkJQ0Wul9q/xt
Mm15dDs1mS9QbCG43NMimfTdzNwxMRKr03T9XfvckwjHgK34pccjdsWyGCQyYNMM1NsaHeBUL+AB
M/pdyND8ZsKptRmbc9Ama+M54TSVgX/+yYmzuqMIFfaPWecmOPkoaklkhRkVzkqcOgjZvQ1NOweM
50G/9H5JNCaKUuzEoIUH+Ev0ICRhlzXs2qjzwPNOYYmE0CGEZKhbtkAOZH5t42gleZG2sB6/y+A1
QXQont7F9HsZMsngcBgOkW1SM3bPY+LuThs3E6w2JVFtpQDdktRV4Aka+fPEsCdCUxfy+HVR3+mD
aoysZFYW/TOgwwH/9gUT8zQheuLIdLeMikrND++rH0lay59XEFX+Wk5UohJ/q0pw+Z65irmeyn7l
ZArwWJz1cacl24/HR744luASfslNARao8LqRSeMUVBMLjTym9+6rwSNQads3cxz9CebUFDVy+CrW
M5EYkcXZdhSEFsnnNPpoSqj/lymMNLnPF/Pub3UwQ1tcQxG8ioabiUuER6rmZjSYog5sFzumpksr
Kg0Ru2UVs329V34y6fAqFLiF0AHpNt+K2y09p5w08Je7XH3X/Ewo2ajNZK7fuARI61pKrSaCinqN
yAW4ujAitIwer/2lNgkVNWZrVSQez53+VRFPMdI0IBfNBjNY++5Upg0JhLLU0DZ3JURQmk9LmtNx
wGOSycLqf4j396A+NtvX+neYYuOyjR3qnlyuV40EsqZ30L1j2tv9nxKJS2o1bRyh3zqgWcoy1XVA
08aEiZ+FV0CdgVQ0rAEMWaPE/UjiNoDdXp7N6Mz8a5Jm+IHQQIsMbOXMe7GsYI3doUZ7gxPAV5W4
SzU0uE0D7YkWsKukKW4P3X91HdBBUtETPYH00u+tcP9W8mwkcB30R1zq8xjiIiZoJEPtNd/jbpDN
y/sJUrxXlD224bv6jC3C6h+o2zgYzHALhyRh5z9n7lggLmTDJ8m2WQnZ9qKTDUSleKwn0kef+INf
O6hzr04er//SaL3vtmzMlNSLyzWc8TmsMCzwxZtim+TwKOtMe4l+TUhrt+ik4LH570ErM5kvzg7f
j0NCCcuxRJnWUuOLCZB9L3nm9BhLRl/1GTcMtFEelFZ1c/vKJsPCUKaIkilloRxU9yrPtFEhR5zk
8IBZze5wW4NtfjC5/TQcXiFZPThbAJip/DRvZ1hzASIqrQjECljM8lLr6kgGeg+2CFHE3Tj0Vbv5
8sg4mHxHHZ6RC3nEuYty2QLvLj1CeqULXup1ZW02BQd9aeWmWk8cXqXo3Fdbroj7myvS83nV7+5o
UHjFv1957710P7gFKT8gSHkSPXcFsAD2QWLeBTsteKjfS4y3YPswFZ7s+1bazrMCdetFOG37zmYM
m+VNoeOW7dliSvt2iDLZvREqgkDRi2hCeg4opjycxV5PoxrmZVCNaLO2aCZus8JO3FfrkE6vv9/t
J4KcQ7sfg/fMK3F/GWFHMkpzWMTpXnTaXS5I1fDeXcJRYRzLLfDNfnQUaI7CRF7aguSH6LxG5U/s
YAlhthZu26caO+th4Fj7QcIs8geaTrmNMBC5oTEIdisL17FJ/0zQ+fAJTgy5HDeUtTSfytcbxuQW
j+j298w3HPcXT5Y2JtEWTDdInW72qjnhv8udq+/Xo571jUmAEr28y1jCefeoFt+K4BRuAryX454G
kHgEgIXXUzOGO2MbGPggtSluAN8fJjNrddxiWMt1nUFqQEk2SD+RVLLLK23ELAcBYKhsZvbrUqMW
L/al6CA1dioRt5dhqWx2Aha7yPOUNol+qLnPEIklyWyw+5sbfYVtSeWRPwbGpfBIEaQIkK44LHmM
g8Q+8pdxUKdVMnwsGi/t9ryJvSiD5gtkZMcy9h87cUz1wjy2ZhRwVMMkbxNDhJjUWiF1iWcH89bC
tVM0JtCf2EbiToXgKPl2RPrliU1QysOxu0MxLtAXL8j4SXJ2TYifFwTubMiCxx+UYD24sPyveNqh
F1g11lnAXgkN++GIRwLvJJEeEtvdVMstM5IP5dj/xY1KybbYRJykpB6GCML8Aocvz4TXuNgZ8a5S
FPc5PxTNdlMnXBtG55AzcPh0/d04IaQHGsyTFDo8zOIL0vw2Vdtfq9Uq5TvJlAwZqZKVWlZk8Eh9
3WetTI4yiitpbm366OK461lZS5De5m1hKyjPBT1x6l495FoAqGEy9tgfHwahJKox1pUz59ycxra/
1RdITBqzg68EqJPrDivExr+UjZ7df/MCtBLqecwmaKmicUUfFaznsfOaOLwt+4WSpxMQVuMYQ2un
UiYybLEEj5aB8/xtZr6QUuONW5q/zVu4AIjSZOgBDHhO/l2AZk3txGlpwedgESrsV8oilM4a9+m1
GhjjSKo4b8qOrfXNlRc6F/QxdsngzPehlc58DmZoyTobbCVv/5uPsvPM8I2RPoNNVfp1aYXTMljh
R7cN8r3xQh4FDgX4je0zDkkaRdONu0AloWkUFUJWbmhNNFTh1NbpyUIjM4weSaC57tID2b9XgGkV
HsNmI5ZYk3vIYOsOpjXIh8aWWK1vLGcNyFndxnpUxT77J/biAM6ush1IkhlIckfRsyvN5pI5WgVA
BNnlbIrTB7rVAnWO2X/HQrC8Dc35fZIYMIumNjrqrp2c7ia33Y1a+c2p3iHpcdJ2RlYUVVKqQTko
0riqVKRHb5eYZmuUIddfFyZOQIxfAP9P34lLj9ukOUD5sI4Oa9ejvBEhDxOBG3I4BpYbsHAT4WsL
c4rRjWYEkFgakcnsRJ3rmwnmwaMMLt3tMvwbQ1PhnhktXs/t/7KRrUScDnr2mbRVHEFXndjoLnyS
xIYPiKQ9YC3nAKBz7QxNwjwYzkmM0yfGGrj1kgUo9I1wkEYw4ySjEa8ji1pYrRfpZDH2sPvJcSEl
3eSM2xcbjgXf6uA2F8Gcql83HCIsx22nH/x124PSHxxk/i3uCXBrxWPN+6mO9dR/3lsSypaCelT/
tqHgGrcm0PlU5//Ohw/ven2DmC4wFwiL7FoVdW7PjilWL/TbHblUDzNbHyFFnUQQTWJlbKlCfVM6
A21SzsJ4+19M8KAiw3zbNJJsyeFLwAhqCIrLkIcbAxBV5rJeDHcFaIOyZmRTCel13sI5NWdrVQ+G
3bD9Q7RTjTQD2fHQnGB2WLU4GSn/O+lXOhI2dbOVABRjvT2YEHtWzt7/kc1spOvnpe1qM1IjGXz7
+Srimo6iNplZD4MWC1jVW37PeA51LOLeQxtiCUAqEzTxF3Wq3uq2NN3B44bYxdawBCsP/yaTHIlJ
mrXxTL+DDJiwtmf/vZqyHiOzumvwDUPc7YCnAFJKr8oWL6VBW1oXPvFafeVULfU837QfmNcyl8m9
fP9XqDU598zfnl/8Y9kHpnEEFRMUxHhhJmUHn6XFZlDywiGlJvgJpst5jTABnC/ptXJxUM8pzQZF
wy/n99zJqPbdVJ+q6elek1lEI1uFie84hwUrGsqXn3yPCi7tGQzFU7y+RH9SW8DJH8IsiOQJs2W4
Ltkzi/el+fwkulDaX9iV6hmLg8unhAM5MjA6rBJcKMPQX/0CkYIZDMRrU9m8yrSWSIlaegiiNe0G
PP/GxtUjSxMZD+GIuzSezNmcUvnoqW6vIBuFqQ+iLyzR78yl3bk9Hg+lcTpl2SODQd/v/lJF50zv
4IjRRChR+oaty7v5GblGAqP+WpPAG1PYuPw/9g7yHtwZX6g4XQVrL4Cin9hxqWHoJUzrR2WWxy4+
Qsq37NxH1HXPUsX0vuKgsTXXavpvYTYdTGDejctEjQoZzX6nuhiMsSLeprR3Erkd6vfbPGJxgHAt
2xODY4naeaMs8/CtIeAWNP2jE6Wu2rsxxU7FeNlguWG1tcVUSG8cRs+Hc87Yv/2uR95lkdoxR83g
/xtYRGGlNRInpqFLXRmvfKHKuX6s1eH7JPUpJdOsHNwyXILhsBLHwsQDry/5eoQQhH7tnkYj9Pne
oQ0j34L+vCOZkfUh+/bpFoh7hS3oO305QFlKbax15ZJz9RYy6hb/Ai5OkN2cfE5XFqAKCvkEr3me
rQipr7dTXtgXHx3ysW/HpJowEUa1w7Dry0uj6TEW2FTS5tc0Dnmsd92Ui3ndH8d+3QkXH6EzqvB3
Dwa5CLhRkiVDpXD93vtJLktqpBKMTjXHK93HwtHJ7H9YfeCHb3v9b/bZLC0R3X6vILIOh6N6n4WS
OMkr3dVOwnmsRdC6EU8N62ophcEd8b6aKUNyGxh+nXbDiEO7mUJofoCzI/4tEZfpBMwB8UnIb5Wc
4Cv5zhDxGDK8nNCGyjuAXwggtm3tWt+Ng7kJi0sMSePPrlvxAzX7KpZZ39S0VhUX3yAlNhQEvcsv
pFdz72xx2j6buGeLrl9+aEHFPRxxscEzpuToqWHCsUQlMgOcLwn9fCVIt5xW7pMb9GCjjQsiM5k1
3ea7+MZDRIO+YvzjXLDA6gWEduAW4LIOEJ03gBJXd12HgQsWTFtsjbtnOWhPPkR5p0uYSBU406dM
SQQMudymrS+Cbl4UyLf2Xv3miXeA+3cV86cLmnpewSEOCG+Oyd63uxLW05XJAIfF5jzf6tioJiwA
IS1My8j7rsjVsz1MftUtjpLtTWme17mxjaX905yaAcxZPVVcMYwRhJgYe7BKQ8gTdiECTYKhJpjr
x1+Z7MQovFzbq8HvevV13dbrLRrh6GSBwqzVf2t+x2vh/PLIaafXNZsbFxfzNFbO1rwQOfltqAYT
nQAFJP/cQ+TrhvmsgAHBUbg+LBHBp2i/j0FvOcnW7+EeEpnuhfnJRGNRJcWvl/tMR+Ilpn0P+1V5
baTM+P6U01kqKGyk/Q3WWdTyXJBSW/MxMDcdSSZYpxU5SK9pnuECzrgm7IGd1Mf+htSMw0M9/Km2
bLjuKq1wuYOC2jacJNe48DVzFUCmtbPUoa0FBnf4wiZPtIAx858yJlmerAhNKtZNJVCJOOhRrZqV
j7HI7f9Et8hFbrd7nuSvmR0oJ8grFshZJPA4wOTXc7lG2M05oT9wbYyyjQ7wPDzNnnpYmpkSbm66
qQyEn0Gd1mj3vAnGucOI1fWHw2XJLDaAQ9s3r0qaImv06sCkDIMwY/bwbNynIRFA0w8QrmhcB6t/
RiMbwFc3Guel1QOzkr7pKnUlTzP2nCGC8HAWY/eA7y574OQ9EV2xWnysD1XAeM6O0K9o78io7p9C
PVF6yB4fZRtbcGjMbWZ7aSxWy7Gk95WmBVtJ2aAr2vATjrTK9Jzeqqveot05maESkqOORoKVABBy
TUpezQgpTr0ZVdqADad58XcP2yQaZVCTXspuTLrsfmhCRmZLis22/JltJdVrP4jAqEAWlcPHA3yh
Mv3Vtcea+wqbbTVi79zVgRcL124uvewMnOQGmE9UPskOBN0lewYtpGLUhc19mFLhhXu6YgFoVzMv
CxCXTkHWHRrIhU/WFc0gMm7dAMACZd9NqzKaQdi+EfWy3vCRYzrVlQWMX+JS3MR9ElZN+cqPakwG
mncMg4lRNBWRK6r+6WubGLQjvPUXttxlHBslH7ga8xp20+CRCJKj+/pVfQHXOUyC/nmfooBlQym3
exlyN4OhBK+FAD7Zi7qHNwEW/vxb95yz/j0XRAKwUojpyXwfbXy78d01cX4pjrJsYxl/3H8vUTtG
HZ57bcfkmt8gzujF/rrhwyHWQJTsR20h/DA55Fhy+tuljKfdbXUyV+qoHUaxfli7Qg6FLGnamjUa
zgYqixmoejco/p/nu7gsnB6xAkq7JkBhUapWet0PL/NBl33IyCdrhBPjAXoyPZ3MBYBhBqih0l4t
7p4onul1vg15CnvBdHlsjiLkZdR57m3/jGeIF8hYHWzLUYfY2wRltXwT/hhUw/AUonMivS5zkVbU
JOGhASNkyfV3UfOANdy+4jKYfo8fs9bbQbGFSZdrLpENxBy9qNpvDh9h6q6A0tmZTBD06UADZMB7
SHpH7yxRn/0yyHTg8UH/p/CvpjaBXmNoRuyA/u8mub14oIJAkmQV9npid7wLQ65J1wlOibCvC6N5
SvsEPM6hwNJvFwVX1xUN7zJTznu5taOawy/tGES1HncZwyifNBHJQT+nLSuoZqbTUzjfA5pTXaOo
pXcNHQ1glMcdXY7+3Dpxyy9U4fbZ/yswDcCUP6HTZFYrfyUywQ1KZDddUVWdEUIKjJgBBHvqjroO
RgOcS3FBIZuufyFqewYB4WFmrW38RvqBejSxpPlDpftwrr3TeoXOuq6arxRvUfPXi42IPXjwCJ34
UiF9bbHI3yik0SQyesWwn9oNWhHA6e1nr1ohU8F8AFCTw2JSLP51TrVm/9pxsv+NX1Neiw0bnigo
xb/CTExZGmISz8+caLO6hs2eI2hdfzHHMEqDox+H6ekkUiz1AJDzefSaIx52J5WVQvnu1q5FAfF+
y+QMQbHeB5C/vjQEtckuhUkVgmWeRsOoh3WEEqpCdCMGHTvf+FHQP5Ss9flcRSKjSb+t2l1XUdFS
7QzF7dfqVGsPeYTyk8D3tNtvKhyzQGV9lZiCobGjMLzFcoKCiBCF5rj6mSmKO70ajFH9K7hvnw/e
6dUsakCZxbmG9bSlkHZpGoLtqmgNmUOcyiovPAK5zaRH0niKwiLvct/Q5Mq0BXw8A2wUE6dqPoBS
w+NK+9HGtmz3kDeuZUpIVkdQ6jKR4U6gEo8X5hil3wx6KtmTG2Kgm1DskcpvVC8bgaHc5XgiXFAv
Wt9iTI6Ao69mchl7M8qPnvyH1TIrRu8HkKz95x/QOXkrONm4qBcngbvtRkOhE44hkdt1Ns4T+pxp
rPK+SB0OiMshryXZ/3BpM805j6AzuNuP2fVDVqZjhQcNguA89VHw64cAPyz05w5ptQtbOxl+EJYT
x539d+HopabBA9ObjqUQoap4TO7grTJeEFDTCuUWEVOIQaeCVxvI2+gEVJGjqMYj2jXiiL1Ib6ev
n5O9HjNkqhkIWvEQis+53eD9H4i4hRBCwqzthtHWuN8sFYedNhVDjbTOFSQ6pJp+yO+zM6J6JjHu
pwJmHtjr3q6V0sjF5Ox4TiVet5RQLldlgsejabHpAbJFmsXa2hThHEd8cr+BWMXy1IiAlS7dxhsf
a3HxlbWqmGgbHGKEohgb46IUXRKUHnCylyD34N6dNOFGUvIITfExV9g5nvyInvwdwyALm80TYmxa
Zq/gHJ5OSytK9G9MJvA/8qWwN4u/CqO4cSppufxFtpfCzcFLYacnExSTh96YZ4v1JKOqakpTPfbt
WLuUnV+lLlVF12Lwv+S/DckswuF0rjrpirGwK8EO7sNsvnvEy7ipwzNLvsO3qt7RUeT86GdF04ai
bBPaG4s+nh9t6bwp6z/NOW7+x3pFbkFhLgygHjGT7S2ZY6/zkLdTriKF/1rAzBh7JnSKd63wOTUH
bjsL9RcFLtoiLYhQGQdI8ehiTo/mq6uS2M7nF7A1Dc2p5h7x6VlDnw/7Gb8tAdVSNs0tKKHiq93I
ip0Gc6ETwZqR1B2hBdp+Ip8xfV3OPv5uV/+gD+/LcURSI1hepcuYEnrzzbEfWeY8aSfqh/izIiE5
oSJRrA1alkHTuU8dF1zrLdaPjvYnmE6J+75cjDIW4vsKT3LUwC1O87G7Uh3SyvfVzjdPj+Ked16n
tRUyrhJuk7BTnEDF/lqZJO5uxNaNom8vyBv8URcqeASQH+bEjfIDNSwLKS1NRk9/QtyMmAxkNQ1v
7n5er+ZzvCFuCbuYaJo8bzP0p9Sx51eR/IB6zKbsN/ycBwkBYKJn1j/3lXEpJJ9bkNOgyFc+KlbS
1WF45Jlrq6E2LGqsASFTZjbys0cvMPrK1S3kwYgFqB8YfIzclBJLOqUf7FVge+4CdC83+DkfCNDL
Dn380JKRBRcLPHRk5zYqRQDZVvge5/1kC9I6yG3X/ul27Ko4rGrhoAYUFDxnVhcjSbZwEp/J+K+c
r4Gl1YBq6Uuvrz4tk/5nrMP8lXgxuRTLrw/bh3ofJFQove7Rqr/mphliYbfkLTrCWhRrwGkB7Y2V
eKpMBoSxuVGW+ddObrQUj20fgYg3kMKUt8dadqxpkn+FHEGOOhbL/Mv74XD+C5v1pj6bge3dLfvF
bonSmd7yW0onQSMJ/OJYEGU03eOke8KoKN50Q0h3wA86844+Ns+kBKj98KpSGhpG1aIgK5fJSGS1
u0coaVLTRLX2lFqLZ/d4fu14vEc3ZKxloaVJvdQsQKcKoVMuN0EV4DiZNpi94IE2tIHEgeaoCez+
l1olysYxxOtkqz+kQVndaAW4uzPIijYjvg+LM4KHbPYgjtO7zI+SQPT8rOclrZNjmjZjSt2jKeeh
rWtYw0eLLHRmGl/hcO2kzzaHlWBvOtEo2PVhVZzFPRq97vPDnbXn7ztXqwpBlYDLXxK8OYfN+v7b
2/urjM8D8WJ5luDCojP80OGPYx0OD4FrFor1ycHlTnivLzQ+chyVOmHOOCfRMJKppCa3JW6vtW5u
PghADAntHoEn13vEAffmDcFvv3mF9PBm0VQdB65l1fAqf7dcsP1xzBVR1V+dh0SR/14Js146BkuO
B4cTtYrxhsj1t+rc/H1MGmfXBk6wTVNz2PkYgW8iGr+u8Nf83Ocywtshc9WNF4VmgC4er+DTUBGA
tiDKMfc0mU/UGEqw36Ilnvv7sioMVqVY3qEbEZeJ0NyvRsqbkGQJNI3+CqfgVC+EXxPRUB5upB6z
e7+ME5vF5SW21ZaG+81bbHGYO4TQQBo6GGs2jh2pWjaHl5X5pMmD8AAUfJEOSJUyYMF/hqSODdZ8
hqt2LHiMC+OlBP+LXtdrAcYhmf5t1/7FxORH6TC42Shi721iH4Gb0p2/+AKEXkUTDLst/q3HLJG3
/WyGXL9FyMZCXYcKNxeKBny3gw56MrbF2H46oW9ERqh0W09RBEPMicKZtaw+hcrKv9vW0Xe8UJX0
bCwZMUNj1CMalbZGeEBJWpSUetwo5StgLD16LFJEgJIMd19R6q3092QH07ZUNM93/tLH537X5V9G
g8X6P1XnFBDQpGRyASGWA96/c0qDrWVimpi7Qpkfd4YfQD8C1jRzFj0v5fKHYneBKoRweab3dK76
ewJyR7MQ0s2uNXksGFR0cqbJYzB76Sjsv6XQSbf+ckXTaRG8cksvkYo/SpWK4E0E96J4WX7E/SH0
rfcpcGywaOgKjqjDWyCSkuO9WuRKz7CHuLM7ECW/N6OumLBI8TzQsWoIJOqeaeV+ZUdkOGK+c7rv
1LXAl4QB2UeBiy4f+OTBit0JWK+GGECZWxQxGLCvixLvFA/knhiTAzW0Yz0pvO3Ru4OLyrB6Qnrz
O6yLU7CMBxqMOq7lm2Sz6x8BEaVzAf+SOqxj+mubWtcdoVU2AfiB54FeU6NRTHeLLYNeUKjU/QDq
pN9Bz5mkF5bb83j4l0ZzPQaJbgAas+/arB8WLS8R9THK5h35p9bjxQWTwPdHGOpfdO2fsNOQPJdN
yZ0Qu68GUmbauc5wlo45javtW2KDMJZl089I4tmZa0N8YJ+0hb3F/gDvY5hjF3F7vBrSdo5q3MbZ
OgdGe9TUYAXNIWqhBJICQ66e27CdCtRLAE/VsrQklx29vjTwQ2t29F6vszptX8m+CJmHd7O8cNZ3
J4JZZxlk81mkn/vWymB/G1XyBBmrPhO3ej/y951JXTX59AtzA6ku5z7N7qEHGJb2r7PW428tUzu9
0rrJNoZ4AVMuSvbCTAxpH9fG8cKR6MuL32UwWEFRxf57tl8viaq1tjv1OV4r3EhV385HdN6A+x2Q
0fJwjqanELqr7ydRQ2LnnIn6HWbs33fnRcWvgLL8Z5gKxlDKhUvaf3HuPdeta973+DsmT26L1i4u
W8HZRJB0KRizGUEpGZl8h6bo8L2hRlwrCwzOhYBxZqzZSvtfxJKjuOZ9MFw2F/HkeEHOwyJLn+vi
SCZj1pCtENx4pPA0Ym6MRcYWijaG/vAEd3UyO74BLRf018Tq0bUFmr9x/HbYNXs/tuquRAEjYXER
FMKD8zo33j8LfYSqqbAID7PnjH2bPcT+NlghHwaHle5jxmKCSZ3MH6RQkpACpjovdpnYG2Hwksf2
ZZdbps8Stf0ukP4x8h26A3C8jvAOd0ySFhCJBE2C0iKdO/GTxDrATkoX02aw8USgHB2v9ylynRo7
J+PuilOWrG9U6e20tjVuw9z93ytItgwo9y3LCmeW8VByigBWJQpEVTOFQRdHNO61isf5ZhA2fIvr
51Ao9D5a1qlatStjLiu/9Pkqo77ZbapfzGqYecXNyvFwBXElUwsI5dxYBT1EWvVAtW/kmiTjn5NW
Sc8S6Kg0e/h+C86nADIwN+Dxqk1fNUl4gPlr4upimVpuc99ZDKTAAmMscIc4OnNAhrZCsUdfUZD6
mHBVEwMaVgffZ9Ox/DtGN5PQysPUSpOhx4EJVJ5vb5pjuCMUZQhCogyuJphgcUvU5oa+mv1KeWoa
dEomcKLE84VGH6wpFPHPU4oCcseAksXCLxp8Bt8gtmgBp9s75IOBWItQJcVM44UuWzPklQVxMQZg
l6BdpruKVlOLKvfcOEHCKWDaF2YIeHiMaKkNpUBWkmcoK+awP3hfkFIEm5f7ehktlXiZt+3AZm+a
H5/xxQuGaRJZsLpULbAWn3SJIT4Qo3b1aztOyEGnDaf84XfVbGLsf1dvvV7OQa1s43l8Al/ejpui
DzURnz+P4b6sBALZqxM5jyyba5xNbR8en/W3NN2bT30FdMvcnCnHww3pOp+pImJ+sDYKP7LU9Gbr
ez/L6FKb0U1lV5p3B010g0K+46dwua+/ARQV9G+vYSqrU81vPd86yHOM/2obxsKbfbNs1j2waRjf
cwABxikIjV9qBLkB52KvRIW2NgOdR3WeVzdGJgCTytU9DwmGZJlAVPC1ZJ1hsRLqCZ2b6eaZXTAO
Kdf/Riwd0Sm5CoeTwkLKhxWRUnOXwZaP+ZuNJ19W51oQRx0UKn0R8u2dqdZDlkoBz8/ClCDhoWHT
p2oh/NKFSxMGUDryFk8V+MpWydGyzh9eZNyzQdROLI+xwUZoXxUoXQ9m6cbCSRLv5QdkLmFhxPj1
71AgJr/5Zux3KLbldEFcM5tyRzLpuNOteCsKamUVeYGwj4/VxZNSx6LCtSjRufbhPZ5iE8jEHuma
5MMAL1/uaGA3UkRdUKdT5u8uotYrpmqkeFAvawFdT4nKOvsGfLjww87QwjCCFlFFxphbAWkHCeKJ
EMOprYHIB/EoYOjO/VG3ZlvGiHi2Vx3rfBqYKkhsH2kMsOniks23K/AiJa0Z1s4YADsEwqmfsOln
kGXW1dz6AMUDg0xDNJyFF0EbEtlp0tQ3um0RGLCKhYup0bYj//FqaVJuLiYDDWVdTlqqZCzKZsj/
KcN50Fr2Qhf8EX0GhE93TzuvTmE3WnC+73sN6pPv7TkeWlXnNwBtovS29oFWChoIoZdlS0aaev0d
AynvoPd1C8MYMhrYgzMFE7RZkXr6HcCM3z6USfF6PcY3w0f+o0bZzFYadiiqLNV7MMVzQdHMdeiW
epcwuAS5AVqyE2hDsKaINMsalvUWyS1XegllhIHnJfFiTCWRfRXbiJ6KOmun63X3Y213vJvONznJ
MWknq5z5zYH35G82vQfja4Iobaj0XjKVqkMhhEwtOS6+8ttoE5KqW68FsADpb2FK/qOPk3D5HdkG
jI5EQMHtPHRukO22/hoJSabU49CaauHYp1z0msGxeBe3C8L2ICLanUzCqlq6BeYP+4XSd1zTe0W3
+ih/pq13Zbo5mx1WbiplQfyXJ5AFMAJLkAXrlym74Sops+aB4JjEsS45UfgidnihFcmIR7mNxZxn
is3+rG1NNJ0Cc8dV0ytimoDY1EKx58aFTyohSKST+EKTqn0zoF758TqoWjXMSFINSafl9JSDSmZZ
8MeRwcjoHWClTw59n5kWP39Y6wRfY25hUWuwktWwS1ymmzGIcQDFlpuE+fYy6GlyoVbKAbm8MMXE
btPE60QnOUIbH3pCbNq1effAsiSYH1+EKH6Z7wr17Np2wO+h7dLOrMtsOlRAb2yYGd6Ofs57wntD
a9aBEIZf0rEm1JyJP1XuBvT6AhjTr2G6i2odMS0O6yNxcYVaGJlm4F6BGMl/JpOVtYlvKfDgEdyx
29VuHmJQ5A1nvukd12p9HBKsHvUo9R28DPzJ0CLCNpQ9gRYFGjQkFclEM642UBYgH5cnZf7E71AU
2nyII+dZ6RdZRqi9BAtAmdXpHKH+mBTqR9NmNsLcULtb4lKmyyx2J4JIDSM14voM6/eWwIQRWDkq
+C1qv+ZkuoHzAu3EyPsIwvnJQCf+MUkxOVqYtnWoLNuFPLStQqpvn9Qh82I9EabXLszBcUSB7zw/
t6vMb85i/rS4X27iNxfVJn1Js5TC4SRAD3hC/Gx9Tg09WAIPJ+/cRf8ImQ7f3c7sz2+dD+jrts3W
rUyLj050hfxr/gBSDwfQCz2+9ofWLKdEGfky9pF2DNgvL/4Q/ziHl5R4AvWVEVezgznVFMXsmz5z
8qBWBLM31JE3XKb0kWx7VvlB/lzI+S+MHUcY+frVmLaC9SuOOsuoJnhrpoE3fsk9W0PSNyBaWarW
EUX2F1NNHUvHJkNW6ZONv8fxzSOo6WkFXOBQQzvWw+C1vbnHqS4XaS8DQ3Af5/Gx5nYDzB5vzSCF
7H0W0pGaDpnnFyO55LZZUc6Y2TuJeMrPp9zq3/gdQ3m5ARFQbjIUFqsVSBiP7njJ8QnAIXAootGn
rpikVUQdGx+Nzshp2fQJ58tBet+xYv/+HrwOsy+7AlUf99mYzpwsfzswH+k8i20AxBlc5l0ffbgi
JzhCCI5QKv31+ZYr2FAFawwsbhmsycN3dSxUxYMIdGwkBTFDDnG/mYALiFrndPRkRl+Dp94G/UAN
6efnwR6ICyAK4N+DSW88BoP8qWO4R7Ug3nKGBVxobOV2alJMTRTjdP3reVtvYRecAH1kEJgKxUgY
rX73S2lrZLz/hy0u6g4IeEtsjyZ2wt2+khvuH86OaFlBmfOVvRC4m24YvibhNQ9/Tvu1DI12AFNj
Q8i9H8JevHm3rMY56PSSZS1Yf3PZYGZXUrrfRndIrZFLgQGxe2d/I4iT6UvuEu7TXPm1/TllIwRj
kxxBPasqerg38R09d+Y3XxEZ2OjbSxTUZ4IoogWOEXe/31HPwf49ORJ9y9ZemYGbgfODVug0QEBc
hj/DFK+bT4A9g6VhPuKVEncCVOWGFhEtzuBJGzrADmQ6ysLZBSObC8z12qdxIhaDEzHlkzvOaznd
wKXybJTaOWPHnvq9Igv3vPvfZ6WBxY80zz8crm2prgX0j9PyUw3fOboNrZ0AyG0WK/5c0q9t83gD
DDfTu6mqc42xQeJybsFeiDb/aMoOB64KfIcLHzVMiM05DkWFbbP2aDmJkgnY2ESLgg5p08SaxPkA
cJeFJhmbIec/NHEk3keFq+4Vo79pZEo0Va4JLiXBtZQTisLn1xSfcICv1oMdLr1BjwBfYsL7Vy8m
qxHyLYgTu2ATvnoKeidNi4C69FjorWMyxuMUJTZWPTtwJAvKAeFLToI65ya/7QXwZEgxyj1SndOE
qAlunJkyadsi9TalpNC4y2KEz5QoMblWCDvOu+vc6ndGGdb/dkAcQ5YaAYHbyy1I1/5ZkiGRZAAi
LX8C0mo5+kkOZZgdFtg7WMqooy3RNFP6qHoiSkXkgo0zTGExWedXvsY63t7cNAxNvgfndxM/MmKw
NoWN/f7BsTmwsDOHL9LwOde4MSPucJDX84zUziw64zcYhsvyIyRquOZAOip5rkEMQIM03CaXvYIe
ThWqobIhu5SMXYAp6XaDyNVdBHikjdp6dChndqI4Lw/jZhb67JdY9IO8Om8clHa5UQY8MncyRwaw
cIbz3CinRRLuob2innRXjL3xwqrryYpuM9T32g+CQ7E4f3dkSDJ5wUJKnQDXjNxSwsX88vI4Nh2e
zzzFfFrz42O7lGfOezWP5fmd9LtAdEnNrdt/dSRGswaMzX+sja8nwqf4dBaxrOlpmFFeEjjXVUn3
KaIMCKyWPTjqp6hdXrmVN6DNQyj2WsBDyn/4q9xIbqDGONB067VMp91Yw2DSh8R+zOWatOY4puBi
1Pc7SQLRqA7iZZsbKeW+oDstj3TRvKd9SKx4455yyXCcTloZKAWNev+4qd3zVP8+hCPqwBxqgLNM
S+qwX56/jN7o1oC6W8tYwJ7yX61kCNjeVOpJSpTJaeHTDWi+mbNKCpWbn8MVDQZQm+QzrWwzBoFp
hwS3CeiAkILdvqnMUJc3Yzp/7JERY8tustGeGfzud8rnHVJ8LBmKBHLav2UgbhvCczW++MmARRgg
c3FcculvmSlcKH4fJrOvhyJuV0Z8gbhDc0TMTKg4fMY2Ty6Uaj0GhAanZcIKFgktA6Jfp6quyE2y
lCyqHFO25JUvTT+FL8NIvn7DnRVSSnBuXzLGOC+pbY5eTW1bNWRv9Nlt5HbKi9B/ZlhU0eoc07O2
RRDo0rdDFB/0/wNW4GUfYAahsHEGyVAgJZ4SnGs4dssnMttnE51yrRt0r51WwT3vdCKQWvxD0HCz
YndFmutTS7FU+TiurzjmFETkMMaft6McH0G26d/NQ3AKYeer96uiylDM6WvyWEnUINAg/Z8/C9F+
CzQEbV1Xrtj5BwGBG9hbdm5ujyzxhjtyfosMb1Ma7gLgcUIsrk+yVxt1nMI+IOT7iZifGI9Y/jqP
kO2KrSC4zCW/NBwJDkeTSKbMzPh0c1Hfcq+twD4uRN4e6iOR1ZNY8QgW5P23lcDzluHEFginiDLV
8QFB5OvRdz2At89RZvf0EFhkEg4nedOsa7j0QYrkTgRMqpFJGTxbXZ0ObBzDBdk4RLG0tfvM0Mnm
h9HN2sipCUtJuyImSvDqORokdSe5FwFZ9zMUrp3Sv3u6vhIr1FO4MHaKA+Wq5/94gFcxMg2qWn3b
M+Wt4/sfCpF/DgmX7X99nHdiTUmcaySFnIM/L9Rf2yqegmLzQwit97lMpcG9BiNNjKrTf3p4UnHV
S5XXpDmMxJoCXNsUyq7tmRxKVfMPPvad7CXisneKevSdbZlWKfjBVr8KCgWNGsFm32f9U5s+SC9P
3SyCbSd/KdyOayEgQkHN4ZJzO3vTbjnGQq35dvjxM9N/+xR+DECHz3sEDJhC7BWipY8wO3DrNYyJ
cpgu5BnrYeyFx5SGC/QMWsuXv9HxQF0URiEni+iDou4zy3zRsXIjbP2BJ9/ZrZYZMQ2E1LZGQlDq
zvWhBAHRHY2CynZPiCykOV4u01rkf6sCRrYmshLSLC1i4XgcrcDjMOhQb8888maBsIp9+XNQMjUX
kJwgbst5j8dYtrcemlhLx4yL1ViDeL+eR/hvPUodW+WbLs5WT+xo79t28dilAeK+aaQvqZq+QmdW
MFBCWukFvYn3gKH/gI1Mq0/VUF/I7qUV8cmEkZ3byOcPSfffIlHZM9F+L7ijykoGDKyoiYP5oA80
2+SZaC0NJVbtYW0Due9wo7CMJPSY4EcZFjJSawKMEh1WnHmvlvjBik7Q1Xmuw3d7YOgEimS5Y5Th
1NwUPAPsGd390HW+Zvj3B6pHkne5Nz3fiZ9qPR94Harvv8Sd140xtmM24J/+dWV0P8vXQ2JVR72O
BsLH3olIp3G0SbEq1p4ieWO4uyfAjzyQ7gTccB9d1hk2BHDpXxrz4B1C9tZxUASzeVoLCreVfApA
kS/wKWVj7dEWL/v/MqovceVMYmKRTUU0mgoNemUo2isqeCbIyXByQIfnjSGhamqFJa33kcJb8LUb
QEShv2zzOSoG/R5JW1tpzmSvFeSXUDAH9L7WdTWClVo/nHGu2KnQ+1aPdgeTzhS6n5wHiCE9O7KK
8YSJyPHtIsMR+oWgqrLcpOhKXr72f35pdLGvRFagde+smd/WoLxYZqhPavOZH5m75o3izeeD3tAQ
Ne7oPyU/ljye1cAK+q/nqpNd0xc5FpVZqwfIDfswDOLE9RjTfmU9z0JSwhpWmxEgWAkYR3gddrMS
g+GBSmPh8g1ThclsFxeOZZ9ZmeYeec/shGYz9mdb8RoIF0TNh3Z9X7FeJrm2hcJQg3DhtQdt79Eo
K5UyeXSC03bXlNOH0lwxhVmQp964qmXj7bk8I300qKOTvWksCZe5l8RXfS+GFE5wnN99NBvdLpJY
K01YAvOOxE3ibc5ltsu6N+cJtUkOGtu/bJreunOCxzi8/UOCPY2LcrbVPKA6MgKZ8N2upfIFdGfw
e0NgBDDgsPQvw/utnWkktRnkOTd8loptU/pUijJPM7Os9CIoXb3SbWqQlUuqke/yhdAyLy6Pnktd
cetjdOuzEXUpsuE4GiUeUkrpL3pDRkI6P1rTVwNkOH4hJE58nQQrVvk05sK/bB6WOLiHSFGv/cq3
JMqrN+Z20LvbuEAQk+xvjIr9k6b/lyfMudcQROALen5OikzIhzILbLy7WPKHUcQ0TLXQurfXrH1L
KqWyxaYyhxA0fgXfseVws0+6fp36mVb6K9J4jwExRMORvLUffunteCJ0+ww1WJdStVaFZmcLt3g5
6ZYCOPUkMVJZdeIR8VZBSLWhk3tWnAHOqBmNL2iCXcuGDpMBHqrV3IRNLfnZUbdYUiNjMWS3Rvc/
qe12UQOyvKuVXSHTMGN1G3AMR/S2EmQcWjZoT+OF5XwxtOMG22RtFv3hkyOtYIp5Tyxg74Bz0zfP
nutMPxoEWW4KOqhQz3eiHriYc0l24nWhk3TjnR58SEggZkNArrTI/4EDU5wVaP7nx85J5WCNkzij
BAgodQi7BML1nOonc9/J1DJw9Q8bW/JVe6Axu9fgB+JhMFNLsLZe183ikQelQiqpoHiE/upLGz31
hUVZ4/3Iajt6C6Y1kzDResXCYoMWvK6qDKdOhRQ3PMLi8/vSL4Jlgm2uYspgLUgpuHSpzDzPc2Gd
V9ieLDK3N9DUnCiOjwpvLSVk005KFOeYj1xtdFic8K4IrUJkO+nXfD+BEcidoN2s0bb8ESwbRcAN
qLA4bmlfTFwk7x6xm9Q/y+ckBcRnBDeQsKDOokSQdDQKxATE9Qdi9oETLz+9d0skEA3S97aQc1XP
8TIInUP7jVO1mOgSr1+S3G6C5vkrH8ru9KrKNgKGDOYdcwtQxVuENnBUMhz9ckoOtRKkoGXoVOL7
F3Uxwe2neEMCiJjmxLzm+HsOrIwwP7WJNGHfyzEAnieXcfcuG/YVkkg3HibpFdiXuhcBFPJa0e5w
pCvvWf5Z+mWl6h175NiMo12wwghgsijY9+UtMurpi9AgdZkuH/u2F6g8LoPYyv8N1souE/ifuqFk
FmgnHxpWLjvFpv+54hWC2ZRc6lKFLSwZdbSWL8rEQXw1rhr+ZdOQky9I9+wgCQfRhvtpx/BHct43
DtwBjujYFhqr/YEeC3GmoIKkMM/yl/NMVE542sWQY7nqCNghpi+hzyxqK88xDVJPmXvfxGE/WoSs
3o8avu2oYcrgLraj8W4+9V6rjCnCuRKZNKHdaC4woX1zig7HOFOXoBtTizc0b1W5OEvYv9PHWuMs
yjav2mXPBZtyHkeOfGYaHphI0DmDmEAnVZRCYyai0YHse7dVpfP8a+DOS7Bet4r0e7JgiGNg7MlC
TE6LFE0XFxf/faXXR3POFAfFex5Zb2JhrDgQsUQQTQuixSWVFtDeLC8fYeMP12uODNE+fkkRUgJ7
XxoAvRCy/kkc93BRYvJg+w9RBs/Lt4Srkvwx7Mku3yhIipq0DAaB0ILslDK+6DhZZ8+lSNMiSuY8
uIDVvk69ZKgCUkjuJ+kj4eo7fA06xUmglRnJiPhnLaUNffvGcuO0Up+g0A8luNMjtXBjf2F+yt4Y
eNpDI/zCUniLo3gUaYso02ziR8xte6vKerZCKCxGSsouYmNRcAiJvAfRsGugtrfS47LBtWLLeoKG
bGk5EF30rhi4ZL/b0GXiu1w7QAVgcXy9bTKqXiSEhx4NYkhpXA/GE25qWvMzAFMIixFC/A2K8vBV
z0o/JlNbmqdJbGLaMa60RelbuVAzyvIVV9sI0woAqOmxNMRbtsFOaYOGqiGC06BvVNc2gYBIkEc2
JGu/ET5pIP6e4RsiwU7vmEdovRLq2xigq91+PUohCcQ0a32FhuwCkriCb+kB75SZtRBTMn6E2JCR
3e45NpFrTUxhkmKXiF2RwmxBws2VbhbveGrgp4cq4gs/7OOoPRY7yxifcoTtQtqLCDhupCNRXdIZ
bcicshRmf6nW4PDboYc2d38vzxm82QR49hlqeVEkLickVElc/m2n0LXGVc7bbt2POURN5HuuB3pk
jmrF7ecMW/qrX/IwdOACjWfMc2qPEWa3U5wAH2pgs/H621VlZgJVeD0t6GjVB9IjU/jXZB3yagfl
Kq9Yd9x4uUIWwNNujLdW3bDQg7NSL/Q3LQ+hz9It47mPNnzItP3y9YibUwch9BCQ0O7cUS5qkONH
KSpzn0BQKh1TD/fNygm0rQwqcKFfshI7vOO3NcXl5dszrtQi3td9c3I2R/o1863nDNOHzn0eZpJg
DT3q9Ie4UQjE+2iDDpInBX6TyCxxYKv1nrNWjye5hvPYhoHsZQBoe+C04lpcOo1QGMY1aaYABIkY
KNldqG3oon8YQZWkq0FKMZrRL+zw8uDEpLZY7czM6YiDPFCw1bj0o6WzVHOBW+Y8SAL8ilwb/0bM
CMW/0zqvoDNwYeS76ZCjNSMmUZnCeOkc12+reByRKNKj+ldklczIzZQOu4s7FTcJJQyT0cv4d8a6
odCgHO75qRz6WDSUbQh8yzjsCG0biiCIMUzUFFUrX4b1o+YxgglfwIE/BzzddX8kYQtSf9y51VnP
RlPTVsXnFcjgKzVHinKfo61pIl7g5zN0CXLzXXfPbWOK/Qa7tQ2rvMYuI5Y2VBXe5y98TYqH15Hd
CLrYiOn9WcdPOluN2tccmNAnbgA6GyUvMMTdWmsSFzyy7NkGgBdWq/vvqFExMKWW9Ti1Noalqk4k
GrDf0Rg7Iob1V++wLrzQdDpP2Atyx4+kudIWl+LDeAxTmNGJCZVDg3uumJGKXk08RfgkyaLo5har
iVF77MnOnwEhAlux8t8hqv9R8ycNmxDYJUtDn3MavqC+OjX5MDr7G84ZGKqBVEefP78TfWwe2XCf
mMu68Ab3cR69hDIhtPGPBoO+98knHCw7iQsq+4nT00CTQk8CxF8ulfI3SZ3ljCLgX61m+w2KO03w
gvA+FH7ACC5OTV6rpBKPA+O9Y7VOtXTp4HVwK9fBvsj4O7LaZ4JseroCYwYnam/ma+EMAOrAG918
WA47i6fQ3xuOltpPCFpdW+G+UiCZNrdEGbkQJehBlUokq5nwXnyq9ZdVyB50Uuna1b1vCgICdBOg
d+kBMnCO9GeGCQ3Ql2KRvAJbN170pILv659uaG1FAQFjpyYOkCztiJD8C1jZvLgzZ1AJYrtXZ3XJ
OPFNNlD1ZontkpE/uTk8cis++lbN2ZY24MMmaVG47fjRpC5Ym63+UoFB0i009eFRm4yHfXuyGR6N
7YwfU/7bLvyzIg/Z5cuUl+eTXB16QJdqJ78d9h1lnN3xbbnietbLuy5PyrNVrdJ1fG+VFft3R87t
o1wPwwLx0Y2K7b5fTUDSa7rJGG/2tOQ5NZvmXS5YvbaW8vK/NwuPbbzxpreuxhWRcnenVdrdLnen
A43ptJB201mbCNkNVoYCPIy1UBsAHsvA8fMQcyNCBAZf2duynyJVEWCDk8Xyy2NOPnpYn4JjHeGq
qLAyJW1JYjzd/YToLZdN8izs711X5oGVkmBtiPU4si2UphALOLODA8htqiT1fACIG0+AGhzL+YKl
sY8EZZds/qZlRMdc6DEzjhvwOiB9s6wmxhRyJLCRXOSkrC6LPLFbekCYycJMFnnbvmUF68CqiBgq
wpD1DaLWr084vtowshLoEIRHNZI++xIA0Gwr3I1/4mwkCI5DB12mJD/mOp8K4xGzETQvufBVh2e+
4pg5tMME/21ZTGmzLZPeCMUdDclY37Jm7z4d30xPRE4r0QmzYgu5wq0PrLAxNilygvNPZ/89TAw8
D7rJh7dt7PRQWfodOxUF1YFEPzyppXhWVysaNSnNF34iVRXLm46XKS+y0SJcyAgVZeUyJCE1TRo1
Ud21HC1q61+YIV22nh8OIIfoUws9qtXPVUGGMS0Q8/bBlA4FlgRQwNLw1+VlPadx3fgaH3AIgEIf
ryvVLVHx8lWbDcZocWTHxYxAQ+OVoP58vohVckOfVHEPSN5PjLwC7bQosz9nzodq0Lz5wxkVeEHb
jQ+C5v3oi27FEPmq0gdz3/nBv3NmHY9ybe3aheOIjfCiHQYZOFdsxXh2gFMfdRAoe26s5BLGrc22
iUJJB2dqqOjyJmHETlGMLJyofuvENvkK7Q/AlYfthTeN/eZ/5r3tBjd4BYjVk4QNbNy+fPqfC9wR
euS4F75m0DQum/XFXwMYpIyFQu3WZ6CNcWVdRGMhE5bBs/7ytfZ5Ty0+e85/p29LMrC2Xc5xypNv
gF+gQ6rfcpaV4sceeDCj1UafuZir+le9zzAtXu1zQTfpWdiHKQwAGbFogJzfnFDnJFRvrzxWE4I1
e5kXDVdHkGJt0SRMwf+dXLeoRzOUUukvlKN2GnbTi56ncxf21VB/iYb0flegwaL+cDQVYJdPiv47
vCfn4hYIkToyG3gLrBhZcSU+ITyStC8Ed6oom1wzn8As6NFeKbzBDc0anEny2ShMTOs9gY+ur+IV
J/T/zkhgPQ16ouyNgrws6CLerZKqkjxV+mG+v0AJ/wLy5sSU6c9ni50rBvowt96KbSKCSj+SbvKh
9nGKOaTplUk5A3oErFagHpln/qIOKGdCajoRBTgWQW4sQHdX17I7V2X1vIw14u99i0FWpb6ZXRqo
uydiN8mtxhegL+zdoqRZFjGd1Jb8Y2NpzwdAAh/yYjV75NU8Jbgyi4iS88P3k2dgITqF7luJm6Ao
nsZEzpZi6U1AVKGSyGd0hjHcZnugo/YMvm9KGQH93qwb6Hs8ydBTCr/y8v2TsMw+gdWw04yi6P3E
escVP4GN6Lu3C7+pXh2yI4969kxBy9OIuuXBevZzyKkgPT0KwcfFF3gYWtHOEsQHnnpxLoTd6o16
0jwGPtufIGwUEQbidvikIf0a3tYDj7Op3eCM4Te2ODlBp9K3Clfll63UKZr5holO5vtshs1xiEBM
ABBp+jHzEyc9Uj9dvHShp3RLGLUZKdINot7nwYpq3cGG07NpPecpnxz+GTFfRlZzVQNG/G3WeVsq
+y878rspxNv7xkydoeXZZ8vP0qn95px7huIOhATQe0iMOAToGW1HGXJbo3WT/5hKiSQPDo2fhFxb
EfPFHvUlhDWMsY3TbdbENvg8ENpfAA0rLMYWNY4Gl8CjJFl9WF+7/zn4sHRkxN5aM1fGm2siL6fg
PJbO7dbMld3p8e/UzfcB9PsMDA1t/nt8dyaDc95Ekye5/mNS/EQSeKf5vwnkup8SLxT+Jcy1L6F9
iHUIzUgMUHjDILud/4eRstwrqKpt6PG/wG65jDRM5H55if2pWsVJ/7UTgYdteXYUdvRiV7WYeQd0
IErSPoVnJ7/vj6cxaj9TVLDLQ6ls1kmUutqhP73KbnhluMF8M867p+w+zAp/Zm0JUfYpTyECYup2
ebfvoJ7C3SeGfFXQ8xI0XwasE4qzcU5/TJz7obynshRQxZ/oafu7SFg0Oxl/WDKmAzJHlIN911Dg
bRUlXpFWHdAN0WdWowXl4cNM5JNclPA+Fyzer4eramgtgXhzpv7ib0kJwdURC0qven02DzTad1Vc
KnJ5NaEdEw4vuLdK9hb0F9xr5V0Al61EoBR1e8wV0oHcNDHN6Qv2SL2f5DDhvo0qOqeBaVh++WFr
PCQ7CQegKezlnReCxwbOcA1EpPTGgbI+hCIxzozAIxwops+yxNC6G0JH+WfqebcGJtK1TanTAejs
dPi5onaAr19JUWsSWLu7rVzaewta8I3FKIh4bB8On/VouUfBlnZ6pG/FFcbW2x4HZPQIKT+uWETL
JWpwHoRCRAJOR8a1GwoKi6qMDMG7t2Ae3BUuATcP8HLDo/cDsoaL2JiZQ5VpijCiwMv7kWsoJp+C
xB62k82SLemas0jZpcccP5CQIFTY2NAgwANuGXP6QrrTX4YCe9qlUhjhW+MsZv/wjrXepJ3GsOc9
QkqMvThH7dHyoKj8OpphhqfG6Lvbwrsgl8QHBzb2bwEple8/k+wvlFhp18fP1TngC1auMVojK+eR
KByMPzI6FuON3dP/kDfAQxDMozxkhhHYUMLZvhnMQCNWKAbbKDsC/lkTJU9qZR3sQfUA5TxnTBjY
lH99ZZYcA42qBFbn/SbM8NPzIG2MXloXePzzsNJyoz6b+hBuMBr2TrrLrS1wrWVIITUUKJSgehNi
OtiJ9doGh9kIQ9SmR379AO/XZQRGfDWg/RspbCTc5qpJHUNV/+IRe3RlmG6iy0gBDStESCFPfOiX
YrxyDw+7OpfqwLJMgBqH7STomM3ox4xnUvE8BL4OBGzCQVDKafQEh1yVh+2shw0gIM+Vssh71a17
vtMTy27SiZMjt43QuKkrnNQxGmYVUBqLx5GArF3vgSgVWKg94nEJjmZUAC0uDKS2trohXquxlq8+
I2NyPrBP3YGY9G003QRv2y87TxPagvsZ3uuSCHy2CYg9oMduUrccjWQVXQ6sxE9p95vlzglGqIP0
XOo5EnsiivTGg6HcBYK6cKqJXAA+5U2nYbVdd1GUBoT4wJu69aIo8JilgmkHes7lkQWCvr4t08FJ
2L/32ZOxYnPtf0SNXgrX4q48GPx12RIGppLOuwdhIp+YOUJK47FcDCUiH3SFyjNBzkVi3UABewA1
uZ2l7fYoLeUdpXE4lGvWelWofMBEevmJiK7LXNxSoboD6lV83yZJe+5UcrpxiXvSKpn9tssQcvnz
omr2pedV6rMVyek/YXYeDb8Dbem7jJNPZcUNvrdROTMouGhy4b3MD0ioeDnZXaHB0RcW02SskaO/
gQEQ2fbr5Mk4dIOYpgFyfk0ZFxTwPN0QDuKeRGWjbPbOpKBa7Ba9tUFcslE11q0PI4BPA3Xh7GOR
vBe9izyzf+KrNBccRlgURAgSkxXqlHKfUgaDp5Vdkkbo7kKljrUD65wzVE7kxhDO3YzvGKqzhjZm
jFk4ocPP7HaicnijOZMP+RxV7shsokSQdOh22NAI4uuMpNwJYXjypdvHjsg2NVdVYQlmJsAPMcmm
T6NeN0l9T2TgdMve+oTiIaiCTG0cjJD91sThbM9xoi3nxCupCkRrP/k/ON9EbVCYsi82NhB7w5uZ
SmV+AhW7iKiL7UBD7pVFApp/5T6Gj7Nj9BuZCyG9/g++hsAjC+64O0vsXB8yW9+GDW69PiudC0FD
UyHnRnq10rtJJQURKOKXcvo0RmoZESqRkgo+U2EnEiKHBPxOpihB2tJh+OnSr2SDFjzyIQEZl3gR
lBfQpX/Fw1cF7+OscDA/+anVLWzv0uMq/KgwgvLz6+qAIornBhEFX2XAtFkfTOZ/eZLw3uCtlcmL
ef25htIJSBPrdxv0s7t28kazlUcofNYcQmSh1Q2JzXc8QS1zBPTteuhW2LMPhguJI/fPxNy9ZsIJ
aa7UHfhsnkJv9OdULQxlzfipBb+fI84/W4Es8GofuN8wgaYH4P5DXAznkDtyE8w/3iYu82wJZPyV
BOf63RLjR18NBXyCMGFscQDh4rBmlF8/zo76eyw6ZBxzTpX31IRfaJcHgzEmr7BuDGiy1hpdYHCc
4Qvz65HC7mZwAEMdb+DTctzCD6r/MkhFlwZlG1Gb9hg5vRvk6c8Xu2CVeBZDgFjXkFmOAJSvDBDo
ql0+m1stN6mYde9vM89bkbHJ43zMPcRpW2zRjfOmjAkz2RR5T6fUdnDQZ8MSVYoln+sHJIe94/y0
S8DYcGaFQ7hsjnnhz2wB6RdXn/NI+lx2rEchCZp5yDlIaEyElbIWbo0wmxHc4OsVchZFuWiIPMqR
F41oHe2ky++oaKxGDk7Jzskc98aNRAgBO246Gwp3tiUNNKmhzpPKILDF5rt5fS10yE4m7ji4QRqF
sjd/ELQlVQLQbv13XSexc4K6c3yQ9LTW8O7AejXWhJTd7CeN0desykAF/LHoFUcy2JI2AOE/wYMG
uCVhXefsTT8xNYjqEd1eCuuo4rxJxIHf8scQiRBUD+BoW585s4WQaOilbJyMQvtL8jOQQNSDOKA9
AuCIVsUCWqM6+J3PbyHpkVzDpwYMv/pbhCtc7Nzqt/cvG2jaFOl089ATUCdqC6lzHCK6utOoQs2z
Rt7LmvlcKrjUOoA7Sg/aHwQYSqt2ldXQGkt9INFujxSkcJVlms5tjkmMFOH6RLV5amXImzfojmth
GA3Zn/W/OVG0m7ioTngH8R3HR+EKJUYU9i8oTeqxj8oHwAiOk+5+ZfDNwH3BKreNrct3JNO/fPXe
Xdh5KORNpuEj0LluexM8feHtlpdD2+U1kIQK9UNj4h68IXRIoPs2Owe0TVfPwnhMO0y6IoAlCRnG
9JkGtkrGSy5V/Zl85F5WI/RRwQqdY2RD5lqcZ+I3CnHCxM0mhCw7EH7Zv0ZCqtRETj49c51rssXu
V3ffgkgJhry+wJVLyFpGMAVQ2IJA247LyYkHjT2F03E5B5edjDFbvLDVGv0QkFxpYBKwmyp1Tg8H
m+Ld7pbXIQOjdTStgmHnwTKZnvPdvnO8wNcSBz0W9LoZ6uAQsZTokY2kEgS9R0GMqxokT8Er55td
psnEKQOyO/HtcMt1am9jiv3Pc5jOcCIwNDuwDYmBIi+M3xmqK/ZIOWPe1m5OoH7evbIMf5lfbcLP
JxYA9FAvyZsqADvasTYLe7PKu0HrmH6fh0Aa/AoPxt0LYxdOdm9Baa91Q6BOPoXavy10MjwdIl7D
ZGisSNnIGWh7PDV+a2BFrHiM4F+JJ0C1oMwp2iLgQnVl92NiSYearsRuIab2r/8jQXKoGaqGL4py
QY1a/sIPu9qJ7/Xz9AWpS+QvVDc+OPSBnk4oDbiiCyyG/35nKxBg+6I7zF3Yv5Bmc7HSWUkRSbey
dKuEcGCQkneweEb6Q/9nzELgP4YiP3ryw5ocbZaE3OBb+4c+map4KSTFL1euphE0htA/BSA6mlsb
cY14ZtHkNwTMIRs7Na548istttVpXjpDyTqQZwCG/A6uB2vlkBr5EWDeN4Gw8GK4xVICtndXuoUk
r+BGsOpvXb01srhukZUz9Piu4uxktJKpdmTRB1Jh91H1j1Nd2/vkVlIArTjLiwjUvPV47Wp0gg+y
Mylw1NADmaRAydWNOI5lis5hHFmiAuNBWY/i6Cu/eu1wLfEckuAcCcOuG8vHa30jN0NPo/M6hAo2
VTID9y48IMStHBRrgR8My+uVKZgXufC1dk5SUhhTm34ig2kNI8SR/WZSiOuOBoRL9GaeQzCAf92U
4ZXNc2tID7PgxOvUG9oFO5rdgc40Ow9huNqHUg+th0KeVvpUjd34se8gg6kXURaAfb5/bdvzwbvA
5W708pPqhr8CYcJAP+lpUpZ9L8gZcPib8t5Cjjc3aB+NgQ5TbUix2t4ZXvAR9YHRUinHHwuWGlp4
7nvVBTbRVwqwiFtPptn2xgwYFNkl2AaVyuKOq8A4Bj5UbPfUPywniv/C0ttzvjwupk8cK5jjunW1
Wd7959vse4NxsYg40e5WByvSGudVTK8HgiY0s3AJEBiO+3nKmtsT2SS5w+ZMZG8nIvXmhwkmnPWA
qh+hfw6q+v17zofrUlnANh4SI0ThvNoOXS5n8nBbEa8naBiACK86Ahg+25St9tdgksj+WIhtepqy
UHfUOaU/M8/CSBJ2nP+kvXwVPDM2o0PdX/+3rahSD3d04e7LuJPM62q2fuE3eGLoq7Ik13lc4VwY
/okCuEEoyZKDIhItyTfSS1hGfQr6t6UTS/Y29KO8kN4RJsCT2EUhjkuyLFwsM0baoO5yT1aMUxNE
r2/sPTP0YI9QKqIQUjj8CQbMUEeIOVNM3LoQf87j2CVUb/DfHXpFCcQtVIiN3YdKemC9dkgNL6CJ
NFAu7pQ/CySbLkQh1hDY6WfJbqULVTTl5okdHyiH5/nDQSNJX801r0mycHC7b3+XrYJg2Lky7cg/
0pnnPUvwO00RG2fwNyAlmQ0yx7GFRUT1HIpsP+OK4Rzq45T03JCQmZwRz2SYEh0HBhoR7po3hDAZ
n/HMX+wfR1gtBKnOdXn1D18rDlqnlkEXRO6W6PTCuntJZiadBdPaMuVg2MCdahCZmlGh21LqhooS
xMAqyaYXnewwAz60+Tdrq/VpVcejaTndidp0xmKgya7jRlVj+rsCINfi+eVWsJ1WDCSe2oRndzCy
x/9WpoX71vB9l7gTYVS3/0b1PxwMAnQl4l9KWqPT4Y8XUj9b/pkJ5f0wpPvrTEbZA1y0Diu+U0zP
RLaftFY+0EoQzmLHdHXltPXUcY5vDtCFM/wHjsPzhYzHG5mlCj5nbaNrpRoPIOqPaeZyNYBA5LpY
f4yhfg2Y4ea+4iNeR4Wh3N/lrmlRknMiqsTOZIuVJ+neehZYnKTEpuEO19SYvzf7Ha3JD4WHcpC+
rWFyzSh57himOSbukUSBLfx+03nYgbLbERwMueVRS6i/QaKmmzd58J7K3LEQXoSlJBZBQD+UY1m2
7Z+GYvZl9mm+M2fGR1odbc+hqOkSfd1AWqOEx/AN+ZL33h6VCBcT/h5I8FgPp2L4jHXHKQN8VJOJ
NsxhizZE6xqz8foFP26hNa37IC1wny5Yy6VQ1Yjco3/M9ni+uK70LNnseQl9F+RvWxozI9w4hlIf
wMsg4dTOmafM0+QW+ueB/2ZElEjJeS52ubXHlzO+a01csK+oSNNo/+YJxi4EwF09UIp8HJrzM+lE
LeFGZ9gjaa3xo5+dMqO/RV7QPWU9Q+yZ30h8shIimZtVsbAbxtGoLmUsMvzk2H+Cp65i7pWL1aMx
cMHkFyzKCdyOWxC2oKjdLkOHQhJ2oj+qGQF/virq3Iq9pT4+SzkqjKnB8nxkfBeUdlK6JMUKwJUZ
ONKvetqXAxlZe3WF5ZneaPbNLGdzO622TTxygZNTNnwlYLSHxZhVKFg6oip84SMHlnponRP9gxWh
EH4AM9t5o6VCt56lJ2BrALW0wxU5jguyZbRI5/bUSbfWlnHpYSwWkLcs/FNZgdcV0qf8ZwsyRXFv
BZ8XdxI2Ny4m+MEhtfAQxXX+XV8WToptjcYEXvJyCTRvvjCo1sc5lb64qAj9MwUkunenwHpD9mZu
550dXTN15MtlZpMOYh+lusqlR40uqNzM8zfCsWWVO2jmkFVVsMyTuuc/HQRcicGAmsag/lWbz0R5
J9qSuLpA+eAgnH88ruLKPl0ca4CTZW/s48g/yMFdoWDS12SAeEe1/xPqwO286GSoE/nyn7VS8H+g
XHiPlQITP+MAwdqU1NTVNjMJMpDqOKH+Qfp87rkl/2Il0hZvcxI6uLrHiFDI+qsudgidPUuOJRV2
bGzXEcuDxD5Y55oag7PsgPDfIb6PXHgmLwRU1Z6EBUwpS3qlv5IYb8xM4LKxEacXT050SV+biga6
tXPbzmFsZx2MDT97m2zE6WEF/UmDwzAP7L5ppw27PLaQBMOn9YMxdw1P+YmANaFUE/3tDje06a1n
DXkVml5SwMZEie4V34B+pVIWduh0vNzErbW1KXP/O9GPvqUw03A4veE6uO7d7/ws7TlVzXQ03NHT
q6eX6Gs3jRAAT/1vRzwQ4ib1Y8QyxJ5xdMN1jfZvuFJ6tI/7P2bf6w87fYOswqr4zKp6Bwi+kDqn
01M7x9KIDv7eWQiyWSdKFEjqKSoAYbek/i3Rz+z+bQ2zdjixXUt9I4q9iWGhFsy6VYFE6d1gvy2I
WdpEU09ogcMPFBGlQ4Vteor6Nc/m46hVxjQyXInpW97iQ/bADDeR5lhfk5t63CP9J3cuOwEQWB8V
7o6qMRWwnuei1AtYgfqzJ8mNea2CVP88KLRIXnK7Ofz1BTeXpFDOzcqAs6uBr/uuDdDuz/fgjEgk
WX0lkiVeRBvBN/kRDVdXk016BWjCw2yPgD4Knau+AuT5sGeeTB+c1Gj3zfopr2EalphAERizKlm8
TEtMy4JllTKrDi1Lhjc5ryXhxxnj+u2DIrlUXV1DTJn7CYK8Zu0ziDlv84Av9xCk/o86R73AwR/g
vl8cdMLXaENxZJxLjLGM7M4iVV/PjwLQf0Ui8Dx5YAYkBZj9KtrrWZPwXOV4yVu5dQ4ohXtfIUiV
8xd/dOePXKGDrEPO+V4kKyhHlYnjKNPRoN+b3xQ/ij4ixZGTUbdBLXbx/qUjnZ4Zaf3i4HSk1WdK
OxHfiL5OD3+5oB2mWAu6Cxg4P0JoTGbvExZaFBoRT/xB6HFa5L8fgjSYt+GoWSdauJXa+E0hmDYt
nDrNCCEzmkPzKqaMpKgHtnvp8FgIZE8a+LWlMPCnUBVrv3ZJhLDAMSECmKgdSJLa+NcXJ8ybvqLJ
zdtH3tE8Pp/katwYuNFAVLwD+s2Ul/V6cEXZwIF+5+A341yv8KOR6BSnsy22TLPSOCUnfiXNg3yn
RZLVlmNkfel/7cuKXHnTTmEB/Ll4rElby9Ixg7PabUF7RYMpsaBI7B1DOWU0N8VizehsXo/NeANF
Ic0v9ayzTpsWdL1C6szPk/v/HjR6I0uvllIJaT3pOe/sl2TJWXcJEY0a3mNt1keM8vJDVD4RaIyv
7pnEC6xQ6bB6QU252sW+jNIBxO6RgZGa0gII9BsR8osHENUTUSFGNYhRsxKU4bByb3Q8aJqJdiTT
EzaWnGWsvMsf6LuHOrNey/0dgRQFajzHKvjc0DyXop5Jo5Oj9K3wRecpTaC0O+HlrdDqF3+OUIcE
ASX91yUeLUktT8bCUhhN1aP8pR/yKHsIz/zaixUiivbhkzVeLjrKJDN2MK8iyNhIFq0ft2/07hlF
MGPNVauNrvGwPDHBF86WO4RvF5y5k+BsoQk5cSi9gQAdYTb4u5+Mmhjmbc5Zubj9EANnjud/z+AZ
T7XSO5QioIAylAM2y07EUpNNrzYz2LfoyqvFDqO/uiSGgN0+SnmuF4HdZbAxtAs3/mFEfWBVyine
P2lQsFxILR/Lv0La1ox1c62BE4kU9hGx0jRQUrscg+qOwly5yLmXvGhMis0EehbPfKrU2FOpl0g8
Zl6m4jWkW39uEALWtE9gNDsL97LMOsUwRp5GthyxWOc83O9gqswF3SqEeTcG/Y/exdWjYQMTyCIL
P/b4e/9RiyFAvEmAIzwOTtYTpmnG4eDKmOlS5y2tJKVb41WesVivDEVVy9RrUIj/RxnZ/p0gpoh4
qWdcx1HEE6kpbGD0opNeYp77S1EeRcALSLP7NXASoVJH2ntr2Bx3MuJ1iIJcLSqQqLdfbucjkQ1h
9LXXfj57WDhTWlsNFaB/X6oUHcDGtQdzU/kD8CSERqunpQ+onk9KyLAcncBZePdGvMHi8dBfKQ4v
39NGp7ZKeNvxLek/sUwY5MI8hic07h7JTSzM7JL/bVaZwpOFe+2VegnhHp9QlUOZMrRZeGcdv8N4
GVXEeFgM8xVBZ6JqTWrXBcr6//43bTHtMBp4hBQHKDij9aSVMSHfNJPjJoX8Ye01IFyD0zL8HUPR
1Um/nQG0rzyl9Y/01BiNdLwU2o1cNAFHX73oCi0VfkhFeKCGQ9qJUNLo7aNG5gL/pqHz1E2J8hek
JF9L7YTcEDCH9j+sV/8QAt8k6op+KbAXtlB9W+yTLqT9rjL4hKZwSvTqN+Ep/6soeynOdBApqqME
RA34uHM8LzPpfkskf8OX5ocoiGpNRkgdUmlyFHFqf0j8Z1b1/KPNbx6ro1kFEOgoJTw//rSRjpsT
DI/xsyxvQGJ+E4WPKEUxr+pf1kmIcegHrqPh5AjrzrLPuJs13y/YaM3BN/ueC8qNcLJ/18siN8JL
ieH8qI+RnWi5uUNJRkKJgpk6MO1Lo8BjEVS4yqp2SDXaFHydoaMbfGxAmWoiOtXENHZvP57SgReM
ZSATadZryZwvF6Y134DzAMMU1KNtSt5AlKlMVc7hHoTnD07ehoKvQt9qKJ2IEaqFa0/9atnJkj4V
748NPN6NN6SMUQTjK5vA18OTxeBFw8BZrgOwAhRzcaBbBv5d9INGwjzIjnxEY9G/qktvewR5uTyh
fmsohTUPcl0gK69wX7rgnicZ8Ns59uqJD+IMHmYLF+1eswY0WnGfGPSzLWNNQ5uio/xBtfUbvNWL
KC8XN1fecBfakFVvtXkSym7VIpoJEM1u77wecOoSDS6SX77UHvL9Unkn1cFNo3RUByZIeXD/vwj3
41TPiufms6A6hCVqbtXnGF07IkvEM0dTPQn8Ea63WeJxIzRSn8nQo4A/AEhBeAhQuF/lqdgEWrRA
oJHY+mLR/mCAERTQk9zHqLD1ykYS8SS2EBfMBZu1+8TsEjymX8HSGcqWfeSEXfKUY75oq0REXoyn
cNUCPczy4K5E/bSreRyqb3uEm6+moA+YFyV5mZlTWakeKTdE+B46aT1m1JSJ62a31pymyyKb5q2D
4jhEz8M5aak2uZ0x1xcsaXIaogI+aBYd/glJWEkF4JlSbSO46X4cnCfP9Z1XSfzEzQdRpkl4lvyw
1SeI/oyQhwm5wm+/Hco3B1oqQVm+bdDWZJx7YOg8CymiT+yU7fEReyO+i6swCf70hd3qk/AtYOkD
zuJVQ9CPaIgKxUgPDlfWTkAjhW/xCUH5ncH+6cnAOBliquhqjaEdw+4iM72t6/liUyIOqfBXJEFQ
Fc5d9kndtTiUFTE88/VrdL0bn5R3TycrSkGlL3NN7B4BSbRZgOQsjCsnguKVw/l2SC9B2orXKS0b
VzSwXH9BEj7TXyC7jNmlkb/iXn/J/yWoXnx6vHnWNWInr07zkbi8CVtMoT+OTF+89rWVOjEjJTmz
Nkeh4JScEMhSTdtbmsmhDBhFRWbDjVT/X3Z/dw92YKTRd3mZB0SY038kGOblBQKuqNBM2tcG8z1Y
l2ZfpzeHJ9Hh8XI11Bp23Kb6YR2uV15Jw9W9oMx78B1S0lb6is70E9WKVzaIBfQtmUzYW8VP+aJJ
0NH4C8TyhIkkxVgsToPY1G1ZYJuKf6XQfHHt0IKYqJfiJrW1sw7BdY6NHPLrciR9NqhQIPPmISvG
egpK56y85Y59NK94Wyvy6pvszzOvwRWYZRbI6vO+D6kOOLpyC6FA831HVsJzQ3awgCIbv8o143I5
o8zn7FcbFF/KcvukqZy5ZVEIa9oXviFePt2bPREr/a90ppITE7tghiQVI6zpdZRfitXdrhPJ/USK
ngVCaCtnIMYZxUfa8wQ0PlwLEVZ/GbhQYiRECZI3bx0wL94ugdUWP9wU8/NW2Chb1RHYw3qZPczI
Dc3c3pzCFhEBljgVbDPFdjaFY+1+pKzlJHSU6dxh4iF2kB3MOTVfmHhvM1H4JnY8umkLiVcxmOot
MhAW3K0QAMrH8pIlbBwJb3bcRi3pirlhOkclzHqQp59lQ3478MlaWz+WAbR1cIsjiKZiYHn9PRso
nxtFUgnmMxgUhMoNh0dgjrNQlJaq1NtNFjptyabgQu+U5qcGW352QOrcD7WxalBgs8+BO7kiE6bb
62Z8wo5ZAbI5QcXCRZd0unWnvZrBi41siUqx0GwJeSe7Bo5TWfAkFc+8UCIVQb/lLkXCfYlJES8h
0G+4pMdeLITEBeb1tWI6uu0f9nbJGq657L4w5Eihxb6a5p+jwQaegICb0bco58f1L/7nYLFN0sJD
OB7JTNYWxm6Bd00yDWp/bFgkwEuM3gNoBWUhLKbSm8PH0/dXagZOLwnp+WAx7yGtwIfIOzdz55Mv
4Go4BCYl7UeOyCngaLVk+01TU3+nrbQQx4AcF+BHgFsFQwm/i1ssDq5gTtqt4LpcHedZmnspHY+3
OYTrFRvUV/6/MHxJiZhtEPeKUcKvpz7+q17YePL8fWOz25rtgQPMT6613kwaCjae/hX8JgtCb3zh
69YeO2RfAZrGJ9XcLkmqrHu4TBydwLlQxVlajAjGkz75ES0y2zde5TzodGcNhZiBQFVltkAaUDly
/vlY8Ux2ktiHT7DBk8BeFodzHb+7P3qwqGKaCttgbyEnAczXoqCSoNLnlChvIAGpiuCh/9iOLe7O
b/VC81Yqnk+uO3f3gTpie7gIPEd0nMVE+ntIeI3nmdUTdb0pFdXSYK0pMnNHGXDcPPNRfaV7whZ7
TycJx9Zvc0ApFDRkq9l7rbvMLfCNTVArhDMfF0sYSGw6vH1Gzn1sU4bvY+VqAQtbCwWBq0lRhGsq
bESnKXaYVCookkMEyYUdSxfJeT27FWURAfTt4f8qcUBlHKCE9OCcD1DGNtPfvwp2NBuGu8z5NOCN
cb/KtONrWoj1jSSsdXazsvijRFG61eyNNmb+CnyOtznp86jwPEUw8g4aOJ6hRE6w44hVAqit1jNB
/a5zDKatyEPwLUk48YB62Vk2cArAVmyjukavy2l/yw+SYG7xHHIzMP3SNDB/p7ooaK2y/uajxNqi
Y77bnLgpq1S2t8WPhHGz+rMgQBgsaXC+cbreKfdHTC9zb3ST2h9Sw6lK5M+EEX6I5XCHsyTtLkXZ
uAxYyiYe0hse0mOtEWdObioPfhWE90WcflFk9XDdgwFjtkAzY6L2TmHER/WpnzsjoAMwz2OXOFsq
Qy/w9p/HW8b/JEYPGOFY+jpwh81EJUAPvK6e+jtXDqsspbDtDBT5G8UOA4NbPaK4XJIarTtKLOrU
ET9BMCRKRMSEqZl0hRaHarxp4gaQQaphPOxcoXsUHi3F+ofW0/7m39y5pZ6Cq1lnOBQU0joKo59q
rbt6g0OgLYr1ENPcWcG3sC4Ua18OYvEsC79THNtQmzVzRYbK/y1kTcoPMqjedBhI/4qbKE6je8Uv
dgg6Mj8PEERYrRfMWASlL0m473CR188cyl+aAVOMJxCEkahZwiVZX7ztkqe9Oxcrx+KBKnXiwvny
D4iiS2ZOoaxyioFgrS8sYuKuppuBISN2CU5R/mSPS16trIFKJIXE+wP14mTRe15NEwnJHXtWAuX/
i9KT8MDd+H6zK9Mrxe5KSyTzGCP+vm2L8E6ncTC7NwmeIEQM/4hQvY3Wg/aEW4qNgaQTgISEBPoS
DBoYThsxUqeKu98X3CXdm6myaxc0kQiv15Ae9hW1JWHzrf/zpsjYh8gBcGCxIQ31sInnbt2Juey7
W+cx21qRPwsKmbiCYQgjzc1AH1LMDDFHJoIh2DNNVAjjUI3T/HjMqVn1MfkiB12KwU0IzfBsaFMu
iszlrIMBwWjZXy5cKZEFDNbf7+wvLfuNBBm592nPKRLbnuYvQjV6jQ3Jcy492V55MN09Qlg94cji
M7yFIcDqF0esX4mWCHeRmkAJjEyjAhE/Ly22cLqBnn1QOmVEQ2XQQk0+ZcwjKTanh67E+EJ9E9xD
LHhRpAtOfClwwLuYlDs5Jnug+80kU5hu7Fj0aNYp9Wj8UHuMqET/AON6AAs70+e0NoVb+FhMWUjs
carbD5ggw7pz3JVZE+YdaasF6lSVx76j8IlbM+ma52CVrfSl1G9mZnbNEHonO2je67XsufWOMYjp
0D2ObopGnEja9NS67Jc9ogrVucQRLco+upttq20ks+gjJyOTsASf5QoH+2kwEI9LwTknvUkPG4em
x0QW3eSZQVGgSpIrHm/ewG7goiV1SyFIP8vMiWSnHzM1ssGZhTTeMtB3G60Xeo2Qw0vTqJ/n1vTQ
I/vZYh1JEVbJ8COX3icTBahhfwB/7pYgvny4O44LYEDZbRfxHW8QrHsvg49L5hrVZYM2VVGpwI3B
YsGWc5vfnDlRjL2TliZX3nPfiZCnH0EKAw2N0fquKREPi8W7FobSEZJVZ77sa8zljoxFQ47eK0oW
gzDA+UPwi208eIguXEEmX+CucsHCiNp0yK3JK3uArzYZ93tcjFnIQvW7pSCAeYG8dUVq08OWXSw8
Fvy7Fylw5XsRx2kX4AJxBSbkNOigf4KzT3YBmhgG/Rlo0AW3Ys9stZ8m59KB6LRRoT2J9Dqe6gl2
O4u8scBYQ6ueDjMXjR/7P7QhijoYWROG+j+vrr3W93ub8TADJnFPKpOM3wsBjBn1244mFn6GJSYa
4vJq6cyZ1AlMfZwSypjzXAdQBKEXB2NhIswF0GIwu02u0RIyUAY6n6+GtI/TSmul0ZgxF6NOUq2t
al6GaxBAH3pl/a3siY+93G37/L3s+1KCxqIOokh33FQ+BwQS9ItY7ab4KG/bfrdrcSyW2kUizDcT
voOERns4U2O5n7+IcOXzF35hChqGK1CMGNJNxmFqt0kBFa3h0JiVA0m+wDgqkhiosKu1LgFcGdya
0pxAKe0N94kAMtHIwXv9LD0MbM31pjwdb/hAe8Iq/RngnYEWtd5odXj2Beb3l45c/0omB4j31xGR
OKQIgmbgEur6HlK5QSlrkxaQLVHFbuUJTkISwAuCwJw+5kbxLFfabGUFEYbYNSEzKf2SBnJpQCcF
qhPuNbHmrAmPaHzR3r7SIHo7nHQJ1Tanx/qr+PvoKm7oWo0ngy+DfbhRZpmUjpyM2HJt5xq6HCpG
05o4tHnjSvfdJIFmOLSK1FggmvzUHSjwQ94Dh8pXt55C0TNQAGkMwvS7K+wJYeFUHgI6snga1uMZ
HZYgwnOznDUgV8rXgmxw/NtA+BuMNiroxWKYgn/lMyNijj5GrKeOUqY5lMSQjP7Ti3wFZWb1/6CE
3UxTJrWOZb/q9VQhpZINskar6/6nw5FujAkujdWZTsnsXncksgjP/0BdkvQQuUmlNSgIDGcNxcoN
Tw1+llffiBkdR+pLoyw7CB4q8g3M2a9ELvCP8Ai/7fdptd2WmscAaDFgakZGhqe0mZWBfcY4hOF3
hycKYafP9OB+QIsDDqbfmdF5jeKUgm+nOnryn8SHQp13HWcnHSu0TXt79H0uhGXVMNVA4yW9+X5w
Q7dfcuoEIG5y1XWFFcU85sgfEpJlSh11ZAn3TIncyuFmZ9yWxZL7mFEL3cC0uG2hk5k5MfkdwS7/
TtUXQEiksfufC6y8RwLxzj2UtoK/Rmtl/GW2I0P8sEmz0WhGjzctp1bC/wpWtxOt9oj5+lKobcjd
+mlaoW6oOI7rDW8yvHFpJ2EBnr+Aj32PDmu9BkaLDkqnvc5oQv1xTEoZ3tgJrsMIr28HbhI5twTp
1EWygMOFQzz85wBGQmCLBfsRad0RADYut/lsDW+950cNwyrz9m7WFjJjLxPi18kcNb5MLrMHRfXG
SlwC8xDh1HBdEAVqE4vteKHkBXv/D/0jG17DoL/0Bqxq2zOGe7aQn6VSeIbUyHcYLUsou6EHgRQa
oOymoo5zNUkE8E7YZtzijxLh8g4nQheFobNfnK1XlFG7FxJJXlgf/TrrjN9NHW3z63j4AdHelqId
lmAPP92KKZKRZm4A9QF+RcwS2r5b/p/Rbv2inHkK8MMhFUPW15A7aUzb2SQyS6GwuYSyKqQU9GsF
gqkix0Hie5BUOhPfFYr/MP3rwregb4okJHVTfvbYMsluxD5naF1Kmvnn1J41gXSvcfbZrXd8R4mX
YM1bfrgsp3XwQs+S5WfQm6SMRNwVMj6TVWqjgQ+4o5JrtPMRSwjzAyd+FH9PzTOghra4HnDz6sF1
SPZ1snhW1VilGbu0aE55Z2NAmuBs0YN6KKWsFLVZ1bxEXboSbZtIkNid9nukU4MqXzuMw5kv341y
9LvdeXh04s8ItirABMIb1B9u3Yc/3oTmdhVdY8cHhibTI5rCdVFydvSSguHhVDmLPEdIY5dRq12b
H8X/+pZDzU73SsuvNMyB4iTO8KoJcZIss6oUA6InkbCiqRdP2yBOpVWywoJKq6IRKZ8+4SWFZ93a
CZgHX0KHjOYoyYSFFT2z6sdhnexc97nCSWoE5RTZOFYnAl8BPjC1U8/Z8FDrIR9/MkI+Ln74AmYm
HhQNlWgnwTOtaitybFlYMqqCTJ9xpgc5vG7EwL/hKL67i8Vql6vu5BurNdOLfLlRZJMJcmFtIbaC
au82AlA/xg8F2eT+3Wv68WgWnt+7NRx4+/4tAaiff/qwQGPTLJhzuvzn1MZykAdhQk94XErlSCAc
259gt5Bz3D1jb0vJa4x6JUukaORYy1BphMsOxkz0nc8b5zyxxLTi7VYkdvr3zM1zLAxiu21A4eiu
2CfypsQvMTSAO3ERGA7FVt2crsObXqQpyGHO4c4/KGpySHavtSjkLFEDmc6MszrzSP6MMdnoFC+B
YxbiIYDJZqpDxYdseI4xpovoqKwvvil6lgmZWv4vjgFHOM23WjLzAMey+X38N6mhnorGbWnMzV6U
mceUPxk0bWLLf6A1A91FJmbK/zMZoXPyC07DGRDz8l6/BZ/PMOBDgujuYtxOpGv0N4X68fzAq5h0
zMjkm4CgmXHjt3dn7wOIzg/U0kM3JpLWLob3VdKYEwYTD+NPmnNn7ZAa3bLtYMohbpp7R+HGVt/s
GKzOINA2rcnRPnonEsC0H6GLrQX5Wds7IxGeitP0lj7zXbCTwzdUDM2yMXNIaG66O/wJqXJ8D4/D
X9wX5XL6MlqKwFaSHvJxQ7aMAGILGrai6cGD3aovCxIR1wHbmFmdx36O0N2RnKBzV+shlVtJ0PDo
VUh4HVDNhY9kwDB6NnrT6SEaJ3vd21y4NaYenuBc7QJWftNDLd0ORFZI1M0+n9CnihAQRjboHXnP
9FX1cvsr2/Bm/ZylAjChI0OyiYFczdOqYxBgUn9LqcB/1gm/lpNqKX4tjUosTkkF/1J5rGr1NXw6
4pi1W/Hdz/M/X883w1yMVASPO3T/YIc7nYOO8bO43TvaBRlK7GfqicQPXp94lyDlMB7dD7rqKUYY
6TgjydicWXfTHfbdFUyW0ybiX/rav4mM7Qk8H2GxrllzVx4uFGKIJ9D/GFIwzFmj152XF9MKNv/D
iymv58jChff9TsuRoQHZcZ92CneIePYcNWjqNW0CbJeEbCki/dSfDkZolBecbVKHMXJTWN/TUkWW
8WjYrZy7arvlDM0AwUWh2IsRHNXr2AIM1Fk4TXEd59zAobpUjgzek2vUm+2huOiXr0GE64HhXDqv
qYdzgBOO4gyh9hFe+jYmx4xO5+3s+JrlPhBvQsEN6q3cbW4KUjx2n4UIKDGxclGZvLT2XZhbHkU0
21F/AN4Hl0TBjQhE6nmPb1FBLc5e/GgNG2xrrfQhyhb8GXO2Gd7EY18c7ri9LFg8hECcGkvLMF/6
4SkyOlfxiFjX8c8T/Nc9RsmmGnHdCCheDKkBSFGp9Jih2NH3OMaPd7rfsCE1YvbKMb7Z20bIcJxR
gPbtOjPiPP5eIii+tiz8zHm6G+hLzQ0H0x5L7gKftigESKQz0/my7Kj7hARKa9+TIQyCf9o4231G
jw5urooSdu6luszL7jGSNhgAY0jfgHI2z78dLuUU5kIX+6F/T8WVZ7Bz/y0jnR1j+Avjc6X7F+pt
OC/5U4vuqftYdG//AHZu0H1clSXXo+0O0qdXChwjfkJwAeSasyA/TJDyXmHJiwRPhgTyv8MBm5rJ
fNdb5q0M4l4oSaVZO0Vygu7UhnrGPUOn7M+R2yOG+E2bEWv2jiZ2cmpumaE3mHnDVtRnYtIsiQp1
PNpuCPU8MWGVcCjQSCiEJpGUDPgwUY3tI2WiaKWQ5OxkAfr7Zln+SR2tal+4RbT6j2hNYMVvkMuZ
wrMgYuB5frTWFDIzofkinTiCdos7hBBew0B5eAuS3N3unILxV888mGbh0GMYqotYV4gC3Q/hatMM
rFjj34SKe8JckX8TNdi3FnyZ7WgrAR4Y+jap9RpPiJ3B2Ny86TbNpv4z1KPp3JZ/j/TdtyieI58J
xiG/SYk0oXH/LE3c4MteNOOff0jmn43akcQGeD2cC3YDb/XPT+hWz4xvNZEKYI7n5/GFuY6EOvKN
7VBlhpzC2Cc/2tSI1qwA57qvl6D03R+vwe7Ie0OtGa6R7UfPepRfUKJfnC3+Nntb3VfK3A4Ffu3U
vYxZw9rUICqC0MZHXs10CTl2gPHMvLvcpapQz7KyQLkUk+tIKcN4macWzgGMgF+30H4kuiQlt0/N
MHqgh6mcYZ6fsbtzvRvOpi7IQzePE9/0vIpqz7RHqF2TjIU/DIQ2o67Cq+8ltMKDK1YXvaozpCpq
GDKKKfIdLzVsgvE9eAqg600ElWq/GYaW8DkoXOYrhZ/2vcMP+IUIFu6N4nwl0EaJH3gTSYHzUqvD
lvCciV2SXXu3Wi6y9124mLNAQHkBb1FCARHBSIFq7/ZaGhXLQDi2TejWeLVDVGo7nlpsijltj4B0
z/LtnbYIAC1C419qEXLfMxqJlbB26UAZMdjFY1GEjwsWYmo2rsNwbdUVnbqzv+WfPJaSQGIJ8uAg
91g3QkkvM5CgvNDMVTxHnPEdH6nafBz/+WhgeZ+kuRtH2NVgk0rpJ0ed4BQhS3gWdbYUbkkRzAce
SG103UQOF2rH/tSlWPnfjoDeM01zetN2sw8PYhTAiaWuVdKdsLn0ydjuZm18sBvag0rhVoV/oWTN
GMJWOGMQXo7OJUcAbeAddIrLZYrfp6ypk4QTyS7cg7a3j1imx1b5wg9ncM8Pcd4E5SkHrW5isDGA
PV+SlRsP1hD6JV2912fI+ALFG3oKp5XG/WP6fDM5yqksckYBjHaT6fkUvLvB/CaRNhiOBIPicybB
+1cCQLW99/3Hwgz9MNBPxgG260b0hxYgbh/4mrY9YGmOysxZbCI4562AatFjoe5yj74W887JaXWU
S6Fwxs+DVcE8hVxgPvhXSk8j7F0x5zIMS/DmQHF7PbCZMp1hJpzR4W+elRZHfQ==
`protect end_protected
