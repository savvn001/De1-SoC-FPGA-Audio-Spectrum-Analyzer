��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl2!�9�k��)3P71��+��U�WMZ6saI�] d'���5��>x�U�fmJ�Mǰv�Zt�$)~S�b"yÃ{�d����+iq~�Vpg�W�Ħk��M\��r�h-M(��(���3~�޿`9=�^�;��56W��R���MC�O����dg"Uf�!(���*D&��� ���ʶK)�9�i�Ǐ��>g  �x~ѣٴ1U�Ņ�Ĳ'�D�É���,��Pl���A��B}� f\�xпF���Y	"�-�r�>O�?1,γ|y
�؋U;�Xl����W��b��&�T��z��,�d?����j-��Q^�N�4���:��q�P�'����p]WQ��LeE�&F	�'sV���9�7e{S{WU ����\5���0�07qp+�[��:'��(oh�<bڤ��eDI�z�)�ea�vP�~q|H��LϺs��o�vԏI��)�h�̙�Z��l�!��&J��U���EF�z����(�e�C�7�QT�6��k̨)�6���MLX�~ej�};����u��_Q�$���ec��D	�u��}�P�t��c�s&��t�?��-UT�z���I%;�vM���5�j�;���V�����>�;{i�y���c���Ʃ�zL%
���}�9�6��^#|)�d~�b��k���|N�<�`��@��t�}�n�Mci2��=$q�[�Pɗ��|�pht�-���s���9�d�Y�z��Gi����Co���Ff�P���L��I�=o�6?¯�)�,֍��/�w���(��Bs����G��B�[_��i�����;!��K�9��!h����x:�w�4{%ڃSG�����1�?0K�ujA|@��_v�$(��=u{��_��(������@�:�5�7N�,ʬJ�9�}��MXrWZu�/k�M>���g��i�絛�_�'����;E5u��[@��Ȅݛ�-��x�9�o.�u�TC�+00O�F���C����̡Lz�����&�8���Z��|����苃}�N 0P=����	�'a�sv��D~X���`YZa�	.��1cv�7A(�&�5߅�O��JOUVZ���|���R��F�'�zn�<�7d������ϑK=j����	o��о� �Wחm"�k]U�B��뼱�J������i�["Z��h8hB���6	���\V[��&���1��d#�7�P[H���QA��V)��a�y)c�����p?D8��]��7&��?Cd'`���6�M�C��̹LF,{�����e�d��� ������r��Ҷ&����6��+����X�n����8�����doP3#�BI�/���*�qv=*��%&�~���'�����}g��x+�����r˷{�m�k(�ç���r����߽��	����y^f�-��㐼�R�7�"�&~x�d�14)>V]�:�j�W{-/l��Ww�5b[�h��m����ޭr��^sxO&.y�S H/�T�莼J}k̘[��
'��z
�Q���WN�T;���/��
��z�^H�f��y�$�{�@��VT�f�B.Z�`.S��e��"&���x#�3ɤH-�y#н�B�<�����I����	�̓�r�4�=^L\�{d,�-���SH���Z�O�aI|_V�c�H���M +��Bͷ�'�����\ (���>=�������>j=`�vk�5Ծ�~��7Y�+m�����Kya_��$t���Sǣ�ȇ(1��E�����׵��P����q�$��dw��$�Kj��U�|�U��v����,������SyT�Y6Z�y��g (L�@�(��>ء�����H	�p��u�y�*˗9�9������6OgKY̝��j�F�z�wy4������=�O���"*g��<�eB&g��A��]Q�w=z���d����}ԃ0&4~T��W�������n��ң�8����m�y��4�l�o���3Vy����h
U{x���?n�a��m�E�^��
Y���n�Ez>4-�|��p_�L ��C���F��|��:,Tر���꿼D3�;��l���;b��(׳3��	�H��x_�x����u��l���t�K�;�d >(�p�T�V��V�-��Y����(©����), t����?��Q��ؕ���2o��R��";�[@`�dPa�GƮ[��yIӀ�VK,BO���և�9@p�̎�OB �لD�b³oP��(���\�,z`i���B*-}�j.�$W�w�	 �\c�xzw��r��5�֔�FF�-��^K�_d�`�d���N�C�H��ڃ�R���7���J����C6���'�J���'��JM��z�ߤ޾��[��y3h]�ucnOv�Edؾ�& ��Oh��n�2aZ��d4����@N��>yɃ������[��En3���e��|g��6����.mt��Û�,��"�ڪ�3_�f��KN�[t�����l��sT��f]�9�1[�:�:'	a�����`z��I!��
�q��4P�f��9Z����4��<9�����6i�4B�:���@nR?_4����O�u�- ;�R���I�.E�)��Aw�g�;���, �fl�ABFڑ�\~��@0�A�R�D�/�C��m�V	w%1$ڎ���ּݶX�ЫȒ��ߛE��h�gi���b~�v���za�"!DQ��y�+7R�0�lDz�%b��z]�ڴ���a�3�C���.ԉ�.�mV˭�r�s����ye�ш ����Ħ�BD���EV	�U��q�SA�{��Ȳ�k��(⯷bn�#�s��3�+���g�d_�tM�`t�D	�8���}S�#�)�1���H��x���
g��.�W�&>Tˏ���U�Bw�������7�iE�4��~��ſ�ΦX%(��2�4�^���B�3�a��f��k<�Y����I����֭�g���=C}j \�	e/C�)�Kz��-u����#�a;#�-~\��[�N�$�k����R*��x$AՑ
y�0훞@FU ���IHYb���a��!��j3��� ��R���:�6|�U��A��BR)K��O�=�D,l3��������@�h�a��{�$�$e]'�zW+���1���!�SKNE����}A�N5f��`���J����7Nr\?�3(�Ž���>XR4�^6��p���C�`f�(�V�qv�ih���'��A :��o�!>�MU%�+�{��%�Ҩ��)@	��}���r�&�̟�}��ͰO8H���ԉ�jH�ض�h.�Vv��������2t�!�RZ`�rl�.Q1m=O.P�e�|CGh��b�ѿ6�P�
Ǆ  ��哼 ��,"���U�� ������̭<rb�pMܦ׍7*m�L[}�����BJcg�6��*����?P�E2�S;��Ci��j���_�\ �?-�O�};��hC���U�fU9�:�r89�����������{���u�
^�z��N������L_}2������HvlWuYd)�#A�F�q�6�G`�)~�U`�1��ǀ�LHK�>y	��F��NM:�n������0>�4CS�.~��~�N�S��PP�c� ��(#,�צ�k�o�C����Y`�g��r:�s^�~[x�>߼��%���d�l~ɞX��(��>���9[<�IO�eN�8X��!�P/��x{���J@��H�0�>��:��m&��ɴU�9d�)�G��u��ө'9�ڬ��x���=Lw�����n���=/�GPAC���N�^=���xO��i���Y�݉1�:홼Eq,#��,B� Cua{�Bt�_<Y���A�e�g�_�YW?G̤I%`dD����z�>���h�N��@,y���x�9޻���R.¡0���@0�_�IgQ�H��s�vs�Ʈ��|�&=׺!P(���������&�-�������F{I۸�YL��j�I��^4X�������M��
��s`��ɇ3s0�zR&p�tvd�Y����@��
�e��ݫ$�W��7T2��2��S�%O��4�XJ�?�S�������F�]�������x��2�D�j�.��i�Iҏ{��|`vv����e������̾�j�p���u��^�%�\�Ni|vיU<�S�I�ᘀw�O�) ��o���I�ճ������J+��ќg�����C|������)�]���f��Y1a���"~e��IS�B䵃3-�84�1]G(�1�=��Ƹ�TH5J�t��U��{�l�V�sD�Ü#��B<�B���"D���s�|	���07zz�`���>����6"��5�|��n"�d�<�o��I�ʘG�8b�Ӧ���U7wc�=GRdš�:V��u�#5x!Rn%�Ȁ8�.g�����Ǣ�2p��F3^d��SX�������+��=Կ�;(��75cw+�EU��o�7���`ɍ�=�����l"9#,��O]\�ǒ���/YX�F��b��x,����7��E�.Edt�#��OM��X�^�»՞�ܔ�K���� s�2I�2��"���OH�[ֆ"�5�3�d_���6"���¤~��HA�B�ֳ���"�W�!�=�޹s/"H��ٷ�e���Na��<[�=1KM�v�H��������I�[�O�b�#'l`�����B�^�!-o��1�1��ʯ	,q���=�5E#��m��"Ǒ]{�M��pq��)��H�U�0��X�J������'� ��7�9���ʾ�dc���.���m��օ���r��S�NسI�;Sk���@���b��<�Qjq��L]�P%�`fG[�.m��P9�o+F�q\�_�uh|rp�-���iY��O<�qi�(V5��a�E7��D/̸�/�����/�h�sX�A�z�;a^��h�
g��21�R:њ*z���v�ı��=�"����ȹ��ǩѬo��nH��a�D��	�@A:̇�Ԃ'͟���,��A(�0��g0��Rx���-����B����w�J� '>�(C�D�����G�C�[��a�e���t!���?�A�+� ��ZA��M��e�R�7'$.2c��5[��&��>�����<cG������Ճ%YG����\Q8�.�ݰ��mf��:��~�S��x��])<�j۫��z+�l�I����j1ӱV�Ö*	��n�GZtN��C}ʓ�2x�g�S��#O��H1^���Z�jB($nO�Lk�`�u��qD��-�d>z/�EA�eS�n4�d�Ia�T��o�K�oHHa=;��,M�#;!�\�6��"�a�t<�_}#E�8�������ä����o�UO���ܢ�'�_���[81���l��E������O�X5�ީ�ؗ݋��6���h#�l��'�S���=�V%RV����Y�hvyϥ�S�5ӻ�*XX{���T��f=�	���5��x�C���W��uVu=m�3��	L��ЪQ&)��/���R���\���yϛ.���Q ��z�$/+�g��n=�mF��o߫��ڛF�ֺ��F�h��K�M�~��<u����I�h���%�P�N��YB������<^�߶'�)���N�(�TK~WA�x�<��*Y8���>�[���.w/��*^��[y���Q�z�b�X�E,�j�I)��4��rq<���/T? �h��H�0�kҼ&��8�x@Y����U7��5{���GjF��B��t�����+oR��P-M���3w�ys�3������덎�_~L���p5�K@�<�&\�Q���ł
:ֽGk
��ɕH���r�[Z���H��~SZd������惴 7Օ�Ȇ��*�A��={V�w��r�����ݎ�L�Gy�JYn֮�]bT@���f���v.N�F+�ϕCO#)%�{$����,iT��7���o�
�jԈ�D[�
I�}[#s9l,7�\-��
6D~b���ܒ��d������lT��������"aq��)�ij���tH����+�K��|�l`dB�R�|�Z��*�g="l1\"���%�	Һ�M����^g�<L�7���q��7`YC0l2B�Pwx>�����Mkb����R���u@�U�է�T��E�A�=@�t�5(H�ʚл Mڊ
��f�.�$C�
�;�ު�Ek�y�Qh�q7�L���r�"��5�S:6<~���kff\�;��D��$��4hG�&B��l�X��9>���u!�*=����t���W$�U�lϿuU�E�,l�\�d��MkFRn�@�vp���ʽt�Qɝ�{�����P;�{���Z�^�	@h������%%����ln0o�U�	��`!�0r�Jԃ�r'�Z����J
x��v܋�[�A���<�2_�|V�R�V:Ŕ/�k��%��aVZ!������C��� %��1-��R*�w�=�e�z�9dfg���L@0�� =���
����@��Kc���#ڈybg\n�@�1�{��[�=�\LC�P�e���k�ܬxG���������M�кW/�v�����~?X�P��cWILaV5�=�Z�����?��Tu�,J�p��,�lM��]���ĕ���W��c#�0Ԡ���]�!��f�  x� ��i{y�ڑ��"^���=]k���ӻ2Y�艌�,�������N�ء�nuU_��m�
*|H+�/����ͩf�	��,4IH�~2T����*!��^��^�>Y�����Ä�7*�6�Q����b�.V$U���	��E��A+��6�--d� ��z�[m����4��_<�@�K�� $z�A`�����S�SBxp� �OS5ƙ:��_�J�V31��r?/�P��[��Mq���<������>5�ϡK�S�i�am��R��M8�9E�������3ǪQW���Ǯ��g�̈���i���H���,�:�������>R؅It��fH�tyQ�t��v���vw����$��c5�������Y�T���o�a��x*��j�&6t��QWf(U;���%5:�t����`G�h���MM��f�_�|�{��A���>Ȅ���#�k���ٱ���Q�$�R/#c8�0A��=�IE1�s|��|؞�*�y&�z9?@~!��v��y�Gg�L<�J1�n���`0�{��JD�|�P����:ԫDSoHg����7��ize�G��署Í��bu��=XA#��PI=�k��D_�D��f�u�7E+���m7��\Ǹ�
`���M�d�vO��T穋�q ����D���N�z��Ƿn��
�Z��Y��s �d�\��]��|la�1_�?{�E��X$2�0��օ�!A7�������P�l�(a<�=b�9C��
�B����v�(�h�-�
sP��.BSw�
R�s|tE&��c'���8x��>�\U��k����bjVۉ���>l밐R����J��AT�Vk��}�����^t�:�4�R!D�A��h�^�fA~e,·s��f�+���?�:�ޔ��-гlB�����$Mx`\_6�V���Hh,m�R#��uo������2%*m���v������F�����!��O��fEh���z=��Kd���ƛ���p6�}�%�D��n�ް��fq4-�Tg�w�M�����O��kA���֎$Z��5�\g1<{nF	=FSxY�:Ut�%�o�4����=R(������Px1}xo�m�K4��r���e� �B��i���Yx-�q�w��S��bQL� ��V��������"��r��]0�p��Yq.�����r���m�H��{¦&����3n�|�!m\&�2zV�%ok�S��w�x׸�hNIS==!�@yآ�8����[AU��Re��-9G���W�Y��R� �	��Z�� ��H�+�8�jݫ�!y����~�yO׳vs�8�e$�?��\��B�h�k��H;2��r6�n[�$8̒���{�4�wdi�C��eq�,jxJ���O\��Ʈ?A��������r]�h>E>"\�1+�$Y#h��@@�ڕ"�i%?��/�>�;)1,eO���D�y�:Bi�F��\'�O�w�7d��S"��hx��g����~k�!d^z!�)����`t쫒��9	2�H�U�N;߷��@q�G���߄&�.1�kl�[�U0o �� ��b�{���IW䌼�]����c�� � i�a�"tw�/v��"�$�mqh�Ͽ�t�hs���WO�F��O������X�,���ǃKq�חi�fz��B��!&�f?v�����p�r�,�ł����4]D=�F p�T7��ȵ!�i�~�s���$vH�UX��j����21������>�*��rB~L�����O���CL�Ŵ��'�?DKwԶ��d���g��L�*i�ֻ��j��B��@E��g���ovD���y�X��{]�x�^�,�6fj�D}s�#�
���*s�ڭ��g) ��۫
!j{E8�h�+�v@�q!<g��_Æ�5YW���v�<�(q,ԅ�
\I�lc�nN�0.����{�6=�TA�᧐�6��ɼ�ȗ+��[�`i���&U*h��*�"
�h���:]-����7S�.1$�H�G$$B�-�n\��<��sj�X9�+��w�lM��ˈaơA�p-�s7ǟ��*�|�M0P���e��(���0�����=�r����c����+ZL�)?��#�����3&�E@l��^_(�70�/���pD��G{o.��oe��`O����'�A�o}�Wb��#���h��oBV�M�J#1��'z����F��"�a�ľ.,>�)CR�P\�~h�� ��zAT_"��w�h��6I����ù�V>��"R.���(Tl��a�����|kx�x
vRW5�:j*�`d��b�,�2^A����sj���*l�DGت���ژ�jOn:l|�,>;��1�B�~�E*In�&�R�h�>��4�٪qnvMʎA�/q�E��o�3�AE{���L<��/	���Dm�?xb-7�L<�i:�pp�������M��]�4k@	��NQ�G3����uO�?�h���e����]v��A-t�|5k�[�G����^�g������-��Ks�rd<��#-��� ��V�}N�(�~���;�ф
�e���"5�4��7��z|��{�)��?q��ćͣU	��@��5�m�Ԁb$լ� m��xS�)y_�p쟷+�k��p�-ܲ[�<�=������O����`�3)%1_?_g��I��C�P�ګ"c\ѐ���gz��g�c-�5}����Cj��-ߪV�����_�o\.����sȘ���ٕc������!8)�r@�]�� ,�j����a��L6�+K�[#H%�G31T���A���m@&EU��u}^FP[(���dG��Y_Տr�&��`<�I>/�q���O>\s�4~^gU/�GO���MfH��i�:���Zx|a�w��Y`�X�rjy�Wﻃ�	I�>�VI6e��l���Y�U9ED���uo�cC��`�ø����l5���˅|R�f|7
ȟ�᥈���qM]��ɠ�m�&N�veҠ֧N��
�S
��U��n&20g+��D���,{<;j���'ߵ�mw X��}��.�O�r�f�3htWq��½8;���r�p2]\,4�qA�oI����ݦ!m� �ޤ ��3�2��w+�(���(v���p��������O�$��UJ� %�t����J;L�=��e�PN%Cj4˘3��P�����dc�E�Z���/�H��҆����<z%�,���B��k8A^�%�&��+�n�1����p,g`��'��5�1gpyB��Z����S&A��w
Ⱎ��'��>����pTJm����I'�'��_�Ek"�0�F����^��}+9�0�8����^T_ޭH[��Y\O�����cͭ ���e!�D2H�
��Od�kv8n�~��iؠ�����:i(��왨b8�ᶣ,V��)&>}"�R�kI���ߢ��x���#+��n��a��z�f��^2�k=����/����S��s�c�l��t�]u2R0��:3RÐ3�i��:%�6�|e�uW�[<��m��<x��Ȩ��V7�R��\�P�FP�wOs+�r2���+K4�=m��(���F^������dx��g
6G��Ͼw�Q
jֻ �~2w�]Pn?���f()���іm`��u[<�|�"�C��!@.k���&Bpܺ���Yt�ءo�MMJЏ��
*�	i	�A�&����8�8E_����U4����}�&�4�NէL�s�-v���(Rf�T�����F��U�^#7_D��
�xsn���6�:�$��| �����[��&3�!qY��Cxq"(ףɆ5s\u7j��5����`~��S�5p�
���]���[�1E'+l߸`5U�P�_,::L'J5���G�n��DJ\[ h�?��
��)�
���'j]�c�}�Ͷ��;���^��A�\]�{����Hi�e:�;;e���K^�2�_����B/����Q7����edE4�M����0�&�K������R��r�G���ʑK)�7>^�[Z��t�s�E�袏��S���>��|!!~��m.���:\���Į�,ãNA���y�т�vW'�r�k*�*�4�e�!q��᜕�/�m��C��g�*_������*�1�H}R��&Ikr�kg*���G��ݗ.�.Ǝ�̳�����g�+Ia�p�����0�CJ�Oe�ȕ$�}w��d�9\�qd^D�����f�]�;��s+���D7�̋;�2zp�)�q)�	>�pq�?Q=hyҭ ���[�� �j��H������-4�E�7���h�X�����g]Gu�a�t=������N����R-	]e�B� ��hl��( ��:�d�h�a���B��V�y���~�i������݄w�}\��ݏ0Nْ��&��Vk6���j���M�;ܐ�7a�h���t��d�c�a�ȍ���.ބD�gH	w=�Kx��<��M���C2E��������e�x��o��~�oʓ��1�?e�dƻٿ$]��S�U��Nڴ���F#�ep�;�	��YE8c=8���1>����~L���IS�-�XR�ɫ"�ͅ>��.�Y��6�%� �k�l���Ġ6�5Kq� 3����ڣ�T<!��2Y��)	.=�LT��G��w6� �=Xw֡�%O<�jt�a���7M�$� ��k�'r��Y%���,R?�չQ��n��p|�os�/��M�w�"�i�}=��ٱޞa��L�+������:��/��x��<�
e�����`��-G�6�nI���w)s4��}��t݄x�d`�7�7z�
�9��s�J�F������E�+/�|0p���`���e��r1�}妷�M2���L�0x�3��$���#�
dƏu���{mX��G�B��1|�]Z,��ct_R���� yr�o���wj�B��V�5౨�B����b�S�梯Ԛ5ϓ)Xޤ�=�PI�6�&�1��Q@d7�a�7'��b�.�^*�V�O��:Q�����m�&KP��C��G��̀>O�.�������Rvr��F"|S�Q��c_��AXD[`���T�b���\���v
�M�j�ޤ��R��]S�����
B˄o��?):�Lf��k=�F��Cꕋ��f�޾�k0�����M/ Y�Ϊ!����YܔG�=���i:�j���4eg}�.^n�\�B�Hh:��V��R���f*`�s����ѧ(eei�Pg+�g�!?%�y<V�oL害Bʏ�������X�>�U$sn�F:U��1�G�xֶb-Na�(L��/K�ms2�@4��2�{��L��~�x	�1tӐ��B5P��.f�c��@	���ʷ1�0M�ʠ���� ũ��<��	=V}ϤV�33ܸ�#g�zp��N^�Q!�_�*?w�LH���Z�پ��Y[y;�G�JW�#r��3Q���hD��GU�:���;�^b�V�}��)� �J�A�ߺ��2H�j^G�?z'�n	��j{�lg�~�7*6_6�t'e�0����j�b���tl�_&A��6�ȋ���Ep��� M��I-H�,p55��x�;�%��~* 5 )DE��h�k���� �R%�Yk�2*}��0�ZR�J�5��;23b���{L�$d�#��,�r�4��xOk!��'�@�M4��@�>�I8�E�S�N�W@w8�	#=�2��)�rn��M�Bc6���b��@��vg�eJ��s�W8�@n!xR�A`1��}�s���c�]j,_��|���M��prЬx��,�V�kV��:z"D`�Ohh�AwD��d����q���55}�n�8��ǘ�<O�?�2&��ER~�%âHx'\�!�d��`��M��H@h�f�d[a"@���b�2n��uų�x-e!	�����V<�o�5��إ<&������'H��H����e�1r+� ��]�lye�

+ ��`��(#ڭ��h��faٽP���*d?nr���Q��A��6)�-��+c�F7U���zE����*.Ez�OZ�9AԞ�f�#�
w 5	[���s�8HԳS��d�#�5�M��
�  D�uwb��)�@�||���`t�LJ�n��8S�>6(?���
�N���UTF�%Ş^�kU5��!i��AE��2�7M:��\�h�k��\?A�59M�3�y;K�x
��%Q�8LVX�6�f��"�
������(�%]g�
x���}�/��~���{h_�i���
4��/���Жe(��5����˸5����S��:��"�4Ou�V���F�m��[�n$��8� Q]��w/Ӌ�:��8�N��x]Rï��Rp]���G�I�Hd���6s���l�h�rYa?5:1��6�!]�K���C��n��.X����_�Og)[��sA˰C��V���m	a~#��R�Cf p���i�*N���^L0�	�-�ᶺ1%Pr��$�As�خ�ɯ�5�l�PKE��oR����v4��+�Yvł�Ͽ�)%�p�N���:D���qK@c �l��o��3�K�"��f�{`�i#�2�1AWI���ʦѸ���6�W��b�Q��6�0mf:h�x;��t>Ӟ����CFV�'�T:,�{��4b���9{�[(��v`����(\��a�nq��!&�p�6홽A�]�P��	��s@�)\�'������>�c&���ذ���fJ�����t�)$�Fi�v`�ρ�@��]"y�����z`(�dZ�ӈ�.ˆy7�8�v�+��:bf�> ��-��L;��'
���o����52�]���[�1J���N;���0�z�S��Y��I�]�ѓQ�:U�}�֞;����h��O�X�:�G;�v���>���(}��z*
 ���	*(X������iM�
�"��r�㢅Ѯ��TM�o�2���լ����wn���E�)�������N{�遲���a/��z���SVf4��r��ӯhx�h�����!�]��Ry�w�_�Z�y"$Q y6w���#��C4�T�S$\������y�;�BC�$�<��P9�����$8��$��V)J�ī�ʏ%hm-ʴ��Ac	댫�>}	�B���vT[���ܚHN�ef�eM�L�85���8�+ �"QNn��H�����4\�]��!�x�
��|�؊1mB{�m~G��"X��+o�0�������^U�n{��$�H;BvSC�8:hʞ��Z�JN�T�b�N�T�9�9+�1�"�m���/�
�9d3�k�m���4���(,j��f݊�>X�#�� �-w��ю���H��U��,&$��ܕP�����<y��	Q�I(p���$��u]�+���B�����R��)B��h�GV���A�h����	cXE�64�X����/�ΒQ���&N;5��r�B�jM�ۢ)מ)>��dz�?��ɇG��P$�&'0�v�7��4Gi�Ń�ޡP�qOV�<O[<6�w���9�������0WA��U,:�p���B7�u�7��+����$��C�k*V���)���o`$Fn��-�	�x�we�&ĬHR��¸/x�,aCmG��̏%的�rց���b����<���Y�Ϫ�/��9�*�~ ���C��q���i��0�ߎ��74&�N\��mb�p��<��B��q��������do"s�[�L�ᔜ��@��\S��.�\g�w��=�t��UaU��X�W�����6�@)᜻�B	�C����s�����|���D�ش�����4����NV���.��;4����Q��i�+5BG
C�%v�/p;��~�w���0:�ĲZ���'/���iWk��H� FI���p��1��lh(oWÉH�YN�$C1b��겙�갿�偙h�>"> ���'[Zi�#��ԫ��7K��x4S�*�$�R��Ck��ϛ-	9Avh���lP���a�W�\�Y��J]������~s�7�^-�|�%����EY��%�'�$������h�^�n� <u>Ȓa\�k	�U	A�H�_w�5�I��f�@td.�-��5N��u�Z̀!N�� ��S�R�=�	[rW��D��+�O��@�7��9t���� �X�!������˞�8@�#��??�`,UC��%��B��Wڸy�1���q�+p�b�&�XjCX	���x@<�����&�E��jk)H��l5��'���v��"U~rOB9L3	��}��:b4�?�%�T7!:e@�HI�U41\2��M�'at\&��ɑ}�� Ad3��E���]��*�4J�Q��>I���q8#��5�ge�g�{�P	�(t���E$1�l���X�b����KZ�2r2������ ��j��<�ß�/QJ1(n6��d�aB���&t�Ծ��.}L�_	Q��qL!*�^��,�߭/�� :��S�bB)�T��
xU&'���M\�Q��ǯ[V��k����6/�U$X*�Zr=��ۆ����8����[X�j^����@6���h�4 Ŝ��:b��B� &i��t��0_�=� ��3x[��s0w�?�x�f&<����b����.�yx|-�{�L=�3�]u�Bv1���k4oy�D��=�mȮ��"��>(Ko�W����-�i���Op������޹s3�[��a'�e�-+��">( �4N��m���`ѷ�~"h�P먴dɑ��P��k�0hC�4�V�1 �Z�]��:��(ZJf�ܿNy�N3GB����p�y�J�r6��"�	_��{X��F'\��Lw�N'������&��oB�%uOb�4�w�C��ͭ�}�e��?2�y�� `�c���@aQ`�h<�x��ƣ��GJjx�%4�_p����]���*iNJ�ܽ�6�V���_lk���dH�UG�-�O�����d�Q�ۃ����^B���y�q��
���E&����[2@?��N(�jI�����C������>#~md�������*��L�K{��l��#���yT�����-
�>��ݺ���HN_���%jU��-��S�����%�b����6zI/2�jp�D%������^�þy�6�Ń���7��1�4�y�dE`�t��P��f�Q/����\M����0'Q�,������h�|����_���;*k��-�s�{�{ORЈ%��;�G��1ۋ�� ����I��մ�i�p_�����(�! �уo�v�t����	(q��D���9�x'�ZsG���A!��	�[�͇�-8��1��<z�S�z��^-g�����Ԓ��0b?�?߆��a��}�z�l�?����˖��o���Fe�b<���I'��![g�`����&�ǻ�k�=��9ŉ���8˙Xx7�U>b���5[�~WD��1	�Y����Dc�e��2>Q�Hom���7|o�q�&�u��}o P����^蒐�����@���`�fAZð�ӓ�
�X�u%���68��F�)E�;]��
X�-�m*�e�M��$|
.%	G�g�oc`?���&��>�"�g���w)
pB�̡1���_OR�-޲@%�O�����&�� ւ~�p�Zh�`���e�/�ƙ���$��r��	�7IdC�ci넧��Lh����,��z�3�'������5�G��j7�aڍ�T� ���%�Ǳ^�j��ra x��«��/��1��1;PƌT����C�I�.��W{���%؋��S�
�h���K�e�_$`������j�1%E�/��}�Y��uf�,���n�u�3N�}�G��bE�l��#T}��$��@l�D.��\��%��%����IʨCL�q�,�[6�U�<�g����E���ٜ�P�P���.r?���3�M:��� ���]A���_NB[hq)�ר5U��{eT��Vs�	B��;+t�֞o��4u������[5P��9�5���Ɯ��J�l��V� ��2�8p�=C�M#c����b�����Ǧ]��\��p�@��+�ƴbܯ�e�9 ���|��6��}rV�5x���n�9�����n����vV�<-?0���q�`��c�D������D���X�e^^��C5t('���,w�j�YA���"1�a�K��������Mf��~�%3��kH�.C'JzS�ĵ��Ԭg2=�8إ�OA� _�]u�>���@Ɯy�;����c�eP���s��
��@�Ҥ�%�g��#�L�v��g��Z	N$�P~��N���	���rBNj�|b�=��9��hP���ǹ�,�J�5�De����UJs����k��{���p"�Ѽ([��7%>`�"̈́�eF�-�m|;�战�a5(�L���4�q�e��^�+1g���=>��`�����/j��j�rU�G�z)j(S
�O� �dk�T��JI7 ���D�����G��QU��c���(���|��ɉ���Dc{��;��I� �A8���ʿ`=�����>$%���E�G�L�@�s���j��kwBV�e"�>Y�LX�h@ph�p��h]JZ��@�?ՏbK��I�U&J8᎒nK���zeY�GB�0�X쫃d�j\����D�����c���*)m�Ӛ�����.s�QE݃��P&X����%�w�B��]�[�Ce�5×7�\�-m
=�!��4�>\�+ n� ��@Z �_�	w)T
ė�}������Z����g�WS�KT��!���S
���&2
e�&r�%�B9��Zږ�A�uoi�p�H$?e�I���VKL��}��^��wl�HQՊ�}覥��NT�@ae5�J��Ø�����'�\3P��s�Гݍ�!(�)�c�a��r�lՉU�SL	�\Q�
�F�y��
���u�Ő�H+�$�|���՗QOJ���m�����Qѹ�5�X��9��m�P����ՂZy�Ϣ6��պ��2`M�ǔe��N�:?��Ul]p#KL�<�� "/�u���Sk:�Ƶ��˹W�������V*����v[ُ�6�ɻG�eZr[q���&�, �ԟ��U���O��HP���9����K> k�N�V��b�	������k�3w�����f�`�:� �F��)������c3�'��0ztbVջ�L*�)?v k;$��|[!� 1;��1�?��%�}^���C��W��s�b�m��T�l�g��*;\����F�?En����A�_u�`���QůDT�^�Vu��%���(յ���"p^�g �;��"Vm���Z�*��r��;���6�D]�Q^pUE��<�u��cy0)/c��^�_�>s�Z ������4�ojWf=����d��֫X�We���3�k/V�6�X�����`�Q�x:tM��[�IX�������H��t�{�^�:�J�$��n��c@N��Swm%k�l�4JPF��tP���z�̊T�H^71�W ���͗X��ӓ+����Wк|8H:%�l"��z4��/�8"����]���E��{���U�{�7e��q-d�_��3�W�+���j鹛{hBƈt�od����B�#ǽ��b����Q�D2�1�祅U����c�'�;/J5~��y5=��^�k�8��O�x1���2�KT��V	١�gKcfIj|L�eĕ�(�ث2�ڌ����=5�V<Ÿ��c��B���(#�҄��ݪ�c=�)�.��ԯ�V�@$͋��㡻�T@Lq��?i��@|�)�w������ ���Ãua� �?#؇\y�������h`��ߡw%�=����&ó|�+<ӻ�zg���c�JD�M<!;|�\�_����1�? ��2ֿub�o��� J<(�$��~��9(������D1I�z��(4��m��¶?T�A�=�x�
�M[�r�� �b�!�Fh-�#��f]�
˦��J/��͈=��,P�"�(]rs��{�>N�a?�W�6mn�.��6XOX�G"��xL���SB��ӻk�maC׭"+��%<��#?����cƨHz�j��;�41t��C3�VG�Ob&�'��/�H\���D�x<��
V�ʓ���V	�>��CReS�G>�`h��s��	Y��*�G�wj�MT ����>��Q�Q�u▲�O_��Y%��m�����L�U���ˬ��s��9%Ƈ_<^��Z�X�)�+0�!"�6�8���(��\�a�ZJ��i,� S�@a�:lc�H�0X�u����J��@�g�\:(��òP�h��8�5�_�JT�}�/_(����X��d�7C
c3����CC�KE�R�x��(Z�0Ai��*wT�/A�S���uj-�iF4�?Ź�(0��U�#��mZ���/	ť�429�/���ނ�'ZW�/�[B���z��b�Bs���9�it�=����w���H�*z���[��(�ԙ~�{��O\�(h�{>`Y�p�^��BY�����p�7dKĐ�����ӞC���� �1H�˷w�1,T��K�e�㵟���������6��T��qİ+�^.�%�ʛ%�k�:Z��ɸ��zg�sյ}{cw���~���s�m��4V ��n�3̪H�5x#y�y�'^crJ�����}!ߑ�՛���a����Abr�V�����;�/���q�0��La6Le�,Ű�S�
L$"�XN�ӿ:��v�.�BIqv?��%ٽ���I�W�,�~�X���*�+���s�#�ɳ���G���lQ��@~)����1��&_'��hY+� ��&�Z]���s��I�?Ao	��^���5{�U�yR��n��~A��/xm'��$�Y��1��`��!��),�g�@�ؤ#{:�^�,u�У��)J�\��?A H1`��)G�]�o��"�\�_칱ν���Gm���	=x|
����f�-�I�_�1x����yw0�ӌ>S �6�F�ܱF�T�m���uw
Zc�F��ۍ�Ɲ�D	*��J6��b�p�&_�S�1 塮�s��-��9����$<}4�1�J��4�Q�	�f���4���n2�))8B�Rėů�� ]���ɯkR��~� ڋ�}Tп,�pZV�ŗ/�`����h��,L�~��?��fj<����n�4��}S�ZN�䷟�_�H�O4Gs��d�Q�	��%�y):���{����r�{��z���do ��ښCVA'�C�D���y�&}�䱧<_*�i&cl�����x>����L�7����N���Y~X�b�K���Qɔ��?jSd\�D�Y�E���_k{�Q���a�� �rIK�v��A��F���	�B��
^�	��IM�cLG_��°2�g'�W&��v�Q�.gP�XD��� #UV	���!�u_Y����R�����&Ɍ(��yj���Ic����ȦO�m�^`$� X��`'Ƀۡ�nɭ�J�I�ݏ��4&�$L��̺�x�t�T"�V�OP�Þ��ƾ�#>�� v�k��=/[}�{�o�����lr/�~���H�8��槪�x�͹�Ο�)�Dj�4P�ƌ�$�%IХ�gҨ�\���D��9\����m�ʻ����?�ѐN���%��9��ڴa���:W4v�ʲ���}��8�1��'�t~6������i��,h��^�"F� 57����%Q�T������>�=�e"�������n{)��T�}T�&fD�b3|П�3�}��cpjĒ���1�S�x���f'�u�� �N�|R����ȈMs'��ԅysY�4z��y�����0�3-S�T����l��>�Qg��s�V��g��5}��xu0��V���sE���˿C��C�K�)`P���٤�A'�Կ^
RŇ�=DA�\�1�w�˔ǎ�:	�}S���O�L�k��G�&-��n��}�STcw`�_�pr���k��|�� !��6\�B%��x���9��"�A���+�4�W?��x���������n��M��yOC�t��ku3Q
���?Q�C�+�ǭ_H��s��}��4��՚Q��k2�Ɔu%2�'���F���Q�Bg�#C�wꆔ}����y��ڊ�trd�V�V�H�*޾�mL�x�?E�^���s҇I��;?��	��S�+HX7L��Op�e�J�\��bV�~!B�?$nQ!6�+�\τ4��~�y+1��%����*�^�T)k�s'���j5�Ϩ��=�P*v�ϡ�@Îm��H´��n�,~�X�&R�᣾�BR|P�rQ|��1�'|j��Xx#�r�����U/�ϼ3c|텆��A�RЄ�nVm�㥺~�ТZ4�(�����ͫ��6�`=������A�l2�[��l�f �@V�iu��4�K�IQr	�pР�+\�K�X�Z;�q��F ��%=PEoE%�ծ|û�1�¢�>�T���5�2�jG�D㼳����=BFZT��M ƍ�N���ą���(�1���Q$�,W-��'�M�:o*���XP"KV�nE��g�a�d�)��}�A6Os<��#�P=f��/��.��	�G�6l��z^,[��:c�G��U0��Сi��we~��R���sn��BQS�#�"�z�%��r�����}��>�Er=O���Ǌd��ZɕNq�3I`����0�v}&��p^ڐG�3ǜ�jɣa�׶x��  ��iD2�|��/�1�̃y~�J���Ǧц2g���<�mm��8D�3/<�㽦��F8�ӣ'v3�ԽX��������L�9s<dT"<�jqu�+�D�'2"��M��	���$��~2
��K�+�x��Jl����	ή�^I�M%���wFd�>]z��ԛ�e�y��=���,��(z*68x���v����7�m�e��?���xY���?.{� 7�f/§���63*�:��'���%B��5Fz�4��f���)��6B8P��I"�%�ȭ#�ǷDD�|KAq��gދ��j��PH.�H�:�������xw��@���6��BwA�j�ȱ�B5�ټ�B�nuj��f,�#��#*��� �`����]�VG*���L7x3��2iKiv�_"��s��0<�+�k�p��+��a�Wo/�6����,0O�|o>�Bj���uq뱹�z��c�r��y��)'4�#�S?Y~�Ƨ�Z��s���Q���l����m�O](��d�>�0�G���1=�?�:9�_���t䳗�?I!�z�(�t<�=ֳ~�\Ƥ�6�)bb��_��O��7K,2��vz�36g��6��d���U�� ��z�y(�CU�W���
jpr�6���c��b&0��Y+��3=��X�%�0� f�Xew@b��*�yގ����uX�٩�[1Šn.����ĺ�v�w�Q�{�so��,�;JP/7#��<L�"��-~� �1=m�+�5���S���s����}j��w6XIU7�6ӏn^����*�y��8#��h=�S�I![�B�,kv�OYl���2�o4��C�<'d�"S����s�$]n���lA�����0� ���2o�,)�B\��� 2&��4�������9����;\� K��u8y���ɬ�z�����,%��������RX�<{�;��h�U�~�
�@`�5��X�Tc]����;:�-����%���E��i4l��+�V�)����W�R���P��m��)�r݊O��LcC������ޕ"!�o��2��G�����1%��l=HE���$��Mֽ�
C_�����[z�KNK����a�I $���?c��vw=Q*K��j��u~�"�wS:W��y���c��nw+t��|�Mi)�a�fh�&��4b?�Ӓ�諾��ty��$�D���=���ߠg��g�h��)����ΐ;B�r>G���T�}��8z���'��à�4��Y����-�+*�l�k1��s�Ճ�(\g�B��Qp�
��G�|�2c?D	>���k��xR���8N1��O� <�G_�ΕF����%���i�Gfi7�l~���p�·�z�%�H�z��ϕQ���뮽�O{���2޸Kw��|e�M5�q��Z�Y����37�BD�$w�^�c5�:&�k�m=�� ��\*mi��|�e�	ވ��8�k���\��g�*��I��ps"���1tE>��%�),��fxl��W��	]m+�~o��k	,�������	��n=>�{i��#���b�y(���i@�H�	�w|o�ڸY�x���e��]�mLЦ��Ȭh�tFo�b�%?Q��D�C �V&����ys��>�Q��x�cv :����r%<��T��lD��0[���U9�(2��@�`-I�����nA�t㷅�[�S I��Zz~�c�J�]Ŝ6x@xm�>�`QM���bN��g�tV��ko._j�R�%�����F�/ˈܴd���<|�ċ���ݔ�*�.�������v����&Xc�BR�T>��/8Tr�>��i,,�l5�Z��r))$;>�;����[B=vӋ���<��_����<Ps��D���줙�!���e�*ќ/��Ϣ�?!odXB&�2��g��Ph	���S��Wdu)g�^i�n�����ι۸|��N��$q�𑹗@$��\�lG�G���N��E@�܇�U(��Q8�����2��;��A ͚�!O�|���;<j���b��V:�M8�����%��pĦ�S�b�V�H[Y����Đ:L�XtIg��VÒ��%9� ׆��TKZ�+즰8�"�Ov��y�7iXhr��4"��Lǚ��)��W_|h+c膂(�Lt*�o���yȄI���Ʒ�����
��س]T��X�1a�s�b�O��To�?w۟���"⅛z�+�ݬsC����|�r�h[���H,5���ٷ��R��1%:�P\��F��v�W
�l�7HFmv~��_���.e5�[�qi��U���2��Zq�u̖��֑D- �V��?t)�Ǫ�`o��d��L�	�=��*��e
��\�d���U��yn�T�@j9��#�,���������l����^|i����?6�5F�n��4,�93������G�:Yǘ
j�|EHS��O�ܞo�ڬ��e���X��l
^�cVA=��%{�����pܦ�����M5ק��De�˲��������>�"R!RPO���+ŒPfk$& ��aj�̒-H�i��Ԍv��d�O����I@�	�����B�����E+?���+�ATɉ?D�AL����Ţ�e��%g�|8Q� ����d�=e�ê�Z�o��m]�$�$V%aq�U[u,�&?�tZ���'��spm|:-FJEq1z����-0�y���*z�a�z���N���'J�$
�q쀼��<E��[U���埱��O��TbN��8�� ]e��=�p���CĊG��s�|[m�8Lq�
T�dZ�����Su��cgz?���>�Ϳ#��D`�WL
aC�%	yI�Ԋ�У�k%��-��]y'��&��o�i�Z���TN�2|�(��h�6�Ş'�o���;�K�� ��W�9-	xlw����*i{p�r�T�u���"�fmuǏU�|��y�q�.�`��\P�I@;��N��P�Yf��2�6q�6�`X��*E	�uoR�u��@4����UE|�Q�@�}o���"����J��Wi��H�D"�h"�&U5��B�=�g�z� �D�(���7��5�-�� �g}��3��W[��)��d73^�l�2��6س/�zI <����c����U�!�M�T��CB�kB�p��+�6�#�">B��nj���g&���N�����}�J��@˄=�Z�CJQ`�� ?��,Y����U�B�N{?��"d�{�J�OfIN����ߌ]G�!sW�%�<oB-�"�Q��P���/Jw:J�zo��dk�S?
RTTd5s&;Ý��+����ғ��q�ɡ�����8�2�O2M��	l�ጩG"I�P��e'���r#�Ao�܊����mTÚI��}���P0���L#�tE������� �[��Ƭ�Tt��2�`C=�Y^F��cz��3#���xxNe��k%�� ��:6�R�����E��J?�*%��Ж�w%�`�nM��&�U�񞪶���	���GF���tD�S��"�|�I�}�2�a�-(���/3���.V�C�+��\�>V�6��R.yP��(��#��D�(0_3��G�2ڏ�=QX���X�����1��)0"H{�X�[��hY��L�'����s�W�P����};�܍p8� C$Z�/��I����-�a��n�T	H	j��;�-�T���&�R���>�K�Ӎ�o��ld������X!�O� -�_�����8��l�L�SpXSL���DK�{�����Ag.�O��d|���3����������X�ĉ�8��d�Jr����tsF�;0cY�.D�/��0���Z�q~5�[�T*�QPJ�@�0����nm0�Ow%8�O�����%��i��5/ڄ�����e��S_��l��ǿ!8�M6,u�6ڶ�h��Y A��5���u���{���	�/
�V� T�:f�柤:��R��u�&$y׋�3lU�	�s�R	���\�5S��+o�.�Gw}��~i̜�.�e���H��4�g+d�� _�f��/��28͂����e�5(��MҺ��Dtl��e�o�{�f�.U~/r\f��>e��1w,��_� �V\s��ŋ��&�g�ЪW��du��;��_�n���P���_$�ۜ��/\,��?�u�W���۟T�6x6�>;��gCU�����|�GA46�{�-�6�����\n�=o���r�� �.o��,�9���c�3^}�x$hq=�ی��jVva|1pj�ˇH��r��Q��R�&�9�{�gt;��o�/G�W�W��i����ƛp�&����ҵy7|�57�����P���фK<>��Xݪ�ԫĳ1
�~F{-E|cD:ٔ���{����9��Y��o�.@��`�V�r��܉R2�2ː�����v��nJ��	@'�%R.��XT�J��5(wʯ�Mx	3�H�Mz��T'����&S<K����	���o�Ej��������3��������.��%v@^r�@������P��� ��f�6��G�Z ��Sc2h���s���k�QB8�T����^��y�ǖ�E"E�}#�r�z��T>s�;v�ȭ��lƍ�آm{$#��6�7o�Z ʃ�j�@ZE��t�t����Gg�բᴏ��#��'��~��߰9ԟ��l�U�|}oş$%����%�Ϫ��l��y~UcsFx��Ң��̢t#�.�	��{>�&͎>`$^��wmpn��ű�\Ő�-����0%��#�-�@�Ƅ���$by����B��w�sM�&-H���a��Y,�"w��=���]�Λ����S~�@�K���e�����2[=c2}+w�W21A7��\�p웰3���ϧҸ���Ƿ���1X�{#�0upZ�^�iq������E�a�]�<5�6�����o���3��|�������}���pXi�4L����Df�_y��� ���v��]���y��}[,.ۿ%�Š�Gƭ$�&r �1#��c]%O�o|�����̱9�S1K7���m�g:����	B(/�kӻuk�~ �Z_و�Fy� ��z8SH��xx�Lc��� �r#�����}n*'a�D�3:���?:�bV��x�Mʜڍ�'�q���ų�.�����"ޙ�? ɷ��� һ�l�aj�/~���rPW���<�C5��w�Յ��оI`"�{s���0�a�f%�F,�{�j��������E��z�H���h�C�`ÔW��+Ϲ�,���(ǜD3=�>�#��;�����ud��^��A�2���T�v��<m�|�Ȋ��N���7k��@i�fu�3i�_P����P���b���\��*�b�N��.����X�+��C-~�I��c�,QY�M����'z7�w�Ȍ�H�e�f��6�6�<�G���%<�:����b�z��U��}�5�JWZ��,����d���!u�*�����;҂F,���9�S�(YF0$���_pN䳲��C$zlQD��Pc��6/�B�ih�ak�KxKȤ�gcݮ��Գ�#̋v���"`��kxר#�!�FF��� �7�x[P����;��Ki;G��%Cs0H���23��h`�*��?T�s&8��׀��\<e���|�a�T62��E��_bX������3'a_��4鷷���:�o�K3��֠[Q��������0�D��
�O�0� {�4I2�X/�a�w盝�͉��E�NIA��!�����>��Sj��%����%`�C�/ϫ9��Qb���}^�X�Uت&����`����x9S��*/������8Ŕ*�Z�m�]�ΉP����������=R���+ V���R�~��T4���A�av<
�rZN��'�[7��	�4������ �M���V�$u�4�$�A@��I�xb�j��K)��m��EҼZ@���p�au5�x>͎ڐ�M��,�����R
lJU!Z�̌x�ZC��9>ѿط�a�2��ĈqT�!�(^TIc���*��e�����8g�� ~߄��m�s�rh�u]��]��_O B3�*:��0���>��MA��������˺A.s$�(��v�_�P��N!tu�Y�: ���&������JS	tFX�
�b#l�>F�=�jں�夕�����p��,Wf����߱$\�Xf;q�'�ڠ����~�D-�7���f�`kA�i��e7�� t
�E�WZ�J%���x�e9C���x+�4�x�����J�+�5�֏tr �S	����$H����PlCX�v�I��T�U�(����З7-�q_�-�ʬ9���Th����PvM�9Y�<:�yR�e �>�8�|�dD���Y�۬3�qv��j  ڤ7�Y(i^�K|c��Cǫ�Z��d��۬w��s>��~"ruҏ�W]*�:��pX���=����`"("��7�X�kk��v:í3��RG�DR{c������L���?"Bk|:��Ӆ#���d�O�Qx�<'8g9�`J_UX�U$o�xy#�5Լ߇�- 	��MH7��_X��J*�ZD6�D�$ �F�;F9��'��>�.DǠ��D�����y���[p��s���W#��b���ܮ@
pT���c�Q���R =W��
�|��7m|�. �R- b�jh*�n:�m��Y�0J	�8ҸsREER�'���=��OO�P�Df�����8��R��d���yK��Q��U�Eki�xvT�Y��gF��,�<D����>�pC6��������խ=j��`mo�lRD=�7z����&cy|���@���Qk���li�)��㖗�I�L�f]�4.�4�R�<:�ځ*�Q��/.A6��}ߙ�ð��[�,)��OWE˕��@r�qx8�D�/���*j���f6���Υ�CQa_��僻�XY/id Zl����s��~�m�c��nE���_S'G�:U���tQ�.`�1���϶�vR�Bk�`�?��<�:v��_t�HR7{.4UzuN�Dx%(�+���
pHhϳ����x2���,j�}~0C����cr*p������bÄ��XbD��t���4�#SX��ȓ��pF�����&<髤���Aөa����ʴ���}���)H��"(]I	��b�ݾm
�����.9��EX�3�(��!�v�.�䳤��c^<Zx��X��,^�Vݡ���|���A���$�*��)��]�%RL���07���N7�
j���kE{(�Jot�����N�%�0�d�ܝ�e 3|�K�C;7��7m��|�h������$T>�%�`�\v������ic% "R��͋�-Z�+�$��樺�1Asl�@I�b�aj��J���������`e��0Yb�F������.��@���-������p�:���Z��W���x*��$�,[��]��m59�#�^�z�^�������<�A�jb� �{��� �����!��F��m7�/����JH���!��(��?A��W�
�X�HE�植r�pa�������l!���-`M�vXzUL�w�g�3�0=�)p�ă���P�i�r�sȜY���jZ�)���; N���V��ĝ|�ڵ�09�8����'h��C��W`:v�%�4)�;�1�bmr�E��or���x�ڃ|���;F١�H����0�gkG���-��N)�.��[/<�	ۅGn���F��M8^���=�8s�n��4� � A�A�b( zS�����AO��v����Ft���s�2�fv�V�6*��z�ΫE- L����0�c~d�jտ��^����<:��.U���՛|�um� kU:Q?҄e+i�ϫ��	���� 1,�����}�t�/�	x�xQ��DK��Å�9+��ܘ7���B��%����(�n�h��-��r�^��oK:�(Ru{䴰�*�EP"HR��yk&��.�S��>o�Pט��8�A�N��A$'f�gR6E/�eU��5?��F�qx(7�e3|�KV���
]��X�erb��;�4�7Р#Et�G�"W�2�]�/3�2�����C
P�ڴh�ɒ�iNlF������[���Is��P��v��7z1G�|� �7~����.C���.�^FN�?�<3j���a>}�	\iOL����X��'&�1x͞
��d��hk��)�ǫC���{��Ut*?��ؙ2��7#�A7�������;��[��TVKQ�g!���Ba�Ԋ~4[:�2�
��-�H���nOp.xx����6�7�a��U#'{q=�C�A�{B@�>���-�(ԕ:j=����W����2�l&����i�ZNfK��.,����"&�x�}oT�4Z-�����ЙF�ʼ��Nk͖{d�}>T���sX0>���?��r?J�NmR���v�Sk�Z����WW�����e\��3�`���c�C�Pܾ��>	lI�WiN4��_���M�U�E�;�c/,�_��3�Z���[4���4x����ꩄBR`b�N	vP����m�t؃�%?1 ��屷��٪[ �:� ��1J���2�g"��x��-�h��P'�},��� hqy�"���弄�����s|!/��6����_�±�n��Р��3��5ٲ�x)z�O����uMb��g�ot�5�nj H������=�&�`ݢg��Hx��t?�6���/o�f'���C��*�y/� �Lt�_'NԒZR�_af���;M �]g�!��k�&���啐����U��yܻdZ�%���S��|Z�Ch�{����;4�!�k�2�����k�Rh_�o#v��^ �IQ������z��I�h��^�4U���e���1��X,"�����(���܁a���hh�)�7��CӨ���N7\��S:V78�g*n�@Y�_Έ���+˸,�;�Q��-<�>�R���kf��.���a�O�˘�mݑ��q%�I��o��XJ!u�J�V�o�N��2U7JT{�,��Q��Jbϳ�$(�]�=U �uUy�z��V�'pM�Q�;#���v�H$��$�u�O�t�P]E���,�\lӋ���ӗ�n��p1��K4;2D$Bn�Aq�"m�Q�p��"\k��H�ḃ�ک�t2����C�5ۢ��$%#HK��;ԛҦ�_D�g�7��W�'�/���<x`� ;�]�7� +/O��W{ fVX0Gu{�N?��3�|V�
�9��*g���+��nG�2�/�{�2����/#=���=j`�0�� >��N�8�Z:�a��"�W�WK_���뜵�#p�Z��!7����ۛ���D�X�-�����,`��bf��a����L� �F4�N{�:9ηJHi>0��9�"z�L��g�6�Ԥ� <ajD#��k���[3D���f�������3��@��	��$�B�� ��S�v�a�� �}Yw�D\\y���t�4��(�Om�.�T�WYu�����	7E�aE���<�5ϼދ]Vډ�}������N�%�\8�-�ƒ��h�C�����S)̻��k����ܨ�Y���H.�]  *Y�UG}���k��M�y��S'�S���bfEk�pF�.����L�EepI�D#�������ߟ�I�q���&��c��v?�آ�c�SC�M������U��.J�oe��K����~�( ��mv��x�N��iN��w�3��y!\#�k�d)>N*�^�!�鉗R�Y�Qi��/��������oѦ���̣G�P�D`d�ۇ"vek0Z'��k�#z�6zx$+�M^�=r#��UR2 ~�6����xEV'����8Tj���,4�q���!K+C�����W���щ�ǥ�v��C����t�r�?q���;��a6�n�c��.�gt��%E�m�YD+��d���E���fɷ���6��E������T4��b���7�b�G����ä�"����]�"�<��[Q�ܱ��2v�(o�Z&����T�Q�>�u����1Pz���6|}y�J_�-tB<�Env50}��	QYR����&����}���Hk��A�R�F�������{qI���Քm�pԷ�r�q���蹭O��-?5���2C�Fοǥ���վWE�suي����5~���wo}�WԷ��+���h��P�1q1y,s_ ��%�j`}ȡ�X��h+�I\'Z�nKP�Ӥ�V�	n-}K���8~��[q���V���	[	�(��s�aJ<�v�;��'E��4�2�0���ѕٝ��4��D9����w�1�au+��g
�`.tl�`Z�����wZ�����Dp��e�ٴ�;������Ħ����Tї��L2�Yzz0^���k�s�^��Z���c�e��Bͨ�0ȧf�j{�҈Tk���`�lֲR�$l;<<Y��e㐥���p�y�����d2<W?WpL|`.^���3C����GEʂ��+�d{=���z�!�)�'�k��}�����[��سl�a��Sp��X��K�`�?�\Ѥ���'u�n��8U������q�����LsQ!�n�4�f|��Q���ǃ���0�ʖ2($���\�V5H\|��Sh�l4����=f$ʗ�oN��@�Q,���2XdCz����������U[� ��P��6�#C�Pu4�|4�pI�Gܚ�A�5�&,�f�1�$u��b�� 8_��O��0CZ��_�-C�Nx��ش�n"��?�J)�n*�{1���&�.�����뾁��OE5��_&E��df�lD���Z#(N���`j�gZ":���������
��}�{�1��'#yh�����$y���U���כg���ɬGH)�(�T��yuo�H�'%̃�'�hn���%`�6�-��v�t�bE8�߁rݚ�Is�X�=`= ���:�r�Vu
G�2w+���!�F_%����M�9bO�D!uu43�я�tP`k�K�W �Ɍ/��
.���Eo��|�4FtOlA=���h�������*e���M�V�*{llGʼD�� VZ��Y�����: ���r�(\��}��y� Ț4�t���V�H;��=�R~�"�W�Ϧ����rL/�|�S�&�ٺ�� e0.��TgYN3[VC���LJ�2���s�9���\o�>����U����/�A�%��W>{�LZ,�Y0n����̬�g�X;`яt)��^�{��(�|z��{p?P��J��D3Z�B/8ԥ
I�j�H�Q'%p=���Z�ؿ�<�b��;���0)���&!(	��2��-?Q�����'Bop����N����N����p ��H���]�˻�r��'��S��)�#�)������ ��������g��%~	�m�لF׽o��}6f�4��39�/j���(W���ovb���|���� Ȫ��,t��`�v�lI�v��c������R���5�y�z��_�f����	)���~��7Fĵ�A^D�%����j�������K� =�F���P#��RO�<S�+ڃYް�0��0k�2K��k�X{�\�{�R��#�lm�i����R�MVSE���SzT4p�⬚uHA�Gפ	�1�[?'BL�0N�>��D��Dʶ��"#^ن�x���$�!���0b�D�Zs�'�2�l�����U	���p�&�Ea�:Q_�P{�8�x��N�DXE�%�@m;�M����M}�S�5RC����gg<��`�io��#�f�\`;��P����7c<抱s4!�T,�g��p�/	�>�x�O�_��~�Cw��D��+���5���9�hz$K�bGܠ����S$>J_�E���һ�v�������o��׻�9ks�C��MVnK̈́N���'рB�+X�^+��@�����v�������=����d`�{����W8�k�& ���+>!��}f���5Rj��7+Xbp���1%2z� �V���<�sƖ�������R�@�&?KVވB,�p� ���&Q��؟���b���÷����~,I05��=/H�h
s� ;��E�q[�� �4��^t�|6tI"fZњf)��.��^A��kO�]�M)�]֨�@�X��M�Q�S2���23����G���3"p�r���&#�|�`�wo�D�"0!���;h�܏�������F3Ͱ6R�w$��4�Co1$1�Y�8���Ɣ|߉��%)�/��5��#%3��6� p���Nt�d�7�%���!��T?ށ�;��8���X&������
�O���<����He��h�C�O*P[PfM	{��ݜfW=H�����e�k�6D����_���ͺC{i�޴�CA�M9�ŵ�/F��C��X����3ǩ�B�);���"!bQ8��&
�?Fc�i���=�s�9㠅�fx�MVSi}3CSWUl�^�@��=툇���9�v	~N����م�d��ND"�XMB�\��`�H1��<}>?���� d���h��Xn��zB~��G�+�h���aBE�ʈ6鶴���?W�Nأ,���8�c�+�7�[�04e������x.�:���v`��+�T����ap]4�����Բ+�M�WLU�yU/
�,���x���1	\��CO�������!&� A@�i��}RN�bs9�N<�fd�U�o� a�K��@��8ĲW���@�U��R��7�u%�[3Q5U��g���\7���S�ݖ�]�����1����ٔ���	��!�Y��襓��.���w����9�w�N ��	������;.�'�`�PkY�R�����鮞�����;�֝1���,��Q/:���aÓ8So�y�~#��]����ﻻJ�����)��p��W��� ��۠9�dy�(���9�d)�b����G4?܀���m6�F�$�2�46�3�~ymv`x \uN�R��L˫3��H>�C�Jϝ��$ƨ��/t{t�<Ԅ��I/���\X��ro~h9����V�\�~~� �^��M���J��q,�9�ltO�R�Ľ����?d��������Ս� sڟ�I�ZgW|�d��#��j�'�vck��́�����"�}�x���#����O���;n�����$��y,=�ڐ:�6 �?������mQ�����8R�*]1d�tjz�$�!�i��_N%���qi�d�W`��DsH)6զ�����hr�BW� �t>�7e�%Up��ԃ �t���g�~���1�X
�w��*ݨ)Z5�?j>� "ko��ζ$Lb͚�q�wj����ڥ߉ޙӅ)A.09��O�^�KKY�(Ӑ]�J?3ݞ��Y`LDthߤu	���rPV%��Q�|�V����@h������I�n�f�斞�]aVfW�UŌ��/轒�,�WV�AB.�N���(l^)���wkjӎ
˭���i�GJ���[T�IUd��e�eY*jOxOB9�(�҄�\\��b�>=��Y��*��h��dBR��2�M�lJDC(��t����d��S���=�2.�(Cp�kOj��L ����q9��YyZ�	l��j�_�A� �+��j�.�߆@fQ��d|H�M�j$�"t�v�o���Sv��i���\er��T����Ui�����3}n3���2�p��sn��מw�_K�y��Hmpµ�� +T�P�97'�̀A�s��:�$w?�P���u9=���ߍ4�S�����7�&�Ւn�����XZ. 1�nH+B��EA\�K���١);^����CY>�ol���)��[�l}�$�t;���c5�]��v�+���2��T�hg� �E2:��N�)X�ڷ�=ΔUl��^D����a�J�M�]���Vr=����c�fw�gm�Ԥu.2��]j����|�ë��u
|���[��leChsZ*��0��rYO�͚�.�R��dV9� ���΄�RA0t����e�2EG��l�dZ;	%b�w��$+�C��1�9�|Bx��Ef�C����IehY��렋7���.v%�\����^��S6���c���򗒉���7�y�~�^^���k;[�����Ը�ʥ��N��gb�\��u�W�:���@�t>�6թ�_�����ѩFk�4�X���.Z_�f5��*-�4aF�pK���er�Gj�(�P[��_�)X!=����*y��L�XS�ÌH��	�UgrM���b��oY������D�<̺���ˢ�q��9w��I�m+C��ƴW��U'��4�j�m�hhR�U�p�X�#nq�@�$��7� �i�wc��V�����`���J��e��a��:����������~k�C=ioի�r�����v��3�������~�Y���MS�������$��3���g�-H�B��zd�xm����FqE�Q����c�~k���!�*�J"�V���w���=S[ȍ�o0A��6�+��xh�.F�1����#� �f��ƞ3���`'���Tg��Zԧ��?3)�䲀���9��rыK'8��yy�;������Mv��:6�`�"]��j�{$u����@��Mt�eq���P��t��0'�O���#����;��s��f�f�,�Z�^�u5S���b�wq�ѻ8K�,`=�Ry��xf���,?#��ɗ5��Y�Ї]KV�s�ՎW|�"s��d�*GʙDD؉�r�0�]Oa ��A;�<���#Χb��T�u^e��8�ɾ���Gq{B���R�n�9sx��_�C�n��>.\���2<��k�x�P*�P('���}�Z�S�E�b���Π�X%?��.	B|�dK��-YՄ��s�v`�Zז���|kl=(o�rՕ�}c�-r��t�o6�7J�V9���h;G�)�ԡ��j�f���;߲�cp���gxhc�Dd&����x�`��������$J��>K��lj��W�{���j�:�F�+�����	�N�X��#_�L��!�r�S.]�Cҥ�Q�������=�f����/Λ��d ��j1��`n[�Km �]�6#��G.�5f9��d@�fd���ɗVmT+V�K�~�V��j�pY���9�!��ϊ��XU"=P�oJ
��L�Q�H99���.?p�d��S_gZj�+����׽�]�����G�C��g]�(A$���?(�\���j�T
ru��h�8��u��7��R6�9C�H3W'�V��8�:��&�ټ_�f�쏕�X�;� A�Dؑ��0�#�]��0������G��d|��AS-��E�ǿ
{~�x)� cD:8���G�T�B[NI@"S,)���;G�����r�׽Ԧ�̰R�Zqd�[e񖥯����T��ǅ�vS�
�)�:v��L��?A)��L�:&�)%�,�tk;�Se��k.U9D�;���|ӹ�݌�EQV		�	�ۗOQ"o(��bu�A����:F�9�A�yf��&�{߸�˟����v�����q��> ����qf��iɩ�?9���Q�6���_���{r�c�K����'k��j�-($�J�*������ۿߪ.��~�AL�c���ġ�X����3$ùJ�'Wb��"�-0ք�pZ(E�B	j6ˢ�&ۑ��9,d�*�0]�Ҟ[�@06��Dr�U%��ވ,Z����m Tq��M3���Ncz��{�8��&,;;�j�}p�op�Ɣ�܍|�O۳=�8�����6�:S)��}�9�����Ĺ�.���glg��]4L+��'u�DG�QlY��7�L����ݨ���,�7'����S_*3d�3�T��b��R-�}TV�dǡtB~���f����V���G�;�����8&��5,�7wug���������N�>�h��8��0B_���C-�����X0����?�o�<򁉈�^ �-�M l�H�a�7tDrk`�8�2v��xma'j! cɲ�fG����8������PIrǫ��es��;�-�Ko������q|R��bP��4	%�v�τ�ߣ�~�h�\��$����f(��Ff�b��5�:�>)'����$,��ތN�`3CO�S���L��8�z�إv���8�����N�&�,�{�s�1���L$,�hĹ4���/�wd�*��f��i�����#|%�/n�Ȧ�Q��"��	�D����QE�^F5%|�du!��� ���בN=E!� �g����j.3v7�;�~��£k�ѝ�7��q��?8�Ѩ`bP���F��x�b�\ �Ҭ���b�4ԡ���Y��fZit�M���jG�z@)9���@�`^i㍁�T�- ~w3�cv�3#�.��Vy�)�A݌��{�yX�Aa�s~��B�|>�L�:z�c=��MĮ���c[�fp4��Vj��n���Q�e�Q1�|�?`;}�6�w�e��!n:��D�d��_�"�U*�U����࢓�Fx7��?���GN�n����@?���Ѳ�p���"|ʣ��qv&[n���=�"Kpw\�<�s��Ĺ�sOt���
�a����4�o�u�vlW�5`c)�i�b6��-9�V�k��Ec�Ny廩��P�RP�r�oD�ջ�ަP�)��^g�Sn�<�y��Y�:>~��e�D_w��Li�'�P�����C)����>��VU㕸 ���o�|��[X��ݼ�+֬���X�<�}����/m��TÚV̿�쵕dlaXo|ތ/UǱ�,?BEx�b���?̳���^�,,y�붳|mE�bX�j\q�Gk7Q���/�;��<��
Z��<hc�2�yt�����䩗��@`ke��m�Bݘ��) �2�mk_�1#�HQh��*b�	�G�8
�N��]���ýQ,N����O"�o4)o�l&$,�N�\g���L����u���~**�u�ъH2RZJAd`Gcs������yI��h׃���F������Nތ���c��U�g� �܇�����`����$��;�0W[��8A�p�?����� �5z,!t%��K�5/e*ձ�Kk?��1�#>��+���ٱse_��c)��JyZ�>�,�&kj84��[�tR�L(2�ۮ�l�����Qd�&��.Ma�9��ڪ��2{mWd��r��C� �Z˱��+��6}��'A�_�ÊQ�B~bI�du�U���U�i�2!�Ҹ�	+��4�Ⱦ��Ő*��z��� ��Ne�h�گ`��VIAa�<����|�Uy2�i���7r9��1�ҷ�1N���L"��eN�9��١��m�uYXX��RUf�мy@piّt�Q[�;�]m&���
�����p�K|v���=��� �P��~�ԩ�<i"Ӂ#Ӕ���K���dSa5�2_hlր�����y���u'��Ж�>�7�s^��16"�Ul,Iw˶��0�O���1�t���Z2���QA#>��В�͟�[#w�L�0��+�	=7C�=�����^ ^5�u�s�/$�x�tB*��#��x~H'QoZ�Ҵ.Wŀ�4
�D�����Q=�Z@*���ӯaPH��7�Cc�8`b��RZ>M��Ky������W>)������"��o�Z����=M!]#ji����,sb��-ؔ ;�薻s����A��/*����ǵ��4��i	u����Mŕ$5���ā��H���r��~"��FՀ���t_)98�b���R��6/�9�3��w���Jg��i��X*s��?�R���q��.���
Qljģ�:5S(�k �H�ѕz`�����3̘��*�&T��_�~��"�X{�%p���<����:K~3.�>�_�)�ذĪ�&ܴT�R��A�,_@:��]3��������,A)�Mi�G��녏� �}�Z	B�j� Zɇ��C�N���	��$�d���^l1���W���)�>[p�`8���\'��\������pk|��^拢��u��C�d�n*f�h.�w#tJa��n#���E���m��CN0H)�U	��lU�)����>����Z��u��}�A�
�ܵ�A} �c�Q��k�CC:ֱ��3�����a2Jk��g��KNM:�u�)�	��,y�0UD���$��/�Y���ڛH��5��8�?��a���Vh�� ��L�]%Y�::S��!x>U�3'��w��s�w���J�R#MD�N��t缣�Zq���@t�*Ꝧ1'V4j5��KB��j����(,�.L�d��$�RY�����V��L�yC֦�#�#6�B9�N#F�j��+�%.�G�������6(��-��w��o��l�g���y���@�5�M�Ca�����pI�)^J���լ�R�^�9���TxP�S��/�:�k5�2�Jh�,�X	7>Bfc&�����-�땕�t�s��1��^䜕"G_�T�*�Ϡ�Ri_Q�+�ӌ� ������V �O��x�j��1��xnV����e�? H�"�B�b����8��w��턦r�H~��72�e�{
�����@��������E� f�93�	.�ʟ�-}��ɳ��-�=�%�����9�
��$Z�`�����)ܮ�j�����
牍ץ�S�o���)D��r�T&Qe(�	d��tz��X�'����\>:�&�V~��A��-m��G�������������"VX���r%RW�<f�Y�D�3�ay�M�D����X�)dt[���yC��Y�zM���ʯ��\Aɢ��U1�o��--�#�Fh�u�:M�AF�}f��1e�F"�?k��]t����4���l{r�|�;�٫�,)�1ܮX��\��@�-i'*Hd���V�
�-r
��v�y�@s��(Y���߅�lj�x�N�ZT	�qȘux����Y��ܱ�B�'m�[���BB����ܠ}�_��^�{���2��� �P��ʋ�pɓI)�V��Yє~{'X.�������EF ��ݖ��I�]�d�NH	�?�����K��D<�N�p��t�r��;{�u�Y[�����5��cx�$7�-�N����8���8'QM���q[�h9�5_���x[@�Z� e���Ec���b�T�(6(9׺�%�cmlx��̪Dr��0D��]���:��������-�G�ܧ{�ni�eOQs�j7���n�"\�%:US��ضY��x6��Z�H�8$1��>El��)P�X�xY���y��}��5Y�~��6�BX8��w�w��>�Oa��6k�+�rg����3� NuD�)E�p<n��&+��U?�b��8�2-��9�}[Q�s%�Gٌ}��=D�=qz�N0���E������ ٶi�G�
���C�.��-,%yk����$q����*=p&���|2�� qd�+#������L{5��#����H��(����b���cL��v�`�t||�H!<@��ƪ�������Z����_�x0���}g�b��FmHR]D���O���u��p�<��3�3\�ЛX+��_��� ')������9*O �{��H��� t��r.&�x ���w��4Ţ�B��k��g.Q�T�"]��*�a�OW�����Xg\m���'�E0,a:�µ��8&[��;�`nu&����꼠T]\�-�ȴ�ҊYR�c0����XZ?�{�d�x���$�C+�����j���rn�kh�*���������=�%Gqn�l�>\[�I��SOdi����4�ͻq4����#��B�7̥���vn[F��2r
��̮S�%9�6Ռ�g��4%�P���(�n����1�Hԩ�K��h���@	�`��'|�\ϴ�ԗ�ܦ��A���Nz6I��'���4�;��dԕ�_�6W�-��!5R7pKй
ۈ�����~���/e�p�$�`�f�#��JmQ^��
`SP�el*p)P�7*�Q3�frT��<t���W�����|LrHY
����|���D?C'`��e�������F�a@�A�����������~~X�R¿���+~���E`�s7R��¹��H���W���A� �(T� �L{�6XJ��(q��0}|#�����c�W2���k��ô��g�B��.��s���y��#�3�jm�=3]�cf�8�'�q��K/i���y\^��d�.��NM�ϗ��ۮ��r�LW$�-��e��$�Lf���ٌ���R�Z�17^1
9�̶M�Oc�9���Dj�b����m/莈��<к��/�D� ͏p�E{��-iZ����(a�e�+`�>��?ȓS�7���,�1[Z�!��^ƀ���L�<=��!����k���Ԛ����4g[���vɫ�M�~�@��qk�;��`��?����I��4IKMR{r�'"�ӧ~�-s����gOm��P������9���}ж�tJP{��H�=c�⣜��_��O���h#Z��~ �_�~�J�����U�ΨX�5v�m�7��O�l�:[�4t+�?긕8��N>KI��+O���v��1�˰��y4�	��Pf8?* ���e�U#)�7�k�$�(�Sp�MtA��Ed~�5?I���-;<��P���3�&�8>)d�L���>)�kh���%M�YaZg�FkK`ss�p9����Mi_��&�p�)��׏�Z�3�R4O�߳ċuƵ1wn�Ԁ�oa����-��pc�y���ƣ��JuqޢNg��nɗ�Tj��]�/��9���C��x|��y�����s�;m��b�ijӌB HS��������8W;�����fI� ������i)�e��ӿ����;ָ_�h�n�����:�l��ś]��w�1���*&��#Ǣu���_NV��"Q�m��f�����	/"��!dz"_G٢��d��k����f<�o����C�K�-���wBp�Nt����4\��j�h���6->0q�L��v�7��7��T?��f%H������\q�J�F�S�t��
a��3�uQ@nO�})��kh��{�#���Tp3��bY�d.b}��Y�h��I0/ʟ3�V>�
6rn�J�r��%6�P��p ):#Io'q�K���?5A��o*�z�7��Ā��2/���7b��I��9GQ����C�pgr(Y�{b�2"��u�>WYϒ�z<M�`q�U�{u�ύ_���b?�F�<�J�xdď�b7-o4�w¼k��@��F�M�&�ƫRu�]�mP�P��C8.�Y^4��7�����
_��_�F��3�����ׄ���BW��b@D&\3L��)�1�u�����oX��n�L6�Q�K60~^f�o���i2=�xG)1��k� �ɡ��_M���MF��В�\�	�Ҳ�RE��^s@���m]^�ǫ�!Xz��5���F�&(Å4�BW��
�	�֦���T�������*Tzj��١n��,Z�K����^~x���(�wlV�0x��6q���5?�4$)r�
1
m8���'��t\�vq��L�O76�|Zv}-��MD �~��y��%��.4��������&�Y��o�4����7lRz�����ന��6LA�#�|�^�S� ���2�����S�Ҏ��4�0��kt�T� ���#�-��Bd����~�}�2X�Rs�]F �Ԛݔ�=�r���F�j�J�p�?e��d�0Q2�W*�D�}4l���+$�HrӜ���\U�r�fΖ ��ufAIy����u��R8�ЂI�v���q	�|��2�6:����ƻ(U�Z�"E��,�L�;h	�a1S��0؂�G����G�GH#On=bɵ�{P�l�.��G��D�|5��y�������_e�:J��3�*&�@a�rV���YM�"V?���1+��f}e����V��#���ka����އ���:l������a��(X&<TK^F��	�ه�&���;S�Mhl^'�At/�)�Fc�y��7���hD��Q��P�Y4��u� ���o�ʯfᘁ�V�Ҡ�k��q�_zl�g�dƟr_����v����ð�E٭����&��"X2g����G\3�s�&�*;h�q�5�$@t�^v�˘^n,�]�Dŷ�T^�@苽7&�.z����N�@�k����r�kk��s�f�.6u+��)�Mt�'�))����=\����G�Os� C�q�,��Q�={�v6�˜�7si���O�k��oFE5!,��~)[��X��k���RmY����i	�ա8%�-�/�p�&�b���%"Mz@���'䌻���������sp�e8J4�$a�&
;9{N=���mU�alͧ���6��ķ�ۯ5�c����WE,Y�3�B��3,��F=��������+�B�
Ó�U�'=%	1�~i�6�QL4?���:W���)S�����*dF,[���i��B���S:}����Ig�u�a> ��G1P]�nߥ�����̤�n�k��`��c���������%Uz��QV,��7��a����)�p�E7������Q�FC�n�`�6L�o!R֧��>�я���T,��0e���G�r%8�S�T��ϮWQ��r� C�갻y�e�dM����=>0 G
[tݝ�c|�X0��Ԕ�6�E����ū�UTuB�:�:vКAʁ����p!�R蕩<��*�j�^jh�����[�bB�ThGt���'�+��ʣ >o�Zd�Z�������&������l���1+6I�_$)9������)!�:��KR�:g�*~���hIckIB]2�8��D��� �v ����	�����=�G{H2<���ش���#��0@k*V���Eф'RC	\�?XY0{@�	)bUl��kK}�X�=�u�Ce��g�t��x���0��ȲD��&x�n@Y�[���_Fz$����,m�L�"H��K( ��H[uZe`���ՇY-�ә��:f]�i\J�}/��n"����-��.'�t�-@��a"�ǵfb�) �W��Ӂ/R=�k�$����S/C?)��@�dio�/����9D�9:&-�/����#��pt?1�;��5"͂��<�@�2q�/�wv.
B�Q�)U~�Bh�1XbP�/R�I^.1�\�$�}�+y�4m�Bj���.ꠇ���.�gޡd����7�z�ӯ�b��Au-��@�Kʒ`�@M����X� �ӊ�;֖��7���W��/9�.j�ϑ�1����eŔ\�C���N�-�~f�w������_=�RFy�o���0�2�X�r�jcg!�Zu(�*�lV(p`��`ۺ�m��7CP�m|.�5�"��S"�����:#-mq���7���%��� ��ط�u0ֳ3� �f�{�)���Hg(l��$m*�ݟ��Y�UM�xfB����XtH�wF��.[W�B9ڷķ��a`lPop��+���@+\�۲���h9w�^_�7C��x�[��~�
Z��ЃN%B.l��V�&K���D�� �K �l��-s�duJ�D��.���+�FOUV�WL�ǚy���9�~�a׈�/tuD/����-Vn(�T��@a���#8e�@���4 F�n�:�M�u'��[��f�@5�K0�E�it��~n�Iڧ�9��l.��V@.�*�7OGǰ-(pҿ-3�~�D3�͑�Y�𝨱� W>��H�*�m�L��Eoe��H�����0��Ѡ4�R�{-*�V�
����xƕ=}��d�\4�p����8�[PU"]z|NY����o�O�d�S*Z 4j�&O� ?���m3	��^b��m^������0O󵻀^	�.=wqF���������E�${� `MJt����^/7�x����	8W!�7�X��k�)����4�T�eh]�h�V�
u�'�7��Z"�m�3+N���)0}j8�傦��H~n4�Ů�S@1<ֶ/+�EΎ���Q�4���L��gfy�ϯpɘ�A[�Tm��|K=�AE�Vʪ�5��Q�-��B��o�to�p�oZ
�G/OF�螌�]g��ټ�A�Pq3�;��@�xw�q޹qx �i�����N�Y��a0�0�"�: !\��i� O[��� ���kGaF�J�|���.
�;B~nT�P�̊��:�����]�*d��a8f�T��)��U������`�f���!��>���3L�|�z�[�y��4���.����F�~��HGB1��.7�Q��k&#$j�t*Y�G��w\������ՠ�M�N� �F�#��8"��9��}l��m���#[�;.tm�A�x������qWw���cu�iO�蓥@e�Ӷ����c�f�E�xJ�����Y]^j�����I��/���݄��y�|k�9R��w5\Z�j�Q�܎�h�6�}�h���U���~}D�����(���B��TV�0�O���QU����H�<&���k��Un�+��>�%�e��Ra������4��?6�=��@Z���P���J�(�5��];ÿ�
m��"���=��~B}�DF9H��]bO�GӠ�ɠ�X:n���P����	���\jRa,����G�0�5^�{ϟ��������s��~=8׷��o���xF�/t82N��v����v�2���]��h��T;O��D��NA�zLb���Ԍňg���\{�5�\\�L#f�'Qr?�w����9�.�U�U��x� /3�e�����g�@DD-�������@(䄊=�K��4OQ�N@�'ʹ4I�h�߭m� ɦ�[�K�&��hB�ɳ�=��5{�J�d���9?�Bѧx8�U����f�.�gF��8>������Ǫ̆���3�0 ���x��[5��)���3��DO�@Y	���o=7u�"T�O5ar�dg���R����鍝m9�?X�z] ��`5��"f�� q�W� �51�,��8g�_@�Ek����CuzQ�l�t�îX�{�>q��0}�j�_8�(f��8Y�O{�>]f���z6�n�WF���`b�B���/-[+�VU�U-=�L�O���p�`�oHF�>�����Ne�<�@?��>\�u��ȼ����2z�����Z-"�}�O�S�'�T�a�J����5��3dE��QwB �`�w�zI��f��X:��%b�$�wt,��|$N�*��5��w.�����[f���|'�tR
�<�_q\;���� 	��.ܥҖf���$(Iq�8a�� 1
U=h���b[����֩غV�=���8��ӼyPN9᯻���%�OS��aU��*�|����h�!3���'��_�BW@�W���Tpb0yR\�\3�s;�t+��}"v.��`ڛ��'I�H��l��elVlA=�ڧ�wC*NE����v�h�zع�q�u��T����x0-t�!ߤuF�iF�t�h#QT��;Z�5(�2e�|�9n'�WR-�!��e���j�Nd��f/74D�����b74j���	[H3Dr+�ᬰfN��;߉����.ba|~U�Q��)'w��j2�mD���U�D��q�8�mb�ᆊ7U�ڳu��6�-�:���������
6;mbd^H��z �F�ʈ�o�Y��KRxt���u���,n�Ʋ$"ʆ���ˎ:���H��Xy�µ�������������4�b�|t����]�Qd��Z��Z�Ǩ�Z'W�=�h\��5�	k�B���ʂM�sh� ��о�Q�z����a�:�DQ��j��6��ա��A�r�������[`�E[�v��;���#��~S��Q�b]
g^����W�ڎ��km�^C����]�|�J�c�n}���}�9�`�:�{ژ<�2�������o�����}}�71fn^{%5��dT/	~T�$�ɞ]ہ뻍�D�&�x�0��?6>��>nͷ�Z.c�i���~"(��x�eD��"�aӲ)��������A�-�k��<[���};�ra!��h�$�v�����Ktx�aҌe݀�U.�� �}?[�Zvu��'��/������>9�~��H��k{O���ƌ�����A��+�ۅ�R~HN�u+~��h���܎���/A�؊�&�4�#Ǚoߋ�2���j�O<J��d{
`9��bص��Ȳ��X�M��2�(nu�g��[Ʉs�T#S���%f
1 ۆ�V���R�J8���������l�c$�i9�q�'X�X�G篠�G�fןeM�P �s�'+�o�V,������<�����F.Cy�_�<,�m�[St{`ꞵ����e�e0E�͎�:yeg�h���r��T�����;�?�svᄀ�Utx�'E�j�R�B��3Q{"=ޏӫ�홮nƛ����(�1Ua�k�ur��]�q\�)l����l�ܡ���E>c@��j|��߾�W�;8��b����"��Q�4.$Y��:��[�ZR���:�5�.��j6㝌WE���!138�$�|Z����c.7M�GMV:��������[;�2�v��J@NG�rJ�1Ԏf;�)7?�k�DL���}u���n 

�g�}��a����dI^41Ԙ/m�w�J�!r�phNi6i�>K����/��>�7	1/h�[���ݒ���_+C�w�X�\�ٚ��ԁ�U�R��S�	�a��
Ï���s/�m]s��Ŏ���s��}�ʸ��;�	6�-�N%����h�(hE�2��Ik)����.��t��a�|�9E�C�qlue�~Ĕ\��*m؂�r�#�4%ɏBq�ܻ�K��[4]����W�����Q:�(��)��i�Ӕ����=4�Y�7E����R$�Y&�_+4�Aw���������ay,�h����� n�T��x�x4���R���W�2'�I<���j�Ð�O�s4��5�Ws�����r�]��)Z+y��`���Rm��tUxM^#n��z�Ni%@Ka���e��f2ڊ����}��'~�}�1>[ƭ�z�*L�RC-bK��unf���x*=MÝ�"�;��#Vg�H��m�nu��lV�5�!��)
�p���5~��E�F"j�'�c�t�����2�xO�d֠D�2|�	��:�N]��"ٞ|z����J��D�I6�?@0%�gTPyh�LܜfF	 4��b�ॐz�7�P3��� a��(D�1�j�l7�! F��y8�04��|�v��Hσ|�,>��]�I�ȝ��;�{z�) y���3K��"�ߙM��>E��/8�/T�!aa6Bk�C7�g��:�\̕v�tJ��{�u9˵V�bOiv~�a��*�%$G�qIj�Aܤq��qX�i�(mѝ�-�0	�YQ����t��¤`Ce� (�!��,Zyg4,�d��\�q8:�r=���6��7�`��P��xpA߅b�p�;��KZ&,d���F��F�G��c����A?'OY�i����\^�6|��k��R�퇟P�K^�`k�5IH��ٖ�վ)r��eS�a^���?�c�U���V���i�Y�;��˶�O�7�7={s�F�0��$~TIr%�Є˲� �Q|��L��m�V�χc��f��e���>��\��^4[΢�*Z�*��1ϕ��=��7xx?_R@֕�&қ�� G_Ya�0��??V�b��O���{F@�lh���Y���0Y2y�N����l �:�Z`E1jT���.p�ԦUI`��(R[M9�E~�=t	�p��Ͻ���`#�#�l�$V	���<���&]Bm�0���f�erM�e�ȓT�^�FD4�׿�r�Am��G�|`^�2�5��DJ����4H�B���������[p�*Ӳ��������� ��]v�WJ6E$��@�ב'�s$S�](̆T�P���F��^q�+��iq�g�p��2h"�$X�
1gp��˲(�U��J��u��O��x�4�3�e���P[#w�MU�4�ɬJ�j4{���!@��5R㍽�.���_���v{K�P�5�<0���	�u'YJ�|M6
���,���{�Ł
�'.���FhH��b3�Ο+����61i��e� )���J�Vw�N�����������Í�*xz_d.+2�=�j^	�U�Ÿ���Q���[�;��3T�9���|i��W�||&�������_< �?�,`�F�8Ct��W�/y��>σ��J}��v�+�OzeÇ�<�??��x�o�n7[��X8Y�V�߻{+�us��.г�)%g���&�7�nm+[c(�7R��O��%�Q|�_�]:�.?�z�(ˑ��Qu�V�i�:����c�O�q{��~ë_u�̮��G�	�.���X�c;,�:��ϳ�$ό��`~`��J�#H&������Y�/d��U?r�}n"=כ���d����D�����!W���qM1���M}�����5�������"ɚ����@zomC�L�N�#^"�9�D7��ʹ��ΤH�H����f(������E(\ɿn�(c^Aj�ke�����ő�� ��<��B�J���A�� � �� e��^F����5��9� ���M�� ��?��ݍ)ӟi�j�[�E�L�V��Q���U��?uʼ �$5��\ڠ �����,V��+�4:��(����-��S�ph�4���[�}��:�"֜-����p�F���2%~�S3���|)~Qs�ˎ�n���V�^A3s��6���SZި!�;�vd�캽U��ҥS#��.@P�O/���L��&�p�����!MV��6�?#��T�r��kHe�s4��)��2Ф?�)�4�|=��1"��a�/a�}&�+�>�� 櫐�����kE�(��As�@�F�z6d6#��V�8w�р�)$ ��Hu����R����d�w��Hؘ^��P��&j�'��GDuUk������YS�k��k�B�Ս��&�O��B@U��+���#��UG�T��r����������_FZ���mM$X�\��m��{.:��9���`(���/G��"��@'ȩ�Wۛ�g�䯻����L���n���*���Î� ����x�M�)d�}���Z���!a�~�t���W��J�l�g4I��f~o鉦��.���/�e6hC5cf�݅�W#$���Ǔ3ގ�5�ަ_�uK��K��P�������,�?�j)銜U��Lb/�+YK�X�& v�y<mB�1Ү
W)|�CoG���0
غԬT*b�U���*}��pZ��Q����-����T�*t�W��^��m��{��} ��Kh�9[��!ς��5Ɔ��5|����DPN���w7sS3�!(�N���L�7y�X���{Яh@�_k����mW�p�>�q��z�^4do G�1��U�/�o~��O���"}y&��F�s�/��v��:*|��iC�8Ui��*0����8���E13��᜹_u�[]�
;�Wg�	��ۍݘF_g,K�`M�6=�\���*�yz�b)�X��������>Ǳ���R!����ぷ�5�ܗ7�����W�8�3���:4@�(5tSq��"Tfp	�~�<A����%�鼒`�\(3C���2V�K"���24��Ɠ % /��ڀ��Y.�����a�U��Ɉ��+�	s*��eƚu��X��Hu8BN�x+��{�b�޻z6�!:o�f�F �;oEw�����O�߽���"(GR��}���M��ІQ��:My�����
�M����m��ΎR)�gϟX����.�Iĕ�t�������?����Cn�t(ř� ���Z����1-�R;���	,�>�G@��Ә�
���*y��]�!������$�E2Oj�8��u1�G'O[�#2�d�Q&�pޠNmb�����Tպn�߈�A��H�2;��n��L
iO=\����\NWg��� �+�Ae.�{ĉ����(-��ϧ��^~$|by)�ҹ�o^	�X*�i��rV<�Zw�����Q�l�����np���P{脑ž!R�4��ϙW�M=g,�/���
^�� ���s$���C8}������)�6�"a|��z���Xz2�7`���Գ�P#Yp���<}���E�Nݓ���6Ѻ��V�ѮX�4O"V56��)��uE��F��`o��~�v|�t��G1��r'�5��q. \�%o�y���P���c/���-�_��OQ��y�i]���WNgp�t�����US����E�A$�%	����ζ��xlR��X����Ju�`�n��)&�q����-��c���O�)}�͓0Ԉ�:7��-e������ƍ��nJzI��D�W�3�6'�]�\��������t�k��"�{'�g�w�kQ��U	S��-���M�@�d��ت���E�9��o��������g�B�.���<�Z�kT��S����1�H4��w?9�{k�D��=e����,m���\�t��eN��&s"��d�e���6F��ZČՃW]܆.Z�b�`�68*\���m<��\_�Cci\4��<�"%����R�yӡ^]�,���^�8�t��9\]�Y(��hAʡ���$�*��i��=�A)��ñ�*>���fb��J�!�(1dk������/���� 5k�ו+�(:��T�5���Н�^Q��%�7`lڷ`;�\�M�ЇW�\dq������#x���R�)0]+�!ݮA����ph�EP_
 �;aQy�t�!G�}�b<+�h\{��Ckn�
�����wd{����)z����@&|� �|�����M2����)/؂�G),e����m�w�˦�i���y s�	�P�<��ɖ������d��|��-���O[�	i����{����f��8����[�䕨��x%�k�X�ҫ�w^�/^�Ϗ���Qd ��
1����1'&tYcu����]���[�`�WN��B:�X|zf{"�/�{p���k�i��!���h�q��j�����������24oԏ�)���ƘcC$7��۹E;���p�X"ь|�VM���=`�aI���� d-�C�Dw��N�_g@�pЫ�� c�	��!�!�����v&��������;�fa�3Lt%$�Vy\r
�q	�*l�Ʈ$��onmV���6����X����V�( Z=�UߋA�^�δ��ſ_j\Zt�b���(�(�0~O����s�|��+���>���2�)����\*�pUII�����-W�Դ�@�"�אDU&�|��{�H�u��y)���H��z�%�v�A%�Ws���Omǔ��B�rs��,Ʉ�Ϟ=�*���ەR�`uv�^t1v$��u>1��k0����:>�Y���DA�ͣ+M݆L8�o���1 Y��S8b_dmТ��9rv$9��5%�2Uv�py�4R$�;<[g+���Mygp�2��8��������w������o�Ő�s�p�6�����_���{T� f%���qQ!�}���2�����%����#���!,yI2>(=-^�^w���IU�\$�Q���"N(ɻ�;3nA��9'��F�b�����k�lw�����U���pչ~�>�I_h	,�n�g� o�ͿUп��O�{�#s�m��d24�u	�G���.�i����O��dͳ��4[��gSZvb����j$�xA��5;Zb��>��DY?���< �/�����G��W���<�G��dyR�û���N��+
���d�5xر��j��ۯ�£�8tt�h��"���ۼ��(b��8�s�X�]p֔� C5#H�mSt)�k;�65��M�ݙ�����
(��^Ky�,�>�#��+� �2�n��}���B��'�P���s)=J��A+��I�x���3�T#8٦ܲ��/�X���o�u�zR�w!���H��������A׵�T��uXr3S��h��Lu���i-Ԥ�G�s�a� ��` e���+]��.Z���Z��֙^�<ȫ̔�~���[�Ś7�6��������y��k��N�s��Ň]?�Go�Ȁ�xa��W����w4;�>��8�������,����Qi�_>���q�||K���\s`����zf����R��%��_U�	�W-I��%��h���?���;���!�+��.ɪV�(�3�qqh�y�&0�wI�X�M��Zt3�@�z��i#e)d �`����U�"�8��8,�N��a�˼�E�?h��*bd������O~� ����ޭs��	�����$>G�|����B��M5qc?Ꮒaچz�9��Gd�U������Z5�����1fHx��o�oQ�/�	�����&�+,�Tei���B�I^�����4ʫ�֊���6/��}G��n�Υ6]��,��5����r8f�f;s�\�A�Kt0.r��V��dm�?�B���I \%�GB.��f��������vfϖ��C׸�i�^��}OPT�P8�evc���H�>�y�8'K���m.�SPj|_!����zb����f0���蚑��iM�4�L��`��j>���{�A����N��������C���Q�ja:��4	%�ƈ#��"�� }�s�8>�nhg�H��`TD�����n�_l��`��	cA����o��f��2��<`�7���O$:D�3�?K�X�G��5t�X��I8v�"h���D�mg�&�i�/��=�n��WZ�ʤ��з��D�<PR�����αW�S��q��(J��W���c�tW6+��P��"GX]��m�ue��NS!Å����5���Z���Z���2�π}3�%�]	j�︗�oK3�P\�7�Ts2M}ݡ�G���bHND��:̞�-�M��0V��oN�!S���*�F�N��:�G�~9G�V���Z���V4�i���i�n�Y�6x,���>��0h�C���X>*����ӌ�n�P�M��~��~�ԩ'O�k�aD���.IE1�6� ����&DqU�<����������^\Sb4�9J�/}�9�/����{4#ρ�����J9Nmӌj����JH�j����Ojl�9R����g��uoy��������_���rt.{ĉF*GE��CUFD4�F��Zo���lFIǕ$�h��"��Y����þ�꧓���R4�	�����u~��H�o�I�m�:K)|� "�UB�l.�J�gE� ��F����nI!Z8	��k�oC��3�>V��n,*c=n��=�^L�%�,M�!���;�r��O+��k����!*)�9�P�-=�{M�R�M��RA�P���}�6��Y��V��	=5�[��U�LQ���ŏ�JG� y���-���r�3�?�t*�.��1�ޫ2���k6�F���W�j��u>�r|
���9����������y-��k%���ʹ�#��LX��Ca�oƞK���f>��0���8����� �Ǚާ�d*�Y�<�څS�����,0 I�;�'��zĒ@d�K�V�j�� �QO�Q(,q�w]�y¨`T��w��!ok��)�g�C�q��Y4��P*�!��A��:�ed��\���4YO�lN0\k�u|"r��&��%��w���x7�^2ؼ�vf��x#G����������k+&򮚕�׵�����.>oz�G%�mR��!D�+{J�2{C�]S�%�
y
X��
�nMm�o��`8q]@q���=��7I3~�������`���"�W�6փ���4@����?��[Z�Sa�)�oѾU�>�CE��nTfH0sރ��=���]t��������(Y�V�=Ui�\	����s��	1l�3��%����^�[�$�_�����]���R����`�{�A�	���ɭ�r�W�������TT�8#�ƨ�}���j���po��["��p桔����S$�q����o�4z���%����C0(?�c���C�4�KRS�8���;�H�!�� B�?|�H��0%���Z{r?r.��ʣ���뜦t�RLXrws�c���=l a\�e�5Y�ɜ���3��p)+ ${�ZE��*�XT����H:�8,�$sB�Ҍ}4v� �A��x�,���@�X����gIf�&�*'��&P[r�vq�۵T�CG��l�g�@�����v���dm���
I�E�51#�+(b���Cϑ��F�Fd���澃����(e�!~m=�������F�j�����p�����MO�\Amo�Q��Ļ��L��w'��C��I�'�r���{�)a�1\�=Ѐ��D3�����%��X�K g�e�.fI��>�͍ :=3�W6���ΏE�R��GeP�̡D;t/�v��%�Q1�ZB^�� V=�j�(G�����d
�4U�L�ѝ��K�#m����ҿ�bƽ��)w�_�{�~�T��	7T�~i6��~��,�?����t�+y�B��@���b�1�G�(�Q�e��&�#^���Ns~a�̌Jc���w���),������m
h.-؜)r��lZnӛt�E�Z:�XIA2��D�S�h��w��ޏc�f�:�O�o�A�Q|Es�2&���а��Ti�����!E�5(���!�@<��\���\ॼ���A�U�8�B�����gfa��3�0բΡ[ՒJ��#�lr��ź���4T���FNvq3&_���u�8���[	-����e2���r����G�X4��ܳ�/c�4�{�V���I�d�;�2>��i8kn/+R�(��IK%����g�����8>	3�d�	[Z&���x�>��BUc8�x
N�`&��c�pڢ*�sZ� z��j�>E��e?��}��:R ����e�3�fl�\�_��xz��v�W544�)V��0��'B�dWo���J]��8cb�9����'n����������z�.������n����Db���<�B��W���/;zF���z�. r�$�SV.���`�#�5��T���F�{N7�I�NCz}��}�S0�We�r���������fh��aY��iO��+,kt��rPx�o<�Gu�_��\����R$�t�|i�bB
6g�U�{Llտ��_���_	�Ȉr*j!TU7,O����E{m ���Sg��y����]��(�Jt��в��[�q�EA1Kt��T9o�ii��VZb�t���u~í�O���yt���9���BW�����aW�,�,}�R�2��3�@��^^O��o+¯���]���jA���X���+.�J�p��k�q��c�x2O��%?C��+	Nq�e[�Fף芛v�'*F�7p*'�ruI=zK��k(i��n����܂Gƽ�}�Ys�b�~,�H@��H����Wp�Z&�ƣYY�\.�G�tQ��*��)SF�۞NN��MU�a� ���Lܫ-��T\���9M��0w [���� �mO��#�Vh�`�j�⿫	>���� >��9����wz6�}��t� ��5'`=:]w�D>��{�]r�{��E��?c�:T^;����H��/Y}���"��~.�ب�X4��_���J�	T�� ��8;k���K��|KlY�2r��++\	9�;�H�Ό2����5�X7+4'��	�nE���387 <��I�P6{�hW9��HKy0�pV[�W���$yJT��;�}񽗧Q�;+eH�ª����$�5�r����w����e�hV�(����Ğ�ݔ���!�iW��Ŷ�

��8E�j�#F��.b���E���5S?�:mA���-q'V�f�����=>�����g��LH���!�kW�f��+"8�f�u�Y�eiE{f`N����n��:f�<��Tg�hq�u}S��p�����D`�����ˢq?T@-�ǣ�$_`>�����/����ȧ;�f�:Y5�D����ߙ��\C�=jp��)����N� ���eJ�I�1BN�f�C# �|�k�q�/��31�q<�
Q)a[^�b�S	#�ZS�U�9~.�Y����ċ�QTm�FKM�f=bm-�̅�i�L&1���4U1�oL��!lup��^X�!�[EQ!�܅@竜��~�a���WXe#n�Ä�HW+���}�nm�2���ΡEP�����7wO���� �c��j�(|��3Ҡ�D�����@�	�o@�b���,5$�`��b�~�P`��H'*voۄ;�צ��K7�����b?�\݅��Ǻ�:�n.*rP����� >��W�dA�y�Ǆ|�0'�n����O8���7۱�iaI��~?�K߿�g�.^��T���,���}�����k�2���%m�P����z$(�*���%�F<�u�k ��U͉h��qI��SW�!�Pv�U#�U\v]v��H�c6c�j:�r��.s��(����01���ˁV�����I3��M��7�Jԋ\��7�_�Ru��}���
5�7�<�c4Zۀ���� l��v���*�8��S/c$���#`���8��whU�#ŭ��Uq���<"�Z�L���H̜��YL���C�z˺�h_ЁP���9�mEA�:��^�א���:W$�>[zJ��h�����5ıZ6Gԧ�N�]���Cu&�0�K���T����-?�1�S��_��P6�� G�}�!a���0A��嗒����)��/̆��Ռ����E;"�k+�m�7b�|�i*.������Y���w��'���͉�^m�J��أ	IE�ΰS��$M�z���B�=����@ƈ�P5NJ�c�T������L��[JD����t�7Ӓg_��d/25����h��1��7�MZ�)ِ�z d�5��J�;�A�k�_s<-��v�o�LUi�!ɲb��%��� ^5���B��+M.z/;Q�o7�5��c�^�j����~[r)|�vY n(\�nmu��+a�_I�h�Ul+���Sv�S�1����+ɓ�ʀ�2�y�B�d4Ԙ�`��Z��y�����& K�Zg�\_��&j7`��ѱ�M��I��pT	1]Q���BǕ�S>�W�
��~�&b���ݖBFvR�t���8}�\Zo4*3}��0#��}����y�fV�j6�8�~���	o�^�4M:����L��@#���rc-���t�������X��2��s��&�����1��%��3��[��v��,e�}���4@訲��yh�&��C�H�Y��I�W6���a�����I��Als��x�c$9r�}�w��Tތ�[eIڞ�՜S�q	�i����:q�U����MB��*����[�^3�L�P�&��f����/�k�6�gE��n|��u��;U�2ܶ�Iɰ�)d����͑U�љek��XB�];�%Ce��.rslc��]70��4�O��4��͈��1e-���~,��:�]mh����8TT�;���L�<��v�+u���+�����a�yS�r_#?U�_E��rz����G�$"�"�V,K�z
@xB"�,��n�������`�ޅ��9�?�l K�}�;^�r���1B��(��V��*k��Η>��Wo1=���KG'筀�-�;����v�3������^�ޱ���Q=�����PU7+���N�샣���&�~�C���Z��hµL���n���?F1CcӺ����c���H

�NŒ1��<i*�k'�ˀt��^}L6�}��6�%��IW�0\N{=�SP��]�C�G9.����:] �5}/
&.娸�7O��	�JT���}�E�7N��ae5b"jEl��&��~-�l�"�j�v������{A �lR���|�41����<��Y+��}���I3���o�5'��%��Iδ�d�3B��hh#���	����JӪ��G�b�P9tfP<v�̷M �j<b��������w>s��i�U� ɢ�]Dy��V>��['HR�t�NF�n<��B���ߐ�Cmfv�
�*�6q�KU�����1����&E��7�5� T[c;F����L�Pp�b��"��q/��	���b~�%/���>�aA�`����E�с�C����/	��� ��U(�pOlԎ�]���$9 �<{m�C8�L1L�5��{��nTO��P%o�&�D^x��Y����$��o���B��zO��(��	"��OF&:��}�(�r�7�7{�sǳ߰����+i|[��98s裎�O`�HG���#KI��;x�㤎⚼���-�zg���&����Ґ���;bC��p��:;��+J _`w�\����rG�i&.(��f\�9��*
W�����&R����٢Fw�Aq� ��Õ�.?�y��#��Ԡ5}gW)�q��}c���c��,�Ԙ�0vq�H{��-l@˦�i++��y�}�@*�X�Beœo���o��޿4����ݼ�VId�k"2eE��q�9_r��Z�g����i0����@��z�����F)y��� �=Oeא9��q.p�$E�:C��dE���]X4(g� �g��m���:6pfT;n���J#��z�K{eH�H� l7�-��[��7?B�C���Mm0���5�		չ�@��
זcm	�BYwsu8��]+�܅���B���y۾�0�
{����>f�P���_T�	�W.8��"P���%��6C�碑��/�9��v�ʃ����;F�NOK�5/�wn���_ Mg�c{Z�C��i`1x�N�FC�
��^�/��~\�ڙh�坺.��U������v�]̓�|Ĉ�;�t:M�4�tc݄#?O����9�x����2�"`�|�4d�?2YZ��HT�7T��%�`>c�b�/�<7��+
���C��Gn���^��t����({�Ι���%*��R.���*��V�ۺ��T8��q�R�:��tH����5�<f� xt3�%�|��Cxs�]>tq�v�Ͼ�g���|& c$��*����ȒϛE�$�a�<O� ����R�=(G�k��|�E�;�zRd��ÍQ~t��!Ԙ9������[Ld�ۡ�0�r=��������v�T_b��[�͞A_��!�*2c�r]i�n֚�����Q��O�a�8�0e�&4T���}��1����5��vܫ4zEƩ�����F+zI���+6򿧳��!��r%�o?���sM�&�ج b�n�o��:��{�7|7�����~�]Z�X�g˛ⴭ�a�u�k\�QF��0�6�{��e��� ���+g�^H���E��`�����-��ZU\��㓖7|��3ry���Բ.���t����!qsl`���%�I5��#U�Y�2"�(�Ki�*�D�Qp5�?,`v��.��o1�	�7.���"l���7x�N������s��X7�b_e�t�ol�X���7E�L�4��4�^�*�
��$�u��=2���8)���x�! �L�
���zt2�xPFc[uAm0���@+Y��"T��|��N���'J�Un�H
�?vo�Y�����
h�~�|�!�~%��Z���#�4�%�fH\!��+��tQ�|�Zon؇#��a�V��9V�_�k �<T�kB8����!�差�{�Do�:�M��%�T&I�� ې��x����!��	�<�J	8�&�8�{u.I��㡾�P���<`�� �l�P��S��L���V�;��ϴ�3̊���L���
��_�Y������4b��Ҋ Tn?ZӦ{LP�x��4���D�z�i��eB�=����,�a;�(�wS�B�~���s��� G
�t�0�B|^g;I���?�ef�i8�e�
-t�q�~vL��xF�*iR9�$+��#A~5*�ˣ�]3��?ڂ���@=g�CU��.���a���L��3>>ϯ�NE� �ct��B9`-�(ܕR*S�h�L��$k�o�������v�3\���~,O[I�W���Q��`|_�|�8F/�9mt���WD��5�p`�=�r����ܝ"��6 0��Z{Z���n�a���0��տ�y�_u�$���Q��ca�X�x��5����hz��g�T8��������`;�{p���υ9�[6B��
����,��GL�|�'�=$��Gd8/Ò�j��/<�C Iz�^�J*i��vW( ,�)[�{�^���q�u�řK}|^L�GV��A:eO��I�����j�G�Z���o�Qf���=����<Qs/[��؀�=�^�[~0���D*i�U��*��L�0W��+s�v��C�X�Sh-81'9������������2�D��(�a�R�}I��$��œ�A�b*��(���z�Z%N7��Z�'��|�{�ֺp��?����h�i���V�[U� ��i�}�w���Ȍ�Z��('I����S��҅��JD�/d l��+UQM�O��A���Q���[�1[(�Z��#+{�9��jS��b
�r��;��u�l;%i-��.
��M)�@C�S`G��� ��H�L����˙�^N����M�2�d�!���z���N����' ��f\V(�F}dm�f����`��6Rl��Y�b������l��K���bx-$]�F�7X�u��)d[��ȅߜu�Z��6�/��.�А�˟�(��wx��A�;tH�I��qŮ�-��̈�9�{�/W!.\�c��[e&��!3+�8��5��W�pH99E4 �x��NU}M۲ǏIEDFΒ(1���yN��z#mn�QdC�fb��L�5�;�G�yI\q\���؉`)۷ ���w�lHJ�ǜ����>�o�c�
j
�Puj������v`�=ח�� ���51db,����;�|揯4u
n��5p�h����W����Ć:��1K�R�	 uI��'d�(%�kИ;Z��NPN�Ӱ���	�4 �5v�!u�R$�v���$hd����:_:#���6(7�m�,M��������~M�vc�8&���iB��j|�1��[?�q�T�[���I)Ͷ��u�xf#�f��^�F]��Z���Z!�e�,|�>�+�.������T������5q�6����q���>�$�[.��M~��Oq�)�Yz�Cw*�I�����z�9�Aby[8��&�o������
� �%��(t��y�����8T�+�������"h� �T�$�Ґ,�:�E��(U�ӣvD2���ĩ��QЖ5���^�d��i�@�?:9x�ݎy[U��L�4M�_M`�Ii��Ԛ2��l�@]�r���u�뫷�B��G؍����o&��qf�6CaR�Sܾ�/�Ǝ��f�v�R3�A�Σ�1]I
4#��'P�K�#5��=��2���fqm��[�K�� �\�?9�����cCƲaSNx(�hPi/��&�"L���r5���܃o-���S�b���vn�i�њ'�0 i�ν�st5�Rҗr�)�pJz�Fu�rl�V�BV: �WO�/h�k�S�*j��R�3U�X��8�o���Cs1H˕�D� ` m|������}�A4m�BG�M��m��z�@w��N�G1�'�$��Ve�Ү�k�8�w���G�T�Nv�(�[��	�8��U�_����c���o�m�Ph�~�g��AXdS7�������!vv//��uÆ'���6��c&�V@~Ĥ	��^b>�2ԝ�����R]O?�"6ϟM�{Ho�Zo��2W?!+Hn�i���?X�-Q���9�n�-,cs��>��=�qM�a�s"�D�����3�lv��_�ސ��©�kĝ�mf�m'F�9$Y�l����ߘ����;@�	���]a{xZ��OF�/�Ж�Pv�aCq�a����>�x�zb���,�پ�r�K�K<�O��C8�8U*����
$��i�PN�A� iT�Ϋ$�+���PK4�*��1�W3jXp-��+ <甲�F��v�EOa��:l�K���k����z$��o�J��a����NKa��-�Y*���(��Aȋ��LsA�X��P�/�F��U��b!�.��Ը
{�����f��#��
�*"9�ت�����[_�)>������٘�} �p�]3��ُ*���W�
7��	�0*���yD��rr�~��p�An�_o����>}�[$(
w_��r�W���_6��:uhR���=�F)!��lZ$��v�s6�p���>�D��@��$���s(�%h�4�k�";>�8ܢ�+z�
��O�l�ݏ��/'�ԃN�x�nH�f�@���S?���0D5�����s���}WLT�_���˧2��Z/Fr]�u���4��P&5���
��2$~�ö�Wo����5�f��>OX�M�,i�m�T��-�K����]?��s���v�mDE��d�*m���_�����)k��'����)V��F}����;B���|͑���O�����_�h{�$Nh1�[�H諯<�uvA!���`���E!m��2r^;%�'A���Yff�:7�+�]�D��3OA���,K�%�z�-V���Kթ8W)j|js�=gC~1��4YzM���?4��R�z��G�S�gC���m|�h����Ҋ-Tm���A�yj�h�Ǔ .I���	X�����f�q24v�2�mf��{bIm)#��q)!%�b�� P�B��p}P]��v0U� �"yfeY9��쾍q�Ԗz4q)���bp3W0(��{p��\��[U�k�x\g����y��p��|z��r�}�j��=�R��w���Np[���A��0N�@�V����of�(kV�힀�A�o�d%�u�Ȑ��K#�ۙh�$��v%J�����\� ��
���ûC>�ǘ&�E�z.��&a�pd��[;��O��]2utOD&�`�~�Q�h�Bm_^�A�y�z��Ը��X���`0av� ����>no-��
�c-G*������'j ��;d�ý\��x%�5"R��%�)}ƁWF~�߂���<�7"x�����X��]�Rߡ��i� Њ˷`1,���}������� !09�����*7"���������j	���> 3�y���R *���T,g�e��Ǭ�@ C�Q[~�,a*9M�`/�+��M��)!N/�=�M4���܎-{6��2z(khv۲O�6 �>)\���j=����	�D���.��K-����V-X������1�9)���4
����twРԏ�>f��������	1��S�"��nxG�Q];9�-RzύP�Ǩ�O힂$�I�iF�*�AB�sy?�IH';E	��̼��^/���Zj��K�@�lm~W&�H�kQ�-�{�:�p�dm��by�M���,��=�]��,!3���v`QM�ᚾ���Ǐ+����f��mG�ژ��kjX�'���=��J���X�Ow�R��Q�Yݹ�>J�����.�.�}��#a9$>��_�U�\������Ւb�ִF<��	H�\8b�T��dP��:\��bH�u�վ�G%.
�.YV�6 �A����]\��`�SR�7�v�*d���H����fq���j�G���Kr�;~M�g2�oE��7>�-���#`%�{t��O����?��vhKWZ�EqM�I/���S��X���䖫۝���iO��#�h4�?Tw���0�U<"	�7�Q��'�N����i�<g/�5��0����3��#��ƪ�r��yr0��i�<TO@<�_v3T��|#,55��7#:�?��7��]]E��䄄Y�[E���`���4�	��J���lx,Q��F��7g �J����ء� M
P]w!VW`�>�hC� ��hA�����w1"e�������{�z�Z*���8B�J4���d\I1��&�+ �Wԣ����"R;r:WL�2ډ�1AD���֑A{k��z��h�g��)��fR�[�)���A�m'SD(WdXuҎ����q���g��Tq��˭��[�����c0�J�p�����^�/��S	����2�k��Д���o��N^����_�4���6$��)�����_5�����l�x�4#�w��zM��M�}�+JM�$�r�H��~
*&��)ۈR�����I�����s�S��o���I��*σuE�.]�32V�>��{�jI�������4L���H�i3����=����&}�քD�Hi=��Q�,�����C���((��W������ܯn�s��|���⳸�@ve�J?L'��b�PJ�
�{/�5��i#�*�F�N�3��?�FM���#j�uÌj�����	���m�����>H����!O���D��@f9�LP��哋80K/�����1\��c��0[�#U�3�0#��YY�]!��S�p���u�6���<#%8��5�q���yS�/�T�sǅD�F5|:���c(��n��l��?�(�/�i�W4�G1��Oz��,�\�3
7�+�Ȃ���$����5g� �Z{pU�֩M|�WX�"l�wZ;���su���uNأ��i�C�VU7f�M
L�W'��oz7�� ,���?�� �\\�y7\���"�a�:JGt)!�j�������=D�Gs�;�lY8h���IiQ���q�*4�ж�q+ACm���v��C��r-�Ux�	���W����^�Z��`��	��J�?{�L�g��M��7��"�G��W+��<'�z�+�;AA8~�_�%l�g�|��3��,`�Xl���:�d��u,Ұ���ɄӃ�'��i���wi���� '����DM��v�F�!�,������2�mIGA�����~�~ʖ�T�6����X�Pc�C�Ľ�P��~�P�Z ����\*���0k4l��Q~}$�2�p�8$�d�xv�/�7�n���K�������]�����꜂�\��s\sp+J{k2IR髀�ߑ�*XS����D����8/7��Yji,�_0�5]�0[��X���9����wWŽ�����֛����Я�D�_�0���B�c�/�t�r+ez�T�Q��nY�1�*�ʃ��h?�X��]�m��C��}j�ke�Z�c�L��26-�Jͯ�u�,�!�'y�Tݿ]�u�T�ҥ6���fZǿ"�R�㘘�J���4Ȓ�ί�n�0��0+&O
z'f�<�����8�ґq��8	�eu�+�#c��� ��Y��n�k���B��Ոʈ�T���?5�Pg������n�y�V�1�;#���8�C�1%6p#�-�f���;�z�#��И�x��U�嵛��%n���[���v�7X��a(HK�S���/nOc<��e��HRW�h��P�%�~/#wX/�%�(<����	bbcZ�IK���B���yRd�
�����w~:����0���0L�W��̇*ڀi0�p��k��͞vQ�XÇ�XZ��r��Wz��Z؃Ǿ�/�,>7�,���
D�J��_�j�F('F�e��$o�ϧԔc��-�m���+�)�]|g�4��� ��uHDG�\�'C�p�-�H�a���� /�q	��z�K�L�5���/]�P�$�Z<��O�LD���+��Ψ+Y�~
g����|�M3����`�# ������!��iD�29���K�}?����3�����~�К�?[�\��̢I..{ń�X�[Ii>��L���E5��ɗ$����[�T��xkW��� |׶{;xx�.��
�-�]2b����7�
�AO����P�|�����-��v*8`�]��������ZMjw@��ps6�;���w�w�a�W�+�V���j,����:(Ώ���y�#�"�zΕ��_݁�����,!��7�Ѡ��&��x�j��m�D�;�EIX��U^����,@qY�Q 9(�AUQ.y	�?0S�NեR�+"<�cz%�n��Q�}HQ̧����	-í�	���"�)���n}Jj�4�<�$w���ҘN2j�5��<���--��ygCR�-����/;1.�m��B���!g��R����Yr*rє�|41�<��j]h?R���3�EǱ�	=�ͳ���� ��S�/��:1�*=�	��}��@�%M��)�d�Ģ�>=��(����<�,ݩ|�T�в�!/� �d�9���G����b�=��ئ�T�Ik.9q�,��h.��j�.���df����KU� KAۯ�e�A�bq�O�;�E��F������L�;���JSn�k�v�^Uwd�ʻԣ��Pͭl�umΚ�D�tlM�5'�{p1ԣo1d��S�ģv�OU�~U|��"��B��}I�C���O����ɪ�h�S��*4-����^�LvuCl/R8IH�*=�E@�G:��K
\�Hė��Y�M���vD�ƥÌM�s��	���eciR<^[=с�����Q��fo;�-R��^U��=ƼL4�d�"8i2�;�ܗsBs+5Z]��J�L�b�υš��d"v� H �����\��H�+\�c�3Y�"�]w���ۛ�k�j�����������sQ� ��ϡ���9%{˵�>sS�{�3\��ǝ
�T�c6���UJF��F�����Fξ�b��<�O�3�~���O}%��V]�/���<Q ����;�f��l']�7�F�#@U^�0��^~�2Lqr"�\:AkV<}�*��R#��"��Ҫu���5�l�ZQ���y�������d%��O�7O�J
vM��ƴd<��h�0q��5��}i���i���io��h�Hh>�B���7~CQ�M���;Q�f,���?=H#&�/�b�Om9�Y=�����mX~��K��E���@�!�ko� �w^�x�;BFn�UMz��]�ư��%o�Rȗ���NA�vݑ�O4����o��,-D.�U译q�C�j���~P6x���c,�r��`��_��@,�1t��+vB�!f�%�J��t�c��^�-�O�\�x���^<+u,��$��[z�L�s�1U�݄l�X� O�
�r׳��\�K��q�|C+��B ep�UdE���Dsz������b ����|�L$��7|��v���>� ��QשU��IZ�Ɣ<�5�O��$ڮ����w$�ӗ�������v��柝�bڤM]��[�V{-q ��~\�$�`	a��h+��н}��:����G���:�غ����(������}k}�!�f�):kf?cZ-�\�4�8��Y	�	OU�t�vD����'��ق�HO�ݧG-ΠW٘(��	�D��D\s��/l5��OP!���C����l�`_%Y��������9��\b��C�<�R�0]k�2vՓnA;�ΐ�	�'����_)7�����=�������OV��3PoX4d�*��^�$*mNW�Jyˇ�ӣ�n�z[e@S5��&yg� [z��X~��yCK��??�yٱ���#AC��q^����8����Z�xY翎��������=���U%��5��;�\$%.zI�;���"fe��(LWu�)��E0��N���e�2���T�V�����X�j{jA%���^��pc�f��+b�>�.���ͺy�aa^�}�`���FmbO�'�<�t)��Β��y#m]PWi)��fo�Z �(ؠ1�O�c���-	���98����ӋX��{K���O���g�R��dhI��tG��|�fݹ���s̈�g��L+�X����T�p��� ;��)��S/:�����@�qÛ�.���@,'+�#͒4��1��jc���x��E����]�%zL�CvQ|��jJ���
4��%R�7z��ew�Q|�
�8��=��N׏�8��x��ө�@���<~P�Q*|�̆�o��K��\\:�a�l�"�^�=K{=��S/,��_����"����O����\�k���/���={��$ĥ�Cw'��Ԛzu���'�"�X[��u��Q���U���A����M!Y�<���N�[��c�јE��Z��t�x�6����#a��Q�>L��'ݲv0B�ƛeJu)���sQ��*�� Q�,r�����v�/�2��$l��Rl]�Ϫ��I����hG1�n�$Jv�e�z�΄~� ������L�,(#��W�j�N�6F�X�$ȓ�J����?���Nz)E��$��H�c�x�o��WF��M���vVC%B����HgMj���b��������!l%�u��6�y%���	�~��(�T5lk{�> 5����C�a�M��)��0��v�Ռ+|m�[|tU�v�h�UH�����Ԭ2���A���Y!������.qo���V�\y���7�>(��b���h�vV��k͋�/�:��T�3���ai��L�9秃�^[2t���5m�vR�:��"�KD-}�[x	m=�M�ա�X;� Rϊ�,�<w#1�Nen�^���N(�j>��3No���u�?|�+��l��ю
%�����r�}�����cj���C납��w��^�aZ駬/��4q������ ���S�6�_l�[!,?[�A	�v�|���=�!T)��>7P�+-����+/�[+�.r�x ���}T�m�-��yQ	V�6��ӝ������S����@瘣3�V�Y�Q��sD�S��[�&
c���z�#G�μ���)��OGS�h��D��K��ɷ�I��bu-S�W�hܤzjxB�q���c(��߷���=W)�'	�A��Q8é��3�D����Ij�_����,(��Ӵl!\M	b�Cg%{~��!����
�M�Ĉ46+�PQ/����}<��~��K������(w�y���62����4���^"�q�t��`���;��vR���{W��ImO�ɒ�pL���w$ܛJ��X�?�8�#ίQa&~Na�~� �C3�G���g�*��T��Sj���I���ذºW���>�c�nR9�To��U!R��ߊ�T;s�:�"/�:�_<� ������U7\���|��!��d��ZT�H�={-��9�8·t0y2�]4G���xO�F�I�Y�[e�;��4n
�|S��p����f��x%�����0ڮ߁��B�o�@J8��L�6����Ҍ��ڽ��xXl�~�7'�F��
o]1⊂'�wv�p�1��.3ɣ�����(����LR��?��\ÄZ�67�$�5�^��D�z����3�.�v�%�T �2���1H������� ��JuP4e���x
:}��r�ff/Ӄ0�2z�V�
I�Z�8���&��l�>��ъ,{1V�Z��4�׆�]˰�%(v�p<��<4�FI�wKZ�����c�Lr��-��^pD���kN��c��{����c�}�e����I�+>�f'�����D*n{S��Nh�������g^i$�H6]B�#�g3,?�Ґcd��r��"�2�W���`u������\��j��:����;N{��BH"�4�&ۄRV�L9K��z�Yc��� �_�h�ûsd��C�.ޥ����3�t�X-N���mމ'9�������.�z72@���Q��*��D��T	n̉��i���J�7�f���bdD�
��g1)�n������KM}�m.���罗lᣟ���]j��|7L>(.b�UQG=�#��ы�Y�n��o�"��{�v�e��QQBh������ke#�tl��\�r!*����(s���oYmmc�o�+n``Q�g�4@�Af$��5�Y�g�3��/�WBJ��U�s2h���c�S���yE�d^wl��h$�T�5[Y�A�l�,�Q-�ޱ�~�+-���RLR�e-��.\!����e�0�����a+��8��Se]/S�(̢r�����d;�P��eկ�1����{� 4�n ������b^�ƾ�5�5p](�7���d�"u^�u*�0�U�2Uu6`L@!�[� d~�VbE7��;J�i�ȍ��r��2⣢˿�sX�
�&(���@{3�86�q��S����T.�:6����������&F
�V!ȩ�m���U����Q��4j�s΍��/w�ؓ��Yg�)@
��S�|�2�%DMh���\���8ɒ�v���3�^2R0���~����-��MX+��1��Z~��'�@����+o�B�y�j��kD�ffa;��f9G�Lנ��C�Ƿ�' �n����ʩ��ٜNj����>%���c� l\s���Bf��HZ���|V�|V�=���`�j���?�0�_ϔ�K���~�ȹ(���Qt� �+��R0�k���vuߴ�Q���f�F����Tj�D�>^���u�mP��oj8���}����4F&1���1���A{	�x� Sji���
�g<\ǨF�o(�v�P�(�H�e�R������7׀�]N.�3ls���	�h�fX)�C���M�"�r�%f�v�z�U�R�it����������-c`'A�pO�Ɔг�Y��t�,.ג1gSM���5�e
��q��8��
M��Ɂ�﹦t
:B�:v}@���!�ms�:�Lۣ�K`�J���p��
4W+��q���حVF�'��Ex�ʝ����5���A�Y��������.��� �Cx
Q	�*�)�Z�ԉ&�dYΑO�5!���>��}zE���t���-�s����Z����9�8(N�r�X<�W7���g٫���S�\��]��m�5k`J��(��VY�lҮ\�j�N�F�ր��-jzc!�2 ��<�M!K���
�Q4n�DP����N�{^�2��������U�+�MCR:�@����!�%�1�8,��^�X �x�P ��Wμ�F��
GDPs�Hq:�O�Z���f�@BZC�R,��l��+Y��Ǣ�x�n��?����Z�O���P�e9������$��,:�k�=ۜ����"���f�a���Ńg�$O{j�K�=��9�u0ߐ�\z��;�,N&�c������&L��?�.��b�*\Ͻ�XKs�
��;z�ω�ȯ�(`�b 3"S����%���x����Z����<2U\A���񵕗�C���@���ۢ�ة�ܒ��������ɝ.��b,=
��}�H��}��߄��g�QL�:,s��<��Yl�;z&ָ*@��@l���rQ��n2����#��;����R�_�+���6�+�4��.�wc��+\�j|+ԏ�@��� �7��!�)��#��N۹�(�H�4��'���R��<T�ܧ>.�yo����ItR�a9�j�4B3�趲���J\˾�!ƸIS̙(��R.�Y�����d
:Ѵ�� ���Z3?�Ǩ`�8��T�P���f	�#b�Hy	E�^��0��P̈f�a���j^�Z�8�������8;�.d�I���Jl+2���Z:�v�-]�;R���B�3�)N���Hnɰ�|��A�����8 v>�_[�?���I���ۯ���J��T��<LVH�p���C�k_����m|u�OE�M����ߒ����,'h���=3wHj�ː�7�/�,4��3!���1�p�ϥ�%�bK�!������m�ЭU�U��o^1 ��QĉG�7���3oܩ�Lp�S��y���)���V�\I�V�e���u�o��x3xn�?}|�N�����;vD�ErS�Y>��@cϷ|�yx�K���*���A=��f��!PDaw��"�b�7�u<�
K�* ��<��*���kP��x?	�l��`I�6�5����07��4��pK��ҽ�cֈ�����&K�BHF�l�����{\�n�(�x�6�)5��,�oy�C���-S�{#�^
��	��
m�o��W�gOO�9j���.r�~�&	��i"�Щ�)Y�OO��Q���*���S���Љ+�I\ꍌC���'_o�%Y��뇺���u���DT��5"[�{��z<����+�d\�����~s��Ə;���!�	�X��� �BO;�p����t��2S�.��ς�ڢ�A�	���2A��߾�7����c�mF�\��g�J��7��h��@�ö�@ʓC�WGR�P ���V���c����!�:� ��Բ�5�B%�*!�������jb�X��h�Sh%_V�	�PJw�A�:�7�*��qޯ'hS��wPaifh����j�������)����=u��,�n9��HC���H�E��bղ�h�OD%�mZ��%�1S�ҫm�������_dh��ڌ��׹�P���Y�oa�j^����Q��[��XL�7T����<!�*��gWdiQ��W�[[Ө�kDp�s_���CQwa` ������V{��ULY�����b=2��m��w,W:�ed����'Qt �|p�\ ���DKǜ�1-�1���<���+�jg�j������2��ې��2�����̖%_8MoyA���	�|�]���<�w(�~�	�6�lK>�㿄� u|ώ�mt�^q0
�1ԓ�Њ�Z}ӥ/�Q����0G�Ό_tU�5��k��M� �:�t�Vb�6v�Vs_���~r���譋�i�Q=�(u=�Y�s Ħ��Ov"qE�(cv���wb� I?ܤ�;�l��b�.{��/3�Ϊq�L�;L�nBDu�\�:%���i���e�*�����1T|�h�6�nor�#7�q�i���)	��/5J㞭O�t�V����<!��5���ȡ_®g��i���oDf�e��ˣLML���F��m[�_27���5�_�R��EGq? ��� ��0��[�u%��c��&K:��"r:
�܂�G�z��Tz�����gE���b&�0�>_s���u�����g�)}:�@zg��C\:&�$}<���-MQ� ��ġ6�\5��{���q�=B3�hX��F�~�'O�	/!�N<���To��;�|�4w�r��x��<��Se�2C�V�|�������H�wP`~��3q5���}9
U;�a������ ���6��b{]}������~�lǓ{����
�:���9%��_/�]@����p3�Jޯ1��8r���.���+�p�VS�(V�����'�ԫ'��w�tC�kH��ɲ����[���i<e�w���M��.�S�� �zͺ�,0"1�S��m&19���c�ZTǶ�ȑ��B�˓�����p">O��u_����xS����=0iϥ|��q�h�R��&�����"�M�]�t�{����#�n5��B��B��q̓����2T�H��{�^�!�R�Nڴ��.��	>�nɿUK޼��D��X�|������(���n�+�AC��WQm�,�u ��$���q%0��@��!,eC����m��'Yr��U��%�Fx6�q��I�����´\���Z �s��;��y��7�uuc��Z�ew���g�w-����p�<��KRO4�wg�I���k��R1+x�l����	p�\׎�辴'Di�u/���xW��P�����&fӱ�"����vW����=#�iH���]��F%�$�?���t @��D|A���73��m�Xpc�y�F<�:�U�ԜƗ*U"��G�]����B7�Өc�	� �5�e^Ge]�c�7� 90w]d�V2 ��?�
l�����m����]۽�� �g*�>�4*�J�(�޶��$�DU=�л �k=�z6�V��PL!�e8�8�Ə�߆�2����oZm��{|Zd��)d] ى���FWc�`����Kw���F���V����@��m��數{��=��QZ���.G�Ez���D�'Ӎ�h�>!t���5�Ɵ�~�&b}eE��d��P�t駒�� �����9H�60�+���Yߨ_*����V�VN�<�K���̼��{f,RݳR���Z�eΤ�Q��:h��~��
�@ķ�'"�C6-n,π�"e�Ali-9�w�o�ƈٴ~-Zp�'�?/J0���q�Y6+8,����B�Y��Rʥ��+I$�pԅt��TS��s(6�Y�&��78{n��XU&�_�lPA3k^[9�vڠO;�,����������ݶ`n���W�t������v���9~�"UW�����>$�, $~�8����D�P�����.c`@����݈��x�
�$ϰ��
�cj)�5�gg'Il�b���U�]7�oIU���/�Fn��)��/~��3:�q>e�/.S��^���H=@���v�j��/�$(��DݜĘ�?s�9����D�{�k:w~�g�� b�u������E5���5v օ��+^Z$��:_ƨ Ş�`�������B9c����%F@Aa|L,윽�YZ'7��������+}�.jOӢvI�MT�%�O��r�K$��/�JJ��!�}:c罎��fJC�_�Ғ��<����B���Ħ w��s�4«u�y���B?ɐ~5r"}\t�!��2fS|�0��.��F�Y��F�����|
���#���lNyY�յ�̛6O2t�]��m"hUӲ^#�
��h��Z���Ң�O_H����W���C��/��d���U>'8�eWAN$����(�D��ĸ���+���mSk��|�dp"1�V�{7%W2�d��t��ݸ�uڈ2��O~��T�(vq��cW�? (
��<��n�Z��tZ�z�7Fo>Mmxv��d��R�v�59C
��uHG�#H^�����&�}K��tE�)���&�	> ��2�8>��%�^��#������UXȏ<����QQ��;��p�/�S� hp@HIK�{�OA�N{L�X����BWU�ʈ��Z��)���[�s��Q�i���W�'[�+t��$�(���b%f"O��f�N/�믲�c8��Yy튒
3��4�:�A� 5x���ON�A�%H�ܛ|#T��z}�8��.�d�ժT��ծ`�C���#=�',&����a��%�V���+������_�X���n�gJˇRphɡQ��@�[�{��N�Ɣ�G�k��I������C;wo��A'2Hz�ۧx�R/Yv���D���;`���e�屐�':he�dM�R���z��z���T���kœ�������J�4��]ʑ�6�7��}������d��_M�c�
�.ik>���e�x���ռk��(y�ˬ�ؤ����;���5����ewsT�q-�����m�yh���2H?GV��3��U냾�Y�le�
���(����C-�3»�Ra�
z���g �p;ψ�y�>!_q�>y�c/?J+r�h���Ey�����,�y[$J �eQ|��i�#Ҡک���3^B�|��,�ȃaں��ΛV/l�;y4w@/�)@8!�m�).LH��R<>�'R���m^ƕ� ���4k@����'e��q�(��c��S��\Ů�)��MS\yiЎ��2ۗZAb����a�V.N��B����5γT�9׽=|{z��X��4��6}���IՠM-��):��A�J�N���ʡ��� Nn�#0z2C؜���4��l�/���齱J�Ì,�c�/l��%���z-��B<���\��ҥ�*'��q��>��ɉP����zx1�5f���$�b>0�U/?�����"恒���фE��f1B/+�5Td�@b�w�vi��7+�vd{�8 �z����5C��.�ޜm��>�W�����Ljx1���D��T3��ާ����[�9i�Q-Ԕ��H�d,+�N�L�$T m*_T�\�&s�'p��C�X����ш0Ψ��Cql1ȓg� f3��[+fBf
D����ʝ:�͈[��t��Y��|Oh������3
�;B���g'=� ���Ӂ���J�G���?-�IpMve���짙a�x��	A'(�\�kc� ��1N����Aqu�����+�G�,≌���M�-/�yD���n��Fa�c�>5h԰��v�T$��7ys@5�Y�����	�$��u`��� v	i7
��[�I���ǀK����O�]!+|�q�9a�B�J��A�Ƽ�ȼߥ��q����ט@p-����YW�B�+��<�h�xZ��׼��Lu�e�)�:��!�8R_f�O�pZ�dZȖ��30�������NL0`N�^��**����ҞI/�2D#TՀ����}��yT$�[�@��*�U�*��uB�T��
\q�ߍ�hH!Z�~�(�)Ib"����Ӏ�$���Ҕ]{�ܸV���]Q�dD�O��=�V?c#^����yy�o.AzT�%(I~��nE,e�#2T#��@^��.�̀� T0 "|��d��-`��¯��|8P�r��@HM�������=�m��r܏$j�o��}��������-�Vq)uD*@�"@$�~BG�~�W��O���+ �Y���۰!hC�$�~f_��L�)�L���2������[wp��*�F�3]I�X�W��E$�{e����2}��<k�qi��<�O���&,c��2�� x���0�H�n�� ��?G��2�_S5��/0h�{eO�Y����DZ����}ý���u)��72�hָ���JU!�b[�{9T��H5V���Q��/�c����O�l���|ң�?	��DF�O-���P�hio�����P��ڌ���G��Vm�|`R�M��ޤ�8p��Y�s%��[��16�ˊ����F~���h�[RuN�odS*��)m��cn��.��Ȥ��KY�k��_B��/�;�8�}��w#ӂ�MN@I�[:.��O��nj����5� ֳ�@K�"��A4�$���z4��_����ڦ����Ӭ�b��8;RJ�Ll��j`Y59�{���Ϫ��^|e�痁Jp]�m�keg��hs�;W��f
�����L�R���^�����tY���5����"=$Ι)+^�e���q�vv���[`܊�W�ɏ.;JKFك0�ɆQ��y���v��f@T��lg�$����l��	��ʿ�*oT�\q��	�"�$�����aA�Bj�:�~l�1�\���
�����?]��j:�D>����`tv����j4!��;i�6�B�;�%����\W�/ጩ��B�ZY�r�'ǶО�����-�Nú̃����W���h%/�p������>:wou�4P�h���9O&�!v^��
N����FQ��4���W�2�7�g=ĕ�d���y߃�e`]�;��*�ԩ~�z�f>�"(���[���
#PjFcH�{RK��!�{��sV�,h���b���^�z�����-�����xz��
#�%���e���7����jԡP �*�.�hY�Wb�)����??�1�Zx��oj�|[+���˥���VGf���Jy�z_��T�P;��,�ڳ���:���Q4#"L���6�P�Tn����L["ū����%��ń0�	AҀ5��1�jok1�<����H�g5O��X�+� ���|��i��5f�6@I-E=�yzZO��J0��#żmT��*�,v����u���&d@��<3C�eP�?�,�sP`�*����M^��y�����D�F��1�9|�1*\����:��4����KXn�M	��2G���ja�y����l��0!��ݿ(*� ����Ԡ�����x�H�h��C-��/ �ɂ�"�	���#r?sU��]����s�Zb�71�eA��׆	�`�����5��2�xL�)�{���k�k>��9+|�^�����zaG��xq��x���P'�#.��/Δ�߬�i�I���a��`b>o�F��uD/��d{3��߳�=�A�H�NPu���v��,�wC�ϲ؞�����'
����NI���Ym���RIe����?(.� �]�`�m(P����Xo�� p��@w�\�z��Q�{�c���>6�l�ʂ|�9#�z��RD6l����^��u����n����}ng��p��0�)��.�l�7+M�X�����$�T^S)�S���u��Q���^�^���$��e;��� u��v�����I8Ưs�CIw*�w�{�X�S��:�����Z���$u2Z4`��}�����w�����f��$�P�ao����T���K?c*:���J?�t���V|��4�u�EC�ud��s�?l�ŝ��0I��g�p��מix�oN4�Kԧ\�`&���������;���6��i�?%��J4�e��n�_�C�� �H���Ɩ�-f��IG[�`�2�t9��{�D|7?�F�.�����+5�P�ܟ�}��Y�yBPy[�_�:#��v��E��*�/���e�\�>-r�H:⶜L�p�k�yP��;�II2�D�:l���2vW<?��jnU6���6V6�3�3Q� 僤��̥�Qg ��٭��H��d�͎�����F
ҙs`Sz�����b���l2+����+G'}`\��hM6���]�T;N(�ն���+��C�%ɷ����d5lr@��9��3xZg�:9��G� n�1��o����//E ���'.R�Y�{)��B.о��-NS�1�H���s_T2�ퟛƶ�z���� S�Cc��ga��q��N8΄�t�/V���Ȼz���k�S�/��R W5pWg�{�^�����@G��Ln��Ȝ0e�)����'��#3Qɔk� cL��隂u�gqN�-	�M�I�H�|��>Ja�׷قgv���l���Z�"^�ѡd�.D"�*��#Gx��&t�^����t�L���6}Lx<~�J�ӥ���ؗo��-�m+�I�n
��)�jɒGJ�/--��2}I{4��T��K_�Ӟ'���g��5��M�o!�ɲjH۳-�@�����n��Ol�;�Ͱ)P��W���v���Z�\�x�����)adp�p�$]L|�g�UWn��*�?�K�U�0e۾ Bi��Ei,?��N��mܩ��v��+�<D{'�S�	��Z򭥖�#(]��ܑ�k��D�CPoX	��L��m}���2����I7!W�ޜ�+)
���=5�R�P^�����y���,��?^���+m3Ƙ�j��_���U���_��z���ڬ�^K����G�v�kzW��D�I�RE�t���T���c�=��G4�3N�k�Q�;auN^�S����o� �%��.;�s���t�x��x�HC\TIEgBۄJ!]�p�VC�?4��l�
s���V��Kc*���T/[�'�͝p��q)7�7�V�zX�r	��䟣Xޭ23l�,���T��v�ę�G��R3	%::��ǝ������Ws�W��R���9��Y��BMłD�Mtm�����~h�7�Xy�E�I���5��W��+���d� D@�����B�E��]\�8}-��B��O�WQ,ˇIr��o��_V}�7�x	���ֶQ����)���G��2��03���]O�hcd���řt.�PN�x�3fqF&������}�^��rxe]Ο��7��O
�l�̣G��tW�#.��;#��-�����#���'d���1I�ԇn�c�d��K����_��L�-,�ϸ���m�^4vb�U؀��I��C_MP���U���3�Җ����S���R� m�w���-���.�����˸��䛐wIlT?��H�۠J�L���m|4�ե2:�o{�ƙ�������Kb,jup�����BX)��q�������~�B�^;P|DY1��ΰi<�$�(��.���p^�߃�kt��-�APĈO%mI++/̪{�Dc5�h�bG���I�A�O-_m� �b+��(�&�ӆ�\����5ٲ�Z��u��i����+��G܋�Y"EZ�G�]B5x$��2��܄������� x�`'�]eM*�x|X��ÿ,�R���/�����Lѝ�ٌ��z�3�	��%{��./��|%`�}�ӽf�9J^�ú|��>$��^ ���)Q���tKVPe�peu7��9�M�"^�s�P=�\6U4)q���f�8����Z �`���)��xq��eɄ2~���4��Rb����&N���\́qg��E)�2l���a�p�3RտIX&ڭ���& A;�k�Vi}��yM ��y�B��Z�$a0�D UD�9
�eо�Nʗ�0�r",���≟�ߟ��Cq"Y�`>�k~	�v�MG�T���m"^�4���=����v������B��
ю/?c�b�~��'��[��0��T2�C�"y6~�K>�^اg?u�S��}K��D��=�� 1"2.�56����'�>n�̙����b�Q�"�D{�4�,JgO��YX�����(+�,�\f\Y�Up~��V�͘c�[�xฅəQy�c�TS������c0бɜx'M��z2p�1@��Ac����68�1K�����/)��������z<)N֤��8�&�R\�5�4K3�Y��Ƣ3��������t����ʥA2���ִ��ɸ.� *��1������a��V���2��˪8��Ԅ�* *ZШE�Pνcrۂ�O�[��S�<O�
\� Pq���¬P�s�@'}���1|�z�%n)�;s%X�4:}������ۿ���w�q����jj�#��H|�'��6�t�٤�G�ߏ� c[�H�BD����恭�hvc��q�����tm��#$�~Uc�1-v��`o���4�".>�$�aeU#�U2�@��pӝjl��g 3��1c�����Aଧ_����1�{B��~w��D�8��3�L��#�����Y�q���Y7)�񰘢�U�K�qЦY�GL4S�ee��z�!�+�0�*]�W��8h�<�+�;E��XI�g,X<d϶^��J����o�h}G��p�E3��L���"w��N�b��W���E�ʻ�N֪lxY(�{��|��b�z}���)Q}2����N�^����E+��."��oy�Yn.jr��qP�^Tܶ�>g<��sX�I�[�to7L�Ҥ;!��݉���I�k�z[-)t�7B�fx����W�u>����R9uy���]�Z�*y��匹�Y����@8�\8L����������1��{�p�Z#�'5Qe�������g��p7��ˊ�Ut�*&���o9��Vb�X3��:�����p���2��Q�^�5W*jO�����l.fp;��G�FV��Ln^=kK�PN��+C���ۦ�N�l��B�����|T�a!�J_���P5Չ8�4bt�����0�=��Oχ�M��מ��
��<�#����N�3�p�����$�&&�W�
�D�/;Eqy��?�Ò�ɸ��Fg�P�{z���2����҅|]�<d�����TrֆxЄ;H�*9���r/pϰ�,6�l�?o'qb$ ��nI0
�h�̪�}�7 <��`�w�NwQ�jX)��/�R^p������Y�� ��R�V�3���A_q��t�ҡ�F�?��@�a�Z][A5:S�����=ݨ�GpF��
�2ڙ+|��@u�h��)�>F1i����9�����<� 5���;�rk^��}%%Wmh�O|C��U�|���9��w�f|t���$&N�_T�H�(����%��Тl�ߘ�a��o���YP�]̧/�����|*鈮��!���V�N�'[�!zڼ�JKܞ�"o<G�\��Q)e����A*`�uV�?Ŕ�(�
��T�
8	�D��a\Tݘ�{�{���KC�\q�5��n�U���ѝ���x�з���n�Nc���o��r��=��8#����,m������:��'^I]i�|��oĳ�1��֝�6�d���9�x�C��K`�}���C��( P�����8����q���+�e�"��ݻ�ǆ��/���B���E<w�3��_�ٙ�K$�4n�5�"wM^�iƥs��ie���r;�]���"�4�$`7�ϧ��8)C���|�7)`��9u�Tb�U�fQ՞�u%D%����O~�"��~��"z?j'( �sG�8Pc���+�z>�� �4��0hU(�忂J�����<��8z����>���P(���� t;2c}N�@oq-i�4(��Q�e�x��JU���{h@�)����+"g���@��-�#�]SXg$qq-��>?1U��S�$q��ԋ���?W�N�#�P�7�6�zR�4%l��>g��������i�֋����u��pe��)~��ě�\A��zY�O�Ȯ6|oKv�0qw�3�\F����/���ax
�K 3��o�k@��N�꦳7?ӓ���/17G�H��ҥ��{y���N��4y;������j-YN.��-�x�aZٰ���ߨ��M]��]���3�'��/�-9ҋ��ھ�>۾�SyL+eڰ��f���^�ѕk�ed-�N���$�HȻ����d���mv�s��������4��тd�<�~�	sܲļ�=5:d�k�����\	��7su�&��c;׫<��3J:⥝Ρ�INUI8d�s�P�:Sp܍rF0��BѺ�3�e��)e�Q$�ܕ��H�"���͛@��/���z�ho2�Y|X������b��;tg�`��4f�Ӓ�xO:fy��8�lt���]Eӥ  ��]{��?<9{�Rt<:{�Z�Ro�Ix����L����8����ϕHZ!�7停¼�+5r�tC�9�grwXRO��_6P����af����ˎ�{|g�	��֜˅֖�'Q���n�J^V�㛌�� �cGP���%��ڄ�����/���I���iqw�����zV��䖤�LI�Iʡ7`�?����FD{7�إ�ۍ1'�������!ؐD21�{�T�D�׭ �t�rAl��B+%�	����)Q���*	%W�E��j橳��Z\�����'�MH�.\�u(Mf(��Ԫ�y�%j���}*�r�r0���	�S������5.P������!,A^���B��M΀y��|&N~�H�3K밤&6��,h���4y
���Ƹ#Y~n���CC(z��l���=狸�H���h�Z@y)�A�r��H���V�t�=j���j�i\mr�@ke)�����>qY?�?�-Z@k�D]�?�<���q	!�EŒ�P�r���I��ۍ�/��P���W)�	R!g�}y�x���K)����1�G�+I��ٲ��]�K0zb��s�����f"��Bh�a\t*m*ZbA���&8˿�$��H��_ۙr��y��!}w��Fh5?Y�	]F��xĸ�p$]��:�#�AT[��9v=Pz ·Ɣ���	KQQ)\�1��@p#�!>>�7��oys��B��Np�'`L@��:��#�h����)/1I&t�J��9[j�wا�2i�V2��g�����i59�	eQ}|�#��@f�/��r�s< I\t��~��2&3x8���>����Ԗ�κx�=]��Qa�%�?��v`"��z�tr�gnu2��%&�ħ�XgKt���� ��������Aˀ�vT�w�V�l�uN�ͺ�L�E:oak=>���Y��\�0k��x.ja���R�EU�nZ,A��b��s�Й2QΞhͨ���.م��A>�&0{yTj���ә�sOrueN0aM7�F(�K���Ty�ߥ
� �@��mm��^:��U;�i<&3��2m$�3����i�Ϊʨ���7�}�Ԑ'cPP�2f���F����ε��Cu�³�U����.ұ��������\�c3Գ����K�3Ok�wl�##�P��L����T�
�ւ�T�4N��y窢M��,9�l��0>��W�@�`�j[f/��1T8������e���z��g��'���>�<��%���S�ۥ]�x���ma�R��eu�i~�ݓ�;h�%�QzC�u�B�<@�x7����)�a.�J��e�E�~R	����m���4H�k_p9��R�Ҏ�cL]�+滬���T�0�o��ѝz�OQ̹ũ��A̖�h��|�1�wZ�]a\}�ݠj{Ǟ�Q,q4��-��8NX }Ƕ��.��ې�da
���"��Mx<��q�TE3���a�э�r����F]��Gy��8�CS\�2B�����y��{�����kն�Sx�(���&�G	`���/��Xvʊ�!�2�:���/Cv�q��k�՞�Lt�nD8��d�K�FE�I�"&��AO;g����F*��/s����RM��o�8�	Y�������7��R8�@�z����_�@<CrW�����[ m�~��(�..��%�t��@�@����C���Y�{�d%*%jk�)O�^Zd>>����i�a�UBV�w�nf5HY)V�	q���hn⠄� ���"�i�E�"�Is	���R���r��%����J)�v��3�bd������`�+���W��B^i�Ǚ#�H6��R�on��B}|���Т$�!;��<�4�z�Dw�d��F�w7>uP�PHd]�eu�Z�Ɵ�jԣ���f���B���ƿM�;����%�y�y��ά�29A��g晑�p�B��^=�j�_(��n�ie+�*�L�(������($%k�_�^�B���jL�=�I��}�� kkZ]�I�X]|�k4��3� Q}M��=[\j�i_P���4X��hXzJ����wb�[�#[@���(v���-%�rN�ӟs���w�
�S�{%��/��I��r���7'T�ǯ�,�"	3�Y`��|Z9��v
Y�y�%���T�� ��\вi����*�20�~8@B�#ֵ�:M�ǵK�TCL���n\_A��A�@��/���M<�o��%�4�o{P6[C+c�"װ����N���� �<�lA�@=�c�RbX����r�&kb�;�����V3�4t&��wB|vR�/�"��?y��:��=�K�x��J�T�̤#L�e�1���@9Y�K� M�ݦ�R��yiT��;wח�I�ۣ�:��>��`�?��U/3�~q���丒�mR�ہ��������19�q;� |��R�BA����"�'�2G	��q��+2��W!k�8����K�\h�%n+rc��a�٩�K��&Nk����9��b�E�P���PI�1�{�p��ے7]+�R�+�u�+�&g�\.�ֲ��zE.���r���Ϸ�Uw1��Pe��B��l�Ex�G�W����e��B�0�q���['Ho�BR�-�_y������z0��f�p]kH�!b`;-tS����e�71R_S>����Y���x� ��R�M2�Y�9��6�G���L��*he�ŀ�c�Ho����j�.O��{X��������.L�=P�0��C*{��:���F,��/��3O/Qcݵ�C���a��Q������Z�ۻ���+������|��B
*��{��Q������O���l����j�iב:v����:�Wd����go�~�׃��/�Q��������3���J��0��2�r�4��P��b���F�L��eah���o�}x�,����K�y�&0���q<�CQ{f%Ax��k|8�Z1����Htj޿\��3þw�,ô�`?�!�d&u��u,���a�J;�V:���5c��2����-��qPU�[��fT���&'ј �զ�h�2��K��r��Z<=�]FY r 9!L}��ݨ�/r���ü�.0��X��HҖ~�q.���Ս�� �iT��LW;�8Uf�>-}Lc�����ȏ=^"H��Jp2}j���կGr�۔8��qi����T�M���K�d��ӌ�����Q�\�Y�q����2���q�������`�B����Ŝ�+F�zZ �h���L���fW�I�� ��V_�5��;���&��נ�V2���Sz�Ϟt�[����-�Q��)	�:�q��2KЎъ;����<Xn�N ĈMj��v@Qɽ��5�?�7��5��]V�;�=��ͥ5u:��@�b�6�_�-V���'���1^�ͅ#��3�y�3� �z�̜�Y:3�Q+���B�j�Ĺ�$��վ��_��pu:�>�&wEzI�.�7a |�Ǯw3b6��Q�'�F�g�#u���݁���M]�s�����}B?���|!d@-�e��x�����������݂�l,��/o�$�3%��Q]429/�����TUw��Щ�����=ET9Ny?���R��Ux���y�}���)�c�
��!�h�j9O��WN��)���L?б��>r���I�I�؏]��^+�����E��Є���υk<��4�v�IQ�����:��:��ÁZ~R�@�q�SEz���|���O�:��D�t�~�!�2��f�s�Y|�E�y��ו����yA���j�u������%`J,fkO���i��!<���/��9�.�F};�����ѫ(��� ��G7��e�������i8��&zUl4)b٤n��|��4�d�ޠm1dQ�5И�9J:��m�������4-k�2�_]���� 7Kϑ �m1����!L˔
��ݮ*��>GJ+��#%^�rȿwЍ�i\�9�C��W����R���L?�@��c��)��iD�$���bN�0�JQ
�D��c�t�`^)������^95���"���v�ۆ���T��FZ���$�O�'�E`�"����I�������bda�-��bn2�@!�sƬ��0�UApU�F� ��dt�^3���(�<�˶M�H����&��"����r�l1GA���O���U�f���\��j��b�%,yC\a6���7:
�zw�
����l��@T?'���aigC���n�|P���2�������$뒜x��t?�m�*��W�
��0��/^�@�]���(���,1o�/[�A�a����k��IfPt��Դ���bb60�2ƨ�e�7_ѴB"t�����ږ�j���&�}K����5��_=, �Q�u+�-�����%2��5Z��1��/���^%W7E�"#�Ex�M���)/���5��V��N��>A��?���Ҿ\��-�ֳ���M$E� !:���5e�����ֺ�{K���3b���o 9(L`��tyQ��������X��%�X�Z׾T ሂ�#�y���I�AӜ����ь.��%!�#rм/J���v�#��F>���������i_/���|���� #)�Ǎ��赖3<�j�h��+)��Vu���Gj���l�`����v5�l�x�A�'Qb��0���¢Wr���#Z�2��cF��r��X�6:�[	��v�D�m��p��Kh��I@}�(��am�1�Vi|��JI� ��9�6zz�#���|��o������x���%0em|�L<��|v��8"l9�Z��CH�u��!��d|�FU��e4H�=����cu���j�������5�����+uzDL��E8lp��NĜ�V�S��,���4p����d3} ���r���S���$�PqG)݌*�Y:P�~ˇ�U��Х�\��Ib/J�JT��	|���'Ylh��$�tp��ܲ1�$�O�o?a*1P�ޞ������m��ך�w|\ql��,7"a��C��c�z L/�N�_(K��G�:Iy�n�" T`�N�)gd��5�G�>4T6ӵ�
�f�u��wS`���З�|-RUy�kY�"=��j� O�Jղ�iE�y�ZM�|�5�,v>/|ۓ����\u�%6_���hG�P���P�����
*	���^|�N�|�wA�W�S�X�/
=.pl�N���B�T�{h�뷴�{Ԍ��c�>4s&�����؝�sK�E��D߼������.e��8�{�=?�p>��TsP~�;��H�`��4�>s��Q\�
&��WlE�`Ixw�>��9,��#̘�
U�Ǩ�D�tO��N=	�O=�!)�k�W��@�¹����Şw�Dӗc��q��]HG�S��.��]�'��D(�}���[� Kx��wSo��`Z�[u�^9e�,y�+�U���$��B���I�/�
��	�`?����5�a� kt5�.��A8�&y��_с(�zO6&/���Us+��4��sZ��7�/�S��L�+������zd�f�ؠ~M���O��p�e��c��������H�����6�+�9���9�W��<PK�8c�S�i8bZl�_r5���ƀ�ɨ?��"9a�Kv�&B��������4��Z\2z1��u���2�a�F�����X��f��k�N9"4l��|��4I�l�,��L^3��KTdv�rJ��@�?"M�������k����GE�ъ=�Ms��$>�A�8��/B�o(���1>��w3Br	��Y����fT�CD*xl�j�ﶥ�%
 ײ��͹�p�� kK������-�� �!z���!�����d������ل��]�u���������3W7�Ē��=����TQ�1��5)�)��KLqw)?u�����y���W�qA�M�"�Ǥ�m���f�ؕ*df�ܛ�A��VmI�Vu��>���R�'~�����ios�w`��B���(�r�8��{�8���?��of�X	���&�������C�|?*����ݫ���'_�J�>�t�:��$���|�)ZVVy�2�ệ�PC��a��9t+�Лh@8�T�ȃ�;8	�ộ5�~�=�ݫ1��ۜ8��X�%�����Y�Qf@���,��˅S�]d����'�k�PTgb�P�_ư1��_�F%�x�ˣh��2���b��	9M��1z�H��J<[��F7�='��(�.�b�hc�u0��������Z���U
�9�MqU�K�e�F5�܇��W�O��#��$R!"���܃�>!�q,�<A�⼔���鯑a~���Y��oD��I�璠EIč��T����L�!\s(��d�Qdq��j�����8`T�l����$���h��`YJ���`���ᅀ�*����]ݤ��&��/p���e��v�̈We2���E@������aw�	���W|iq���=rb�C�J���6ŲrήkǮ9uBF�W���ŉ?���m�8�����2A�4�N�ō�),DO�o�D��K�æ�cm$<�e�����Z���
7��m��	A�5���	�|e��&|x����%04�Ȕ�l�ϯ�Xs�Q����a��$�s��7pVA�Ka�= ��:��@�D���lQ+�k� ���R~�Ѳ8CVu��uɒ.>k�$ ٖ����]%�2�1���>������� 0��\Kii�"B��&�Ќz����$6YǱ��v}��s$���L�O�:�<�Y��y����&��_l�!^?�d�^��T�@��9��p,��h�5}�ys�l�߹��<#+�Q+5���R�E��:\�ͽ6�V�S��ݵ���
+Y@D�'<�t�d���2TӉ�r0�ӌ���ێ��|.�b�B8�#+�w��r|���b� {�.nipa�V_+����w�q����
������e4��ɽ�l���mG���Ж�ii�'IG��C�^+I�I�����d�Z�Ԭ5���r՗�22��ܑ*�` $���jX{Ç�����O:���	���{��*���:X��5h���M�.%����O�� E� ;��\�)'Xv��¯.N����?��|�{� S�;�D��E���;d��$ğE'b0�����|%VW�ws������=��d�C�5	؋��ez�i��4a���o��ʝ��6'�u��P�Ⴜ��.`��ry�q
^O~`�;�`]��'��fnŗ81.�.o�`a�&�v������:Y7.�(��_�M����+����V�/H��,V\���H8s�7?Y|���!����+��0�#	]9i�L��֖;zUtG��|4�&�{z����)�N�j���Ǉ:�x��n���<@�e�y���T��զ��qS[��!D{�oC� ƹ%p<�p;�!]��^~Q>h��%�e�l B��63qb%V���T�ِ��Ç��l�<㎪�sU��0m�Cd:�.��i`S�~"��5�YB���������p35��E�U���]+;�"`/"-�j��oA<'E�����ʏ� ����V�煈.�*`lT-���d�+R�F�
 ������%~�'�,�jy_O` \����Ld�8m��i��}���_��g3d�C�R�薂��Q���z�0�(��C�]���4|��� �O�%��'�
&�g�� 6 �1_^g���.��@ї3��,� W�!���g!���ֈ�DSS�'�×���wB�PJa/����\�%�����Z`͕@�%j��01V6��&;@��"I�������w���R]�������3=�@BβX�t��
|z�t��8�8+7�g��e�x@>�8o��a�eҁĹe$?bS�\h9�nO��fɣ��ѧm��e���sIg�ڻ��5& #�!�KʉC��ˏ����B��"y�. ��
�|�,�X�V�XhM��AǱwCF��ۊH� K���e��Bv,�Mo*M�d����2��5OU�~�id5���Nq��3�5��1J�B��d3{=�M���	=�U���� �ޣ9�ƙ4�A)�4�e��yXI���1*oJz��'�x�c%��m�F���kT�PJ{3�r}�M���P�0U?2����'��Xo��
���"�
©X��kq��vepU�1(��T�{�^u�[���s�������l!��c�K�11�#Rҕ+d�X�
��ķ�[�jǷ��@h2����٠�
��z`�m�p���ViT�~�������]^��/E	�׏!��S	"�T~���2���d#� ֋!_I��h����%_$�KJ�D�����Q3[%����6$)edV�����H�G�"������_w�93Z�d�&/G?�q :�l�w���Wz��b�VN��GY�
5  a���዁�=w}}e{�I���3�Ίfy��t�l'^�3������1?u�3%o`�.��w}�X�����[LD&{��w�{�V6��k�zS��ރ�Oja+���o�ʱz�G�5T��f�ϣFe��:���@6��4Nv��lRd�l#��*�z�#����7}��g;�y���(���(l.�?W�{�IN��E�"F�Qw�Ϥ��_?�&-�!Ir�����ֿ}EP��cG!LI4i�>3lX=o:I�Ǐ��6�ks^�5ubAm�X�J����;B�-Y�g�QLdS��=d� �n�*<?�*�t�bcs�ox�ڍv1��-��eF�kb�}��$x���_���^Ҩ�0��|�.��ٙjL�]�!O&W�S��tp���(.V���
�Â�g�E�4��y0�˰�X��=!U�xL��-b�iB��t�L��k��^V��c\%�gQ�����g�`ۺgl����M\�k�*�Ƃ1�V�;�t/�Fu���z���o`�ٕ���2�?����5Gb�>��Ⱦ��6���	E&����&N-��Ӭ����FZ.�L�T���`�j΍������ ��?�I�GS�9F4h�p-E��^�(Yj�Y�]���AB��@�1I5��!��3�~�����oc���9t����#��V��������`�OВz7[]��6�v�(Y(�Uڢ�=�ř �I�z�i[��Pd��V�3Lr�ࡘɆ;�O^���b����ߛ�2,4U���XK͏!��B ������O�uk��24�N����ͧ��T��*����[h/n���ɛa��vPת�1s���~U�! �Qt6�D];�$lC'D����Q�/��d��x`wy�{W��X��WB���}0���f��Ҫ�г�tJ�$�`��)0#Q4E���B�V]z�n����(�Y�!BD����Ll�p!�!�+� m>3E��אr{~��ٓU�I�'­�HY���@��M���ܵ��
)��czWJ�]��Rf������tǧ" %ֿ0g%8$*��/n��f��&�.���i�]��wvM��&����_<�RH��a-��i���o�&8(���,[��F�
�#|f���yn�qF�2��9�z\�TT�z�>���b	�����|�������]PȤ���g �q@+J��1��� �.z��̡Թ6�ѻ��g1H�	�g���é�ﴧo���D���5�i�;҉A�&3(��E��6S�v��3c�L��2X�������0Z*|����Ƣir�v�ʞ5s� �{�2%�rX���NPצu��롰3�HG��M�p�"/�9B��S�q��/�Wou��|��)�q��� 򈔭�T��]���d�q���R�n�t_�o+ᓃOx��)�CG�x�{*���V�����8ߐ�!�0S�aP�{g����j�"P�DV.9�|<�Q���ӱAs�����Ɗظe�ݹA�w���������E�B#V��>z�q�2�40t�0���%���f����!S[�:��s�y�您l�;�W����>�	Xӂ�⻔6��O���۠����i�B�n�o��5�Q�9؉A�T97�j'n��aR3T��-�s*�}��X�k��μ(}�*}�x`�R�݆l·h�58$fi}�ԁr5@��&��0��*d;~z����zplc�l@+C���4s�0,&��s\P�t$o|����[Eb��cG4�����*��q��v�F�!���qÀ��#��p�@C��^xN�H�E�1�d�./���h>�H�<�0,��ZrzRz�O-�����$ߵ��DJ	����H�~Y0�:��	���'��{�JVVc�ԍ�a��j�e���e3��D���M�bco}7g���<�s|^�T`��s�]�
���	?;�U++��}�Яɫʺ�k5F����h��M��
Bn98�r�'x�ȕ{��-M��J��v�a�9�g�EZ���Pp�;��}��#��x3%G�V�ы|�zR��Q4�2eWl��+���
�G����9��o�}��0�
�vU���Zs#�@��]��4�m�g���뿿�6�ة�:�@�&las��|��=�,jD�=���1�1��gEcKG�8�!���St]vs���Zlz�y�m��i�NѮ��r�7^�|ѣ����u|l��i�%��a��Ĉ�3�Ě(�u�-2��O���t�Y</Byy����^��EaQ[�ñ+B�V�J�S��ɕH�Ʋ��jM����o��,���F�2���b�Y�v-��ď�',���<�)��pa'������ZO/��A�%az����!���K�n��>,vVH���1eA�"�-e�{���;���z��y��-)�&l�VLu���
v~Y��F�ي��E��X�v�n$Gm�d	l���u0���1�p���:��^[7sH"�IY�����9���nK�EPؼL|}��4��aɫ���
�B%v�)*��@��]ډ��6Rj�6$�X�����Ԥ���{OM�y �<�*�t�fʮ:T���:dG;�]S�(H��s�v���ҕ�vI���b5_3!{�e֤6�����5��ͯ��K;��i;X�YƗ�(�xe�q�	ic"x�S�٧�5���l?���~��u�A��.�}Ӧ��{� �g�xi+�:�'������Ϲ��Q�ָ[�5�mΟ�������d֮N��!{8
럔�ְ���:[{ q���a��<O�e���U:f+��,;���Oݥ9>F�4�������Js�M�k���рˉH���+]!ܭ�(U2#�=V���7�bB��t͇�ac$y����D�7*��d��"��u����1��C�N��*,��d��_y.Ҟz.W�o�͌��o���n��6����&���*�o�p��k�z��x���\HO�a��8�����op����zv��
��1�����@�!f��R����#H�D�&�*���?:gj��B��	�U��P$Z�{
�஗r�{fOv!q5�z���.7/�=���N���hg���G��3!O�PO�O���J�s�wa�7 \E��i��)�&���~ȫM&߂���~xh@��{1���0D���eP:��9߇�ً:o�ؚ�3�����TI]l�����Cx�5�ے"��p�/�3/]=<@ǳ;��x�`/R�ᓕ�ƭ��&o�za#�˨zs}y=��<��ȑ��}�a"D��V{�*aE�#�jb��]I������Գ�_�K��tܲA����*��GA��׸^�����d�-U�F�qB��p��}��t<�D_xѼ��b�[ܗ�X�V>�����Y�O��R��QN9�j γ�}za�1�=^�2��l��}Q��-���q,����03�Q!�m�E7�Fe���?�?%���_"��h���Q�j��w�f�;�3�?fbl��v��O�����&�T��+I	��q�NF*Fm<{��,�!��Oaoa�7��1^[���y�@|����x�:�/
��]��w^�?��t��IV��w,��ϕ��q�$
+ �qp��Kc��	�CQ�k��N�r�%�3���zϐ��x�vr �x�*Am?����6يdY�ڹ�+y�)�s�����)��2�b�[�T�������"]H:��uU ���Eo_6j�ڲ�wC��I�|�ui��*iإ-�L�N��;��c�G&���''v�5��b�g�c���h��1e����K�,��XLn�-xw���X&Z�_~x��� <��
��@�x/丸]�t�ݙ�b��@�N�h��;(��ĵ���u6�5��/r�����2��2���E�:���ܚZC����E
���.6�,\��1vd��ƿ�[�9�ȍ?<JFNs+s���zD5�pY�u�
E�(6_�@`BLE�j�#g��Q1A�^���4j��x&��
��$�$ֲ��a`7nf�D���BGw����C4�� �56���@N87M�Y��Bu����B�r�Aeƕ�>x�U����/����˂)贎�-��mG��gB3l���o�Sj���᠝�^�е�TЇ��f!�_2]̅DL�� ��K`xK�~�5l�@h1]�����rW�A�90+��a���u���ZMz��^���1�����l��ڮStކ��e1Z�����akV��|��~445u�G��4�s�N��%>�^,TW������9f�Cn�\FN�3*�����y��K����ũoYٗ.^Q��U�{ӹ�#�_:fVl�b=G�m����Dr+ք�POw�y��1�o��L1���ϝ��Y�D���,��,@#�ai��%��\��������y�;<|1g�P�X�R��Z)f���'Q��R{r��=$��������=s���(�=T�熎OuL�KI�4����|�B�F��+t�c1�ͽJ�U�<.�������q4n�|�匨v�5���<rn�N���Mo���`�ƣ��ӕ^�[�_�{B+8�YG`	��B�v�F��z}q��J�=S͆%��[���JК a�?�����x<!����@>�Rm�a�`������^�s?;C����f0�P��5S���Y?�O�i��`��i��nB;&�a�Ɖ 㗼f;{���w6�����QywHrD�˄���M+�z�Z0n5x�_�g�/R��2Ղ�� ��&s�|�7�.N���g�#]���k����ЭB�W��
L��Z��с��S�F?�8UL�xH�q�p�5Pc��'�uKM��r̮k�K�͜j�����j���/q�|��N�x$坿��g(��z|S.��\T$����9P����a�dm��c�ρ|���ľ�Utb@�Ձ��%��>�7�3]�k�7��<��X�S�
w�� Ȏq�v#�6���>��f&)t"N��k�&E���FQ4�Y�w��J��UiC��p��#�����@sppt�dt2�X��+��=H�ZP��l�Y��_7<��\�x��D��e��9�j�!`b��7?����5���S��NR�+-z7v�1:����y�$% -Wݩ(�Q�6j����h���.>y���	�;s%f�࢘|�$�S�g�_��/��
u�=���� Qp�P������ER�6{5��5u�8��\�wb1'�8P��QQp�ѻ��l%��	��kc�����z�N�K��J��Ё��Z(�4�{2'.Z4�RwAd���[��X�hՊ���땀����4������iפ�x-�	�(�p��z!�ëR�����ւ�	���Iw��o#dW��p}p �6O�J7Bgn���%�-���o����0�}₳J� �1䬙]��`�0k=�*���[.��N32�}�W�	EXl���qy� �ņ�s��cl�=fhO��I0d���:��TA[)+�1�d���2��Dռ����U�6�u�#�.j�Ӱ���$6-$&��0��(���{k�M�em{	��0���Cĺ��&EB�k����y�z0���B�8��gj�Z��X�ay�� ��J�GT���a.,L�(!�J((P�ơ���CʴV��,�^�7h#��y̦��Wf���TO��t#0��6xA���c4�P�O<���>�'��	��g���2P'M����ώ�H�&�GZR��rJ�����W�34��R%�U��ѣ=���|D�1��]=�y�\��g�D=g{˿�aJn���_��Q�KN����q��'1EPN�q=��޳J-W�J���+i��� �t�5ZO��d4u�ʴ�o�$��֮t��~��踫5b���~E�:�I��ݘS��!���n����mo��@�x�=-��-韆��3��fJmH���FH�&L-�����{dL���CK�R�[�����eadh��xC�Y݁�ύZ�&���@T+�(��Y��oA�O���a/Aq_sҷ�a:��.�������9���`ϤE9��l@j\���$��oB44���۽��1�RP�V9K�N�2p��+5}�~x�on~�e*J����Nv� ��D�*=�>�n	��&�9��(᧑�#��&I�\{�+�Ѡ{myO�<
a���:���%~&p\k�$����!���o͚��|QB7%X�6�C�A���Zw��f��	&��/b�� ��IQ�Ϙ��(v��=���(���@��԰�_��.�8���3K�(h�O|pi���8�#t,����A�P!Wi��#�)���5H�!���~8Q�Q7�����;�i��ZӠ�X���*�*[D��jo�r�M�I����R��e0"㩙^ij�j�%&O��gO.��F���3���l��AX�9//Ţ?����Qg�p�-
f-�␜Y���|�,���6��=��X���}�h�u�D})�\��*RQ�%1v+!�V\��7;%���� e=Z��z���T�n��f�!"��o�/���Z��q��}�	�O�� ��X�!|��*Sm;�b�n�bA	���c;qx���zY��������B�sJ�ĵ��6 �Wd_�����2�f�!l��tԎ�o�+�>*0�d�1R$dJ�D�Wx���j�b�7���'x6Y+sZ��m}������?�u��Dz��i���PW"R���{G$L�n��ݴ��]�����V\k����d9m>��p";��J�w�v-W~3��&�
�482��c�ѫ%a(<l0��T��=�e� yUB-xҔQ�?�������.(bSq�IK��7��J-�Զ���3�b
ƾ��	��c~� ��6k5̾!����%���^��a����KG7��R:�_jd��::X,/���O��Ґ�#@z|	�'r�����Eo��]*ʻ��f�W98��j�z�ZZޚ?����΁�(��܆]
�z.��z'����6y.�m\K��H���.�H�Na\Ɋf䦦�x(��[<��/M�@���͙݉�\g�O��B�����N w��1�VE�)c5�j��2�7���چBխ߾�Ο�7�s��<<�B�$V=��`����^�&�h�\�@�Qb@� �ܡVKˣ�țmq7B(���'�H�/�gi�*�S�ɷL`��v3�'-e-uԞA�n�Ơ�z]1�e�'C����<�����Vh/�&��G{���Ά�3�2�~)����f���	�\���gNq�:��3C]����h};��J�\��m��R�*�N��\9@'�:�\e ��E��:LTN���	���d�(rd��5hCv�#��������汤���tFx ��S��4����J�b,$aH��q.w��TU��Q�Y׬Fw���v8����EA����%U�m<e��z���յD��Zv��,������o>����-�*%k�i�t.�N[D7�!OP�y1D%�z��+���I�E1~��
i S^�SO�^����)�2b-ץSy��g0�PV��s�s	莩���e��S)�R<0� ����΄3	�3@O�\��H.�1=8_2���L��f�Z��8uTL�rع6�?3*S������[����V�R= X�\+����.F6��ga1��<%{�e�����az�(��p���Z�^c�!�\jm�J�:p1ߪ_�Z�zжG�hyM��:H1%��-�4�`��H��ڂ���d��	n�	X
�SY[w��MzD�4���U��o��e4��V'd|�I����+D#�^���f�\��3$�3O����3�Il)�Q�i�����!tu�1IX�UPh ��_�5���+��׋bJ��1D�%{��abrJ�5PQ_�7������)nv���d�C��k%&�$źsⱱ����\�p��j9�o)��Aoo�n��5����9��L�i�sC=��э�x������8"h�b�k%Ph;��l����5��������2�E2V�w�Q�3`�s�3�:��'��D^s��Ŝ�7�(�`�v��Px�jGӹ��>6}�/)XA�Op�d�O1���0�Ib��O��s��N峢�oE�Dt��"�JsZ���Sc2�7�o�6�/b�%�Q__���ĖJ�Џ`��c�L�����D?��M�w �@���$��NDQ,�$lN�h\E���|�C�Yipi=��&	0D�a�5�P]���E���RM����i��sT���_G<�ۭr�T��
����D���ݺ\�s�~9�J�ԬO��U�U�6v�HFyG��Y2��W"CC:s&���\<SOZ|!�V+E)�7Jh�X^l_��SΫ����QV�1V��q;?��*�&�^3�drH�P�?�^��:��_8O������D���1j���^v�D�'PqΟ����ڗӪ; ݬN�	L~Y;	�0��Of^�Dz�3'�@��9�K!�:�U�O�vŹ�&����9�'����SY�T}�<��i%�k1C��Ҥ��pQ(�%~���Ж�=�I�����J��t��4���}��ё�~��_�}��씠<C.2#Co�7&sf(�3g2��D�@�ӧ��u*�*��Q���UVc`X��3p8ͯ�4�}g��VJ8������,�;k�"$�b݊�����a�]C�+[���b��e=����~��|*���D��yqs�sX��n� �+�1�0�>>=R��%ʰ?�;�l���B��m}i���o]>��	���v�d��;
{�A�v��,��ƭ놷y�T�������~sڔϣ���K^>@q������9�,\�#�� vi�5<O��<�%����C�C��QbXn*1{�QuN$f]R0�)K�1y �� O.��6^(��s���Ջ(���l���ؾ�e�Id�@�H�����fl��b���{����f����K���ey�G�CP�A��)���ѥ�A�m�'>����-�ߔ^C[��Z���jJ��!�z��i��x�f4F²��{�fd&���`[:#�KA��q$��#�~j��=y�o}e�L��yo��c����	[8�H����D���x�S�AzQ�m�&�6S��!䈽��B��+��x�����ս��<�-'���鎕Sg'���<7�o�9��Ӌ�!�Y�2�������p�U�0���W>���
�G���Cq�ҁ�璦��
�0G�����o={��qR��?�,�ɲ����4��4~����p��F��1���s��t� ��N��d*n�2:���bOv�ޔc��Q?����Z�"$�>�2{���EI:�ϭJ`����_�K߫��N�،��]%�7��̃�� K7��Naږ�Gf�Z �2����ȕK]p�y�{������/�����mڤcQK����ۨt �m��¹�^ep��`/p�w�-���j7D�n�٥��ݯѨ���qœZ����q�V}��3N�Y�(����k�k�h��v[�s��7g�ƾ�7Qd�׋.� AKfL��<$���9�
R�*�Q��J�PΫ*�=ㆫ�<���UC�x�ŉ�6	�>����2mˇabuf���љ:n���=��οѭ��(Y2�4�� ,m�[0h
��9�&��DO�Rf�x��R+����d����.�g0�Q��p�دg��Mˠ�D]��r*Uc�;ҍW˅����^5�> �5y5���&��i�j�ڸ�Ņ}�^6�b�|��b��E��Na{��ŵ�,�sɿ��]��耺1�������sd��iq�!���k�����#�1�+T8��?	��2D=-p�R��M��`�9;�������x�wL'e3r� L1�憓��m�FK㥃�rGڂ\kY-�~�V��y4�E�7�����s-h*�^O�U�Ň�j6w'��Ih� P�Ȩv��"[�����v�2������98NR�J�fpT�S�����Ñ�������{�G��b�N,���38Y�v
�����	��y�o� e]�jl�+�JN	:���ҏk�%����N�}G�����,�"<�|���k���ګ���,&��<� �Sˆ��@q	��r��T/0.�6�n:lf0��'8lq|����,����e���-ÖNM���5�#*�+RS_y�~Kʂ�ڤ�m��a���,��EX����$�f.�I�D9�A0f�/�C��1L�i�L�5�9`W �R�E�øȤ�"t3�/����(E�/r�X�Y�� V����R���DR�P��<�neq�hEP�n!��.�;�^���]��,i;r>߄[ ����#�q'��z�Tb��]�2e�질��	o:�\wj�襜���+�Fd�|d{Mq�G�Fc*�K����������r�sF�����0ON(yoR#�Rg][����-���s� zW�Y�"�wqmK����p7�=����A���̖��2���zʖہ_;ѹѵܶvdD��i�7���M�����sE�s��"f�G(R�2��
�|�q��4���(OH�_��3�y���H�2! q]���C�!Q�`u�A��S�_rn[ y��H6S���2j�P��x���X�q��aC�B���,0s�[����T������}Ģf�A� ��6^=��m6�+!~[���O��Dh\~ȑ��V�J$uN"��X4!�XUBМ�X�� �UpC�]lN=�����:\�/�$+�Q���)b!d�X M`x�^�/:P��Ӟ2�|�ek�a�:�TG4S}�=	vظn�t(�ka�RԹ5ՙU��Ē;��S�+F��T�s!b+94�J̑�������\\���ڲ���K�02���^o�x�]l��թ��"ۺN�a���k;����a�L��2F*��5�Z$�����+�w�4�g���Eŉ�>���ǝ���֐"\��i�U�K�}�ƣr)�;�CD�������DP�=M�� >
vڿ�����p��G ȯ�,7�Q�KS7�;9XK�H�÷��r�� ��%l�P�����e�b��X��)���'���Y��3}�W��p�3[��E��g��ҧ�p@��hD�퓰�38��|�%�r���G��T�r�1u��,��d�]�&%V2�@a��\�����ye�8r �>�\���ᓻ�1s-�8��^Q�֔;H�,rm�-�G`��Dܑ�i�r�-���#��`O��.�yU� �z3&^�TG��ݼ�z͍��A�3g�o��hG��u���9�A�!�!�:��h�U~��b�}P_�S��R����`��5	����	��M`nO�y~%���B����/����g�Ќ�v
�H����k4F�f 9�P��� � Yv�U��U��l��1����J<��]X':�7#J�0G��	��o����VW��Vvܬ1@��04V�վT:dg�:t�;�s�K�tC�1��4aȀ�vX�3�χD�pG����ͮw-��&���ٻ"�ٴ4qAZdt�����B�0#�7t+-��?Tb�����GH�e���0}i��k�&L�����D�
{Jëu���#��e���h"��}'A���u�yܖf�ug{�yI��ʈ�M��Q�C��I��`�V��8hKq��_�l
d.{���=���Y~�E�e�}�1���}8^���C=P�g��o�vX�lȵl�;�G�-� �%�!�LV3EIdO"���,І�|�$�������b�e�?�ߓ�$|!�9�Rl#�ѐ�^���V#���:z��]tV1��,bX��Y��A4-�Ugl�5��>f���FG��[��<-sΌK�V.�p�.DH�6����*�#|�Z�F��I��j�|l�Ӎ�aߴގ�F2�_7�,������'��������k���x<�־�J��ފva�n?��~��A{%�W��v����1�
�A1���9�5-(�o��#n�I,�-J�X'�čR�:���/BA�6�Ix5��u��ж��7�3�m��
��)^X4�,�-�Bi��~�f;�4��<�:��/�����n�!���	���[����6�{�Qklڊ�ѓwp�0ѳE�j5va����(8&� `�@󇛆��&Y����N/�	��s�yhY ��gx��]9bɽ���0�?o��e6J��;���`SY���T��H)�:v�aɌX��ӗ��F�>.!�U�K2.��- k"�(URC�e����jyf���OwֵiP��T�?q8uAg�>���CI��݀��k3ŗc��8N�N�U��zzґ���h�; �t/��3H���4�{�W��_+���;Cg��>);�/㦚C���vw��e�6�D�(*���Id;ʴ���hc��PckSK���7|��������g��*-e������v$}�u_�Jda���>�ܐ�n��E�HHk�b���VB�<�\8�;9cJ�˙��7���5�f/�v;�n*�yt��42a[�*4���F���D.�L�P�C-���@sъ����I{7����3�A�_����dh�z٩*����Е�%���=��v�1ic�@���]8c���K��� ��l����E��؞(y�|�jm�^����X�G�`����M�N�@'y�U���}7�]�%N�'d��|]]�Н�̦�͝C����5�Y�9%i,v�/����Ս+������G	�ڜ�_,\Xb��M�A�a�sݒ�R�6k�&�r>�2$[�ᶽɏ굲��QL����-y�Q�p�G�z?m��K��B�!6���������l��_�γ��5	w~��#��Z�����@�>d\�U�]Z޵�����B������f��e����d�N�A�j�#ԟ�(�I��	׎lY�D�(k�3k46Т�/¹W6����P���oFa�l�@ʮp���¨T�?���o�W'G敳Cˤ�"/����M��^��w�CuJ;�#|de۷Nx�������&�0(�i#d��ek��L��d!�z�N�f�Y������>v."B��r������w�N{.��}{$�3�l�-�J|������0 x�Q7G툟��T�W�#%�6!�p�?��6#�τ�[D+�ݬL�	�>&}�9�c�����cG*w��׾�D��}���d-F�7%��.v���]<`t�[��%�s���y-Ǎ��@a��#��~��L E8�y���|U�-��A\� ����z|����OJ݁X 5����W���t���5ǈB�b�[y�c_x�OQɦ iPި}�Rc��i# H�UO�C���h��YƋ��X`�7�k�bD7j�C���cZK�BYA��H�)�
F]�&����T8xۧ�|�X��N�Phv���C�4s����oƁ_8�V�00� g�DÝ�՛��F���B�0��ܿV���7�:1�*��>�J��*t��/^j��������T��&8�>/��}/Yd
��usVN2���g��<
�ܥU�
$�@��_�<w���y�E�`?��j˲�rJπ��؛�@���\����͇7�/+�mՉ�Y
֬��FE �l9����\�;�����s�x�3�Q`��5L�榴�J	�cty��
	~w�L���f�h�p�y#��b�uH�p�e��Z�� A�̥k�G��&脴������
�;R6]�����z�*EL��c���K�! �HƂx+h�1]X	7ۍr�/��S��ץa 0�mh
wD`2&3��4拕eD͚��8�����-�ct ,����K$����a����/�P�e"���B��IR�\> k�INIm�̷�M�9ze&ma�,/���c�/����λM�
s�Խ������U,��``6�&�����^?��1���`=�����y����M�{H6=>�Ia��U��2z��Ag���@���;�KB��G��Ɵ�{��������ɌP���W�嫪S�vU��3��6B����/,q��>�X4���Y���z.`����ŏ������JF����{�ަ=�:��Vf��u��8�i��-!�XHx"��qe#�\�V(����M����+����}V����S*t����ί�2��+��G9ʌ#��~Ahꢕ���fG����q�)�jP�u ����b�u�&�/�0���H��3�ɸ����L.0'�q�����Ce�Y܏-��gH�j=�qB�L�#ǜQ:������u�*�h��^���$��� ��f�	��LF_�����[��w�%=��VZ�w���GG+.w�]�`$A0'N�Y֤?��]��P�Yۄ>��+hO��ܢϝ�4�D7#M����/"����'���jD����-q���78�͡�2�r���u�-
���}"�;�d�ϫa~b��uA�.�G9��x�x�]�O�hy	��T�`�K��Ū�y��qk��+�^��F�a!;��@c�n��*I=,��p�TGY`2]��Be癖�`�m�,�J7E�?��Ӛt���Y�#���OɯU�-I��L�ݘ�B揓:~QD�ӣu�5{�ԉ'�Ή%�ub��_�������
�}����iXg!�3�۔�4��B׹Q G�D��߾�V"-���8秙�&cr��!�"q\���|�8<�N�U�K��ϖ�L;�Q��%4�ݰ��}��>���J��*��֯ܨ��@�������V�/��N�w�����Px�B*��hA�C2�Ǥ/���`��Q\�`�vm�ݢ�-ْA�ax�SZ���+Y����D&���J�Qf+̞N��Tvwq?m��C�8�5�P�ﻃ��~c|�W�	V�0ti��6��#t_ȖƐ� )��̰��o�`��9�*���ˉζE }�: �rC��B�#u���� Y[�?�(ay�c������^��*���4&F+-M
��nw�V1S��� ʨE�8�_,��/�X*HC]0/�(�\*�h�=O�gx`�n��5.k$<}M�Mm�<�jE5*B!ɻb�S��'A���\�*���@ۡ� �Q�`�q�}$@K-�*v`����<��iX�b����NMY���S{׌$�{h���ʡ�"\�=�q����,�]^lE��u	��A�e ��<[,��,�sWq@Cn���K�޶�[k�C��㎝I����;3��zۜz��� K����]��xYba�
��zq{�����tO�p��P�.�1��9���L��ip�4D������JS)��V�^�#���$�اN��5՛��jȍ���c^����'�)[�<Fa�L$�K���M�RӲ���!4rcż�؍���c�<5e�川�0>�����m.jT(�Y�WD��q��u�/j{&���߆��Q��0���dW9,_���`���U�4[>�y��l��wKk[���f�4��h�y�-�����
׳�V��t���&���.�S�w�tr��}=c6�Dd��PĦ��r
����x]����3L����Ƿ�ظ�_`�T��
uj#dpFIAt�Y�g�r�����ܮ�@\.����J:�oOV�@����t`�?y��]��hn�Yo�̯���%ֳ�H�����J>Yw~}?R��8�*(.�!���xx]*���q��3��c���Z!:sp�:���!B#�1�<ob� >�H7�x���@��T�h��b�	�}�E��]B�`LVx��2~��ڶn���/�!�t��%d���3il���Q���;�]<]�q����]����ì��]Cdщ"�H�,:�űYnR;�/��ڰ�� Zz�ߟr�f��I�ɦ��#��aY�/�j��f���1œ.�� asTo��kʵ�nz� o�	y���t�!��6�o��'��֑�ϫ��Z`@^���E�>�������'��>Lw�H���P[���E�� ���Gjf�eu���i>F�6�gW*��p?��L�!�r^l$�P���>��;���U��{�1M���q��G�B� $_p磁A��]Ο������2�dv%��I�Hg���
&I��7�4��e��%t�cd�c_bNg1��������zRL��r)�a���O���R�_C|װ�{�~ߴ{l�}�����.�'G�}�I|���`IK��+��[�)�	a�[�cMV?j�V�_���o�,t�$�#[��!�R�=c��L9,FA��]_���6-�%+�L�l<��X4?�At��FU�ÍV�A3iם��j����b���7�zJ7�Q'�~� 4z��o�ۈ|����rb�,6�N�U�A�]���#�n���fR\&4�/KK^��I�(�a`3�s�.�]�2�\�=,�z�e������M�P@!Q!H��ҭ��w�5y�\�l�a<5N�U�;���}?��Za�l�ݗ@� )���<���)ؕ��I%�Ӑ�a�/O�R��� r[q;N�Y�~Fˡ���P��0O�o�#�;�A����	,+��</�T��d��TVA��OM��jMn��2�ם�\!���e�1�"�����C����xˉ��0��M�Ы�$�c{Pĺ��D�D�G�V�b&�X�2�bR'��1��G�?�k�N.We.g�\o�ۊ늮�D��S�I���ۦD�bQ?�d��O��������S}�B�6\+¾׻�j�2>������4�>���������=5f$�\��2�bVI�WKo�� ��M���s�g	�ur�W��4��(��?�[
���:y߻'�L1��$��b�Ǌm�n �<�#�iǰ�4c�Kd��<6G����pz�]Ǻ��<`^eݥGA�}���0�Ц���V%$%��[�9E���}Z���gi9��ܷ�~N~��>�z�S��E���$���=����с��k�w��.!��ב��OZ���嬿v�H�S{�G>ڀ��Yf����o�B��ƬS��L�&�~����:�d4w�;��Y���Xw��Ey�|Q���``��8�א�l�ǋQi�W�-o���ש�s����;H���h�W2y��~e����o:[0<��#�� "�J�����a�9а4�����6�N�a��&�M�����q��xTκ@��ߘ�1䁑�>-ԖO����'�f��E�����|dPEd	r��,��Y��g	���bD!�E��ѫ�1���Z�S}g}C ev�~P\\����ɐ�ɶ*D^�2��MJv��ʼN�f�م�=X8���N������z
���گǾ��:��e�xQ��`��ӓ61��3���Jvu�:Z��,�~�:(Hе	�l'�9��.ք��)(�i�b2����c� ����BP�`��|<��r��q6��<���}7���ԗf���#����u����i8�r��-��P�R�M@�%��0��;ŽU%���25*&#}ġ-�_��֛=��v����AS#��W߻r:Юv'�7�o�>���Z�8��y֌$�X���/�N4�&��s-�q�_�8:αo��8�����v���NP|��4�o���]t�m�C|�8��U�8���:̤��e n��B{v��/y�cP;��hZ�>O�:pɨt0hd�2Nj�����_k�y2dx[u��p���x�񵓬�c�t���F��xq',N�R8M]3�5�;u�|A�*~:f�X��f���w���H�}/�ޭ"�I��9��Vh��j#�Wc�0�y&�,�kvf?�rő��$��E�������	��u���Ṽ�&Gmje��abD>5�n��:y�臡�h
�R�<��\N��gH����_p�\VgOM$Y�ԁ*a��L��YXV.i��\���4�>��M��e8v1��S�����8�G�ǽ���F���/�Pb3�c��'�м�F�T&b��`���G�������|�iq7��9��A9�f�I�ԲD��^P����m�t��ʕs ��8���r�_3�F��2o�{l��� ���������d���P,���Ȣ�N�vH}#�1�"M���*���W�!(3��Ђ5 Tm�@^�� 2#a<k��T�� �n�Ss��a����o�M��6�?�Jc?lK��f�dC4v"�����S@��^���L9)i�U��\�{��0RO>rMt`��:��ʚ�(��ܗa���m����7ᦩԞZ/6��U���Pr@�{v��/�P&�-Un�]�Y��{}'W��QLUv?'Ӏ��G�Ͼ�����eI�RLFjD~*�qZ9�X�q71ֹ}�v�%=m���,�0��-�~��`!�:���\��j��L���L��W3��撇v��71���w8�߃�^gg�ϔ�4ۚ�"����ܕ��Vv��o�FOd�Ò����BX��A�EKp��]��^'G�T��-�:�B,V_��#;{妬�8�|&�=u�I����*�f�H�&�o��'�D/%[sϕ1U�9B�k�5ʱ,ݿپ��ּz���t����F��.����➐-��&��WUN�Z��Q�m��p�7Q�Sw��Q�}s��[r�_�K(}I4�4�����hI݋�΅Be�z�C�c��ums�h;��8J�C��"��غ.�O��R��G�S���m׼|�Yd(�5���)l4�b'~��6n�f�2+
m�T�֡�&@4�Byڀ�'�n�8x@� �M\�>�P�WjL�����y��?�&�#��b>%�`lF���#	���1[�@>3�%���=�������'���b7��G�ePE�$�ˉ}�F���v�5.1R�O��xgLF��s��<�_����ZXP��(�9�no`\Vz&h���j������"�3�Y�[Y�* �/��t����(]�c���ci�l���o��21LԪs-�I�!I�w��O!� ��%����fd��ri�4U� \���Q�`�_"�y��m�f�抅g���A�5u�k5j�֒� b��E�_�Q,8���w��2���%s�a�Br�-��`�<z��"͗��I7mr^WW@�Kr�Wjg�x�[�Nn�TE�^�^�k�V��=��������?���F��O*��r��V��0�#�����Xߔ˓m.n �O�;(b{~�ژ����<v�!�����@N+���s㣎|K���QL��|(�h�P���Gr��m��2��]@��_�M2��&�� k�Ga��U>����^�oM'�C�[KGI�@/�t[���8�q�$��E����F�M�;P����g��p��R�c��mp�XҖ4�0A�*�őތh,�r�@&2�b�,}���(0e	p{(L^!p:�d���y�����O�n)<̢��+k�,�-���g{@��2
F�����4�z���Hv!#�l�>?9r��އLO�+���x0�p���CtOdDz`�+��c�x���1^��[�	&�Ϸ�c~f��\@��7'#�fq_�ك`��B�,����6�p��9z�ǖ�!){dO���aD�)Ϳ�zݔ=Q>��%�]ۮ��(����q�L�`�6p/З���@��-R�4f��|�"��uW	�!m�W>x@qǛ��ʣȝ+� c�tF���V�,W��i�[Oy&&ä۞RΚ�q11�yP�Zc���T�W�:��$i,P=��f���{+g�֣ΙV��c�ۼn*�q�|L��R=� �.�6Tl}����64.�O�]�v�N�5n�6����l,��t(�ٝ%3��ʷ��lY��gD�=8ٸ�y�Fvٱ��~,c�F�q���1f�ЊC���E��I�L��l�Pe5���ǟ[��������8���pi�o�����-Ua�h�v[�i�c�M��j�t},��,��'��uq�%R��C����vc\C�|�g�Xu���*�,V�ڨ~e�=��S}��J���6>�AQn-8���n�f�g�m��>U�Ǹ�8�?���T�(#%x�1(�_���'���s�w8�@���D��9�PZM��-���/�DZ
,V��&�Mp�S3�����?���T7#GP�X�MLި������`���15tg�ݯR��G��gy,������`�b�k*'j∽�uS�^������ֿ��Xr%�,zdc��c�3���tߘ}�	�瓞j��Y���
�����}ϧZ"�֮oW4�V1�UTU��u?a!Jx��l(�-�LD~r7B���0��'�C����>V�6�\�m�6��apO��v<&�Yd�[I�{�k�D�;S����t�D�ǵ)��Ϋ��b���g�T&����A�c��j��c��e�5�Y9��j�A����'ѝ�h�2:@�is���d[>Rc�O���m�����Xlf�����̖����W�o�>�i����G2�/���a;�M��I��Ù�S��e�
�*���
xGA��G#X�	�2��ɳ�][��Bnjwq;��Q�1���=���*��{S"<g�q ��oO��{�tY��6���E���d}�P�oL��ǐ�Ȼ�4G�X��޴�� ~4����>j�!s`A�9 EF�E��ky�K�Ѵ�����ɅF9�yDHnP]�%I
T�����ǲX1����F6�����TTqvy*��H��f�LB^{�̪%tV�5v��D�����|��3?Eװ��ՇG�ohpB��?u��ު��`P�_W۰,�fI֋YE�f8~�������%�d3�����ᗷ(�0�����RT�nR O��D�"�M�$��P�a�:�[��"�4�P(hs�������a���K)�pL�"��\]K��J�ȍ���w����E@�W.-ʄ����YYxH!V��_5p�^m�!vB�����+����1j�
QP^�L��%��K��F��q��|��Ԡ���
l��]��c�����5���b�n�RT��Jd�CS�mXoeݧ����AWF�KSM/S�#Vg2AL���g(����9���{}|U�?&������$�G� ���3M�����{œ��k6��B@9��N��e�X��X�)}G[-�]�h�w�"��Q�=N�]�{u�49\:v�iC�Ɵ�_%��m|}�UC�e~��I�����Wt��s?�݀e���F�k����t��+)�feu�#к%w�@~cN��"T(뺌���N:�3$��i����+w&��ۼJ,����`���od`���c�T��8����&= H]}bV>Xq�� ����^�3�I��:@%-5�M��"��Y\e�.�v��a�	�M��c���T�PL��C3ɶ����~���-���^�,�ݒ��8�(����z�9��l�����6�?���'��\��D���w���+�����C��*U¬*�����&w'����#�]�j��m_�(�FI���?��%'b����l�;�E�(fյ昚Ԩ�:�{�e�HØ@��.����G��~h+���G<�|�����AF���%���(�o�@�и�'��D��}����y!T𶁨R��M�S_o�X��o�$��{���6��5syvi�9��IPS��l��y�5�j�؀|������n���%����XB�0pyS�f�B�.=��x�4"	�	�`����@��V�-�~q��php�Y���^(��1.���a��0��:�b9F�2w�!�ދM�Q�1�CO�W��
Ypsy�%mb�ojw�!�3�GW�ۿ:���ьf�en�x����1��9o7��x}��,�?��[�	�d>�O�FA��(��4q��$�f����Ț�v���et.m�x���W=�v�?�.g���(����=���3�CFM�sά.I��־'�w�`���e������s�}�JD��}�����Ȧ�mK`���v����ڠT=�}�h?]�����+�x.�V�ou�'���n'���������-������X�@�o`Z�ؠ	y��$U�^a��`8����� �r�?�V%5�/3�#c��ͤ`��5����	D"�7��U,tf6I�S�Hp�� �@,��6ܥ�O3���lX��Wo��)��5<PYB��B@�V�f�!����WB�lF
�����	ݑ>��}����9�6}M����e��}YH�|BN��z���u�-�f;g'	� mS�v�>^s����1���N@��Wh��`$���h�ާ��a-P�'�M4�;Z/�+ۿ�i7�dy�[8$#�������[#1�@�$Gt*L���-�q��}A�x���ެU�48T}h���m��MB�VҶI��W���$���s�C.F�L�8��1�?I6�5�RD<h;��=��Sխ�>RoO�9-���鑯�L��Ȣ�핚F�ƢQg��Gâ-DUde��x��󗱐Aʠ+ۂѩ�':��z�xD�$aD:l��/�2���(�%d�IP�'�r�`)��)�X�O�SEf����]@���g?��W��1�}�Ƕ�Z��4_�� ?.\0��"�����7ZO3 bG��^�L!�W{y;R�H�t�jEt(�OHC��w�[LC�W���>%o7�R�X��oT���q��2´�����S��c�Z�5��u�a�SS��"���ϓ=�>��b� ��n"�.'���d��5�1��$+_�>�n��k��\�����TͭɶV��I�`�q:���2���:T�x�eC�������j���v���=[����h帔uy�����܉�'Rj	��=�8�ٷ�P�/�^�#�K$�_��������V?����ۯ)�ē(8u����CfF��q.�������f�ֻ�P��%#S4��e�Yl�I��#E�����%�M�X��m
��1���us>GF0SO4�����X�=��ED��l�T�M�Q��yR�G�E�Ag��N��-z-U<ȓ�u�D��
쌃�s�*_s��!�� �m�x�f_�ܞ�j�i5L�f������!����+��IC��6L]��O��1 �UN�wG�O)QxÎ�4���ْ�Xœ	bys�ז��Q. P�bM}S�}ɦ��15�t�b�/~��M7O`9N���S�v`�j�&��__�����tf����yܰ�^@�&���^J�~�x��2�֥�����/]�?��Ioįg����[n���n�r�CnCA�N�tȹz/
�:��<*� �3_J�0�Vo�CDm_�l��?Y�$O(��0��r
��KLt��
�6����V�q_��p٬�v��:F2_*�eΧ��U�f�T�%Xsy�z����N/8Τ�fP���O7���̱�=����WT'o2���}��Ş!�	0o�+|�)��Wz��/\���U����IA0�J�B�>^���E�y�?V��X��\b(���m�$c�0�q�z�۠��K��`f���٤�lTlTl	C[����K��}�4j�]�Jza%���H'?v_"ުnZ�>����_Rr�C�u�P	 {#s���� W˳j���G!ϊu��cU�z��C�����ҙ�(r�^«ʂK���O�hb�yc(Q/d�G_Y��tb){eF�r�l���//d�3>��qK8��o0ӱ���Q�l'(�/EK��X.�sȑ�0��;v�r��qp�:x����ʊ���z�G4�Gk8ew�"ɏGĵ�]"Y�{�R!��c����q��4�Ht�`�^'{	nw�**gQԆ�F��%@F;��ӺP#'��#9���M�]��)^��9�N霻�-�����/��Hv|���V���F��
���\��G<���1��">Ȣ�٥��w����+�ٻ�p�@�I�L.�LP� @�D�Ԣ����^磫\H4Z_�c������ڶ����-$�adY1��iYrD�v�θ6��_A�(��wW;͛?t��Y�D|�'C�}��J&�d�|\$�:(�֊(^�o��Wnpq��zQ7/��'�!��b�L)m����jy/B����P�+�x�Y��$�8�ʅ���ޤ7x��nx����d�NP��'���jH�٨�1"�ݸ�k+����g��V��=�\Qc�i�nl>s���z��J����3k/�uh��%A���By��8���y��C$7��'���E�~p}mH��k=y
	��������#�������43�����Q�$������GB�FS[7��|$S�I��o�%<�S�ӱ8�RN�\�*��*�Ԁf~'	F��]V�͔O�9�:x��h{JE_��g`����)x���o��p��ng��\(ec� &�����7�\	zK�f� �9� �P*�)/I�g@f�ᮐ6J��/R�����;����[�m#e@[b����E����q�	�VR(n��Cqd���/qu�_�m���y�<(5F����,����Od�֜�|e�h��转��ר�b;��U��NT����&J�F8�Q��)�zA�����v���0d%�x�+k�0y�;�u�1h�Q������#�ZjMn��5蔷�}� YhO�}�ļ�G����^#G���-��J�ā~^����j��@e��\ң� �|ŕ/o���;���ȹl�:�M��Odn^#�cP����J"����ߺ7��
��_`Un��E����h����=�C����µ����~��6���V�(�@њ[c_��N�+���ha@��>�t�]RK튤&�Y1&}�Io��=�9��"����4�X�1�W��[�#�������-$;�����s��?юΧÅ�n���I	��|j���_-���\�\Dqjx��E�+��l[�` Uw�r:��i|}шȂr�k#E ��*��԰u�Z�9z�jf�sG?�M��.��M�ٚ(F�fg���\~��3O����7��4u,+G�K~�{bWփ�o��i={=��=�c�E5��a`�'��#���j�Zo4�*�7%�����-�f���I��˴zE̋�w�I��������rP��!7��ZE�U�&$M��=�dVMG�iO;ѥ��R�t�IA�ؠ��+6�3蟧��{$]P�����(�nCz�FY�A��y�ѯ�,�7��ҔDM��_�/R,��³_������2�N�_!����,,�-��w�q���H�Ư�_l�Q��yl��E�9�&';9M��4W0��+�^�㭢	S�&��A���>�AgG����n�=�ŴP24 �[{��_��W�B�n�m�,�jNK�!'�ž�����f�����6>m�_�Q������0?l����Q�H(HTf�[�N�7�R]2Cu�`���Q�����W����s���������*j�� |���'���f�RA~��|Fj.�/���Ղ b�H��Mښ��j��!�0G����Id������l�����������ӫ��&�ro�J��]�ޢ-�����ju�b@��W�8�>�U�ã��7��M���{s%�����Ճ7�����?��,�;W�9�z� <'��&���S�	��J�A���1�8�S��~zgnT�+�f1X��0�(*���������|���/:|���Nc�snE-�\������^�E�t��*���u��:���h��}/��b�|U��=G��r����`�`d
u��*������q��9ѹ*X8�v�ݟ& k��vC>g� ��j�)Ҷ$���ة����E���%_��%�x��v�������o������j�l����uh��8�'U'�FLb_8�2��?X_PUĪ#���b�k�a���N��ny6�;�h槥?�6/�t>Bf ��!��m��(Yz��b���`Ě�����Wu^;��K"jf�g�<+���`�]�"�/�m�&b����(5��uH�ꉎV}8��7#>�Qy��%m��Q>� &�xq�J��)��� If�ܑE�$������e.M���W���|�,�0W�wo���^8�⊨2��Lw~�����_�Y��żs�}�z�&&�a�k'�H=	�m�o��3g
�4��5��b=�ع5UN���w�|+���gq�.�$Q��e�!D®)������pR��R ��d��e�b��gN�>�����Qهg'�M"�Q!�92Z��*r\;��?�\��#�,s�i:ְ�)�Y�>�����lw���8���ׁ$^~:VP�����Ɔ�2;���lbݍ��ʏ[��3[�`��ix=�����5�f�Le�A%Ћ�滧����Rc��F+��e	�,M����������u��?�R�'K�b��}��7F�G;�$�V5�}d_B��=X�l���=������܄$�'A�a����"�ZE�1[V+bJ�,Vvb���@��A��n)UJ���C�gW����հ�SdMEF�%&m��t����y4������	[�$�3��B�n��o�(S�9�Ǉ{��Tv�r`y�A��l}O)N�tL=d�r�z����btO���$^�e��گ��f㐪��l�^$�:�l�>�1���Ȩ�ϜXA�$�N��|1�yXA�䮌>�CFŞr�D�ٹD�T�TY��@)rI���)>��#1(E�@�bD.
W_����2��T�A����H]���q���������'���.��[g
,:=5QAbq�8�b��7��Jh�;^F�t�$S�Fh��5