��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	:��Ii?���s��w��3�V؆�͙���d�;��{��A�,\pi��⼅Zř�Sh�8�'��9C_mRXy$�������a/��2Hd���7�AxfQ�����[#�I����5#S�N�h�_\�A�Ԅ�!G_����MV�;����N�"��J�'g:s�����]�j��%�j�Qu�������s���SM��g1�Y���}h�w┾� ���H?zIH4�XjXWK�*ѻ�������;����7,yT�z��8�I��q*�ڨ*��-
zh��ј��N�Z���.����CC��,i�lL��i]�Ĺ�!)b �!5�W-Zv��
x,DPg�	����:{p
|���X�ޕ�Ƃ_|.�K�H �t�J~Ӵ/�-�Ex����}s��(i:�e5�m�gߏ�@o��+� �$��Ln~��B�>ҳXO���A�����ܳ�7l��	�����#>E�X���#�.X�E��"�#���E� ��L���ˎ�o�<�Rj��\4)�:qO!��bS����.P��Ի����o\��6���)@���u�+�>/uz�H��w�1�u�R�8�<�P|p��kQ����<t�+>��"�'��'0 �o4��5�ظDzL*NМ=*��ܱ@��1jtz��j��,�!��鬤����x��1�:��S��r�aړ��ıJ��3<�7���U�!>�
��;wIǩ�B\��7!_jn��K��80[$J�.�%-��8ڰ�Q�JW9��T�V���r��8�K����t��j
������_-�{��R;��K&�{��7�L��p��r�	�y<�]#3����1W�8)M�����i�jdJ[��(Z�f٬��e�zp}��3u����Xg@���6&��z�L�bWFbޗ_��n6me��Kk)���n+S�����v�Ƞ�z�٭�.��{cR#Е�Fn�/��0�����uy���Pͯg��l�z]�X�3��}��L'�*ϵW ?�֨I[>�"nҠ�,[�Z��	�){|l�bo,`�,�ي���s��Q%��'�8	6wh^2�� A�8:Ag���uَ�,ġ�}���O�y]��>ky�i�d��OY���Y�y������l�����8&���7��=�@d3U�i��gL:䩵�G<I��<|����n\r������E�˾�~�8k���d���._rm���ۿ�nC7�&n�zg��H{0���h�T�~�b?M����YRȃ	��E�Rz�^����8��`J�8�x�cG$�xL��$U��3�:�>�M������LX����yR� ��CS2m�!e�JW7����� ElL����f����E�v��M�qۙ-��:���W���#Y���/�͂gv��U�j[h�i�����u�d�!�����K����Yy'�@=����RM�f�{����FE^L+����%ٌQn���8�����R�6�lΏc�Ac�z��T��0���"-����k��Q~��>��S�8���# o&!{v�������$<�Ql����6�a�`i��UߩHt;�:�!Zoz O����H*:���yߏ �?.��$��W_�.��p�[r��ů3��S�#r��痟ߣ9�F�f�,�=�󩾝���Z��#$��N+[� Y���;���*����H,2YGd��\�������W�H}}��Jh=�2��V���M5�O�,��y<�=R��o��(U�F;kK���:�O������=gڹ�'5Q�tV�I��}/�]>	�<�K]�������=M�#�u�Ϝ��T���	(ʯ��iLEt�=���Y�=�j�g���C�q�|�ېY�(����*���M4�i�7��o
��#�l��,������	�=��l��\\K4h��1;��@��:�C�>��<��!�	�M��0k���;Ibk��є|��E�n�g�(mqv!(���Pv�3��?*��5�E%��#P(��i?�Y:��p��=�M��a,F;E�
��k��S��q�R/Ę��1ёNڿ�;U��ؿ�1���G�7�n���L�ީ-{�� ��]�\r��*R�2#�zo�u�-�p���R-Zg�_d�z�]R��1n��t8�r(��W���/]�n>2���G�|J���Z6}�9�:��
�R�.�J	M�v7{8V�(˷����Zv�s�F���dԏ\���yt�Z�`>��
�W�[x�$���T������D�e�yfQm.�J��	�ρyr�~_'�����f�b���n��62Ј�����H�k��}>rOP&@8!� ��}Gz�n�O���<���Y]��:z�[�h*�n��w�o���X�eܭ
X��B�˯�|0�J4_�擸#Me�Ef�p��i_��H�\x�33�s�H�6w`���0�,V�>;�~���/�)�O�5����T�@%���r���"��ۛt�J&h+5�h �����*�'�p��M�IiD�a2��o�%;)P�[��x�Z��X�g�.��J,D6vR��m��#�8�1S���D���'��;����?��QN��E�k�bDW%�K��Kٶ7e�b��0��\m-4��9�y����Q���v�\�m�{�X���o�_���a���w�rkgQ.0?P$�Lm4q3Տ�1�8������&�YW~� Ouy��G�Ůw{{̦o��!��J s}�gLc2[�%kYd�"�	���q�t��R0K���l?��B��� V~*�bO�Jچ%�U�����H���'��P$]?i�Q/��T���ڌ~�C��D��=�P	��5��*��x9�[�I����J!��'@��J�n��*� ����>D���J�����i�������$��kB}��>���.|߿��~���n��޺�%K?�E���l��jyVEQ�w�R�!�gӧ�A������ꥯ�O��<6E�5x�s��fv!��zC1����G��]�fj��aj6Н����0�L�{��Xp���u�l~$����ݧA��_P�,�˵U���.������Hh���#].(�g�h8 T�خqy����&q�6� �z�ܱ�9�@ò6j�F��ɨ�LL�1%j\��F����W��@j�@T���Drߏ�/� ���a����������W)Ľ�s��k�s��"W��Y�q�?���6S���ѹ�~���bh�z��5����9�'�2B���4 cN�ol6�%�� ��T��O�����Q7Bbűu�9U���ĳ��;�#h/5�/�>��u-Ov�쁾�a�r,9��Oa����r�ɰ�#`��A�X�rҁ��v~j�2�*�#�V����w����ȟ������xV�^j~;�����~[J�i ���_�;d�z1��ȗv�J��(��lJ��ϓ�KK���1
�_+	\�����E�T��4�G���[�����Ϩ}n�����^>�#.8jP�����"F�0���s�]���|Y8#��M}*��Z{�6�9B��`�a6~�"B�9��է���ɷx�Y�֬�Dռ����!�F�?�2���L�E���Q�d�j�Մ������U�T�������)��c�.?z]q��m)�E;��L�ڴ[Պ7;�A�wb���4�'F�+�!��N1�&��We}ܟ�9���G��N�ܗ�=�FfVK��0}�~¥1���{�U��'�������7����B�y3��Lă�XԸ��i!ec)!�]�d�eo�޽pϘ���4�)L[�Y��Z#j�J�}�4#��F&'��$c��3�k�[F��>1
��SpAK��L�EA�LIcj�3�/ce�Ä;�h���ڣ�+K9,�b�Ƅ� <�M��>0��J��ǽI*����Ux�%Y��S�	���������.���b;���_�4h��Y�u� ������+���<y5��p)�X撅��q��*�S�VE�\2��Zh���,�`�H�;��o�K&�G^|h�]5õ����K���>�&�o��R@�1��!����6��ݢ�=i�,�o��11�+nV�h<1�c�f�Do�S©S�&�K�'�=�i��Xkb���Zxؤ��>ݺ�gT}�R�Njӣn�ڪa3��Z��=ӄњ�A9$\w*�6?0�DI�/D����^�T*��_���ECTU�@��w��o+�B����(>t�ÍLjp���p�أV��`��ji����涍�G���go��B�@sH?�s����M�)�{�8��Z����ZY�2���:v����������>\<����'�@n�j�R���נ��������B@"v,U
��G�^^Sh���ޤK~9���� ���Y���lB��f��wA��!gˈ�A��D��<�.��u-��	ȇ%\_�XM�F�M�l���`j�MC�&�'��%���=���Q�����}�ض�e�����ҽ����Cs� )P7W����F�<,
��{a�w�-���Xٿ��4T���5T��v?d��f�HD�ZYA��<!T���N^�#�x�5����y�X����H����v�++q���5|���t�ڐ��C�M��m��RM�/�F�ȍz�$O	< ��s�X��d�-�X����.2Q�gy�7���G�
��	��aRDokJխ\:m�|k���@22�^��h_�JI�!Տ��12wʰ6�a��0G>X���e0�{7*x���a�Zi��g�S+�K��W�+�"���L�ދ�'V�Gn �ģ�i��Q��:⡯�۔x���"�+b�W$2��V�\�vITuf�Gni�����tT���,�٢t겧OC8��=�B�|i5N�}p�g%q
�����lZ��-!}"{��Um��|聞�y�^�l�$]F���:n��4�)l����E	p�N�~�Rn��O�]Gw2�*���m��@�aw;�-�K,HuA7��C>�K���m��[�,9��XZFO��I���n��}��H�O�]��mJ��U�3x�8�O���}��.��6v�7��<�������use�C��Z���?���inY7�7Y��90d��>���k��bPx�p��f$5����e��
K5 �=�����B��O���Z�Ab�Wbk,�"?�d�n�F����s��>��Hܶ��e��EA��5��Ø�ǝ�d�s���;������).m(�R������Nc/
l����bJM�.�n��1�k)Ӑ�"QRl�,a&K�<�fJB���������.�0p����G�|v`�O~i�m��:3I�]��7G���*�Jӿ��I_L�~�Xd�6w��{�cE3�Qd�攈�iB~�ʼ�U �R�ǥs�O���-�RB�o'�;rb{��-=�&����KC7�o��<�l�O�t������7��!�ω�e�/��3���v�-����	$
�s|u���<G+=�[x���	L ��q��l/�3n�^�֝�8Fy[����LW��z�/2�����0��e��"
��"�����λ�}�b�j8-�'��|�ҍ�т�X�����r�.eQ3��G�o0�o4��6�-�5��R^��v��M,��%�¹���@��h�3V ěɞ�4�&ŏ��G������t6LW@ԑ�+��c���nؼ�
Mt�Ȫ�2�UN5s5���LH��6�\4,t!!�*A�	��v:��8^B}�+Ѫ�b}���}��+<�L�5�� Գ�C��pd%̋R�S���WB�z_B`�'�ּ��%��'Ƶ��|s�']z �Ϛg��9)=�����H���[�9���vT��D웫�@L�IOh�tI�������5����1r�;�, D���?ή|ȹv}����-�"��z�������[���s�u\���_<�:�R���6Z���_��l����E�j����P�)��
�d�p���J�*n�h�2�O�P����S%O\�sX�c�Ά5���	����to��$፿��(V�i��m�͏����}��y9���t�0�:s{���#��ѳ��� Xop�GM��W���, ɬ��������7�6���~��ߘ��@�H�M�B��Ϝ��=x f�q����C����ֱ~�$r�����uӭh������6py�C��g�W�	����
H���� a�ݫwN��fe�����ݘb���|�h�Ҟ����pJ�6�ĆR�VcGHF���n�]����²��~�l��������!��w_`��99p�)b����1t����r���u����Ų�g~���N�ŕO^jY��A�٬��O
�����ƬNį93f0�Uu0E3����=�2�� �����HJ@M$�Ȼ=�i6�i_��}�w���녲�-�t��ƌ����(�@\HC�P���Z��c��,;�?�HI�Un��!N��߮��:�.�y��!(0�����
���I"?�--'��
��v�~�.�� R:<0��*�9X�>��̞�����vV����6*I�7k�N�$/�m婶����\@� P�Q	;���X�n�
��/f�eb����������#�)��GQ��1�R����kU�6�^��M�}Q\95%��U�|%�8u�'TH(�y�㪼��E����[@��\����$&�W0� �<��B"D@Bf4��b�P8�ZԳOh+�I�nt%�p�o#�������郲_{�{5���T"&f�Mu�H�ﻜ���%Lz;����}�ٽ��z�L_��t��߈U��.(�5�j�K]{z�L'���7{�
���(��ft7uQXG��N�F;��;dm�1�G�����,��9����՞���fȄ�+��ھҟ��QCN�֭����$Ɍ������}��1�`7&�H��:�T��*F^w�G�̋��j�V�w��1�ڒ��I��7�JV�9;����(�AG���*C�̦т��e�L-��tgU}�ݑ�w={��d��zm.�B/+��R�*@�+�E��lE`}�}1�nfĶ��Q5p�=9<���L �n,���ZO�[��P]����>�l�a=r]+�*��R�9c�P�zT�٘��s&��\:_1���4�P|�W�1���N���æ�����8Y�2�e2�ƖL2��p��?��
�lzV�&�aTOf��@Hy�k>|ؠ4m�&V#�=��3EY�C�ވ�L�sL���D����U�X����.�̻?H���lgN��xq�Q�*o�f%��G=��l�Yh�+�S�f�g����1�s�=�+"v��1�� P) PNL��f�����NBBWC�G���ɤ�L����dZ�V�$�U�B���
�1����+�q�Q�W&���v�;̺^"�1_����Þ%F�<�Z?a�5��쳀Q���'C ��~Y&.1�lp	h0�o�}�uOHY�c��V�kC�3m YΚ���a��R/п�w��<�M��^ڇA��2�H�\�	b������rg���d�p.�!��I7� �Ou�=ʿ��
%��>���%N���,K^�cڂ��:�<]yl�}n_����t��a�9���dnNh��d�+2y,	i�)��V�v��
���V\�bl KI�%YJ
��=+%OMGlt����e�F�����f5=8!(e��<]�DT�/^"�w��@��w���Y.@���c�?,8"*���|g�&J��;���lC������9�r֘�o��)����J�v?���.3ǈz'.ʮ?�n�{��v�?�P-�F��t�$��������)�z��+t���3�A��ه?gg� ƻ-�NG����N=~����(CV��A�o��lJ�e� b����}E'�3�a��B)�j�FV���N\rI0�>U���|��9��W����T�����n㑲���n��\7/?!�iH�[;�,*J�M�&5	���3��Y��Y�D��q���c�m
yZ ���[U���+���L &�P�V��lL�~�ԉUE�@�D�N���d5��t4�~�kfw�#D���֧���.x2��U7�H��0�Ʌ�7��?7yF����}���[�<=���З+�P�j��^�P��s�	j�[G��}�S�F�h){�Z�饢���sY�YX[�.�*b�ԮhT{�g@$�t��8V���/����U~#ҳ�����U�&�q ���`�v�`.C|D`�5*}ooOo�<�/ .��x6.J9���E��V<%.��#�ܞ��Px��^�l��k������B�����)P��-�AK��q#ҿ/A���N��?�"�͡����i�$ ��.��w���h��{쬥�o�U���y���Jv�c5I��ȫ�;���%��)&�
����:�n&RQ�-5%P:J�^���I�����Xu����r��Vp�!tZ�-�����Z©t(�XZD�W���._%���A���W��ꋁ��������D�M�X��F4#�F͔�I�"�;�+ԃ� -�~=���]>�r�ewߟ$P�֦���q�	��uԳ1��Z��_j�;?[D*���2ۚ�����<.��;jOZ��ޗ��I�g��
�<��X��V�pw����@fu��@�'����%1�b�V�`�8]��i?R��Qr=��8�����n|Ar�� �wV��7JX�`HR�D�>H�l@s�w����W{��~�kF|-]�<��W�R�8}Y�7P�ͩ��{[AM�c(ߚ�g��g�H���}�/|��V������	|DO�}`V?{<�S�Do�c���3�ߌ�(V�%�݀_d&��$��[R)�j$9�g+�;���� 	ty�H�Ae���#��}qP��O�R�Y.�����}U���������r���?����{k�)-Ҝ��|fK."����'z�?�_3�����������q���*��i[t�a�������������l�8���k�n'����$!)�n����JEw��B�g^�d�D�� �g��,~���W��wG Y<�gf�n��<�1֢�J{Ef���K]U�����Kp̋NDA�j�,��4��ͩ��TH+����;K<n��O]�Db��.�}~�슇4̤�v�� �8	�fJq}�!�A���b��}�q�����D�M՞�L����Qvy=���d8.����u������k� �XA���p:=9N���C>��CZ0`_�7�ke��$|��A�l�2��iǵ��6FK�9j��BJ*Ю՞��݋�9>R��+&~��JR"5;��N��������`�����yd�nz���G ��Ey��gl-$�;��E��׏�	gV?+�aqN5^JVO�*}H�|�|��h��n����K�.��0݆&� %��I;�D���W��#K
���E�~�p�t��!I�?��w�)¶|KW| O��iHC��R����
����HK��X��)����5���> �W�/V��J�ܛ����Lh���X�!�`hŝ�����Y���(s��[�"8`+\.�+��c������U�@f���a��W@���)t:�������*�$ؚ1v˔/}��6E�@C����j̊u�W�܄��z���J�;�ǘA z(Q�Z��=H
�3+K�@G~��6�i�
*��ވ�̲1�:�N��$�� �t�_J۪1����Zf��(�.���)�$�np���N��7W��v�r�I-;qy�&�]�KW
�|>B�`��3��9�Jo�
���QD��`��µ��?�~q�W*�/gC�m����6��1ʺ ��J������~V,�i�h�����j�^��#��+����hC�
��
���$vL�f�NSW���@	�05�z����J�D�SeߙQJ�\O��N
5H�|n����1��x�	{�ڨ���gK����J!�W�45r��!�����=%ey�����a=���Q/��YKBgn4�Mݽ���m�y*�z�'\��·y"����N���y�f~�>Ld�i�l�<O�}.x+qk��x��٘z�����1hj�����߫�r3�@�ر���
+�G����A�K���Z�w�&8����d���+�t�D*�g��z��T��9��>�0��#�f�W�+{Q�P���9�7Ttx�k�����BV3Z�!����^o��3Ij�S��|��q��҃��5F�+F�Ν>*�z�QE��i���sNK�(Ì�s��/��Ӕ�g�F3rw8��8x�'�K_F��F2���\���ЇW�n��v�qo`�❲}���M >{��M�ʤ��U��_�XF��y-���:f��gӄ�z�Ȁ��=u-V���b�!|��W��V�a6�X���i�b��_�����~���K���x�le��=U��%�T�O݉S�K$^h���l�צ��u��4���y����Q/��p��@v]�'n�����W���h*�k��($G��_�\S� ���XV�Ţ�Eb���^���"�C�Y����a�A�N�}���0EK��̟����q�>����%fioq�|q 7�W�	h��Ѡ[�麭e���Q��JF��[���)��)@��-���2t$�qh	�(l[��>+7�'<�E�Ġ��'P�����^�P:�~�6�X��?_���:�1	������0+g��q!(4��^��烉��_��נQ��xo8��\/����-�@C�+�݌ƍ�I�H{V�M@�k�=e�Mo�I*`��5���uZ�T�{[������q��I>���Jm�2Q�67j=6%fE���U��ko���ۙ���Od<��	�"�2#tP�z����������G���8"�'���4W��Kܝ��~"�":;T30L����j��:��'n�֒bL��̣��#�#|$�@ǲh�ܶ\'prб����mt�q�Z�[������>IC2!#�3���DmZ���N��;,_Z9Qޏ��+��OT&��-c��U���dph�R>�1c�4�bI���f��7��[�v^$v�P�l� �_~�\��t���V�ä�&�,�x<����WÇ��ʝZ�j��� ><�7��kӚ O
�
tCT�7�c��I����Й�!c�6�vBC.UH�g�yi�ڰ��t�����	Z�p��/z�������E�T�ۯ��^ ��
��k��X` ��bwl��SM��TG:��k{c���PC��gt��?�O0-�[DE�|zG
���ǹ~��D^�&C^�������ȳ�J�1��7xpC�:�~&��ie��J��
�\B	/���9>G6m��2���p�4e�ٺb@,Wuƙm'E�Tr_@����o�&l5����a��֧��e���ٰop�9X�kC��՘��yb��"���bXT�#0^�18���́���4,���i�	����{1Q��P6_��5�?�N��g�)�ů]���"�Ox7�G{��SeI�n�Ȥ�"ķJ�l#vM��$�^�Rs���Q�utu��n%�_��E�����k5(�̥�h�֪S�2�U����P7�	.f���h��mp�;�>Z;4m��n�o6�<c'����h�^�[fi�1��@�쏨�އ?jK���t��y���]�9Wb�?�ڥ��[��mx����AB�̃>���9��@��i��_4�����6�of.B���E~���*qhø��&��#�+���Ŵ3���6��KO�ebs��F愸$ڠ����f��v��t�I:d�W��=ۈz�Z�>������ߠZv倅���O�������aq��HH��g�R����r?�'-ǻ`:���o�?�&�����<��m�P}���r[bsH�´��h�{�K� �X����W�4Ю*�Ca�<h7L��]�5d�,��+@K�;b����\<�j��o<����X�G+`��(
���y�ק}��4l�"��>-e�.�������v�j��|���mO��'����l.R'��n�s�����q��H�����*V��'Q m�|�J
��)~Y��\u�c6Yt�5�;ȏb��{ �`�6�����K3�5�����@3ۼT
��p?&�A!b
=/��k�`�V
!0 �_R:�JI��� ��)r��W*��]Mb0�JQo��uQ����^w��!YF��]0g���3{X"�S=��@��^��2�ß��Lx�$�DFl�˷��.�������x׶���^�ud�_����!AP?	讁`0�$&�� x(ϵ��׍a{C5o1���T'v�����v~���]�*b����1�$�g[rI��q� ���G �ݥ��@��vL���iN�i��|n9R��M�-I4
��:��l��$)��X���՚!\�Ƒ���^�G�R�\���X���9v/jl'��$�߲PM���w�m����rW�ؚ�kl����=�~.���	�M����xRC*L���_��*�([n]]�Uv�|��pk>�WKʽdu]ؠ
�@�[E�w��bԭ$�[�o���x��x��a�gF�����@���(أ�H~k�jr ��������6(�R:u^�k|��Gr�'�6����Tq W)lR��qV��t�n�2��'��|���C	�$���q��,Jq��Mz�=�f���n~1*%������˪
k�Mr�s�Fe�_q�L8]W%���n�葖d�xo1saie'��Y�Q���*z�n�H��j��*!��h�y�Ł�i���jԺ{8K�8����
Տ;���1g��_�^������m�g��/�.��L/�S��q�2��m�M)��m�b�A��P���N�t��q�B&�*c�\F�F�l�6���i�����u��!4J8�گx$�M0�=n��g���Ū_�Z%�/;���� �z�.Qrn�����L��Aa�4��G�8V�Cwty�,}�<6<Ύ?y�Vr�V5"�~�)�{��xTጪ����ռ��5�N��'�������ϐ�W$�7�60A����O����Jq��F��� e���
V��x�4��W��A*���{*�ج��|���A�4l�F�(��nSg�F�ճ��*�>�EZ*���1�֋�L��q.�Fo�J� t���p��#�a~�?{�!lʍ�א��2Z��;O�����_&j��!���	:"��R4�;҃Nb�m������(4.6��i�x�V�^f��b'�@1����Q��+�Ǣ_2���2_.�9v/���;%g��['g��tJ�3�ޖ�^��|��~ٜB���Xf����딎���ղ���f @S�ǰ�����`��� C�1*���5
}rq\�<�Ϣ�*�;5���!ô��Yd�h a�����c� �A��~��\l�(���w)�Aj804�i-�F�G���멠�6i���mc��կ��X\�y������"��Ӈ�¢�w*��`�X�L�@7�,�@� &���M�d�-{�/�O^F�E�fuC<��<WB�1F�r'2�	��s]����Ҏ�J���oѩ>T!��v>;x�$��8o32�^�Z���o&/�z�v�\���tO��ׄ�۔�ԗ��ܙD�U*�f9/��O��|� SL;*���4���G�uB�]���!������.Z��{K��{�9LH��X�fڐi��� ��d�';�&;�F���-۔�ڊ����d�V9+)�d����yx�H����V�[��̏k�+)�!B<n��?��}�N�z�~޼
֐���T��a$����葅,�7����I'�������N�Am�U����vp��`c,��2��Z�|Z�Lv�;o����s�'�3f[�魇��K��::E],4^>�P�n��r�w�bF�ݸ��)�h5�W���Ia���_���DYp?5���G��.қ+�,��kb��j�e���?;��v��Zk�"؜׫ߧ��oYUoڃ�i�Ϫ:0,yĔg�s�L%�s���=PJ�A�z�IN�3��Y��~t�y1�4��:ڲ���4H)x�0���Rc��E0����eU��񺺋0�a��סEL���Ft�R��
�������l��?�NW�������s.0Y�%�aF�<�+�F[��[.��02���L��r��C��l��&���%���+���c����&R���	������9N����2�T/N��Z��(���m^|�[��CKs-�K�	m��,]� 0F
�<^�h�	����aF�[C�"�8tgJ�Ȉ���W��@��v�%�ٶs��U{���x�p�Đջu���._�b�)�mװC���`t��@C���[Hi��҅x�����[�1bk6�7`����.��x(��ޞp��5��Y�B��yݱf�F����2y;��Ө��\�Td{��g���yWDzv@�uFy*+��V����%Z�0��@�Pۗ�RU�z<���zBq�����#�}D��RՈ�"��*�uQ�mz�zм�;�\maR�!3��BwҰ���}0�',E^�<y����D
�HV�]�����2��_�5ޱ�L��N$*�,�����2&���_xa3�}�q��(�욉�?�/j�f-ց|��,P��\��D�^'g�u�D���G�n�UX	�W;�-��w,K����xRY��w�1���B�N�~������mki�1P�3E��N1'N�t���JE��bw�E<���y��]�L�E>�.#�僩���mZA��03��4B�x|:��E��pm�D���S�S����*{�9j߰��^d�P}}vU��!�7.���N]v���	s�p��-�f�h]�9����l/"��7J�y��H[�t#����6�ƴ� {pW���[H!���gqiO~D���q��������Cޚq��"��H����7������s�Q�9�;3z�#TҰ�&����'e�w�������h�Z6�FPh)Ee�^�U@~��?���,4,�9�\]��掏�&#��a�ŗT�=����g�ފ��Lj׻DIE����G�^����S���>��I�_�H���,V�2a꺈�R�z������̯W�l��͝+׽v�w�+��t]��s��%N�w��[���iqW3G� �x���/�BW�B�U,�fR���)���䯯�n-@uO�a2��3��Ȉ�K�a)FHE��}�p+�,߮����f=GP{ch����^�x�����Q�ͬˊ��,<�د�κ
,�2���f��R	�q�"V�>1�a�	H^S/ �.���BS$G�|k���?n���W+�׎���b(z:ܳ,;�Ư�y���l���<�G�܂��W�p��#���@j�!@�V�e�$������dywb�8N���6ONXbq1�� ������V�CJ�Dۆ����?���(7	4�^V�,�#w�R:C?��,#�T��)&�R$�v���X���9����`U�ح�4
,&��ٙL�\'���3*3�Qs�n�-&�w�a
�Y�?A����P��j����3tA �[l=��>���r��\�L Q[����u��/Km��59�#���*���˨D����N�O,>m�J�L9?�L�]c~�b*�b0��#��"c8҂�#8��r1x����o�3��-d�0 �t�:�(�����U>�Ҥ}6Ă*d I��_�f�+�ϐ[N�X}�Ǝr�9�ʍ��$��71�I��y0s\��aAx\���gq˟�5��:��ۻf��`�ղI J�0�jἴlUa�M!���d8u&-Z�9ss
�O�=Q& L��ZJ$�]��c涑ZRoM랪�n̑x�|������#��ۼ��T9�_����4�-Fƽ�ƱbO:/ߓ�g��p#���]!z97�JK��=�t�����������:d��M&8^̽y��۲-��r�I�|�f�>��.Xi�,M9}�*�>$Z3xh�M�\հ���i"�\���t"����}�������ےs�xH���[d2�8U�cPI��V���2$W�<6����	��}����=<'Ԩ��Z�o�^�3�t�^6/ͳ�V�cp�n��%$��b�/�\�lf�M�c��Y@f�M/������r�ƹ�uZ�N��!��2?���V����'�(������
����A��2�r����"��u�]ӗj9}I��}{�g�Y��,�vj��>�Ι$�#���h��A��$7��YY��4 {sA��,�KRԊ�]`J�E�+�e�N&�{s:D~y]:�/K�j�yi=�{�{��Rax��54EKL
�*��E��	o��Q��6Ǳ�%J]���mdCw�9����I�^6�����H'�@*��"F�C��N,�lM\E�}Q�J����3K� i Z��[E+PoM�9�j���v���ɖXG�AM���!G�d����)ʼ��c�y�J}M��#����ar��幙���!��t3���ԔW8DŬ^�X��)�!�t�!�̞���(��A}+��n�㢥5�;~-2�����Z�U�{b����\�D�i��}N��l�e&�y'��j�*Yc�ǭM��uԖ��ޖ�f���O�_�;�D���a�����x���7<u��K&��-	t��0�
�iee�&wå���
ZbX��u9�dEw~�i}5Y��j��J+�V�V�H�F��#�W����dd)�8縒xj��$SIr��/FHEN���Z����B�S�m���6�@m"����, �����4h)v�S�ƾU�n8�9j$�b��"ʩq�!*��^�r�c(�X��_S�Uj\�����FB��zJR˪0:0�OfG3��s��:��bv��\�>s�$C���������e�Ss'la�m ���0�3h9��;A��D��go���z��`�7��/l1�O3�����"CP�&쑾�{`?u�0Ens&H�"�8=�g>�����5�>e����� �B'��[dA�o�G�s��b���	1 &��'�gJ��#��.�F�#�W:,qX� ����U.�r([��"v p��J&u�m�[p�ٺR��#���j�Q�ˢ�dU����Y;4���s��w�"&{l�_P�jR���l#�l��ڙ@����9����5�f�s�<;b/(tFW����Ŭ�oa�+�}�_��j���~R#9J��ǝ����.�ZJy���p��Hp��ߋRmb��vI�����g�kĒj�hV��ff�A0'�@�2�ixJ@�k�T9�b*G!�=���3����7��I�,Q�?/��9$�+*��'u �IK��.g�i�7�i\x�ȇ�m�up��
,@�����~�}k!.Ǵ�7S�ב2G�@�����9T��Ԍ ]��~�A峾XՅ�ҷ�)x�嫾)v��q��h:ݓ;]6�7�#�r��()Xή��W���G�䶊t݆{�N�,�ɰ��<�7Y,�����Lt`6KK����Y�������.3�Bџ��03�$�v�2ʥ���m��I�U�0���lR��ʾƄCfdye���	�7�x͍փ�L0��wC#=�G*o�|�G����g�j6�����+9R� �b��{t�6��B����!�3,8\���NH������D'z��p#��q�b �JIk�#��*D#x�x'e(��a�=��3��Q�=r���2_^w�♴�9���˭�G��NK�����4z�&R���d��O�%�|���_)w<��k���L�	H$Yt�����ǚ'yPb`�fvi�y&��<S�����༇	!����3�P��9B$ '2V��h���~JK��H+XB����ZQ��Z�1j:�
D(�}[Kk�ޕ1=���n���-b:׈���#[��yrb^�La�^�
,E�q)�2bX��RgO;JI�.g�Bh��݉�� ��*6���!��>�[�e\ ����f���&h9ԏ�Y/H�,ę�`+#���Q����8@�-�2kl���附�kY(��ʽ�U�9�6^�YyG�Q,=}�]����=��Q���bm:���wb�`��������1�(�m]7���~��w�owT�o���2��uy��a���!A`��*��WѲ�5�"��TG=x(�p��S�9a@��P��}�����Ǫ2�����:$2A���x��_x�1{�:�ȪXl"�;`M�[k�Ɇ�����8��]�Ƨ�J�JQ+�`[|"Qeңx���_��\(Tu�w��͈L��4.��_���A]��ɴy�j̔�M}w5i��/�v�nb{�+��I�:@Y$���o�1���x*��m�T��rEȸw�N�%�D�m?��"�i�vԮA!�c�B2&�k�i��(��
��`4��-���� �WL�ȿ^U��F9�J�ڸ��&����Hs2�{Bj�G��,����;��+2~�Ý��j���v� �gl<'���%��i6h��ʁ�1�!5�|���,�;�a���
�Z9�� �{�� �?�^ſ����1r�a�>^ �ʵSR|I4ˇ�S>[J�D��х��WS��s~�����1�q�Q�K߈S���r�`�ӓBb��{�t}�9�w���_rwh�=�OT+57���l��'���\��&��V�t`e��w�۳�,(���R$]A�H��������F���S��f5��-���v��Yo���%�D4� �^,^������i���5%G]g��$����J ����U
K�t�zoers���
���v\�L͍MJ`)��#h!]�lf(�>�@c�3|FN�]1��`Tp$��|Џe|-�P�Z�ET�%G��7Hh.���JR8��>��s>�uOe�B�Ix�U���˯d3���Y��|����q}��P&hX�����Z��@X"D���.%,�@�z��(CLD�^�V=/Gr|��U�W"T�־�dG��V+P�J�"�.�$�ƾ���'�q�50�@�`g't8֐9�q��d}Y.,O���:�.C��G�:��㖃��v��7���h)��/�U"iXX��טgyt��5�3�!�;d�rb_�]@��P������Ľ�K���lKV:C�*+�C�S�m�ϸ���q�W�X<f�_ʦm��ppwUա�LFj�祫�Ŗ���J�>U��A��t��8=���(�z�������4�?���AE��I��-}�,����|���QP��a��
#��	��i~a�uj��'�����c<d�AE������`�(M�D�۠����w�K^1����3�۴���-� �����,��~Ұ�	���ˤ:vَP�[��v�uw+^*�t��f�d0PY��\�&1)Kl�����?�L����K�������&0��@=�k�U��xә�i��B�kB�'�*
9�R$8�*ڼP��-�	rK��#���Rj�KOP����Jq}E�z�?�W��D�D��IX�Ԡ�� \i7_eɩ)�o��9~sPnL`Z��Q�-PJ�s:�%Sѱ�/�J���O�MS��\�:
Sr@ɕK{��o�8$�}l:M9��];-n�>5I�ǟR���,n�W�m�\����C�WT�Lb��K}�O��,@=Tzғlw�Z64z���O�ĭ�X��d�J`y�-?�X����L�3ݍԄ+6>(� X��;����ћ�fA�ۚ+�ϡ�q�.��@��Z��)1�E�3���o	Q{�"F�!NY�2�n�@�ԓ �+����r�v�7�	��-�x�:0�����D��Ů��f��,�ws�H<��\���7�@1���Mppm�^󕲔"�igN]����0]}[O;��M�8�3z�'f� %^k��sO|;ΕB�_R7�mq�/A�C|<i�7�H�5B���&U�\�)�`:��D�ϛ_�ҜϏj4��}a��y��m0�Fu�T�3�Pȥmv���hl�	�98�W���s������9c�������Ri�������#����s������L*T0>T�۝v�$x��?&�HʃswK�����ibD��ux|R�p@�w�,�}VO��a��Vs�2?�p=~� e�:E�	��ۊZ�nK��-Ҥ)���5���l��Q��ȷ����Y�8m��w-mX���4X����L���ȐOT$����tSi���C���V�e?y����#F��.^��,���s�Ĩ�Xp��
�:�	�B��H�1z[y5��E��.�����Fq7�ф�
I/r���Y��Gy�G\X�/U恨c_���lO�A^��$o3a�����K05g�FV·`DOo�j��u�� P	 ��&'7�M���y��XL�rE��t=�5�}�A�e�j���{��M�(�ʁ2R��*���Ф؃�C3�~2����T�u�u�^ȴ۽4���s�3��QH�)�=����Q��ҕ����T�4��V+>�Jƀf��\,'�ťT�?Hf�N�_1*x�}��umIu)�;�)Cb�GE�`V�B�3�I�Ǣ��e����5���g}��H��
_� �9�j�FTwF8V#��E7�=�%h��g��xv�<E�z�Y�쁧>��]<*�]t��FF�9:]x"~��	��޵�����Mi���	}W�c?����K��n��Nl��7��U�F��PL$�q����������}���ss��R"6�Ȼ T`�Hv���.SI��?o��D;Jtw�����C
b�m#���d�o��1e�P�+~���LHb_�ӊ�u�12�E�d>D1p6J���^��+w�q�9V��+>��xj��� ��N/f��Nx!%�|�Aբ�]ʲ1{��6"㫘�=c�Qx�V���
�FbK62m�"����ϣT����Nҥegv`�e�6����ҙ�q���K
9��v�q����!(i���&b�.�M��f^�hG��:JQ
��~$,���GG3f~��ז��>�'�*r$��]� ���,�N���97%��G!"G��ĆG�WF%�Yn�$���\�D�QrB��2{����q�5+H�e(X@���E_�zvm	-�����g���fXN>�� u��_[4��E#��|)�C�DT�8~�&�[��z4�T+ⅎ;%U����3�'�*5�P��V�m����{}
�J��Vy�<��]D0ಂ�T������.�:���'�;���n����B��+�������l�1��n@���@���v]��'/$��b�Ɇp��{|+KD�,�1 }A�e���L�3��Q�I�`�d5��p�@ N�T/&����%� �m���x7��^@w�f1�Q�\u@�U��vq�X;w�[��ʺJS	���YL8p��6�Z�E����/���o����/95m�v>��⴫2[��r�N&N�`Ք�:���p��� �*o�AL��*�N��^V�J��LԦ�0$Q A�$S�yc��yQG�&-+��ӂ萭��k|�m�S��k�0�+�~�~,����c"C�!�<�$�T��z���I�wcD���ֽ�i��S�k��[�!e�N�h �r�R�������Ɨ���î� �Jc�R�Kj��[	����S�s%)�� ���;���޼}.l6�D�jEScm����a�nϮV����'�$<���¾@�}�kNN@-��G����͠ �L"kP*��Y��԰���?x�mtW���Le���s}/��Va��!/r���0O8�����?R�)�����H� ��q��t�@\M��NS�귾Ə������:W�8��.ˎ�x�y�0��ЖL��&�������zK��!ըI%(i�/�u�G����ՙB5���)��Ǭ�
��D�߂z�\J��G_,��g�?�<�+�{�a7�{N5�%h^�Vk!�?Tt&	�k� ��j�N�.�l�Zш1���qDk�$q�?~y���%q�V�:��U�Q+/7�Z�l���T�<r�*���l��	���=�����T`�8*+�?]�3�c3��y�	�Zi�̀؈�s*��8�oO�i�S"ޒi$	�n��7��
��*�ވ1��;f#'6���Ι��1�M)�z�{�meg�uZ9�x�t3>l��V��:�;? @=��^�m{u��G!�ce1ٲ2��
G�/FP%�py�����5<X�9̻ꈹ��bz����t�� K��gܻO��F7|#~��i��+J4�����js
��>�L�u�Q���lGNN�Y��l���j�wn�s���#��M�����07�V�;N8��'�JY�����)@4�Q�ݨ:�B�]���&{/��&Omi��'}����/L��9�JԎ��Ш�χ���d��-E��3���EZ��僓'�0zR8LY�A�zT���>���P&kJj�ny3��B�K�E�� �`�;�R�i�sx��������Ta[0΃$Eg�z$8�[u"`�&�<�G�}^�4�����>ԣC�(G���Q\Я���|T�������5mh'�n��;[v��f�f��H�,�'x�:K�n���[m����H�6Lك5�O���6�-�%c6Z���U9��7�޾�4��CD��w�)�z�8��<��f��4�?��H�����Gwi@	 
�px
&Ц���|���D&UL�� 5i�+�
�媞p�k7�\�2�PÚ�rryQ�[l?dTz��,�q�����`�U��Vi�3�Nq�P�� '.c�e&B#Lh��!�UߏR�8����j(� ���Lz��[#_k^���OT04�� ]��jwPM��A:%���5d!^�)� $�-��j�漟�*�i޸��P�
�U��%�]3��i�������:�&'Ƙp/�>lK÷��ء�%8��QJ���\�\��R��=��9�ﳚN)cZT��aA }�4a��������Q�}�E�̾�:1��GQg� ��pA��t���Mӄ����J�e����-}
x�#j"�ʾ��'殻���>�<�w�B����:�: �����n4��LUN��A.�8k���GG��"&rbt|�� T���K�	���EӁ�!�uL\�9�=��p���=5��<�{��Ϻ5���M�N��&rY�'����n��W`m�Z\��[�M*Q�&����;���y�"	��y��Qe��,�_����e�C�Q{J-���`�2�;*�u�D�T) l� ��I��<�k�a�����F��v�뾀GU&k�	�b=F�-���L�+��7��}x�(�܏��Z��5�2G��ve���FE#��n�Dgte�?C�	5e\��4R�Bڏ�Aj�,GyD�崐�J�f2 �V�?�7 ʋ^O=��ڮ��o�Y]��w�a��u�,�!��Mz��3J_���:�����F��w����T���fC~HT�83~0����,o��T�t������l�^���Ýpϔ�����O���KD�z�J1�Ep"+Z�XX���Oj*^L�����J�|5�Q���̏��΁N��mO�KK,Օ	�5�0/~�*ӸM�w�!d��7��I���/�.8#��'����x:�P��T£꼝;�~���X4��R��\���t����� $I�[�z.��d��KT9[�6�.MV��tYdI���_��EH�P��Jtu���/��撊H������T?��)T��%� �����zh]��t��"  _��匫�C�\�d[��j#q��.}������������B�2��&Q�t�Lo��ɹD�kH.& ��	<��/4�L����{�+���$��1>�oa�� g{�����O����#�)e�Y��M#���Wy�N~n5u��) ��.�J&I	ɺ=�Z���a͵T�:�p# p��]�ޅc��Q�����l�,�b�e�0�R}�tn���wav���N�l�<�󷱳����H��Ɔ�d@���p�봁ʰrq/*N���%���֢�ą���RpQ���"�L�W�>L"$b;�\ �����^�No$�k����A��aQ(�4YbH��0��:/]�=��2���K0sF/�gў�
xʾ��Z2�"��U����f�����2%l�.��V`~fDþ���N��U�bp��4VU?#�n�����[��d�����y�-���q1������������J�N�In����ii
V�4��:h��6(66&/ U~M ��e�����m",��Y�w���t�5ɑ��%�WD��(�f&��^�g^/l5�c��_��ku��8��/BK�|8�4p!�o<��(��0YAQ$�ɔ�� 2�	�Shi�������'��~��B���]\�c-��~�(�gǑ�kp�␇��,����7��I�K�.�2 �Rx�*R�X�������k�w�/[jF�f!2����eh\��E�̵�{����i��M�AM����Ր��F�g �����r������p���0/�����8�	��6V���w2};(o���>���6���$!���)������
{�!M��)�����<Є�\Y%�m�A{LX�VY��\�*ې��M"=N{�[�h_���^<��Ֆ�FIF� 4�@���߰�JV��f�T�|'�x/R�K��N=�qH5ȇ��N��Zm���x/�w+~�6d�|�N��l��vC�U W9�������� �\0^���n�|��4��\8�Ԅ˯ ��KȨ|!���s��oҜ�׌�^zv��@�V��ܧ�?��s�x��_ �Pi��;�@[�}/d:�i+�5��|p��F�ܵx�����p���~h���7�/U��/F�%���jDA�1�a{������<T�omW��.�����o�����J_�GF,��^��	�HFQ�OY��fg�{�:l,�`�|�2�.��OƐ(iL�ξ+��e+9�|���=�3�*����0�CD�-w�b�7�$�u�Q,5q?>ͥ���fpg��q~1_��1s�~����(TC"a�P�%��q-�f>��Oc'f�$�s�5u�O�Z�:A���қ+�_<�<��/uoQ�˫g�����V��u��?���Ί�_���HnJMԚ	]��
���1�"��v�&Q���AZ6����!�x;�N_J_�a�����-�	�r�AT����5�[����SWH��ϻq�ܚM0]Uk�����Ι���2��q���	lZ�ǀV��}F��Χ�G���2�9;��Ԩ$\2c
N�@;E������L�%���T뱼��p�����G��~�J�F��'��CZ'
z�:���b��
�t>͹��&�˘�)NGfC`1�ޖ(��vp��T�� �����Š	�g$�Vh�;{g�ș���Q�УL��8�e�2��I�|3E�Q�
!�`b?��U� m��_/2�����agpb�8�����Qk��k�v=�=dQBi�~�������f����=
��ֹ�_f�p�~@���(����0��Y�k���U6��_�yg� ���ѼڳK�kP��Z�A�4���R�,S�I \��D���]+@�d��5�����z�uÎ�-��Z��A���f�o:Pmi �5�cR��O�/�2����?
",=�T,<�������,�����\A�3QL����w�������/��g�t��9��<�W7'&k7��[�" Լ|��b��j�9�M������@V	ŉ����]�8��~��Jwe�6r���>�����DT˵�>��*�^͵s��![�>��7��4��YG�W��K��Q��y�qB���Q`�����H'�~��8}oV��/gHΏV��������D�tY��;�����/��*��w���fu�e�lJ�/n�*~Q��/�U�Y����I�^����ې�f*��.�ohaG.Y�)�fB����m�wb�G}�?~)Ł�.S̓"$$�c��/Z��9�)�����B0I��Y\;S,H�ڬ�k�pS
c��B<�GQ��X�!q�h�ɥm`�J�s�����0Qo@A^��,\�R��(s2y����<gA��{�!�A>q0�X��g{�ݓ`��U�3�DJ⾏�2��O�My���{x52^��hL �r���p�Y�ذC��}��HHU�)�V�T�NY��X��A��[, ���f���u�:�^n�df�q�}��[o��ʟ���:V��ʢ�>�I5�X ��4�L�^��
�!o�.AT��z�q��ա���1̞)���B���[�t�xH_}C��6R�7$��'*�M���5����C�y��F��b��t�lY��~,T䭻�`ќ��e��ɇ�N��@�o��h�@�* ����v;fk�'��Va�|����b��kN��]��l6�	�!�� =UQ��`�	)ZA>�k{�V�?�k�[�}��#Y�{���<���pN~{иD�n�%^R��u}�Eyؾ��&FWE���c�RB���[}��~���v����JĖO;T�h����!2�y׹kș�y��{H�n����:�?Rt�@���������p�#㰻�	�`S��'�_���BN��CC��S��'QY1����$W�����Um5�!ѓ�t��ϧn��Jds%��D��I�0d�N��tд�C��'�����ZV[�ͯ�;�BC�ń���ѭ�2?i���b�{
��!�{�ݐ, ��a-�ݱ�ϔ8\�S[8���u9������|�{oU]�$�V~l�B����H@`��j�\bD���oB�����dBB�h�j���Y)�vz�W'{C�u�3q)�V�#��,�����oD�a���.!���������~,���:�g0=�ϸ�,���?^�hn��V�!�J�L+��7�cѽ-�kWZ�W���Ӷ��"��J��;�s�����H�� &��mŻoܟ����b��n�KtQ��0K
�7x�!H^�HE�k�^k��n�><�P��'����	ãN��ݗ�u�v[��b0���)U���k6`��A�L�}�ODC`����6b����akۀE�7$tR97��s��n~��)
����i?n֥3a98ַ6�(���v^�2�B�$Hsf`t�	Uv��Iބ;��2p�%�栀`���d�F�N7n��P�.������d~e�)��p��䜇4�q�$Eʐ|@�3�(��yügk�8��[>��l�K���5lS��p�x��đ�E��y�ç{�������nJ�ze$ɳ�Ҷ���0=ǔ!���F�/	Ȣ!rgS��`o�<]�&�,(nsN��p�P�� ?;���NBP#�n?PV:�x!�����}ņ�m���S.k�)۱��=6؃��q[y
��p2���w��򾤩R�z<D���@4��S��K�b��G-ow��ƞK��؏������V�Cp	$T�P����c�r�ek�����r37�Zs-�k����y4���Vɯ�Ek��/����x�0R�׍��C6���[O9� ���/d^vWb^�u�;�W�y��S��.�vOF���T5�t�g�d����t�Nc("<��o5��b��W%-� �@��5*��vq鳚� g���'�����p�Y����3=o
�c|D�3)S�ސ�덺Ŋٴnh��k�t�dS�(�|U�CI)$T�J�<֫��a�aS�ũ<m������,@N:�分�~��f��1�xՉT���p�Q��*�Q�2�����:����0ii嘚��e��|�U�������m�5��;9;��h2^6C��Nz��m84d�K�/�[�G�m!-�5�W/ʺ�?rˇ�Z[�9њU�?��m��
v�X�z��P,����*=K�}�V��x�$k�3Mw��@Z���m��h���F����_]��[js)@�i����;d�V��+'�gs�@"
�g�c=�������X�2�T��j�y�E�ymiC}<�2졖����"��O����=s�\ǭ��� �0q]'�NGXg;�l�QG,�ᕣ��Ԉ�d=8�y�9�!��9L~}hp�dx���Q�:֮}I_3 ,˷`���-9'r��'�CK��@��+o��E<ņsc=��;�Z�S\#S�0�w�&����Z�"N�@�yD�F���QW��A#�0�x��d���N�J{ҫH^��R�n�,��<������q:G�f����'^�A��kM꽇R�n���(��P�%#ҷ�|�~�B�@��%���Â��?�N~�Q��px����L3w��������h����o{�n>x�σh|69�d	a&<YeND� l��vʒ�I��:iU��m��k��b���H���KM�^1;�M0� ��9,��ۭ����|F�F*
���'�Dݩ�E�v"y�b�<��uE���$3��K�>զ��%�/D�4ZD�։}qdR��
d�rK�h��l�z��|
����]�Np�J����<��
с;E�	'�x;k�x�0�og�>�z٭�[{��S��͇�Q��O�j	!@��[t	yk%�m�H!*Qa��k�*:퉋cf����ߧ���}��<����Y�?�	��"6q:p�I;�y�;Zo#�Ϥ��zl0"F��k��D�	���CvC��Y��_'J4�"�!��!q�����}|��d��G��Op�ݭ��1@z��n2��{O��>��C���;h��㡇��)�C�>����2a
��x�`�U��B7���c4P�~�A��!h`
v,���NM�ixkd�v�@@��=��WF���b�1;ڹ(��}��_����>��-����A�X^9gn|F���< a��x�ָ�z����*� ���U{֨Tn��0G��-��\ȴ�j#	��e�L��ܞx'#9�IA+~�H_��H�!���pJ��!�@ہ���╀���CQ����N8!zMa�״� �pH8����|�p��7��Z�(.���@��
�c;Uբ5%����F[&-�dLL(��{�(��ķ2a��\��"��]@Qb��q@��|�0���*�)�b�wx���%b�Čɯ0�y���ؼ�U_����' ��5COb��״V!�[�I���Ɉ��\pB|B�^�[-ױ4
�6ƾ����'A�V�4�#���~z���	�b�E:9�d�Am��EH�������m#�/�֛�iB<�Lby��H#	;� F��_+�{m���?�2����7�AOׇ
�M�k$}
�G�ؙ{x�F��%�73G���A��r����Xg��o�e��;��7��x���&�^�<�A"��;����-�8Zw�����G����$4JH�`�=އ�o��I�H�M�5�8٢lx@���׌�s���>r>я�G�qe(w��]`��hw���:������Cg���g�g϶ּ��Q�Y�|��X
7f݊��j�Y�}�F�7Z��5�=���*��w ��bx�M;sT����n���7!+����n�W�q��U�L ~�&����-G!�Qrg��g)l�g�w�Up��|�x8�A�C,�4z��x߱��_>�Ov���*4�a�˸^az�:5�L��N���#k�?�����n[
�g�r����=�2����IP��]��	�w���e�Q�}~�')��#'`J���Op'SBhы�0�
�y��/ �n�b�^i=٩Dtz-�鿦�酾Q��ۇnc�)�_��.�����*�8���F��<�+KF�r�I�\�� e�O`���[^wbf����,J����eM�~���ަ\w@}6�C� 1^T@��T�:ur�VM�ьb�av���x�@�-��3�-�!����{�]��~� E��[�����`6��07��E��O8x��8�`
'\ʓk��	������ҥ�U����L�g]�;�Y6I	O���*��P��N�����M��o���j���B��3�8�e &oԎD��bЪ{�1�7��US�%e>�SA 3<Y�����U����OT�-l�4���UE�S�w���U�0�XK�"˅ ���e�a'hoTA�	k_C��#��B
�b��0'n`����Y�����e��'���堤GA�&Z<�z���������o�'�I�����H�1��FW ��M:�����d����Gh����6�{������duD��y�U9|Ex�ۣ&�Ő�p�������z#�0B �i��a0�ԙv���V�>�[6�%��?O��/�+P� �
0���� ��_c�ȵ��4��C\1��YlX~Q�!������J�K��y��n�8I@������ܿ���3��7r�V�����cP3
局]+�>T���3@�h��V_Z����j�餙MJ���?�������h��(%Xrֽ�g&
�2aȺ�S��2[�{�g?�Ӓu��\��lқ0[ =8�����۪��ѥ����n&W@U�1��~�\[T��(���β��Ծ4@)BG"�M�U����]�V�g)Ó�3��0R�@�	V)�2�q(��wc��h�
��x�����T����[�٣�\�yG�X����*���ѝ�Q*� ��,%�F�,�s�S�T��!m;�G ��������n�1e���b�=B���P��
�T?`�\�������Xt ��$�xaD�e;�,i$�\҉�Z�%����ql;�v���_K���E�@|ưҢi���t�m;>��*�!�a U��tru�� n/z;j=�t�v��{����]l�z�Za3�_�cxr�|�J)?j�A0�w��Pe�ȁ5bwv�<�mL�ǭ��;P�w[y���: �v�N;VV�{�m<�dU|;<�Gٹ�p��K�z@��؝���U���r���%|�;�3ƚæ���A-)�y�!ND���ȳ�/#���`�G4�6o�oMV�����]e�l�K~�/�..�5t�ɗK�l��&�&7�"�	g
79���	"$�����q��;M��M)�V^�39��nb�|��p����Ɠ�PՉ��5���ϧ,�1S=l���L�"�!�$�@�YDĶ@���I���!\Fj�LʦRSI�Ei�=� ��,8�E�dS��at��<����*�� -.v�����H9CW�h�H��LNl��%����R/-���K*7���X�;��h������iBӥ�u�C�/��W��Ś8�ӗ�J
Ƣ3 θk;ew\�8�y�<����q�� �	y�6j�G��ؚ��+��y;�*�U��C��"\��s�dJ������k#"�������a�Ʊ�4�$i�3�e�-n��_қC�����7}��h��:���b�B�a��|_��B��R�Sy �= ��/���=����0�1"%�5��7�i��'B[�9J��s0��i��B���j��(7��c��h˩�c��e��F&j�H�*�=��"P�%o�,�x
4b��/�i�����>Q��%�b
�Ȝ�i<uֿ��i���l�:����KV�"��a,�o�����倉�<�/��	�̄Xy��cr	�C��ϙW������^���g���*-��5�K�kW�zi�o�G���V������e7Чݾd�RX{������O����xn~\�85u�-�}�!�J��p�+8Y�kr��e%偘�Orb=7����[QP���#��ڤp������$�0nwT�d?�+]�L�t#��8N�F[��Len?�!�5�[CWõ�F(��}�i�Z��G�ٵޯl��b�4]��]t �
2��#�mB�*~�%�{��R*�H�A��¦�4�C3�ȋDO)Ӎ�Kȁ�iF����Z��~�Zi�XX�/#��\��?�2�7]��S�+U�٘��̽�ɁO ^��D���0nn^�, SN*�.X�6�� $p��$�j����I��̩NJ'd0*A��=ך�6�� �ˏi�{��Y�Z�u��p	�s˶�C>�.s�f?�k�/��Vw���؛`� JKX�;�&����R��ړ�Y�!4샅���5%Q'�W^�d9����4��h�������L1����g�e�2,��9�5�{l.�r�v���'��A���K�v�+~�DG��&�DG1	�з�p�8�)2�b�����N	�d����+kp��O��6��Ev�m��X)�������D�F�xi��,�O�2Y\�8d=�<�|B<*�>A�La	 ��@�Oi?���ߑ@<88pk���r��fV�c�����8���;q"���B�,�#l�Z��S�B�G�WWYd�j%#m)������=�>�A$K)&'�s�Su�/����C�k��tj�v��+�غ�k}o��o鳈�ƽ�4|-Q�`?O��R郦8��PSH����n>�d��r��4pQHߠ��2�?z���|�h�2���X��Q=�N�&���q��4�˛R���WE
,R�řʂV��øW,`����	1�֊"��OrdM֯�3=:A߲�vV��qדtd@�D۟�(��s��:%q,�I���wx��d�)�Y�E�ӵq�W�7�T�h�1�FE�خt��T�P	~K5W}�q��
T�\�&-�����8 ��Zl�i����w��7-�>��Tò�r�w'��o��\�}���b���mX��kQ/m�C���b�1����l��-�Z�@�q<�kUT��ݗWL�e�U���mT܁�WvN��5^	�.$��	��VV-6����:v����Ȼ1����D�{��k��(�������䫬f|odq��6��ȕq��Z
�cI4a�[��`��*b[qj})�K���"�OqB��k���չU�J�_9 �L�q�G���҅V�}�Z�<L�hb����R2��պqO��X���ai���8���-��Y������4�5��,�?�7��)e�9�7��[տ� ����!:R. 쇋�S���=��\i�D簀��(���VI>2;�c]�?���P )n�'"��^����;S�1/�P��q�`��W9'��!�z��u��m�j�(i\̛��O��O~�(��p��9g�V.,L)uU�C�(dz�Y���\�r��YW6;
]8��0�o���:Z�-v���B]�KH�G>L�n�4�oo�$�9��S��P��k`���rD�/eboD����Y���EcY\wּ+��H��xI?~����x��&�%ǌ�n=�p�ڎ���b���pp�"q��q�G��L>a��٬e2|��d��ua��`�Q�!���R.�0�qzM�ј��7&I�,�2�g��������k�RJ�����Tw{x'U�����?��M�*�Į���B���($���r�����jG�1�x��#"	Z�6��PA�w�q����)�I��K��S��z��l��S2v���F��n�z����ahd5���Jj�Aܴ��|�h�k:x�Xs�0���Lm?U���-�P���J�pY�Cp�H�����-���j���5*)��M f �Sț�DrCY��=�u�bՑ-�6{J|o��/�*F��ȾO�E����D�(|��]�&�J���#'�2�[�nV�4�0��|��)?���:ތZ�����Q�e9���S��:XMg/���A(uo0U�M`�>���S>�ږ�k��EN�ЅH���~��[���H�Y����[�?F�^�O�j�%̻����ƱP��U��Df�Pt���~����Ⱕ���z��u΍YQᠩq�w�n�o�k���w=�-qdW\"�ʶ�ƯJ`��fi���C�
�#Q%p��X�G�Vbʧh�i���O�H>Y�iB�l�&K��O�G�E#���聑p�	v�6�O���a�q�;�z\���C�NI��nE�,;^ =x�1>Y�"z1��r8r��sE�{��������@K�`�:�9\�c��b��HaV�ӽA��lp��|��X:���P{�eߵcH}�H��]��w�a=�o���}6�ST���<R�>��%Էy��ݷ̗�$7��(��w����zyIU�;�ܺA�C���E�yo����+R{N�@`P��pכ;a�K>�e�9��q�0�EL̋�`͆����9L���v��3�"�p�<%�Je��o�M�wB4J��5f�ޤ`��tz5>.z�*��E��8�6�.3y,�N�V�yL�{g�T��g��@0�*«��ڍ�#��I�A�*u�[��8*�_���w(?b�����W���5��������V�SVL�fW]�{��7�#�l5�]c�1m ܘY0�<��+K��Lo���l��r�Xu"��0y�铬��Q2h��L��"�ZW>0��=�k�-8��V��6+���H��c��N��$���ì�v�<'�񜊀�h���ɥqX
A���*�Ї@_� �AW�����htr	P�a7��`�*)�S�CwaQ���E��4kI� ��!���\����kzm,j́	�1׺�>��wؓjmD�,9{JMG/*N_ꦏk���!1x��w�!:h�hӨ�WrJWq��t'���2kG��l��	�M��S���Z�y��v$�V19�j�S���q^�5�.��G0%��<�P�
��O�n������O�Fd���k9:���Tg��9�>s��f��ԭm�I~���I_�����0ϼlX�8� ��-Mp[v���p
`�z5����_-�fz��k�ë�w������[�F�
ADLg�ai��E��j�'�N\,XC�]u�Y��g%��u�t�#T���#Q��T?{�Q�1����㋺��@��~��ncn��!1��؀HXyu��~��RE�r.K^R��0%���'���r6�}>�{�p�:y�aaf�F�d&�{2J��.SR8�����裖tu>ē�`�(�ę�2#	gv�Ī
������O�Pڟ�s[%z�����6�p�?(���ݭ�`�aYNA/g��G{�E�'+|ǭ	�q�����oG�W����`S�y�q0D]��Ba.�NѮ�\��[�ӊp��t�� �~���>ki��@v���a�����Y��#3#�a"��E/(�D�0�g����9����_~���W�%W�X~���b�1ڝ���b�X%����~��"|4�]M�
cHdG(+��s�8	L��9%*5$�P���
�c��h�$[�(��Rp� ?�f<��7K��YH��k��t�-��i��W{j�}���n=^-[��s����~G��/ޚH��S��3AM?:Xu���E6���F�Z�DX~7<Ó�����\�)�.zW�?/U�i�ŗ�W� D�b���/X�i�@���,�ݐ���L���R(X>)��QҨ�7�l^�=ub�;4O1ښI���CI�B9Ov�@=�}�3�)<X\m�X�
�bJE�;l�3`q�^���ٓ�кF�*l"��Sc:�֫��ct>i�e#xw�ڛo��1_ q�P뫆�d���S�_���M��΁�2��)h�w������/�;���Y�7T���mS���b��ч��A
[��/SI�E��%Ө>T�0_���R,�`��!���Y�'�S5�2tq_K��8�0zliA�i����R��W/m�&�^���)����p���TQ��K�F����u�����'�^�w�3��}NMF��t�e1���}�"]g���&Jz���CY�yw���T�3����6
f&W��t�@���#�:Y8�����R]m�s*���0��xD�!*�[�*>����.�DD.�Y���]�_ݤ;���ML9��U%�C]��E�5ʚ���5w��wvE��Sr]�`��)�q��&�4�FcEzLX���E%�c�.'�_��iUĢ}�W|�X��Yț�.��|0<@ԕd���)��N{�a�V���u�a[��Í��b.��Q�rH>~�%2�֯�j���L�D[�*�i�� �&�)�㈩վG�~���0P=���/�o%�f����BH�#���Rm�N-�a��')%<3��wx4qM�D�@���b�ou3�;"�bq�B�$��J"��e�P��F��փ]kC�+�w
���'إ�ぼx`XV�c��&�f��SB\�i���A���|�$��K�U���_�1���ޕHѱ�K��.�<	9�P
�PG�w��䢭s��Et�BjJ5!;EOc%�B�/}K����B
}b�苢t)��\E@�T�UK�T�PK�h�+�����)̮��)����%כO�\����+汭��5ri�H�0��!�3�Z!�̜
����O��9���������C�ņ�D���9\��|�
��WV�
p͜ߏ��~
�B:?~�`b�j�QU4�k��eN�M{������8��Kc�Vl,���!,(��{V�<�����h���x*�$�r���y7�K�sK\
���)���՘HQ~���dLM�ܰ�Ǿ`	�����+	�Q7�4�GG�"�t�n!��M���&) �Q�&&SZ��i�	�N)���l�Fcj (����%�g�q�ۆG:~(��:g���N;�~P�4O��l�*D.�D2��M��'m���:�xP Ɓ� ��K�Q�~&}���c�$����(3�X2�*>��`�`���&mL0 P�f�\����������2D�PM����zz��ko������/��u�L�:�7�9��0,XT�N���z|�Cҝ�`;�����;'�6[�($��aMd��zH�0!��%BA��J�q�7j��::�f)|X%T��U,�#��i,���#�$�|��X|5b(�[Iؚ؁z�LhZ��X{�S]�l�?_
�r�;�ͬ��t.�$�D�%o�p�����%�S�WxJ�vC
0�����Y0"Q����2�D([y�rZ���G<}�F��0j,UM��yv������K�m�)�َl6�S��ژܜ�3a��cJE�O~�i"Sȅ2.����)�yQ%=ێݪ鰥1d�;83\
�-���*5��3���vM�Y�S)4W�w�pK!2�F90��'�ʦ��~��xr�`֋��߆Uw��;߹Hp+\��b������%S�t49{Ek`�;�����-����`�,�y���Ft0i^�p�[��oxm�N����@G>���śOm2�1
�@��s�lt#T��M2:�Ux���د�ٞ���
�M�6��H"rYlz����_ ״*x]�Ls�&ϝ�4H�=���f��(��c<z��U���*�u�K��SDg*���*L��>�y�qӞ�:�B�S���E.E	fc�U;��h�������Z���F�.~�=v�nb����[/�lk��H����M�-�6ϥ���ƫ�� ��`�,��YU�o>��+1x����T�!� ZFK��dU/�����`4��S�Z���/-K�\�Y�+s5��<��hQ��c7�����|��zi5�/���[<nn��LR��LΒ��PK��f�|#�!!��M����H�봿/���i�}҄�9��i�P�;uN��
�������	�*���ֻ�R��3׫����ls�^�
Ѱw�]�����ٲ~�)�W�����Mtv&
(/s˿��,�컕�ř�r������_�	�DQd;b!̂�T�`���B��������Y��[�n-�٨�e��z/��p�G&%<��n�g��1�}���h[:ܻVB�x% c��BIO+(�����-���%pܝ���8NVV7�C$f14�b�ޯ����+C+a�c�z�O}�{$��������m�h���9%x�\7��9"�N�c��U��K�)���WQ����G�"�%e�05.�!�	����H������>��.�� �א���W�.v�h������yPݲ�-�bP��x@��=��O�񙓱oB)`�6�R��ݻ����z�h}��o�8�n�9�=93˅��ܕ5��R�>�!zkj J��ّ��T"Z��D���kA{�B��[c=1¬�	U�I�/$g���E-�x����k,jL2�v��-�n	v�5�#��}-3����0i����/���˩�.�rzM���4'I�5J�ޮ[�l���R��ۙ5(Z�~�3���x1�[�m֢>-�Y��f�$�\��Ͻ�m����F1�C�OL-�h��'���'��$w����t�7�G�l9������6F.��/I��kjyؤR�$	�l�+��tO�w����O'��z*n�����E���n�.��<���bG�wf� 8/S��ݽ�Xm��<�AD =�T����YxP6�����J�p�y�.&i&��q�;�߽LE���{
b3$~Z��aFK��H�e������gf6_�֨��%Oƻ(��"��Ds�|9V�)�t�M%#���6��E]r���Q�4m��t�CA�?� |�̈́�3/K� ��*罐J�!���AT}ڈ;p�D �@�MՄ�$@��+M����ك��~�n��l�.��Pz�x��m8�ҍ_9=ḥ������%�uH�J-�m{VH>6Ĵe8-n��䖏�P�t�1�wwY]{�O$o��&��۱��\�e �L����Q��%�N�̇+G�A�TC����mr�'������=T�#Å)O������)&�'O�����=O3a�6ν�ӃQr��&��]�lx�l����%Tv�7���ΦHC˱zGխ"MN�;�
�dN���X^r���y���}l_g�}V!ՆE����"���cu�Eb���&K;�s}�Į��:�G�Trm2�y`u�4n0S�����X��H*@�(��a��i�o9J������B��Zø�m�����g?�Ro���R�k��-��|~]q� 2�G�ب��	��(�a����7QGp�x1�TJ���Ƶ�p��?��SW��<��f�Hc]0�e.���(��Zc���"�k��9<PTQG*�Y�J.������� .8��QW|IO���!�W$�c9`/����.��S������a}h�E�$��ҋ8MɩB�\:`��>�׻)��bH���ߏ��^4�"�O�zr�����h�M�F]�~lm��˂����3Ϡ��}�5��a����o�h9P+�ۨ��P^��k���h��\��P�����㘭o>�GRF�S:<e����{��8��8��������i����8��
�$�X�"�jJ�A�}��P�=F�0�S�Ln�{.�gC@Qtcpj�8x���ZA8.&&�tª-�"T�U}]
�������� ��Ų��:�i���*���:&�-UE�
�i�n�U�ԁZ0�V����	Z,�ax�g���H�HT/�P��%d���}p�"�u��h���(%Ynm��9<�J�v��T�&�"�� Cql��L��8�iorh�c�zj	4��Hjt�c�N�X��A9;"��AɿYuD<�O(�}��`q��4���>�.:����6�rqu��h��%�q�A�ܰ)Ɏ�Զ���ω]�_�؜����1��1��/���T	�.a��J�1�n�9�*_$�uН�_>�Њ�( ���_`6<�$B���Vc�_�d����vQ~cdK;�*<���[u���D��Ψn�i&�߭X1�>��e���4���P��������Ig�E��>HR�A*a��c��1-)��c"�
������� �;\
$m\�͌�#l�̸4��?w�^�_�r�D&8����w����^��S�R�(R�X����������R(�����̥{&�I�a����W��ް����i�����s�4n���w(M�!;���L��iy�J�E�VP�>��o�.�Ty��.��@��@�8�w�-�
���n��J?m���p�d�ܽ�>#_�|�^4�̎@1P�4�!�тp��,�F�T�(��~�hf���vU��X�� ;���whT��`�gM�td��A�c�� ��V�<�X4`?��V���z�$k>?���ىɝ�}e{��s��ӎ�OXc3�Q[7��,���7B��x1MU�Q�n)7�d���N���ۏ�,�g7�M�7g4�迱�
a|���w���13h��Ұ��'"�iuy���"�"�C�4�Z��Jh��+��nko��1���[ ��f��z��ށ����%a���۝�(k2������tИ�8�p���wEy�S��ߙ_|ɣ��;�_�"���K9��~>j� �G���,�[�q���nz��3g�TUzO��K��`�h@�)����[�G{��N��?�+G����vx;����[�Y7Pk�Jʫ�e���Ĵ���LNm�s4*�y'��`8WRd׽�}P=w��#���D�Oe"�G�#[�i]�]��f2j�o�.x���'re�0.e�'�`��:X~7d�r�|��no���,��=��kd��!����0m�w�79��d�&�wJ��x�-]�8��2h����n�W�6��V�t���AL�s��Z��c���I�v"�Q:H�h��
o���E
2���L�$e�q��Yi�V�_���s�n�ȷ���P�+EO俧��RFL��|��^� h�}�Ȕ|V&L+�J��B�NVд�yz�U-�G��|!�%��{��q�	�O>R�R��j�I��C-Z���r_�B�͐�?�߯���g�8����Vp�}� P�����Q��'�p�B�IW����4��f(�q�[[&.��v��C�b����v�S�?�>��/O���4�d`���9�01�/���j�E��"譡�Wt����P�! �~�7�DzF.�p�7>��#����}=��eMQB������q�.j���V�У�u�J#A�,�����&j9�[�ۖl.m�<O�:{�	���>���p���eo�g�8�l��ۼ�Ћ#����Rr׌���FbzP���-s�0�i������9ֶ�޴.��5)Q��E��j�C`ތ��G'4��0�� �zs���5TŒ!A�z	U�^M^�8jz���W�#��4�5�R�sAQ�
�9Ɔ���Ph4�L��>�c���x�ӛ�ܓ���[s< \,�D�U�5�72
�lնC1�\z�4��n%����]UP�3����=�g#��y�1%���_��v��	���wo���W�2\�������k�	�ɷ넳��a��zr�3e\��LY�E�n|R�|�p��n��vxX1ό[��	���Ɉ=&��LF��g��G=?{oo.�!���\>�:2b(d�駯)x���&�����q��WItd�XK;1Aqn������s4Q��gUD$��f�8���:�e�!�* 2H���|ܒI�d:�/�'.X��C�)��� ������K��1?Ю��-�r�V�+�'}h���	������G�<��E!�Eޏ���cü��ֽd%:>e�)b�@��7	 xFKq���j"�Q��jT���*ِf*�~�v֐xp&�B{*tj��\A���l�Y'OM~��)�y�hA�Քy��KIc帀�+x���h���1��̎��_����A�;��{+>F� ;��������Y�`Z��_���.�v�m�t/�E�@��Lo4K@W[])x��'�~{��W�*[tO��@b�H�\ͭ!$�ΓK��y���,%�Є-4Z�7�-�b?����e�%��厥��N���󷏕 ��1�-��@;��AU�EV�-c��d�楟g+��)�M�j��n6���->׊Mc<��/�m��y��k���'	-��y%l�����z-�Ql�Ml�l���D��OG���[�AQ<Sڭ���x��\�kZm9��d���A��I����]�wQ�C�kO�:\��/�,0��4^oK�ߺk���z���|�����;����b�VH�3m����"p��D[�q8��g��K�s�v�O�e 8�0]��?u���j,��sp�;�x��+2U���-��Et�ck��|�も���۶��%KG�<�ŋ���L�؆��D��4��h���
��[��� ���߃��L�
E��b�^�X���k=IH��ۄ� ��(d(+��Fh�:~��!
����z�����Z!5�3a ���rY^��ѩy���/�^��$C9%h�P�ms]�%�A�/�R�
��z�Ār�4uI�č�t�����͞� �K×�Vk�6���zL5�{sP#R{�&K��������ʫ�m��',�)U��D،��ϧ�c�>�7#i��T"��F-���5�Eۡ\7��KV��v,l�喨�iE�<���N��7�?��>�8�#i�X� 䯁��g��p4�A�)�s��cEj�|��:�̵�Cf�!R��H�<��[��x���2u����U_�gdڕk��vJ���ⷞ-b��+,�ǊZ�A��x������i6t4ƼxA���Bn:�.D`�tX��1R���K���\�����~s��=�-E�_�N�.5��qNO�_���&�\[]@=!��?;�F7+����T���n/���Mto��z�B���Ȓ��EW+�-��$%m�`D$��^R9���|"+�Hl��w�ka���Œ�����8���e4�Y��=�x_/���&f��hb���;{�(�����?9h����H�^^:76���_[h�,�qRF�������16�r��6��^6V�E�)o�`=�j�V��6jg�*�1BӁQ�?Xy�n����;�:�O��]@y�Y���jo:%3�P�q��y�62_p����t��_]v��L�D՟�<o-���imUPi��=�y��W,��f�^0�'��h#4ؚ�3���=�>v1jE7���dFhԼ��!�2Nw��!B�v��&��aL�fE���+3�Q�;e��^v���'A�x��V�S��\��j<�C�ԥ�I�<g���m��bYotg7S�[�64�{#��R���t���K����>�E�/��2�d�2�;����ڌ�����L�=r�HU'=~KF�<t	�帮in��+or$u��N=��o���za��-���k��N?�~�n�b��(.r�7��4W�~��	�d;�.��{(օ����,(>��ˉ�-(��q��r�o���n9�`��o2���Ww�+�f��(x�sߔ��k�IW,�o�Ȃ[��Bdo=Y=�e��M��.ޒ�z�����c�ak3QN^g���vϜ^?��%HƊ�J��U����e�gz�֤�-ꊒ<JG���S.���F>�z��ዜK���QgR�xw���H�.Zl��S�N���M�<���LX�IV����t7d)����F83/�ז��I??@�=d�(s�& ��6�e�|��B<ު!u��8o֡&���E���!5���;��ET6�v&a��
���oT����F�yf!�N�&���'w���T)�� �h���Y�}�iԎG�d���ݷ`p/����+/��!�e�>e��9��9k!���C-����� ��DI�^�p	
�완���%'	Mht��*���(~�'�fp���m�)����ig*�*�y3z�W�(��q^�c�Z[6o��s�!��`dŜ���O�����v{�|�R�=#���G�	%�8�C�x=P����B�q��}P�U�ˀ�c^������T��.Υ!yX4�Y��i-8�G�;6�zz����*:��@Kp��}}�ZYp���~a�*%X>���2ZǾ>�!SgK��U~b-�*�Z&��Q�q��q5��E7#�)��d\��k3���]3�_��%�R� ���/�\lyJ�E�HN0�#���g����Ο�`&��X����#�;%�g��3��k�7�&*a��s�؂����grR�ʴT5�:������D�鸃sl��o��(��<�� ���@A7�,534�M�Ʈ/�7�\����B('�Xr��X}�	d��w�������k`��[J�	�]* $_����j�V�Ij��c��]��r����k�j�;p��׬0J�D엔}���ҏ��CAQ4�~o�g��I5eڱ�!����P�Z��b#= V���Ŕ駶�@���Я��Nd��og�T��i���� �/��<^h;Kl����ZA���Gc1�h[p���Y�dV7_�����1Q�^�}�O�Eu�BS/Z��ߓ�3N{�l��WJ��s��-F����\�b-��*$���P��)�1�퉴o��v&��[#u�#��v[Ɉ_xV?�u��⇿
P��Q��&��o QZ岇؄2�^	L]�-�*�IV�T�X�K�P~z1U'��Y��[��+����|RU�zH�tԺQ�')�}��1��0�����(N�m�om,�4��	�}�#.�\p��8���ݜ�ڽ(5C�RZ�0f��Gi��"Y�$�(��C�iU]��b�G���ss��𧊪	*�p�LC�y����$���Ş�k�O`�UM�,���x��(�$|E}�q��Z��RmY�w�;*f�ON�-y��	�$���ˑtǮ�%����/l�/�-���r�>��G[�wc�N��N�[�I!dS���wљ9+X�{��zq0�p�%����Q�$�?ɲxS0B���͈�Zq�S�/f�Y�Uxܕ���  �ş�n6��r��d�����D�1i�x����x��1����N_�
y=����h��V".��@��]/C(���w���tNڔd٫$�K���}�zo�>��W�
��n[��*�YX<|��}����unC�b�Z�p��>L
&�p�2��*�Kq>�"�I$��	?B?bE�WS�,^f��F���*A@t1n�qM��P����m�VA׌�4.p!�R���H�Wf�jC����rS
�>ԓM�ʪ����xoP�,�sO�;�x�s��ژ�f��{�T����H�[wgiu锘?w��'Ū
��@q�]F+C3�/*$z�q�b�勓�Pcvdr;���vV�arP��92�
~N�*XP�T,_u����e&ew@;�xKb�]�4ѣ���Q�y���|�𼹶�� �(������)f�ߥ&�b�b�|$դ�������Xպ�҉~/ꬱ͙i�z#�!c6�k����?y{�s<�AP�"}�g�!���`�3V��~4L�0?;�Ǳ�=�$B�u�5s�u��au1T�O��;�������t�w�N�!Zx[ES�4:|�{��骇A���n����i�*�..9�N�N���$Io�����Rv���7��F����&X��|Bw#;�h�
�m74Τ�U��ˈ�j&�rU�p���g��uJj�}N��}hi� �rYE��^�|&"�����}����^E`�q��U\�6�f���gѐ��&�7R�L:��<�"�*�8s� <#�қV�*�3�Y"��l�P���W�)���j�:v���.^5���ʩ���2�{.����0D�[�?��֊��M������)oI�vT�ru��釀�\f�ԛK���頑��܍D��5E,8���rX�gߨ�*�`��4�LW܋�WBȨɵ��t2Z�Jod����K������;x�v_'�� 0�pn!�ƭ�NHpL���0�^4���w���1ҙ�L���=��C��%ڇ!�چ����Ƌ?o}k�n���`_�p����`��tȆ� ���d^ ��������t|Y�K���%�ߑ�[3�QG�*�]�x���[.2�IP�r�]O��;Ä1w���a� ���-o���$��}&�Q`-�JU�2�0H���G|6:|J����I7��l����щѹ�n��zL.�#�k�3N_)�bM���>��$��T�~�F{��Ӑ������ƦKW�c�٤p³���흴�"ޥ�̠R��a���J�n���.g�#Ƒ�@tci�J2�b��~'��f��"���T�BČN�����PP"ᑂ�)��a��n�����w����|d`�T��� �f�?��z�dV�؂H"�����΋I�t�=c*��9��ui��bC�U�,T��V���8���:#�S��I����m���Kem��Ӟ���Gk����Pƺ�Y���m��V��t�M-��)�⯟Q�dBa�(�������d7��`S��rhY'��������5�� p�ϼ.A�0���?i@��S�F�hz埈�����?�'�V0� vˆJH��AI��oa�����b@&7�L�D�b�1���n�l.�S�P�XknH6���Ӡ��I#̒��$�q�B�ֆ������_C ����}��V�+F�$&��h�q�o�ݣ��N���&ȡ���<�@�{m��@�0��d���PDa������END�������p��/򙄠[[gx꬜��hW����N<�X�A,�M�o��&���P�����VD�r=�lV���#���A>?o5��:�D��jV�Y羖!+���b���֟��CrB��W�Y�°��];K~�s��5>%��x��u�������WI�M�>��̈́❟���K�;�� z��l��f�E�8÷T�_T4.�U��[|��SSR�����@��R��0e�I o��ڬ�E�@�%N&�����0[ w������0!Ԙ�/�@���Y�M��Ű��׶��� �&��xh���Mu}�^��a�f���I��m���u[���?/y�,H1
�2)��,�8Mw��Y̮+�5�,�o��)���c85ͥ��B�ԃi'�#!��	;``����B��;��G��z # �fL*���R��L�
Jཤ��\i R�#�nA�R�iUT}�̹��P�!��VG]S�T�x-�,��J�MIqJ�ǵ�L���Њ���8,q��6f�ȇ~E��q3'ݭ@�2
�i
�:��b@�����W^&1c�x�F��iW���1�o	��T4���乹�|�ܤ�EJ�-�N@g�����a����E��%B���� ��&$U�V�#�}qyOr����e*��?��;=�b�2v��	/�+��4V����I�˛V�Ԓ�f�I��^����:�d�+M�Y�+���MD倊���Â1H(I���W��O
n�}=I��HV�a(�Y�h��,L&H��Cq��.��(�e�ջĥe�ǮwV��o�k*}�E�"�l>o�J�T�:o�XC�/H�@k��.�	7���El������qݠ� �Yr߯�"�����=<���/���}%����(��η GYk��ܲd��]�ދ��; Bi;�z�Y��ǵX��xu���*�>���TV'����v�r���z�r?E����<������'C;}�H
�!���+
׫7Ӷ)���?�3)Hq�XȐC������?���̍��u�誂y�h����q������/���	�$����_�V��r_5�%y�S��E�9\����en�y���݅.g�z0�c)1�G��u�@�D�
"0��J�L���cz(@��Y��#x�A���`���L
���u�B殉���$�є��8�<�/�S�'�xBZ(�r�Re���{�����ShP('���m�'��-�̰_{hf���',+4R�Wi~ ��P�V��b��Jj:3�2'��aW�m��$�ب;V�pV��F����=s9ryx�$͆q���^�{R �L�_Q�ݦzͧ�r��"��4��
H�8��}�櫯������i��Z)�l��`f��a��n��g�F�:��ޭ�:����0����=B˯��E���x�2Ē0��	�W��iO0$8B���b��l�^����l�bz˚����n4`prf���g�"MsJ2������r�֨�I#������F��ߊ�pG>���ۊ�h)�D���^!7Y��{+�Pm��O5K�d۴MgƎ����D..�W�Y%20��0|���`}.+�Rb9
�y���!����w\�3��bt��VwK�OU��'3���`�\=�K�������X??>!���k������%�5ݺ���P�`��>'�Vª�ڟ���C�a#d�+���(��� 2و�js3=�ȫ���]S-��xu���=��Ii��;�>h+uhnz6\�+|�ڋs�9�K��~�N�
�JʙC�Ҥ�hk�]���]����7ճ]F!/*�;��FӞ~~xVU�ō�1U����j|�|w}p�B�w��W��$���-��,l<j��#�D�w���;������?�Ə�,0m1�X&�r0�7k�V����:y��V�t��?J�ª�����C3_�7��>N�%�f/nSo�p����X�zu��)�2���iC>1�Pv����`�7�7I�ji���nQ�`��˓~5I�%��1ǋZar���+x��;��gy�P�����a�Ű����+����Mjs�8"��vG5 @��u��
i�RE��
��iשXե�B�#���D��?��)�j�i>�/[�Ute���ͱD��+�=˛�J�?������?�4�s�d!�$�"V�a�\M7��|nb������vmq�={��({]�w�W	)�c�e#iw�vt����[��Cf>Y�T��9�\�������6
}N0~�g$f������+����P���j�KX{�'��纘8��*�.��M,���D��T�������g0�H��-殒�k[m�6�,�+�7J��t%�jra��I�\��1�pզ�k��[:0���;�4H��S�H���yl"�PD%�	�V���|}��C0�e?�aOqi� �cn�Ԩ�u��ט�s��#��´h��6�����!Q ���^jr["&��[��^W����35
F�,��S��辉1P,K%��k���:8���$�+�%��7^�b��V>6bq�k �ƴ�~��5Y9���?ؒ=�W�}��Y-�U"�w%�:�R�RK�iG(=��TpqX���'��Q.�Ӱ�F:�l�d�9�_#g��,�{��WWo�_ �m)�pM4>�>�p�$@����,�ꜿ1qK(9=m��F!b5p��?�[#�X��5v���o���XZv_�t�[sِ�҇�!��=�Ѹ��,WC�I�f?8���� W�ƥ�[�/�-ɚD�W��x9�jY���t�CmA��#�PsW��IZ�%!��Ci)���薔
�s��f��nv!�,Da��ꌭ���C,�]����R�x|��K;�.�����r���`\5@����O0��âH,@G;L�jγvm>%�9�ֻ�/K�D|��4Z���T���p}%�.<x�3��v�I�%��=�y�<�M�2 \kL�����J�\��t�7"�tp=GM%�W�c����Q�J�J\��3��
�FDؗ�������
�w�I�b֝�Ѝ�n�52;�ʞ�?�_�Lx�ZT'90Z�������e�T���
	Χ^����n�b%MKNP�]�X^�&N 2La8�T�\͑��^?f�sQ4{M�BVᅯ��٩���hc�3�v������~2�FR��)�����J�*���	�����S7�:������M�$ h���9f�,���B9v�>o�hC�
lr�6.jp_U�)8�@W>��Oy�R��Rni��Z���@�� �������~��
���s��Q�fk̫N�嫫��fR����I��@�������BH%��esJ܌"��al
�&�/R��BbI�)�m�d�4.�m�1ָ��O�m�%�v{�4��]��ohhsQx�v��e:��cSV���>D�,.0�S����ǭ��d��'u�;)�]���-cEOr�.`�)���}0�7-/�#�f�)�0ޚ4������G��ں"X����fq����8��G���C�F�h�{$�[��:�J~�*u�υKV�;=�d|�b�I}�:�|W�,fzЫ�����hدD��h(�n�Z����(%��c�Z����T�#�2xR!vDE����<&gk4sQ�N+!#��S�Ĩ��k��0 TIͱ��u��P*2�K�f%�J�h�GX��|��e\�vi��-)�i���O��~o�3q[��a���	5i7'����O���0ѡ������&����/�F1�|$4���ӆ.�fє<I�����m���uZp�t�%q�ǀ�r�� Kw��k�߇ɢ\c�'N8���_%:,�h��tm=��2��˪ǈ)�P׃O�b�3KQ ��B�����L9�0������'�]��F;��R :��%�Έ��z�?*�ݬ�E���X�M��Ҵ,��'���|t#��֛L�_Z�<2ޥC�;��������=h�+��b�5����t���ܔP Gwځ�r��d��g	[*�?zH6�?K&������9赣��!��oN^Ѷ���}��-�Q���;d��cXB�h�n�c��`m��9m��B��s�?�O��@>�cN�Lh��獧X�tw;m�ܴ�ګ�C���/
���n�\�6bI���C��A�	�ޯ򑻟�{��x�i�c��UX9\�� ���ھ�$�[7�%�����R�]S�r/���o;E�qy�
�:� |S�<%s&�oW(b<y�뾎w�������OD^���'��P�_ 5tP��cB>b��l˘�ԕ�'���lbn �������@3˜���w,o��t���t�ﵳ��C���T>>��DqȚ��~��Z
���I��E�j�R��<�[�O�s��=oL���*O�MZ9=�1x5YB(�fj��=-�ϴ���K�~��:��f��:�����s�[�����σ��d�R>B�Y��J��~��������=�M"C17�ŮM�q=�C�1y��n�߀������Ы�(������T>��8���BlGu9Ñ稔��ڃE`����j�K���ACO���3<� ZFuw��w8��Wʵ�����I�}~r�\Q䲀(h������5잞AK]s"6z���&I!~���6' 7[�7��!���0�� T�P$�o����1��j��{_���b��~h����Um��A�6��5[0\w(�<���$�p$�chp��L-�R�9��J|rL�|���-�F�s�}�ݕB8m�x�^���tO�bn�W$T���ٶ��&�P i��%6�>,�4��(s�f����e\ԝ����j�b_D��F������Gs����m*�?��Ib����A�i>&�4N�=5�;|s;���K�L�D�����x�e��cD8�5�d4�xɗުu�(�5Lr����~�+��as������|����W��)4��z �~�	�M j� |+7�4N\qm�����1G�����t�Gz|�����ey
��FK4�ܡ��xu4��9B(�k#�Ş�����wR��"������^~��6�#m�c)�ٛP ��+5$�� $$QIC�z��*^t��AW�"~'Z��ħ��&c1mag�	�F=d`�k�7O�k)�l"nXs�do�\�.r�߷p?��������2@;�(�נ�ܔ��oc|L��`4'�g!���a;� 	�r��&��'�â�k�0L33'I��9�7V���0яAdv�a�\�g�3��N��`E� /����V���g���/�� J�y�����sY.�<�وU�;��0�J���ƍO����0H�~�d
��������pퟟڝ�ɓg�<�IO�:���nP_���t�0l}�9�DhZu`�[#����1�����{�3ſ�Ï!T�p��q8k�h��LC����c�aB]"[YT�A!���f#f=���4SB����l90�L��V�<�C��b� �que��(�5^�a��'<�F���q��x6�ʢ$27�����F��X�(8�o�rU�0ۤo� O���dSW�zdġٰ89��N҅���,P%NO����@��F8�v4��@�3h@4&fmyn7��Sך:����_36C��`�ו-��ţ���FS^ʸm
�D=C�.5Vo��[n�2T�%�g���g�����/�E��k��R��o�$�.�A(���Hr���)�1��Ǭ䙬qu%����M��'�RQ��.�+�}V8ׯ%L��膠��o����2�Ͱ�Q��W6���Ku��mO�Ӭ�L���W9��u$A٪S�34Pp�����^7�ص&��
���/�	4��a�K�*�c�ƿ�]J������^3�z���!!�L�r�p O�w8}�M�>��\�Pz���x�b��n������nPA�����Th�����*�+��u�(�ݙ���`�
lLWL21*Q"q�OP��&�����`������6��iG<��/������ H;Db��~�g�?�tg��:wS7-N�_W&��k$4����A=��^U���U�Eho�X�>�A�$�0�J
���MK&W�����]�/�[X!�^��qbm�Z�;�?D�W|ag���Q��ݻ�w�IT#�����'�M��0RK� ��