-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eKo6WsVKosS69HnBQG9qKUimwEuCgetliV25nwnC3lPToYUVpWW0LmtAl6y468yOnQEZIiewhjaH
CPBjJgDfGysDHKaNQUTw0hvpwwCh5e/ir39RfW1fPmByY7ztDoUxS+ohJqoayW45MmsIQhYFnARI
MbMZhCaLzchJD7XOdH7rs52uvJ0/i8i+sf1NAjQsizrmza4v4Med+VkIzXKuTNlP7Z+SPGxFkZuA
ty0nOoixIxVDynx2uFDAMvXgoxfUUwGp5IvjBIw3CeEtpC++rrkdwLOSUV5Z8d7G75F5atLZNTkG
S1HpeJU4Jiqf9a9Ol8T9SeRkz/qN499WI5as3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
RMuiWrVsElA/r/GOpcTEQfJr0AWOJwSxXNbRGMNgFh/yFgdasvAXPl+k/SFFOlr0E87O2HrWD8sc
BLacn24h6NwZGsKvKFe+oDlD5L7UPiE8sLXe+DVXayqJL7EKN1/B0xs2nR9mNerNzeRmAxBwq9o4
m7U6fcgilSDejAzdolzMuyJ0Lf5xx2CIe2+IVxPtRBJIU9yA1XdZA7TQuxd2Omf+SXsnTBaHSqrg
1LFF7NeDwRj9duxwMXcKadYqqChTiYPW56KEmNyjsOWN/cIW7wk8V2ui8N0o78S86QisYHvj/5TA
qpU+RY8FqMdo7vzrin66AuwYmTTf39sZ5tq0l0MqGqltF9Ik0HLnrKlFUM91SvHWFkpPo8+zVWM3
Zz9m9BrUImXpJ7uRMNGou4HnJAhrKdvevqcvMXk4RVXsd4+mSWYrDhGUsthf670dL84KVp1oJYHs
f4KteN8DgPCkN6LFQ9UAlacrEITaxtpicTUGsIcf+2DMA/sU95IfkkYd+IFeOmktadsVG3Kk1pVb
NY4GXdGfSj/DbvdlPqXAzFqYX8L1socGUTszTNH7TuY0dU0dQ51OdRRofOFrC1NOOWCZmAgyeDDc
87tu5loQMNQsInhINvRKSTjO3rpWTKeGDR4MjOsHI0d/OlUmjD8EVT9fNotltJwcKmh0uwp8kfEE
yhMQtjk34FsuZcCaWbtEik3xZhzQlrL5VJiNCCBBt6HGTHmh6z4RZLctwLNT7jIFbN83zt+MjKQR
Xgo6e02tpmUcyroESoDtqcx7++6RC/HYfmoRbc8SDlxVcGPv6LiYn4CdLuyZKoa5qtxzjJr/xazV
wnu3zcmk+BVuZc/x1GZlvIbvAHTqnKiPZ1KW2tIVuaGwKfvCfn63DvxI89GdCDFZ0OeIWRHCh7VA
DZ21d36YAExoY8Op3pCZ9fX01u870pF3oYrEYqX91cxQjn7qOsvZ/kTIvvmvBYFikZ2OhmCBRBnz
ddAi/fXR2QfRfEcHaxD5QHZUaiV5fgNfkNIwT8N7NGJuzJi2N/sxpcafCqZ3rwpA0hAayFcGIBjx
yEFXvLjVl88QwhC8vcK7aJv9oG0cAuD0qYw2HQKlQ6AH1iC8bTwSI7DrYgtCsj9PgEBeunbb76tG
Tiw3AtzOGXCkEooV65J9VyHw6U8LNq7geIEpO1D/wULfy1Js7NCANYUMhVtpwM+m6+Pf74dZNm0C
zvso7ZdCO1bVnum110gWQ+Md/UlsxzuMFYlOjiXkWc2AbHRS7/R6X4B0FjAZ+KSS/r+4WBfnCZcm
iq8mg0L39Aej2zxOUQBPp2YyYmpsIhkVVXW4UTvB0n93EGV49AgSe3cau/ZLPyOJ3kIV9hQ/zDvP
yr4aSzN/u6l3xa901euMWxqV7bsu+Rv5RhrbtPLD5ADBgKeSsXWZ2oRR/BI+B7dYF5+ipUoaooqc
9W7Zp6EksHinCxDsv9fVBKcj21OfhucDoMBVXAPjdaMck3KNO0ocQE0VQV8vyx1ADdgp8yJaAbzN
nliVisAqUvJsH4Yn4Sxv1YWf9ucAR4sZuaaKpkRBZ8I7PiGM+GMv+zjlp/dr/7tZTHmWuu108NeT
5oU5Ssgp7f8KRAtW1sgmUfMGx8953MivgyeAo9YU6S+bnyLzYv3Sm7HWTC6rcuzmTJUIh2NArgZY
ayLvxFSiYIzNCl7mapMZsg2aWcKI5R3wz+cPb8c4UFSEAq2r4o/vb33iA5sR/twckGCwCjcsjMW4
MWEPPj9nS73tb1946vfEXfhWuCxCfr5+zyr+m95hG4j8iNDsL0MH+RQNZgkeaTelvhyA74eawQai
/cFZPV4HbXsReXljcFb31wBY1MMeEhfXHUON2K5/PfcriUk+UKLLrAiOrtaX81eu9B8kcBrAES0K
9kQg0OBYDG4P5l5WqKub2IFWvERk1zXH+H8iAALtckDgUYrMC1fmlNJBlnyqF1DAk46fLgfD9ezh
CqQ9jRjjbzemhiwM8mPdXyv9Ue7Xt7RXWMjtrq5RRVKfbEksRVLISUuT3ZNuDJT3lFQftibUAkLR
d0zogsaLB/aSWy+Oo7glUwYuReYbMNRR9a/yrGusJDIdfXlfb7NTgisSgvuKLajuemexnnQoKE/t
ri5mpGE8RA+yeIvEgL+z9FIRyNNdgKgP4tmSUGS8IhB6iGjEujAwHW51fO31LtcrupqeLA0iG0LZ
hlVXP1HOpzYidWX1e/qXiR2sDpA3WlOU510hj3qVdj2dZhOm6AGcDfM1vzqgumZpHo7Y6Lf0KTqN
8B8/HLE5oMMzXkof1n947w1aWdNOsiE0cU2WUA1bKjk8o9x5x1nGh4kSpjMEx/5JHPmymwpI9Bhv
R30XggxXL5VzJQDcHcZfJAb7dMKJuOvdyAxlCQpcl7o10LInWIGBohwlt6CcBxiQ4MJCxLWqiAgt
ttFFcA/6Pbvo/vGkIxzNW/MjyPl/O0+nGo8giGO+GnmwhaGOoL+zrlD8cym8IJPpjJVRlVafQ+dD
GBNEMDoRY2L4xxpFO1SkZeNUsQY9vbvb61SBgSwsyzFtM/Fe4Xl1Fee7rltZQPJ0i5YHuuujuJ3A
YWuBvMSQwkMVoUGwgXXyUYucgM1EcM8Y9iLwsFFLsE1uCTWFbfiwe7HKRYtdrf5W6qd90cnSRTWr
SDVO1wQovY/zKw5RWyfE1XVLxalli2NrfAQL1ArEFMX8qBLsixJ5X4PpoeUusQNM2IP/3a1unTuy
cUH2Cuk+fhswILV6yMFR2sKr/2Fok/7B0WUV/Lx9/Y2kTWTOpyXPZmOvpNolpQq7StgTRdAcVu6g
w+yPv0wCeU+vUW+lFK2TEe048TyoxzINZqudQ/zp3LU/SHqRao/5dWrGPujWYzX0QSPAo/cbfwrY
nR8pCkgCA+qlzyGbI4Y2A9W333zQ3JmtDyRvZeYPWuGHotGZz4qu00bcQSta3dA3FIRZni4uiyzC
0Rp3i8riFiIyrXFw7iuIzRwoHpeMcKlMcD0d9Io5zrMfyADS+3hS/EU3Nya38VK06IjXbX4gGCHf
lcontSJ3tO+ynAP59o3rw+3fn1Q4skpfRa64AvDPX0HOGkFPM3qkq7tIAJ8GjZTxK5GgJ+OQSwft
wqyf1WHZ+DQOdV+BHb38sZagGkF22A/IPnCuFT/QDAT0KCXkH7l8TKUo+p6c/DLQU8HwY/MiIWFu
tjVAD7Z2EY5gh9Cu/xZeaHtPiKoWSQ5itIqY7gr1VaprsbwmW4+5SXw3mWWYm78QcXLatB7ub0FN
ptRSz3ti9mPSKA0Nv9H39vGHnhEZxLdGtYbP9gPPgH32rsFO3qsyYtD5d4fmnqBwrVmDxoitEEg/
6UJolcgiWOVDfTX++JHnKofs2GwCo/XvCFjmbk7FIvnf5BCWQl3pfEdYnAHYR/V7YSyc03F3T1tB
qN6bLWAhhor3dnchc0RKPl+dpUPBiFXwpFhf+pB86Qu/R4ycER8JoHkIb3lEdIOSgpa/Dm59MCzI
CM2FEvHDDdpLFX36EtOH67L/yt6ju3E/yrg8AIVwAj5uJFmwtGc1J/ahPqyejuZMXayII1PDZ8gB
9m0KVUd7B3WWCaOWhcFikghe3vheTs+VvGMDf7oeU4LmB8cOix8ko7k4S20f4+5DvkTK7UqysZwP
olhIbuXR/R2AdQ3CoS2NLDOq2GCbOEufBMiUuUUeH5Gobtdv45e/MQC+nLtnMB0ivGAXmdU2Vbc3
wOXTcb5RDpMqLAHFthvLXc8GG7m4npyX9KSVVakwwDqLWg0sqlkUg5nLMVXakminVFmA+6qaMWOh
NlViXX5Lb7gVFVsYIY5LhAADB+Iy1LnocjSnv4ISUQd2G7qzVLjmk85+KonHk4htpZ011Yr9/Xv+
XX66vPEf0/hhDL738J0CIG1UxRvpih2Re/qk3wFlJoOfWuE9a4enXS43ogN1j/Mhu9y7/dmoOyWR
2KkKy4avHAyX4USXxdKWJTmj/JznLVN2NaxNyTcBlnNnwJNViuoP/Dpm5kAYElexe+LAGxDKCkgh
YLsomyc8Dad7afFFJW5olX1ZEDSjoKBVbE4ZwSdp13C/uhWXFnrl7T5q6dRP+HDNF7jzLSgwL02O
hXu0jDoeUYNBd9ZUVzUcBOkgYtBRJK6mG4S0h8iLlT07w9zBcGb2wpNxgyb3HXUdC3Q6azFuxVJy
xy8xVgEJphGvH6dvT2LD2eg5BL6zLuDiCJ2mexL27RiyC+G/O7bSkWeLMSc74tzYrVIboStf1Bmj
Zu59qTWPtKBXQT7C3+o6fR2aXcE+qK46zSRNwFJmVJyPvdD7BZVAgirWwkeYYNXQFEFWqEE9UWZ4
GLxKBYqSayEr2HaRoWnaBlUc5KyXAlIsV9gvj97GCfehc2AOFElTQyKb3mUS5dZ0F3PHWeXkUUVY
FDuCjCwY9KrGLDonA9pVep4m1eTRyTjDetbeRYakJUFawTua3k5vkUuO9hyl2vmXfgYNniU3F0wH
DjoCupzq/W9aNpHE67fhzo50QAoPtGrPGubOH+2WUphPcPixyZO5EcJ8IHnpJ+y2VDhKI9FFxQms
jrImw1czeRn9iPdlQwWq+dH4ubltiryIAnuYMTyMQxaFmnDteDWviARwJJRxAK1WXTvNtnFP9gSN
sflSPhO0FdkrHE6IzAA1Bwjfq7McVwb2jYvm2Sbd2dg+AEdTnRqxIJ1d1d2ckfjai6D2tmK1MLPU
dENgEEYeFIuxtGINdD6sl8gIGv/pOYFHLXWK9aJ0Ws1kpfxHVnnlNbOKr6KxFkBgMpaeGSmBEMHu
3Ahcj5W2sa+U5GKNcGGMG0Iu0Jb+gVa29JuGAFyjU7Z94tPKRpL8Qg7OSiqplNa/rIyG2XChbnYV
fDCg4jIKoAAYTPKgPQ0dZhoyW6QjtzpQoEIfSKazZ41QwODpvrfoOuz6wcH2aE2KEE9HlBYtk5tQ
qoXfZr9kflsehxbWEweMYsaJFeMlohNDMSStYPYJ8djEDOPeGFP6jJUH36Gkznoqi6hKOWOZOOp/
Co3Bzqb3ateQ+SucMhMfnTXq2TtJPrbQJXSclEQWXbtQI5StpzLFWcJPtwU+t+7lwwx++ze2HfPo
gTH2oIPtk7ELCoqvAjlJnuuX4YjeqGhun6WvbH14HoeD++aE5Lkwx+lDnkvM780yI+GMf5Yr5gKa
r9ueGx5by6hly7iMQn1CBempLS3Rl/qyy2BfX6NyiskFATyB7pBkChNDSAFNJrL5BZvKcHiejMc1
pe+oCfmUf817upDBqdkfrQKHwASGfJAmE/rKnCfnr+hJX7k1XJbwbHpgCm5McdOs7ZX8cDlXv/6K
a7EbGB3rSy2Y9hIjCjJkknVz/eztCcibPekfekIAy6vHowpazfOdYFMQerI5CfAV2YDV72K1K8nu
R43paSL+p3r4TRX/I2pPYicDmiqnMbLGnxUGQGk+HzgXLg56qWZCeyVi3RCxLXVRekcPF3Maoo5N
68SS0KEl5DooxHIOssST5WpEvnNMrucyQCpu8vFLPKshU3Ie1b4nagEs8M0n5ziprhis7sCqNOl0
RESEVOuguIamW7853J6t3k2ptAsYB8iuOQZlay/yLdRe7jjM7LrHBY2zitfJQ7hntCJsmiEm/ima
MCAtm4dXlx0mocjGYb6+tjL/pfUwK+DtVXtfUE6Oh5Ff7sToDIPvB12NwFtMr7GyfDchjUZrFVuW
XwGzX9m9PdZhz0BLEomq+Qm3WTIEUu46shc432SqYBF7kFJ9bYSdRrSAqRXuFJInuiWdWL/XCRKG
YakAWup9tbA7gdv8dy5qAQTyUtKzmOR+RCn/riGO/Ls+59OXRTKP+Xq3Jq94SfMlj9PqLSqg9WY7
qPBBPN3fzeJFiRV7w0W1d5Ppu9DGwS811oIqXqTMSgYka2SMjhFV1xAA3tgQwranlRFSfELMb6CA
1nYQG7PXmgrmXbHXPO2buU36G9+aK67pdhtOs4FMCHAnt7HyybdoBwFJBD+NJwDkI2DH79IkwrWV
Tpdl/bPHtzblknNaWMTbWPKfFasVsyhqPkr8rvZJEu6aCy603xn6EivNHrxVus9WGfxMhs77jEwF
RXoVlh07BVk+tKqkmbtRPdbikmaMLryER+N3w9Ny5G1ZJ06fkPJkreNtDwdDmIZ9XR5ujZ1bZpwf
qsxxRH0HZghIVqks6Qmqck/O5BlFEFLawwVX9+irYyuItWfxJO2R/vUsvFKf/JgIqKV4UlwHXSVN
j34ri0F97b3HFWouActtSha9c7qIU5R3g1a6wojiP7cOavfrrvfhp9DIbUTvfQTeIyTg+oCkhVcm
sF6SF8fWprMudkNWMx6iHsubu/ZaC0McvuIOdzUA2reWyvpEdzngnlAHj6zkrb5h/Y7jZnTdgefn
xyJ2jNUg6n8JiRw4P3AP9lYx0bo4kZEmiCP9ALNGwxneZOPON7SSpMyn2GYr+BiF7qOgmLG/tpXl
U5dqUoFbods+oDj9jGt1MP31fnH93TYkWumuK7/raY3EjEuD/remUpbSZQHPyBz0TLdhE4iiA26U
UOOcjw6ZAxt0jdt0yx+CYQ3y2/FeQd1P8M5BSYK3fzU43DJkpAxYjNULXNoyH0yyl66smUACtGul
dtnuhxrriaXETQy60aHqpZXDZ8uoqlfqQycOPW437u0r2quOYCcngjelzZOVfz6hIKRS3DYNrPus
3PcoK79ChtF1pnCRGp9BvZTS+1kbkcFKOKYc4fRrr1MRcO0z3xeVNfmdoqJH1ze3azGGsnOzV/7x
OYidt+nEn+7m+Dm5tC/DOXQ7W02cc4mOKuBF5J0l6ymx1srtpCNmrXU32XInInEF6CJUEQbHNlGC
M9uBuyWfZoa17/URbRttZe1yBu09TIKBPH8WKYNsGSZ4d/C/Jfx59t5/oVMmj0Sdi7SuWw/I9nkO
eiuEC0kqjWiE+0cig0h3ueOoqhyJrJOm3Hz4aAdu35x/TXm8M7vhMvcZJXql+QgAh1m38Oor4Y3G
kBbbcEdaQ1vWbnJvP8SdRZLJmPWyGqVALMqqnv1hcaXyrtf8Xw24hMl4yP1forRUnQBS+26k3MGH
raqba5timSESE037mbU+GDqFRfGXujKGXU62l7V15lzzBloEl09afx+nJ9gcmz5a/IMYyC0laCul
7AkPAwbxClmPcuw/hgHLV9nHVY7Ya38skYmsFONuHkNeY5D3VYNX0qbywWkTwQ960+hxraQgtkG1
yM1NjqwxJxUEQIvxuEeU0HO/Sogynyq1HLia4cvOChbYOqll2qYpWtDbMwphJeIMipDMmVphBD/S
ivddCa765uJ/kxB1NDuzR8sQsB1M3w5+uD2FmD0zFZmplClWUThuMASZu5q8pIi/aCndi8eiY69p
dys46d9mWJvWHRljW41VMUJ/bdxmWXuRXgFGe3ibVxSDOqZ9keQmQqFigCV0QQR+gDMR+6Pot4kV
q19H2sdeFLfEDbuhkxOmHwAQ/nVWH9rvdH3yrDHilSdX+p1FBilvWHiFfyrTNHAU0VHYsK7dgJcj
tGcaYqFsGdchkLSS8Ifcyn9X3pzxWL1kpxEtFaajrtKnelWd33rSB4A21FGuZIAe+tQskv5iyZbP
UJZbUUt8FzvtOIzgb+pkhYJlekNaZEYBwWqV33GgyoVUigEP4i1xmgiP9YE6i9Grfy7aDFky9/mT
Hl7dx2MZRENSK2h+OC7H7mupnWQz/a5KOA7+oZl1faQOpg3bOsFGjmfreAwJc2xDshmy6z0Fb2rv
bNljDi+B8/ambsqXJ7xMb6iSYWhnxnJTTCYm1kxqkm6+9Kpecmbnjja3tM577NAsVUF1SniL5Vnh
ZqxZr9Atbd/cqO3/IS4P/A/3gla+qr3Vm16PxhdekLVg56Mo1odvveR58QBCguMaHxQTA+sujBjh
NKeNKRUQBfiVEhyb9oh3R7PgU+SKRcZHmGg0XcPW9UPDQkR7+3BQGzbG5paRGHolHq6P6zAROVUj
dqnKskxSe0yCKRU7G2rRLyLdV1vEUyJVwpZhiTl4B20U6CyvVfG0PoIx/HM4vr/58C9LG4hKd/OX
2UHlRHDis042XzePkKeHIpFnlffdDqMJIlj5jyE9uM2pMl/do9JvF9IPfuxqUlRhN0eBYDp4QPt9
2WF3j+FMal3tDK6b//QCD+o+XaXck0wiQg4HkDg1iIe9st0fAv2XZsBuopFHjpZZv0mUYZv3RFrE
bpA5HrK0Rce9ihllMG7UHa9xoPU9Ld8teHARiMwb/NTTN6OLPtU5IMZf5zVjS0fsAbMd6liXMhth
lNDzuss9t8Ctcya29Z1oAYx7bcVLN+pmeCOLa47Daja+iSpyVsBTtvdNozWaIUgNf1m2SbT2hdk3
bWhNLXfepYWO4vcGuBLnXYzZ5EP9L53XIOnPXLYDJGU0G2az65d593WW8kWCR6eZwClhOdeMwYp3
JtCxI4L1ZUxJILhpQVPEluAgbaOM7M9rUYKen0oGs8f5+ncAeJiomAoiECdx1O3JQITWns5tc9e2
+7FaUfyWf2Ev4bs/Zi52xgGSq3SAWrmzYl9EJbAp7pk5w3URlYUtRZofiUEx4JqInJYxBBZSK2zG
eL3m/YDYwJAxPGZz6Au+u6rj8ZLpTz50lQl0jSJFqEd/q/fvORDmCzR21UesrB2z51VnKgH0D5K9
fKJ4D44zP3J/QZvHkHajV1ZXhtAHwdp0y5AOAwnWuzctmnos87ESV1iq9hR/52Z+JVhQeWwri0o/
tOM+yPX3EJXmLoF6LYv/Pflj0ky/4GYObGhUr5VDPV511J1055TYOWPbFwDJaAJV6in40yBxo4Yq
2UTYFH3cQxqXm/0dW8q59f3nbtykdvUSY8hxLVh4RK8sYOUwn1qgKqylaoiTAJwWer680P0UeHlK
dgWdd7ZYEMFzcvUPpDM77QK8cLn64haGx/eSRhMae4II825rhSiacT/jcbD+OLS4LO7r2FkZQpIU
4yKdiP2Wvyl7CnPwZvthKjMQgmlZPzNy2ivh2RDGlKS8LUfx+Iwf1T+HPTjTpCtwMs9oMZRTfPTf
myddBVpuPKrzkQsJpeV0bQ2Z4UqgzsNZ4/ofutdzVSlmDyOPcM5NH4WXKcsLrURReue8IPfGOnpp
zPW9lhHNEURvWXIWtj/TM02R8BXsylAk8UPYvQUWf4/xAcFoQ3AqFZIGYh5UlPUOzb3+reIOyJmF
YXjxe25D5RrSdOaoBvXM9Lt4RoR+zLZPoUQigIMrWHIUJFGtbLEabiNoCwCuma0Z2eSK+LpjTOuA
0jHpaca5qvPc+B9j+v5XRthzU/3WYZXc1FaFaU1UhXfR+2pe56LBTBBP//VrK4CQziOm283TWU60
UXdUs0wkRdkD5wc7ux2MXxtl2LmEjsBj8L5ZHq+kaY9lUV/RO8/kYGSA3z9XgvgPDx0RWkmGCeZH
xArPyBHjZoRGCHJXjpmfesu4nfEzKygAPPAUPerezm8JxevoUpEXC2gpFjepT1spfWZcPcz7O+xE
WxX/BPpL85z3MiD/oFf3VYYuH/9ctJNKMclSHwuaLdV6fJOCibICf+/e3LPsi3ibSfGULRaw76dS
WPwlM4hrJQHOT89idJR7AzUKaTxd1WU8X4ryUEMwbCTFHV2L5+1VynNXtqpq9m6M3R8TzFFuJZ05
pZPCBq63BlkiKxx5CWSMsYxK0gJ6dTWCzsbnQMX9jjtMF0Fo1yZNhmzZmBCjlOROG7m+PGEO+doA
rNwxAuUp4HpbFtGx6ZO17dn6nUBBzPGY/wZBTqirF/2sIJdX3trjsDJyO6v4ybh5IFHeEFGm/CcB
TrkYG4rh9ZA/sZbQUB/vox+EFeRWdZlR2DVM0ZyQYXKB59kIddkwBmhdX3QlI8+8WbO4/S0uGcHt
i5KOr0vy+v/V1KVQHI8qDUyjhAbEp5Z4ArugpCqnMhjI9enGhnye2bRnzcMWR6eUaWD72Ik2Vny3
kjbeCvl+X5OiBBPaiUhYiKoqOjqQI2fiKHFumJcFld762RTobnmIk6t0hGOGe0MApX90Ky0ZDYh1
oHqjxfT+w4OZniXy54DG2GnDNGjh2e/NhYLUjGLjHn5Y5Yq11p2Vl6iZpjF2DRpG4505m1kfUYgd
1TPZOHfuVOc779r03SqiOZAQ6umDLoaRA4WjRMjpL/S49eAGwr4RaqKP0T/UI85lfDi2qjIXLraH
zl0Pk7ejLI0E/fbNLLk/VakHQmWT1hgZVYdhx63HOoaYOA+O+GH43DfYD1No5JE/oMKSbbn3DzRr
OHUUqervTKNi4HRw2hcZJDAGD0dFfY+la8iPq6c17Qtc5R6xaOHwNajjOvJf+1pd7nn95fF4JvvC
0gMtk8YEgBElA4EP4zXoAThZetVBZmVj3T6NKMtvMzHeBJgewncOOYy2yHihLJHtnqPuhHvjfLx8
go2PSugLe6oeWFZp1qe2i6K3C56KAv1ivwOmIrrxnxlLkvq3cTEt8li197FttYuwcAhp4JaU+FMW
7VhK4i8GuBsU+pBueSLGVd5DmWklJPvw3LX2yUt6hWuy98tTqEcWvWRi1KuF6q8lvNGbOvrtHdcW
2qHF0/0ObuNkhJeS/95b1DyTVR1n6bu/glgHdOQqux4bkfltdtxZllb10gRM8JsxEsuXsFyf30Bm
RkXKM3cK0AT4SI6vNUQnp4uNuYodXdVKJjcMINkwwGHpGhwq/eH93DhCBuOmm4EYIyzdtZlYYqF8
JVuxkY9CeTD420O6omsMvaPHRbU3neqYtNZSLLFkJyNUeGP1iGYsJFBPNc+0zvuADimLewA3neuy
YQitE+RAG4mNaLckkgtXyhPTvPx5k1SXNFga4dxC8n65okZEkTXLm8zyZbRxVAXXF6LiZxDnOwkS
oikyM9X2D/tIrmFL81RhSeUo/yB/NFJ4YrSBi8xT6jpnJ9B4hz1yWey6xSNq2pbGx5pc9C76r76z
izn3zIoPwTbYVvIocMj7Jo6crl4XlZ469IiYN31g+DBlCwiIg2TBManSG3wzIr/qdgEytTn9vwii
yF7aTsyriMF8uSTpISb6YGIKVHqIYma0l3uPDayZ5nsSW2pOscL3JzHN9l1aRMOfsT6vBEN0hPy9
9Bo7XqQ/mJRTXUSgoSJT/CgKaxENHoiSvdnPZ1KFCSH5Po5uFQSLT5Km9Ufm9GG010Jty6CqksMI
uc2WIpOSuD6CwNGB+uktceWQhQRvOgT/uBA9Zz8GM+8CjeUQUYIwefNZVQeB+AhDXOcswBRQP63N
VCz2dHxaZgUbI6qBqdC0eZ2xS9hM2r6MP4rUNdZJXzx+HiKCMf5mAAek80jmg0mf5P1/vk9gwAFQ
3DRfqH1EloMTJA01A4AQmFUXcVR+7+yWzEE4DXn3n6h8Fd7OmYJ4DbAQUzveJxhSddT+O3HysQ9+
otb0LPezAaHO9AW5HfnCpCVZg1j7x+/Jmc9RWgpdYRxHzOwZ4Dk4kwYs8QZoJSGpAIXMKa5zv5J3
PHM/4n7/TMHWi6wk/hZWV4v7BaDr156BKsez2/+Cca8D+adhS3nbS7Z6FjtkHMKgz3DIiizfTP/4
Hl/5Bj1sy+bpKjrlR7nAhjxG2NbIyYxjM6lR2BeUrJXBVWNc/EDrDR9UYTH6RU/B2VlEbr6vJhHs
ZjOt1a31NNIv2E7skEVlVOON/1hk82D5Qq2MJGbgROIdmr7i3Nn714EtQ63yRowWG8W0CfR/U7Z4
H8nTqrz9F18jLeTeROohijJ1ZnGmXdxDOEVzj1cVFiysq73QBnROwALvgQ+1vv1vA9JA+VGRGsPE
4BPwAvYMQR5HatSunphbcIuXUteeLoEIJ7rjBIJim6qY7tqzCLVfcbNAsB476l4QQNI3O1xwlKGU
3ItO2DMkCpGnORnYhWj+1bXH+1wcTFfWfxrzp66i11f/nJXVA2rGeZsirEg8fdY8F9v9lhL4nlWy
p4G1GHaW/YPTMQEFJAxSd6u7GlN4C6tTaIGsBx8e2tGSevaBZLW6cPhjte43tXr9Vi++OXgXQ0ks
55AUE+F2jQEBpkEFt7dIYux1fgGr8vvm4Q9DgcdXgcNlsldHu0F+h0PjlqNX/ldlGVyj6AcQpMGk
Ph4XMNp6+agnpyGARI8HMJZJ0F82GRhm57usJ+/Sn/zi5Yl8IxbyseH9/Hahp3JGhKUVhlJTalkD
yJOb4NQvd9WVxznd7uQ0zBqZYVt3fRJ66rwf2tYv6zHildkyc4NwIUB/mMJnXWGzzlZw1Nq8mVgh
R9M6vvuDj/f1Y5GvIw2lIeJesimCH8goGnM3bW+OA6mNqVTwqULU25Iqsg2wXJV32JFwTgHlv78n
bsz/yb4poi3SRcdqE8YdgAJdTE+Sb+X/Zw1wD/9m4kYDmredd73BpR8sgRPddkT1ZrPzrlyGCR0a
RezL7vakhFGSi0VtYh8W64airCScPam5UA+uAVfLODgURc3fhfHZ+q+Sw8NV5ySH+UhAFXpcK0Fv
mLH+UWo0x9Z5HG6c4sLlfdjlMfdAVwlCdoW4+9Sh7G3jwW2MJL00TFX9stmVuDkSUI4Em7rHhxXF
ZS68AoZ3k7UlfCpJSIW+MNKPbdMuYUHyd/C9Vrj4YT7RkOF80PqAJen9wJm1VVD/UXdmZg6QZ0D1
PVnmtwdJnIl+qPRbA2+wblNv7tpY3Ak6xSBgj60/KReqDt7DEgUnW91JAbkNMhh2vXw2cG7+qVI4
QzZjYBuvRBaFujPU05SDM40NYbTo8yOTpmEg0tauB/LaEiZ0Alj3mdZjRbMkfxSl210FBjv5gP3O
jdgjk3+FEH598QeMOMht+iH6kTOYiALIZ54PRcLiMx7d0+jjUJ2kqvSF3hRGzXBtuoDXWHn3oNY2
v7C7wzrOyFL4xQau/LFApTSmVLymWDz/JtwIUSoz02CLcMdsF2eLerbn8WWJ/zuZuB78flzog7Uk
uT+iKaLxw1N3D2BDZGMndlkq82X0/IBDYDBBUJb85HCYtc5xvI6doqV/CgPvNDa0eOetJ1GPAjh8
py4fLeZ0x5hdIAxfACjfzhpE8ILsC55siszHvOIww756LW7APzeyXQaNBrpZbO/wNYmaGYXvVjpe
73dEFhU1LD0CTydwmruxP1GE8eL26Zib8I6nMhO0fJHMo+aAMJfHRPUOho22lHXX8LFnaWxpzYVV
8S4WlgHjQpbb+vO2lHFi5DEeZ5VkGhM5xEzEob3rho+vjXKWgr41DWuuhBY3U+DBhxnKN8vAQnyD
9Htn2hAzKkQEk1cJpI8w/7OA7xQAEe7NyM9KVLsd2gW79JTaokKhwVGv7Ne8AQa9kK+y9Gck80d2
iUaZ6mtxQd/kRBOsv/7tCsPaeZk6Z+Ck8vE8x/tArPs2ERXz3Z/hQWPF8hhGYmRZ14TLDIgNieGs
+JyHwIVtOPaXD/AfIS3TUzTLiWKFhbgX+vrMxMJZ3T6bonnyiwEsaXVUiYmAvTOAeh3INKAolgSt
MeLCtxou/TVTIKGac8hrQ3YZjwDNSVcPGBZ98gjBC0QdZlVGmYa+CbNEU/ztKDS69Pn1FhQ7NkMJ
SOcruZYi599TMl4Wb9R20kxZSCQ07eLwtXeQ1502ekbFvUSDZSqt+6aFHvsZSdphgbs3Dft8TIyt
evHS1qKeFzZja9FtZz8+XmdKrJO1i/cCFVFrtrTUYo45JcEjVg+i3U8X+ZafvJzBqBj4NhZ23lCN
l1SX16VYc67YeXikBjh3b8/3ANAM0u0LOddzP1h3y9jDhElhsOk++ryjb3xkacktlXB7uq8+wHoS
bJgXhOyc0c63ximPVO3sNWfRhl9ou0AQogaQOESYgKWoHUheGg8+UU5I54QAaurpdtmKKTkczExs
ikN5SaLoDfGTKBdUGAQBJKok8XhnWjq7XBNAfDLvMor5Cl/R/AiJPVdjx9SNqnDegiAkoeRBoFHd
1jA6my2DFXgTkO5nmr4fv70IyckLPWnzgQAE2CpxHAdXRi9LXHGW5VLEDWiJcDTs01owU3ZbIrHz
64wlJADgiGe1HUOYJwUZby9uj5SAH8n2m5Ubli1eerABZuJutZViO8AWJIJwAm3h87tVhL0Whq0T
aU8Z1Yky/vPM4zmCOFym67+4nwqkzokKaBi0U/N2rq7t1QWnchH1vJoXeDWRZV0sHb2c2/KONLmE
ZNe8PwiSEOqpT9P/YoHFWjszS3bXKCqsy5chUQ5xrD8pv4BnNIkl9IFHSaL7BS7qDqYMxRaJpKIh
REAFttTU39xV9m+nADoRM/X8QxGDqlqkganZNEN814i3/Xgzc/K1E6khhVE+Jg9fbEUYfxzIwjSC
6TaxKk1ErGqwtRb/FqfwFx0LUFi8OlFsgsfHjAJb8YET1KyFyYO5JYwi3+irdLmfs4rp4DvR/X2+
Pg/jSZbimDHxaAo6fxTlvJlwJrxVxvFgNOE2BMvppLE121BKSnUd++Y1mSwOiWhMQLW5eXb+N+gq
2JRIwYyFcIeFzE0lHluiLvZv1gX4/NruNhxYlGvs8SUAc3eXfrwoe0lD1jsaBFQzXNn5GaxLcSc0
kJTinxs0/EAbrH0r5ArS3b9voxlnE8hsx6IGUz4b9WlkrRm1UwFa/K3nuLLA6+G+kX6Q0CcPLpSb
ReuA+zpX79CZQhAI1tpo0e9heDwjql0SQ06lNE8HEjWCtdjya3p3vUTgzmeT5lR2GLxHcKpuPBgw
y7DDypiHhilY573JDNyE/0LCc7+L976YdTdT1Cii040A9lIPOm2eSw+0Ii0JTvlDjp6MEwnAya0J
nWczUXs1tQUS3KPDnTI16JJJnABlANHSW53KVBNcf/6Py4639UNbOLqjFS1/6lFdoSvjci3gygIz
IFPRfcmXSG0HBxCoF4yzubbJ1PcSOehc6ShZqiJ84+gyhBk6ApfHi0In8mkDqFg50hxTehVSNSqL
EOGWCLbQp5Kku0VQ9/FCwdMVj+cRkE5V5559bPktGXnDMdnw242L8gQTxWJBK1eOXofWMv8yDMir
UNma2pL1gAViEVC9vAeBmnP2Xd7C+rsdLV8ZvByR/FGsueJEh7RnJDdNhmW5bB6Du8ikf4PHCfbZ
SOssNgS4rZJhiWKcaQj0Xjvt1WT5OlhDdx2/pHLYqzxRhMBzkouqDD/wx16JCTNUOjbybEwUkub9
lhHaZlKm6woGuw9FEiyhWpfNCyTP26gfpHamz4VSLswrP7tu+8Bt6qHEEzWlWYQBukqeQ0gjVlRI
VIYzBpKdIZRA/TGNOZA6FbyIaXFQV9JfyFBhhI7MKmXiJkOynOYe2zUXnAJQLC6VeAqe4cYNlr4N
X5ZT5s64FxhK+Pm05QWnoNJJcJP03S3wYlNK6sRkAe+0iSjCnhAV5dkXvcs//I/Bv/FeYxyqlWgt
/yuZDoKVGVSCiK4OlxDDqE41Z6eyPomCkoooidVNs50RZkKpFrFy/P648u+0h0/3J2JFNQ3EQe4i
e8a80P7HIOx9/UHa/jH/o3i1nKJ296QwMLnvTQa7DgRfOZpy6rnaXpVtTY59iVQZdCW6Ckf1npOm
VTgYpljKqsfUUAxio7wd51c1zB9Bud+mSEh9BOi/LZDvrrH/ofWNhSJ5Z70YKm8N25RkErd2HKyg
+LeyAPg6KNLyNcEzuQL/x9Q7QaUtgCHIFuflokrReJqpZcW2Du091dQPF7rbbLp+gb0qwjZuU04N
B2pkYLTK/gTbxrfrewr4pUYsDNcsz5aX0L045v70WMmo2i1m4W+OUSnobMbjyG0f1KYIsxpYoTAM
A/K4j6YOpomtxiwv91AVIn9Vf2R1ymly15+vwmmXKcfAclKw1wdQg6D+diANZjBWf6YrIOzDORzE
Tsvq1C8NCNyxa1mEKt8tDHiQMhNNt7WDQQ43ALfoy0Sz+7jNPhcvJNRh4b88J6umFJsw8nn1pMSL
y5p02TA9GhlT9yH9EGpA43m0I8fOYR80IEKxj51iiiBfIK+7uiNHMUq+KR244dzq9/ZbfxzXSyKO
r7T+64UTjQ1oBRRonPPcNBUPHNFib2Ye1abhMPAT63LDfFKAsKo7wGjDpKGzjPHk6e4q5M+Siwk+
RpUiyabS4pWqN1k+6pcu/rZmwgH43LH8qWwM64huSMqwpxUOihG2jtD/OmEnDjJczJKX4TFvovI6
xnkhsBiQUxqaxO6/S1WokUHOOT4Bv6r1V2ENl4vw8xKNQpAGKVYjKL9LQKweYUeuS0xcvR8qFf+Q
1pv3v0+zMP4om8X+Eh94OA0dzSQ/SsH5g86s/4jgV1cRIlmRSqyd9WwCcVbyvCnv/RT+tDP+P7JF
rykf+83Xg/BrDkJ1zyNAO5ssZztU3L7I7HAtb30qbSd845boUrhNd9brLukCbdutuOUr4XZ/NK6U
mfZo+zwT7G9V5cTe/oxRZ3W1/9bF83UsbssWA3sP/jD9tTzgiD5Y0wcUHiGaBQULTpqwhipbzuyX
rivasWh22F8PcG+Crv7FPyDatRA/PnPS9sysSY9G9v0w7c5lm2pmlOYbzZFFbyCS0PN971aBNE8M
DsPeB0UY/SflgjvtR59TQbOhgyUbjFhyhkUToNtWyQRRq/PaS0SHT6wcLuPzhBiSmJ8XuwK3SRLm
cB6YG9+ztf+PSElCJGusxM4rRFW0+pXq7mxqM03sR7BX7Kay69WETmJ7GTOUfw7cACyaOyxAwAvp
j7PTcb54UbVKgX3x5QHrJGE0DV+Q7uHVK9k4g+UXVCp3K3CAOjkhz5csrJmSOXPRzY6CdWmERnZ9
bkATMxEklwriTExrkrG+E/s90hOfIB4UQFruVRLL3LWZcmd/ZK/hCfzBL1aId0HmMexq58S0VpQ0
QuzLanJb6uiqft/WN/DKct0TQTRIUarcdo1f02O5tlEOwDCChqmZnq9THGHnj+BRaEwGx7yCx03d
wBjD94mQtcjd9D0wVWUv9m3ANlx6yvPbJAszJmY0J19hr/zfjdzua0OXtsVjbkO9UsBBVjhibli2
EyYeWrPk4GmOILYFQLcJ50954a9mwwUR0GnwU3rI7AIzJyy0tn9T9rxuSqjCuO5chfP4FU39wxh0
JwFxGbnr8HEvSZNj3gTsq6TkI6XVQ8jqtt6t7rtrr64B5fSxtEUqVJecGwWa3lTuNCtYOZx/Lgt+
N7PB9QNWmo14DjebDzsqBJW3EnQN/slc9rlmDn0UZqog1fu+gxA48Ev0UIXAnfUVaI8qtdbk7ToY
ZZzdf9iJupf8hcJk8Gmj7yoZaijjr6wIi4aSRe6yz7BRt9o33Zwir2YEbd/w4cpfLLCeuGbARdYX
N94Y4TG36EojuyfPy1c6EdY7tW/csoQsKrnahqhGoNVrL7kq/t9IiRbnORD2s4jlQBRRI5HoW6If
Py4sZU0m4VJjHRzi7otBzOcFfVJ64VlC4vuoeykgECkWEry4TnriLJzQAjR8aJt8iXVLWo1hm6hk
rSbdF6laJ69kguHqHexoq8NY71KXcPDn9JMvKv1nVoP539VJFWTX+y4n73sCirMMdfPehiq3mtpr
3BLtZiyP6I7vQjwZyQJdwQtd4hvWoPGg/8Pe3bDrcSYJRiA3y0ZLpYwvXTHgdyz72ImlGN71z3QN
bkIYHYxKDf3OFedi3wgeNU1b0a2Kf8ge/nhy/v6/+I3n2tFEY6YxgRa0Llacaec7xnEYoJUekBmz
b/D1HVESlKQRp99TVWg7O5ydVWr9OequNxNLvtDJvP8ac32MEkDxzEzVqeKG/v+h7NgjA92ojR1K
h4wr0Aod7XXUj56mI4l2Xve/eKEQLjiJ3yd6OlzmdkJZvIJFv+jGM6Hvz5Zj3aG3dH1LCnBSyuA5
F0pDUsw2OM5xxnReEHfM5pKCPfNpHHLdie7wZKuR0S7aioIo5ghASQO4gy5unIlLChwsFTbCIo4U
W7CZAqSNS6wb/cgOPnOqlVsA206ez3PaMpOW2Q4hyCaDyrA5jJo80kipVZTS1MwgRR5PQq21Ohbc
ua654M9cc8gxLJXjbRyZRny1x3MCg/1FS951xa43Hp8tx4ObrDU93chReOTdyFXX80LkNzPR5PIO
RFha4wDijLzxtFE82XpZC/CB3uvrdkWCYd2e67Q1y2wGFYucJxnB4RuZhRFPnLHjLisx14Lt5h78
dL/K51EbQS6p62rk9Vn/nOyNG2IoaNinAPAh0TaxndENbOI+1QW8O2n9AZgql3wFl8IR6jvqWAZz
/3JHJla7mBjG3o8sNZUT2Z9pploPBnz2SwsK2mbtOLEZW5IVaRFGivkze/aD7zdm2wXlil24iEC2
Sm+CHgIBwd6Af09R1DHtyNrpWnSJ8JPY9oxEsMbVZKQ/BkoYijKx000vSxbIyPFRbgROmr2JO/2z
X/fJH/BkaBi9f4bfgnipoOF27qcHzj6e1fBn+2ZP5is3ySnmvTrO7cRfQpWfTISlwByYveivJbjx
UHzmG+YtyAOGRBumjSeQl7N+aUduoI4KOJQz0QsIIDDBjVADK0FhfXouF5ZLJcPopURucVQ/Unp7
+s6STp0qrtbfLPK13+NpkJQvd82PAAexVlmZ4ljmO6/qBG2QD7yLYVw+Bmggg9a7Vdzobk+ZWQSx
sOfkNbeef7kyuemoqZsgD3h14YSjUehF6Iy3Yhwlfki1y9iHLOCJSm1fQFcdt6MwQWNlheJ2krei
+fMwsq94cMJYrqwApUuBZyt3JP0IfbHBDOs4e7Ox0h1vkNx39YAFxFCTF8fpDrFy1VxcXmZ1hyzJ
ZaS0Swtp7lfeYcp3cFeF589pZgLm7kt8o4ViVmdvOwALyG0tYEhSYsTySnmtqUvb3X33yeS8qt57
P/m3W1WZepxC+zP4WU3SAgIhpLI84yN4iQdCT00TEMxZ/4LrHXPCsKKTkHeUtlGictewXeFugun7
y5i94mc0Fd03dFGqjzq9vGH02CYPz9dlzMCpIcqCrUqo3d0/6lxzgEwOkIkTC+G50y0NsdN20Rf9
3mR9aOMQz+IkLY8u8fYI+nRiPtv2ifyCBPipflPCznTFpvwzNuUiqvXqw+EsssYDQEt52E12VmDa
R0NWWdKB9pYipVsgZ94Z/2J2CU0pGvFqFd4viF34hGaKo8q91kuI+LUfj9DO2qEsDFrfzm/433Dl
ADu/QIMkzwOH9AkrPXOqBkrOI7SAsXw59wf0y0ux0mbf4wISBIzMbiRBfY8fmnWdPDn1wA9NEFkI
UaUaXS9Zdsq395n7JEkW9iCaCA781Fmk7TnQj/mdoazn97fA0SvUHQ22pnN8+uCD3vtN9M3WyDbP
p4eQOZTLCWjxXEK8cZbjXQgzXBefXBQTWbuNZFgShU3S3tfUauzziFiJFWOSv32t74yL2wOY5Ind
wVb2DhEE3qU2rZUHqfchQbmjgmdhcef+xAprKvcYb7Wgb6fHi6GAeTp5bBrBr0VsHVfApV7sOkrF
3xjIA3GSlJvI0e1j4jP1ftTMy2F4j26G61f+7M6uyLVV7ijEObHpRcUk+LQW+Wd1D+4q3iLDSnSv
57h/rjpJFbN0QzdFgWq7K55gW9xQlUUcfo2P1Ve2RVs54410BqRbWerhtKRwj56lZCUj2WYLvw71
N+GpIFF7v0bBJgL+SbVzL9QvpGndrNrL5Pkts0nulouI+ws5Oe/ieN+0GEa/qIJueCn9AZhl73c7
ZoH3kHrY1n3pkZzGN1bGan8Ax5YmYwcyIMeTJE38/AfVdIS99E1KYvOs4zZnk0GNqib9RGKiFNc4
ia1p+XzxVTCwW5wiFAsVNAjYRoeVasrsyr22pi/uzx4NRzbVEoc70/1KHRMa4ge3NZCLKJp9TMlT
scD3FOHUYWGiQ1RDXaOkFbZS47shwCj7XR52PizwRJox/dzqWPXC253m6qusWDzJa4VuUnzAdR4M
QeAxRZOjjmBD4MxjpYNCHi8PGDWOiq2DNXm0qt4S8Otfl5N5akxVk4v1XODe/Dav/zDFLTAIuGct
V9H4haSdhNzfQq2NepbvwMNBYdZwQVk99d11BRYrSXkv07ekccLhmovb+PLTc1AIDfspN6pRF3kf
GrZBxvue3XaWoVWgfKFQGgiig7gGJzfolo/SUHh1aByUCL8j6RpSDfr9VtM1b5jAERVuzs4Z6yeT
drizWZQCpXHabxG6MApy6iLhJhd7FtjgMiY7lgq7ErL+oq6Rn2foGe4ICbsY1VVDdc4TbcfgG75w
WmD+fcdIdfZt9uLC0E9OU+szo/1GmhKtJ6RKQRaEYHy+ex560H1HGq13FcZpHRGIQOL8lnaoLfXO
AQkdv7HJhV02uve1ZrmyO7lJ1kCwE4rMLfobytZymQB54rOcv3TH1v02/EyF+hkenqdtg3LHRMTn
4PYhFwVz5hm9/mFYBIAFch5KURGZFoBNpPP2IxPviCSwZebWCb3niQXPZAYxhWjxAn9Go8fUAsq9
sfWa6rojjeQg6K/jPlLfaOxAT+yENY2ARkUD7HI07Eia9fA7RbeytA1SOaa1s1YSAfUfYA6v5j4y
Qgp8eC4GUmjLCeFV7mLHHyyoOjQh8QEHh7nTazMDo/Bd/zNAi7Mlrpn13cnoamxntpecRcssOflh
P7+bijCx1whS/08vrWpTgO3qybJCYPew9oenskrOWbsjj73pm9whxG5sSIZGXiFRzWUHChkXKO0s
5ZQCj0Ib9txfrL8nMNX3+66yXnbXhykJ9xZFYpigEaFPtoel6g9Ct65RRUqnrR3BvJsSO+8/+4AK
laff6e+Zs1ScuU+28n+urcg3qgxmZfhaKH1k08UDmHajy+kdsciG19HzZv3aTU+DBP1JW0JRA6pc
9eZQqA8Ze9UuklA2fJ65/TXb47FXqKaFLJUlKFlXPEpC+qQp5SykDA+aaL3hpxNVG6Gcc9+HiZns
Q5LBHaL9uYIRHXLUXyxPXju3yeZ6wpuGSPQShMMdjfyzieyshajSqbzA2QamFKQOvpW7OVXw9Tb4
QhcFpcpnSk4i9BBBnnVCUwnOVxG7oKkaZiFMT/17D4tFQ1P+Qs+kXrAR+rAQxx5KAWwvVD7x2UXk
8vErQ3lHJytGW9gIQHBcmeN+hZMcGLsW6cQiS74FKQWNYqy5vvCpyssFygpReniIiNfCzDAYA4o9
4b9nWNoK12D8vE0JrCd7ia7dNsu0CHGCHixeuiEMYwgcviaY56HIzphbB3MxSQ8puKzTU11N5V8j
7+40ne+kLz3FKd04fHLWBxo9GDNsRn1eX57MMMMnQzO2uLPso7brTXkvqWHZlIDglL93ysWr81pK
GcVhUY1DHKNpyyvF1Zqdh2b+reLgaW4PIbH9r6+aiSlaAJZ/qq7C1OG2x2KOWkhEnTq9KjNPFwWa
uefa2ixr70IjpKCqcBAt8ZgLOn5pbzURgiW/C6WgBvTJArjEQq5yBOWz3stN8DlZCT92oZUcgP/g
LkPAccdKFW4EXlArAkoyZq9Y410KMtSQwbGdIhS+IV/JB9JoKbJtcPhStkfO5gdp5H7WEPC0jqsu
CFcxtYj+VG7FkFcqPgHLzifLUsWdw1P/2YILpL7NN62rb6y9n9uk3fy/MUbXp2lWN8ec0BrbSgh3
RZSYroFUZeQ7prBFUZqyV+4/13H32jZGcxczFaoRWgoWaqIH6VFucGn7EcF+CQhwO6Y4klxMASz+
AAt73+bRs6uRDQpDKxAsMMFRapDQzN7iusCgbAnxGTenW0vsJlaQICwYhYQrT8oNr65+YfKlf0f9
d32s8iDBfUucNmtTGiRoA6Y+Yepsu811XTwEqwOgSDdtjpqboOInlrDWMGYuaYrKVNtcXLg+gTM4
+/sJUidmXARVBBv1T0uOXI8XHwEhJE18Qb1xLi0C8Q3zkRcsjkE06X58UBX7DGaem9Uwu6HEfN1u
HxkGeCjqRoT0FagzAxOx61ggNrqBmRVQ0z+rCTsE9YA8NLCg0z+gAI4/WwkgYLy1mj+odWVWWSUp
9phWczdO5AeOTfVN6FYzZL/4qCG9C1C5YyVv73lDu8qOwmxMnqFLexzdqKO21jrUMzfc6F7IVvUC
pdAfD3CeZvjVinRp3rfBs1OShr0Q8WhsgkM5hNfT5If0iYvBEhcx0A3FoJ7z74Qyqy4n/E7FCZZw
gff9FqL8QNdOvHypsUoyRLFPyTyIpJrBWbU7iqfyDXX//d+yq2ensodtxIGqFuk46+t/elrCCBOG
XKzpBJgeWbWy3TUNpfRmX398i5ElQd3V7wPf7HyH6AKTGMhog9x7UvkT+8oB9B5wVvar4KZsuOAN
r7DT041iqdHSbAZFn6IINLKY2Hq1lzZhP9RL5fESU4N4xrbC9BR/xLIaEURiiEilLjenUGVaVz9I
rbYWlpOaW5x4CYR8VZ1CdeY4pwNi8EEOGVn3FTGjJT7EA5H4uvqjRFn9uJ1TYUVjjIrm+AvobeMF
CslknHnzerVM6X7DebHPLwvczxUF5XDWQMH2WeuFGVa882GGQxryWWsutHeZHKZo7AjqOGTy3WJV
OT8iAXMnkRhl7A0R/AkF/excWf6lLM4z92kzkHuNrSYdqG8IIDQBTTuzuw9h1ufZ7TJ7bVanPG2p
Kp3YNrv8ERQleJxms4o7z/vdEvoI6h0p3zExxDp4/OcCv7WwOLU2DldSzO8ZvbHw/2ia/21854No
j0/jjV3KlLDmFjzHWlmd0pScOuC47LVijGSXzYLCt0KaLUoxjMgqP2dnge9jO7jXeMfdt5ks6F+8
FAED0vLm35xb3zkuqZ+n+0hv8UPW8UKVwYxzuZtACO5f/BzP6ixLVdcZmat1jxIpVTMlharkomKZ
Xw975HSI7eTo1FXS+AsVOs4Kf21o1KzUp1H7/BudprHkDmenb9hjSqwDJ6SwwtDf1+2blm+uZ7xA
8zq/ui0hDxRMqSle98FJrd5TM+mAvyWM0uajqoGnTTvyMKjb8e3EbcrFo3+hBqUq+qenYXlqdF7V
tl1CcpD+8ekPTWhwUyjSbpjI8yWYaoO5i0Yz0u04TIZRATKklQsbnMn7ooVCEZ5Rh/9KzSih32sP
QiHCoPp3Gelbq5ofaa+1htLzZ4t9WYAysTxoI/kZSjLF7INigPLaG7Y0ySsOzhqLrce2OdXx1cyf
YOv4VECD1fTbgpkf5jF5kIZ/f7XbhngM1ujktuY4B5TACiaYQte4sQT7aFPTd11VYN512sCG6e9K
ViECnyJJqzk8XEHpQNmorXsj3aBxex2G7k5/33yXOIOyFHjCrK8frY136Z5jkXGiC0x8EfYAzdCk
bYuWNf/7PEWV9bykPp274qjSvi4D+DoUteqP8oQgubLBFxV/vfWGgV/E68+8PnCjtsGYpbrTkZSd
wGWruWQYNN4LqTSDJGdmZm0SddGzqf0OW0JFjCQPXGecRNEIHkvXIIz6rzMJoKXhGNMq9PRcjZ9F
zhk39eAm/lfY1b00qJvLiuk5m3cPR6qW1HhTtFVfrHw+MUXnbNkIdzEA6mkaJgtr+A+MEs6aabnV
fMjHul9w5ZQdd3cHeNkY9p9Yt4FxtcGvK5zCMQquuYLldAvNSdCDGe+dsBqV0jknLWV6Bcplkj8L
9FU0bjMqjwtZ3jTQSP/CI04geKDPB5uqzOtFlqePeO6KjrPExvg+0+NMPOHQV5ldi4KtgX7f19aj
dTje4O/irIvuvnklx2fg6HqzG8nXwXVpG+gDpGyCOyK4xMybWAZfxeScqzOuQ2mAmD5yPu54/QTi
kl0MQElA9DWoLe7iSauAkwlaJ5lMv2IqGxQD3NA4DU5rdR3J7sszgE8s1609hORL0ISP8tKfZRea
VoOEd12ATlHMBgg4roXtyor3tmeH97cDqWNF3ZrIlquZ5CTnylcOTIdvamyFk5Z3zJjgLPh4apze
GLLyrS03li96CWq2OMyagLbbPWN88PqwBE4NMzjUcRxJjtI0V9fhnRRRRMTqXQu5r35Faq4XuWTW
NWpLg42JBBanI/3/orHWLabptikhUPbgHKu+gbO6BZKapyqmmdziupcLT6okbabUlBGRlqE7ZyFw
87D3aKcVKeag7pPYdiO1uz/qMF9K0cwQq4+V4fdlneQKNR2jAslKboqK718bhti0dCjtbk+p8J1G
YNYiWrRzw7uTpDVikvEIoQbOKUbUgYMa0NCnJsK01xWfwwvdOoYsZtTC4VDwJhTnO0ev9taLpGMs
Nj68exJglqPId/ddxkHnbgLUiFh1mHaA0/gq7hEHnummcdMYURBmpfuNSt/7IvRKUZ5hYP3ANbbt
b8Bype7EOjaLh/JvNXfITDbI//6g4vK5A6QoNu9rQzFMIlW6PbOLZHvfQDrTVS2jiB51ddqQ/glu
UuTqaUnqJiVlOYUEQvTpU6vK8pdXFvu+y/XSttb5fj/8j5TLKL/OOCSGNCcIUZ5oy8GLU6KN/4uF
eSDdt3e2M5G83uL3MWpHuGwrwmMvHb8C7POdgfJ7Ae/5IiF+/846DiGjNHrVum5v4a3CrZIrLtW5
y9Gmblm9M2Kwf80LuwyBcP+4RuOgxjcwPlTBh9rz1i4cXnnLo8ViAaPtS4ArUW4xOS8ESIu0vE5H
TVltfiEQgCi8osufZwNrlOxXRnimq6RBSyjusBHlgKkO8zXMD/NAMuuiH3dZYTu//IO0Kyzrg7Kb
lnjQRGlaGvWaNF8f8SrgZWXyFf36DgvCNBo9m+IKfSQWJGVpCjuQPelESiCHourcAnJaWBNH1pVc
fOpFVwfOI7cjFpU4OoFS4fslOeItHRDa0zso/pNVB/jQ+Pt9JnD17vq8yIT3LHUIqGRDcZtEH5DZ
6BvOlMGe5bm2tbna+JwQ3dWcp3eLz8PF0NXS3U3xz8KHQnp7daGAQuDY7pQ+7f1DigJ8wuHVHisF
184tTnfYn1QoMBqoXOXbSZANJLR9DMOshBGHsnbnWzEH9GUEKBRbcN02iZn4BKtcmFQUNYiY1tOo
JTg2ad46VUCQo9FGkwU/cN69OHU+oqeiP37JtDksGU3uLQsF/sfOOYnKjGkWS8eqvKNViCHI4aoW
gKZobBZiBorHONXHrzZ0Shry41KPKvclRuOhoSVYLtkuCSvYmvn/u4uBGdARZKMfyKxLGEZe9Uxh
2lXg37XppnsgYjMtH2sVyObPwTUhTAIVSwN2qQ3GDXPwmJ7qpR/5FM/PoFnZD+52C5b3E+iP8RiN
TAtr9QF3LBW7T7KuayM9LXwPLpiAHdEu8xfSVm/oIXOjCI11PtaJ/yrDnex9DQcBphjn7ADHe/Qb
GuGrsK+a1D6LOjUUKan719/O8iC2bf7IGhiYfuYYwU/Cr9d6TMpHrVA0IL/w+BcJN0OfYcD1fPUE
XZcpoN3R0oVZiSlY3qroZ+9AwOAUdKUk+hrfdHVlfkib2Uh4F1if9zqniIH8V0TdHZ300uAG8Srw
vVCxvwf8FalUrl5VJL3gfz3H/cxvs+8aXZI7ADniRzGbWRSrFIDz+eMtrn1mDcRuTqF2J2eVAyLJ
u93wigsCXGpTKY5jCi1YypMHzT10CNth66n169W4OQTtsUyPft8kMq+6r/y87l7GlRjGQfAHz5Jq
lmKVXOLfAAqFOaNXzUnePYaOu/i7XtiYQ1UmEkPiRZsLcvrY5VvkIzzumzNR06QLMlfPwLKFZ49F
YsU9vObH/PNqqpexoZT5tsu9D5hcx/xTSOoy0IoPaRrDP5D3X4rLZ0o+GV+4R71KLDPp1lF9pjuJ
/Qkz/eI7jxnzFFY1OX5qWM+gfD4Eng6Jw2QNEKK0LX+QKzJng7AeccXqmJajg4OVYJZrd5aJmU2X
oSkNT4nHqH32RJkyZB3sSrR1Nsjtj/BorelvlmwKOP9D4zjVXRVp3GMx5vQ2XrHoIEzqPoM7u7vS
qCGcG9D3hH4ZZMITiPxH0KuetEf8WM02S9oak3dybSWVaAhG1yCS+4Ac82MjnOVZXP+zVTVwPX6r
IsuZ1rxWgQ7QQoK8lmzVbQWKyuOPNVC9R4gl+P+GB3CxWgGru0wicwv0Rvj9oUoBNiiohNEKIdhf
zN4L9xFlUFyt1fe5eLpbNS+HyEuWWp0VAR1lrttG/P6FUBmxHdGPmsOUEoqUUwXT/1PZFwqwMMTG
IvaejOtA2NzOpwPkmz3wwPvhvkjUT/1cI4+tGCQIcHyk88fvJIkOKEcAXfuR39F8lecLmMJnPqxL
gFpqSPPL1DpilZoSbbI+bGnqhECUqVWrbomUVPjlNUUJ5A3JZsfu9USyyiP46/g674FO02+oNQ/J
qcPIQJuNg3sGO3NvA/7u/DsN94jCpNP85krSkMTVbaEYJthEiCUcfeux8O2m6sC7n7IQBFcSaCIw
rc8S4hl1X0aHC9ti/MYHGKH7up8UgJrtbTyp6WJAuQpFUo/UKur2RV8W6H8b9xHlF7yCVutcB7JO
sjzscvwetNYIDCRr3FsxUko7SCcYvmFAAsTdGdcijTcTrnaNpqWRF827FnyEUuzylPSXmdxSJWtk
aPfpZQFuxCXtUlQBEhSSCdVWOGxssD9BY5Az5ZUmHTfFOthONYePmy957YlrthiQd/ozSJdZxUMP
E477lR45DiGSR+t3D0089yOu/MiueM40pWIpGrvHtgIfoIOsYjyBr6dGoKK8162ONEfj9HmCSkKr
EJOQskRQP4EBnbfAGWi5Mba0Q+wtewchDusy4xweNX6gaEycjwlrpmatoc8znz634DkviBHyo4i2
0LJ5MRXPZD09W/nygWDwqR4Xgraz15C+6uQyLyTfl5+juvTpZr4hVvoykc/grn2FVNV8GgDSwTtq
LLM3KjBfYa9T6J8+2e6Z9uzpgSelt7DKuYv4kCnzgBM/Q3i/gwZEUBgnH0WJU+i7i9Pb5+PH5s8x
Omu5bngtJF3/nAuRRrqqVz/z4SiB7yFzFPbRyTAp23/C7WzhsTluGrUZcN9n/jCN/nvMQobYqyay
LeMM2LpS+6ZGVrCZjOXrMJ9S9JWO2PI/YaxXFWCGdxYl70Jtp4jpLUfkEclbQrbFpUQHcJgjElpk
Q462RG9nffhcW+4UVuk2azaP9bPEKWj9V+lx9FTxw30yGBlyj1/b4PQLW3NLX6rCPRp62rFS45l8
1C8roQySYqIP44vHLgxXvU3UBYRGssI5jQpNVqm6sgNl9O2Pjv3pWy5Tt+rbIASq2Fn5Ind/LIgo
vIEdmdrgLruHP4sUFPGJvAa67AIqe0xOBZWrE1vQeZbNwYr/Xl1VOh8/zDEavqgomV5hdiyurzoq
2q2/1WehDiU7/11nl9htdOg4OGsPjYoslyBW6R5ovlscOKNSLc7l6phoHT1i0a3nrsotYPGQCMu/
7q8308qxorbbhL7EFycPVdbXfthEEMy8mDGnf/txKRUHwax9yUIY/eS2ZfiPAcSBrDGK1jXFgn9t
RpEiN1yz6gLuzsDswRj+o1Sdt/XnVXQsDiTRrooZBGKPEXtRyybHRm4X/kgfLJKFwYlKtcE4kHfE
OE1XBlQWf2fffZ6HBzbO0eAt0ihSy/4Ww3nrTNz5PQ0CTBooCGw8DjEJ8miDK9cx11dhWD1/eqYd
4BU9ogRSL+RDpN/s1+Mcmn0p8c/9xxqbwO36HPdN2K1PZ5M5V4qvh57CxhmeuBr8BPtn7xXtxyY5
IsXi+7qe78HKGwNOv64zNAhmnlxb04Jh/xQ0HFhi+apQyxyi1SyzSIYUxyNNKzKchvoK6GYG2Opx
RPVwYnRyLVkAMhOWoOkfwo+5/zSy8GvzMIW33JBwWr4sUlq3nEykTnj9mhqwxOjK+vket2wuiCoB
kvTz6CIUx5Pu6yh7XACGmIeTjwDzGr5wteMlbkUHc98AS9y94tvo2DdqcfsQvQQxDa0ELJ/o74vv
zWFcMjQQIwT8q5oDxtvxEXWPlS8zSQn0d9fo0tnCQqlK1ZzvaDpMcA8ADLOiIQAjL63zIfm2i9Og
euFUaoALMViI+LgO+9LLFv6qmgy15FJ4vOaWEHp6CKWp99mApURUzNAh/ohazx0IZg07cuEmfdQi
t5dKmo9mTDHgZ3un/fIdPpENHuVm8ovndIE3lRi86OvEKJx0cy3+oBuSesa307kzxP3Vd04PTAWV
5IAHsvcDiqZbkmKZxOJZ9GFBZloe1fSlJfDDATieUwDqOg490x8XTLPfmqOkZNGS95XrQLGimm59
i8Wh4eATk+Ok6Nw0f7J5/yjzkCphokQ3MeSUQRrq6w1uuudIUKE0Hgxusw8a8qEVFuLy7iaLBRuS
MYtaHjCeZI90MeIjHkhRIQnCYNWU6zlfanZbgT9AMTeYLgGXJ6xEgVTn+TaNnnceapm/EK2l7bUs
uAjfpQMphUH2Liup5eb5Fjuqiv5rjtzTlUkRS52NJTrQsYhtShxiDAkRhNNUFjw8M8+MH8XqEi4V
usTN5WAAd1vSzBU3sIVAvG4XtO+B1+jDYrGFuwrD6V83mtj+C6cURb4lOofRKT4txbRneMA8nwmT
XxuQ9xgNJ8vNqKWCrCCd3A9uHzAN4GqpEnesdXJQ7ZNPRF9Aj0MnJvIRMagb1zEFp8TwdIX3kTkM
T9qmq/ctqNhV+SBUk1Gif9TXwERh4ehIgc1LdiKkhMIpMbq3JSdOZ/+4jm2qh7jpdyIThrM5y7Bx
N0eDCdQ9vPgUqElBDUNr7VZIovcgPi1ZlExjKHdpnwopwgIRZVLShw94vGRMCRR0fcKc00hCSc3O
eLVOM5JqJ7zaZkJNpj/JA54YLqsvYUIcgSPh/KxrcxqLBwRXWzFW5+4il2kaHgN2VNIK2yZxX3hm
4ajJuLHTqMBGkZdOYHQfq+ZBHwZLtgKGs7jnC2JiQQ++F4JCXNWYrr2lVmJiGfBG1VoFDIF3Uql2
zqHSYtp4ex0qL3t500jGjWV9Et5mIucI7OVwvdmfEYovIO22J4pIeYRp5BOn803ZvRgggmcGkKLB
CWiPNG9QKQ9VcvQK6in41UJm8cbS8Oxy7wU6Pap27MwLsI1v1+ncRT4LSVCWQGDPKVO5OBIKTMUX
U0q0ZwoTnPP0dS3eZQm470APlkMrWr2Cye+GGs2kGk9modppmLqCq14u32P1qgrCuai0iIK4Ln9O
8kmxlMflPSh5d4GAvyAeZKhY+V8Y4eRmCY+57nO4FuR1tMLM2Ez0cMlVsXjm5zZuNNOo71dHLDyk
B31AU7sizfi7p99JbqbWWM3xmMG30qDRknDx2LLwlL58CEUQjaQxC9VOgzLJBht87PDOxmaTjLVE
A4y7AE0C1If7aKUlbGPUVFKHWN335YeDoQJYHBA5YKGNp6R0rkGAg3JYV7xzvzaW9Yr0F5nm4w7C
hrxXXaelqi+pOAN3RxHrbsFF5bH3LT1bgZGZMstnIWCOQb7Y4SCBvLysRw0ceuVuUyvAwncX9YRV
25o+hVu1y9JXQ+HYrGWygUSwNt7lwK+Sy7cYJh0uoIHOqCqNiZ60g17sifi+MYzxA8baUNpMt0kR
rKg8ZTVDwT9mzpAPzVLmjpeJ5NfBtHwi7n24xBBLfxEUD9RKLID0pmYq0wlMFGLPPMdoi2RQd959
EOtG4tmn/QC0U6LWvCaiJp0m6P476iysJcbDyfjNXxMRwd0smwBiqGDkUXlNE39a0EFKObNe2ZDT
Zt8McxgvJk3KeZA+jFL0GxDZWPxrI/nScjuvMavCcuD6eUA23dEc8CpnHa07s4Kc1NfdyiPHDe5R
ltfPScb8FbMVt2WAdmjrCv2Fup/+FKf2fLaDRTWmVgTZS+jImPyuV0JVDfHBLz9RIqPm8NUG3COk
3eGbOsaoerFDUt5Y1onJMjGex8bA0LLyg5bTBzk9/RDuTd8UFZ/FS0HQ5XoejpL9skeLvsTNAONK
daj1XnnNwIpiBazR7fQyyK7EvpKu8oMB9uCfnLeHBS97xjtcEKENAWHPEOlZTg+Arp/mWibpLhP7
Zj5MLlPzfIbFpimuiysOwkCmtRcZ7qLi34i85/3031ZaBt9VTVesHZDGaO9ItR+YGt9EwLLEsVrH
PWcPe1o6Sm/25w91Yhh2SIDzUSfWb3S9CkaNRZ7n+JYEw8sgo91HulnT7pYB3gNt32DolwWf7c+B
/HxpFyJGY8bJfvXig639a6J2toKVG0cATogAUwtXNx5zTDkZotdIKe5CoYFoeulJxZpeYp1yr2M+
ounoPUPUlVeE/MnEGJi33R0DDfZrh1Qpa22dVq/QP3N4CvUKUVdXZAzCRA/p3AkFZLzjEBgZKgh0
p0L5q0e8gVGo4SNIYqFtbJOLn5k259Vwdyd1os311h+XLdRg3pAPY6ttMNBENF5YylBVC0a+d5hS
4VMxeSUdvf8N+8+ILdbDInBDn/YO2KoDtObfcgiecAMBcT8hF4BjOtwn4JWtO9y97RvVhPVYnU1s
pE524xJt53/f1BRNVw5z7u0dSHFMHXN4gIVOJJxY0cc9BJfmZumCj+At53IKiwCfl25P4tXzZQpF
MZgCCj1UUPAy/9205frBW8HrAS7wfm2I6p14XM00acBZqVd6xu3/drEGaPB79ZEsm8BRuYWtG5ue
CWx/4xn/RV1K4KJpvhPQxtOJ5Db05ai0Jn4uuvH6KhzuXqFUX2nf/1WtqPxg2Z/zML9BX15l3vhN
4HDI8XUCsDjEAQBKrOzfXhTOrCLnCSlnYbx5zJsSbd1S2WfWyH6buaWaa38lreDOARMRvG/rTEju
ri6L8iehHJLgPOVGP/yVZFf4Ax4SVnKXWrcZrM/lUMmpGGfGURjlVGC0Wiafs6biQ+Q4Cqq5RR8Z
44YKb7a+8LJSFgL68rhYOBEt1Tpzg4D5jx1y0bGzI2Cr019pJRZXa94nffZurqss8NZ0FeBs/j1Z
VzTWKz+fqm8feYGJOUTs4bHY+Z8xj0TuYrIMv1p83bQDF/8HT5WBhRjvKkgyLHVCE2CBsf6XdXAN
Ku/muuSXT4LIYDL0wLHiQbynIxDkTGruXt6r2/2S7HoE/v/of4dJG8PG7fYuLfOYZXk9401anquM
T8Kr4pRwuCgZWF3IIe2O6U0hal3tJLW9lFAHIeq8Y+/RsNyGb7UWbTCYUPUUfDB8kFaLSr0QZCJD
nGataH9NaNEy5dxtdx3+BD3mDcaz83FebSgBeogpcFxghLDLNEEH933uKdoHQYQCdtaVwP9XYlPM
s/2Zi+eNFA8E7VVaP+LjNN5U0Va1jLk0p5f4WnZNOQTdX4lLUF0ZFJoyWDI1WurK8qbGmPjg8Mho
ie5Ok3wDfe9DddB1Y50o7AbbWOO942WTFitgWPpcveuH1TEwpKe9z5ibawovYl0Pmhmxx4E6pVb9
ylCVGQCRNCZDXhnDCnlHkNV0nLvAn+Gq02Mphg4aDCZQcNbbnBxeFIIFI0sXP1YbKpfs/Em2b3yB
S6ndISf5igbDOCyVH6bZ9FdLEsC7Px4VVGzxSDlOyKora8teClWbLZzbrvP+gjyAXJTqy3i1Q6Z6
xSsMy2VkBpOnZ7gcwnHtI2WoSRXIJb1I/ptUQzAX3gqQ4Q9u24sTDcgXqkUrJqM6b+ZyAuX3/Hlg
HzKDiSN4jwopq0Z9sz9Yd0RDZSKqbXNn66r8cfmsjh5BmooacsYGAbr25piwggBH5wcsx95q6oKd
Hc7GQRBLH9tQTmgLD78G/K/EVIDQpSaZEkiJJ20KHMj5whil7CaQKr9OuYEGCDY691U7RtbAzzps
k91Yid+TmF2kNu/aKTAtu8AV7Ag55guHJAPBfMHV/vXDsGOfRbE8fEn15mnlR3LqJpFR3Q4OnzIf
VKoqsgXoQ5+UxNNrMK7ExtJo14zmahvomCUK9vZxjY+SPEIs/Xi+rxC2OFs7R5zcYsT/mRkq2Zs/
cJjPqDDWzL5n++O0dnS6NF1EZe1UjG1O8naKtvido4RuHhIHy2n4RL478KEy9tbFE2ld/jjDWwfh
02Yy/EZElz2L3Dy/lhughihYDDRibqY0lhUGwaGuthjfiR6VY0pZ9jXQIObyGAlkEmmm9o+N6g5s
Bqe7XXky8IkzRlWKHWDgPCosoPa5pvifjE5l/GYmP6d48Ubp6HeDLH+0CTXo7Tk3PIP8jAxLicAP
1pvnA0vG5zRDOlTfuhtjUoK6eo0BAjdYAixrej8mfv/W7CNPP+0WDuw5jNcLW4aMcJ0LcXJTZ/7z
kduP/liZ1OBuONoR39WI5lwxw2UpXaYFLgFTdAc0t9pAbBvq1AWNFIDLycaxRorcDaOKf5JayYcn
kPu9cCoJa+0f2sEWInsaX4ukdX516XvnksRGNC4j1AvvzlOejG3CaGMNXAgLqcpz8d8BeF7iPvaK
f9YOLUxW+uwQfTPqHhiuUFIaY3cXBWzfDxO6oZeuN2LaWYGKKgyFprTG5ec2vc07HMyQ6Ubkubf9
UzvOFyvTX6p/arwndzoEOYJJgajmsFCKrwadS52Lyc7lpe2hR/oMjcNkQt5wgNuIr/z1OxdpcUpn
PGNusUNQM4HRoAWzsKXA+IO29OV0UEf3c3hPY2uxjVWy/pt/VCvRfeBbhCD4dLWGQPuaVc/JHWlF
zVMbxJJUpHIG3TzPkyDYEPqhK7fnwRlt5jdEdlrLlOufscdcwPxH/OAw4eeaU1MkMvHj8l/EuHOc
yU96GTklJcU5rlZ19GQehYQAWkDWuu3pavVWQIiNNzTJgu9M8XELoKttzCViEHYR3eOAYtpVSGj5
ylNbWtPpi3En8dfYdGgnpOS8s0ZQRkBoQFvFAp9mBfajTaQECW70YQh9At1caahcPys+oUBEoN5Q
1bOrBd0aAvMM8lkCXtok5YwUq/YJ7ypxHotRxu83K0GiMb7CWxoT7SVv4xoHNx5xEEbiYi8cCBkF
2+XFKrsrp16DKtRwlocRN0TYMEMqKo673dt5A60dgUK/oPtXQPrhXMEMvPSTXm8u3ReqgCCCqaWs
CFFXb2Y68NqV56a4kZD4Sdp9tf6DYpktPblMSFKxcvsNLnpof4AU5dFvfxkwPq9eSGhorFYzBWj8
PtXA1Kl5HXZTND8rQ9A/2hrlJI+MJf1hxejDf2fnM4I/TME8nWljz2BxmVlE9EewuTa2DX02j80W
ObSKoiS85xMhJ+tWkX/ACwVyYmk/Y2Mkx9rDxxKDCU9Irc3Ho9SZxBOkSlJD8jjt5DCCXA+mofj2
rX/xEV0/EgBLd7inimijcPMhmAxMkegUhSSCJBmXNMcFyryrsvWKoLV0M5ck2eEhS8cUXIy1PnHM
bOyRZwuUtBAgxn0HkL4lQ/xq4w3TFHPaAoMTJ4n6ejrlJeaBsGc06J85AbgIgl4MJlha9ZGwCkbF
al2Cgpp25ceLOFx5R6E/F68YBjmiwszIOCxNwno5p/gdwwOz6hszEVa2ISJSk+RsxWRlrmnx+oLY
4AzVYkzJTb8muph4PW4p4h3//p5lEio8m/BoLZlwH3Pljn43CxiiHZNBQ1zRjZskcWt/XhA28qlE
M49AsU52fMRe8hZsNUb1HI6D8ZLVSeSxrT1Tm1gik+dwEqZdkZzXACp0waDDy3Wu0KiTSpGq3y8e
SVaNY93hdOlXrQMBrpqAeh85E0lr1QBmJTFSV6jBbvXodI3q2iwVR2v9gvQzetC2znNUdx4U2OPp
Oc24FpvUQk7tEAc9I90fb7u4+wwNXPvhPB0Agl0GfPhtvFuZ7rPLEJEZVc/ss9xSEe0T98oYR2nJ
y36pZIyS9tUjqH0Q+vMY1Knf1XyGmi6l8D5CZ4aUhIZFB5w+GWkRbc8WSThdDAzSfQNzaj5hBFuQ
nyMM6v7Y98QNSk+1EC4QB3Ngl9lJpuw65kz8oOOaYg2w3vHw6BsVOGQy53D8zkTXw44DpWd/72lD
k73UU1HGHUpM9SR9mE3Q8N/N8eFa3MnDUfCtktFpNkG215AVCg575FvcoI698x8+5qeAEZB5hS8n
l+jUV/VcchDKDK0Ms63nt/+1QNx8UqB2fmZgsAfw+y1mvEBKgJkUKVqgtJ93E0mp5uJGckgZt7yi
nzKOs81RpRoQlMTS5CYMhLnLUagwF7rfIVFyQoWFBDTso6o0W3GtSUYqT/QP1Jr1oSX04jHcZfii
7gNuBk6Qnoy0eVD2LXWg6GXQrFqGqz7SbDvewK6PHyT+hjyI+zANJv5XANbowrqsR/OUN9PLzb7d
M3JdiO7Mmq+GQKvl14Cqh2i6bc1KMi5Mf+cUcrh3QS1wqqo9LFAhpmKjSQB5uyWd4j6Hw5mwE9Qk
aGqiAsaPUtbgo99daotlq4DR4oYgAtlP6oNb+mGakKi0ork6fwWSDVbYrRufuSzOXZWfSSz6eF6Y
40iNJwOzMOc3yTEzS4mbdtyxrBU2r/8YzucS2kdbTrgMdjcKWLrJ1BR2XFQIs53BTTFBbYH7mTw/
jELWVVz1/jmztH1rJ7D5q1kV4LBmJCSClViH0Rpl8wxxINNPAVqkCNVdcPT9lDkcKMDeHxmY4iHv
BSGVPue9RaPRbmWqgELA3qOBSmablohjphxW37QqP/xP71J93A0nMnullZhGzeNOoGf9uo2yxfh4
88MHQ9SIh0Y8vv7v4N9bRoQ2A6sTKFi75KXMVG7LyP2oX1VAToo4Yr/FR682IgtPqRUthL2BKeT8
qeTFooOeBgNUJEjdm8gYip5YFydd59t3m/XTyhUOuRrJuTayVfpgQ5mrb1s+NRnxoknN+MMoWfbz
X5ThTK/Sek+Qek54SdOi81Cbd88YuPwImhhg2SI6b0aB9Eq9czCpCL4rEoRVatrswNgvu5rf+ta2
ZwF4LrvM3Zha/TsfzvXlI1P1+h6wLOfEK5O2pElzBTX89bm4f966rAK0+g8vgMZ/AG1F+9QyJhvS
KnIGKeSlgAkzv408ST8qXISM3puVY1Ipr9TnpWPjP89cx332qbQYiomkuzi4GWbpJhBV9tB5ACnU
3Sj5wtJR993dh7pUqG99IvzoV6pYbWtgT4KzCUOwwz2BDUvkh5pyNbjon9fdTPrwM1KL/Y1dT32t
5wggU0ZOlmsmqDCwa5r3pyjiD15a4SHMUmNIZl5uwlqNJU+Z+CXrE5CU60tnhkLJ7d/rgGDZpfTM
t+nqK1Z27f3c9fU5qhfUZbybALD9gPNZWNBsgb8sFY+jfWe9ONy6GFlM/c5ieBfrIEeuhxkdw5bt
XgvWIhfRkELHK5GEDrm5VtAn6tZ4tDp8Ei+JTfieV7x0cFK8OIFvDIPJJUIRJjDXlNLd5YU0q5K3
ZWr8B8JXOZjWRXQKQ9RUvqik1wAY4zOsBztDE9bS3j9I/2Dr/0VWkpslDbOxFvoO7S/RXCcluk8F
v1OXgtOrVebKt9GIIWu/EPojMHAIs71lSdgx5U1mIPcpkkH36deEKvqojpbqJfq8lSv/XniEptsR
ii3ZMci2sWwkAOUYTz3cHPPHfUkTQ+e7Z3p71ZPmZNIhVb3DI1Mwy4bHBEGl0sOGS3vHEjqtmoW8
axQkrVUQQSQy2Fl/3erU9fswNUkEnWMyKpKD3wCDXlIHOCWfxk7h019tLJwlMDEG1qaEiHRIXU7+
6G25MuL7qmAUKGRQ2FblCHtSuy++jk+ap52YvsxrCNlfCGx/BkJ8Nz5DhDUEC9sDU3UUeMQ9utTK
MJYhpNUgSxeB7ykJbxWJ7iHgkJ+ObTcQlvoXRSCGX/lhkIix0LZAZOqM2mjrgbCT/rSxYSs8hb6L
Nt9AEcEk28PbNwuRECFFEoESDQbyXlVWMmR4IcCjLBP6YrLR7hvE3/LUmEDwlleW/vjpi9O6W23M
4jfX0eXbiQySjqrqqNL9ixK89j6m3SVDXqzSbaTnHTgZdMgpq957S8zQG0CW+zxUIvVryL2tdAzt
WQAbs3E5HYmvlTKrxYRjT9qBDrXRqwaekqkhRawSzKpUBf5MC8NrU+wmU9jKKa1Kdw2yce7JXAdC
NLcIMTjgL1mCpC5rvAf1xLNXkJ33WKG5Y697f1KtHQWg0mL//vi4PhfLwvqU3PlCV7Q+ewyjs5Gi
q2Xf25r2jaVbJP0BXHcoujSSSlyUb0LaaWixZ3JQ65ox
`protect end_protected
