��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	� ' �SR��(X��6/�mf�չ��R��n�|�C�1�"�1Ɂ2$�Jܕ�'��J�#�J_����?j����Ǧ��L4� ��y�O	e�{G�;n��/�G�����4����1{�N�؈��z����5m�����P���pb��dA�Y�����a�?�4#Jϛw����})Ȧ��*�bd���!~
|�G\����n��C�<�u�\���4��vz�~Ѽ2(��hw�Po�X�g�b4�5��ı��/%)��]���k1FླjBi��/"V�����Z���p�e%�bN�Y޿���UC���noV: �o#�@��񝘈�~yf@�o��G���-�T����z��I��Ft��c.B���p&f�ޚ�<;h.#�%�G��w���)�^���J�6��3I�F�'��4.4����rh��}�s�)��Y�?Iю�h�w^��5�L4t�"��-���?���Ϡ�L4?eR�g��Z��=�ן���>��T��P1e`�6bu�:��<!ԡX�Zb����)�k�>���a{���/���jf>h�J��d��;��o䞉���b���"6<����������p%�{ю�ѹsS�y��yj}qR��=��<�t��w7M0h0M�.���Ř��c`In��M�2�DȨQ�NW3j�.�[x;H�<I�}
����'���\X����{�DoZK�SI|öbg��0 �Ce,K��z�ӡ��Dy�䥜]�g����@(��G &u �<(�>�x�r�2	�W���!Y䵄6�lw��Mճ] �K��%Mk�M����ǬZ#���evf�ؾ���Yhd��ǜ���<_��~X:x��D.��Srr\������6�!��}/�,�ch?|�nlv,�*Ds�������{�ǡ�!Z�%C>y}��!C��PpA�P�A��O�`���7���q�|�T�EݲqdFLP�2��j�Ʌʞ��z8s��	�B���?J�_��Y������<��Q���_x���U�"�u�xl�o�5����}���-ۀHp��zP��Q�����o5�*�����p��=@{ڱ"xVx��9�g]O]H �����)_���b���gp�d�B�Z�]�@�fFݘ�\���d��j^r���<*�)o�Z�6)Ɗ��!F0k�[J�$���3K�ʹ�*z2�F�ح]��YETx�R1cqBĆ��@qV��J���4d������
7ǐ�D0�mJ4]�4��T�i}���`����W��ML"@��p��F��1w�UĖ$4l��j(�)_x.^�ϻEzA����ȁn:��d�@��6�u��,�)q~���q�(�0z��==Q%�%S	L���4�ʂܬ�T��^39W�8ܐ�t���ͽ)�;��x]|�U�B!��Z�w�@��4�s��&ÛI\b�(q髚�h�� �O
:�w^0����e6f�pƮ�m1g��$�ZC��V&��X�����!d=b*�A�e�g�_�G W� u�|�_��4]��uD#ԛWsEW�E���i�^�@ծ:�C��;��l�|�Q��ɤ�\8F`���~3o��7���b�1�C����&2�|{����:�����		����BOb7!y�3��-�fN�<�JH�fB�p�+�h���㣌&��d���'%<>�ü�>1�W��c£4D�]m81��̻�Ѐ�O��_�D;�����4�xF������?A�=��>��s���J[���4D�Sl�>�zaA(����L_j"y�AF���X��i�H�>Y̒��ɱ=�%Ꮮ����>"Y"%IUw���*Q"/(0F�K6j|n��5�},�娖�|��w�F;D@�-��>U"HO���X������lC�[�:F>pݳi�������%R�X�<䁃�!LЇ����$�Ntq{�)��z����1��`C���y|{&aG/��g�P���F�Z/�@" ����3t�u��3�K[�2\H�t<?�w�Dͽ¬��2��%dwB���,����؄�ή����X�~�d)�q|f?ĕ�v����1y��jvq=�C�I�P�l9}r�������[,��|5���u��'*��ׯ��&._-���.�u
R_^�����v��>{m�������4���(4� �`��V@�6�m�##�$.��W�%zMV�99b��?��F-�v\����Ul[��\���������<H*?Zw|g���Z}Y���ۣߙ�T�o�}��,'J�kl:�w����sʮ���;\I�Ժo��d��5+J慇�25��I[��Y@�D���~��9&~b9lS��*�ӻ�I��h<oL�k�nn�3i�ŅIB��`i�S5�ĕ"��|��=�Bq&��е����AV&�����E�Q+��L�J��8W�X��{)3y��,dM�R��0pG���P!�qbk���0�&� ��j-��t��$4L��/"y�0���ci�,M+A�E'])�Z��c�Н�}�Wq��:��6�v�'�WvO�Ο%yOU�8_򼐘���ߔ��j5#����ל �8á����sI���S�ݧ(�?�p�>�R��&���r�s�ޫVYPzh+��x��&�p�ϸv+Ɣ]J)t�����P�]�I����P�ѡ >�����[�5�(�V� X�fA|�๩ΰ@�Q�����
�}1"�hр.�����"�^�T��%�Dۺ�����Y�]<��C��yױ���A����g���s�k�4([\�ހ�E
:v�P���>?t��·1��$o�#��N�_�ш��/^�����㭸^�G�!O��MZ�=���E~��l�;��{�)��A�U�{V���4y��t8�ѹ�Z�ie���M#�2�~���������Q;Ӵ�ԗ��|Wf�A�+�u�yZ7��Yx� e�q�!������Ѐ5pM�_�F�����BM�ĕ���o���ʨ�b�JSN#Gf�����e���a�g�3֟/no�ˊ�XӍ���S����nr����E��ݢ0^�O?�RX4���T2�Qp��v��σ6r�
Z��ٻ��&��q�VħN�@�Ln�@���%�R9F�V�in���&�DO�h�8-���<�O[W;n��9�E���^e|�I�~�[3�4��P�Py���y���e o��>����"�9ନ�t��t��#��$¶I�l{3�!�l,��:s6F�6�v����U2�G�O�q�:��ج��9�w�L��J�v�:
dO���Dc3���*�H?R���F=�|����m	ͣ�MB3Q��������
3e�������+yom,�M�����!����=TۧYv���E���f˫���k�>ʄ���7�3�}b╊1�"�L(E%C��ţR�y��fO2�պ��<�s�ܿ�	q+�*�Ȳ5�i˯q������p�S��6J��zSE���͌9X1���Ox��`�=��!��\�H��
慼? 1-ݞ�����0^0�{8��:��KMDyD��xo�&f<��]���?��|!��&0$��, �\�� ����fc�j�*b�D�Q)],��1(��mܢ��<x,:έ\|:"4dqCg��yT�o�g�X�1�j�W��7��|��=y���/��%Z�5�6�[/����wb�K`�?�Cb�:���~]����д�C�q�s\����̍�rF��R��j�R8���l[���Ly�y�U��� "B� ǳX`$�8��F��o�3��bw���4����-Ҍ�lk����������b�	����0�xvҸ6uQ���cN�� %a��S�ѳ������P�>�~k�X����?U�C`��x-���i�V2�a�Mu��[J�5��?��Ʉ�
��<�,+:"���H�Б��,�R��$�ZB��]�M-7?C��U�%�������:�`�2��
_�hD2�?����O�)W:�~��N��ڸ��N�'&���W��Gi
���?ÉJ��6� ��؜Y&�`����#�oW7�gP���Ő|�!5�1=��9%.�U�$|w
h�y���|��A���Ji��:`�F?��<{�����Pya٬Q}�d&3���J"���I� ԍ��N-x `Y�	�U���N�\��r8S���p&=�L�;�h~���f��JN	w�UbY.�}k!�0�
�g0��Lںj���
��N���̦��D�P�xA\�
��I�}�i^�yx�M=����b�A�w� �G��.�����1[��Ox-mJ��m�U��H�\�C@D�Z�+{�0�D�F~Ú�����Ɍ �c8�[�����6m����㵬��H���bՌӡ.H���7C�y��c�1lZd�"F_6��IU���T_���)qO���0��vw��	��t.km�m��c��"��3�!��2��uj�	~
�9v�VO����K`��O�{K	�� �r��R���`�G�O�#�*@R��D-���d���C��V`A�%�誷pA̳��)�Kq�)�$]8�X3���R��������Ɠ[�>x�[.����x�J��p,Qq�LR)��@���]>U�������5|	�����lG~�p}�g��'����,o��8`�`њ�?�����Kx�]�]�M�OM_�<zXy�B��Mq�-ǔ����N��J�����9�iP�n�͓�tZG�uz����|�P��x�(:lZE��j.��)�1m>D&Z�E�C���@�v
r /~{z$���]v�7�Ǜ�&�Mk�)'+���ik��d��%������?81�H��{��uTD�}��cw��Vg�ũ��c��Q��&��_��Rq�vIpY���4ϣ��َo�*6n��:�|]!p	t�;������/Z_�iy+�x�M�Ř�g�D�߫ʖ+�T��u	&�[ha�������Vj���A�?��K��R\o*A-�-�>�"���XF����f���$d���zY�:�0z~y>��굯)��66*o6�[��r�>xE$+����?s /�`V7έ���}�Ҫu!ַ�q�ǪA!��:�{P��\�%���z@w�~�gܥ��o�g�uȬ,�#0�c^!V����|Ȓ�Fm�T�-q��sLL�;(�7�YcCL����M?��+̀���T:�~w�O���E"-��@MJr��d��M�s�IL�f|�pi�#/�NJ�$�G�j�����L$G\6 V��2�++bO �P�a|�+Eԩ^ST�#�X�����e�j+&Cl���ō�)\��"m��~�'<mݐ��Q[z��&�AĽ.?k��#z8y#�
^�n�N�6Lk#�=�{�1����>5�v�`��h�d-҈μ���kTw�h�퀭et�$MT���1�h�f��9«��<j3ƷZL�y�~.��%�}LSs3���/I�/{�x1ɺ ��Y�3���ѹ[�ќp3H��XEߖ��ur!{MK�JV	�P����J�!�
�6��K|D�=Z�����$����_tE�fb6;�]V��&J��7�!ٝ��Ř#wq�J��?����=������`S4*���E"1�����@� ��O��}5i�÷�s�Ӝc1���DGR��7}Ļ>)y��U	�;Y�6��Z~�E�tytu�Y�YC�:�<P�Z� �T�����i�����j�W�$����%N>�,m\�����~���I-^i1�/����<5�\eBs�d����׻�F�)�03����	��^�Z���投�ɘ�M�R�# ;�B�Ў��B��	���N<�""o̰�e�ar@�}"��`��Ȍ�a�=�"�F��F��+�QKӥ~��LZ��F��MX!7�����P����:�Y�`�r���R~��Sj����4Jx�҈�:-̊�\�D,G��I{"�0�C/�a��W:xRK���K�$�y��mq��!r��x[w�O��Ћ^:a�[��,�F� +&S����*�	��~�5������AdƖQɻ)l�:/�0�mrg9��h�y�o��L�S�|�_����҂���� �M~�)=�fu>��0*����M+��P�Uq_�#W�o�ެ���L�{�$�3�8pe,�fTu����z�!�&�^~C#u����2 �h�a��^����r�
6��8S��� ݏ�2���O���0TPԙ���q~ٔ�h����<�_���jf0��×\x�^9��UM�ɇ��B�A�>�J�k�r�e�ꦴ PܧO����L�ve���� }�� G=K���݈[�������K��z�6�K���y�x�a�����oO�GR�jڌ7X����l��U͡kq�6���h�X)�f*XW����eF5�/ ��Ψ�ؽ�쑍������E�tè��%_�G8��?OR��{�'�p`T�
�����Ԣ�ӏ�=���@�#v�ܘ4bfa�a�6�tZ�v5�X���<��dm����@b>Lr4ّ �rq��a!��gE���~��U3mR��v��$t47!�svU�#��O�z�>���TyŭwPM1r����ᥟ��*���9�{~}W�\
pFu�Y.�kx�a=���R�r+e08�[*�Á�As�z�|oRS�e!Ur�25��5f�َ��/.��PQ������<Z��mΧ�m��M�e~��l$�������<�>rZrݾG�{D����wt��	�\��Mg�G�Q��i���o�g�93I��fܛZH�g1�R=z��J�hn暻2��.R���.1� 1��IT�;-Mն$^�?�?"�1�o�ā)��#�<f��Jl')q���<��jtvc�Y�����p��ދ�I���)2������4����X�����
3U	�]\1���6?���)t����H�<����0V�a�@p�7%�i���lX8:/�-�FK��� a�8���y��'(͂֓ޞT��	<S�8���1}�/ �݇ 0��٧AA]��|���@��HI�$Lt�AHd"Ad1��¡��ަ\A��&
�%���
��>�x?�6��rA@n��q=Wk��L|b\��ٿ����1^'s��(	"�-ް]���n82��;�4�������h��>2���6��[5-9���{�J�y�(��Ǐ��M%v��Lbc�`�����Z����_/|�`}�I�89�%�	]1�p=�d$,F	�V[VFp{�k0���<+��P 9��Y�ߔDgr�Y���N�ޥ:���#�=�G;� �g��#MB&�q2�Feq}v"���OW���"�#��6l+�\{�ڴ}��c���^��ƫF���g8���F�QJ��t�+��(:���9BR�X3��j�oK����5~O�Y�0�=�ܘRC�3i@(���@_D���!y������iy�ʋ�9J�<�
TU�R�ap1Bd�tk$����?"�\�lQ _�ӖPq_����Y�,Tl�;7����Y4�-"�6���J�"���V��:�a��h�r?PI�\� 3����8���8<F{5��J��n�%EW���Pǖ��|�/$B��`6�3�v�I��ņ0�����aȹs�	^����Hq�
i�@��!tiц��8P��
f����4�h��A��#�k�c�%LYX���5�z��>6�)⽓�u�\y����OLnS?���C�N�xʡ{�<[*W�����1 o�d�(��0x�#��� W��Z��h��ԕ8��a�gj�@@_�������O��@��~�����I290J�����@�dj�V� ���U�#�=9�Y=l#�j��8iG������]�s{{U�Ͽq)����̮��UM���T�	I!'����e��dY�~í�wP�Oei�u�o=U�{T�[v���4�2����GT�(]Y?�-l��:�@l�O�E>bp	�f���5*��淺P��M2��W�D�9��2x�U����%�~Y��	��H����� ���݈;^�ņ��̘}�f�4G1�Z̳f��sƸ*�[��9���, �$���F�o$�҆�>���s)�d����Oϻ[�{��@��	���A[�M]^C����U%��_��{�?7r���@y�p�!�|%,������c7d��A��u\1�d�m�y%��a5�d7�l����׎rWE3׹��3v®ϥ&�'yw������/�J�b�y �GU	�=zk o�tU���N��"�;l=e�~wa�]���[L�b�}=7s?��=
�yo8�am�N	<���_�%\�s�d3'N��o��I�X<xǏ�V�������tZW�v۳<��B�vOsx!�j �̌Ό���s��ѽ��K�M�/U7�X6	 ��H�C�#͖T�����(�Hrd�>����l�7?g�v�W��`�J��T���|)���0<{��)�'
.x~� �|[�`��N��+O@�ę�(L��_��5K
��DȦg�{@Ϊ"��ʝt=� �����:�#{�a� *8^p�2���o*p˳�����Vs�6|������QX��y�5[�}G�Y�n[�]wT��D�t��g��E�\�Y���/��f���](e~Yx�H��kd�����Usɋ�k����+=<?P��k���o]uX̾��ң���gj*�qv(]���tV�m�u3Y֑BF�m�S�mT[�5��+�O-�ր�J��U.d�/��Ѿֲ�1ɯ��b���Y�R ��o	�.Ƶ���ʻ�3A��SZ	��b`v,Y����mχ�$�7g�K�A_$Ih�����D�tO�2���}�:�n�/�17G�Z����ͤ*a�����ʚNq�7*q՗*/6Z⮚?��Ӏ�UA7�wGO����K��K�>�) �[��h��
� 8�у�^�hX�m�t�_�| �j����I|�tEM�l��*��hL%q�{z���G�Z�\ߩ���Џ|��O�2Q��9���	����~b%(�Wy��;��,(��`�ba:�܎���3M#DJ)���4Bh�4�	���bI�������i���s}�ˋ�dG�S���{ț��V��ȷȧa=�$�a;��j?�Vy�F�y4��[Bp���L���������^��g�:.;��*��Ք��l�Pg���Md��es�������o���ЦB�'����:Mr���m��;�װ�J�;5x9��d�3���}��9�Ի{�߃Hś�l��S�uW������(��0ʉ��Ubh|�F+Ƨ�����:�m�'��ؗ�뫾�$�L� az�/��������t��'��.�?�>%�S�W�ѻ8�"��	�x��@��	
�]�<ꠒ���XH��/���5�OC�Q�e�(�Ąj7zs�Z���	�����#�ܬq���eK"��۞4���39e�v�,$�L�)�ui, %źg�w�)A�4��i	_;���J��r�Pѵ�:W ף����@���0�F��	����U/)�\Q��^� h�yz�Y�&�-�K��#�c�ޟ������V_�?���H�n���)�M�k�3��̝�%��P����.���)�G[]��k�Ïq��L%ͮ�O-��:-))ҏ�o�;��A� ��}����2��b�<��Kj2I_���4 �l�<]K������5:,�M=᠟78�r�/S�lpS?��ի0�`8*V!W�����^��t4��t%,=�G�S۔������@}�ܢ�-%Y��Y��G�x�R]�!;o50���1iC2�ӗp9_�q����n�^��T��Uf��U��Ou6�&3�K�~��#�	H]Y?�Y����X��,s������uveol��^w�օ��I���m�u�Z��x�5r��	DDX�p�ǃ�d��p��Z��i��Թb�{M��gڂt��Z�w��Y�K��,��¾��Y
.�!����]l�ق��x�|�9~:�d<x�N,r� N�Pk��Cڥ�eڜ}gMP�����[^�{�Fd���,y�[�E�F���m��o���c��6T�-�����2j1��٘oJ����Ŀp#��Ҍ����db�;��k���~䍋��G~�J��֥�1� �
�=_!�r��x�"8%�Ɇ�̢�Y�\��G���A�*��AkUZ�	��B�����T�n�����0W�2�;O%i)�?��D �����6�"���.��>.[f	�k�*�<A�F�3��'P1{E���1���l(\G0����ہ�U�����$�֝� 1
̶纐�����3���o��v��k{04R+��&�j��ka�UU�-�Ã� Ԍ�/g�4��	}=�Q(T��_5D]j�7�Gr��B�ih��3���N%Y
����#գỒ���8;3,��F�q?�pZ�_Ҷ��RV{C��1q���	+�ȝmb�	��d����nǥ0��	����-E�&O�5^�v�u:1I��yq:���M���k�
ے��\93����n' M|^4!m<��B6��k��Y<��Y�g�a�!'$ڂ�صr]��Cr�ގd��iDi�&Ѓm��(&4�^E!^I"�cʆ#XWM����cT������C����+-B�� �N�0��{� ���ݙ���AƠy+��ƚ@��O�$�8�3MܛGbhe
)�j^�Կ-_a�D���d����^v�c��jgh���ŵ?G �Gt���?�2�@}$қ)�7��0l�%�mXC��Q�Fm���+�$���4�%�HBŔ/Q�T?�è'��tM�G�E��	����&�����)Xf��xQ����PH(]�� ��I�_��Ԇ�3�'��!=?�U#�${`0��Ҵ���9���Ů�����c@�J�wi�$��fW6����lL��c�V�qr��d�SHVO�S�TTʲK�2~����y��4�ʔ}����_�J1�p0�L�M	�t������Ƹ�{�B�y�H���%] ���
�4f&�Y��[F��|Z<�c�vݞ�mBr�
�HQ�>��4>�g'���_�29�12�U�DF��ʨi\ˡ<b͕���7>�I�/t�t%��9�GvE�L"Ѽ1��~��I���f��g�X;�v,Thߌ�	��f��}4m�;��������� 7��g67�b_}u�5�^46Y�,�]��A���}:	H�h���pvZ�]�!���`���u�hDh�[�+(R���M��.U��N[oMr/Ι¡���6�h�ϧT����E��Mv��c�6�E�s�R���4	bLݐ|��@��h�\�1�K���w����G~�J�V��i�D�T'a6+�^<�gX��/U�|ތh7�iu�g�@����8�}���o6��JE+}���#7�$��GeI(�/;�-�kaz9R���G�x��"|�7��.R/�]�\vҳ��?yP߳�UC6o�k �ꩤ&J?)b+�ז���8��$y����Za-p�L=R�7 �����$0��4&H���+�s��ތBK&6R[�r&���k�TJ=���J�8�$�W0o��پX0iO��T2� $��J��GW* ��H�-��D!:�l�vD�g�I��q�������T�&ǿ��gmốZH;� ���h���PL�p�&wN��Z<rʉ����Ddc)�v��ط����<)���W������iı�Ѷ49,Ͳ�6t��p[����W������* ��� ��m@������ɳ@����sY6�'�d7�\V0�$��"�ΡoM!��U�����[�/�LX��@�"��W2�Dp��d����U,x�/� \S���Āu�*06zoT�:̿�ﻉ��q`b�0��Ɗ}s�}�9_5UeQ�S��l-�v��MMw�9�Uwmh��PW������EK���r���ՙ�DFMtth��R�����T8g����l�^�  �N�����KO�<z=qu�o�޵���d9C?�vt>���~�����G�oy��RK���BX�1q�K`鹸��${'�7��K��~&��D�*�^���|���������C�ߢ,Qe_Dw)�N�,B]7::�>�:�����|�c\�.C���H�G�xh>�!����M���U�q;�4�;�{�!������#�������ض��V	� ����= ��.��P�xȜ��47�����_}z|�B���v�W�KV^[��U� �^j���C��������T��L�v��RJX(d�9rOs!�����ߪ�d���c���s��9���o�w�йl_��j47����Y��N��n��QP$��1��Ψ�.3��KU�80^���b���{C'U�5�?j?�E�`�5p�&�P���`�k�aNG2dKW\�wɟK��Sc��Gv�Y�Ķհ�4u�Y�����m)�����tL	��� �iWV$���0tP�.a�OC�9�xe\�ԕ�n4Pe�h�l]�x�n��^6k��1��$P7³th2P|@�&d]���J��;'&"%��n�Qo]�&��1d1ܘ� �]�_i����dB[3o��d���d�X��콀o��=�Rp���:�f��������Jx�^�؊~9�\��,�tk-���|����ا9љ1<��ʬ��G�q���Cۅ����ZG����|7&��ɣa���5
5��L�W�����_��W����GuP��0)^�&�	W��ظǺJ_�Tv���]�$�ֱ��w�����;�����@�G�՗������H�9�N�<R���f�����1m�kؠ6�����zy��o��6��~��lf��������&��~$U��	)�N���%1p�����Gb��Ư5��n`�"Q��福��S``�]�&�����R~Zx�cAC�ȣ���q�YGT���k0�%H �����O|p&	�p\T�F��0!�k�u�N3�����P]���� �����W�"^��VxBH�5�&����.:�?����C'w����qo,P��6��<�%U�n����)�893�m���Bq���s So�S�)8~6W����������3����,�4}-���ȿrO�$'a+r��mr�@��9��ԥK'���U����(A��o`j�ق]��P.%�<mlK��=���D��T2&��y����%k$�ܴ�}�O3�k��-I�w��me��`��$��$C�1i��tS���A���oj��tLڠ����C9S9I5��q������/�<�xq�/f�.���9T�=;��,�$Q|��538?���׶���u��b+Z�e�&*��5:�K�eb~��|L��weH�x(x �!�*� �����d���U�4U��,����ؒ�|;�.�'���aͨi�wN*���H@�T9M����<��f�斌���Q�R�јL
��%6'�1�K�bY8�(0��:�*�6okp'�Yg`~Ǔ�6��˫��6��%|�J�� ��'�Z2.�s�y��b<)#MU;����]ټ���t�#��已��\��le�%�z3�h�Д0C�
`�L�۪$Fz<a��C��eZTK��`x�\��J�����3D�Tr���u��)s���6=}j��O�o�3�3^�u��M��c��WY�u�k1��x��ۃ��f�����g{je߲V��a��-�/��uD��� i���-�Q���V �Z�2<��D}
�Gؕ�%�:�G�Kq�b�e��M�3"N���ѯ����=��1��R6�K;�v;,AҺ���3$�8xf0}�����-\T��WŃ"
���4=}4z�����?���d����Ϳ�cd�Rկ̛U&��D�o.䪟�m�G�H�$Z���H����
�-c?��#��Z�)�SB���Ș�fҫޑ�/(3���1�[��{�*S���p:�d����A�ܰ.��ʴ�,���5�NYɈP�B���,R���㭌) �?�dȭ� ? m2�t���x>j�����H���8�Ibve�-`"�@�VlTX��xU-9���3�,=�},�#�[Rq���p��=��� z��1��#pP<ƬB'w�p�����c�NAib?5��k9����%,9'5.��o�& �Yq�9�Ɂ�����ʹ_ݠ��Z�\��o��!&�g��~nҵNU�d;��q���k��'R�&�v�����,ؘ~�7�Oy�t3�ƱUAv�B���D���c�^*����{����� SЫ�Ɇ�g��µ��_C����c++�k�~�*�� ����NZ�~�MМ2z��{9I�
�(L7�/��y�fX�"��h�{m��}h' ���.t��v�z2	<R�p��h|؎��e�N���lm�y�����Z���_u#�׏zqD �����ҜӐ]�6���ض`��Υ9��ew�(����di")����#�����v$7Rw�#K��.�o�bl�R�����wX|8?5�q���BW�������z��g
m�:�4P����`�^ ha����Pyj�x!���da��-�(�
鄀�" +	�T�����:���7bp�ȢV��!�O�h/Jݬ��JИMg.� ᙅRD�:��f~E�̺cH^$�����������KZ�W�L�"L��Xy�i���6G�U_�(��Io�p�蓍�IJ�X$-ǓRpe���p҃���I��zceD&�����,F0 �L�[Hx;�G�oj�1�����#cR�.]����sM��I��LX����<��Sӣ����� �@��k7��P�t�%lo�H^�r����Q�JѢ ��`1HD�3�\���$�������sw�J�$�eP"�VF������',؃�+��s�'>�Ɓ�k�Ç�HZ0��r���ͪ�l_����?�B�>F?iq�2?�Q����X�N	вB;UY,�|}��A�N�Ǽuwg�Y���&YY���;���xx��x��[�1��œ�"V;����%�#(�w�2�4lW��� �0�������Ǟ!1T|�Q.�s[���;����Ȫ�JH�*ױ�)2o��t+�>ec�̇p�	K#��IҰj�����em��I�F�l��3�i��ғ����^��ʄU��u���M���՘�� ����R}�S#�/�Df��l��;G�k%���3i��$����Urn0�C�{���Q
�=G���1���o�46���i�y�Djv�����vIj��-{�q_<��p����C�7��M��ْU���FkB�!�w�d���>doU�qy�-�seh]��b�$���$@�ϸ�؉t2�G�s�u2���A~����%%�-zFl�/��:!v�t��o����U#7�ܩb���_�5�ӎh��懶ι���1�Iu�a�ye#��k@�{�Hç}�ޝ����Џ�%ێ6"�����7���z��H.vc��v)3|�$/�lG�Xe����@�g�����+VW=9��#�@M�C����n�`�z")��J��f�+�+�c� ����w�S���O�:�@�Vc�։@#u�q�4�cZ�Mv����I��������4����Ɵ���[
d �O���������e ��Bp��~=!.|)�3A\��a\ ��j/a�j[�/�y�~�#O�~�g银SC�5&9�O�~���s#b�ĸg�EŜ!����c/mD��c�g�$��eŕ<��fta}ڙ-7���$�1\Sa��%Y�����u`������/����ZB�����	y"K6�Y���s��ן��y�a���A"t��*P��S#�.�k�7B��"O�T���Ĩ�d�4�Si���>6�D��p���P�[��Jg�l�`"g&�^��	?{�1U��M�n���XT�|]��Ir�������:�$�+=ϐ�v�=�߬=&��B��v�Z]@/.#�)��!��2��&2M�vTV��*�kόZ��@r2l՞S�8¥Mg��"�ª��q�a1�k�&�(��3 ��C{��}A�\&b�qa�f^�#HӠZ(��ٖÀt{[R�^���-0F_N���>n4����t�N{��D�6�V���_�.߷����tot�~w�<B�������g��E��곮}�F��bь����4�i�.�:�vz�O-j�Dܩ���s�j1��G�t�~���<_�fM��������pL�hg�T)�A9X�$���l{L����"��cf��"Њ�6˥�C���{�d�xAx\w�I'�+��R���#<N���m�q��M�����g�KF�߾�G�_��ʆ��(l\c9�I��p�H0s����j���	�Wm^0`����Ȑq{_
�8�!�˥Ý�*vO�_�1L�~{Hm���r�frv��،иL ����$����vn���δ8g�%��n����7�نW��("�M��]j�5ЉF��h���h�<�R$ �wn��B��Ü]4Ք��@^��
�;�[WoJ+�2�/��p��:��H�]��[Ŕ\t~zf����U�)��7�.��m��.�is��H���SeF0���7;���'W�����YŕT,�&�@�S�X~dE/�&�P��e�֘�Y�nɡ��C��s%��BX�4�q��<��8�,�<#���,Le�U��iF5*�N9�����,<[��w:#oPWC��_�F���%�X�.�]�!@���oP���Q�� ��ULڞ�:�4?�R� �pl����5��ׁ01����?5�0��xr�nZ����5j�|znI��X�t�WXAT�_�r
э#���
ÁI3[o�c�ͦ�B'ަڛAuʺ�w���.��u�y�#Pu�I�C%DԺ�w�g6��lN̮�e<�j��S�!���RVhʭ�]�[	�n�]�����oHV8����ҕ�ۃ׀H�qV��UM��FCU�V����P�4�q�+��VHE��ljt�t��U	[m��˙]}��bS��>�	��Խ *?EE�sz�`sx���x�D��p�(�)��V��.�@<�|L�?��ۀ7�+�T��8���Ju>�3	Ɓ��Bj���+����]z��W}ڝ���-��~[�A�컐n�]�F����p(魛��X�����̉'*n�ϛ�N5�xxҼ�3����=D3����bٟ�:y}���D�"�=���*9����i�[�qΜ@�ZReU�L�d /p,\���ϭ~�����1��+� ��P���r����x�z���B��Z*C~ nQ�dc��]��@�����U��
���0l��w���Qk���is��ҟ�Wo׈'�?u=<WH+j��Hb�Wg��
$��Tv)R��љ��Γ��R�t'��'�Y�� �_q|����G�)��;k�ub��0d����<�e[��s$��EcQ����ǌt�P@Sϛ!�g�E4�L��j��qN�!�ؠ���6X2�ӳ�GE�%wH�@�+RJb2�׼.�{o{]���L��o��Xv�}�gA��	!?'nC'((s|r8�E7�s,��"�Yr,K?�A�p�6&$��0^����mR=�D�:i$g��:�
���vhS����ɔz�\|�m��HC���}>�Ck��U{2�
�f�#o����|��Fw<
ܗU�a���4����`n�Ghk&��+�W���~��!�?(���f�KHl�A�\�7J���c�2e����SX܇"L�i'��s�w��o���:r|̓G�È2Z���t%2�':Q�٘^7R�8��R���Flj���@X��J��+�`��ʁ�>�c�l��H�V$��[���a��_�di�胐��=3*�#E��j��1ȋ[X��h�I-�j��҈�`W����]#����_��V�v�7��	��N�WyY�b�T=���l ��U�qD��e��7�A$j��|�f �~{I�e�:*��Y�A����<�f��dR��[�Df)�2�����J���=�T��mc��!��w��L�^�o��Vƍ4�i��T8 x�V��]#����w��b��"�����wÂ����aq�Nb�	H
�0|�5��&R2��*�6�l������uOI]��7��ň��W:e�hZ�\�����oW� @~��0��5X�|�(f�N�<��E�.N�=���� �s��t�\�79+�K�[� h������9��DO��L�i�;��]�Z֓e�A�g�\��7�ɳ?w�bjoW��%{��׃�~E��n�
(�ӎܱi�O_�i�8�P�Mf��a���ܦ܃��ih�)\$Mu���]ñ=���,X�n�4/ �<�����v"zC�����>s{�P|�m��y���ט򧪺t��t�K�� ��l��|Y��-��Xu�x��J2��n�+/Z"v
�r߭`���=�x��8���I�Vt�����,v��� ��8��R�dp�K$S�� pڕ��o���v=�Ļ׀/!�Nɂ^��T� =.) �ū�j7�!n�s���s��e�0�@M�D>�U��u�L�(�=���q�h�6���7$d�q����a2��ל0��2�Vn�#X}p��?��	�Vb�����G�"����ƌgL�y5SR�*mgK�V�I>��I��3�Ɨ��lOGE�(!U�L�)��'p��:#`�ʿb]ӠȬĈ	��~��I��:�]���N�! �r�/�J�]L�
lm�u%��q^ʄ�a�*�+���t�&��	 s�(�Y.��A8y!OF��>�3LM-W��{"�q9"*�To�u�!0�;�Zoe� ƕ/�#PGC]��m�:z�� BC������p�6?w-��I�RY��M��b����pL��gK�I����(��$Y.2,{�Z������.�����C��v�U(�[w�����I 7y����m�x�@��T��]��e�s����Ԗ�u�8-.Kp0]���������B'�8�Ú����&{��b�`�i������65|���m�m%��>�>?i��E���A�TNpQ�e�ᘧ���y��?v-6v� ��|�s���2��BQ�֓.�(����7JPR��I����I����x���ǔ*	ܔ~��Bh�p�;u�U#/�@�7}9���_�כ�u�o��!Iڛ�)�9y�"�.d`Q��}���Z�.�	ܦ*���M�iH�p�r�ny�A}ƸU�n}u��y���&o@���GT%P��7�z��3m)Х�]XĬ��6˶	�7����^��k,���8cO ��`��J�mr�2�?��?�TL��t���s)_�k6<U���u�&���;�Ս.m�X��x,��7��Ŵ�׿����Ԅ�M��_��溊w���SvJ���<x}N�o�0'k�d0\���\�Wi� ��M�Aa$_�b�k6TKm�J�E�K}����<}on�4��f�ȝ4l3�+��PS`y�k�2���oY�����d/ز�ơS3 ���t[m�l��y᪸�] ��5�
��|E�������a�j]�Y����<��%��)�|�i(ִ
V�8t��[!�Ƭ�կX}}�f=B�[��2P����r+�y�_F��.1��f��@��E�����k�/U����#�������\�P5��7�
K����+n��nV�j&u�iT']��=W#�|#��VFo#������� �`�I��&y�0�zXu�@�5���h=�hZ�a���ӕ_E��0T���eB�4�۶0����������%,I9�l���� ��?�`����;���z#61�0%>�U��c8(D��1>���\d��n�(�2x��4�_15�l���	�Ra1	�e#+���4�XXcL�nzg����O�?���ثI&�-���gw	n���5?W�'�vx��O�������>�iw����E�)�٫~RRيC��Z������/��C1��^��Koҵ #����� !t�fZ���(d���;�_]b���G�=#���O�j~�W�r	�U��i[��t���1	�m|5ã�W���2�P�'I�
�?�I�w�� ��?�9��̕���L�9���(;��[UK���}�[���K�0�}1�`U�[DN�},�4څ��������!:�R�
��3�yV��q�.ͳE;v�����(������t� �[�,��ވ�rl>��������G%�h�NZ@���R��0lC�'���(Cy�\�Z#�܎�4e�DV8"�jr�}�������ٜ��� }��s��:�͝I���
k6����j�v]��&�1��Ĥ9��^d��:[Jo0�[��sm�
Z/�x'���;�AZ��Oi��!u!ɾ�H�ϛ��4i,�T(|��)�R�Ʊ�o�U����w/��Lv�	!S1-l_����h�/k�)�c�Z�*�4L�>�
��Zn�\a�3��o����6�r6��Z�\Srz�ۇ����M��L�^o*M��q
��)+�A��y���ț[��v���*���b��Z�X�2��77!%�x[/mT��1�cIU�Ku�a3�WC03ت�Ϡ��͜C�z�q��"��Tl�`5ӿ��e�RTZC�_�� ��-�1Ǣ s��=4+���xe���i�����8��|�u�W/yL��	�.�t�0�ՖVAM��<|A����"���f��{_�?��w�A�t�D.��1� ��
�;�%tA٤�8��X3�uM�6�w�>��v��w78�����
�L^&�1��HX_`��NT/d�/ؕ�P�)y&��JG��c�}�6���xg�:��~[�5!��׀��27@����9��:m�n@dwY��*��t��1ҕJ��́y(!�2>��I:(���Z��39��hC��"� �����70b�D�ma�ik�y��Q{^)�
��� ����0q	��\n?-�Q��m�_�e�
`��*2����C�í�0��t�d�}���~�B��`"� �9,�$H��������\.��;|\6��m�~3�o�~H|x���6���_%><P)_F�r*k�`����������yuy�'��OdD���*�޳}}罓����瓖q4��:'��=�[�,���و�[�NN���&*zLJ��m��C���N�1�q��q�������I�|��g���*}?�HV?|5{�7B{Ԧ	ɰ�x�)І�5�N�12&��`���F�;���6�g��Ȟ9j/��f�dEa���5���L� ���ڗ����Xr֤��|�M*�����Y�x��X��x��qb�E�
c��هs�[�I�q).,�n��U�C�!�[g�>b�N��xD'^��X�i
2O��p��ܖ8�[�� 9x[���+�)ߌb4H�oPƂ���5��w�L�i)���1��cA|�\
S�u�]�m��e���ٓ�>�- W�J����P��	��V��|��P�_��RvuYp/�	�D(}��׍�jW!�-�������=��>���.ɝe=-eP~��^�?��F�*�?���ݿH�LFH���c�����{���?ѹtr8�{�0
�(���y�(�}3v��~�K�+�+/K��*^0��:jN'��S[��L7����rޞ}I��~4'!YH7����?����D��g2�&�$����-U:���.;pQ�ه�PKm�5��TG�Xj�n+aO�}�[k�/��c8ǿ{݌o=� ��-���D8J�+���G8b£�U����_��(���Y"(��N��~�D<�z{_ꪹ�`�L��n*j ��{�o���4�Mp��?_���L�lXڂ׌����}=��1���
�N�iמ�����T+M55[�):�y�-œK@�
��;�w[S҄kYI��R�;П�:S��6�Фd�^�������i�?�wR=�����>�H��~�m����/, oD�β D-��2�|�kN�4�qqUW��VvP��U�4��ԋgĈ������=����)�6���3��y��;>�P�߉���ǡ��:D�&�t���u�ɧ�U���@�y��ݔ[ŐA���h0�����2X"�'ih��{&�_bh�� #,���2���r�2���W�S��ZM�R�R�~�+Q�<$����j3�+*� ������g��F�P�?K-y�����h�7�z��2v�;��r�0=Kr�5�xO����I[�7����y0�v��;�5
��,��n���ff���<万\��ml�.¨����f��h��>[��.���b7W�8Jrܸ3CF�D�G����U�����lF?Z=�ҳ5=����:X��ݵ$[I�<g<nq�5��vY�w��W�j%Tۦ��b�wÒ$�G���ѯI��軛IO�&r��q��[ʨc��o~۬^��_r�ԁ¢�_�����pzr��Dto�����@�$<*�>�X�x�B�f�crp%�&�[������=_�qc�;�zz�7}��,�j�R��]܉�O�����u���h/���7p�[����
i�."z�$�@e����0E�����(X>`^�6=�-�T�{�t�$T�p�G��G|2P�Y<H}��9UA뷯g��_��b�w�Վ��?���d���H�^V�g���ѣ��2���ŏ�A�`ē�s��7�R�/���a{��[���"���(��S;�O"��ȅ�0����z�M�J*��*�h�@�&lc?��л�0D���U�y ����CbP�1[h�x�c�>���2w��CL�زq�(�_��'/^��rN�O�!{?��4qA�uGRl�̭l4�)+ŝN��5�QM\�
�S��1C�q�|�2���Dz��{�Vʫ#q\�i�Z��H?�M��6�$�&��
��bP4���9�e�UԌ��~0|�P�h�%�[X��{�����o�������	�x�a�D����*H��9�x'����qy��K2������@J��QB���3���J��q������J�]�����X\�&��%�K�I\w��A���vu����޻k��%�'�-���՞�t.eA�f�0z>Xv�"���0���sM�1�7��l@����i�<�	�����Z]	V�#�pb��������_��25Ӽ�@�^�-��xGr��"	F�M���&n��?�Lj׼o�Ђ�v$8�v�+�ϳ��C�F�~k69i�m�r�Ɨ�m��jY��XY����0(~_>��<�<�P����B�����\�]�=��� 2
H]�I4��2�u�~�鏆O2bÿ,Y��3*b�ebt]P:�ǓL�O
���8� ���;��~�8��p����[�RH�/R�bbó���G�ͦz�q|N�Y����+;\��I[�wY��A}>��Vkd[���M�])"�`.��-R��9�ex�{�y�j��F:ӽb�f�T!q���UTҐ7������Ήa~d�W��{vV�*V�t�߃A�Oh�\��	x�������$��|�M����4#ғM��Jzp�OS�˨?���(���DNf5��ۥi��Ih�1�$�:Ft@���66�P95���l����T���p��	�`�dw�<��
̔ơ]c��pݮ��5k�������jFC,�1��_/$TH�#8,��?�Y
B 'k���+�B��#�
D��w<��rH��>A�*Y��p��1�u���K׷��*���\��ԉ�%&���z�Z��F���-�!����r=�8���kw�!ڬI�jB<F>�;
�4�(%O�1��F�S��nd5=������:���#n��p�����[���L�Y�@}�}��"�0�e�.z�,N��ٴl�P�&0�C\=t.���A>���s7��煹!��V8���i���ʱ���� 
D��q��7;�y+H�ِ��90�8�U�q6�R=�%1[HU�+�h�^q��Զzn:X~V��J�P��q?Pl�m�KХ���tm�A&���⾅��ȅ֮�'�b)����"�,��q��e1��5Wi$�ᨂȂC��2&D簇�2e��X0f��D	*��L�E��������G:	����|��2	H���Kx�L��_g��$| �oB���JDO��Kq��`:ӳ���{�-ػݨ�Gi������+�+<�ѶE�#�n�Ex���t>�}��d�=�
�Z���{~S֦EGb�6�S�<}����ԡ���0t�m}(�h�f�fZ��x*��3C-x��"�'��}�z�v����<7��x��4��>�~���sc���3�	$T8hf�[;&��>}6\&ĵ�p@�q?�`j��l����
�ğ[XB5��T'i���i��'�Y4K�'	=�
8�Q��;Fz�ln��&(�G�Z�DG:��y���v���[�?3�A5?��#y n�iXڷ5��E0q
��Ͻ�I-7�y����'8����x�,p"�0It�,%4?4&
�b�\�_�k5X"�!
��߾���AL}$�k�O�nk�m&Rf�}�Ղ�D���|�Acr�n�gA�����f�Cm�@�E�R���)���HޑF��"z7ҩ�ţ�߸N������C׾�#�� ��?��/������$��fx��%�;���7�����n,\S�<QU|T�UN'��@5�0E�BbQ�[h�~����.ÄT=|K����>1X�{� DZ+z|qј�B�۾�-�L�{�����tj�p��´Έ%w���=%'��)=T�H���~Yl@����tأ�5r�}įŤ�S�d �_���H��cʁС��i�b�fv9���
�u� `�Rҧ��Yn��\q�)�d��fO���݃{�%qEZ�h*c��p��N������S��#s�^�p-�� J��+
2v��2Boɕ�RA}��72�?�޵wst��VƝ���0p�k6"�qm`�&/�5�v�M�8�6�͗��w�_�z�n�6@�R��$V�!�W��v.%�$�Tc$=^X��>� V��@����>N�g�'P5�P?�DI��w�O"YD�]Z2Q���sj����S�:��}r)Y�T���r�,v q�X`c4ӥ��R �g� ��UWX\�*�ɓ3�H�Ɍ�Z 2���k�T�V^���^W�/V��+���1%x�z8���%�%�2��\Y��'nX��N%Jㆦ
�bZ�k$	Vp�u ��Y��A���l3t��`G�OS�'^LݱoCd�0%����jL�2.:���.?&d�<k�[��y��x)ģ�?�䬈�k�sG^���e̱=����u��}��(��@~�ψE�2��Oȵ -1���"��ה���Ұ����	��<���֋�)C��:�����w�ڼl�<��U�h�}xp<������8�4)Tk�nf-�·R���X҄��ы��|�8�6&���SLK�����0KC���5D�p�ڬ6���.�K-��@�I����>�N��p�[B��c)���~�C`���O 20�wEW�{g��|��6��x��?TǸ�`����Z�*/�l����+����GO�J���Z���f� �9�7��P���K}_<�`����֭3\Jy��7J�N�����T�n#����(fv���M<-A��i̼朼���tʺ������T�Bwj�G�D��I�qr1��q۾�_S�;[]�~zۍ	�<	kg���'�ځ#L&@�єX��_�g���]�O��C���QƇ*pو}�J0�>���&����Ճ!b]��'3��-� �EQ��AVo�34Z�[�)�]�<��(Aa�!���Y�h�5l~���	C`��ǱRo�S��lM��E6����ɲL�X����kQi�&I�-��6D	��N	2���;!�ʱq�O\�֭j� ��`}أC:��4�b{���R����BA��\�CJ�=9�G

�|��<����tB��5���N�����p��,�W�J�N��h�5�*\��$#D�6,�ش­	�h6Ji^�[�>W5��䄫�R`�z��Y���.z1�|��4�1���c���[����Kƶ��.Jb�(7��Z��rd�<�Va̜;�Iߛ}�_4�r���ζ��Ҳ</�L�Ievy8��9l7�H.J�&-�H&{�"���FPI9����+��
@As.�I�j�ڻ�K�ҝ%��6_�D��.��'���hf�V�����M�1���� �"/b��iۇ��i/t��50b!(���K����Z�^�q���*k^�� ���D�(A�ܨ�g���w��,�D�Gx�*�����:E�/G��`gz��a�'�7v��/�Vz�U�S���p8:�����9�/4�|s��$������_��	�SZ��
F
������;���{��/�� ��.k���wWe���.bs�Њ	������hW�N������H/js������㲸M������T�Y���_D�����/J��g���o�䱮k�F��
�9� ��Y�*vd5�t��䂑�5D��HMM��s��?ٸ��aŔ e?�?R���[��?�����&�צ�U*�����	;M4��YXe��O+kbؿ��/6,µ
g_&�@���.U,�I=dU-56�,�g*��O�9r���ٌe�my�� ��x�d�z�jW�Mu�
�92��O�v�yա,�͊Э���e������G�t�����KR@D5O��\�&-�2�"4g�G{���c�D^J��ߣ(um-���SJ<�Ʉj*��4��Q�xҺ�K|V	)�ū�B|�3Ӭ<�la1��� �CXOi�t9D�X�����ש��n�S[��`�B�m,)����$���i��W�D�>�g+8c��$�eyR���q3��D���������,qY&&� m?��ʄH7 �0YZ����-�N�Ԋ�/����lT�;����]Θ�RTe/��=��D�P���7)�d��VώJ���XW4n��L�e�h���mM��Y�Կz'Y�`��9[�_�1�zҜ��Nj[��"	����U?K	cz�9{V�9E\?x��Z}�sx3zJ��@�����'L5�^w�)���f�� ���~�@��բgY}���5<�|��?I�d�!�,�(�J#�N�
���v�$~�-�c@��C�?j)N;X�T䙞c����ࢽw�Bꏝ��=�W*R���@j��KX��oȓ�f��(�]5���z�}^�-1'�x�XW[.cNyy4��H��2��T�e��9>R?�@`綯V��ï���)HғcGc�Oҋ�3�чQ�Şe'Dh������/��|��(D�A{D/PW��}.�)�qX���Mu/���
".n�HzQŤI��H���m��,��PV���Wssa�T�c����;{��H؛���d���<ZE��.4������C$��D��H�,����g����+$�i���Rp�ԅ����FY��+�<S6�+�s+"暀�	q�)f}��=�n���`f�|ȸ�P�C%�=(��Y/ Y��� ��9�H��J%���(�A;�O��Fq��n�L"c>�����M	��D�kb����a�ς��")zi�#>x3��+��RA ���ؾ��x��� �#�NE���D���aӐ��t���Z���2A^6�T�Ăk�X��o�.�%J��X�2��A�_��J�����n�wչ�Ѭ��k����i�Y���X��G��,@��"���WH��a���%��#���i�9����V9���E-�7$I�C���mo�ߏ��ag�a�O��?�I��?QE����o��/�0����!n��[��sBϨp�oy�J-p�!��]�<�fښ�x2g�����FV�ϫP�SE�u���w?���O��0&�SG�I��o҆�N�	<��i�>����!�{�v�x��iJ2X #� ��L#��Ֆ.�gD��ޫ������",0ɘ%d�=*@pb��� E{��XZF�@��%D���%�Zb*'��M�y��b�۔|(e)
�-wn��;�:�w�P��_7�>�;��I��oE�TZ�$�����&���b�;?��:�f�?r;�۸�BU�XGRJuq��FAg�$
���"<�`8�A4>|�q"e~xi[�A��`���H�XDC��K���rN�Z�E�~|������Ѷ�U�����L�4�y`�W�I�W#�>��!�[�M_풊�l`v�� [��*���a�K��c�;&��cm��	�\���S�Dgvx�&H�jI��y�g౭�InX�>F�mݬL5%O��1�Νg���}�H8'i�� �߫8��e���hiEr�[`Jc]���$�g"u�j*���LMۧm	�t�/�9��#�Mw�51��5Mk���{����R�SY�_%����v�O@���n@��?�\2�vyaG����G��e0���Ji� :���eT���v��@�p���Y&"6D�/����C�����p�
� ,��+�)�9�*���G�]z�����qk�2�EVY�nբkj���,��w�ɴ|�%dW�ދ'�`-��3YYfĝ�xf�a%�p�n-ҽ�>4�*濈M]�,~�g9��J��_Ua� $��0��<[�_��M����#�d��?Uma��<�h��wW��&�?��0�a�0�VO��S����m�۵�YUi�9Z�S����q2n�I��8�ݙ�p�pS�p��87{��S���ų�i}���I* ����'*p08>b4����$�I?m���'�̈́R�=Č/LN�@�|�lܟ"�xپ�k�ȃ�/�_/@s��lm��A�4�c�W	���m?�jr���:`������Xie�����LU����˔��aE�H�Qخ�:϶U��,5o�eFM�<�ὰ���doB)�F�N�=H'��5��w�!��5��:i�x�J�4�W�� �1SrԘU��5	�~ܸ�0h�5�?��
=�����ݕA�x�jQԷ�h���R�a�����{Ԍs?U?_�묳a�l�����K@��g ��d�_s�?mO�܂��.�	0�!��{�j�9�� ���O��_�e*�j{�9��lA��V�d�)n #hI�'�;𷧷y=��{�#�|���2��j�C�w:�{����
��ז�D�y��E�t�����q�i��Z�||��'���-m�%��)�¯�Q�9��߅^�ʷ�¤&��_~ᐡh�*�!YїU�p�3N��{���$��+��3�
';-P���D��[ <�	�6S�]�txV���X�3�a��9� ��*���?NȮ{��rT���*twC.A�B��A�JuG	��a���~v����4�B��:V�����\��C.�+�a(9������ 4x��r"�o���
1ߊ���������Ǵ���K5w�����NLp�+��$���3"�!� 
f���o�{CH��sQ��I��(���,N�.b���),+ݓ#��
 ;����*?��M�
U}����?U�->�'�<諧���~�J齰��k���m@�SY:D�Hp�/[�,�mP��p. 9�Y�+*SѤ(�kt�4��W#@��M����vLm!�A���|��Wv�k�O3J�W��P+�1s\Տ�k�M	<#&`܃n|�E(��kT�~Fy�UӋ�)z׼]�w̸�̵S$8�`��J^�?)�Q��T�=޴�C���5�J0x�R?`�_D�n�\�jf��8�T�, F�l��g�d�Ϋ��[m�P�"t�9aG��ȩ�ǂ��1޲���^lOn�z�`Rww�A4)���eOXȋ���oe�[��b���������C��ŏ/� L��8#	�Ë�r��h�ɪ.�i��cq��l�Yy����9+�_@��-m$�$�S?�? ��L���
���ZؕA[�i!��
y�<�*$]� ���M�3/�k�����d�(80�gH6,����Ҏ����ʀ����������X��[�2�ߵ_W��uq�`[�*��ʐҏ����_�y�۔�1�,w�nDxڂ�^/mUX@��j/���2�t���!�;���΁dݱ&h�p�����v���7�X��}}��-;$�	�YE���85���Y�D\��tc�d�����;�U�`�CgA���v��1U����\�C�Z��X/�z �/��UU�<:^&iǯ� ���R|��\�s5��	*%^���Զ�m��	��*�V{
C��Ҷ5Cp��w��J�z��{{��k�:�Y<v}
��u*K4s�O�|X���-���Y��d�6geW�L#�!�o����w��ۀ-z�����8���C�w	��|�LO���e�r����e�M��6	Pg]����W]Z���jY2J����@꫁�҄E�n�� C 7��&�5J�i���~sD�ŷ�m9��wq���xv����ȚM4�`��#w�U������b����K,
2F����u��ῠԝ��R>+T�:D�˓�±�& z0����6�r*~:6Bf�H�E����(�@Z.�#X��,��)w5!��ٸ�����&���*A�Z���q�a��h�RE���׮o���+���,1������pF�S��%얡Ӹ͟������i������*���1��}��K��<���P��iIvbޮ���<���_�5�X�����h�f���B��6�M�@T���	~�����K�Y�0�ٙ︿[�U�>�CS�p\`�r��@@�a`�G^�)�SL���W����ʿ�W�r�ik~�<Y��kJl.䌫�C��?*�Ǣ=����7��Po���֯�'���/H�JOn��3NV���YyP��x��1�j'�������,̲h7g��3�Y|Sa/��/&`�2f.Y�J�|�q�W*�3�\zJ��602)C�Z�Υ��Θ:�������e����%���U��{$����Lh�3�ʢ'��-�k���j�Cl���T8��>(��9��B�Y��U�k�V�>�O�\{�^?�Ci����f�gi:i�q��p(����p9�[%�u�l��	G�#h�_�F���R���P�#dY�a.��`�D���q*mB9 ���U.*�+)h�_ JRw�����S���Im��qe�����Iz��F��2�f"��ke�l���A�f�mm���V��� �:����o� l<5�;�����>B+?63T{l������0��O>v[K����_�n0�T�Q�
��I����¬j�w�����ȯ�B�Mb>���V-����De�-�O�U!=/��fj�%rb�5�<�p��gR� G��s �w��0 ��|1��%��t�\������B�S�7ޠ�=�P��!vW�(Y�|i��D�S��7Emy�`ƺp
�➍�����jg�そ�ǆ��X�A���/��n��E�ӗM��1�U
������D��d��ٝJ����n���5��Hh5U���+�6R-��]�E]OH���L�F%��H�~��GK�'�O�2Cp_|3uo@��i�$��;a0d�$7<�Ἲe�LǮ��"`��Q��r'��g�p�%Uv��	�e���]�CEb���T=<�n�y+9i�gHԈG�jy��Ω'}�5X4�mk?��5c،0���얥�̨]?G����a1/VQ=.V>���3�H�A\�U��p��S)�v�E��pK��Z֩I�P��\љ��F�(=zH-��a1KO
pIQ-�O�'�ŝ\�A��Y�ӌe�La]`�D)N�(�$No�o���J�d�K:-0Y��Ze�����HD�B#���;���@���i���l�r�-�����c$=�IᎫ��htv�l�`�>H�E�EU�*����v����_`Z[�� � -t���he6j�v�RP�gi!�,�Nն�`�*���߽w9N���^��Z����n��F�h��{ ��.EQ/��S�汧�Ɵ��>9
��,/ؤ�]}���ƏB�	���K��L��Jۂ���)�[�+y��(T��&B]4��i�3�L ������C/�Shk��F(,�������ߔ7a���:��l6J/�Z�~Зj��VJ�_CC/ �9<�fl��è��	[���Iڲ9���:�zd��/0��T�j�����DM5\S1����&�%�=�����pj�n&���V�H�%�"��◶�unjHU�r��{���{w(�P�m.�k�j��m�J�^g(��L��Pj��r�'2��kmך������.�f��ɒ������^U����B:<-�`'���p�I �T:����� �p���q��jF?5�i%T���G\)1]*՗hk�G����3�k)���븓�%Xy
�,�E��(؉��]���[CH�<��GBEh6��P�v_��Y�z9<U���/�"�?��R�vC�
���!�oHEj>{���~�<)�sb�!�j����/w�hr�dΦBۘ���=谱��mյKݜ}�ǌ���[IƏ����Q�`�2���W2�4�?�m�R�����|��A��e�9w��
�A����W�N�
-ZD���\�& ~*�kuxf�]ډ��2~��j�+��.K�ff����Sd�ߕ��梕��郆$YH��TN����Et(�A�Y��e�fXE��U�ո@Z��[Ds��;Qi8�]�{�s�'6���J>�+N��)ɋH��v��~��'����6j]�TK�+(%�,������9�e��|'+�s	�>��j�,�Nk�R�8���.Õݢǈ��=䡹�BI�8�����q�m�ĺ�EH驱wY�9��8� �iv\Xav�|a1�T�C�a���Q���ؚ>�/��B8��$�y�b}���ꃾ�,3^e�R̬6��b!I�����k˿�,g �%�QO�En�%�_a�E�'<B��W��S���L�B���«������KQR>�_����j�N����$�9�:�z���C���f'���A��1Ɋ���2岖���!�Q�elv�A:�?�]�[�f�}_����)�0_lM��,�a�M��a!L��k�ek2��:�������~��W��������Z�[��b}�=jߩ�Cݪ��'Q�~�h�ƽ+a��c�hTl~0�����u&��A��q�k)n&�y��_<7Ͽ�Eo��G�T�~-Op
�ߛk�|�D�35�{�-)���x���=r�$ ���amZU+4��fȺ��-jg�f�Z!8ѝ�;4��&5/=�]�7���(Oj_�d�c��� �?E��g"��E�X8�Y4��Y��,�&�v,�0x�.D���������H���1i�l@�i����;y^؄�ʄ����%��&Z�a �����:&Y��@~��V�Jة�����������M�#?"nS��f��bj�vX}��n�$���s�>��3w�d����Nm�]��'�i��f�ITd�/l��pLZ�FL��*wj"\��8/��o"栂

��;�9�gN	i ܜl`��av���	0�A�0Z�j=���l�I^`��0��i�{�s�"��|Q+2�Ȕi�ݎ؞?5(��u䔯��sk���/г�����d�?*#�2���������t��^b���7����t����3��1$6_�­�K���PU���&^�;�s���H�ҧm��0l�.X	X�q�ΙWT��y%Y�y�
�,�E��s;��q����a*��=�' So��eX���I���W.;$�KD�7�S���?yp���؃뤰���"J�N�pr<!_2��,H��C���P�\�ԥ����r9��w$3*�������s̒v��4[�������x�L`�Isś��Ro{�G��n�Gi���h���
��d��Z�C��ҹ�"�x�;���3�F��̕+�}��	�UU������O�O���S��ΐ�/�q�����A�j���W�G�Հa�#.Qű0d� x�::w�HN�j���<n���`��=���d �H�&����_��l= bE�_��������
���60t$��)x��6	��n��/�29|2v���1H��46�u�`�}±?g��(����*�,��w�B�ө��S�;oGѮ�S�s�
%{X'����)���� �քX�IafM�I��X3B6t�D��-�Ȧ �N;N�)�������J�7����׸{>*%���6��j�wjB��a��᳘j1dQ�(xqnCCj���gx��"{�$)�A��#�/e?�G�ԥ@f�a���uO< �t��r�O9��c�a�1�`.F<�M�ú&�E�^�4��h��n��� t��tJ�N9�wRf}ޙM"/%���I��sL&���a�jIÆ J�����2���3��B�c'�M��3�ut����݅ 3"�7l������5F�_�����o�ț/q�A��y��؉y�mG5,}�����~���C�T�=��Q��d�F�a#�b:��F"Yd�7ڥӖ����Lƺ�rL[ym���.
�E���7�g� ��\~�:I��i�Tj9��ݱ���:�O٘~6����#�3�Ş�F,����Ǯ�+s���w�����E����k|Ԯ�X�o�p	� �l���0J6٬�=�e>��P��Y-u}O�����g��{�V㩪�>���fm���=�>��H��Y9��x�g"(�5��_H��UkZs�@��[x�J�Dm�|��������h�f����I�KDa��͕Z ��j�0�}<9K��Ý�����Rb�p��7�X)�r� ?C���|t����9W��V�夸C��'�_���X��L�kT��Hx֮��h�v:�%��U��Xw<���/wf��_y���F�$���N��<CjB��b%�k���J[�5 &st�&���S�\�lǈ��\q�Q�V�g�gr3��﮵mYb���������l�����H�yD�ppӏ���7uX� "a�.J�p"��y��H�R][~h_c)T�_�$c���@sdҩ�_\��� �Qb�܄�pO�.ilڵ�_S@φ5��R�Z�v�p�1����[
9Y��GM�ĖDzV�hf��
�ѹO�����.��C$��ī�������4AG��sM�ǎ�;Y��O��b��f�擒����V;^�d�qAi6{����w
��{�q���h^),愑�+��f��n�\Q��� ���m��aY��i��m����05��?&e���t-.���^L�$��w��mU��|S��M����׏HM��ݲȌa	��ƪ a��� �Dnp�n�{�7�Jz��5�|�Z$W�2�?!����\�fr�a�����v��*H;�G�ZC�M���nM���D�<Ss��ׄ4�o����w�4g��`CV�,*��S�����!�������.#>r�D24�&d8��{��2��T�G����lO��?�5�B3!��~lH)�N	2���.΅�,,;`��#c�P9�X�a5�+���6�Ef��r�+�!ch�ȟ���q{�,�wRE"��7���HmA��Ҋ�_�}	�k93_O{� I���qW�k}7cs�,Y�V�umRt��^������i
ͳJ��K.Z7-�ض�M�m���~�]D�B���	z��2����@�F[��=|�k�T�Ky�{<�o�Д#���|zM*��X^f�X���C�r��T�X�#��Cw�)��,2Gu�
՝��t��AfC��{妰m�p:|�SI���4�|�f,J|���	$򊬛#�I�{�tas�4����d� �z���r�j���	�=�z5s�����M�tQ�+�e��Ӧ�a�c�%S �AS�#�%��u���Z^��ZfH �x���$o� /��K E���>PYa^ei ��/��U�X$�ea�T��k��5�tnՙg�q1]|!.�Z�B�����$o�ɞԮ貒r����f:�^'Ԕ���u��T"�S�+��'�Q��.ö&�hV��r��<B?��sDb>��ab���o�g�8A�����D$��̡�(z�%�8�8������������	S�&l!��'s��� �7c;������`V���}��1��Hu�Pܽ����⹆}�\�-B��XF��ZR HZX��<��X\)�6�=�l-��$�?17��@���<�S�PD�U�~r^<nJ����P%ۏh� %�}�����G���J��p��Ɲm&&JO"�\,Y�x{����\!��λ�R&ý�سs��	���>Ȍ��"������V�ϫ@n'��1	$,���mR�+��%^3
8G�yu�Bw~���0si�,��дlG\;X�د��6|�Q1yGs���l�08H㕼�d��H�GR�\r�)xX���O���݄��U�S��Xx}é�{����6*���c��uɛ�u��U�Zu��Fu�"[jANЋ�j?���|#�ð�߆�� *�
�@,Ew�@k����@_p�J�2��`�o)<
mJI���O��~��41�o�
sk"�G�A��#��Ue �r0E� �4']O�xP}(���,�� m���U�!����+�
ᣪ��
�%w�EU��4m]ṡ��] ?�0{�������E�V���P-���@r`����t�$<��d
B�ax��԰=V�6���p�=̬������2�wl�M�5P�#��a��@?��2���[!�k��#�Gv߮|�~�)U�*zw ����A^e�����ڐ-aU$�C<��-_.�&���mx&�|�D-��QBL=g��b��=:U�� f��5Lx������J��<T~����B}�!b����O���ʇE�joQ� �>{I�G5tj��͂�z�)�u�-�&��q�K�ݔ��#��,��y�0�'~32�[�A��D?�u&(2�uƸ�}K������׺d�yM�]v���HW�.�����8��ՁDI�z�.#k>a#b���G�:�(�=�����-��bv�3��O�Xa<�\kl�d8G��)���H���(u�dx�sUz|�*�A�dִB��n�����a�����f-�M.0��nM3�_��(��e���ӰN�û�M6��^��JZڒ:}9�
���XKЕ��|�n���(�-�s�bЫ���WJnj�\VfO�I.��0��"�ضv�����U����0P�G$����H��t�[����m��
:�fy�M��7q{��c�,��?8�]������P!@{�hZ�Y�pm��;�$G�x���/�wvm��wr�Z
�#z���)b���һ3?`�4`.x�µ� 
��[����#�0�*�v��7�U��G��#��6e^�π�B�mǔ[�ȺB/��u��d�#�#Y�ե�[;�`���B�2h=�䲂�䱰M�5�� C������88,��%��"�υ�����Yg��/6HGc���6�ap�Y;��u*XPt� ���5sMHL��z�i�*�Ay��[�Fg�Qv�
}��;�^���.kakHy�fU~�7�_�ӫ��8 �@���a�S�:0=嚍K����7�5nc����wDf�Y��n�hD���@��Od��_V�B
=�H5C�rU�t ؽl�d�2G~�����Ֆ�wI��&m]���r�51�)cp�U���]k�,���!��Ry��A�5�z-�ҫ[�xD&I�Yj=��5���k/�ͽa��T��J\�piY!4cN�J�ƿ��W��Bq|��ۂ�O6��E�l�r�P�H4)�leH�iO5�q�/��f��%�Dum�p c0�,Cnc�0��M5�@��_pI;AIo|�x޶ׯ���:@���������!�
�f��̢2����gI ��y8LYBP��ğ9�j����Π���RtN�ee��YЏnM
���ɷ�R/>�~\ 5�K�jۀr9
f܃�	�U�R�듫M���}��:d�$���t[�3H�C��J�B��������и�8p�&�}�XeYpm4�vػ�p,@�os�e�	�\�La�*���.PQ�]B����d�<2b�)�<=�-<~��?Je���. �9680+Cp�
0�%��7Bw��H�1�Π�6(x�/+��im�d�m�Jy#d:�;D#��yB�TgZ#�N�{��H�.
Ӝv�s( ~��,��>�lm�s��������)�=���x��݅6��}�F^���Y�dUf�<����-Zt40l�͛B �n\��)���l{����Şԛ��Q��$����
�f�`���ۮ��?:ˋ����P��{�ȥi����N�	��p�(I{9�GTXc3�1��̀. 6X4�@(`�O�f9��$p��=��Xɗ/(����I�0	p7���D����ل9�ސ��g��� ��f(�Avr��;��p	���-�c�J�ſ� �S�("��#�J���6�����Y�T|�s6��ۈ��uC��N�t�N�Ol`?u�;焎}�Љz�=_���/'�c@��ku���S�L�z��G�D�v�8���.�ܚ��넴�[uQ�%��Fms̬�(���+"��`s���u���a�ɣi�3����� �kiP���X|�S9����^��n�G�`�p�fΠ�����"��JO����Y���?���R�>��,�w�h�#�?k�=����d�6q�|���A���YY�N\cy�h�+�6�/�#�ֵ���od�)��=�8Ev�=��*-Lb�����9x/ƹL��PJ�B�;Y���1U�HbJ����G�;w#�qR�=�[ ���$ \z:;<��z���IjJ�i�ZZ����E�M�-�B[������L���P���Dg,Ws� ���t����]�U�K7J�ã��U0	Nc���U%X�ep7<U��Z�����1��F�R��3��~�(���@!�u��"�!`%a�3�����$eE���ү���U5-�ES��fX�&ِY����.��bbk�2C�T�s4�}��iS��8o��+�.v����U!�o�j�Oeu�d(x"c�j�=�Za�Z��O��1hN����n�Y�L߷b�� vW�`��lT�9	M6A�&��>��R�?�^��xLe����=���>�hx��Sc��^=�}����=�!���|���!�B�$�Wi���ͦܸaY�V!J\���ӌx��P�,�R:K�g8R#Է��U��Y�H&]� �uH�TѷH���Y8��$\�ً�p�i���Y*��8�����q^� �?��O� -	�9�Z{1�����7�?���6���6I��;	 ��D�z߾��2zs۞�s�H�寪�t����y�=4@lՉ����OSB�7Q��C�}��<p��.'��gBPܴ�O��\�eY��@ �֫C�c�`�5���su��q�bd�x$��S�dKŭ�]G���݂��rq�x���]��]���w���S	��OL�-������f��{s"�.����LA�,�Z(���������4!�r���7nr.ᐢ��:�r��+����L��Q���j�R�uY}��q�/�e��f$��H�R�?�a��X�~��߱�m-J�M�&�hط~�B�U�&a�ާ |_Eu�ԕQ��b#�
b����J�F����� rOu�Ι;<sq;pD!g�6ON�M0k�����Й �v��!��b�P��-F5~���Se��6��Č�"X��9��&��
ɜ6���������g���,HR��� ��N)���65p�#�C�]��J�M5 �_τC���lu��h����ӴE������/SW���}�>0���4=�Ͼ�i)��Y�:�{V���;�k��B���HF���К����H@�3��4���W`v�ɴ�ķ��)�i����I}����:��e�s3�N$��6��qE�箞�xB8ԫ�xmm�8m�v�;�Y���n��ѥ�I�h@�Z�nK��"%�h�9��eH�l�s7�Ǒ�;��P�u��!�n7ng�p�T	1���h���QP�L���t�+��l�[I�No-^)�m-�����i^g�I-\�('�h������6_R�0Y�$���I�\|��e����jtŝ������/\�J/b�I9/B#Ki'�}���=;ګ:��E�`�M��m~qkI�B%���B�<�1��S�jv1���St�I�C���&4��7�}��HS:���?�� �PW��o�4+���g;��T��񉂩ۼ"��d��w	���X3��a|�;l3^:��[E�R^�\Qu�|] 93aZƆ@1�Y�q�}e������}�}�4H��2Wp��.;�[��ž�ffo3�ѐ�wǉ��3�,o�6�k��o��ŗ���X�$����Gtbۍ��4��b��@�6�hl�R���0�W�-���+cv +R۽�Y@h����R~�v���� 5G�g�d?����~$��p�v���1<T0��c��sp���$Κ�C[%�OaZɭb�%�D��_�ҀR�N7s��I�i3��$Bޛ�Z&`��_��o]���޼��s3ck ߓ���K�gY���D��Nv�z`]��q���^g?��~�=��g�����J�pl���+��]�X�q[N��f!z�ɷ����2y^�mKM���?"	����1~��Ƙ2�3����1��:��U�0���-R�Q�|:bHK�W�,dY[�1l�XM�-��ؒ���ߕ����f��Z��E�"Macz�Ί��,bſW�X�*�t�ݍ�[��� �5O�]X X�h/_�Ӕ�\����#��S&8���9�3�>I���[=f(�V[LX���Z�¸vie�
�!cv��� _E"鲢Rc��w9���gʭ���Hv)�����.\E6��7�J¡Lew�KlD��&�Ϻ,h�ک"�*���b��b\W��?'b����xB�U�ԭ~4�M�M�����X�����&BA�x��b�\U�W��ҍ�@���ϕ�s�������v�D�E�G#o�~y���Ft�q^dֻ�1+�Ic(6C�4=6�	����c���v�e1UpN�i��W/[�u�A�a� kڱ�����6XHA8�Q�lq���/�$�H�2w�Kxw0Ͽδ�����E�6��Άk��^֤��̨nH?�d͒�L���-,P�X�
�G
�A�)Q�H�#�=r�T2#��f�# �ä.)�X���d)]�>�"#���x9K��z[<��1w�f;��2��V�Hʚ���dE� z�{N-��u��Ti�CWu���?��ۮwؘI3��<4��)1��S�4�2���2T����Bw�c���t�^)�0�}�C�[9Q�v�FN3����?�D��_��ق���|��\}������w�Ĺ����uL�V�����ĕN D�z��=�,���O�����r,|���Ϝ��Q�n�A?�@B��3���q0]��Z�-^���41Żv��]��*�#��l!����zv!%hp�52����k>8[b�W�f���]�����g�̽���?���oҎ��g��j1L���S��lᚥU�r���'Jo!�n�mٯv�A�Ӄ�b��V����&�+K3\y]��O��gG� q��*y�:D����[�l%�/-��������8o��%}��Xb�2>'��6�8"�n]��*�����	�	) �.,�D�
�g��܂tR���CVP�;���J�e�wsx�`h�c�l���� k���2fW�% �o<�Zed�nQ�~0q��U�.U�T��n�*� �d=���y�g;ԅ�O� ���MV[w<y�v_G0�]-����	[�$M�,o��	s"�������?��:i�o�R��k�-�/���U��Ԫv$ N�F��=R���:J�D[�S�ȟ>-�[�Ȧ^'�,k�<�~�V�#>ڰ~����Tg�r���2:����k~�uɫ0�������h��-�4�+��u�@�2�c��r�T@e�W�d~z0��jU?W������F!V��w)�F�&ר�"<gfy�.�8�-�V�j��k�z�̀}����/v�\}Q��=��⬣9hq �i���c-�O`�G�п�
\a��F)Zh����a-��c(Fq:%#��,OBiݥl�M�C�־����{�]��k����œ�����HR�/ζ�d�sdS�Æ�cg�"� ::oO�����]*(���9�׍�ʏ����:&������>ό�nu�!kx�qI
��?�a[ٖ�(���/�Xf��ÐC�[?�-A���&R?�ubt���+��b��1���P{���WZ
-5d�C�%x:�M��ɕ����D��jD�h}�]a�MK$��2�Mu��t��f����
&�$R��5s�E��{Z[n�}|4",��[.֮�d��&."��U~l�>W��g(ݐ��c��{	%rBvm8n^ �
F�(s��t:�K��O�^�aү�B������=��a�dlR,�`���[(  ��\���k�hb�fU}U�;���p"���p��vy���w��~� ~�&�~ �j�E��i
��#�WQ� q��T:Nݦ�������I9?{b�6����ۯz�6~�6�hY���C�8�~_ ]��=�o����d��l~�	B5�6�����`2����٩�-��8��4~�kɊ�&���c��_�\���@�zl:Yg\L�}�$+�;�T3��Dþ��k+����]b#�93����h3��Dt�qu�P@����;N��]���+B�25e��̩�܄(,4�p�Bʱ\�̟E�wj�+�hL:��o�)���9 ��	4�ڗ6N�����4��*�_>�ҫD����5t-Ȇ�!��,B���V8�B�7�yyS�f�����L!׏���6�Qm@d���a�@}�W�쌸�f�)]Y��|��8B>���*�?-�EG�S:jx�8����g�k<��N��Ʉ�h����΂���zXq�@�������)x(����C�O'��U���\��|�y"�8�O�z�u��ݦ�@�/f6QN�S������ƌNPM��������dL�0_�\�E�^��,a$���8���I�f�=sc�.�z/�@����꺺��뛩Tu�ZGU�H����);:�]��ˌ����R���O_��5b���c��ʏLc(l�h���&�F�����G��¯M ��������LT`+���Tzo�@#�#)(��u�h���g�\Z���I����z���r,Wsum����lE?�z 
��j���30]Ef"� ^�uP�����V��g- dk4����`QP�e�a�3�:¹Kr�[=~�I��W�GdM����A�&N��(��E�k��J&/}��j��|�J*E�1��C���x��e��r��?՚�.�*��rJ��W�`͝:H�I�z_�v��eC�V�,�W�9�lF=�������Wo'��z+�/�K%2���&�@HͿփ���M�R;Enq��n"���o��}��Em"|�pq�S��\��6M�+y����>P�)
��(�y|)r���|1�~I�o҄�kؗ������AL��7o�9���@�M�~��7��P���ݶ�(T�75>��V^jиR^�nc����*�ܼ�<6=���z��� �'��C���.�u�s�S8h��I������so�X/����Nbc��V=�j��x@M�΅_�Bw��h����E>����Cʩ�N�{Y�S'1�s�	��������<u�!3�7���� H!L��� �XX j�Q��As��f�]>Z��-��R�r���7I����0ֆ�ÈaH��Cc�j$�g�y|��c���-=k����m@�A�?�];�L���c�p��<,n�`LD����4%���@��{v:Ȝ(7h��tQL������l��RK�m8�]�C�1%�k��%
0e��_����0ko(�n�Ӝ�g�L����;w�GtT>���/eõ�a[�OX����V"n���)�y��k �Xr�(��]��aމ�qćyÎeY���ת�a:��4����V}��+)���ظ�ok�п ��=�7�Qq�����,$�tx�%5Yn��a1���N���������y?/xWW���$k�C����5C�vჿ'����8d��d��k�_y���q������)�K�Lq]<�'�&�:O�pm6�_W�5�1�'ضV�&���%��R`�TW7�pTHE�݊GG�hO�/M���]�����ͬ�)�TE(Π��&���������W3���T5����!�f���y���	[Z��w�B^=@`�!���_;�S	�^7�7Q�)Q�لt���x���I[`F���8` ����Y ��c ���neL$�9X��u���,������p��?R8���S�UD�D-{y_9:{zL�t-��Z��o|*E{�e���ceI��jn�	���9�����`}Y/4d�� �4k�����-���ܬzBo��g�����2�=�z��G��O�vAa˙��%���+d����D6Ɏ��o�g��9?A?�7���
ū`߄P8�b�`6eo�w*��I˕�0��^+��\��
G��~t���,~P�"��Љ�B�x�w����ޅ1ڬu���Ú�l���T�s#Ɍ�dC���'���o�b>^�3��%��b���e�r��;��7��(Yl5]!a�'���$�pō�ڙR��27�d���Ph��`Hv.����bR64���//��K�[����t�	t����cM�>�u�+��Q�
1���Y9w��My�Ԏ#���9\gFld^�� `��|Qd�����}�q|a�<b�GO5 �ɷ]�d�j��H���
���e�� �}�xja�_zHwB�,ߌ�D�ׇ�����/��r.]��c�)�J��G�A,Hl�TC�q`�k=O�ʴ_���? .#h/������ Z_+	R�ֆe���{��F��z�]�!�� ��Kc]O�_�=caM�Y����}��sU2)	�,�h���	u�#�b��)T6�ظD��B�B�oN��ZDj�+~�r�v����H��=�� ``G�,$���䯪�
�N����ֲ`����3����N��l��I4�"�t����gX��&Vm=���O�%6Ɯ�X�����vmj?adƷ#,����gg�uO$��Q����D:u��l�U>�{}vTj�Q�.�ѳ��y�SuA�)O�R���MTh�Ʃ��AmG��Dd40?���t���m�717 �y��Ӥ����<Ѩ჎ƭ��s�J>>�]�iq����NG��\_�2����ٖ�:�R	�M_�aV%B��R���jn\�L�8�Ց�%�4�&K��a H�7�餾�fdw�J��&&#����	�Y���j�QϮO�"w0��P�n�>6�g#X�Q�����Q`����e���'�Cs�v8���O�(�u�i�=SNG�/�@G�),{��"��ȥLX��@�z��W����y����$t���,�x��=��հ�;���p�f�M����5o����#��+U���+-U`�tA�zzd�m�X$����*gq����p-,�\����xo^��^���IJ�����)ѐOI� �e�+�liS�ُ�2萦uK0/)��)b�]���$r�e]|�V��0��D��9�,��"+�w�C�t��_����#�����FkV�� p�#}٨b�K�۹6��f�`d<^8�x�e,ڤ���h:Т$rQ6�8����2�J\vZR&׮*s���wſ�wK�����e~'J��Xb����>_��Ӏ�����|pW>���#�i�W�)n3-#��� 5�:��-����Z��5����B�;�؜�ASic����d,R��/������3��v���ݍ�t������Ȓ/��*p�w4��+v����[~��!���ԑ+��[�&�/ƣ�(�o��o���<s��{+J���"�Yգ$�N2,��T�$����5��-w��\A|��^�frQ��9N��}%7��6;^�+���$r�q :O	��;%���+�w���+86��!l�+KZ���b7f`Vﺢ����{�FN�%�������G��;�]��|��`�4@?#y5m�����vNI|��,�qwF�_V\ ������ۨ\�ƨ��{��a�8�lV>��o�*8������5a8�0H�$�5�>��W�wDSl1�mE{Tt|2��!�v�h�p�O�l wYA�����Yv�����UD+Ԓ�`�/������}C\"��1�,�u6�(�e����qI�#B��]������0?�[���Gz��Z���sX���2��a��#�*�e)�ǯ�*���Ki+ѕ�OnV&��Ֆʍs�쇌�ϲ�k"(UG@��5�pXt+TD����g*��i�~u�,m>���XQ���;h�sބ��Vk�p��r
��-��h���-����d�=�F|n���ujd�m:�""'�ȫɨ��c���#��]AX|{�\)�;g����3:�>�]-y!��ۋ�NH��=�� �J՟�|���
�]�Z���cx�ȳ�'j[��u͐ŋ�[2H�7��B��������8��Z�Iк̺)����آ��z-��z)���K[d�� I�y�������c./�U,�r�n���Z��Ϝ�M�I����������;�JLi�wu�[��J$�Q��/���� �^�[�L���Z�Pq�}�c��2�F�A��8��ȅ���tLe�3�i�����F��+,������[���'V�i�0�_�{i=������Vt��y���k���M� ��⡃)��q��-Kao��	��3V!�-�l�������1��u.�l��l`i=|�C�Yc�Cy����V���]������.��.Y���B�y�#��x_.�=�lL%:��sF|)Ղz>H����qc�����H��E�ݯ �p0��9�,G/��?�v>,_�G�~Uux-5�ם��O��n.j,!�7�x�h������$�B��ʹQ_0��}��˟�����Mn���d?���nP��*s@������_</#��U���vvI7ܐ��m��O?!�I{
�����P�����W�4�x'�����=���%��y�f*�F�mG��bf~̢�wٶ�����(r*����X �M�[�;5!'��a����Y.��?���pm�W������g�`ay�%5�w�#t�F��8�֦�\[�ŉ6�|���wY�%X	Q&�fOKf��0��)�]�R�k)BR�HZ9�g��$G����0dzEu� ���=O�?��Ԙ�U�����CT�l9X�0\�H$�����>��M�6�'TLk���b<�s��yk�ܵXKr�|b{��DU4�,Ι����|�z��{Ê�E�l9���%B�|�/O�_a�%����!U���O:� @�s
>}����>��Jo��+"�s�w[�f\Y�2�P�t���'G왕�"�M� �����z�壀��r�
ۗ�L
�3���I�g0�!~��ye���]f�4Y�ܳś����ɽn酧-Z9���,������>�e���ql�g�+	�͈�'�Y���p�(��P
/�cڨ1m��ZU��>����x�4.w����
=�1C�͊x�V�hձ�����ܪ�R����;oy &j�}4��K͞>���*����o媾��g�M0��`wI=�f�t���`5�OZ�W�3E�xx����f��@�!���-���8�������EA"�(��y�����lP�2QD�%=�jG��)���7\�2�oV�A �<�r>�]�J^ɂ�;�B�q{���q����H�5�tAZ+��&�Q �����ar)I���O>�<d���4��"�]'���C,a[�!Y�~&��?�X��m�[yK�W2{��皃�L���h�<�˻I�މRѠ� �C��U���_�[��V@�2Q��K@<�����Gp�W���a��Y 0Y
��,`P���)_��|j	��>�j��PM��lЖ�5X�B�>#�8[ٮ~+ĳX<�v:�a��V=p=Ի i�C7�ٲ�	h#��RA�
��_�	a����smۏ�> ���v�ˑ��ebQ�? 4��s�mc�G14?-�>�sj�ϔlW����(e����N��}B�c�I���@�G��O���l9��%$R��/�8����j����t#��cx���`eȼ�G�M���OŊ#��B�{!醒�����m�¬yV�)M��n:�=K�AꑍE����ze��w��Ԉ�(<��۫À���,�u8�V1hG����߉	��7l)Ӌ����=Z�t
����o"�Yžd㐄��H.休�7#�f"U�cO�!1J��sҭ���B�@�P�K�.z\�?o�}+H�3ݑ���O$pe2L.�$�<��>��Fv�:�n��N�m��Z�騫�i��PeUX#t!B�~�Z�Vo:�\/�6�]��Y�@�.��1SP�~ ��>�{`��~Y�o��Ύ�K@�rfG��gg���E*6�Q���\���3���7BVX�o< �@���}��qy<�-�_bTS�H�g��]IU&�=5ڌ�3.�e�`�6އ� >> ��Xf܏E��.��8��~z�G����!<rx?b�^U�6�1���sg!�"��	�b�>-"���Dpհ�S����MN�3{��0H)�Tt�IXn�ww��-6�DG�����$6���l�Q�۴'�!���3����QE �Ws���5��X$6�
Fg�����A	"�u���Q�qL�>ů@���$�u�*$�����
'�	� ; �aw<7A��E���,�k�RU�}D��Ʒ,�T�K1	)��t��8Ҽ��<YLc��0�[�<T�}|C���H/��f��:�r�!XbX!3	q!F�<�����6���`��ڹ24��'ծ��ٺ��s�}�Üi�0��z�y֏q�>cM��O���
b@���C��D�j�W��Mz������z��a�FN[-A��T� u��n��3O��,���b�RŒ��F2r�YLdr�k��J(�lXufp���U Hב4ʶE�qcA��:?ⳉ�u���-(�݋!�vnˊTekR]U����4|ل	+
�]|vn e��𥬤��P�x��-Y����U��0�E��%�����<*
+�Bbr���$�옼D�OS`f�3�5ʫ�a�'�sI��ʹ~>@��J{�.�t2�3 Y�%�~Al+�;������U�sE4�3pRJ���HR�w�s�Q���1�%�T-�~�;�zxn�c�7|��%�5������W�/�{�xmڎ�[�-S&�|� C&� wCSǦ�hX����Y��iZ��6��31W��*��2�N�il�{Z���a�.r�������n$����nom��gr��76���9��8*ml�v�����-����8�`��ٲ�d�	�V�[�tv:��VYL�ł���d�r��a";dl�،p�G(=~D_w��c+�j��b*���֡�~k���/i���;H5]��|ݛ���fٙ讠�|^Re�F�N�����H���A��;p��c:���aE�)�7���H��z�7��Acjt#��oNc�(cH�<+2K���!g8K�'3���+ν�,��M4I'SP�b�ɶ�}YwҜt�rXr����D�Z����V�?#�0��}>N	�J��X��Q�>�1h��7���e�c�o�[:h�?�Ke���F�C��,a*G��T��f�Z���~���=s��D$ϗr%��!���aA>����'��I�Z�Z�@Y�7ҁpb^�e7ɓI�;>ԟ3s�j��靾�v�EY�F�ۚb��K(��>��K�и=���9{�g��k�������kڒ���8Χ#��`�X;Ɓ�%f��mz��y|}��Cx]Ӹ72�I��m��}>�
�����(Ĥ@Q6w_�e�T�r3�A���)Za�!�"Ƃ#�mغ�����Q4�/����o�_�-j��gO=S��TB�#��I�Ȳ�0,Ǿ+L p�R��#��Ѧ^� ����o��n	�z�0�vҗE�D̛k��;n���2Q<nsD�)�ڂ-'G����`t��V˃Y��3l�zR#��7�٩����6џϙ�V��*��{E*�{Z:XX�@�C��(�'���Z�X`;Na�<Ģ���m�O�K{D��ɵT�TN"���[�j0�;t4BL�e����u�#G!^Tȗ�j:0��K�ٹj��Cp�u���9B��R�ų0g�
P���N��C��7���W��O�A�b�'��'k�0�3Hڳ��-�{��2��� �Z²��1�A��;<�,��习�o��2�6�9��p]��Ѡ��n?i�u�������@�����?ޒ���&8K����i��!m^"]���r{�B�$�y	�VH\)���"|���^�ױ���¨��M���
����Wo�hv�^�ˌ'ڟ�]d���1`d3���ܯ*���8YK}�5�XAQkF��rM	�U=�����2?��pv����gdq��Sm	��)/H��y�dN�E��C�bRq�|n��P�L���S�i|h��Y��|Ĵw�W;�ʓ�d����ȯv��/�0��Aގ;2]��R=u�ޥ�
��� �j���
�orn�b�	<g̻-��bk9onh���7N1�$��1�ܑ�����uH�'P]Ƚ��h��7ӎ��a.q��┕%u��"�KeUn�����V�}Ām��u|E�@�+Ƕ����r�`�A���6֣N����S�m?۾Z���θ�Q�����Fz��o���3�����*w�*=�Ǻo�'Xv1�7�Lʟa ��1=��g�n&Ǜ�4c��>��[�t:*���=�9��T(�5�/[%7@��_�3 �V�,�B�A�#�XÛ������I]�&���G"$P�9g�c�>Zb_F�m�dj�]VI��=T��|w�������;���3#��x�t2c�`~�GqbȪާ>g�!���sd����\��4P�Ir-��)T/z�y����Z=��1P?T�S�t�lp��G�%��b�� ���7��1Pig;3�q�gZ��gD�,�R���N]�K�+]�[�16`!�;̃��2Zz�h�a��*�׫�� �X���#rr�G�@g淈%4 ���G�	��[X?h]�ٓ�r���bv��ӂ�*���<C�����d^v����d��y1���~k�P]��g�&���tq�VtLg���x~'wԖ�0�NI�Q�0�؄Wb	�X���L�4{q����k�XŬ����]ZUK�EZ2��.3ΐ�7t���Ě��Ԩ�K�˳�į�7�iP%��P���1tL��o��-����:����Su[C� Gp]���H��ur(2�I~��
O�L/_�y�T'r>ٚ' `<�2�y��9H\Jd!�F����U����SA��8M��mpp�q��D�@�wW��	}38�m�w���)�8.��Ic4�	[�X�V� ����e�����T��{��	A9Ɇ�p�󃿆*�VI�汦'�)��*C�s���e���l>/���H�9��y��� �/��{�(L�J{������PWU� p�̓~�ֶ�业g�zS�į���5�P�`|� o�xFAr��9�>ф�{�]V�ƅ�c���z�n;5 @4�2]M\��#�b3
�� ��]X](����7�kE��O��0�u�{/�rs��4a�Zh0��Hs��3�'f�˘
6����۷�ݱ�=x��xm�Sz�2*l6��x�>�T���CP|H�;�?��򴳯���&�6J:�=q�T��ɛߍm$��{�~��W�0^]��bJ��;�)V>�5�{>�#Dس���?XQ����^�M]S�4��l�������M���JO�i��?��+:7���,?˫D>_\`߯��!�x�V�/���mcvL6�M�NS�A�o�X�٩�4
ϊ�@`a��x��d�����LW4@��CZ�����Y��fGŅ���;%��§�Z�f7b7���ߜy/�E~���a3���������vo׈��˰�m�|B�#���{�Aj�0��#	%yl���X=)�����
K6��9���%"��뀰y����?�X��0�i�wap� <,+�hwFs��;/�А
S+cߏ���/�"��jN �[p��sRM��I��3(`@͍T������`���P�O|s��@2��5����=�@Ҡ��WA���+��S'���Ɇu�)ޯ�F:�}����98��~B#�a�գ��?/�1��]ĩ�bH�$&��P�(g|(
�fM7�A��!Bw�}LQ�Y�-1���,X��y�Di��%�L���CT�gIDG�����*� q�d�'K�~Q�Q �䔾��zƣ��rŖg���a6t��x+�ߒO(��4�TwP���Z��C��jl~�� �VX���W��y�m&�������^Nua��C�2s�S�����Ä�J甄}hV�K<p\��U8�H�ԛ^ �
��h6?	�V���@α[ߎ���:���W����a�(��i�*��a{��]�� �o�%I+���ӆ�O�hw���=8M����:݊�_��5��/mW�-�}~�q3�6�˾h�^
��X:_A<-�5�yӓ-sgA%��ܮvq"�����!�����:61������V�z�	m
�m���T��*�o��g�p��aA�"n��
zn���Ȳ� �R��� N緓OL������F�ɾ�R��Y�-!:x3˥dGIPM�~^E�C�L!/V�v�������aD��7��P���I/Q�N�:�̌x��e``QS�#Wz	�x�}�tn��,WL�����JK�j�����(
<^w#��(��Q�Do!t�%�nț�?R�&a.g3*����Ax�w�I�����C٩��,v�K�ua!X�\
w~��#<���e��o�[_zM�����\ڹ�w�7�7x�ٳ-q8� y�4SM����W/x��o�������d
�H����lp�8af�.Jgs3ey"�P�(��@=��G��ģ\�������!�O�@v5dGDj��=�����c�����HD.��)�e5!�5��>�i��i&�<�"��Q�?�?H�ʿ+ڜ��z �S�6 ��ن�H��=�)�&���?Ԝ�B:�߁�k����a�]���5�&�I�щL��ы��e��
�d*⯥��W+~C(vb��h���g�+�h�Eg�j��ƽ������z:�*�	�S�̜h4oЀ�i()���YF�O��k����y���&~x��)��o���Zj6�WjN�F�!��r���S��F��ap���|�N��U���	~6)�F���0=(�O-�Q��FM�����D4�$��I�G���H�m��Y�P�Д�RH##���4H����P��+�c�f��b=��_D)����3��W�ܻs�н��1LN滹o��z��2�?˶����՜�]䩺���H�d���kX���.Y�g��Cl��H� �NvG@b��c�R?��v�nSC\(�$��~xb���a�*[�#Tͼ���$�Un�c�0��ɒe-���B7�GWC�Ń0��ӭ0�1wP{ʌ]�_X9�'cu,�i)�͵�2�[�k���#��xHqaM��qI@�pF�X�D��[��SV�)ɻ�:Gۦ�&<��(	:�Aӥ+�6'3g�)о�#���']���J!z#��!phH��|[!�k���ۛ&Bۉ�P��h���arh�Y:3���S������ih��g�0���M�p8��_�O��V#k��;-��";4�*�&�x��n���zm곓�����H���
���v�G����16�����5Y��?i����z�)�������xc\ew5������d��|�llS��U̾�r����&�������bQ��C#�E:�rVi�����Ú�e[�޿ �\V;J�)U���M0�nzZ�`Y���ã\�d�L
 �o��.�R��T�gEQ�|R6�5�2R?	z���%���_��
�=1���[��H����L���_�1u�
D����7�TK\�s(�9����mO�ma&8F\o��? �1�����%B��[?�Bm�Tf�=Z��'�.�4�N�1�$�a`�NУS@)���n��Pd�ͰL���K�ç�)^��B���3�.�.�����'�u�`ľG/�X}f�&�,��&�U�RF������*{$3ޯ����wwp�]C��m�QF�̊��AP#L�p~���.�#f^�g�,::>� "EpM�0@/�
��_ݛ�o3Uƭ�o��EY���v����� ��ĵ{�~!�����В�)Kq<�{F ح䳾�y~nN�y�I����ǜ���A����@�Sx�y�1����E�3ҍ{a<e��:�ж��o:Nڍ���:�JcB��:M
�[���KX���k���#�����\V�V ��Q�]i��i$6�m�+Ëj| @ G��ް2�&j�c(6q��C�5��e\�k��ss�V�4$�[z'����R�F�������{	�X#c6G0�1�:��3���ˢ����_���|-Yq:\=����n��� ���
[Q[�o���WpV��1^��~���4����9�G���"Պ�;	�  �in�<9w��!S�G\�wXxd��B�@$��}�6�}��E>p��6d8���X甾��wZ:����.�-��q� �Cຒ�7<�$�*,up3�#8Ãy߀�|&���:��&�v���%�J�F��6n?"�.�i�G5�ͱ|��e��o��Ȣw��n�?BƜ0�^R�����7��	;���@#{��\�_5L���|W1�l�Q8��(���Y��]2�=	�i!_In-&
��9�J��+����qM :L���8�'� ��m�C�Q����y�7ʬ���*�<��/o�ʪ�v=7��'�5�@�oV�1��Ǣ�sY�I�L��;(nQ�׬�!Fs���@j���N�v�p^�b!�N6S5����c����B��7��}GI�\������"�ҟ�}�H�*�_=�8��ZDN�L)��׈�Zo�
��v\o��2�\��|���K	��!�=�+�S����=� 
-�<��/�s��x���d���4���<�&5��a���(�o��wC�\�|���,A�tfH^��P���QZ�jy��I^&sD�
D���
��@�T%��U艢��x��6XZ��`�����qy��MT<����U���[��Q���3� h�~4�}z��~h�F�t�!y.�`�1i#�K2�U=)��&�����X$;̸&u���ֆO� =]���X��(�Ȃ{����� �gtx�X3,Y`���4��b0��0��M�VY���/1x��n��:�;�_�����ej����꜈����G�ƥ�%Ag������]X��+s�ګ���,��'^��G�*o���a>�|�K�:�\*aX�w�e�0�|z����
+e?]�a4)2�	�	����`�;Z��P�´&*Q%�=�^�&_@R>��L�D΋�QD�K: �#E���S�I��&�����w��7��vzS�'s���1bE$�q������S�0�lN�}�o[�-�.
���y�'(�\�Z\�-#��f�uXe5m�S�S�����yu���A�Cl��ǥ͇$�dMу$��s��b��խ"�=� �'t�B'H���Hd�s���B��~�;�X;G����$�g�Q�)N^�F��T,.��E㼆��-�:̕1�ɱ�6bսg$�e򎕍w�*���5T��mN��Ӫ�<��U�?,ȸ;��:��m:��4.�_%��?���f��e��~����g9��eJƾ(bi��1����c� P2z��[��ܳ�V�#x]�9�֧UN/���$<3mD�$�'�s͔��^R&_���S�.�@�l���\��:�RFS�>M�j��G�0ik�����dՂ;S(��˶�Ω?��!#?qzr��9�F o�`Q�h�hz|)�53apn(�$�w
zW�F0Uð�"��*�Ȩ��پ�[]�3���S���!�$���a���Mv�	qcl�?�t<̱��~1�\�a�~���j�.h2��.O���+�ݔ.!A�-&;�� -�aX�m!R���:g,���y��aI�2v�>��\��7ճ�Ne��51��Z�ӌ���6p_�-������p�#<�6s���VʨH�?�(�[�
�3Bu��@�u�Ù��X�G$���-FL�# ��ÿ��f䢊X��ؠ{��2����b��fC����X��A������6�,}�Rz�a_�!� ��R8�h����$��e�|�,�כ�w������~�p:n���ƣ��$K�8��]q!k�<��yQ!�C�b)C8�S#�\�Z�q����QMi����x�L�gmR	x�Ŝa���8|��t��/��]Wx���l��b�D<��~�>���_$�����I���<,�;������ڷ	���Mњ��Hr��Jv��^zO�L���#��qB��/� �IŃ����}�޻*3-CK�K���o#{Q��)[�Ȋ^�@�1��OY����V����=�Pt ��`�gCѸ���x]2�Z%:���uo�A$Կ���}`�Y��8����E"OG��Ui��<���T�
4�߳&�Nd���Ti`:u��MvW���N}|s�,tl [) /����Ÿsm�v;��ЊHӈ��g퐝;�!���.��K��	��<hbw�F,/��@6Mt��82O�p$䠙ݪaO�N��u;☽'n �"�~�U�eQu���7���o���^4x����h8��t"Y��1�7�2m���g��Y�-�1�B��
�Z���F��H����gm��y�,�(^��;��'"�;2�jzJ����&�i�����M�^� .n\z@��M�4e���R�t��2��{�����_��`4�'��n�&{��=B�ns�&ӝ�E/6�����ȳ�(K�i~N���K�!��7��:i&g�ĠK�����&�	���D�a-c,�aB�c�GPqi�\��!P���'�mp���P(�#�!�s7"ך4����_���`R���Z>1�F�s�k��M�s��Fۿ	y��鯓�C�j�t~XS��y��d�s����q�]���kr������Ed�_���r�{������׮Ȏ�[�	I�]�;g�]�/�91�}�trg����Y�cG��k� 6]����S��J���8�P�h�Dm*,���pzϋڎQ,ًt�P�Q;���Llv�V2=�#��ܐ��G�d.���S6h:m�BF[��QXX�K|4ˢ$�Dϝ*�#X�t���S�ˢ�١�u(eޱbဦzht	Yy�=���?�t9Ba�L,T|M�a����E���ӣo��%NL����HP��V�vRo�g2T1��5�)ʩ�*f�O����Q���9!��4B
yd��R�>��YZ��Ig��(t��$&-�҃"�=���<$�R�Gw�t�V�J�,�����ZO6�gJ���)�"Z�}��eIgQճ��b��4�T�lA��Qp9J���J��$1�'������|�J���P�s~����_���%Mw��5��?R@=�t�(���%��\��P6�J�ĮA]�1��H���l�B�ŭߏ��S�ɒ��#a%�����\��~�XK��}��7��>�ޮ�%���D�yㆵ#ы�:l~�SeR�;5�B�~��2Bx���6�K$���x�&�c�B�nk�Y�����6��*�n��O�{Z��߫�_�xF��)b?aN�}J�.d����b������V���3L\��{Qps�H��@�	N�����k�2����2���:p1ְ�}��j�Y�Q�^ V���fp�R����	�Q�Cyq\�T�P��wh"4��n�B�|��"l���l��pp�����
~�G�!��8��@G�=Rt�G��}�j�L^-SQ�D����3۽�P�c6^f��|Kz8x7��c"�,�3K�C^ԁ����g6�xAh���Zǿ���B�"~Y��t嶽l����<��&X�Twl��:�|��A}�7�F��?T	%�~ aݕ�k/���0s�!CX�A
R��q��9���/��5�v��]�S"�D9jM|y�����h����R�j0Bh|W���������0Q)�ވ9�6k�� (V4[��R��@��g��q�$�̯븴;��N���X=ͱ��o%��<�$!p	y���ls&
�.���3�2m���DUR]�o��5���杵Д���v��i离�%H�t��k���Im[7CwH���k��:��vm.S�X���:@q���9�zj�h�7����xxl�h��d*�󪟽����ˈN|� �W���j�
+hU��ה��lZ|Uql��b���(��:�=)�ˠn�v����g.�uZaq�b����W]�l{R��;�GӿSALh��Ћ�/(��mL�<zr ���3n��T��$7)�����ǆ��9�TP��ܰ�#GS���� 	(C�k�_���h�4J��t��!x9~�R	 �8��O�t�#.���l���6�6d��2dB�Uj�8�V���-��Z���ڵ25�v<kf�aM,B��3mF������]A`�*/��Rh�Wm�C(pm9p�u���5|�R�י����5��I��D4��7`�~�Ӱ�}��1tw�X�plp�V�1�5Bc�=~��HI�URGu�~���5�0���'��I�� ]�+]�θBE�a�eݥX�C��a76	M�h�M�̥b�<�����,�$≬(��*��0�+��R\Ƅ����8׶��tAم��O�pf{v+��6ʖ�i_�[}=:1��V�^�?8��d�nj$7!OTY�W(�p�#+�@���oc��5YЊ��d�X<��
�6��/���{v�g��uEW������T��j�+��ٔ�b����"��D[�m�)��5&x�H����X.����c5������R߰�UcQ�Y�8�g�����qq���;ihV�q�Z�!H����8��8�Ƞ�n�:�BuXf�4��}�'��u����e�q(9�<~�t-j��#Y���L0F#�/
�����
�<��L��a���i���0�t�kȑ��`��xhԏ&�����Ex�'�j' �!����Q�c@{�m�n0�v�����8�}CL�{}�%܍��a���i9\�DB#A[-���k��3�T#m.�|LG7��r=mIl24�ڛ�/u���� 	�V��d��]���t�n���r� *Xv���>�?�J=`>�$��+�c��lż/;=u�BA�ZV�H�g�1'���U�}�a� �����G�����.�	w��	k)�uT�I���!�A�(������D4-�_�SD�Ĩ��Б��Z�k�����I�+WHH3>�R�[$�[G�?#T ��t�� ���g�Y̮k���nՂ:���f���QE������r�q]7'n:W��bW�$���hcz䣚��z
���)?�oR>]bSE���ݹ��=��1^�h��+��w3��2Vg�R�o[?���Y��w�SWW?��������(�T/�]���<��y3F�?��e3`S*OY���8́��
e��=�|���)p�S�:�=��J�?�UUK[\�wv�u��6]�J�d�opݩI�jĝL�����6���S2�a����H�YI�fSc�S������û!9���PJc˶{�V��ZT09������ᝋ�-����K��&����`����L����T��_ _5��y@N� �)w~T.�K�Ҷ�i���cn��(Y�VD1]@��_�� "h>(J�X������'�/ ���d)�imr���43�T#Υ�	{O<��~���1���HeFǤ��צ�wU?'�u�����2<�UUm��x����3�Cޏ^3�y�"�m��K�_���^�5���N,)��5Pǔh^?��95%���n��y���Khj"w��i�-�Kģ�e��|h��VoWD��'�����}��ܸ� E���쎁���k�n=�lDg}����m;7O�`P�J���([%�8D���,�(�4��)���ap ��RW�~����Y�_l�вE�L�_��&�	ĥc�H޵������
5�1���/tcxP������R��l�����͝T�}�d�`�TC1�z8�N+z&��˨5��T�=m����"��8�E�� ��T+�h��@��A�F��eA),Ǡ`�mYX��.+��|�.�p�"��	�"ԙ&����q#S�X\��L98m^��)��l��+����)zz`�j���C5���`֤	���%и[��U{����<^r�u��6�T�y��z��: Na$}ܹU�wa3�\А��cE4��+�zb�r �:<b����b�1ŵ�3�Z�ܿrٹ����6s՞��}]z�Բ*O�vҗ�s�&��Q�#2m
�H�	 ̇迯��{meD�H�L_r�$>�a+�]
_	���Ui�n���ۻ�N�H�.H�Ȟ�7[o�/��\�ը���V��o�kF�d ��4������R�/h�(\ޟ��N��o��:��Ţ�)_���-o$��>�G��<U͙�y�������F\���=��O�y�!�ꖒ�?�����}ъ��m��/����	q9���tG�M�I����M�D�I�nN4�s����%@�������,!f���n!L������Ί��'"�F ��p���$̔W�ι�*`��#Л��q\�(Z�A:���m��J]hU�k7
�t0�e���x���H��K�݃>)6��J�m I�J�mx�������l�f�/o�P$<#o
�G�=�1����ns��D^SD�@}܎%�������6	���ʟQ&r�@
�o�R´3ƛj��ZUv|�6?�O�Bnd|U�����z/�B��D	�y��!)'�w6�SU
d�F�>�� ��
K�=������ΐ��S8��* E��%g] :�C]�PWj��+P���='�_N��\��x� �p9{y0��-��zKm^������7�Õ���~�e�v�.�Q�\=T���$�Y)��'��V��ə�\��񢍰�Яtq<���E����o&��3���E}qf���Z�+f[����EuGDe6Q��Z��9ms�7�b}��z�J��t��&Va1��ύ��Ǵ���n�Xp-�\���㉥��WU\��h�h�<��s�B��Y���><��s-�z�B?Q����/��
�J�c�m �9 ag&brJ^uf��2�s�c��h�Y!Sk� ��zm�2ֲ�����H�G�d�\��-@��i��;�kp�{8q�5��F�K=;����\0U��[��^s�#J��0V-���8�Y���D�:�!��Gy�����f�7Ĉ��C���}6�P|��^kMY�2�/�qr��p��?3ɋfk_6���N�n��ȗ"s���*�s�5�c�ˬ� A6�kJ�v
�$��J��x�M\47������ꨣ��i��n��ǵ�&�C�VE�\&�,��2v���7�{��l�&^G��L���=�����-fVp~���w��t|.q&*��ڠ�Fx@��}��偮W���_XhR/p���<k�$��Rm�'���8[n���,&�q��,�#������2Y��
�L���R��"]Ȉ��uUv�رmrfyu�)4!�|����ʡ;s�'-���t��;]TK\%]�M�:Z�I���M��hh8O���OZ���;�y�`Kx	�`J�!r�	.%dݬ2=������\��.�ӳ�%T�g�&�	U{ط����C;�{pVˆs��b�쁠����!�Q��IC����9�It���q��%V��D�-���|GS'S�4�
4O.���7f�C�[j�&�Wf��%�jܘn]�wV�/G��OG�y�a�s��D%��`ӣ�6W�K�րd�ֵ���o޿;���i�	gJc`h2�
�h��U�����i,&{���wy�8h�������"RR��n���$�͒�1Q�#�{�uSY˃S�{���q�e�Jo�8a���pu��lk9��d#�W�	�B��h�sn�g��hp��������n�Aa�3]"�4�;O(jB��3��?Ovqn6�,��dEJ�����I���ژA�9C�����3��Wsv�$h����
�� �?��Z��I���A0[��� �8�o�F;M������7�hy-c|x�q�e��:��^� ���c_�H_{9�)*?6��?L����Ӣ!&�N��m�Ny=��� >�X&2�X	v���5R�u~�6��vS�S�op�,%?C�����J?�>�̄��رO��Ώ:�����H1��0�K�k�9Nhq� �I7��و2Jj��JY^��}��\d��B�������$=�N�����B�-w�>c3_с�l�M�]��-WV�v��|�ȵO� !0n���	���Z=g��<s��EQ[Z�/�(	���1�Y&����g�����eS�N���ؠ�UC�Z������D@'XޚN*������Ų��#�Q�-��Ɂ5���������� y���Kc$���fiL%hI��a�ӾV)�|SI�.`�����#qnu�e)�-7.�8
�>(.m��FIG�R.�i/��<(N��z��f��԰o�q`B���&��P�|�=�'���13�'�84������{=1�e�e�<蠒�u�Ad��\�1����ٓ��L���9IH��6'vRPUIy��|Sl��?���6OA�ǒ����w��a0�?ҽO��(u%��ИF�Ⱦ#c_��w�J�[���@�j���j�Ut�iF�ȁd���[J����*�T�1�spCEZ�1���0LD�5�T��M#�Wk��ȫ�@i�VI:P[�g(;�/�$/_���.��S8������ڎ���M��)U��Ũ��e����d�T����:����{���J6�@kH��.��B�:�`(BP���� ;_�0��N�:4��z|HQRG�K������,%�@�K�ڦ��~�ep�޹1�Vb����˗�㥴ӓI�z�7г����?F�U3�f�v a�	�	��R�����Yd����:�����	���M�!=��"[����z���;� 4�����8.�p���mgRZ�)qc������t��+\���-��`�zY<��u���/���[떦� �ܯ�pP�Zz����_��V�J<��x�����Hwa������S���4� ��m��_勩�I�vh���LE��Z�V�:���<5wڿ#Xr���#���K�憋�[��{����A��b}
,)]ky�g�w;2%��0���v�1�ǿ_B&P��G�ZP�yB��B>��CS��ښؠ�H��w@����.8c�LIjG�tLӿZNǳf���y:0�b~����v�7�ɤ���as�4���?���N�� �Q۱hẽ�=]um e�]uH��|��0 �4�<���C���8�)�� ^�|wფ�#5C]�&�&��78Q��������'%Ɯ�{@��(�W�Þ4tr�*�9'hG�Gid|�+'�{C��0�H���q�}u�~�h35�38js��Q��gNͭb�w���������κ�CC� �d/�]��'��
Wt.`�����]W?c�∏ӫ��Z���ݦ0fCUk�]�����x� ��$j�b$�8�Z�2&5�����Q�m@�I�
`i�h>fCȔ���Y�[��s�]���`��x� h�W'7��q�qs�PS\�S��G]֘��Q�=o�*#����3�g������|2�ΦYllX����<h�C��2�n���@���@c!y	������-IN�����̏}���L��y�R(^z��`���,�������$��YNQ���5t��]�X
z2뼟
�*r�0��CHq�0�u�gdF�1'��2��+����ts.�P���N:�I���>̧6���0{�뒪i���#^���U�,�0�:I+:u)���M���"x��V��f�6����1܇Wj�G6+Fz$LnMR��s��GgL��xT���c������+��g:(��	:o�u�e��[���Yȕߑ~�r	Y�GVɬ�c�6t2K�d1��ܐ+�X��3-ɒ?��0BK�0�o���t|�P���Q��m����KN�讕�_��5̼��ܳ��Ԃ-A�������c�N!o惜i9�	Gœ���K�	�.�ޅH s��|��:.0}e#�Ӌ�wKKM'�����g�'Ag}��e]@Ŏ���qC}��Z�)\Gm�N�X�/e� }�����'�����k ǆw�j�m���nG��o=:y�͊Mx����<ĀLS�8K�'-�2ֳ��˱�_�2���7H��� "��LyX�Ͽ��2&�0�?��$��*e�J����tu`��LQR&:[���\b,��әp�0�"���s�P"l��)Mͯ���;��W���X�������Y�Ӆ޾�w�\Y2v�DjJ�R�Ja�t��n-s�@�'Լ���'8�m���Q)?< W�����t��	�u�cTo�%��N�ͪ�{���˱�y�L�;��4�P��(������1�uW4��*��Xix8i�2����F��K̊���������w�"�8)��E�N����~��/�Aө2_J�����u?Ե{��-B�u��G��7*ec�U�<�U\�k��0��V�색��Sy����6̅j���+ �n|��ֆ�f(��&u���!riX~[1 ���Sw�4@�1�����$�㫏>4Ѯ_��&_�f�t��D��o�E�"e1<��M5YEP]=@�i>_`��UO{��=	hM�O�Õ��0�z�Xzam1!e�=I!�6�#�t�b�4�k�[e�rp_%�U蟰U�Dl�Q߼���!���r�1���5
�}�V��l����N�.(�|�.��¢�x(hݸ��_~R�����SǊ����]~��[@�G��i�k�h���(iV!\�o$Ꮿ[q����\J�%+^�F�3����{�|�����γ3�AFǁeV	���kgJ�Dl*�����G��0�f�h�z��2�����ww(�u���ҽ�z&��	�0���y�e����z��h7�'�f�P;��o⍘���oͰ3�.��5�����lrt��#��IY{w���A=�7����ب
tSX��	��c��웕�|	 �Ķ�Է)~�ͮ���%*���G��
����� -j�M@���<mVd�b��آuD�����q�1�F�q�}=V|�Bf�2�.��7E�T��?*�����&=��ڥD�z����,�״��6�&�~��̼��#_�5y��sY��%��֔OC�G=��W=kğ?wu�t\�
��> ӑl\�񿤩���V#LIc��U��Bt����$w�x�dm��
�%�{�??��'���-�>�Lk�Հ�_3�0v�rBM	�y�B����W9�W�m7�&7E�@����6�4O$��ڌY���v}X�����CU�{�N��:���Cl��z��{%a�?ϱ?�h�����jcM�Ix��B�9ՇR����~���K��HTĀ�1���~�]K��H��t��'񵭖sοc��}��/.�_�s]� Q.�S�?5�gQ�(�o��}f�d��E����{�k��� qG̐(���G6���A%�K�ɶ��c&��ῧ��߾�S6�Q�n��6��kN�uctݧPq�愊�nB������k����)P����4"38�������WKv��1���.R{�"z�S�8	Q��q�
L�F��_��9��y�/KZ�g�G=��7`=�"� �#!Z.f�1:Q�f����X��uG������1�������`���;��x.)�x���F�R���41��K[����U���
M�'myՉ[/���iU�>9S~U�l�o���?��<+Y��ͷÉ�� %�S<Vg�w�o|cJ��`�T�m�J�Uo��h \h�*Gs<?DSB�O��}�MDHl_.��~���:J���7�dz�K!1k���Djf���C�D�x�{j��W1Y���	,p�|��kܷTNc0��V	�=y�ﰂ�_5C�]�yA
 �g��ݪ�5�-&�͆���(b�R�ҰB��'���Kc��Q�3�n�sh�e��t7`E�V{s�m�����B�g����@m�i~◟*_m^�_z��Q�S��).3�?��o�i�����"��Z.���x;�H�1r���Ų��Y�e��:�jZe5�`H�	�[��U۸d�����q�w�i�p�= "	#M�L7e��Oh�?ϖe���JL]b��C���"�1��]J8����%�\��_�б�����&�>4�h"��x�r��⧤���4vMKl�*�Q���3��l&:?Bj^v
���g�6n�G��\M�"��K�>4~��Dˋ�"��`2���u��5�+�q(Fh%yg�S��8�W�Gf}7 �A�f�Я�P���P5%�n����,�+�_����.Vmk�5� X=2i��Vn�GbQF}�a�������(���E��4��o�L43~W���f�cM'��OP�c�D��5�\؂ ��3��>}9���rtwz�F](=E_��
�[���%
%�3��jB��������Oc�HHk�ϰ��]�����}��1^_��������k8�~"袑^�,�z��:^���iVyf����}&cf��_,�������T���E�ɫ'r!h�6:.i؛b��Z|ǯ��������&w��S~��|���G�)B��C�ri"W���b�/V�.�<��9�Y�@���Z���k��0�$ޅO@��zD��ky�9$3�H�����ՙ'������"�{/�4���\��u�f���:���E��l�(��[�qQΏ��܆x��}QhcS.P�HM�����3���[�L֯�0��VA Z:�g