��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	��3�A�D��͡�k^�e�0棎,27��ttcqkqI}i!�0<fC�#� V�g�?������N�@�	��/��"^P���PIp��@ u�ҫn����g|�a�@��=BJ��S��d���\f:)����n�fJ�l�U	�'�L]0u&ձ&.�h�i��B9s#Q6~�����I�M�&7�;GZ|%/��輥"���!�A[�e���e��}�"%k
��~yؑ�f�RL�B���s3g�C��?�=��+�DO�u�M�6��%"M�d�N9��m����0�k:t'U��S�W�^�5g=.�3X��z�Ǌ�{ׄ&N6\|�	q�9�X{�ܘ��F�����)�"����FWa��&��ƴ��,z�Ә�����>1GU��� Q�m�!������bX	�����1-�]"Ki�;B���&o���>���c�8�E4P�����~���2Ny�ߑ�E+���z��2�d}I��X��V���-5����CG����<������n&_�L}�RtٷT:ϻ8�o;Ȥ��K�W��ޏ�X˷ž�i	呆��q��Z�x�<����p�T�g-y�^E�qQ����\!n����g|�)z��kW8 �p�h�Y<�C��?:ėW4��\ڴa@�~�Q������݄�KZu��8�.��{��B�\�4���m�K?	��̰>��[I7Uj��T1���0��
�BW^�C��J�N�,�ۥ*8�E���, ��e�o~է�tF@�nw����j��x��H�� ܴG�N�y�d�c���D$IL����ɍ��"�P9+ B��;����CW��*u���l�%bM8��;U]b��E��Oxnl|�j�����n�3�W:,��]��!8��N#����:��ԩ���|ǩ��#<���7���~�"�H�n=����Y��pk3sy-z��V��ò�:�t�"�U췜�>����A��g�(�m��Y���.�s�ѵn=�����W����猐���ì/�Q�<�h�Ǽ}I�%+-'�����@�/�i��lJ����Jh�l���5���;pb�yUkxP�[����Q�'$��A���ߜV�?��f��M8��T^��δ`���x�*��@��[|�'mjA���l&�m�	�#T+�EZp�.	���U&��f@R2��I��T�JA�k�3_Ƈ7�|{P��&�������#mf��+�aCc�����U��_�1-i<�R�va�밧t��'��ۜH9]�u��bl�3_�y��"�;��<��sG�}^���ե[ex���nGI��M[!��)�1��S��\�x�c�� �G�4���>�,�E,��"%���\��v�DO
Z�����f&u�����k4���@�X�!�"B� �3}-�䒞����T�7uu��F��J%�7�I�:?M�W+�Y��~KɋՊ�1�HL���9Z��0��H��U���.����`�r7E^�3<t�^Z�I�k�ﭼ�J���"�s�����G5vzq{)C���璧AF�UO2B��<���,h��*��1�	��S0d�q�AՀ	(���>C�!��%���gc`p��[�Jt0�:��$p-3.\zec累�l�C�Fu���mׁ>H&[������|��t��Y[�||��F��V�Y	���L�jtt����F��3iy�g�,H�)֕K"&�W��X(��Zܓx:ťs�[�z-��t�өK�Ҝ�&N̸&�ts��D����=qET�,YΉe�6럅�C�:�F�@���wFN�
�Xj��:z��`����)O��_����'���hZk�@��*��P*1��=p�0��=@��Yj�j��J&pA�*���*�K"�q���]��[�JA��ȼ���xir��~�A�� O��=�E��"�W�T� \���t����1��e�F/�4U�����
ә"�l"��<dդ�я��F���(Ɍ��(�U#���ߊM�����tp��^]���Ш�m��3B'2fb�:����Y��������l��U�h��<w�2���	./X�!!P�S-����M��#��s������a�d��4�*���dm�n���¥R]O�T,�|P,p�T�]�eһ{�=�~h�&�UAQJ���F,���,A�/�~]+�-p~C7>��3M0�"�.��'��1�n⼼\1����#}��/���"���+~��X�:++_��+�B�s`L�������PCa*���� ��l!w�E��cp+SP`�]u!�z�퀅�Zտ���Ȫ�w=΄���>���&
��[h�T���q��&tV�CO�IzV�a�YC�����6����9"/R���n�k��U5��q9�;{�bI㿼Vo<���͋]ո&�ĉD������l�_d���(-�]n�_�G�\sn�U�C��Əw>�JW��A��;n<p��W��.�UH���
:'_�wd����ՌRׅ��o��rq}R��&��U�1�:��m��d���Z�t�i/h��h�����c���w�^�����vu���}ŭ4�g��!�uJ!�O�h��l|I�.����Q,8�@T1C�9����\�V���#-k�2�_���:�'��L��bh~�0��'�2{���@kf�sio��܏m��=P�7)�~�C��^����|�B�W렑��C|MT�j��z%k�<
q9�qxa�����׾��B>y��A��b<�sz�������z�cG��jE�
�VL��P���3��D�Lt.�:E��3��AV�V��>zN^�����RN����5l6��.'?��m�����H1Ȳ����}UM|g�h!�;�᯳QS�Oc�Y���Z�@�=r�+l�3�5���p3�Q�^��%cf���F����H�Q��H���m�ժ�d������l�t�lH����C[
��*]���O������q�����0'[����� �z�Ag
1�I��ۋ��l��3�r�~���d`�g�v%�V��[l5�BT�#���$H�(M���+p:��[�E�Hؠ��e�2���Ʒ��B�'�.�� '�9�ӑ�> ���m��N�6�^X��#M~{���C<��[1������l��-��W�[����ys�Z��/��SJ����!�!��t�2
E�M&����G<[�������)L�)���:�Ч����Wo���A����]A�bɫ��(!{^-�.[qE�C~�+6��g�e���Bn��=�����c$�M�<�U��M�,���	!���oN�)�92��ٱ�{�Z�{�/�����^A��(���FN�M�r�q�����zM�P�9��Ξ<��pܽs�w22s�,"�i+xh�a�R�������ߥ+<%��A�6O�PQ������j��rx��Y����ī����D
/P�i�o�2X� �	 %�RP��o�LD$�n
ى��G=+�2\�<�il�G]g�x�'&���>څmm�:ӂU�aZAc?����&Xq�	�����1�JGeE`�Z�
���	<�ڴJn����屠�k����3�glxE�mU_�zr�D�Xݝ}yi��e9�����]σ'بK�Ѓ�0yV����Nh%=w�l&p�P�q��,A[���c���Zz:�7���)�lޜ�Ӭ+��<��b�)渟��d�������L��R9�(��<���팣^gč�}=��*��@�g.��I��ã�>i^�6��d�"�|M�?����������J���G�)R��B��o~�Q�����5��L��Z¨cdI����ɟ�`&���O�O�N'	�ɒ��E���>��/{8:��H��}��>[XY�8�Dn�c P�)��b��u%�qg����XI�Mÿ�"ےK#��(��B*e��� �N�.��W�I<K����0�¢�����¶/�s}�C�n�=�p�{�D�̊����"���9W���E��X�Ӧe��b|�zY6��w�v9�V�ʦ1���S@N�H�p��;���F�R���w(c::ކal�#{�vM4!;K��8��P�@֥�G��l��*���.�n��st*:I|� f�����fE�	�����:���.��p�	�.4�~�����21�ƾ��h�l/ �,��H���Ł��i�B=?Gީ��nK(��	2$	�l�.����Ǚ��-SH`��{��g�7$��� ݷJ^��m ��� zCp��ɤ��c�ĥ�V�ݣ�̲�@UI��ɷ�oSh�I�>�w��"c��z V����αZL�!=��NI��9���9yv�)x<́�Cw}��쾯\=��s4��{�U���.2
e>� X+xOuӠC\U|��� ^Y��v9�O��l}�<k��d�PiS�Tj��sƢr�_�a�H�A?��3�ou-ϻyg�86�FX�E�հ�w��6;+�����D1N2E�(J����V9�6&���E6^g�o�����i�V��>M�8@��;�����ȫG�_V�E�f��+�9��BH�r�1���r�M��}�Ʈc;Xwq�rU��,��! ��Svl�($ey>z)T�^���?�5�w���?$Z�w5�&$��Ϊ(��w��c+��GxG){��qO6о:���9����<��z��M.�z]���4�ʋx��cLgA#\�ƾ"�	t��=�Z�����T���CbQ�K�}��_�]�!vC^ԯ���*�)J~���_��SLɸ`�3XjS\̱�|�r�:���6��%����������$$	�GDݹ�b4�(Z�
r�HkJ�3j�WoCx�r�\=o;"k�JU�� &ŀ�Z�7�b�����]�>ٷ�m9�|'��ȉ0��q��������o�@|���E~b�����<˰y�U����������|m�5/ZQ�6q��o�y������.l�4�?�&2�o(�>$-ĩx��Տ6=M����w6rXD�Ƣ�YQ��=o0��������@T�]Xձ��ʛ"�r��ּ�9��;��gU
va�WC���]�Ə�	L��[q?��,or3�q����_�/�9���_oj=��}6�T�\�ړΡB��1�C06�?�"�KT���/��Ń���@�3z���~�kG!�t�	��շ�$��g������I='2H�����;�������o�dK�=2���D y���t�ye��һ$4y5�t��]�����7��SW�L]��M]o�C��-w��:��Ŭ�E�O��C���t�4J���iɢ!)��V���6	��}5��;5E� Bn�t��W�t�Ɨ��;C)�����>�ճ�3�T����غ&~������p ;o'��;ܪ;K�vvd~ڸq	'
M��{4�K��=h�Egԑ�Z��s������^i�e��Zи�QYh]?��2�{�u��I6`3�T��";�\r�`��&�-8ٯ'X�.8���E?�L��p��* �����[*$����&}j0z2Fߦ�6��d���	�07�G�!���o@�Y��p��omV�]�𾆰@����Vᔜ�R�R)��MB�n�ݝ�,.�/i� ��H��i��+F����jy1�Z��=�2U�������6r?ۍ���ݎt�ݡ��H�Y��1��j��`Ä}��ڎז�q@��\����>-�g���/g��O�z+��M�����[�b+V��H��r�9�vVh�R�螇���، >GƑ/F1:� Di�����@�]���D�9�^��<|�r��Zw��B��M��9Q�¹L��-&���ӌc0�Go����X/��>HJ�m�V�p��!.�.���������CS�B��!+�'4Y�ab"��;ԻS���WR�����n:�&�(Fl��O�<�b��W-�J�R[,V��	�hJg)9RL�V%�ƽLId�h[�.��~��E4�330V�ލ]��>}\�;��2��8��xF*�uӦ;o���@\��u҈�:�U,���+����vDU�7Q]N��m��$Aٞ��'�}^q��S���ĵ>�lS4�Z�m'�m�M{*�V�,�i��A��x�t�
����b H�^U)NF�]?u#�������,���L�k���1Y��Z�%.�F�a����\疁�*���[�^��J7��DMؼ��a�Zn� w�1."K5 ���af�3����4�X(��\Z���iD?\S���kv݅�9�S�Qg��z�ֹ9'�Z�� �u�uw���#��ހP�\���Dd6jc�e�z���-ԏu
<GŎ�8�n�:�X��W�V�6�`�P�,��7m��c�@ϒ�ѥcul C��?_ܼ#NR�.�V�h���(����:-/�v���VH�	��!(�XZ��P��GU��'��1��?���.B���F�[nz����Da�l�|��I挂[)�:���ҜŲ�gw�P!�����L�����8�-�uރ<p��Z�"@;���Cin9����&%�?T�y�K��X?��B�| �n��YH4{�<�lvw|�����]M�z1$f�?\��Â�8ټN����,.=���zF�(��QҤkr��X¯�����d��CF���-�R �|J��fK�s��c 2��ϖ�ǩ�R'�ʵ��4�۔����4=������-��(/,�E ����}�%l~��Ļ�ȓD�o����E��l�U'�k'�c+��s@�"�����!;��pƫ��OR
rL(���Ԧ��������p�9�P�^-�N0�m u���Fî����ӽH[���FWh��������s��_{"뤽vٯnyYO*�l���̞ ��yqO�<�D��?TűA�bi�\x�B�>�R޻�����'h�_r;�����q�����YV5�W2��v�����M�4��p�9��[Uc�<}���3y ���tf��+�ū�n��r����Ì650=M)G����ֻ�Q���$���8o�D��Q5�sy��D3XB�۝G"s�~��8R��?z�;���o�
���{�t�{�Ƶ���L�_b��P�>�ˬ��3�4E��n�� �b�4
�n��}�AO��:H�ʹ��nj��u��&�X���NG���2�d���h8��r�Őh�����L�)�ll��㼛.C@ tA��>�S��p
�ad<{���n{�zk������pM�y�JT�� �R����H��z�E�����i�T�=��9$�fY*ᕆ���ֲ�
�lV"@Yⱐ|=3�w�$g��~�Xz����+~����K��e�yߛ,�v��`(ͦ�uټ�^��h�-��w��<q�-�wv$�����uA�a��q��r�F��~W��^��b"�����?#2��9��n�=�0�V������P&��|&3x@C�Xg�r���9���Gl��������%:u�|�`�;����|d���j}�@#U����)�4��O��@m液��\�*,�O�f��j =�F>af��M�՗���傂�
!Wj���_�D�7�B��˧�_��3.Djg��
�I�%z!f+K{�2�.��k�rA���@�j����[ݜ.�H�COz��v�\7֚6��책[A��X�є���q�ϝzvf0Ŭ[�"x k;���~]�=ƴ"���{s�r�4v�I*��)�U�����ǌ���,y.�'�^#�]S2����	_�C�H��]�jk�~Z�A�C˹4Q/�I��K���rW�9���C��c��O7_~ଆ���{�7��-��S��ƔM���W���� Qg�0M��b���ڨ��yh��r��i\ZЯ�1�L*x}L��g4C05u&��R�_�Ȧ�[�U�Ɖg������v�K�����WƜߕU�ٸ(4���wu�_am�E�^>�Mr��恭Ku�J��'�a�����