-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Qk1EKbjkkTfjQo9E/CI9/reQUPTm89DHyp8VkzG7D5mvttD+k2vFl2AN0Si/KTaJBdKr3IrNgxyn
XPY3cCEyX2sZZHCCkYLeH/iepHi09A4Vc8wFLBIOZ2C+Kf494Cvi9+H2ZYtFyJQYh0KlS6jCk+4/
/0Dnbj4RJhrhPvWpSzDFKszLqNF/4R9YYHSQdjLt5pioWRbFtc7ZeotV1jUGPJsUFc9ojXO37dvK
LUzLwvHyJ6IXBJ14VDkWJgZ2iwL6JJySN+Uv1ZzrRk11NQOd2KyNqOrY8237ce6gLRE7Q44QSJXo
aeJIP1Z0Fg718v3viStkuh7faGlYWEsI6vOu9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
FWUzaKnAZyI09WelCowwmtaKDT9dx0Fmlh7bFodgVRuC1MM7U1A5OVs/mu+J2VXgfsXyvxSrYZNu
lyKPJrUVTYO3nqSI/ySK0Y5z9BLup8s9jY0nVkeWq3Fy9YvBeZNmy4GvMz0JTjp3N8HhuLm7HjsD
j3zMEhqsxQOGkpgcWi0JWlt/tXKQNRldup1ekSuBV+KKQDfGdo52p8H3ThuJi3NzE72dSD4n9vSd
I/4Qg7GO83e6OhHkiL9LLHs//NbfD10pIiuJsvI3APCl2eXBfnsG51S+QzbfMXFEX07e49DyC1CJ
GeSzv90bru2zcNkNBVJ9R2oaF1swD8V520niRoe3Fh426dTsVhvI1SlpW/sJ+NZggfEkF8oxdJHP
fYrkyU+bv4QTT5dr/hHSQc+ect14AAbbLwZc9ivv6ABDG84my0DmzHc+l7uTsIfFxoGSnXZgTK0G
HOJT7V5PK2rY1b6+vSsI27sv6Ae1saaKtHqcnn+If1n+32qckUoodhbxsxbGmdhKTykZs+HAOwSS
6UKaMD/1zv8hxbRk0++16Np7kJdSKVEylIFv3esn4KRQRnV9u3QWkBxk7AXSCyQL8uzGX8ZWd2Hh
5kc/zxHkkCn/kGMwIW3LRkpxHL7UiB17MIpBRqd5F2DgLwqqkBURnr2XSSsjvne2NInczxXqsqYh
neLl8tIOXFd2/NTW+iyyDSLwRRUZd569v4Lq4ifnDuMCg2BFlg0SgXEArmTcvtr+3cH4CGJXoCpW
puaHIeaxPBagGkeicJwx4CDgSQK6ImHTEg/Ww6N9mUp37lXazFWhLrM41MuyFZT4BDMB/0Qx2nu+
adwNFSc443KLEUBWun2GMKNWa49rrvjwUUFb4fMGenZIKuCRoFVkHPHZN/Je49PUKeeO1Ghjhbg0
WLH57p0qgRQpXBjGnwOTKpcs4aRpP4fVmpgaK6o3rIL2Y2Ff+7O40aYncLUfvwk7voov7oCQv5vW
ffOgIY8aYvzyMjqjPx3ZXjXBHGai9ZbKX2EzaXFhxlgj/bUCytB4c6D9kKNVlXS02D+71uXTnRQc
gXcsnGAMJxLgEmi0eeSDGCZH7kps4PJ7nG6MELIkosRAKrf/ofL1wpCsZYGRXsGEFW/fGRuS0XtS
hm0e71WSH7eIJaLWk1BWz078lmeHjyj/Z435zPa8dHIBR6hS3fukJBsuqgz7J51mcnqzsbN7E1KZ
JyjGqIEpHKN8W6QILauTTiEbjOh0Hl4x/QHJ3yE46OBhd49lTvoB3AMvN0qIKbmuZw0n1pRXaPcU
CAifqOqxHfu8YSv7O6C+dFceQ+Y3vVMrL2uc/0s/9V13mRGqIZmSXz/rzf/lBzyYs+SyPnekPhrO
OkdWBzA2aaHSTdhq7oJP0J9whzkZwYb24yyzgcOF7a6JRZUjJFteKBDF2qsb0GOIOyQTZyvCE9nG
0GrHceW8gVFBT4/FoSMc2HLv9LuGPFCaGIJ+fr0YkOngGCnNf5EQ+9tuH6+LYuXOOVKbexPxn12k
/dKZCkHe6r1+5RPOQahkq4kSEQrw2O/JSEwNaUwv0uvaUgTlIE3gIfYG0xHhBCrAx/1AGYf3L0Jb
f/ZfisEOBZqPQqz45svAuHo+qH/BWhEDUBlfZFKhbVuBxbuiuO0G0ie4MHoD1HXs+oq/S4gUneRn
ykcTZPvbnc9fnNj2HIgMViRF3IjxisQkU7FFW3nFaQnBPzWS2KPBYn9SL+Mm1r9RcnJCpcK3AJX0
64kNFaY02MeyaUkPKcZphTa24Txv/hj20UbfrXklOOXIa7Avjh39+VXcha1zD5ovzek27oautc+r
NvW4rH0CwRxjycOatiEKWCKoVIEVXsdt4gS7i4CaXUVx2NgrUcRRfz3gRx2MdYGvKcpRoqr2jD81
hSFRR1/dDh0vOvmFT8fNVVFixhoHpBWxB8Ko33Hd4xKComVlDLe7OR/RJ1/7pDNQrBiIvHcOqYup
0GbTY+LvhJiWnD2lJU7bjRnD10Levql89jNpmd3fFf2Wr+hwo36zltCOmlp+ShV748Gqstm/ctxR
mlHNW9SDoRtgZABslXOVO4GKA13F8/BxQJuaEn+BAPDB3YsdNlvhhQGLkfjidd2TGhAc2hTUSwLb
QxxwaiOO496LjIu9+Ao3Vyb98MhPYBFQVXBlrecYGXJDAZ5iW7C/G0piEGjAAEv6I/AoXSd7we2w
zKmWwMxu2OkPcQdyY6qmb2ahNuXN/tdJ7N0coSPLmGXdA0jTfzExFI8corp2EyejnqL11rMmIzEG
6ZWmq0jr7f7cuVvg1LpLvzW2h0nGIL3frz5qoWjVgLhtuUp1+4gSnrKUsfIQjuTZj5TTOpS3DiPF
5qTD/VC6w7LZ4gbT3qzFSxEnBG67pJ4rpYLZFH++kQMetvYu3VLIbpdJHHI7FGhjJSTZqr01b0Gp
PnQZC02V2QmyGyGTk8d8Z5+g2qtQzOsXjcixZc89v51zazL/7aLJlTDSTAFb0rjgNHkl5mZH2oCI
Rja2zIYaLGwXHSPubivBd3JGRi1fJcNJAl/CHAxIArHy3voQwfT7nPfooHsv0QjehZLf0CykgJbg
KCHcOeB+hJNhmGuylRa2jKnjbK/uREpq6xsEFTJiBhJP6l1wOTxF0s6qrb9Wj3BmdYMmfVuIVvdG
cAvonNtr6xLee75FvbVpD6JcRSE9q2Woqd4yBNnPn7fYmK6FvnpX0eOFUPmLbPNojDUEIEoBr1ff
QrvfVEAQo3kLltfcWhH3smcTwgvjP+PQdhtpIm+EuwlEi/ILBWTtR0+3pHd8cvE9wKlghuKYNXyM
aHRfaM25T/t8RuLdPTRojyD6ZJEXF2oYVYePifPvlLQVbmj+kAWvJAoSqLD3efr2NBINEIbFYLOP
SWyUUgLv1iMScnQQteIqqE8REwGkHpOENhZOfyUWK9WCnbz4rktnY8lOEo0xWx4PJtdRhIIav3jO
VXiNV7cBv9AvTYWKvuvfNJWpYIpx8zY2QSSxYC8x7+wh61IErC3+5vD3ECg751Dwn5WAOzqpr/Vs
s7S2sySrlYtZW2OBd3jQj9HnHvILu+bdG/Klt6iQDEZG2Fc2QYsizUI1jQ6wvMbb+O2EAArrjlo1
Pvk4lEdpy/LD4B6bsp5PBi+yoAj0DCIaDPaiQiOZmjdKTCdHN8IMJwgEHDYksyTmB6e6izWLyXAR
n0R7G7cxjuLj9+CMaoxtwT8SOVyhkCMatZFFbrNdgoBLsBX5hwojVhv33QOJmttnZRXnXcG6P/hP
Ov+XouleKS0Eg9Dgnv+Ku8oEi2+0XpU1ZAAHxVvWGGxM1ubEeVzzZByXH9HMDrjTZLrRqWzDT+Au
lJaptJPFhGlWHjOlXXDZfWpW/kO1E6KtuliRCFztOeS7orOloFEK914mqL4qmB/FFuN88w1of1cz
SImz8azPn33l2cNmctryrWHv8LllKFirWiQpztokDM4hgHlZwMhlGEdL4v9ye2WEngze7PWjFvuz
SUaB/7fBMSKuWwAEefH1xvEKT1Sh+tSGyIcX+65e5VzygmoC5k1DMfxdjNDhqb0aPzzeF1gBs08k
X9lilE1rW8p9a2hIKeEi47VWeZhMzGeFdhjYLeTFjhBQBqy0wKUNuQmHQ2eBMow5LdQSuMjnFISy
ezpte7G/G0b3e4JNJmmvBdW3fqGPZgjbHjj8KzkA4HSBv8OQE72oROLUI/WOSuAdN+Wyzcyfh93B
SrBSwqLYvvB8cmHwgAcg6BzylXRNwd9po33D2foeq3O7zij4s9A7Kt8zApMRIBdmtNdZR0cDcsGt
RGqe7gfUN4omqJXkQi9L+PGWQT1xwgl2uBMQSeg40WWe0o1QTCXuVB1ZkYNLNgEhQh8xK8XIJwZO
/HlGm5REnuRvF3TX1dR2pq0QxDhF0GPvHcsG5d14MXA96woYDuLhavRQqU6yU8KLN6PBaBrOtDix
4E6s3707ZFVaPJ1ASs00fR5dcOqWCvzFN2DDXzUfJlob95qeMs9bFpI1oxGZruuXF7Pr9Mdhd/22
Ph3SWfXjUyu3rYdypP5q9t6XOa9Qpuro5THGvpOrwlPL3rk261b+tAbmnrUzI/JbhJT9RFDE0pBZ
FNyUy6Qx534uHKbYWEQneHyeWICr6bceuSM7SZMkgvtuKv/yjjXKYHUxABDMCs4EL9ppaCh9iUBo
p8yYVI1x44DbhghK0xcNLnfl/j/7Yt1c91T+d/fgy/YzZo8wMy3GhzYxjfZ/fzVb0SVSWGPDqNXU
+swizPNR3JX9FIA0LgEZSI/bzOqQDqAkmG1w24gOvELOvmJVUkxg2oqtYXFxaFMXNadeb4JvSngD
MHouR8pSQstBcm43pMo6lO7Ec6M46ZkaoCKtpkhgXNOnuKUiGMYyW52vAquQsVMbLZLX+5/AESWY
HTyFd/2j4YOqRq3OyJ+9kRLWIxRLYdSfvr/b3mE7dbIceDZ/VwvkanSDrf2M/I4tkePioPAHL0r0
Gyuh5fuXVqTBqktI8Om1i1709OSSb2B9wfbYfKm/onjL1LVBJtlFN1mkR09PKQb0Q8aQnzJ2akx0
QL1FH1/PDRbD6ohKMXTbcMfFX5rKbXTv60uBbYSOrK8tdraoH8cA3vjEZSZsRd+nBmvly6kLFQO0
VeTmcGrYBDzGVXI5f2gv2X/QQaqXJlXrPBrQJZHVhWcIUDhzaB0J8ryo1QSzWiJYlZqzUW1bLFV8
z1tPl1b3/Z0cBbtR1DY/K9U+ubITk/QCSYqK4B5d61/ajclo3ck+Bs2mQTEAD0RG9bOk/BiARZ2o
62I2KBpK+KEzpJhytRmsCx1Fj5GteN4bu53Ebm/b3VaULNJSs5e7f1DA0POpO7u5jVC6WZ8JV5tz
HQp2P/UfTTju6ILK8krih8BAOg6EVLiVHEf6VCnA0Dn67/ziaR7FYyeyKxXMFuuGirC50vU7LzZn
/zYxZIsJz1Oe6A4H5YO/TP4L9qqK3D/i9IafMFpmy+YH2MSmFf6/YtMbaXyswaXZrwbfjzF1cROs
EyAZPl8u3DxvlOSG2VeS3Lm4ICMcrZHmlfiWlv09j+lrzlJGe5300XOgb93MbqEtpEgVOtxDm+Wt
8kICohAGhaqMDwnMiLdmn7q72Db+9u7lhzvAku9QCjlxnbmEgHeE1eZ03SIScKwuGO+PjtjhbiBj
wVB583+Z2R7Edyrh/yhjC4oBzKmUhTivN1yW8pxYxeLn13flae0ijvD0nDguZgG9CKMb58SS8VW2
lRufVFiUokWayVaCC7BjQdUXR0MLycN2n8jUXXH/NUVlQj2AN2mSfspJa+f2i2woT0TGPKx28vHm
T2Ur/Fo/MFo+snBUxcazbOyFCL7vPkqKxgvIzCHBFNSDPBKiEILcGPE5wjRiaFEHnTj3IZc1VMpe
KYlFfBJtxelFbA3xbRj+3Ai3HCBjq71adNNJJ7m5eGAWZpgAN9Cxl2KANRfkhxplXvwmqJMMUx8+
Mu3E9c/wgsJkyHKWefqUi9ApM9MiiYDwDxfsJngs+kbSDPHkKL6PXrSDx8s7eMDKb8IG3ajRU//Y
shocKD6U1ptVSCALXwbUUmKl40rK5UYEcVqTmoOy9BfmpUuLtw0JofDsHP6owuAzJwaWmFOfvPio
43h1DBGgkW9xZL1Jf7xJx97gM9sSf0g33j4gvdrc61deM+sK6QXe0XOECxjAX0eWV77enOSdmmSS
eGeyJMbYYYKrYJt2GT42HA7wgWOXWH6kH4w+mtZKJK2MlOPxJ7KL9dFbgpBNlDqgRxzppLDEvTNg
vgoJQNxeDd8jMIGSvRu7W2JNNcYvtSHkM3vDdGoAV1IgtKG8Utc3cQ1pUgXUS1wpQm2YNUOXupFP
zhYw0b+207nUgFFt/rGlkMT1cAcOvgDTqqJ9mM+jT/CdzgZhkts0goumBjnbfdCE+Bb8gjlnrNkP
iUQA8jEaNgU69iyzlgtYImCq/DKNyQu/84bIeGcdcWVvPjjAKcM1z2GpjrlE85AJ2n9iaRXEYKAw
DH7zKuSr3VbEeJM4IbS5CwEe+U8M6KzbE7a12d10+Cshh86iMv8oSqaNMPIYdDVnsDAl6LJF0qfM
PnyqEHHV+tlqic3IFSVJHOVH4D2z6r/5CEKzo6fVA6Bvn965jz8r+cr6IEZ8t7pB28rj00ezyK5t
en9Z01toMDGank4xuGv0GJlapGngooUuaN3buLWkL4s4HcSrxt7p4w8OQAQcDvWvutMJhC5tl372
PjNCmRNHQSCI/SnezO6VzG0bi6r2EP3HBhScBu7doA0PKj3PyFM7YVO0GjKw0GubPhvJkBLUbupL
SIXVS2Iyym63d2wRaMWCAXF43Gw5QGeCwOjQD+cAStYUi0IdE6BopyibRIjNq9m6e03CDiIARt/D
bZc0BmWIK5oBiy+qACKyh39bjU8ZkSRWdD1vTedkuR9XGYA9ZTZLuf1Sh2tEQwb6nOE5T2R5OJ5D
WH+yVqdynJK1UbVqshQE3961qnJqC3OXA51fR4i71HtU8tuSmb8o4UOl3UJH2tUieC0FWmZeLVxy
JIS+8uxcu/OQedWyyrpaoyz303q5JxW2+W9jo8zkpaC/1HvmxeP1HWZ0PJqYPB13VurzpdWlkpD1
FSY1PH4WPP33MdAgJy02CZ3iAdo7dbNiFHTSEHggcQO9LQzAd5leWyvptLnaxDPmEEz1Cv0ZerMX
eBSTvcpWwDSaDy+AN/Ef18WaaGjPod+mwyqhsX8XVWDQugd4hUow5jeOe/+Qw5nZj6VOetQ8Fj/r
XHpPHkk/bombiVLe6K5FeZUOSx100JnWtzYxwF2iB2aJg40mIfaqTRuFbXgAhPkdX2uQGUjuVN7J
x95s961KlUOX3VwFJS0ND5Ti+FP1CIIr/ftqqG2uTGliHrf8odxIxG/2EQrsFLR/dIFoXADJy4hH
Wz8UsBpZnQqFXi/lVEF6dTAtUI/sokBP6hiqkpAxxBub0VYidpxCTheMjoEzpknf3/N2CNsxrWtW
otmfawKRi+elzeGps3cV+bdwzOFKVU4H8uqgCXFKr6TL8WpxyhTW1gDr9rrG/R3NQTGDuVhtI8gR
Gp5FfWRiaMSSJmFN8dOQgZ+mfFnKSwlo8eRnYdDaXOrZN2K4sRpahYEEiLHIKBCOC1TP8umwjQ30
Waf6mcePKqAn03GQJvFhUXgUds1zV7ylhimEkbf7P5pKcV3GTFQV8BqfJJlEzcalId8A3JSxHUXW
NHbMi32pTjakauCZRh6HYS6p7/O+AncUR284hjGmsRw15mz1yPuAzq2LCMtLdrR1wAzO8ZlV+TvT
G4Me8A77dY/yVDmuu/2bDFtBV54WDFGN1yvtjHV7RP/zyk0abIns/fIkithxyp6fjnAXb6AVHwb7
WHiuLc3TB8KvaZkEWgwckPUw7+VKwuym37XaS9HoDwxSgFkwkqNDy7Bn061eS8AYmEsnITFHvo4i
z5Lx1ZpeRzuPVSHd0emQjAKvniX3KPhEe08XZoJR8lRk/1qxn9z80g08+5Wi2o/9Q7kGMYs+5nfG
jPk25jbe7tTSXbnzWqPM9WrDfNobkAHALpD/MOQueelcLHLbx/CwIySsLDCZq0vHSs9wL/Pmxwmy
dIMtblneAKy9JGzDqjTQRNoy24EumZ/51M5VMx4Xpvcf+/3Uyo6h9/znbkmgFagM6WdkOPOSsxAM
ZqtwgSrpe5LwFrhSrYcG1/7yehOwhQZCCQKa4YUJV8bcOYXI/E/qfMK1fdATE2G3KH36ewb5u6G3
R7LFlNuZXhsh+zxQ+YAK7Wm3/BJ653txGDBiLMbpvx+7eSpWBBmHJHin3A4M43Puw747v1cSgIj9
cOP8uvxKhXwC+SL0VuDP6G6C+Y8SywR7TzPQ2uU0xlZvs4vmCCJ+5rxSlRkG7ClnBTfosvQZAAdr
ohWvHSPeNqGVDDhrgI9KWleWRZlLEGkXSZAbaAOG6nhDqQr3skLfnWB73fU6Co3sEJWh18RIF0qP
l8oVrlTlRhzFIP6FjKES1NRN/L4KaKijPH7xC9UK3cVYRkl5ClbVxVLwl/HdpBtpnd5PQTlCtpRN
oiLoZMaJ7FVktRtvK1RzD4tExewgCaU6xFIiy17eAZQ+O60T51kwc6jOgjO0EcKR97pYPIXGdc9V
ktD2Dzb5PRYgAfyq0IWfDmBU7QniYDGU0VK2x3tCmcqPP3Q/4fcXs5jlET5UWVVP3yclPu0HBLMg
XxqbbXnvDqu0v6lEp/aSFL234pP3CNHQfmz3DHQAzrejeYi7ceCHYU0GhbZis68/2gSYzgQTwVn2
YWpusAxZylGZ5/1E6fdkS1Ez+LCFWa9mFl59/lef9mgjjiaL8ovK7PqZ8AeN2FEYGt5O6DsLXqbf
e81F4VNw10tuU1r4hsbb1VrHdqAabqIXxGmTUy2hVOZxwyHDPQF6XM4tcfkEzepF4mbItQaKRLhT
UnjtnLC7Kjwm4J4ZgncwL6DCRC2O2zARMI8Yaeu2N3lTQ+oN3zKInGUxWRUH+3KtYqM3KWTQ+e1S
veaVlon6zaWOgSjcXzX2Vk0YZV5ayVx5rQ5PZiFS30oY5cWMChIIVlqqs1aXY4TxcpJyFjWDUT2a
fjmAsfmaGzbEgu2hMb54KJER5uQHjlvJBBm2nHU1tWdi6IEkS2rfn0oIHF4seQe+1T/lDW2ZK3Vy
rDxKFCz/AolZBRQgBFRCW/1DOo+RIwx7M/eki6bxGtfohOBwX7viD+PW6ikJWkFdKDt5jHC7Bkfq
v8N1rL3OO4SWr2i55UOPpHAdT7X2gYHo/+/XV+iq1dki2pfeaPwGoi0Plmu+ok0ci/sSOVX026nS
HA3Ts/jNGzxK1By88z4e+hQQ1yN7FCT5jVFfmGc8RKXEf/UccsYIbcUHU9WDzlZlmLmvApPHSFz8
dfEJdyOG0mwcZZip45jzVjEzKr01qRBqP2baRWCCWZARZTIdZKGVozfPBy5HRvdwNXRMgtFvR3OZ
7MD1ah9FLWbmBZ0F2DVGz2jHylfoNcP+LzYctPPOWKcjJ6/T9qrrvLqj3wD96pco4YcEoGsUQqbE
E2mv2LMMpUCtKop061SU3d0MuT5yQhNt6b/yZQTG97bmvQieIEboG2m5BeXjfLpXk97tmwd1481/
cyGOJIkE++nsbCsxf8aDcRtp91MKkk9ISjZ6L78QZQTA0oscZCsNu3N8edcPbbQGsPCEVjZp7fUE
drx0kvnu9/z/NkF/rxqx8jLfqtVpwKK/rlgk94ZQw5lxjOWdgjSvJi/o/jhrNcgjS2w6peoHTZ/Q
V/uUVVsu9/Ug2KigYZch1uZHsgtDOLDbbd4KDlVk2ZJ9ed4kWczt/d3etR3hVov2aQ/9QtC+5dm7
bJCHDlT9M9oPF5vceCJm1h06Laf/DYABGbTGe78Xv6yDpoRZEwEF7SHe35eBOyCocsyugMYWbhn5
rR/WUasJ7LSvhvfPmnBC0f8usltW6OarESDMia7vnFWsJ5xQ6gu27nl4xFWsvZ05EH8N4uDZxWyb
M/GXOXlbJTgEq9/PvnJI7pKdH6hwQDSuzMDxPH4fWKYxtmW9sf1uZJFS1XiLIybpfC47fjoXlY/Z
BJycC3FlZLa8iRwVf6KVw2AFvyuL29A2FhwtMeX/iQp4rmY6owrsuV2BBnOEUFkOh09TLzobvf/w
IF2FG6N05D6UUIj9GJYmF0z6YpXJEhnoiatwxGMt3cbEiTe+BQtSYUpxt6I3Bj5qGOF5XYES5X2A
Nz2ViPgThEtwzWEuNZoiNhoGRoD/cXRKTP5pi+VvKaJxFsMQ5ucglrqu6CQ/DJ95VuAj6eth+DB0
02DwgenVymESMB5RgzVcPpkzBjtSvDeIkmzAbUSgsYCg4GK6rP30XCc9MjxxJXRnNhxg+LyQzZBI
YXKJx5iUoAsheOkK28PBqW1KtkCU5xuMncNT5IpX2uDOxqfg1UeDS/Fg0Xbk7RlW52bPQsu+fufH
RpoqPScpmDdCNnhxfY8zmWW6wHdMTE5N/wQ8ojy3RBIV/CaTzDkDNbsM14PSSZaWTzacN1KL7Fia
82ba3SLx0/yaHOJdqNDpr8far8LkeRJZ2y9iPM6AabJsa8ZZTCZJFxwDHzr8KxLfq2/eSPQt/85t
3CiPp8hQua41UqnEURrllDJgtB09e7AWmkIlKQkm8NjyVeUN6P+05SJOAvqgoi2pYMRioHaJ74XV
BuJRYigPPSN66DHHcEhr7A21wboN+7vNgWkd8Oy9AuMjPQP1X+b9Xo4xE8tH3BRFob9DOvnSlpsH
2A==
`protect end_protected
