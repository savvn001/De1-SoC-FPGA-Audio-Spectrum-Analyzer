��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yli_��#js~
<�r]�72צt�-I]��&W�pٷUT�O#-�@^����(��|Z���7�yH��=);TP �7	�(�@{s�`���������^~	�_Ȏ�U���}� �v�a��cįy5�Ʉ �̑P��W�V����;@)��c٫`�~F��YZT��x}`QԷ֎7к>��ww�m��ӆ��)k�Hx�=;��V�ֿ��|
�X���vb�Z�@��ߺ�(�V���%�k ���a��FK����J��6��Mc�l��e�d�"⚲-�����L���5#�B)�g.�	W�#���}u�Y�ɉb����V5%���7�����	�'�D��a̕���_����� t��Ş:����=�M������?mQ2�A����!���\5�c4Lr�hD~�.hV`�E�\����h wѱ.�U���ttG %%Y��'d�у���F��7�;��z���>=��d�Ⱥ�0��a���������T��ϝ�^�R�
i��{@ݦH��o��ToS��O�C��eM����
�����^�3m��-˟�O�&��e�GPU}}��qH?�WV�g�J��`mVPܱh\�Q@�<'֐7"4DWW�����wΣ��K~�Y�tbE��;I����diJG��h0�3�Y<;�dI��>:	�%�]|�ҪV|������H���]��cfb��a��bx&@ϭH��>��=j�c�-��3=��d2��<�s�1�
fH��������E�?x����#�2gq7e�BDB��[t֍L�1ƕj���5���/\v��W���BB�:(���ki�v^8�7�[r���xܝ��G[�r��QΚʜ4��}�b�f>��A��-��ﶭ.t�O��%������N�k���Ps�$�[�~�93�����g[;��$��4����kx�	9�b��PK�M�S%�5��Hf�F�R�{ᔵ#����7�R<h�x/�!�" PR�V벙�y��"(�k�Tpr���jU*�+)s��F����cnE�\Ek|���smK�l�wM���0�+L���xI���H�'�9�%�����i�F��@���!��)`=S��=��Y�/"]�B=Yކ���Cf��`�H�/�i�k�e��kr�d�>�L8��<���xk�yC����6{L��x����4	���"�J�Zq
���A$��%7,j���'ٜ �W��w6����uUVn��]L�����ZX�͢ #l��18��Խ�OZ,F�Mq�ᩛ�� �;�h�;��=�}C2��JE��i�f�H�C]J= !sN��&��kEPRm�Srs{iȌ��~�nι3(�y�R��s�'���ʦ+�#%�L�T>ݪ�ޗ)�+
Gq��]���`�!�F��*��71l�:�'Q����t���֞P��`�(P��U�E�#�����
$�A�e&b?�G�6���a���̓L��r4����c�9�5e�>���q>}��:����>����ŇJ/����S|l{"d��e"�&n��j���5�\.�qωM���]a�`�f�v����<���Z)$�S��7C �@�_M#高j��A�����=!��+�o�r:�U�oD(�2�P�Pl�Oqgu�\��*����;�O���0G��b�'���4R��&�_&j4ǈ�`�4ɤ5�!�z}����]�V�v`/�=Z�33�a��b����/&`����[�'��@§��}񹮜��n&���nOM��fkr�PU��������7K`��g��L�I��X�
P�S能�m���%�D�#�B�ӐO�L�u����3���/!B� %� E��'>��T�gc��b���Ӳ'a$�,�:���z������U\�I�.����~�-��(|��Q)�Z�,9f+Y?���?��a�0{\yr9HV�pO:t+^�����p��=��U>\�����T�?L��9[M"�Zg�#�(ɀ��]�Ē9��}Zl~�40"�̊�k��'_�X@�X췦�1�	��tx�Bc�WK��~�q�C d�$���c�L��T3Ս����NU�Z�8��� ��q-tߺ�C�_(S?��2j�=�� f3����A�Ř*i2��0��xx5�9�w�~ec���<�7.�S[)�@���y{�Z'���1}G����2��~���#��ۜ���eQ��=�᎛�@�|ڳ�:$�}�Π-5���1p� ���9H;<�=�::�dJ��}.[<�����5"3M���%�H
G�xg�g��pzMn�,Y�H��D�1��v�B��o.����;�2��ք��9�f�@�B��ǻf!9;,)]G�*��Sa,�7s�R��;wM0����9���ޡW�6�{������m|�X��L.��,��xYs�މӔő�`��Vo=�oH��}
�B�D�ⱪ��N����/� \M����{V��L=��6Xx���u5!�CCcAH�AAP����՞/��ݛS��e���q�G��~������DvF�·Y?�Re8�͹'\��9��	�0>�,\8��8q����X�!D����\�U��椡dK3�ǩ,I�������X�H�x�0�Tn���|G�:�^�:�ێUi�3�yeYƴ>��&�*���G$4=����\��L`��a���7sm�@-D��.��`Z!rR֐n�N������$�t� 䄻��J~��T"˫(L�wN31t�*f</�P�]�Z9�A��!�(�9�Ey;K`�����&�8�6q��
�O���dt�oP�rs-�<5˽����Ph�(A���]��(ۃ�,���J����b�ڟ��!��~��d7X�v_���@�p�����u�4�ڈ+h��Xh,0�=��c�*8�Nq��4���7���j�bRS<8�*�"MC��U�wM�C��K!Ñ�"n0ı�@��^gW��\{��M
��8�)�ʓ�'
_itw���x'P�I8~
����盍�GRգ�l$�<��3��=z�@��\h�ȶ{�����b�[�Bm�Q
�`ݵ��E�䒋�-R���4;[�P��,:��g��;D@ �f���e��$��fi�=��=�