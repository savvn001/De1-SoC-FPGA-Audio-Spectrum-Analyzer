��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	)Z���'in���v`t(�u�ʗ"]>'إA�����J��Af\����8�6"��XDd�Z^r��n��lUG��>NBK��e��K�ɮ��Iꢺ��/zDBG�tuT���a)�dg:&�s(�;�+�k�k�^$cg�]�_v��p}{1���AȚ.��=W������(����H*(�����p����n�BT�9F���ZIKNsOҶ���w:�A����_�ڌ������zt�U5��gU�ޡ$��!����nʉ��~�n�`}ȓ�	ʣ��i${B�xAi�w�$�fkk��eL7�V�pa �5�N�z�uA��>�;�C�&Y�z-4�I�,���K��=G^��@ ئ�J> ���7.��LB����X�H���
I.��$O��T�pt�`@�ɮYg���BYn`�J�)/�®�E�q���մ�=�[�����P�IU�����_0���6�Ya�RT��d�t�ܚ���c
�8{:'�������NvCK
ג\rCH��`�2�_g����]���yzɶ䛴���^�A��-?��$��L<ve����wUo�B�܀�_Q+���<SBs|���6��_6�ڷ��?�t�����*���I^o�?�Q��� e��gy�z�����fG��u���k9>iM�rqt`0-�p)����x6�pm���I�e�W��p���0��r���Z;ÈDA��Di�-�O��՜�Y�`g���b��ak��_�e)�b�鍚5[���T��+cB�`ߋ�T�*r�R� (�2uGur�z�-Ў0��s�~r���r{���V����]�VJ5��0X���:���݊����X�ㆠ6	���*����c�c~���IC]��h�c���	�g�{{r��$��E0:���
�!�������,�!pf���A�W��E�:�Ol��-��h9�Q�9��ȶ2~���>{�[ɚ�=�(Iu68\U&�q�/� �0�}ﱺ�C�F����N@;[�	�u@�N��_Es�p���w`o�[�5t�j�/�u���|�f&�0|Ua����S���J�]�7�$3g���fg�'�	����#e��_w�lNG�l�����N'�E�y�S����_�}鏟$6�֯$�BM1��rUO��
�w��<�G�9�z># r���k��5;�'Ŭ�̬7��S���HQ=�_�"f-��o
1�뼟̆�KlP�O�>��rƶ%����+��2,;�I�8O(��{R��>�z(�A�-�p�wr��vG9Q �泙	�s�GY�Q�*�j,��Iw�S��d1~���\���@�1���`V'm2�����jo7i�Z\���~8�C�&cў�t��R�+(���U�05Gd?3�DV>��8@�P�?�U�ᚦ��w�|]x��m�JJ��j��R�D����0;�7)���ӥ�*.ZLpD�r�k7A����}X�N{���` �j��/I�� ������� 2�l���:�w��
���!s����{}�2��ܔ]�҇�\(��ְ��KL ��v��L��)��6gwW�wؒ�E�PX��c��
��U�Zrk �j�:����+OE��D��Z�Q�Ȧ������*�g��!C��AjX�b��3�"]�
��4�#y򄳃������2�����6�Z��1���^�p�pF"S��v�/	�B/�#�:����\3����?cݥ=�R(���`ғ����S2T��v�SV�O��ԎC6s�٩ܡ���B?��E�Y�
Ԑ4�b�۩5 -�ufRς��B)l��^+eIÆ� �O�%��K!\)`AG8`�]�j3�ONх�t�{�|�����4��Q(��H ��4��JΡ"9��~rJW�J���fE���X�غ��S̔�
o|��?��J�+T#;
!e{�]Hnۄ�o�\��҇��1G��p���)r��l��'�.?���w����v7��.��ψ���ޥ�u�E�WZ�Eq�����&_��Am��z��~�8���I��T�:P��M�Q��'&��rި�b:y=ٴ�1���UϩQ��-JJY9��rL���+�IM��F��XU��6gv ~�`sh�ʄ|9��Εf�oyu*-����tPA��v��<�� 0D��^�h�����0Ysa�̘�j���1-�n�#y�f�\����B^-[z�K�{"�~��?ϏM�l���ԛ�w�PGͨ�$��_t��ԭ�ork����q������GR�1[�X�8��P_�I�j�l�sR�ȓW��*���	2	��`u��}�9����A����׊�o�]VY���D, �e_}Ʀ��'��<x�:��'�KQbU��F�Y]q ��N��N8�1�;��~�$���4�VO�6��1����Y����4Y��Ā�|��m�A�5U�E+�R�R?�������3�\�qQ4�GU�~t��/.o�P|K�D
Iz�@̃<�DAc%}`�L1�
P�钺]"��y�?�{�bC�ѫgZ��C��g%sP�5��˦�<n�{v�o�HH� ��r\dl.� ��.m?��b����B�@���f�A*�a�I�]�~�ݟ"2�,���=�tW��Ng�磁=H#����|uU;���৮��G�!W�M�3�J�x�!���ddC��[��3���=7Հ]6�8z<�m(0tky�4�uSCf�k[����_���UoP<���*���9���Ӣ�A	��ʗe�iI,�k}���k�7R���gp)J��k�-|2���lܓ.1�X=임�7;?4d�|�MرcV�!��0��,�����	���1.���9�[�8o����|b̓�c�!���J�e���
V��R�x�郴.�@���ObܷPq��ZYi"ޚ>mb�n+ !����iC&{⠟d�4g��I�������h�,2�47�е���4ER
@�e?���I"3��-"Xų������Yܨ:K~�/��x�F(���wF��v�9l����& �C����ԑ���˷S������X?��<Ȥ�R�~kN�@�W-/�g0n��s��z�8,IA��=����u=EW8Z�	3}��I4�T�C��y!�B���+Zn1� �a�v��[�d���d��f��֌��p��O���U`��\��?5U;8KB�=,n���"ZZie��l����ΉOqA���ς��WeBԵ�������}�с<����.ɐ�쁔0�R:��tk�U�sȯ�����E �/��4Q3n��f��6 5D�?�!��I����T�$1��KE"4������j�ڦ#Xi�k�
7c�,���'la;�)ٴ�l����yq��.?m�~'�(̷��x@o�f��'�ǀ{��sT�V��3��Ѧ�Yo=!�'�c43���i.)��ꬿ��[��O���w�e\-A� B�3�L��O�u���=��+> �d�K�1��<��ݑ��hP�f�M?x
� �g� A�T޼3��j/�ӳQ�=��9�:H�m��A�wؿ��lټ��"�2�>1��W��h>p�,"��Ǣ�m�m5�\6.�sk��u�̜0����pv NOOT�`��7(7��!�.�O���ۚ�z-���S=�R�æٚV���NK)��c1n-|Bi?n��
J0O,��}���3�])1����+��/a�z6w1��&[j�eI�~"gY��t�����FS���%�y���ÝLs�ɇ䄴�P�b!y�W�3���&V�@����1�h<�8[�w�����\{{�� cԂ�i7�(7��q���%��;I��I�x94������W�>�m��>;�����h9���M�~k�	�{F_��ݼ����I��[ҖiX�!�[x������F�n����S�<|���F����ky�*�]��W(r/B)�O���þQ�����F��$���/"�ႀcj�B���n�8�r	z��h��+˷$U@q�ƞ��z������lU�8���h��*Aʻ3�?2>����V���6K�!��P��,T�!w���+E�KT��^[6���:A�G9/l�������h��X�*���ت
�����
H�����Ղ�oxu�*��p���$���QM(�i.�e{����!N?����!����˺¹�`a][�O�b��zmd-]FW��O���e���z��~�?Y�o	�4�R1�	��ƭ�t
�����.��ߖ<�I�s4>f����M�t�+k5zG;N:�`,g��{i�,�jb��� [Ì_�/e��T�����kp�SlC��K_�C�0�T����S��@����s�ĝb�x|�/U����0�z�P�b�C���L<�"�.(���׻6}�"Y[]�du�� S�/��T������(|���f�hF�c}�5��(��U��̠�]8���G'�{t�#�� �&ƣ�eBS'���^�=��\Jt�	����5�|hd{�=A����:}��:��p:$ɕ^�w4�o�迗{�L%X>𘞛��e�#�*� r ���8i���;��x�N�����'��<���?mj!a�� �\�;�����(�j�~t����6���č�.@D��	��3Ť�!�n\�B����$S^v�@�'qԺ�]�3q�a:
D)������E��ބ{���se�� �H�t�,E�?Jݙ��|������� �����F+�"ש>u�{�6�,f��\7��-���0@J�`�>h���3P[��:6�߽��ej�0�Be(���]_ܑ=ʆ���Gg�݉��n��m��ڇ7�������]�|Wp��*��f��+���9Ej�_Y��~�5�+:�V��|��-M�"� �܍�:�)�8f ���˲�m���Pe@��߬����ܓ6~��:!	�r/�e����gW���(�6*��lszf�3hH��%�j�a�B~̻�o1�GL�&��,B�T ��������/+<}G��xW�a��(k����W[��"�C�!��c����>}t��r�^�C��澼�I+��F+���b/F�`j��8�k�#_=nlk���aR�JP�>�iF� G5�9G'�d��"`��<=�ަ��([�������ռÚt�B� ��>/r���"�U@�ӟ:ԧYt����:��;rY3/��0%u���1MB?��l�%X\~�:����� �QїNy�(2�6Q�C���d��m"Au�!Uǟ��Ɏ7�ܷ���D�b�cd"�gx��а��Ht��L_�TΖ� ܓ�S"^@���8����"y١�Z)J)�X��Āߓ1��Ay�g�?�^��(�۰��2���?x���5Xf�7X� ��>X���=זĀqдk++�����yGҰμ���#1GOi����~RU�{-����l�p��M���%)1p��[	hp����:��uL��O�"ˡ�&3��E�-m�@��_B�e�*X�Ov�[bUY����k���\�e��^nN���;�g7�GW�D���G�-������C����eM��r`�CKg��W*���������na�B����hg��dyeĂ��$���*�@����#i?�]��s������N�Ic|��S�/n�dWc�y�����b3aα���-ޅgWR��}pI��W�|����]�HA`�-�İ���dx�WC�����H�+��z�zA�iM?����ַĀ�$/�
`�O�� Ƣ=&���t�����h.��yIĴZWbi}��`?j��?��1 嬜sU���(Я�T����cլl�pmj���ٔ?�p�4�f�A��quC��/��4��b��; ���	�G�jбA+�S��,ب%��s�}��9u#&�P t�7q7[�V��`��H�bYHO��+ˉ|3Fm8�ۉ��!j���He���bS@Gd��� x��z!POV�����%��Q�'.����~��@���L[R�~���?�D޸�_�~�#E�N[x�EE�a�a�Y(��Q�131c��-��m)V��$Z�P��v���)0-6N_rR����E7$�cx���R����E������"�{w��x�jGu�Y�*�4M�?�q��⮛� �7KG�$B�s\;_@�:_ܩ��,�4e�vlZ�k�HPBU*l> H��Vz#�-�z\��V�L�\�R�5^��4F��.�IyN��Z�)��j<i̿)�����\y*��-L�r�xg7����-j���U��|�A[<�`�#
͟(h��c-M�̄�[y�;U�5!k�j�N�\y�Gb��L<^��0���Oq��pS� K�/��8]t����Hq��i�®�5	�w%,$�C���<\p��/�N�7i�_�f��݋���D�Q�pͨ�O���"��!9�M� G�x���M��?LD�e$N�,*	��=�u ����17�S��_��~�mG�VG�ϑ�P����!����U|3��Z��H�M�t��Z���N�L�&4��u�Tf��2;B���*�(�
��x[u�|'I�jsaR�u�4����l�0�ެ��\X�o90�ȫ��n]
�4 ��(��e�?�5�%��j��R����Dg��RHZu��!.�̢��9{��Evā���wk��f^D�s����(E��O��p@W�0�	MI���8��������>�$�Q�u�=��<h��I-���rfP{�7�ʬ]1���7cQ�%)��I�v�.����K�[�~�3$� �����������Caa$c͹� v�{mր��d��s�XM���V�v�gӎ��q����N1�"'\f��U�+ayʐ��yX��i+�=��!OO�v�a��~�U����t5��*���&�%h��۩B(t���C�nn�Dkhf����=���fM�f����B����%�5I�x�Kk�:����o���"xEtƌ��{$C:������J�qM�"$HJ����(p����aG|�<������|N�:X�#(�Gƾg�$t���&h�V�wS&��z��| (j9V!|�b�W�s��`�n�@9�S�5����V�j>c$4.!������t��oCV#2�gÙ�iI�X���ü�a�[K���ҍCo<�p��t�u��VF2?e]�t�.���ND����l+���?ؖ��h�ڬȥ��19������y�"ԁ	5�A��Ƌ���V9[������V��؛�_��
���q��a͇��䂈h���5"��� ���](���V-��Y���Uh�?j��4T��� ���%|�(HQ��!S�q���@�T5|�H#�.DΆ�/xa ۟{3����sfO����]�� V�z�� i��		P���Ak�Z����Xyr����\�G6zV_������m��J�p��v �Z�N���3���FF0r�qw]X��B��˶������Up��}�2L�[K�x��=(�#U�2����v�N۩4��9��#a�;�I�-1�ro���ݐ
a���{Y�'�ԓS��e�%���<��H���v
C��um���H���W��t�r�i����1,�@PË�� ������/�G'�CF��w^"�-��Q3������/%`���ݩW�[^����V���N1�Ŕ���-I�Ta�Q��ύ��`ӓ��Wڤ5X�>9��L8����!ɠ���R��ܐ�0�2?_�U�����]�lz&n���m�m�:��a�R}ѺH��e�rZ��AAыGX�׽��;�J+�Nh�`����j���?���Y%"im�5�{�m�);Ǎ�H��	Sັi]�rT��F�!��)��W�c��a"AA��M
�_$�xZ�o�/�0)�tU +�7�ø�� %H
�M�0����؇s�R���׍&�iYSIrL�#�C�wbA2��UHP-��/�G��NfW�����QzP ���vQ��X��C��~/��sƩ�=�+S	s��_��0A�3}�`ܞ�'�����3e�(Ibʺ6g
��A\�L�s"�NW#XȌ�t�ue�=��ϙ�>���Q�B��������Q�$����$�pt=�e,x��F#�\���%2���Dyx#Gۙ�p�+�qf�-.��CE7���J����,iXX�iV.p�D�%}�~�:* �dט�u	�C^t� 9,��7�kV���4[�^!���Cu���mI��I��JFb����<���I�I-��4�Y��j��L.�s؄���R�.$/T��X�Ьiɻ�|��K5?_�TʘV{�pReQ�;�<(<2H�3Ꮀ����"���w�M��IFA����[˥�����2g�C<e�.��phӤ�Om�{�yh	\yg��.���3k	��������y<��'q(�0Q�ԣǈJ��1#{| rQ�-_��G�gM�+�Yφ�;Dҫj_�$�&�K��w\J	,���4��3�&o�Ɛ�}����=�A��1�u��/�׊���j���+��m�q:]�t��<��<���N�v��4U�4+E,�p�c��q����W���Z�Uc`�A��sߎ��_ z%�#���=9O���W&���J�N�0h&:쪊>a+�����Q
�{�qh�9j��f9	� �Z S큸6NA��1�G��|�����_���pg��ۍ.$�aҰ[�A�~b|;���)�@�v$��!.@چa���B�1&�M$)�Vo�y�Y���[�f���K��}�`��iYV"S>�H��up�DQ�"����8��x�.&nTv��0��J��qU���"h�_��ѓe
]��}�Z\���G���#�&����|f2'������X��p��	��:�L̯���2-�����
zs��[�#�ǒ��=Z���}B�R@��|q�}'�a{d&���9�L�8��Ƶ������Yvw7X;G�>��G4��A�G���uYt4A�jB�����p��JS��
�hƕ���m+�%����+�l}Mt%�����K=SOyA]F���⮎�s��ܬ�2;V�7�����`�"�["uY�H؊R�����>B�S`�)�U��������4�R��k��e_W�='~@���
dȳ��)�~Mrq��뫗��:B��7��rp�4��SN��u�s�#_w���KpE�>�t<���{P=mǌ5eG�s�o�*��J��}c?�&݂:ǰ���+6��u�ʏZ�;S��xm&�T��T�al|����w��ס�Luf?���.{�)�N���s���/��0�M���T�o�`>����!�Ct͔�#w.��m̲K��TM.O}`Ok����K���A�U��[b��%�wX������F[����4�[V�钖�f�dT$W9.Q���p�����mކ�y��0��|f��O�v���z�s���	��#rڙi�
�Q��!��<�+6����),��U?����E����Y5]k:|ޗv1�R $n���P�pe�.�;^�D�|rYw�즡��DӕoՕ��=	t+BDw����)]Ê�ȴ�P��,Ρ�.�]��4�8�(�P���=��k܄���Ѝ��U�R��ię��h~�ꛍ$�P%
��+B�r@& -�X[Vp����u>�!�}�n
;4+1��m}�m����~`-�β��l�#��3oqvv����V�F��^�~H�5໿)��`,��;`Z'�hF���r���
C��!̜�`�!�6�/���b(p�wd�_�&��k�|�)<�80k��<
r���=����{"tZ���0����&�*���/#v�}�>�n�m��Z�l.��р��6Uk�4<pC�Gv�y�����;yK�_�@��� ��y��cjF���GF���.���d[p��(�D�m��v-u��Y��;&/}�=U̙`�@4�~�=��_�=���0��L�H�w<�Y�|���$S�ء��%@/(���[�89U��:n�_�^��
�+�%��` jq�P�\�$��3����\��J9:p��E"�|[B���jp��]0p�u2�D�(i�6a��n�)j'd/[]��oE0W��GUѳ´��mY8�#�(���B��Ѕ'� �$��(�v�d@h��I�):�Gכ�Ԧ���A�`'��~�P4�p�ë��+�$Y����d�%y�3���jsr�[�qx\(�GE{ܴ6FT�ɥ��=�?���'7��Z�'��W>�����1�6LC��`H"R�i������!��`�R�Y�T�\cܗ�O�,�KGjE���'f�,�C�j[�#�|(�9���+�� �Q�r�*1`���o���Q"[���	��I��b�Rb�*||��?J�{�Fq��B�g���·�$c+��8�ě�ܵ6jн�O���rٿ��`�[)5��Y��2����k�렎~S�3����N� �
�
c�QK���M�����ʚ�T��(;O�+m_	�J\0��Mk���i�0v�S�*�9����d_|�y"�g?%5��֔�r�z�Ū�ҭ���}G�Q��_4�W7g��#�q��pk�d���A�J,~	v��c܋8��0�H>q���&�3c��P���D����{�k�!�b��v�|��v<;e��##��tE��Xf�ٓ��+���ͭ���l�	�T��� j�O�3Jw�i�\����m5PQ�0܂�{딹���oM3�3��Ժ �,��F��D�sR!tŒ�b}��Y2[���Ʒ�]W�q�A3Ϥ��������/TC�U�P� ��-S��)Ѫ[��$=�~g��8�!6p��朩��ߊa΢�O
_�f�Y2�-�ū��ޭ\y�;�ɐ�[��m}ۀyY��D�!�B�v�+t����d������F**W�����)�%G�N�_�~��V�Ԅ����.�b��I,H���B� JxLԱ�;�R@�D��8E6�6լX�K]s'�
s�ne�d��l���;/��w'�y�Q'�j��J{E��htB�He���b)�.��gcϟɍp� n�|��{�1�F>��c��k�]�qk3�D��G����mQ�J ��qQ�a�
YUV[
	�QQ����"yd���X�K8I���S.�?>�U�_���g?	�{����@<{rˈ�'�Q2����:�e5OHB_�:�PVJ(�Jqa�>#�'�XX��A&�<{cܛ�2��8i��}��c���	�ù����C�wb�9��l��|��'kP�]0eo����@n֩�@h�H�i���C�m1E��*��p.`�p���o�?la��mD?܋��<�tf%0��P����ᒲ�5�-�����=�L�էͰ�L�U�[�M%a�q���Fd�7l�կ����̞�E�� =Eד۩_�C��� �sv��?y@�0�b��%1�ʉ�J\l��¬�$o�ҋ����E����xw:�V�)Y*��0 ǥ��^i6NdG�`��)k_�_��c���V�2AO��i8��KH&|���3MR��