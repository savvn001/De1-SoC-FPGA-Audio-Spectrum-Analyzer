-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
02h8L9tx7ORwxnoXTu5PIsV5izkdG6DEZCa3nyRNgF3fOvHFyXNcx3Y7vQw6f5DDqj6D5LrX16Ve
NlQk3jAf9s90CuP+vH8EPNEDjfZiWKGh5VDz++N0+Et2gPeBIYpas8j8UGhGLDYdPqHulHQiW2mx
XQfQcb9pMW+A36NDRuMY/PNf1H89JVER3Izv1R10DoyBn49BmOZlHu3LInxGmDrB+dwHt/8yTk61
FMaamxxGFGMs32howkH6HAKe0MET6J0zkp1Py1+pVpW8dRJL9s/3XeRlab4B0YWDCU6Q9dCe02kL
J1ioYxC3rtclVj0GDpd6+2LsIMZ7RakYVczYMg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
dozqCpCwosbRAPYfJqg7qiC5nYq9cqSdAmnxPFZn7F78WDOLoJGpRYsC50k4AF1rx+/CKd2o3XnZ
GN88+KeHfhN0AvcVyq4CVUta0pYm0mntbja4EycDl+1U5eTc1Bb4Ppehqo5XBDnho8/jEOHoyKUf
dBRUwYAdD3stKgqze+Hya25+9UjR5/Pqa9rlOpR3fED9TTjWENMwab04iyivhe7g86CkDVfuX0Kv
Eq4JxLEXu+ul4RUGNb4c58ZPmDdsJu3gpGM/fkaKukUPGF7+dgja7pB2Xpf7tF1o3OA9wx1ijsRn
QJLNfEhBWCclejUQoAFf/HK3ZmUGIcu8gSnwz4EravahbzqFgYIrgh1ppjTDCFeEnc5KIMsOGpnm
FjGXOKWeHOMMdwsIkg5zcnTo7t5qwBPygGa2xMuqy9orIc1xuHuEmRJWwuKqRSf98Yu1grIPOveK
vXuDMu/82f03Kvi/bUP86cfvNTKqDB5PrzTGzFvIrGADoD50Q/rr5H6ewfuKE5Z+6ZlRdGP9dshg
N5IRA7sNsMW1yoBUq8OyM21qrKV9GpT91dDI4mZK6Qz6Mwn19zo8DWIxsZk9nhs/gCLibNGwf3k9
CY/AN0/6UnsjcA6nIHlmCkrMEIGNGYBGkx0AfSOSywBT79lMdz/WiigxjS3WDNrxWGsSUnq4ntQt
NScKv02lQwe8INqarniBHVQEy4fvIDRB+AAkyVmda1eFZwXnRDi1bGi9NzXJaQmvChbu+0wSoRBw
FLnuOyGW6mszM63cdiEgzRo3tLttKu0q93xX/9j3/hA04wiDo7qWOJaRaq6CkeBPeyCbHbtj1qED
rn1q24XS4KMqu1baZGFA/HBlXSjYHi8xRPSp0ApFWvaTHZebNeF4AHqpNTg30RxDyzWANZqUWhrq
RRXpOgQi69F+tfp5mGc5KuxqJbNrDQpp1AANIo+elraieqj7+2mt08CRoM+YLMg7AcWhusXYG6yX
0L1PpJCUaDRaL3zwISzV/1TOXKs20B9RL2jGnVgvQqlOh5MB3oqwFYaWjej1EGwS0trbFLzPlJ/n
RwkS1TUrlniNRJDLphFEcwnUiltn2yEyZpwBEtZhZeRGV27sK/IxRvJ6zOiPNR/VLDkLRDl1BiWM
dzIycOCeJ4mhwPNqjBTFAgNXCix5IuGV+AoteKOILT+1b+ssT7DZBLFDa8YmfYnurr5qrzeDau9D
sYn/aMga0YZUTpTk1ct263yMIEQog58Se0GUR3aWwZC8Qo1gT0YIhaJgGi0ODFsVt260CTUxcRAU
jT57l7qqpAL1AlTUr8rKeSvsMHw4vV4/qi1Rs+DWL10IUILsDvFowG4tTTv8hIFXIh2LqhKDt2VX
DF9Fk5Gofn6D6Y/oRQeZB0PDG3M+nvWwLR8ocqxGaF1EfXjGQsrKAzVFtU2iF8F0e4+4fTIKX2o4
EExjtn8sBzPH0HDBCMVE6vjda7eGbuPfpgCV+NoqRqAgTkMXzgZ7yeN5UVkv6eGmR8RYtsrYX68M
G2OgTcouy86byXH0tDVf592Nnv3lqf8T2gttZoQxBzR/PbxJp7972dKXQdzwI1s129yiVn+slMJu
2COR9kM4uo3TBJn9GQwNqY60CL9zXrcuZ1p3GihM1W+gfjJQnNZJ9iAZm/8FLMSmpkZLVafTUjVs
aGuxxPF2o9vkkCmra5iIdcO31jqYrMsnFm8ZTzwZiIdczUGQtmhlBNJ3NFqqp6SDQ8EHziypuqt8
vdOrqDOg5dExtyW7KUHXbB9OAPOjdamEqfxwvrCWa3NpMHM0S+qZ6khfHZd14rxKbi2so8dhIFmG
fkXX9ovQAZ6pwT192rp3ZJR/Xf6psJJP3U6HL9c/zzlu1JmG4HrsfhWBLldPDTi/PAJwCwf7kkvY
rwoAW/EeCKawKI1lxmTbw4dk1zOrxUsLj7fVHvDSH8Pz4dwc8hb2v3pipWUMhBLHB5RyRFC1Wbnk
wuknLgo1adC1xpmTM74hkls5km++P/3FgSPiX+KwVMym/tlUlegkyCBMtI7bzGey4M0Sb+YSkwMa
srpGAyrhRytU/ycciKRruxb0QhEZl88ZCjyc571odWg2W5rvmrm+jK58DQeizyiAh56jDxcBTiA2
L+o9Inm5Kb/rO0Eqmcu8EgDPgGrdBnX2iWc422+Whn1ollt8PFMjr0GinCmFEE/HXVd5femq0YKb
A4TiNEFkzXhPGS/gVAS9vSbKLVdM7lJuOx+nTit/nR5eX+Ju2COu+2ANEbJ0YNMhz/JrGh9iuIYp
LrknsHjwUGMlZjxe0vIQsnP9aCvK1Eisk1CVEVPCotYAUdYbsFaP/CdhxO4hN10iosmVkiOp8DLb
13bEWHN++dS4QhYNssxZHUbO32KdyKc06VuuQRWU7yiKuG+NlGjeHMNuI3onf3XW06TJeF+fAIUs
kOdadF3uK2coIVPQl+5AQI91k8DFafhrPJa2e+JLIgyUiM3KxHyyNwS2hg6yqqw9zHEYvwCktB/n
7rvfwd64JZd76FC4bTpyfgFsNpCwGijVdItF+vKu8qIof3E7l7IcJwG0VMKK6j7S7mlNYXqlV7pB
zfNhr/PjFQos8ws+enhC8bInAEHzeuazDM/EOSyj+w001EV/LbW9e1NL4EQEA4dPZYkTN/qcoohH
6ILe5KWUq3N6qBwuyVVGs0Xg/tcaqjaHTsqKL5krnuNwDcX8bAggRkWqikPt6CJR5TOy4o9B+A2E
uqDmfBnXt2v1KWOcmZIN3E8a55VfseTRTtDhF9j2TVI9TySN1esog0xezMW/JkpnGu1SYlWEv4nY
buYMRRJLk3IVITU+p7iE52s+MMwKW5aqR4+mFz8XXBQoR2QP75wCxFywcjeIxQaJk6Rml4fg9Cnz
Nc+FySJe8Kpn7UFKgT/A4hWFS4+yIexm6q5tI5bEuspQVb+cFfLlT3mRqesrknmZ4f56ArDKRz2o
8chlMKGoxtdVlyL1FX3Mr1ZVEWIUYVEO6U6y0MLB46/ChXEtPNy/DHxfB9ed9wO/zRQyc7IKSZKM
X9/mIwHkgWZtbqB5QzAFViRpH6bZcc+NqOs2mal94hfvwe7dTMtbiadO2+dsRaq3bvigskFaQk5m
jeX4mYC3Xakj3o1Fr/K0c0AGQzvrtllfOcxpq2irvlF3lJCx7MDGRHc5Py7C8ykXwYrcs/qlEpgA
avggfHxe8FItZb0f9W5Q52KypljBko/fW9gpdJ5lpbw/DaaLw3foalWe5GICgGTXzTIvRKBg/wEV
rN1dg8dNz6BQ8Ocy3HhI7rJsEpCMgmaDklaFtE2xExJFeFILIGCa1DzQiH6HEY3tZ1Owk/UwbFo9
bypf6gOSGXsW4w5HZwhCrs8z/0I2SIvsHY7Xu0DUI0jwZ6mYVT4O3dnTI9rA0eFLGS2AZblKil9m
sb+GWxk3HVc9unoz4fzs/Gj6tdpOnv7gBcsByf/ZL/VrHuyzWLEIFCEUhdJYTbQ53NAeQLs3dg8Q
dAEk94mJXIwAgJN7GTetNauI6d+ypkEPzAGBhsj114w4j/3UqExIdSp5l9b1OPp9n2T0OKrsPevB
aeM8B0zc51t5Sq9lgFCkKZZnWt7PKEe4TXCxawhyaZUZSjpX3/tHZjSxgn2sNW5RbM5nq8ulW8rq
aZhZhm6cBHccT8I5N62I8wEI7Ni8CMSsHwCVkVaKZ+cChgO0Dbmhp2R1WfD+S1sSF1FuOlrmacP+
l1CNbwxcjVckab+sElYylD2OTiC/zDMDc3dxMI+tfxmchqyfxQ69crWfQaj1KSpLJZjYPFxgBF5v
jYo+FSyJ1donJb0Re8Wa7OSb7Xl8p3+di4xvMXth2v+6w8A1D/Oc5H797eXbeMfgf2dwV7imH6O3
/FA/8jToLxLLAtHmze5uQ0rZ2n+MXIuoIQASH0MJ49qzfpKTIa6Y2VDRyRpDFXEoZRkWpdejXe/Y
IUaGz+k1/uekgvZvrfj+1NxnoqiQf0ORTJ/9fssHK1F+8tTjlWOABh+P4xw5ANHel5mrc9ZM/ZAX
77UlGeTT6elm/9B8h2PiTxYomZovFV+rDonAsfITeaC95aUN3NiG62+u2fw8CuSnRWuVHSPMRO5Q
857oMe03Px2rOlrAS4Gc9ZzyQrD7ZqrRlS/OO4r6jLEnX2qUWIcAyU9auSC8PhGsPyacl6qTPCI3
tqHKEM8scWPTspYBLuGPHgwk3xynKByXDN4QbCQ9savX9rw4MUNloBCpkse0lGbMCOvS5759Ony6
wetilzKCJPHuxpB8f6A7VHI3DdZCUVoPGwtJQtISnR2e2QEq470KQ7SzTkt71T06DNgjiAGLZ9nV
OOlc4pm1vAjZRj6nNIn6St1eDjhhERc1OXWMvJrWacHduXZ+kTveZp5x108eu4md1mCGSCy7Ij9/
SSRTuueJDj16gPVV00/z1QYKXF4v2lCfmpacOcRT+xNXM15xFDTsFjzg08Mrp15QW+ylAm/OaX3C
cqlEcShUo99sNteejmkVorIuCzxucf1ch1Nv4GbL9a+Kpf619vgK0uLhgsa12Cs5BBNl3cFHocSv
cxi4eKJ7L/aoYJg5o60v5LoAH2QkM3ucE2RBkG1hItk2PqljGvQrWcSWk81CRobcWV8AG3wxIymj
SVM8M7l0BEazmZNIeP84XOw9cm7FGQgxJ5/FprEBcVgonI7WOIYxeBLahxNVjsYzzyOzJJomVTHy
2RLVm8kgxB1UWXs8OJhQWy66FUm8w6YPGtxjYv0c+Pfvr1audRnoAfKjtbJSBrnJdfU+7gJMJsff
f51e2v8nIM/rWUo0gx/Pl44TPkeIp6CeECHydSWOfKOxDyVldSzPXtDJzfvKDLEOYLShTw+eXh/6
Nko9bY8nEJFXgkHiJ4DauCAmaA8fFbN7wxrWbchDOxCEovoecm9Q3ZOvfbqBZKAQttI5b9/dKwGd
DV9bLzJ1I09WKvNHCP5oKyoZX42MUO7pWC6/w8HjRSX7V30zV3+d/pTv6pfp+8BLZW/DXzM7Dw9C
Wt3/XqiQsoPIEKRg523YGXQUu3THxv5UbPdKi1RoqNp6T4+cbM8waHV/VXCuvkE/N68Zv/O7L7aK
NJnuUUg8dwd50kju19i0Y3TxDLHyaZx38QrS9Vtcm7aU3SEO8OnOiA2qoueLEJg5bSwkR6GAH1uj
z+OoH2pA+ntDXX1VQ33+XhW75lRSN97mWKs10/y3eZjFeovlwK+g5dODBgzzEnphwQgdGnYMBods
ovkka42TGf6yp8pdegO3HESwlIqZfcFWH8gbiTYXLvoYB1JMeQSglgT7raM3Fps35XwPu+Mf2xVO
8g4w2vvwSE0pjdbzhN2qu9yiJk+BGslEg4XiJ9tppxgzWbXiQWW+ZwaJcZKRoUlRh0swfClrzRpP
nft710VF684kkUXn8u/RbqwoAMSFGd2mzCbObIN4aCq51lEg0oX/jWYFFHslf+jWdofMb+4sfQMi
/M/EMOMVwgxheJ/0qRkRGUTDs498Hyyol3J52ApLsEWJVn7AgBDlwAtLE/gSKKgxY+77ozv2TF5R
RlkmNomuAIMe3NFBh8OOokQpJXuiFxi2HMUVMDEN3s8ldHbJys32gCq1MF0kX/g4PFtiJ8ubzTZN
3fS1Ll5WY/xWvocHXeh/E3If1uPLJbGJ7Juf5vo8MKge+ZAl90K3d4rjhcsQcA9ePihZThodevFG
lNORWFyqZu1pH6G0g7YawZ+d6+MwZ2JlGlerTb75BzXW3PNspvTzGOuX2vpNejD+G5yZTLJb8Pml
LkQYrfjCLgiVeNozimD/VfqoS7e28caueH+IqR02QpQHl+ZPEQvmvTsOJtxAw51dImsW2O17InQe
7rOjAL6FiIRL8hI2hYwqw48D/i4AAqe8ED7379ZTgWuqzmuwBNGGGWyCO9v4/5jMk3ax6AdvQJOA
YidJYagCY+GV3XcHTrfTZnd7o6NZylvP8cb2X+pOijc5hb8zIpo1i3I5S/JJsPkPCwrBEKV30i9i
GbB/UAxnr4uWQwIpdZpH+0X29bwiAy4WnExyHfj7vo+jlltbiVwvYuOmtuHtMihX3cXMUmH/Ut88
z6rf7F29YWiN7xBydciqG7yoJjfuIEgq9c4gXEQG19goAbiDMn1MN4BD+Q+4hlBSFkCls2WeKbVh
rDwoNMi1QyCVt5484DcQtU+DzikG4QgMNUDsvOaWdJa/bnYYiDv78tRnRKMvTE6J32JgddTHorBR
0krnbQ2yGezxBLKZf7FzrS4ChZOy1FbJS2kyeHV+PS414IpABiW9CVqLKkUq/+73wnoyOXSOmjsC
bu7eAqExuiLqVyNWNpl5RF2UYf+UqmFbISG02BL3m27dkKQ1Afcdk1VizDJOg6VzBHdXXlHXl+jz
Jxm78POhR94bPaytGvrj2RYCwA72v+xzGYHdEgVCOlWkT6o+WEeO+wse51GdGB/zk+TCZ+Hd0qMa
rOSli4hVI3G4ytsubmURECUE/ogdXlow0BgXu/6V/gMQRHeHcru41cSFrspErbFIsQlb5pOdmlf9
GOpF+Ero86UOw1BqmnUxMaNmlrKNKCZngStK4HdrY0eHcJaSqIqjeB9ZHZCMdBrM86eot3xpNkFJ
0w4YcPAL963ZStYdR/jjWBV2lHHywr73T19l8F/D9fijy2UpuSxmdn5mvt/708SErPl7q8PBgIki
mLwH5tclpTDV3bkVHTXvewBIqNXO5R+OMi4vnFG3DaIdpPokB/toRTtxhgXUy0fPnXA716zXE8jU
p99l7CIaqEtOkOxMAjQbTRrhastIMNBteThKjRCg+a/zL8fKJFFFpnysq7VgK5SaxHcyRdvbAOv7
i9AZwe+kQ97BI63sT6+T3u7pcBukpbNUxHF3DeNQvL4Si8O+h7ztbRDTbr3epzBwteHSB7h8RUA/
Yn4si86Bwnq6iaM82Z5Si1wPe1dt/O6pAFNKUys1HsdbDnrhetsdr0gHVm/ekU9fMzdNaNu24J4A
SIPwMgJiTalIHtXplT0dC07AOFs/6DrCcL6Tj1vnL7CUIPpyQYtegxtcpeNcqVqezM4xHc757YRE
cMEMzhWmYzYIje/yEl86Ecx3wUXhyq+zaZCpsxZjI7QOxpNzQ37iildEvOClhh97zLQBJWcq3NVD
9MmkUF3fO6mdymK1P/KnOl/NK/bUidJfz3cj+t/IHB977u4cy4hSWTkbrAII7xHzcs3lv9slckrC
3QTWdPb0s3JHdweS6xJopUkZqnfLmsl1zRkZCMlaTLLae/KU2IphwCI1/3gsfTfbuYdn1kv6ezQX
ZzGQvOFkK9dxRxPZUVhFpTof9Sz/VH8WCcl4jAlE0yj8S/UzpZTIxRf/y0pFkVS/ancHvQRz7R+i
vHtM8X9Vygq3F1YgZIFrLxfzA8skH90JkzaXCuReXfJPaCvtit1+gS0lDtFo8qBM1fMNFpY/PPt+
b5iJ+YnJgKz0zTM/qBEhRq55omuOXUwABKnzfFigsw3AeBxeaedrQKtAEpYLNz3xGHZzLqQQVhA5
01U0CcvXlSjuhXjV8yGgrpLFUPC2E296d/lx4U5vykNq0tQD3Y4CVBidXo0b/l97HjO+kJc/6TlU
fxA9605jzLWFWaZuw309BViDaIYtY04iHh5i0dhjSod1kk7mQBrdyB22Aed0fL/7/G6cfi1OwyoA
o5BNjGslvJgRB1tJ5O6pLEfRlI+o7bqJ/LeGEEhhcBxDWoHo+CEbCKnRzSbEuNQvwsxF0dXQ888B
Bz9mlQg4lHv/0U20i/Kqu52I8Qf8U5U3lIq/Ze2NfJ9oF6kXwRfCrh+X3V1M1m26J9OPDv51svoj
dZfMudP9Jcfckj628HCujKXx9Lmuumr68ZviFEctAj+po9Rh3d9M37lsGS9wDNBUDPLIJNaRlNi2
AyjVAykabsEUIzgAFQUwV+MH/VaDkejK4kC3KBqgjohwyf9Lzdn5YGQ7QJ9HCHcLgMDgVoilK0pt
ZaOwEvknPkSuZ8YGWOIIoaR2W2uENahbFEd6dSR90D5GFFhHVKCYgo5RdQiMC6nAQXTQ/R306+rb
W1MUPWf9mbqTa9Rzd2olxFMeEAixHdjtzy+4Pk/WTjRQbVrpqt1DFac5sVMScLvkN/m9cIldPP2m
mn97/pC5j6qfPisXGndXXrV2j3ZzdnFkQcxj6C5eGbbtS08SFHn2JX9Hq4apfb3fH//NOG0wMrm6
V4KL2lsIZ6hG/YRmgPC/b8nbkZ34wq5/+N5E6RSxcUGZDWxFmKs/tSNUCQjiBrHk1TRWDt6rseQ0
aL1SPdZxjVCLxSM+WmYKdI3cwtc8G0btDKUIIwjtxPTBBmyZvadeEWJsCxx/0kxKo+zdSymUwpQ+
CMUT03fLDsG1XTdYvb7DtP2+XoU//XhpYWnLOw2W8Z1KgN+1ROGOsBHxfW36cC17QeQBvuLzpRnt
JMgHIWed26z0k4bKkxS/uznMCcTib2XjIKngatl2lOx7G37p1wsFY2qUJ8184F0HyR5jrnd5y+o+
JSWO1RjrjhCAtm/Yc67PQ0zGmN2PkOisxTxWjOG6XB+Lw5ENnyagC5Aiak9/GXlPpGF6YWo3WQSK
rzgmB0O/Pg6VjwTYDSpaY03OCL+JWg75gEO6CWdpINOJg0Ct8hUONxgkQpeNM5zL/JC0jj3wMRc4
zrs05kw15hMaKGMDOa1VN1rrNvg4QyrAlhRHkAkeZrrA711Db5q4xvJy06RAEnwhExJ5Wx1IfOb5
a0lNaglR/Yaijirxrz1fnBs3S9D9LiXhmcvc9+9XcjrfOg+Ru5M++Ft74KbRDWWc6sPF+vV9iHZ5
r/QdiG4/uNXGeWhHd3bglSTva/kiAuO4iYoHslMS9iy2jZM6fwk50w9FM+L4HvaQ3eQVjaWCkFB+
yoRkCar/8NtOgfu2IMGINi2+wya9TtIPMIYGW7brsbZwbkb2YHG5gifNzWU1qNhJXFzfZDQsTnUZ
VqbUT8zraEQYIMq3sG4ltAC1KqplXcCXNpK7pymODhOz+JZ6Oj/5T0K/4kOd6SmPsEdGGYaqFmJR
645AfRJ3UgF/oxpM5iVXZEgixOAUFC/4W84YdujSI7y1nhYxa6qKbg8WleIGxBWvcmZHBne7qm6w
yX7NUzu8VcGqvF6BlBQJP6YdU9L9bQCOp6LdwPH7f0GbV/wED3sa30rVMhFlNUKdSOpzdoTmPg2E
Y66JcHkd9t67a1iWyq2B2qeb2nePzbt8Hri7tQVOkYpiXtWVgb1mj911eHFAKH1kCzlX641arPJc
f9Po0I9jqnmQJfoYEULhsr0yj3kdW4s6j2ETpUr8wcOlpqbPB8oJgRIrMari6dib55jhPTUKcs/b
qqYI05ys8N9T67FB4+PZHNvQr0kCBvaBKUSXgRF0nZ8ErMyvtSom1SoyNMZ/v9MNbnmCin5mBYE9
ZfggR+lslxdwIkKTPtwMKQnWlGRN9qw7GIXeuMc1oKkdPxXwFQpl0W2Ivc8zcWnCzSYd3D4OgjgA
AQpjnZIgKe027klJYj4qrDGhh2b2g2CgkerMubH5LLpFbil+JMLVT4Vl7D19SstverQ5J4hqts3e
6REVnvmUjk2NXRhKoT/oezYG8itbiAzdAo7ZRpiO0DREy1Be74EqEbhI58NBvMkN3yg5sPv/wOtV
FEUoFc/QwC+R8YAML/6Z5Eb2gttMPYjZH2qSUzaXvu7vByzpLrW8Hnbp0btuDwPICWK7apxB7GsY
dV87rKLpr3n3bd6oZWu0/wh/G+hOyOpsrYG77HyZ7jr/r/BQDggg6Nx/GNsv2YhKIkUQJ9+fvH/f
S/lsTDVIFgC5SDa5NfvEgq+l3XNiQxf1eRgcwSkEExhr6/ZPKygbWZXEtkhZ7jjrdBJG8nKIqDo+
3BGkXaVwep4jCnM4tMwVgb255EB1onei2WPlw4lCGT/HFLhVjwunFhckv/fdPE9uB/4+frjLL6ci
kz+01e2x2EkjV1jvzT/iSoZ/UCn7dFt3rU81nCjJ9F5nf3ALCvs7IImGV2BMd5OMEAAO1DeHsynK
lF952qEuKnbRirhacSyLNKxuBOb5qdQJJInJPIwWsUBH8UyluV0bFI7pZFeo+n1B5n1s81iYbipQ
jrJPv/PBPtjMATaRgstI0/Fn+HiqO5YbTvGr+qDqANy3+SP0Om/ajnbZO5EdMfR0GysN5/G87pmo
Eyd/FQtjvulmaCnRqQ3Q1Ma5QSpZAteRtBRPHPTjJ2P+Brsejsj6ERiQYfXmWvl6g7QmBi4GXYER
gvHqKE/xsvsy6BcokJdr7GCvNuUfH69rf6KdY7TKHTo+XmdPeuUeGjcMu37JHEycLvgHpIsMxJnK
uKi2A+IlbgLRDels0SoI3zIx0JU3PUT4mEIw5VLsEf9riptLfXWs0fq91YntucPSPyujMcCuwOPR
qESFulF/cAGCID15dPd/aAH5PiX2MNfaz66iQ17RGCkSGkjDCGv+phe93nPtiN5qp1UNUwxoY1Vt
Xu0RugObLjAU2xfPpDhGtWu36XbBIdgLeosxe2XTy4phdHNSke4ZtwUD65tvSMV5VK9VITsvCoXZ
NHiOZpN0NAoBd7BDI+W1h5NrhOyJF4ezhe6DJpqus3v0cnUh2L//urCR4Ty6AU+wXwF8cpM9J5rH
enlkpoAM4C4k+KyQkv3ADRcNZVRODKRoXajEZ4Vxi1NHlvh7Szggql0qEMzhd7i9/bw2aP2kway9
F68cMfqipco1uopHLbfOqbVv0TsK70m2TVtCv1nmfnamkuRNkB3xoPFX5dXuCDphNHTWL9CVykPn
l7BITMNOtQeOBLZJ0mi7n41v12bY+2S8SKiKZX/CLL+Y2Gofqq+6cFreeeM20BNwaJPfyT5XbzQz
8YZPsbVLwb2fyLxEajA76hG0QdUyMxFIxE6EvRLgmYbR+OLaLR7rYnhkTGPEPUDUlYQrWjtl1FPN
SxLRiISmgLq2XMgl/1Yb+LGAxuiU9qFSkPYfGZfyCIj/r3CjoxRAOJhL3GdNlB+aIhcG3/adZ/jT
IES7dbEGm6mWjDG+kgROI2b1iaYH+7oyESf7j1Ax0EgesZH7cEEPFsojpi1cMX7nl2NBs+dlx7NK
oirnoKj/Ss2oa+6C5RVh06gF5Bafg4cmpb7ZT2xIwVvTdJg7nsY8AIE8CR00C65GaR/fOgFEdWhS
mb8FAkbeTWvYhNCI0dT7PtlS3Baqv2bMW7+EYLFt4aVpKXV7LBLF0csyBIbWvsj+d4qZkyccWtM/
Co9IWoef/UvuW+cz0p0iE9ZXZ9nTor22ksO5IXVOeDPoBRd199UYEuszTDZ712H90YkXAdKYp9No
oLbF4YgS0jv1zfv2Nbqu2ky3cxPsigwr1IqtOrVVK6oVRdyKgp9JYZPV0wR0bu9UfMfAmag6Eu+D
XBFYXgQjEC1khpbZcuin0Jr/4VlkBdmjrp8FFztbBkLlO8NHS6LlY3EUOBdIttE//ofLCCDfIVOK
Vh5ZF60/S3qXMTMNFVCHILM4E4MtTsoev2+PilEVi/A2mtg8oaeZZz2rut0csWhr4eE1eWDPoXAv
4ZNLbkrUdJRpdwGduVUpnahWeL5pliGYY/PyPP5FrKrESPahhUCKUVUsR+pHEUiUqoMT3l8MtpgE
IG2WZvHZOFDmJMcSCb4epRcOnBx5IhtrwhwDQ4J5igvoKZLTv+45c+HhDkgz+Tk2DdX7i0d6FLje
HvbSRpwd4Q3UCBZaanU/ewsRVHV4AIYsBVopcGDcei3C4YJsiQud5lE69OQcPzN4NYi4ySMp5ClR
LxWlAXLEwYXdIE9nazy6YMJzyeuFhhDTsSAq5P3xfVq9PUjD8UnIzC2BLiZjOqFkvYaYqTUEB/mP
Fdqzl5Liacn/BUf0iZnusRUzEwxlsl+ZA0a53EE1qe0gvzDW9N2UZMRWG0DzhA0gOuM66KmNE9w3
+E7em74ybvZ0KlPTjDvjlPXkGChvJr4BGY1u+JfgiD9qf2O4EE6jVOLXwBX+zasbM06VcoX89fME
YSx/qio2phuRn1tqfM2jNjPc+ihDJCEmIg4sqZ1uhvlluGGQRDNZRtEYmvkEwcQKzG0CKoYzHCUh
LPZBKSK+MMUDqgYPWRkA2cDW8BN5b46qJDM9jZngTiujx3bCqGRQSD2epnFbVoyowJi9iZzKmch5
jrOVQ6pQwfrs75Pnr8zkbXwJExlGgU/NbMG3rJfVv29GbFcD8YgxX/mSEJKdCYXdGH1kQrEei1iW
DJ7LKkofapihTfG7qPaUuGF7OJyPxwUZBIfsABoqHM70u9esgMOcoY0OWtbUxDEbKyN8L4KueLFA
IN1pMW/Rr8MJ4XGIHlIwZdUIwJ6zkoSWeWSDgfi3C3VIfpGUTRUjBLlMeTp8jNjdJBQXV+2T4LSR
h3YuuHO5f3s60CcW8FBZBegtQZS0X4BfTngOJEvZMqrZw2bxFho4S9Fv+zgoNyOyjiz4SqDKCdjF
Apeb19FUTllz/X3BrfJL94bpJcDOs532EUmQoL3PkDF7pbYn/3aTWrB45ojZ81nKVH7VcW4BPBDI
WV+7dZSozheZvzHBxdG42VsNfksuSHkjSOOg4l9f5sMJ0mW1anbPqTIMi1nUqubt6qAgywAStji6
8B0tEWHAIl0YQ9Trz8oCMWKogYi6n1vvM5QWEmaOHKbUZVZicHbtU4ZQIBQBN7f4b2l6iE8U6GEN
E2WUFeufAWJcJXDfsNGlEjWTtYSwDEXDVMWaA9qVgSHA+ewYdfRIu62hE8hoh47fPjSZ8HlqswfU
m6Cnw1P8VdIX4MNudfuSVeh4a1DyDEYKABsChe8kYtbYF4L3txz1LhuH7I34/g1A3Gdi0+R9vaHS
M50gGok2LnZL02E0HXzLiQcg+6F9p1JQAqCxcFc4ILewEmphnvPHwZ7tftKl5dqmWFsSA6dMj1En
f9dgfytsKJQD9SzJZys7kzdlTCMFUzXyBFIEYk/6r0+dVmzP4wqXAJRgaZ+gyWjUvQQbDXM7MlJd
lICF+cJ+ijmyKAh3WVySBNCF6hnMLr3NDFFtJ+ALmI4puf8lHxn934+i3Y7z9EU3jL6cU5YBKR20
/mhliCXLpZzpktvrWv1TeOH+3s9/clCRMMzPNTZBekTCHJ4+TElGNHs6BPFA9DomirD9cnF8+0rA
fryZzN4VShQyzokyE6tk8DuZHR/3XyG6nGr6RHOhh1Xcl3lFMLR0uWxngGJWXh7wsKptiOwZjynL
0mp9Ri26Av/FACWO5YhI4nfk94Doe8N6pwDqKzokO0hjZKhwZRlKQQYgFqhd9wiY9E0XbaPb99hz
WnlYKnX4ubi70Gp4fX5CbSIs51JcMRfpK3QmBjoROd1wAPCZBu5dIzLvukEk1fc9zzcmx1F/hkhv
UNnp9Fj+DT2JebzBO/W6nomLZ5Xj9/gYww5RhjY7HIC67cw8Kzq46u16g4FfWHtJduiopMiAinR9
LntbtA6VhKEg81qev3/hVflTWrleaaKPNGyet0eZBHRqcGpqw2zA6eWyLL4TYDQ6XjXknMqrgF1a
Tqt4xXlUaISoVHBAGiuUNK7Sebdx+oX3f1QqvUNjs3QZXfU99fE6Bgu0axWOcAK4Z7G74OpCy6XB
KcQtQ4KAaJ6glVFP6Yez7vGQUsSIBqFcHKCln9FjyOySVBzO9iTiWArw0f0kro656l0yMJdSogVZ
NhB98l1Czji69hLDmVYRRJ9sPwyC6oPDtTbZ4FMG6c3GHKrfNntQK2V33G8IEDYzuwFYFnKXDXw9
18MPS/FNU3K4qj/jKk4PTouHjcy9BmughGE1C2GJfglbK8EEbxah4DhVfRIrEhr/c9510N53Pef3
1FOQDQk6I9WMoUA2knQ2symyYKVx+PQFkSCyMw+7MwgKCiTh8VbBIZwrYf4mCMVzwpy3cEHSCFJp
1wX4x64zUEE32LMJUwtFr+CdD4bjj9HDXa3E3C9vwJIlZPYtckIW7/dDx2V1kKKlZyxMerl7SS/D
zIAoz2tVatlhpLYP5SgtkgPU2EKBS3rMTRuxNCjpIJTUUQZ/GyK5Scr+su+Vs/DHBdNGof9dmRpM
g5rDf33o9Cci1I1ztNWv2u6tTprwVaECoRv/JFjst/pkq2jk+Q3c7Ur+ZMj/yVn/rTm0/VznrXoz
xg9+kvszBqx2O/iKEbJcrHL9WYJNSlsfDcc/O1uyhXfBWXJErqxBHRPH+1zaT1HGokML6eyBqqax
ixDxzO4W9aCxFEVq5ofh3fhJOJS62RaSMmGuXTgnqxVz5nh/7ruTwLkZlKNv+E9QbG+rdxDHbXNM
9kruD+iTt+MkGPwaile9R2qL+zOEw7ioIYJQnH4t3hfWKMPsPeOHZicy3R+vx7GylSUfhpeHbOyQ
j9uB+ApVXruhAoQO4jaTXkbl4Of7sbFTxrFOmD09UhG3AO9ywJp3ag9K9DWkoDwGb5VwgHpeIWyB
cED6GtwAr6ZES5necGnKtguFS3i7VzfDeQM6zpsIYKax7cIVszeIz+JFbEI6RHB+bq75a7tys1Gd
xvrxFwbNR9Gpg/KUr3oDq94Rk9cOlRIVHJV7mRYa6Ob3o5Nrl1s/5Ug62keWdPPTC0xLHVYDHdgr
A1SiB/J2HtLFFKZK4vKl46wQrAkpljB2e4GOPMBYP4Q8cYfxM1+kEAtFNRPJVsNwskPzHqj8Lbdl
rLIgZcuXaswVAZzzo3KPd7uwccbF9tWeMMNkZ7wpdTD/KTU8Tbsz6V7PAhpIUKAzgw48V/cjcMxo
I486O3pSUy17gWuY2Q+Ls8r7Oyc99R7+H48OJZw1ZwmVSWkueQ6xmff6z7kdw6wiK50L3iI1KC7m
fajGeOdrg7ATa8j9A5WAuNB2G9WHUBpRtiNaw8PEanUy4Cvm0NiYc++FxS3NeRk5G3ts0c0pxvs6
UNZZ8Q4naesDH4GJ9OveXRV3UrrlqPToHFdmmpoPdCwcakeiS1VBBeoj++2tqceLpGOZ+kCf+wlI
kguITsqGZRZxbqwWFpe+YXW2iDgFH5EJpeBUMf4ZJyBQ0hhDNg7TO2zsvfoAQ01TSrf4i+6JYiqE
ANEsaG+9hsMGLs1Sny3f4/yFny2KmmMxHMvK2hNIraqu1jxgDp9K222Qa97kQ2DTVMP5/0c+6Eb1
w3k1t+9ry9lC5soNh5fL9glgSdIfKFwTG3BwnylM/WfWafV9Ek5eFdphb7JmA/GA7Oz2TCGLPBjH
lXJompUWvtrP3jt6Ba2MZHDDT1PuAwTFr02CG2F2UgfF0LwabGGulXBhkixZq9mPk8Ly7RJlRJqG
NzT3vqtKyBhP/bzeFWdZ+A0avOSuhpm5V/51Ui4WMvTmugpmjz8zTzu36gF70Ded7kHtzlFjJ3f6
4DbZX9UgfRifkcNPJeViyQu1J7sfcyMVkpM9/14ITcdSgR8uBO14rylTw9Y4JlwHaCuasGIN/Iwl
WesRdQw9xSP+wBpL/n1KT9o8FwajftqDqZYoeTrDjGDOO2d/HceCj4xDpLunf15SdLEgDOrovGzg
ax6DUxmX75yzoXooM3jB1R/j6TE71GZrvZ5HiDcIK2ofERo0OS6AvxDHt8JZzRNNoJ7xGfz/5huK
NR8Wkm1so2IuF2MFgaioVvqjda9EpNgfry1Dp5SF4GTp7Y9q7r6F8yHVVEGt4ionyX4TvCrAslDe
jgE2KgQSivhFPv3tt9EzNEVyRkNsNwFoamOitLe6QTVT+g2lER0ZDfgvCALIfWoHD+momE+XV5zh
hCT5b8F9pr/akf//7YOC6sfmr2Mj23A1GeVAzvnqJ4FwC31Lw/P9DN8JIFqiDuP62dPzgbhDNxYf
3/Y1mDCo0luQkJ3m0tubQAxCbB9DnVQzLlQkiAAqHyINj7SOipcuVpJOZy/Y8pOfFAX+2T+my8il
BO3kQPCFCDa092uZqwXz7l7ctYP7oMjaP1aIw83Zgk65CmYv73R8sl+MBJBTxCgtE0OXKVOuaSkf
hj0ATXMTF15S76WEV3yWPYNkU7Sc/8Dym1GDvHHhBMjUJdfdsdREFKaoqnX3PMj+o3bc7azDN+62
aKHfgDZDe31+U2f/X/gdqMiiH6fiumXnHsvtm4iRgHcu+4ZFZNtBCuA0sXm25eywXxfvFcH4gMQM
zkf6/vpgIEIaLdN/vH7bHOQqzFZRmsa9sxJgWmJL7Px3vOn8aDJeG701aQ8rjnH1bQT4fVAnkHbq
88In337dO2zeAuBjn0gqcBsV934rWZCYN6Lhf5iFxShBqQL32HCla4S4jv0vstUQKYGUgHARARQe
1ajQl2yYJCnYcJ4/3CzA9i1bq9FXg6CDK/YtUqUhsrclMYvWhZgc6+juVqAhNaDUDphbTwd/sf27
iQZcR8F6/cQGoJL1BLI3S7tsOQTxcS2+8Cr0P7KxMf1pEz+Yc/dPCL6hiE21WfhJa7B1LJPknmZQ
Q2+HFli7Yqc7Y81jvhAfsXG4eTIK/wTfAea2ecXuT5wmSx2QpqXxXRMZ9zPVNrVAKhTlZRdOmVEe
meaApI+l/NgU0mYAU/+5cThmC2LwF+Dp64V/mQ7y1u1q5PTbwjpXoV1Puhg2NxU0u/u2ubLrgw/H
DInqTFkA0SAVtCdB8wQE84Tj8dnv1QAf6N6nQF/xxDxm7cUQj7WBwrCpN7XHKX4gG+MBjzN2t3dG
C/tXZz/LhOZZAJGFLJpLVKdgNFIW1wZzEo+uPhgnHxh8AZBcSUDXqu9Ybw2sCiSRQ044IjwsJp6q
K70TqXrDRreUlxQrDmaNW3KKdwsV4MR6ZupBAKtJR5JFV+AC4CPMmdS/u0qLwxT4ylAABWbXEZrT
pEQuCjC7gb8fzX/f8KQHowMzNLckyZo6RMnRnLZ9nna25UjZK4MQmfSm85Z6A0d16rP/fL8rfAKm
8IWWeif5BO1SaffDJP3268ABPYVfI6WR5d6Qm+BtDJc34hokKnsbUP9YjeVvL3ETuzhBBdu23PEP
bFwsK8DWQCsieZREJnQjFgLRFhDK3/DogMMpQNPumuJhvry4Ov2ispsD2fwVXKDQuZY4L+xjoKUQ
tVd8pn0L1+yVIEJiGfIfAPKHm9xSwsJC+WtkPjAPyK3BxOkdztWpwyr2Egrt++iZa1R551B6yXNU
5NwtZhzqma+V04oBGsNZGitS0HJWD7qd3P63EUMFGW1H+MbiYM78ylq0bP71AK44mxz2Tq2AbACt
P40I38F+jFp1DAU9uVtnOJGzhssmLOaRxjFiFVS7E/LrMLRTYUFshnpRyRgrdk4eoRH5cVYlJKj0
DKCh6zYCOx7MyT1jvkAlEFiQ6JtU
`protect end_protected
