-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Jt77rXZps7F3UxG5Chqtv5PLXs0AC76eMOCE6/R9RxlRsO8GRDU6I0cxA3Z01U7PPyVTL8TEYPQa
ecLuaArLAnjl+26ZXHZooUJGYxk2EK7uaBT/wDbFvFwveJ4+Tw8RDiX+HplhPybfOH45VGdAJBqy
TX1YK7V0yYlaiXVXwHTRtu8glQrOyhg7hy9FYzniR4jUbt5vR0PoNWi7Ka0A03uhnmZZTRNIwSJY
ioFoPEXeQ9BCPa4UjnxW4ZsgSkRFoOaaoNIEP0zL2p7oLjePFQJDUaVmOdgxbK+6pD/MwbKguA4p
tj1oobzbe/24M2X6DaZusJXOAGS8ie/syqvkfQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
TVNrdHEvut9Ekf9RTqmvuKcQ2SmRswiLAgPr7h/+8s25XGWdHYjob7MOK6vAKkRSCQgticQyIO1H
YBRPHOhp6XkglUCCHXcGaSp75dNBEbM7RSrlU7e7ckHhdn6EKCU6n1b/Yi4et6E8JkJ7cBCvBWbY
guIlQyFR5Rin5KLI222seMAHjwbD9+NtwpOHdm6N8ZF1hMH7YwljDUv36S2aFSvSEYLbEPcTOn07
ZVeDnMU7KYgLH6IKpr0NmnkBHrFMROUW0d6S815htbA+bdyejms2eFHyodN2wxh9OV7P3C/KIh6F
v9dvCpdBfu3azSHgOLcJnHX4Rq3z01VAmxOpzkc6f4mOJCC419yT4nBoO/D8X7Szr6NFGx68t/ts
OqYKGqH3hU15gqr5FESkvy5/RJPdoKpW4COG89wZWISdcp3TXwyyJZ+VZiQIbGnM0e719tgGTQBE
34ycOsALdYTUqBkwbmL3Bf9RvYalbRd5T6c/DxyvHzVyMiIOLojV8uDvIMG6kJqPxvB08K/4j1Ez
fEKiuo/ZTgUSq9NgTY+HC2V1g2N5efVwI2RN0J7tcnuO5AINopZXnMBd1qmLd91tbnJ+2+1gRo8N
QDl/FoHR18p7CtmTzrLABj7sfDaLCmSOvYtcxiJlevNBwnFpztIIpWcq3wDyadxgdso+2ShK5OF+
qqOc6ba+6q6QZM81Vnl9wi7NibDwvSfutGCXoTDqb1T+6Rxqq0Qi0USbh1MJJOzwvWOfzf4yG5H5
MfphcvzIEBVm4uOKVfXLk/iFC/aaNvNUw61K3zeS4O0oeM+sZG0Kko8BKsNi2XwUlQqkqIxk0mDD
CxUQhMYNynhQ15Akg4ADKpwu55SvAcPkJCzc3XJdQTPTSKEMqZP25rLDHMg+RX8DptTAl32LB7QN
zoIg4D7a8LvorNxvGsB7x35V9/c9lUXyJitcE7v4BdagFUPIntarE41lYMcs91AIza+0KCI2HNAh
6I1QWf1xhbd0zP3/LaaY96GOBe75zTtwzxz49akxNXjM63JWL2X8OI4mbL5u6xQpcMV9qbB6JmtI
HZ0uzhP6u4A0e0692woenCc3s1hruMbGChVhnyju3P3UIWh69P9DYhKJO4gkpLL2xcm96fpwcaT/
bu+3JpC8iWUbYxv5LGBhP2xT3WusKKgSYokjQ/9mdhD+NlkJj7GWiVxGduj6DZS9DbYQHUCM73Co
fEkC41jneK22wrfu0NIRh8cvA+nWmB9eScqFse859zPP6cfO0EK3CyRlAXvcHqAuWp/wH2kE/mLh
EVS4IGZFMDqs4cMiYtbMaELUpTuEyttuF5VpPs8oKTNFSV6cBxJZu4PLEZUeKeYs75DoR1PbGYpq
rpXtxHnFgchi7s3tKbZ0ibvFz5wbOiViF3/h5FqWm8dRaksm8LXKQ1LwTI9fPAmusGQ/fFqwe+LY
QlZGrvuIv5hZ+trC3dfDSMawaQ+pa+GcKwvt2f8M4nsfivs+LaMz8C6DJrCe1X1Oyyp6rciFlL6I
2bt/91hWra3fWTtCnMw5GuG/MVmjh4SuKblgl//5feME88qWKsvekwu1W6e/rrPJ2FdSY/XvHYZd
tkxoSAC2JgNR48Y0rWULP1uKwtClIXirqXYxkLqw2LfHtHhz55MJ3fJ1/7b+SYGpmUTa7fZ5+jzV
Y1pICSWu0s1JM4jWwfJIN3Y/Z3H6o6avedirr+2TKvK5bP1ivgeWySbO2tCrkOa1T4/O48yYVLpo
Cp1jA9Xma6eIBalvxnLI94WLsRy84wp7dZByOjyLOKG8CGkI3K04w9/Y/3/OfBkhMNiMSZyHyPNu
UMoaG63Ux2KJf85T2MI7JaB5oCCufVey1gcd+wV26dJGgZUdg9Uy129E0LsjvGWOnYKZZsBoM+nx
6OZfc2a+2J1/Hia/yAFuuqjaRu469hDMhy20mOVpgXBYXIRD2J/x2lxiR1MofWkiusxIq4V+Lq74
qBodYh66DmSQzDmPbWhqQ4Zh8S72Jjauwt7P6JqhfcW88sQYq6zcU7Ewr+TKmFGuhH18Tk5KfyG6
UcjaG/mIKFcxG8WnIKSiClnQi5Nv5MotwyQr/rIfg/NEYLeitGM0pB8YF6rJrm71dz35DGbeYl5P
ohhyj+IC3wwA2QiERUwprzEZuErHqjfSXkLcqo1Fgwh5jg7WjYmhgA83lkEbz4G6MXMxTMjVSzgp
Q5ETH97X6q286GnMeH0PsN9HB3aG92754+KV45y6ukhxdgBxBMXZMh+zy7aw8c5HuYx9XgSa2V/6
Wo2KGMFvz3DD/19Mv6aakc/4F8cR2AO+OotDLouHhd1O8oECOK+dUbpkWq6qHZ4+9yltjxADS7Me
0DjHqtdSsjcDhJkDlKCr/MNu5EW1VprswHHnWgo7hmMEIwkb/bAg/w7IBimwOWShBA4OkpqHVJjv
ugnHQDHsSqpmYn1Rz/VQjd4uaEZeB8FqW/ZbDKrCti8qaAYbdP2cxdXB1gATZ4T9rYdarPOChT75
c0ZHhiNnx2jkv+03/VM5qE8r8Gsir1qTHuw+R7bK4cOlvQZh44WuaKCYhqHbbRrpf/uUIaqjKT1i
blx7WdEilE0XEtWtkDi/s0nbn9uxX/yrUfIL7uivI6NSI7c/F5OmrJJkC9os3/e5AD4jCWut/26V
WtFVmSWUEAGsygI1uqq+ByEyhzI4iAGarmlV6EV5mmo1m9bw7f4+It8AQ8Kgfuqm+18PKmIAwMYv
cLx82zTO7F9eou90sx+liieQqJVVSj8gNVZFyI63b8HH+wwlxGQjYX2lREtvJ4sfDrHos0tIHR2K
o8EVANTWJtuRZRIWm/oeXpz80bS/RZls+1gqzUIQ1AAfsDkB5QB3UnAb9p0/DTJOveyMZtV6CTsd
r3jnJm3xFJ+1dtrah/m9LB/XnCwZzLmThBgTR8gT4aRB88RDQrZC9ahBjayW2ZOh5cMzOG1WpL7X
ye178H59yo0ZqO2O/DHUl3ogccLx/DfFWSSIesCLAwO42gtdz2HcXso3qYuiCaJwgLY0F330qBqP
ROw8gj33t+t1VP0uYKKoQCcMuHlzWRXNuomun3qdzgzQaCqHD0R5H8CZPe/qOCImC7VTg96fCXVb
E/qDvke7LaGqzT8Zftq06ompgtrjD8afnplnyzKRbk/5/92uwWHOHoVw75wtALqhnGz3o/dlsV/S
T3mp2e9SpgKZKlWQjQyjV7hJTI+1xQSymX6vL8aqW0kQWwQytztlFWxValgGrFHyNuGkToeXJZc5
Rtdh1ISNayPoC2nFaiGek01JNnJZ1xSkvD+SrW33zhbUMsJolojsRYMDNbPsRglnbyT8DjMCVQaD
EOXNHTwTciWE75T9PORBaKZAj4y7FXSKbiRJgSc3L1nB0fWQNF/7FjTkAXj3dJJwH5StBx5MLC5m
2pKz5IWaZ1j/ZXKbxhnUsVAKfTTuf82d6aJ98U4Xr7zbgcLYC5vYWHUFrNfq8Wi/QHQsQiNb3Kng
j04d9kUsrUP+wJV7Ugw2VKQcrEQ24Z5bO1xzs998Sh7EAXndN0dcV5zKTSyedAs0x2Hs7pNI/S19
qVebNPsvMjXgJ1UJf+EtvLawtueqMAXQ4ZkbQh65nQgJ0tctdPPWFCEG9CI7AjyiQ8hGyt4/qfb1
gmTHMF667eh1cHTrmKeTMRlWqaQvrYsDY0YQjnkyj+zBvWy357BjcwDrlXE0X5KeuI89ciF6f6uL
4+05P5TQpApZiww9z3Lah+jyFHNRtuoP7iAYNAZf7sTPM8kvoAU2D2gc0wogRZMz7mvjFVZD9yQ7
exG5nyWwfp5cDsxMosl58tQ0AGeMgdq653Ah2pmQbz6m1RI2WDQE8dKV49fBu+frC5cT4p1IaTtA
9l6ypKPUaKJ69SoTnOXlyhkOx6juiR9aq65f0vAXRnbtJLkxEiDI7WjxUWolHBm13H0Gc2PhIO8M
kQG/3yV4SGczXrQgOSSKgjqyPf7HWdOKmKBFqHR4C/0WEHarVeqC6fCBpK7+WPva2gS1ttGni4o/
TLfCA1kcZZLCNQzSR0TiTL1RCibpquI5zj39qvI7uAt0tkXdZxJDYjBAfyaLKDseyzjij1xvxQWD
Pxcg2OzvSpJM1FwRHrhW2iEI9BFoRTODTg1x9oqZqhDbwrXmsGj/T69VT5h0t3DIDwa+Ec2hs9t8
eL1C2gAyC4MZzeDs92JbK8PuVwXuNOTiahsL6uqEhm9sku1PHbx2XYs8V+WpEWV637AZnRNrsD/x
hfXKo8PnQvRstn1U7mmyMscyiiy3dNY1fF0qpP1qx/KN5sc7+fG7vDb5/i5eHLsquFn8lAyB3Km+
r6oacmeBxTbxDgBKgCvuwR3J0B2+v4g7YDyK6UTDmUh/AvABBqcHymqpN161ix3rEOkmiOvaE815
aPM2/AGQZqsj/hlTRGCnz7qgpEATxVwLEKEKl4xTQMoAAyiYnMGqRCabPrWgEuErDJiX6pkx1Ojm
ROUD2cdfJtzNciZKkZMXSnHsstMPpVq5lomPWCxnQic2IZy5hBxCkSE2hFb/eIBWOO8OlsDRagfh
eFh0cSy6wbxJxZ89uYlc1ZyKlZRgjTLPa6Llmu02ICg4tVPVcCM/HEPJwSMmmw4trbQ59jf9Lo9g
NyDKst8Bb5dzxju73fpxZBBQrAclGu+nwrV9P72zSL/Wmekvj0jNpQd2eRK0+fdr4JyafYO+xn2V
X/krekQLPrVvN527MyQ2Sef92mgZ3g4XQCAkBVkFQtIzJQvHjwHyimr7aOnZjcckuJksJzVeqGFo
8O4Vmgk2h6sVuB4B3BvtPHFcJBrD93xlzNz5/FILz+D6ZHsUmxC7NL63VfSpopckY/SkgMIkTIeg
7tWj1pZtS/xfSHNT8F3Gsd8d/KMu4oIvmhpwpCFABGm6px/TGHtoazzVNbdWjBUEYDwYbAkfV11V
CY9OQ+hqf1oNcyt1XXVyVGuN9epU5j5KSbOE/4e1pu21mEZUZrHxrcl5ocBku17EBjoBRpBmTR7X
O1GWJiKfnlx26Jp4E4THSnqyz/V9bxw8QueJcfHF6rXW9ihrNTERsHrMXHApj/G6Xig70NpQgDOW
iBRpas5JmFvPPkye0jU9FZmGwIrhcZUeV+XyWn7BPWgfNpHwc93Thm0/NLatzAEQwLuJEnwzf8Iw
QoVnoJDLsg48EizbHuxVcAkn1T+HwdUF4CG8mxWilfJcGHDTOKWViDmBcBE/65d4Homixypo4hQL
0TVZ3O3Un9sA6fTK+OZsjt1BHKMbWTN5RFltEUyE9wdtVnykZwwIjr8RFU2g/KFA1ve5sEUDEKoN
qvEHvWv/IKQmQpPV1Xh945kD/yEb7tOOvj2g2K11ULkYvcp24uBLWuS/XP27z18kOrNYwE8eosUY
BF5EgfNy8v+JzI1qu0oOav07Q+k4WExuIVuBJISAAzspbpZWOgfciQxb0H1lGtGEUyCC7Ip6F0t5
JQ0qv+BuqlsSeI5N2OOGXhbIg5zIuLzg5SKTduegaBCFKB9ZR3DqHcSa562pDwkzQKN0CwlvA5ms
qtpdnPL7zwNl9u+7N2OUMflZ1i3hvF+uoqQaRcVMpOsy+0aInDoNIiR5em4ZKkZey2bPpd/OElFs
JBg2RfJq0A9Ucu5rT8CrFevZZh1mnG5eC9SQiQDVNpI45roTnZxNAVOMqYt25czGoLdrHRJfU+8d
/LNGbNPKaU1/sRlWUK+0lJgTEvz8AdcsaIip1kZ5KSotEFHmsiiq1CH+qIdExgbmW43EDdx6+vEl
+eApVQqrnRKGeh+nxnjo3VFsNMqIbJOyLazhyGkoo3fN64JMgIvpJxv6qRvEAZMwRML3o+fPMUUE
+BU1KCmyhjBKTKMeD5BQ4NzV9/46APxkZ5/iA5bcy32nNfuqROesBoOMDepnA13TJBj4d0DoDwQc
7nY7yRC6NLX9wcuDwN4f8vOETv4ZU0NkRSvbfcLtjLapAXfNJkJ88vcLnr3uDbFfra8CHNa5zlH8
wDlPOzC/+E9oVI2ozewkhtvw4VM/i4nyszxW6MNwEp8aQJLRYSW80D4FAMg6ZsJ5TgFmDOT28Rvx
fTBOmX+RirQYjPuGOvzv3wcijzbDMWseI/elsP1QOjyvJwQ7I9qYQPTdiI6hr2hwGLPR02+WF1qX
HRrdN3Degc+Z0jhVQpQd/WYk8rUwO/u75CGzYh1F2+3rhxuvU2mirR7OCtOXwYPS4aM/Uw/UPpcY
Cb5/8ItDETF48c7IW1XvucWsOg+Qx45M9ge5L9n4nfgzF+WcD398sfxSA3z7JiC+PeJWzHWdxmUP
dQxPM0taTuBwSmMGYG3YzuXRiIgNT4BIWo6/uyYauBVaE85KYXoUF2Aadu4LdNqOGe4eCK4STxAl
/UKCtwJIrvJDHniMfKmz8GYvb8hn8XVaQGDjzGKcjU1cU7LWBVJZsOlcWFzYbMNIYCGnSRhe4fSG
KE/dMXuXwaeBAG426Cq14dEASnvr+GnCTqPxoRT2IKXJ8v7Sc2WLzkYZb/QXs4DJiual2+EhSWaS
TGweJOM2+1HJcS/nyAABYyMuT4mNYgH+9ob0sNtw5cFkEQMnt1MMWfjoNVShdto7M0KVCP9a5VUQ
91HyrjhB1kL9B/IVoaMcty+pD0A/eGc4SSOKWbvkV3tcclbg9a8g1hFcG+9xQhq/tqQeb44YfQe3
ik/j3PIj0Xt69KnOQcLkvnP31gwToAb4hu8RulAKjRrRWpEXmD7aCUL8KmmEp87fKww0pePxJSUu
on3Rrdkzf1wHKPistPzEqu90d5nmfiuFKs4z4JBvX7FNsPunJpAcWp2Leq47MEHeSzk0wJ5Rn5m0
d9kj1pyzNIqpq7kdQHJWK2n13n0X/ArMvCitu2jNF1EP64UoRk6bl4kmshczPIiW+L5Zl9dW/ZJC
zxIJ6m+Vh2WXTOZMw+pUWB0hy+W3dVd4m7jW5is6sfK4Fpawcs9ckHHufj3YjoO7elK9Omemy9ha
NpbWz97e37GNGD1dcZExPMsMHN1r36aNOJfxKuMbuVYeyF9gkH4u7hGYkgFOUczVwFk2JGYiPTWc
ZLhxpFYJbfHIiPWN25hzTabhO7RL0p5amdbeX/EjMd+RmvG+H2wuNfsOIqfP7hSz08Ai92phlzJl
RUYZ5vPhe+hLOCnPyhp49JSnAdrdHUf1u3JcAuPBlniX+TrSUONjlct2O92UXP6Nud3DcUTmsgWd
I+yFYN49VrE0LDKpe6gpG/TB7j4bytR2bHW043pOwHFgWrgXCDUNMA8O+88/Yk+gIamn8d7BPHbc
xxHs7M8RAAqmn8j6TJtglipcuM7CbChDnj1bdjyCOVUalJpAuihf9yRKy2eQbYRTK7t6sWiwyXgT
sALNht0nyAhrQYneY1JOmffcyur6BcLoKQWtcT+1FHy0EFyxHIGAfccghJZdP6gkY8NOw7XhEfk+
VHsLgexZmLyTRqycWmDJDmj/Tg+dXlw4B4NBNZgpgBrQHDvtlaUV9ewZ3ppFOfIuDfjqglm+o6DB
DLiWdB7O6OHJICD/xd0eU+C/e65rSzs9ylY7hW9jeuQ1zP3LO2xRiV95LWMjTzg9jBRdfmzOtPae
4nwX4XgrVAxeRSPpTM9oD66qbgVYjz5XMBskpWceBQ/XjO8klaZqIy6RcrASeYGtpk79puGuwFnW
HtzshWHhzVg0aCPOZ4u/yfvjAlNdiZ7fUY276w3BSbt//Pyr+KOKivGbYImQRm++rDjKBQJw1Bhd
QgL4CsmASgRUC5pZccBV8YO9xRN7Os5LjWmtEhYl/YhwTHJkp3XO6n3NWFE9Bom7+dARvbZx54z3
M3OKxphURYuOkx93x+ySpQH6i73AXAinTcpZDbOk1QsbXxx+HAnkyR2FHRymissZ+gMQGEnSCB3s
RvhG3SAQBNxRhjqDaw4wtjAn2nh1pk8gyRSnwJTN0MPi7OUeg+Kvm3rJgjdfvpzxZR7aVcGNp7IH
netG4ko0/TFVdaHC+1WpPvQGZa/dB0B1AWcl0k4aPjumCkvrw7yu5tN2Gt9f3ZjNJPqZkwo9ju3S
+13eYgeHdSv+KF2xoAqDyscCHc/T34H5Q9rzpMj4Tyq9sVHNxzH1YtU14685oq2p9FsAU8+9T3zQ
8ZtYVmGrFpfSQttax4amIxcVLx4qcHDJADe6djmQJ22J/Kc7rxS1dZykAIntZPKd2/QQ4dIHiNwp
toOKcwC3NwxL+8aRxweaapJsalGh2O/pdKc/s+Wa7BmdsK9/eRQjrL3AwEauNFzmXiPvHAJZsSch
7g9u76uPVa0BjzQsbg6lQzBmGcP/i+6KRq0w9zPWagKFqibmCA0mUfeyClyfX0x0R5g37y5+coVp
EiAR6TQyUTml+Ptop1VXbBhb6HxR0ISVkuEzo4HRb2cN8JZf7WI4ubMgufo8LL4QgWx6UwZ4J/8J
kCZwj9Z0BO3nWTDIg52ZXOFPgcH4w6QyyAbzbDM26AubRCPrhnj0qP6kXs90o1+mUUHBtfTXN0LE
bl+mWJ00uIs3dBHb4EAztaFe5cSPWZ/Q4QqtbWU6vmXV4taC8EYv8enaCXDoYGy1y335JQjqtW7/
j4Y9QlUhWfqcf8kChXMv/2sp9nZ756SDWsWpLWZ6lSmoaWgk/wG9lUk3vtcHd12R+heH1jNZK0Jt
ufyoM2J8LbbAYuBrIEBMEnAsJ84Sp4Jw2B7TR+n6L3JU2TRwKl5+kGklVmEePefe4RvjV+t/DDay
c246mbh9D5I9wuLn4WtLds0gNsga9SLL5VqEnK+/KRvtKo2b/nVWmr6AsEsea2SdX8kGKK6tuGYw
g82VTGviHlnul7++A1otrEfvwJ7WE1JMYFUFU9rwydv+euC4kw9tSzetaGYmINvQgX2RIa4juwd9
sh6Gh/zm9HwPnBVvs5mWQL720cLcsHSCYh6I6EWkVLZXK+ZuPQu7MgyS0pbS70n3g8GbWBkiTVec
QLfl5AmT+T865G5qkz4PZQbTDtaEzBe0FJiyogiYAl3SZQRNbLl/cEd3nMaFBFAG4GnKFupaHxcV
CcqkHvX/N2x1aIdgrtB8qhWxvvHDrAMLYsL78+fCLxt5GaEDmXPJgqf9VuJ7wtE9Zw3dn0/H5BEz
YadNd9y6gt1QBHSdiWTgWs6J0ezJ29DRUQZdNzzPa6Wt9RbXYke0Degan6R10b2g8JmbvfPgGJ7I
wJJconkgJhzQyB52zcgX7sGf9u3kkgO/OnlYy+Bjtt21MHsu1aqR2zsOVxrz2JrICvl6EpwEm9/r
zRDsIcZiw7cupM/9EuszT2Yn6450oFn4dW9tgPnBF+XcN1ZLBhhI8X5JpKdBBbzOIYiysdQOyw08
nAdGA9D/osanldH32xkF60918RjomfUj1VTFQP53kTUSbmFyECfozNfILliP5LQqmNh+ymeSAk0y
OlInv47TaBkOcPPL05wJpFV5eussJLCQ6yN8+zRHxJzdClve0a4a3Qqu7Af38JFFSYgFFvQGmX/c
IOUu1r7PE8UGFb3bbmPPHEKlTPRiTUejzdZ74FfCl7pF0MojohU4Q3dp1pYYQYqEYa/x2LqgJV4B
pP3WpjxxRUQMPgz7U3WSnG1+ZLAnCyhp4sq7p7kRaenC6k8oaQzsWiRht8DfmK4qqsXD1kdq47oq
RWbrZ95gLcsC8fA7LzGF/cCrilHxhZOlEUgeu98X8YMEXICLdrDoWcCyKrMck4L3eRssZXKNpz/r
He5KB7AJXgxgPqq6qbK459m/aE6ax0TCJK9astEy6/5N0jQLbIbPDMgP/YYQ7pHYjU6fz7W/nKRW
WqhbvnHKyHIAZza2SWhk12TN0uLn3AQYxXHZ2u0Uy9XdSIlF072Om4YKnlygWePemX46znTxnxIZ
w/5tzNYBXOTwNNfuAHRyVsWay9Wq/iiSeDc5KO561vydYyLO+elMFsf3OmRrN0lTGuiNTqXdUScR
7UnCVKe3Oz+sc3XfkhXg/qkE3OliQ1gO56YWD7eZRH7lhJhIGqetqAIHO51I6K6VpUMYBLoDTAE9
SyjNyUBcfnthMPZWXVDfx0/2nsnIxaEpxTXWMSO7ByBw6bqSWED6mbHhZFaU0CGm834koWit98/z
Q9wfl7fMW0cNvF2yE163shPkGm42gyt//Cx8crlUjEni/g/ybX+gJyrDcJofFfHpcMUnw7da8er2
Wae4WAd5p9pnWPP7oZRUEIQzMs/eXCyv0EAMEvw56YCeZ25SoeenHnkjGYMVH8kf0e/A3afmIeg3
r7gQYIQdI9l1960kBy3dJhDSyw/E3xIOYpRLgqrZ8HnICAjYBhzK034CboOA/lAv8LiWZRIlj5rp
CQR1D616zSvQFVhzMcmqZqt9PZcSmEUJJW/aRMXbRTxFu9LeMsQOmGHZo6wJH4DgbsonDPvAOXys
s5mrAjQF71v1PkiGts8R6GIJ96X9SP/2PeVZutNrBmBcL6YYAuehUMeoMxkNg9EFaHL5IF+z+i8k
KyF3jB7SKn8xNADznfk1tXGpKpgfDqLoa9MAL3b4JbTLHEgnx4mLiAUhBe6nZ51ksWjIidIgVCh6
NkvJrw8pt8FSfg9bRrJQdcQJPndfqvSxlHRYQ9D91tX7pot2888BUGPFsL8QtVXLG4BCQfgJH3MO
En6IkZLCgC0D4xy2k7MXfJd20WE9qe7ZrN8cjqNL5P+K2eK+1vSwGxKY6z5mbNo/C2H+C/1NbsB+
9FyBpAod+voAD4A67v1ZqrPVnPsQeUXWIzelzufQZjcyhg74xe9HLVC4TJJydXmG9mkdpU09DrEw
kNXbo8pgC+grYKC+6FoLCcrqWanbCyN/h0qqQB/ri0n6QbTs/Hvu2ydQQsyhGUdWL25J+0GYGJLt
5g47ySTfyVelrqJR8r4FF8byKHJABQSrjjLQnqKhUXSstM4b2VW5vdOfrCupFkEjP1a1q4o3FkfX
ESZrHG7LTb7OdN3/nMQnIlUniLkXJPq4DKo/Nq0LgWaJXPdLP4us0BLYQVPRtVRStDF8yB+SaRza
zCjnnFPba3GaP5yfs3bhLevkwCGAX2mw5jGWXZsQV7rME/Mvh/s3z9xcOLjabBPmfhmNImTBKTbP
f2qLAfrGpnoM7fYocCUvsbFnaXqEO+EIlIDVNqPLNqOWpi3HgY7rdyP5w4LO8Bs4KxUP8dlEfdTg
u2nxE/Om59PsP8wrllc/txLV4TgbUacjGwvtg3BN6ofr5PQDW9dS7G+wiAmNGyX7zH5kNyaNkzS8
Gn0vi1NaEFiNpt3nU4Smh+scS6jiToF3+VNxuYjQ18mxgrhJY6N16gbeSfR7hrIG0cjsy//8yw4g
KBq6oquFU/ipddlExOXYRD35eB06bu+G+yLFq3HAqva7CnMWVQY5Y9De4hpNElHuOHVeH69FBlEm
mkqrjBiLt5KcMvtabMLgAb6oOAOIqrrNjJ/TTXDD1KCAcmOLjxlWMrWk7/PeXbFck0YEnx5BlrpF
XcFQQDtjlSvAHnPCQ8VTYYl2UDmYyQZmLoAbbHUIAAo/tkE7uux79pOqyRob5mlHkmEKWsS7M2mm
w20N0ojK4aZth2GWZHaBhBwFBFaNGbQ2FbpTALngmsowwFGYCiGdkXlGc0Uxm4i2nIbycSQcvCPW
Ty/XekscmyrUBgwkFRAxYlCig7DQlwrFK3Ay8TlJy4LDEP3IBf+IET5dqBceW26oCwX2c6HJLFfR
fvM5gZNrYFUWgUzbabEhzhO2VBqhojd2ZgFYaOre0/thNG2cTJU1kSM83SevhqZA5t6T6IFaX0qR
daENtDcpyoHpF71kH/7vcwQw5EZUv84RSaZUR10ixuSv9yVX6QiOOHSDjW1+JAjI31qbMmiBFqbf
RosqdK/EN2hji/jAE+7D7wpzaHFKvxoBayTMSPYzQdCG1lRFDbUp/7lTArIcBOK10iVFEqDpayHw
Qh2IxbwqLgih3ivhBLDHiOiY1F9I+9r2gwbTYd7TyTo0L3sMNq0iq20rq97E8rJuYIfM21Gz9NLw
AFhdsRe4QgZn3vPGSHrEORH9twgHnKeeGc3xEGqH/m4P7TxwZE8LY9m7HuOD4VSfFSFbB4gpRC/z
m0/7yPa9i9SE9WK4KkHPPZDPbRg8pQpYrR0WRe3pQwJtyRrarWBb5zaCub2E2lZTswkBPd9oqvB+
s2sfgV1pwd43a8LbEVEic22zkffiP1Is+GAKK7I5y1TnwCKGN937bd9QhcbVF+2kJgi2CQGpn8xq
dSQqxTDwFzQA/dTRQ0zh1bjBcG5cUj+l5MgqldiwiTiJGZ86L7OdA8a0fnngH2nW+NR4pzRBN4SW
MCWQBZRhP1IFKhjX4TysKgIX9TNM3WpAHHQE8DjkaxhafT08lGoPS7IushxH+dTIOPRV3cVnp0HC
y92XaMz7HaMCOmJXdGcg6uAzDoypTp4/7ejtahJ7OoKiUCjSK8ZrQLTN7hUR/I8BQB8Mu5o8pOKz
cqh8jwg6evcemCKBatT6brTuqdFbgU72n58AmgJZqBZkcPNANeRQMaomtJaslSer791nN9SaUO+u
aABquMXlu7FAkIYLuUOBKINrraCqTyNFVUz0/HfW6ZoKzVAdUPvqvqqe3M8WyVI3TuXZnkwc5pyu
avEQE1exbssimI4Ad1N8cJe08yuaPmU3bqeqg5lMjHpoS5PVIqjByObmSxC7dhWqvPTfOrQgvCP7
HRDPourCWGPSALP4HaC7xLFWvxlmQArMi+GDkEo+Fw7BaO2vg6CkD5XIpeHu7ZxRlaCs4MIosFaf
Q6Mw5v6U40ZrppdwtirJrVn8Lto1NthhWAPOV95iqCTeas78du4jk/cz2RbNxaDIxRPCBvfwrfsm
FUJ+YrMcILxOHZSnQZQ+wF4+mw9wLjiz70rmYXfTHBMn4iY0OyCFQRaOhBhGwXveVO/Xlsa/VdKa
5FPbyUBewYwQZ4rTlJeSpopXzEhLkFPCEAr/NERHT7SX2a+86GPRDATXQYRJhoNrxtLtHt5JMyPc
TeB5h7O/ndZ4jN3QQZni7tHLTFrL/4c4CHBYhKro9hfEUcZgR0hZhGbSR5kVr4twjgCZjK7oNsO9
EEe3GyZPGOd88CYzeZC9C2R/OVjx6DZysjBYMpwjYGvQwaZ/rmAy/nhhgswNZL597hLGgy4Ql91R
MlhWcm3OJeDI5T0oHdeDTwRisrmtXE/Bc7n262ywch0n4/eDVednvohienVpVLE3j8C9cZuLE/y3
AJqqcPrxRXu2LDcktdqdLKIo0MfhMZ+mCM0R+p9X+qCiXF3eCrVpJsdlW3224jriC2NjScB5BMRg
ESzM3dV9bAk0rQpjDMzLjzu7BOhnHjHRuDd1ljMhNbQhBtjYFSlOPaWrw5nmghoOp+jwXQSSmm5D
dQlVFnOOdsl07C4bJ6P0OC3DU+SWYGXvhUNUqzQ8o0GF5ia52wrRX1/HKsMbz6U19w2MTYGptRTM
Q9rIidwibIbVnvmBbNpLWQZXAa9PNvji/1JWSwFFnxDhr/YyV73NbpJZS1KH0EHe3FNUPVlBQPtI
dNohiC5xq8ki+RZnWlu83gAxtPUCxBrTL5dJBYomQROEsO7lZKGGG//0AZR8LNaWy8m3NOBRtK0I
IibSviiBN84rtN7dm+mUPtk1kmU46jihZmQxWuxKPNPHS1pqpS0c9QkOssVvD37uUh5EMMCD9l0M
/xOpk7F73c0wumGucmafHDdCIY2XpOrJ5a1X3Hu8w1/th2d2oi4m1ggTXHoCCbvqSmuBU50q3Jb+
025ksik8jOsyVa2PChAvCHHMisGVrBQiqGz47NxQ0xAvSDlnHaXTn4PDJPp0QyWfGpXDMaSW+MYo
urpWRgaXOba1tZFgV6WJrLG9ghHXG9e5sIpshDXRneM+TRnUliYhvf4ubwJYg9SmeOxP8+nQ1McP
GYqg+pz2dHIkrT/881Ek3SXWo1J0uwPJY0DBXwW8p8q9YuDgF65edIOTgWM4HYltJpZibKAMMZSn
P2tv/r8CHcKWykkV/Yl63BDklaye47npZkQZBdr9LSEtDLaaL2WXMDO895stFbIsurWoZ3VHY3jL
6iHWBPRT2dItLrcrWHLnG0y/caMMFlJJbwPDHJQOSw9t4z6rJV+BEfuzLCQCYsQbiWtKRvM6ZYLq
EWD6fKWYayNxkDNup8yKsO4y4oXjeSHvk6236LKSeCXpZnDHWUZST9AfEkplYlKPuemCJEnfP3z8
bXevhg47pwuFoBnCUAOtyQ7CiFHJzWArw5h+rwcIIcgyl/w08wZk1WKghyCtYVDW1p0cLEUZ7NLG
kLWjj4gyw2fwM2lIYEFGxu4A7jvbP91E2ECF17iC9m+HHT6z7vIGQ5Ru3Dhdxh957HZi7G3pveR4
fCXjGfvGZoBon/ggzefiCcNeQh8lOKDtpi6Y+t5RBezAh0ADOsb/oXpMZCmLCgn3lZv7z8E7B5qI
UvrwDQUbo/inRjmodigpWHBRRBGuyTsWbgfwsyShgBeKC1jeX28Gva24Qpt8stpjmuhuu0g0+EE8
URB4NVS//0uKtW66yo21aDhq8jNv/htevRVldN0AzjQ6VXBSoOtmIDKrND27lqHwAYJiFjbyiP+i
oUQi7tmON9UuF0M2IjzjShx0J3M4lRRgeLOtGiuR5+68bqWPzsuR+FpwHpZrtFLRcXQZWiT+ZeOR
C4KHwncDMfcF7iEhDL/mkE7v0gm2KwY2CH8CanJH3xr9Zq6kFiIJfI4WbusiFu5mhr1UoCTGYxz2
RkwBi5KQpM1pD0N6lSuBFSo63FjSNKs3kAOBuPAv1M+YKKs2A3V2PZOgmhBzz9AEL6hnHjvSrEUP
NdcdzCi83QD7hI2vlZ0Jg6xySfuX8NsJ0xcGUYKsJ5n88QpsGSvGloT8Rq0Odq33c9msw/mDpMXW
BigqTAvRHVU1v/sfMlCwnYQxWYcEwxnJozZimJ75JDjZoh/rM8AR9jrIMG3l1KaPkoDd6bjGbpsw
+rg+pZ2vrfKKwbC81+4faTl8lSMuEK4jBtNunNJNRtuKxWMhdhMeWI5iMoIC6YA+OVph67xWDG9m
BA87Vg0R5MJgUN6hhRfA04yjiDDKu3lwT/O9se6pu3yqyjikj3jeUhi8ltSxlKJ9R7Au4j9wqtbs
Qgui650jg0NK2SmZTbkyZ1k90m432/gDn3ysn1npKyM8Ohgt1RKB4J0ndDuR2Boa+gAM09gCOkGr
tjO0Leci4Z1yiaNJFZikTorqypKZ2d3ImXfI+GjLg3YGvmFFWo0s3qLas756k5o1EC8clrGfcOBZ
muxviWHKF2ZpExgJk4E/2vreXlyYh1XYlOXG+fIm7tC3mR7WVtepSpGbUqumyRORHhMbgfRSvsOQ
aO77ZXkjtOWyPVo7QfChW/Ljdm8O+LYI2J7+HzL2ZVGrZe2gj1vamM6wh095zUJ7CSf1KGCWdbE8
DNbjeeyD32TyhEoIRarCv3l5ZtIlucm0aslvbX2Xg0X0DNqeiJNr4jn+aPRf+BPBRvV4m1bWjvWb
ayt8/A14PqAhTkbZ+PRXmPTz60QrVhLXKiJ2oZFjTnYFsuMojxKRgi2u+hkFjZW/kZnyc6vYravs
/PqqTMpAZE9aVUQlVBnDBXqhMyjFGnYmeeN++fyeb77uRRpFSsgyYje7atdfxkRZSpSCVfg3fQN3
Szs+MiFceUuTg5gnECccB4kxsDoGNPnBRLIoikM9n4K18GyjZfHz969+y1raWMq8e1zd4sxgu2+u
/GoIVYOTNQ3L/5zqOH9y0hGhSETrecCt4y5PCG0ZMDKx69CegBVp0MWBQX6UA+mmyiDnlY574xGp
AmcsfH8VHpqOr6x14Id/bWXsqbfPzhkacTac/NOmm2v/ar0grW4GLHb0ppFP502hHGkTzhvPw3aK
urPMRqFnm0n384bbq8GYK6LsQyMLQAeT2VHRwf+4mSV4c/MD9d+802LMMP0Z3eHfLFVDe8e3bQoD
ebqLPuciVSTTLVZJEzKh8JSalUkcNpm4TizDr5DZ3c0/foBe9FNGo0RANrazCrZLp8E80+ZLwPl4
ZDO/hoRoFBJ0PKONV2+aN5foPrQPWtbj+owXJjtFO/StJWgsyjcpSqU5HMnE055kxZxXYL694var
9JuEL9UNSfMq2R/eKO/3vF4aqZRhqMY6oobSmU9b5g5RErFncu+0RxMz+4oeAdg8hu4vqOsAlFCw
aHa7+B7kBN2Uq0PyaKBRnTlTsSjFULRnMnQ9bGwdTXhSliMAI0KNlhkzMPtzGysEvbqQ5bvz5PIK
Am6Qtuk/4hixcnNLOYfSL+RBoN50XSJq328mmYgzKdiHeVgugf1hBnFoR+hvLa2aONFH93yy7lgc
+finStPvW/a9xc1Hv00WtMvxKW3RwV89jYvjKIEM/r7yy9eexGw6146CZCYyN4XwEAoxM85TfPtP
a9Ly4JlVqIeYfSi6BZkcASnEWBrrEzLMUPGLuGUR55RKKP51dRpNATDDVyHIstFOUhNaKPwmZ7+H
e9XWpcHHe7WCZM4GU0WZ1TpxqINii1uOteHXCYb5/g/wsnDeY8xnvkRPjk1KU8m0ojypeiuvIy9q
xuvN+qf4/wdgrZqNZ/XeUORNPZZgnsXGyc9oiBUIdWLuulU/9cCKHJYDinqEPA60yKQm9sVxYV3T
IFcg6AHQdPtKPbBrWTGH9gG5Lo6kfvfoBDRZyXjCnKl14BRSps3xGDo3Adi8H/g2F+TpIicJV2Z6
zCrQeKznfkIc0b4VntaeenhjTz7zIaka2+WjHTIsbHlRwgwuKUMxX46JKJ699fulmSXoSMreLn4i
wc9KGWNwWwDva472QpiMGJVIWj0XAFLZ4sWnPVDTh/UTPF8Oow4ayg/jfbMMfelp/UwOknmwq3xU
nF+aVCRlCspceHQ3XCYVrmdbvGc2MFzQKgnh1JZnlCP8I81824eToulBS3ER1vqJaq2jjqa5dPf/
OsWOHeIJUyzitkOCluqRubE2M2ANZJnAGu/rJSo4EIqmWaUQytqF+6wQq0hIDNQ1ggfFcdRfgQkR
XjCz2tu5FeEohryi7wHegnjI001UjY/9A4B+pW+L31N95ZjICY1xvlO23nu7mVISxlCupekNGeMS
buiU03DPOp45rCiQ0LvjB1CCLPp6Nklk9jAgMyR+gt/s27lKVVWOQfAx8HkdfnNHlyHCLoKShJ92
G7PS9LwU3Fs39hC2qgEx8zzKPW9a58aRETNnkPeAmstMz46C2liyudfloQE+9lgi2bDPgO6E4+Hr
BU4ShYP5O8OLi0vV3wae7JWuj/BIS40TD60ySoKgl0aJnJHfwe9r7fbo1TaDjkHh4L8wLkbSH/qG
URkiiDhNcR8wpicDIzyBEm6k7vCFv1Zu3AkNi7JQL1I7AaoyChdGLfl5i0uzjXpQADXexCYSttHK
E7jAYPVcEIzgRZ3xBVYVXZufMLCjfqtHoKvHEifYCXR62sd8gP9aM+lnGN/XCiuS/kv6FBa5IBxQ
VEeJN7Bddrr42vJPDLGaYJu6yIcwcCIZfRffsVwV0xE6J3gRoY1pZm6TQi/wyun4y9zaAaCpf2PG
e/mF9ZKoado6aBdnlo2DATLYOD1D76YHKduO90XraE3ZRJEdqG7KzevtIhaJXnqeR0Fv5zWc++9c
9wKIqRjUYsvp8q63L3F8GCDf+pyEWSyAn6+fi1LfsWb6AaRQzCgpW17dlCznOmzZ6kMY5vt0y+yL
wrf8rOOYufrFCefzjiNCcf4AsIYgHr+jQXtR+ak8DlP6EV9x4Us7i81nvjd4r3nPu+C/GvDEpQRt
Sj3+7CIO8hLLBJTXcNuPEEaiW6xnETRHBEcj5CB683AxEBHkus3SJp6Pl6o1DNQol+EEDfyQaNGY
y6/9dD5lkWwNfssVdo+lRGVtAdMVNr9Z9IMAAEO1ooMUth7bDURF0TQRGH2emeaPJ95ruXGyt4K0
HROSrrotv3MYCAv0T1HB/xKMaJVL2hThE7lo7J3vMaYQ/1nyH9y6DBnWxBXLWE6e8S+P5hPhDJ/q
x/ZRzWiEwF0DZAkcCe7/G439hXOXhSB6y12nlcIn8TvX5rg6Bv8B9kbscuyRHdX53ZfVVbxizGC6
DpHsPNLHZ79lmoBrLeOlM0Pzh1c8nkeoQe1jK4uGddwJNcWA2zfFQNtqAeagmuVAJQ77eVcgxe7y
tmQTJ38T5JD15o61SYlkAAiiiZEOfqgomPao38dskE619zHs2N5yjGQsi2GXcgW+J51mWnFxaxC5
0TJekQr7CSFWP7hi2TDpsmf0BdF6S9VzCM7fmE6XJiqKrgiDxhQFjF4x6soNUKTGGnp9UgiuDGqq
hfzGmQdk7Xp3C09C/vsK8fLGpfaC8SdPNU9ZQ1Ps/RSevbNc4m0UQLWZb29dm9ldeD3IrTXrZg/j
vhMaEq3vOxGDWSiIlmfhIv22kacUwXRhM1mCyu4aadLaxM0dAzjG09GTJsp2VVDBu3a6y+/6+SFu
tLwynwxeByxrNRINGcS8s6NUQ29Oj5Szp3ltM7ds/1RvvulYPRE2hE0iH1SluBbRNR/nZXDx1S+q
cNY+x/udl6X3FsXqf4NNJJqli8hZmSRFh+vQ1novnU/3pkBfAPxhc34ZLN+TME43bOVVLwz3GBtu
s2PyfK4He9rsYuPoRD07XhOJ/GiG0pwxZm+WVET6Mdc1qwj0RwqzVBKrWgrmmKAABY+F11uCavqp
hLKMBkcJdo0hivdnDo1u8u134lrQUeDPrUI+nIRx5M3mO8LavxOTnvbFcTxNonYGJOo9SU2s0v4s
zjpv7kU6Ggh7RkLoiLI8Q4nqSUNhwNfJZxH1MXSSEBoQjTFoCSPgWhX/Tc1KFeXTnnSUtMxHfO8E
qXJ9maNdNQ2zIwIcHwDkfWLWEXzIuLXxMAIvlyJR6L5zY+u8RhpknUQxzsNHgFPUaHqcSQuet1a7
FUNV9m098nzu1D5I/tCic70U1WS/fGXRZpHLSmw5K2qJ2EnJBptcNJ6myJpQfIeEHaJvgIXcKvcK
YLSwOyVARUtamCIMih1zJ1rCcht3+nETLWWqsVoQ/4yNW0di7OJrlRJysSM84FQ+yPpEX/G+H0qM
aIX1N44QtjyZ9YuL017hkxNmgqiHje8QaqCCNPfGOGtYfdXfVb126xYNcUjbFCJCo6+jDyJsKxsq
RleUnwSDbC1obc5YujluNC5pS+SINJry/GB3GNqtekMoSo9wCvoywI2cNSwA53xcO7Ojbphxj18f
zoK3kqeZJdYyaQkRWTjT+L0H+dzIpIepce2NeFG+DOoc7LrV18D7ETkF/CvdVpUQlfl9NoEu1F9D
voP785yaVZAtcb/BJacvL6JeRlGwTEBLlX6po2CzYqgVbF2DYU7Oi5t8yk8GLR4baa3r3vE6cek1
UxsmDHgkA4VqaUWcYvoboOIzmHLF/jUgZFk281V2amjy7WwWSyC6w4M0TkSo6p381aCfF5xIlpgr
XHUdxOx/i8K/i2697zJnJU9fOpgN5J5zap7906QB6vlPMGxMdrqkXcYwcgHLT5d2ZxtEiLRD5qQn
+RbSV5S6mg==
`protect end_protected
