��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	R8��&`XAw���UZ��,u�]�b����3��jWÚ��=:�(�/� F����"�K�2H'6{~_�s謪P悤%J�1�h�\����|��? �ת�Gj	F�ɳ��j��/n��xK}a�=�7�"G��;�X$��>�a:���m���2�1��gG^ EY�T���SfǴ�9�Eh����R�R��o~ V�qH�:HޡG���*�{�&2Gk��QJ#=)��,��k)�I��J����o�FG��Yj�!�j����@)�-S�����t��Q�O_	�qZ��(��p�6]��e��{�%����!H���һ�K�GJ�Nd�_˖�ÁWu9�ꛆ;�Qdc%�q-� p���-�"Τ)�Q\2������*g�#��K�g�f�dl0�]5�JDp@q I툪��8W9�`�n���B�A�Bh~G�^
�\���o�
ɀ����^�o ��R��;�[V�z��-t��2��y  ��$�`�I�p�Ajq�Ք_W8+ B�_��&b�j�w��l�"�G�4X!Iv*�h�O�p��a��nN̟�R/�^��ս݈�DQ$�i��q����t����hְ0�㯜!�XJ����t�uM	�l�-sg��j�+'�0��:���W6qTHO�֤�.µ���ib�������R��> ���-r�C�9�7.Kk�b��>�1��	5�����jc���8��0F�b���X�{��lLC\C��`��߆�4g�3{�1/���_�ǜsLLS��K;>�*�����!g �4�!�B�ѭ� ҂#[FA�4&��ĳ-���!A��8w� ̀�Yi!���h\Є<�[�:-CA�_�'��Vj��O�5�dO%�j�Nޗ��m�z}�%�j��
L7��eȜ�M<��#�"�)Rv����zDt�J�`'��G�,Y�dy">�d"Q �8����ʡ<NSN�u�i��Y��%���u��D�f%#�1����y,�k~-
�Rߝ�[+R��
���~�6s�P�ԟ�WZ�+R�9.�H/
q%S �����EH��LP6�Z�G�wUo?��5� &�n��'�e�:
J�[��P�4�ԗ�W��4faggKY�f�B�������\�4)S��qP?N��JV�+>M������yU�жW�����ʢ�3�&*#�`�u����ÎL�����v8,+�	
��+wR������H��di�E�أQgol�#��+�b�U�L�
�Haó��+f�͕d��݄R��h3I<gE��9�_:��1��1 6-2����&�7�q���@@].@�D��K�&��u%�  ���Bu����	��4�s~S4�)�U#F2-�T�����g�\�1{}�E���}G�a /`��p[�q)_'g�a���}T�6����j�4����3��"%K��L����x2����J�?C�r�R�g�9�4�\O�l�.�6�z`�T> ���c�f0���RG�}2��r���e^e����G����2ȅ�