��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl����8KCE�=� �<DC"�6傋�	��I����G�"̿?z�1c�y�^�&k'�#�b%`���m(?Rq����Z��r-�f�a�
�Wᢗpd�f86،#ҋg�KpIWkj�������O�(��)��F8�i��A���<�ѢtL0u���g�в`.2��~^�[�.k���bIaN/÷�φ�d]���+.���1�lf�
�G_��������F�C(�J�K�wk7���6�i`b"����J����k���8��Y1_Ⱉa���Y*9���ܧ����c]���5��ð�����IJ}��|�3��1f���Wua<�dv]���+p}����&=ɷ�M�@vy�u���$����x�S�a�C�
77���t:�W�BG֕��#��t6E�+����&�A[���W̉!��yğ���^%G�Wا
x׳=�Gq����f>m����S�rN��#ҟ����%��--�kv�218������ ��Cһ~hebei�a�AS<�ˆ�W���p���}���o����wQ�f�}���~�C�.J�����x�����9$TyK)��M��#�m8��5	J��)�{��~�b7�e���Gz�W&�g/QM��Eڴ �ڑ؆|��Rik��R�oa��SXU�R]dZ�I���b{�cƳ������*3i��5�ĳ��7�n����bi�t>�}[<��j�\�/PcE�J���)F�;����f�c�*0�z%�ܘrQ7�f�j/߈	I	k��~ �̮=D{�L��o���s�m̥��9e{���$��ᦗ��`�7T�7Խ@��-��'`P6ssئX�%����v��<WOEvt�CD��dj=�����+|NW�uc!o ̾�G<Q�M3�m8�v���;.>�;�w��&ڸ��M���%��@ѳ�'ա�`�iW�F��m~<���H��̥kK����D��%��5.������o
�RY�x�@��E*Ge��&!�L$���a	��+`�u�1�u`�h}B"�����8܂�H�Czѭ8 zP�y(L}��T5�^�1u�cI_`UW���kۥ>������_0^I�o ���E��O����[��gG�z��Ї�x0���D��8��}}nT��������hXEZ!�J��Ǐ�K���U~�(i$ر�/A����.mfe����Q�l]=8Z0у�dc�uz��Uz$K�{�Ip�b�(8+�oW�M�j>qU�2�b�X6�i���p8}���o�t�}��]��k��
����f���a�+=o���y�"������rn��!K�9]�WD×ߩ��b]X$ڕP���4�L�Qp�vG�N�����yp�}i���n���7N���+DD|]����S�"'3s2�#<#��#���+��<g��h�D��s���@PEgf��S�����!��@�$�?�4�|_�h�\���(o�\s;.C���˵��F��q�:@�9�k.̄l�0Mp��#��M������f-26Ufo*�2�/�eF���H�Z��1���G��5[zd�N�-:6>皑l�RYDk���By������;?$���P-����sb�x�֛�
����'�����=���Z���DB�|�֑��NO���Gh"�c��!�D�~��T��e�Z�����XS/�E���:�-Ua���J��V\3׸����E�'�.�sL%��;[h@�N�F�'I��
#�:9��2�t�aU�(��\����Qr|�Tq�^r%��eء�����|�3�'wV��	��:,�ӱ]C�_A��K@�Th�1�] �蚬ݢ��� J7��eMLP/��R�*$
c:n։�(���̘ܽH�td�_wa-�H''��|��[w�))v?����yq�ڼ%�>�grxy�$ndR��W���K�	��%Jm!��/L���VI�����8�m���Z����jA#d�.��)|��>���pw�#BsB1ŃѦ���0x_t�����f�*A�WYt"��c�a?XW ڬ��C�Zx7�N��^Y�Z5��)V|u{W]M�$�.~����bSߵn+�	%�%�����c��p��������1v#9��Rc�/fvt�Z�IL܇�L�w-�:(����'��1|�*��n.�D�;ҸB{g-^�FM�0�Y�N<���D�H"qG�\*��̨Ne���u��)?��7�Ճ��Z4��Z]�޵�q�݆���U�0N������ݨ}<_K�3|&��R[0��57��6u6x�k�>qϜ�G����(�������ZWƏ�*� /�!�8l� ���q^��\kBi�(21Jic���s}�l[�Fcjw	BVP�[�4R�M׍���q��!#�'Z1u�E��^�v�	,�rw�1)B�g�0�h��!N��hK��C(ͦ]8�^�U�Q���6��搡z,��J�w>�!�i�+�`�v��ު�p6J*�II�<�b�a���}@	*��@��Vh����#��Z:ɨ�*)�\������Wn-.5�7ܩ�d�mQ���u����-�����5qq��ў�Ʀ뮺4�-h�W��h����'<g�:�_[d�ݾ�]b�����e����WX�$��	y�p�Pq�mmFܫ������^�)�!����=�88_���	*�IQ�.�����Ȋ�S�z%���[Ճ��8���'�=�Ҍ]�`��7q��jF��y�IZ)E#��zϭ"P5&!�!��?�:�$Q`
%bF�/����G(Dc$�
�Uk��2c���Wl�B�O���Em�a �=�ASjj���on���#f^�9��![�`sK��L4�T�sk�|.+p����ck�r�����}�ŶB1U���~��--���N�9)�l�D�Pr���ILT�a-��Y��#:�n���#7��d�_W�Ԯ)�-��0q�+��GR�=	(�jnsn�[���r2l##�Hu��/t��� `qͫ�X���0S
W[y�d?�_ag�&MA��6p?�w��.i�-8xS�k�Χhs��a��N�������c_=�S�>�'V�����r�.t��ᐕ�L��J�&ӷ�܆U C�JO��A�Aë�fS�5�;=�؇�C6� ���%��g���٫B��l��&�_݉����j�#��@Q���p�K�kJ�5G���E�K�ϰ��RPC啂XU*_� �r �ɔ�
4zW}~d�yO��(_v�^*0#l�g2Qq�iI)��Y�T���rgG�8������4ߑ�78�|x����MMmFY�n��Ã�ꀟ��'hꖮt�6W���)�{D�_�`�"�_3�+�{E�*��|�P��g���l�bIÏ}�()Å2z�Ӟ�Lߓ>~W��V&�dn�W�WNwSʮ< '�L�Σ)��c�'���f7��=d,Cu�q��kV����`e�Q޳Pm��;�'�
�[v"~�^���8w)�9P
&g ������n�'.�P/����6(�}��Z����
!i!��������������\�,~�jI:�%���{D,}����2%К����O|���%ٿ9�� B�n�ܤ��c�b��:p��[���o����\�MCzJX���%�(�:ǚx'Uu0����?��XAW�G�묎 *{r�����YfR�� $�X���+b0�t>nU�=!��0BnZ�e�`��k��0�w��j����#8���������� f㏇�4���cx%-��i�� �����\�Lw��P6��%��2���_B�����P��n��>�/w��;H�9I4���ϩWpig���ft����!��wt/��?~YS(�u,�~�n�-����h%�ʛi��^D�ƥ�����a��=v���3�12F-������g�ߧ�E�o��D��l�����|�i��%�?�ݱG1�/Օ�h����1��R���Չq�� ��ձ)H[��,/�I�Zen� Y� ��dvL�yƍ�@,��k�:˶�:�*E�W�q5S��UX枘��H�'C�*/P�`��	�A��RH��!����ݴ%�|9�憐�����a��7ɰ
�"UN��U��g/K���#���2�ذؠ�3��LeP#k��}������F����)9溼H�U_�8w�2�2ԩ�K.>�+��ypͅ|��t�b�Y�>��S(����~x���(�Ǉ-3/��B����{�u%��f�fPS�_����w�� �Z4�wdժ�c�h�Bξ{�QH�/�?!!c��{gOr��&q	d��)Ǯ�v��e�� �zX���7����E"x���5��\1�@ʧfl���N�yPG�C]DAz<���� �?�*�! ᷛϝ.*��VMN��J����|y_ޝj�w��VӢe.:�u;��yB�w����suu�2e�?��}������;��z�^�|�5�����H�����3�eX����c��Y1̀~��V�qV�4� 7�^�d���3Ԫ:�Y�4xed>��圄���*�e�}o�B)T|�!�!*�|�e�^ɝHo]�bt�,��������K�*�f2Qn_8,�<_�`W��lA�u�jE\<,e�(%��|��7�W�H/��0��}��g&��/̐�q�%i�s�(��g�p**�XD��V��N��l�[d�o�A֥�)f�=���«�(�3Y{@�g`���x�&��:�D���|pul�k��`Z��|?\x~��ZT.�t8>b��P�Ƥ|V��M5ߟ$�s��D�4�����T�@X!A�Lj�� \w%��%�-�!���p�d�	��/;�H�V���ȧ�D���L�ٌG�
[��#c-"�4{=9��/���U�^O�TtO�W3�_�BĀN�dP�P�������ً�DWx�!]60#d+��E���3H��Yqރ�LLT<�$@� ���a�"�\l��Ś]�]��]K��p,w
���U��r7c�@���q����Ť��.�La���6�[��u��W��w�R�N%��"PT
z�F�r��g���Ɓ�6Ƶ�:�)7�";"����X.4�y���]��9遈�2�͂N� ��`$]5-�[��n|Cy`�{�b�kL9uaӥ[�r�b�b'_�� HL�u9�D��w�t9�-��j��H�p��W1�`H՗�{��*)<�#p�	������)ͤՠ����?����^q��1m8���|��,��>˛�ɃAc��'�"b&����[Y0�y�*3�y#�+'y#)t��e�g��β>��O���a��tb[���I'ŋ�<�����!��ˀb�̩���I�H<�*װ��J�/߬���)e�rK:4�`���x1��$������c�F��%Kv��f��k������x����r�l��b	8����</�ܣIf�&���j��==��2@��Z���;q�B�0��%�b�fu[�=8x�N̆9a&��䙃��> e����1#��o4$+o��qՍlg5V��kY�=مq���k�V_�dta"�"
,vp���ٽ�v�_Qj��a4�Ld�5��y���J�pيuA��w:8�k�8�؎a��=,;W��� yѐ��H�_*1� CWP/;�\U�X���	nk��3�)�Y�l���2�#�`PM�pl���l��
�Va�O���[J�ك�{ ��['oyP�Ңd�V���U��&��� ��%�29ۓ_���lSj��C
�>w����VB2��a{���Y^��R)5���w��a{��,�*In�j��ݎWn^�@x-��2R�W��ˤ����p�G�8��Ł�"θ���򔑭�X�4����=Z�:=PR��ꏠa8I����;��]������+�����Fg����*$p���1�˳�cU)�T���- :ƕMi��v���o�=H���y��J�4���ֶTۓ�M�>��30c���o�K/��8�2J�sM�-9���S�5^�p�x ��IYPl,��kP�_���as��oxY�4� ��b�\��V �#H�k_(}O^'P)>���J���P�8�2��$҂�M;�Ag+�^������[e��R�OH��5:���$�>0`ر�j6i�C�r��t'����zx��U�k��s}:B�o�;)*���A���q̽�������r'l��Y��<}0��ĉ�hR9��;�
?���#�|����FO�����~�����ﭩr��FEt�޹�i�Ւ�B��'��}�_xm1�P3d9y�t/�Χ�ҙH�M�f�#	�&O�3j��X\��ml�c@�z��!������!=�z;7��(x{!뿈�p���N�9ΐ�z:ȷDЯ�Hn��@�h�n��0����M�m֯)l��q;���ődz9l��@[g�@Eϲ51��O׫���#�$�zgg�e'�I/( ��<ߝ��m�3k�@�k����S�U�������V���f���|�j���+���u��$3�`_f�Z1�>U�jĉ>�F�����=E(��i��;�3"�� ~cJ^dת�zp�ש�\�����޳�Ä�����2��I��B�Ik���^~eV������Q�ΐ%/�r�H��D�Ȩ�U�?��f��6C�00&�&��b��FB��z��f�L�{�M���V�L�^]�[_�Gj��aP�����t;uݼ��lD���I���m*A�m�Rx�[�x ��$�
^�����)�x�Ș��� T ��k��E���r�􊝔�b�޽�c���z5�[�B��w���mе�U���d�L,*���ҏŤr^��_��+���Y
,�� �
1_�W�۱�6��hro�O9�����lIX�d�����f��ܺ��/X�E`��-,��s�b\��
;)�{&�I]��@��
�&�[/�~j�f.�##�h@���;��v��>D��A�l�\���v�4;�>��iC�K΅�;i��A�����A����VDO��.S�=�0�S�b��L���,vIT�8z�l�x`ب�[HK����Ew��� л��:|LZ�N�W���5�n`}E�$q�8}����l�5��ZM[�}�N�n@��W��]���C3�1[�^cV/�Pw��0�?�p���n��֥�G�A�.k���L�E��  �L;$�:�+}�6n����;� ���֤�Ϸr��e�3��E]Ը ��ϵz�:��S7�*�͝�!;��3lhqm��=���f/aR�t�Ri�r$��]�ƫ�A� 0��+��X�zrn�D˾Z:��^Dvj,��P�ě��Z0�����y4X\�NX7A^���f``�Z��}�7��\$]��O�ٙv��O���T�_��[7�_����q^�&���E�/�N�XQ��0o����� У�Drc��w'�:;+L���� h#!�"��'�iП�ĺ����UF�΋B
E�+2�z�o� ��e�,�g�?r ����9������ԇ��@Mm	��Pc��_�1^�;���G�H���(/�����K�)4R��84W�X�N!�����������н�}������̪l�����}~`~��
�J���7N���>Y?+P��qSx�,��i����8��@�}���e�s�pV�!!�a4����N6��b���O|=C��W�:*¨�@<i�'�!�2�	�y�_j��t!�c��X���Va<�R��ʉͷ{{i�7ML�S��I��[���l���ϸ�#��H�I�&߫!�l���s&���6��1���Lvc����#L�|���ͼ���Ikz��$�eUa�Q3����Uc��QV��b��خP���^�8�?�$��]�/��̲X"���׫za?Z#�D�1_(Nz��ii>}��sR�	p$3��UQ�Ci�C�v_���&���� O���;K##�r�\�&��2M(�ƥ;L�o9��dh�i�r@�7⼡b.*��*U>�P���U�� �0kU��������L�ʋ~�9o[�/�7&&0T������#? ���E����}1�����T�bkY�g]�yC@Fh��t��$P4܃����aʧz����)�����"gFQ��!X]�a�N�U��܌�z�dn%���9��FG��Z�3�x�h�ۍJ�/\��'��}�O!�����%�E�U :�+ߒQ@W��������S���$m��t뒽Vʿ���WȞ
m��H�5�ϳ�Y���bw���`u�)������X��?�D;���(nMI�m�� G�������q��i���!�Ws#ķr0�ի��w�ބ�p[}|�tzV�(�gn�F�)wd�z��Cc��8g��И��̉�l�myYR������ �@�I�Z7[�x2�ah5�`z(KF7[�1�A4�������&�"R��ѽ�Ϙ;%+T�3qB7�:�p'�$)� р!���t��g��-oe���ҖC�� �ԉIo��k\�פ��uh
5�P�\|>�M�W�����I�%աz�4lF#�F�;q5��8���J��bKg'���9�M7�P�� �nI |v�	���ݔg;�c_��*d�6<�Z�
��,�f�a���@����K��0{29_|���[����ؘK���xG��cz�����U����r3�
2K^t���Ia%/�WV���.�;�A8`wk�3l{� ��ZoDΪ-�wT܍�.SbRô �͋��I½R洹�X�1TI��}��U�Ϻg�����������A�]�0�4�d��10'#6��}�����K�0D���˸W�����~���nP�����Θ!6�a�P˷�J�*�|[0&)�g�o&���ɻ��e�2�ٌ��6��8��A?z20?_�̷�ܓ�w�Iu?Uəe�,��{�&���ow���S����K�;�~�5�k��0��t������ߖny���O���転z�&&�!��g"��h����0�0�/�5��#V�";�u����&C�Uc�*W�T�ʱ$T�Eu �K���\�I�s�Yպ�d����`z��H�2D��/[d�~1��4���D��?�ݹ�8AޡHQ��-%�S\<x\$�����O# ���;�L
�@�|8�U�s-G�ď�'���e�Ud���a@���~tg��i��7��k�5|?�L�@[���Z���A� �b������o1WwaT��=O�(c���������3�gF�k ;�1�v��NI1��ϙv%sL��cX�+�ED���+q���8�Z }�x����$sCqJ��/9;nee��ۅ�OU���̆�p�<�vN}z��Y���;���b�:����
�M)��x�d�B�J����}�'�BO�Q&D]�B�i�t�]�N�uBD�p�\���(I]���'Y3v���p�&����*p�	��R�F��4Vh�g�9��¢V��+G��fu͜d��z�*-ѵ�V.'�d��q����е$5����CPY����a��� �;u�nV�^��P�}�w	W%��*i��YGpfL{���#R��i���T���j�b~�*P;�2���i�
�#��^�r�B�{#<e�����Bu+qH���J��[�#����RC_��rg�����^/�l\6���ޯi*H9�6Qg]7,ȵ6�d�XF$ohM�Kb�#�}.��	oN��H�D�G2t7�G�$�d���L|�_g;�j�/�zq����f�,|>Q���eV��l8ѥ-��aF��eQ�^`M�v3e�k����4���x�m%RK>�Fԛ�sK�V|]�hGP���/gR�����62=Y�� xI���v�r������a7n���;yf�o�i,�E�⪾"wo�}:Z����CDd��jy�6g\*���䢪$&��;�ש�P�6�������8ƛ�+dDvX&x釵�������!Wi��t0%",n�㶁��W;qE� -s1h�qR^}���%t�T���p�&�՚@���bw|�Q�.�<*H6&��-.��ўU�E�Q]�̡���rՏ-���tr�7s�[���1�<�2��XH{�:;��2C��C�@�O�J.&
yHpױ�4bgXq���C��u�9&sS壑w���d0ؗ��\l$�}>Yg�=�\��7���8����M!��K�C�T�:�G�����$P�Һ�:��i�A�G�W��ą�Iv#�4�-a��tZR<�Kz�0%)@G��nT٠]`W�,>�pAZ	W�0y��!�H+��Tp��H��/D�nXo.�.��P�6`]�0>>����܄�-��!TKN�f�z��ʇL�-�d�N\�_�.dt�(�I�d�V����>�t�U������w$B��2�*�G�H�� �I�}����f�#g���J���,���'�]
��u-D,#�����:�'��l��Z�d�60�:���\=n��Qe��6�L�h���n��{7�'���}5h8��B@_T�u,�M�}t必m���Ӆ��� � �_%a҉�Թ�ұ����]��vs'�[Z��C���ι�Ѿ9ĺ�K8Zi.=��waOl_g�E�v�:��w!wt���^���i@���XЂ1~{�6~���;Xj�ұ��H���9�����]F�w+�����r���[F�ګ睦���d1�G�|S�`7-��$ �y%ECoO�M+Y�A�#���a��`\8����8x}�3&BgI#�
�T��Z��ͽ&0�(<)�@�w� 7�B��YF]�Ԇǥ7�@Ǧ�)w׉� �5[�l`5�V�N8^�\����$@��!�x�)����K�Ce�}��z�wj���s9~��(��`3�/~n�Z��z�ּ�YS|DU
�8z0�������C�G���z*j��7Y�lxK�Tfr�J���5��kAn`�,�)dg3S]ΐ�noO���⮾j��+��k�丐�Nظn�JD���ɍQ���>���ȼזW�N�i����*�7hw�ŰK>�_����ߜ����yn\����P��Ϧ��eL/X�	F�:0��A�c{pjf�|�<gL�Is*ǭ[zZOu
Ԗ|�9�!g!t^��RC����T�t�oRJ���xK�3`����:�fP���{\�@�jjX���g�-$a� ڎ�t�� S!O:�Ѥ�G7k��h���0���
�D����M(f[Z���T���6E��&�z�]���^"��@K��C>9�Z����dÜC�[�x~G<d�[qfR����%6�3ù�+ۛ(L^n�g��PR�ؑс�>����j���]b��j�+����|F�[�J�>Qi]T�K<�Ʊ8Ãtn�+6��hVd�9��9��طt��s���O+as��EZ��Z��C�c��O�`������'B;o{��o,h]6�.�j����C�o=�L����<q��j��h��M��H�����;ؽ�����%#�>�@H~�w$2m�OQ`��NX�����-�$_$&x��Ve�H�F��"��[��#*���_���ɯ�o����G��A������:T�m��J�\���;Q�\{�Ä	�b��a}X���kCh2�;V��NCLRnڨ��1�j�XЉ�2W��vm?,I(/y1C4��1^�{���7�ʃ���A�<̂Äv������t-h�����DCo����(�������K�D��G����G#�:�0�(�E�E9X\q�/�I��KD�$���=�b5HJ|]��is��I����[�u���"Bg�|m����~�i�19ëׇ��@��#[�;�Z��߈���"��8)n#K���C�B��/�o�/���YP���O�
��~#��^U��Y����:�F�H�� ��	�G�T*�@z2��BF�&]QB��ӵg��K��<��J=zw�j�"�S�j�Ȥ��2���TػM<�O���걩	��ɟwG����S�πĆ�*����G �s0�aJ��m����O�Y�̫`׼R�F�u���I-���\&bvq`PH�(j�f���o���_�d_g��n�Wa�]4Ո�F���L�kU��~�O���[�d9��eA���ے@�􀗔��l������R��5���`S���'����/���o$�b��1J	`�-����6�L��'��\�w#('��CæQ��Qb7�d��n'��bֆH��DΈ�0hH�����r\YLD�Oٷm �$#�*�3�7eQ:�Y��u�Y�n�6��ᦊ����<4��y�@ ׏3>8��Ω���y^l?��2'��:�߭�B��A��-��s�'wUDx栎+̆ u:V�[8���*5z� ׊�|���4?bA�G�Bi�~Ċ��1����ȗP�� ����J���a~�`F)=�P�4��:����C~z�L@���۽V�,Pd�̜�
�A7Ϻ|�:�zޙ���GQ�Ϲ���(m˳����/$+�A\�uwwa6_B�#u#~x�ZL�݅���ˤO�.UE�DƪO�K\i��-#��t�GWRM�l����J;�k���/�sγt�%|�?�AE$�Ҷ�%!�u���fO�|>��4*��k��)����U�2�<0��v[J4_ú�
6�?y�;%�(6�3q����4�R�Τy�Ji���u��k�`�����<�� �[�Fl�0O�r��n��w�O��n.���`�H���A7��[��E�3L��,��'�@�E�=8QS���-�3`���VG���H� ���d�RN��j� ;���S-J�ö0�W� �9SW MatiDM"�藿��xh�r��%�J쎄��p��u�ɹ�N)Wy9�ל���V�����2�֧�����'�^�T&R�'43�p��˒��]�`}�l�l���$ɢ�S�5�?�7��Or�ì����a�+Ŏ4���gR	v$ ,Sj���!�;�@FR|��\ �ѷo�?���'��ܥ�[�l��D�]N��_�$>�����*�X�ڻx�٠�[��!��~�-h��U��ѲK 2;��
��0#�x�c�{X��&���J+���Q���Efs=Τ��B2K������:��[�,��(��H^�
*S��L<:3z��u�#���:���y��|��= <�:�pC�J�8��mҞyp���$� z
�7E�+����_9��;�ݶ2-��M����R�9�p���l�BW��F��|@#)i�H�^��wP����^�#B��=y81���Ci���I�g	Tom���2(�X�4گ�����h(�ibrQ&�2'���0f�@x8߅�|bҤ���f�9�|�P�q;8>�5 ���[���V��VS:�(�Gk[o�ʘ�<�1I5�o5����$JjN���KB�������)S��ƟO�Kל �po8�i�E�ɴ�m#?�𰞰eW��H�S�׆�ɖ�xS=�����Yby���t��B򠖲�AEFo*EL�ڛh␰�aG,p����W��� ��p�<6ח�>"���/nJ��[�B���������E����Q�o"e^����1d�WX�e�d&ެ�xa�C���G-N�7�*�u㑭�o=�T{��W%��e~+�G5=��s%I�As��- �Ic]�6�*;���%@�(+�#��ւ͢��'9�
�����ooA3�
8#��\�|�P����?[�b��i|aj|H�vҳa����~;Cw�����߯ۋ%<a���q�<Xx�6�`(!�-H�hگ����Eb�B�M$K���@˳=��ח�	 � �U����a��h,�A�U����ҁ-��ECU�a6�7�a���{�6#�1U�@ꋸ���S6҅I4%�}��"��b���W�� ��"���b�	�Y��S�Phz�y�6�b�8�g��30N��,Z���T cc���c;f<S�Qʐx�x�[8P�Px��;��Z�B]6,%�7�̇TIc~k�f�a��,m���6+:jtMǊwMՙ�zz㯃ө5rL�L�ls��K�Bwˠ�^]Pſ�iT�]d���$F�a��a���7~����z����a��B��}G~�&u�<O�et�)�#'���|�����rfU�c�f�����'=F��v��ZD�p����edK�eJ�����u�T�-�ז3VG�jX�i��Z �t|�{���y�[L�6�e��T��MZ�^��w[,��|�dc�@���Y�=�Y���e�P·ؠ�#8���O1��_UԗSh���tK{��B����$\N��u]E��3�N�����M���X�����_��p�J�[f�Q�Ծ��*7�O����L�P���J�{BA]�+�J�����=�&�������U�*�� Ә�Q2�����'i	�f�4L-�Aܥ�����X[գP���֭j�t��gX�BE"��!���/uKҲ��ɌM�O �kz�?Y�4��-�$��H�¢�V��B%y��r0��t��h�
b�Zv�#�Ɯ��˸ S+�`�{�/eA|����s=�o�����"Ǖ!��p��T�r�I^��z-�U ^:j���S�S�r�,���f%��V�%�� �O��>�E�
���<?%
��?�P!�dN�v�j�bP�~qp��tH��NL����q�QZ�2�C�kˈyxyZ%�R���n�ߤ��'���\�:�0g�Q�7c'�6PO��yl�%�k6�Գ�� ����N&���&#n��1i��Z,Ա�8'���?������[���/	��-ݬ㺚��c��sx���8������J>��8i�G#c4�hiz������%W8-��a�����<��g�y��x۳h
�|e6��o�,����7"������1�kI2�g	�L�c�=A}
����䦀�2�s&R턅4��6�;�a����zH��f��jI)���|ƽ�U�l
y��	��#���@N�c���o�2+�+5ۭ���'=�Q��(��~�.��	&&��B�Zr�L�$s�p �%N���#�z� �^�9���q2-��r����LE�{E#��N/�M 5�K�ȫ���$$��-� �yc�yv���fc�)'n:�牬�4�jE�q�tթN
���<'NTN�^��s�4+3���݄~�Y��VJN��w�9����J�"�>=8���3��d�p�mu��5�9�E�)�N��2E��}��n����F��x�e\�PƜ6��i���G
���\h0������T!�W����M���?H�j�HgL�e�'��Y�j�^��M3��
K\��y��	Zg�~M��[+>i�ǲΨ���~l�=��:va��M���0�D�/����` ,�t�/o���&���<����?%ݳzڎfO_�b74q��B�V������I��9]J�q� �Dwhc�C���|ܟ>��N��n�i�۱���m����w�y��~d��%�3T߼4�G�9:4����':����V�^��҉�Y�RUq�Hp��ϙ)k��2�bK���C����>&��D�TG-��\�u}vɩ.9�]�2x�` <����ҳh�9��@�L�ֺf��&䧨dl����~��c�>��{�ľ�j�"h�L�*g���.���u�3sMX��*"/*���.4E�\��63�r��lٛ5����� 	�#� �%��y�=��#�^���g�5��*����O��x��	zD [Þ%Ѡ�B+j�A�iğuV��A�ɱ�l�N�!�R�YS���Ő$�!��S������
�rX��ޫ���p՝]��q�t=Na�¨�\��t\�6Ԯ��NpRz(%�ӵ;}�®�<\xGN�]Y���Մ_Q!��e�� �;|�`N���GG{拼��Vd�x��
�3��ԷݺF9z����I��Q���?Q5+�����.����Z����`����,!G�HYZw�zR���:�ľ��T��j�E�!�O��w�?�M�},JX3�����Ѫ��
��P̟����y�3u%v9k�X4.M���
	���WO����i��t��pA�Qƅ��	wF�7���ٓ�oM�Y<�i��hk6� �B&�c���
�)�ޥ� ��5j��*L	R���B��=���cQ��D��[�F�[��%້w�ݻ��l��ڝ&q��bP��_���j]tgPk&	��D�T���I!zl�o����B��ǭ4K�ll�E1Hs�g�	��ْ	M���aC�31uQ/b�,dP1d��e�'%�w��hŭL�}-A��=�l�y����Oqbg� (�%�>��e�cO�QAd�*�X�\3�S����O�=�O�mՐʈM�+��D=> ����D�V�T���3�~L��t��/�?��ޜTp�2��l����q�H�??ٞ����N��1���k��|�q��w���3Z���x�@'!�)/0�+L�\ɿ���i*㒎A0���`}x7�u��ë�0�{װAWZʍ�S^Lwjն�,�KW,��d_
ޡ]���gv�'�@���8�g ���n&��ҵ� � ި���WcNjq)��Ls����~�h��/-.��� �@�#���Q�W���o!����o���}AB�,�/m��l��O��\�.0�y%>¯-��o�H�u�uV�l���7m�l�i2�E���a-�;��n<	8�;*��jR�U�Rƚ>����d�=cӎ��6Ђ4�f4��<��,�VrB�!ޓV�����XUK̮�{�+s �;�Y/q`4���$���<���L�^���@�Ҡ��"���������:��3�P�h�1W�Zյ�}���Q�"���v��Lx�?[��������Z)�Ɛp�F����.nRc�r��#/�$"\x�@0���f���*�P_�pM9[��I��&Z4���;�!�(>�����;R��2��w��SI��0ƫ�M�'@�R1a	��(���\��s(w+hDϑ'pF�M��?E��f��n��\oȚ�Ǉ*�o�s3 _�CK �nٯ0�[#�!:{�9���g;���D����l��A,�W�G,��T����HD�G�{��S�|�4���-=AO�>}w��U��pS5�^7����}V<MfM��DښX��k��[6�TP����-�&�V-^����i�8~��$����PI����u�h�E?��~ �Lp�o_����h�Y��*
\5����8?�/|{^`�|���5e�Q����#r��<��eS��t�%_Ex�:@z2�g�Y2��� �~)���v���By����P62NQ�z�8�'˺N1���F.BMl�o����S��T�>P�(g@Q���J-K�����%U�}?ՈHi~����]��:�"�Fa�	D_���*������L�S���6��ճ��/��a��q�_�a6*�7�u�W)_��ME4f�Y���J�E�{BZ�㌄\�5�t�0<���2+(y5r�F����TK;�l�d��U��S�$#���<�E/&�&��sH=�M'��#b����9S�Ó�zD��.X:�ll���0w�Y�vU]*'0�t5�j-~t��Q��x��ژK�+�@��ϑ���д������d�2�0��G1HP!ؑal�C�z6`>\�_������wB��(���ܺ�iwЯ�M^2:�[q�+֛?r���8�$=ʊ"/ĝȮ]�4��=���D��t�#T���g՟���'3��P�}��E-�܅O�ʪ��>٢Lk��q��uO.1���+�NFe��X�H�X�H���h��nH�;gJ1����4�b4�Ղ�3�6>���D*݃,GM�@T|F�e}u񒐗��E��YN��x�?�"s7H�n��ǵZΥ=��s�L������|+ƄX��b��o�"11����jDO��V�H�f��٥N�'�KH&�Ə��k�Q�(��n :�呄K���ކ�n/z�~lw)���+�y����M'����тn�2��_r0_ۣ!/q�֕=oSsn�,��R�L��[�q!�s�Cu'3��2� ��;gT����?�����h�*�'e�<��[t5�_\n��!�Hq0 ���j��8����l��?H�0ʠc��R �"�����p�9���u�T�R��m���:�/�J�W���;{!�a�hPj#7p随��maAZ���lil��W�4�g���8�
���t*��e]���b��W�v�g�n=�w�0�����X�-�r�8SB܁�[3�b���'K)x�r떐bx ��ݖ^��:�,̫&L��K�6� ��S�����ד`�0j_@�������Sڟ�ohv �F��+�9��2R|�<��T�4�;K�&ŇT��n{�f��=�wt2�����U!h��L�ڨ?0�>(�^$�}�؇,F4��1�������z� �ta�ҵhٰ�*��q¥z�H#1���jUZl�Q���6H~}iv��~������ �l�\y�^��c�I��-A��fǕWm �=Ǜ��`ر=s�	��D��� �]���o���E��gk��N9�f���	L9��M���B��v��Q#�p�|��a�X0�3D4 �R �X~�wx�����P�����A`��D�F��'�Ư�t�",��x4�yp����4ұ�:U#���!d�r��qNA34�N#2K�r�I�Y̰�b�c����ن~��%�F�A_ G6/��T,�o�?��߉O�JUW�*��TdG��|'�Q0�e^k`Co��P�դ`X!or��3k����g	AI�Lo��AcI�BFoo��7	�iM8(�g�dٚ������1�U�.m�E��98��6����@���? w��K����2�ϱ�����B�1�� ƨ�_�,���in���E�����T֦֔9R�>y�
�h����k�/^��L�vŶ�"�D!�@�k�l	%��Q����e�/�0��zD�?Z ����]�Z>��J$�b�4�*�{�dd�j��5���N $������v�������q���9�iM�r�
�+�u{� �s����}��W�ѤX�J�H|� ���Y塜�z	a�������
(J�^	��"|�2!�AL�sS�,\��v&�sEG�5K����$[}#��ìS�Ϛ2O��@��b ��ї�Q��R�ݢ�6®0X%�8�(��a�~�I�S�p7A�����h�=5����9�.��Fzk�^�0�N�����li���d­����@+����6�TA|]���"|�fd�#0PxjŇ�b�B��In��K=�!/'C�9�l�K>�y���eX���0�p��w����q4i�e���ҷdLe0�	�_�g���m�nf9����Ya�'�:C��6��2�0ߝG��Dpםl�#<x��&DV�������Ye�3y_mrl{�^���nR�}wЄM�������THk[�&3M�y����w�Џ�d��g�X���|�ΒP!�}�O�H:��m�u���m��� ��k�Lh��%i>ә��|�dw�CV��y�}�GV���dÞJs�j��ā��b0T�C�aA��L(�����*��]��=��$gu���g�FM�۴Kcc|�	Cy�J���tP��JM��K�A�5ю�<Ľa��o��,
��^�R	cv=(�q�(����*�eK�.�~�w�0����*c���[��d��8e�F�wi��'�m��e7lQ��&2�׷QBz�Cŭ�.��B�3��2&�ivn������U���������{^QBI�\b$&�Owz��K����Q�y�>nѣ*1�Ns��d���:������#�|�����.��сU'](�CP(OuQ��J*	AX�z�΃ V�Ѧm ���G�A�y�:���?���3�iiP˿��%��3RwP1�� [��_j/Z~��d�}R�ţ&K!��::�魶
k�9��7�|&��M�B���B�a����S�#�w\�����"��
�v�+v��8��F��Ȓ�a�	��q̨��DZ|�H(�I�ͻΑ~%E�DZܛCpb$�H��ۋ�v��7�8/��Z&f.i��	d�$�!i\C���^Y��o���R���#��R�CF⌭!Y� T�>��Si�R'+G�-�q�A��U�I��=މD߈�1����@�{& ��t2w#>��DA�`b�ŉ�뙻d���G(g��:G9����؋�6�h�j�oû�Ŋ)�Ǹen]ɣ7��j(���֢uc�s�az��=.�B�~���*W�E	�=Ǥ� �����6��Q�C�ߓjN��&�|���;z�����U����X��*�H5�� Oԝ��(�����51ɲ�[���8jw�N�m~��̒���$�{vi���b��-��h��������f[�y�*]*'J;2����T���?Oy��j�B���o 0�)<�u{e����Zt�X<U��ѓ������`.*�\!��jI��L�/�둘E7����m��>=?�cԑM��0ChLo(��>¿W*%\�l�*�XYԽ��^���rS�꺺~�)A��6����4�r�>��p_��t^���a!�q��k��׾�ji̟߲3S��3Va�cl�)�/@�w�G-�O����4;q}(Ǻ������p������*=�����M�J�4�|�z�k��Z�i����0�t�ʚe��0���Y�{8��2l�B��	�������Rw����h�o��5��#�D԰F�e��������J�I�����x)5L���o�a��������;.�Vw�\��d�M['ڤ��Ng}%/Ǖ�>��q�~��8?[s�o2�d:Z̑��o��%��tI����*�AZ�H��Ofa��6�jӻ9)}����b]*�����~��A"%L��������t<#Ps�&����}D�yGw���"�b�l������ )RxB�����"�ߘ'�f-Tw��ZIw��W=����a��[70&A=5��S!����r�0K!����Xo��CD�����LY~��H.<�yT���� ���!��ȑ?Ҭ�\���v6A�!�j�EN��~���C�UA�����{�k�Y>���p^���+�n��h�qɠ�C���?�A[2�o�.g�!Wk@pЃq4VPHdlD�U2:��u?�l���*r`�x������6ՙA<��'����_�a�Z���fH�����(W<p]�$<x�̍@ޡ����D0���3�;����6 ,՗�������kX;y~�e#N��$8@VC�U�\Y�*��Y�(�)�@io�ZݣEO�z��~QX$ �ӎ��>.'9����@ϵ�:]�z��w��K\�R��@Ğ����)	.�S�ȿӹq��o�E����/�۝Q�\�p�:��˹Ȏ:� n��ɚs��J6{��*Q$69Ͷ�X̔r9���:�?$w�GW$3d�f8�i�]�{\���%[�ŜOi��_�+�<#�O+�"ذ��v?3v�����V�,����B4/s#Q��=9�d�����a���n��+�6�!$�qn'�4��"����> ����ɡ �YRₒ�}�>9�{]���."� &o��l�b=đb�#�"�7��,�<���!�U*8���H��e���=�^�r�ʋ��P�g��?	� �a�(2%FT+����Y����� N"�E�tK�eY�N�%�ȓDV:>���V'|���گ�#� �򑾗���u���� �r��P�hd��
ViC�e�;�]�����\.+{{��c��V!�zi�'tz"`^�tt�㩏k��N�Q�`"#�&�A�0���nc�4v�^�Vm��|�������$�܊$;�Ĩ� ��l��3Z���4�\��ZX�wld�g���BD�0�0�3�"չ��Ŏ�G��C���k՛y���V��� �63,�$=�j R�a���"�PV����^��~�-効O��L��M��D�����]g�>C6���=T����8��3����(&�׽B��(�(r�`鍄K�(�ũ �I=E�� ��,�A@�!�����M�Hm��M�r�&z,n?�YYV(�|QŲ��r���0�H��1���l�p�/�+s��3���g*e��������!tY���X�>l\0�}�u�b!�S"\Ud���ttOW�2�0�)��)ZR?��Dx[�9&���c\c�憜�2-<Ǟ*(G���y��)��a��7�ݝvk��y�9SV��5��?Z�ǋ&'�.���޾�;�ZgX+�O�d�"ݍ������T�uŵ�N�d���-1k�@��ߡ�{��	��up0Ic�����:ؕ���U/�>�!��Q�S��e����_-vW����3�qR�h���24�_Z%�#M�XږZ��b�aM�)�|��#7+�hD�s[`ؒ��"xu���Iւ�K���epT��Ö�R���Y��5�TE�H�".�))[
I�멺��KzH?�m���,��o#�;�3��9YOa� /��s�L�y�"gT� ��
�~�)d�H�������d�Ծ������&�y�����+��>l6�*V-�wN=�������$��J��.�)���u�1E%��K�����sŷ;�8wC���"�Cm�q^��G�X��>��~O��3���H=rBљvW�X%Q�����jRG�<��
 o�	�X��
�.����Ե:q`#G�]:M7I���\o��Ɯ���%���vp		f"�J�NS */Y¯b�.�_��@�ȶ'�S�9/h���, �u�zJ�����s��&Qn���)��r�Y�!�	���Իy'T�ӳ���b�CScb��ա�5N�ŅY^�=����������oc��A�l8׳�#f~�p��c���sylv��y��V3�5bOCCXC�Z�>��mP)��Y-So���j>O+&�Pۘ��ed[�Y7�
v��Ϻ��_;�bB���kB=Ck���I��sq�cן��5� B���?�9�j33~ �P��?�Q)�a����(��*�P�Y�Z�̤W`�M�ބ�&�U���|M@;��Z��kf1ˏ����-'�Fȩ$,�	�s9�P��%�ι6i��|Sb(���&�е�6��%�oC��>l ���tꜤ���<^J�&A����:��?~�&MYā�!ĕ�����t�h�^�M�nKd��̦�M����AP�#�W!$��?��B�L�EH1ʒ?�	=ԍ�7Q��.��?ۈ�:�1��}��3��N��0}c]%��M�]�e���:����c&5�B:U�tX��²�O|Z��j-P�Wf�mwG�;����0��/qq����FS�J�$���0�쪵 �W)\���9�id��\`��Հ��8�?~�l��7y�,�?��i7=�ҵ;cI﨤���w$��?�S��$<�H�#�h$`A���:��ӷ��M�5	%�l�P'����q�q���)v�h�؃׽�}��qq��Z	}���U�tJ1�B �n���;��ZM�{-c�.�ߥ8�񑆉����='Q����\���H�~<��C�S��3,��>�9��=����#�p�bt����������m���ʭ]�������QY�kS�j5�6&Ĭ4-�������CV�p
p=�	ɘߣ_Iq>��@4]ѹ��*g��>�s�h�(��2H��$�ȄӵU�>g��/� �W�%���Ǵ**d�d \���u�Ҍ�}�n�WC��3P����X���|�n���v�1�܂;(w���7	9����b���vΤQ���t q���n-d���ou�%~�\��8Q�, ��b�Ō&6{���Ki�>�9s��{^(��sx��"I"3)��>�R�W�_��c�׎�!!�l}��/v���-�d�_�_�o��Zx�kd��0}�3�9HD���L��/O����0��J�l���;�^�v�&fɪ%��3о*���n��.f�i?T���C���G�������B��O�Zs��|���i��E3;�� ��2�"x_�W M��ZQ�6z�:Bҵ/�����-�|~Ϻ�(q∸��]���l���'����,��	y�HN~�^်3��@�ɴV��)ڸЍLA�ؓ!=�8�{�֐�ߛ�l��:
N�X⼖�BS
�V@:�Q��u"7v�t籥gK��)D�I �X�(��Dg��ܺ����q�j|�"'�X�)�	B��������_q!>�H��!R	c\m�{���_y�i�� =��u�'��W�0`{H۷;%��ʺ�õ�e�#�����V���y7�`=&��K,B��,�=��+ʉ00 �ӫC�)n�JT�g[��[�áq�xo[������� �����T��Ii��}�ϕ)���_��kW��ZՊ�Tٟ��P���R�P?ďa[U��R
���`�R�-2ކ���� ॱ��>�5�3Sk��$�CO	���UEa@N[��9b��~��a<$�̂�f�~��N������1��T����/G{(��x��v��ݯ���q����MY2n���F�(�|fC��+/�����*���H�T���>��+R�! ����x�;\x�Mr?`�*�s�U�AB���K�ۇ�g�ھ��|y�K+0m��;um�n�?X�P�������������}b��cUo����T�aP�a��c�W��p7�@ݦ;�Ğ�bo�9�g�j08*�rBK��k����Xݻ^�j�]�?V2.��]��VA�9%5f����[�������˂Җ�[�'u*��H�(ۏ���;(
��1�}�9�泧�����E�ځ�ʎK�!�|��7b �Ϩ���=���{��P���\�QGʳ��Ϙ�.?�9�V~��d�������m�Vx��]�&��3������tn��L@���u���G���܅s{$c����S������
l5�|Q�N4���ƮʨZ�:�k{��Q�iq;�Qick����r`�(�D��Pg�c�[��@t�l y�A��96x�L����G>=Qa�>���K5c �����'�����-a%� p������h=Ҡ�(�u�p�4UN��.���Gl*Cv�ρ)�Td���ө�?�U;�#�y�� �ז��Q0��'o�82��д�X,*�-��F"��L �;C���K� g��܍�s��H!^��IWo��b�fC�����}A��h�>�����U��c����]܊�s��O3��*��E����{��AV��2�~q��%��8�s��F�����l�҃|ή�]��L�����M����$+3;V����TgW����8h���0eiU�3b�����W[8z z���5��^{	o��ň��א��<d�r\�;��<�I�>Q���,��K���Ϊy�����q���B��>�m+��>Gj��y�H�6��(/�
d������{��z��K�T��Ca�G����� ��K�t,��
ʢή+�L����}V��5���������6@m�̲c�R��;<������}|1u��v�����^�2㿜�>Q���:d���ʵ��7�~v�рUʪ|����]=e��#��r��SީaL�ޡ���2�*�+�"����bw*���Ӵ��c�B@��i��jVawҋ-��O��3�k���� �11y� X�"���Nu��62����ڟ7R�	vl���-it�	sm�},w0W��P$�@8�޷b�����/~�],"Bԉ4�W�D�	 (�v*q���3z��md��yCG~.�¥BAw`��Hh�P�v43���Ig@D��Bܸ�&�L��e6a�0'_�*�M��f[�}B#�
�E��{'�K|�~�S�L�w��,!����t�6��֏Y١�+4�RH�ו�����K-B�m;���JNB�E	��Y#P����%��ώ��0M��/C�޲t]pxd�&�b��
��dLhI�v":�B7VJ`�����J�һM'�܄���sI�GD@�@�N�Ĳ��ANǎ;�5�Dx�4��#u�
�@0��z\J��������j��z�-�+��5�W0�e(hx*q�H���>ۡ�/H6�Wې Q�H�}%y�0�D�����p����4[Sd��ɰ�/@3ё�oB(W�wH���yI�mC�!�SY����CTM�����t���K�3���p����	�.�7�-2��b��(Q���顖���.�a#�?h��9����K��Ŋ%��h�ҬV=�O���u� ��O�d!�d��Y�6��{�>~��0݁���y�g��>�y���ڈ72���*s�.�����k<�H���UI,,Ɖx�h��F�B��g���@MVµf���ΎS |M�@����Ob �Cw��]�N��C��fR��^7*M����}�U�B�9�{i�x<u�&�N�|vB���˄o�7�5 ���K��t#�����*}��Onm�'ny�<����i=Y����+P�W�z�����s8�ph�Ȑv\��*��L�'¡T�!�b��#�{�g��A�?�Ʃ�؀z��ۻ�f+��fAwN_��V�͸F��_��h��%�U;��j�	C���%lCjD��(C�G'C _f7�̸N�I�����J%}����c�2I㬦�O��x"��UI�/P�HR�Ņ(�dآ��au�ޭ�#���`f[�o�����~���wc�@�:PT��6���S=ƽ0��äqi^��D\V�<��A�\��aw"(�կ�S��7��z��0��!�a�t$�u����CI2�=r���sɎ�۲$B�i S~Ԯ ĺ�0�@V�� ��q��m=�ff��.^��5iB0 K�B�#>��hڜ? ÓS:ӿ���V�	�u��S����_�d��6A��'��?�t���ڠ^�z��1�fyu7�(Q����Y��ݿ�Q�|���_���q�s{[IA"]c��*�שQ%��]�kR�\�W�]�|�g��8�Dv�;�n�*�nrr�r:p)Jt�|뺂����lV�goz�m=�(3a�E�1���QM���I�;6ß\��)�V�"f�HH-q.0��-��⛹}@u+@K�2��;^���g���Ğk�=�_KjK�a' R�c$���Q����X�9"��.��lsM��9]� �m�_�U�V������`Ln-��T�W�_�f-a�-(�P̭P����Q����vlт� ���af-�K#S�<�ύ� ��wh�oZ��N�*0�-�G��
��s�~;�+n�Z��;�J�_�WJ�'�m��8�1�N�k;c���� ?g� �Wj�=ޕW�]E�࢜�.6�Y�25������Of��@���i�TMl�IL
�^bp٥�s=�<���in�I�@��D?�Q��]����``�T�ȹ�S�/��TE�4�A�n���t��n��іB�[�8������v�U/N�[�w��ѕi�j�ص�AP��A�̌(�5�2�&w�Y9���v�t3ǉ���U"�	�h/��X����Xׂ/>��4��*]���t����S�鍘;�l?S�j�P5ȿ���餿j�)�Z�C��I����z���%DДk˕I�yɈ?�������r���ǋ,Q� jE���h���G�N&��d��a��I�.�	��f�oG����Id����IH�9�ni��?��QBX���	��/�d:�,:: U��b��(	M�ٯnݡa
�V�����u�[�����֜}�e��7�=��04׽(��'\F�W�1G~t����V��e�k即N�R�R����	��u�8&��H�?�*�ȧ��`1�o�"�j]�u�ZG���!3V��FaĮPz0PL`X�'�Zu̕m"H����i*}�{[,-��a,���s�}Q�hiu��y��w`��6�{�:+t�u�ȫ w�m�l�p�ރ����z�}r��-�M�xd��z�%�c��#y �,����D���!:s�,y�)�$ �K����l�/g�ؔjT�lL��]��n� �x�Ծi���i��*�m���W��1V�Z�S��;d`���=��/����4 (��r��h���[K�yV<�_h6	��F��6s�ád�'��>���Uc �}G���C�?�W��A Htd�JnwiZ��b8+�Q���/ӗ䤏��a(!ѐ~3M�.��f5�cR�PwfQ�����E�gU��~ ��<gP�rB�|�Zp���k�(w5��袗�p�s��`+D�ݣ�#�3�b�_����.{�~�6����U���ٺ���ɽ��-U$�T9�h2p�(��Lf���k�Ӓ1�&7s�_�:�v&���w�Xjn�QJs�Zo;A2$�H.�3������g3��g��؅[�܁�ؐ�".f�16E�{�ejD^�7�����M�}E&v���a�)!���z���9�Y0�k�V�S${�6	Ifž�s�3()p�
��n�:n9�G����Y-`!Xv#H��}o'�%�tƭ��o8��kf���<�3����QY�r��p��J�%D����	)�V��t�G8\��,8M<)���W�U�����S*��􋅝@���kKWr�נ��%�Ս�d%����5'H��͢d�$v��H'�ہi���`F�G�M+�d�`
�0c47XJ<l�1P��Rg&�[�Y�����x���m߂����`���p������;�kY�ll��u&�����T�>L:{����_)΁�0j��(��۫Gƞ���x3A�R�A�^'��c �fF^`�޲��^%#Hv
�Z�"�U�i	����C2��2
t�NC�fV	��l?;�am孜���h��n'=�����C�[��p1{�B���H(�����&ܾ��*�T�X�L�d�6*�I%W�� �� J���#I����RZ�C�#z��w�k�����A6~q?�τ��h�͏����T��I^�"&h��H�u7��=�1���#Yu�ݣ�9/==�I?�9E� �s G��_ՁS{���kR��O��xmY��_ ��Tj���a����p��v�"hs�+1�YݞwB��'9X[�߽�}�7�� ��Yh���s��x�E3����>� 4#xH�')|pJ��#��-��p9�{�R6I�lN������j�[ aʽ�0�$�`%栕��� ����U�p�uū�IX
�^z����(��4*���;B��5�~�Z��V����q(�v{48Mu��?�O����d�ƅ3嗲�Տ���e/�ů*��.O�����4Ę�ƪ�T$�I��.r^�҃�N1���������ýe�:o�(��B1��r��*�V���*>���M�4�v�˫B�~,m���]�����l��[;�D�쪣Iʎ�G^=��R׵4iE�| 1���Ҁ�gFs5�u��b�y#�ּ�C 嗫wº|CƄ]S��3n'X8�v��.b� �i"�	4{"O�p�I�*����T����d_U�u<j��Ӡ(�n�lT;x��E�/G1��l�9E3l��������h�'�Q�V8�7���-�bB���):���(�?�s�q�Ơi�Y7"��]�A��X��B��p _�sL>H=�k��a��ɷ8�CȬ�5�R��2��0*j48)��l[!0��!�.�2��C/*
�1uA��Z�+����G�s����H���݀���8jkaD�p�������PT���z?$��m�W�y�����z��L���[�کA�y����=Mީ�v�U�������1y��dJ�w��]!�����-�^��Q�Vh÷�B56>�h��*�JI��T}�G]����d��{^���� l/"��}�^"4���\P�3�PV�9)+ฬ墤Ҫ�8��s��]�H�����!�5�ess6�z�	W�ɪ���^����oȬ���4�ƨ��K��C�A5/�"�eEa��h��u/�X����M:�g�J唶D*τ��Y�<��Afmʑc�KS?>�w�dĘ�R�_���G4�n�%g^\P�N�X�F��S�MZ?���w�B�Q<��#�������������!&��%��f&�K��m��B�>Z8�E׼K+C����@VW(���k{���x!�x��P@���~���S�:vƞR7^�����+W�tH'Y�]�>3=�~{�7}$���Av��䀭��z��:Y�G0z��Z+���'2�>�/�|��9(�`\�����N�$L��Ƥ��|}"8���B�j��<6� ��d�,�r�Kd�.���W��t�$'�VE��:�׼�D��V�/�m�6�\������|�d�l�����q�vķ^m� �[��v9���A���G���
��y��Ys���5�[�Ԩ�Cr�x���T��j~V�7���6����*�O�y��Hɭ�F�������;��:g~� �ǷvW6%��?�hl�p�Łw̏�PY�9Vm/�6���lD���H�[����UwS��ZY��W�#5��%ن3�S(�Ɲ�eX�fD.�Y���6ٯ�;��M�	]!�|	}�!9�B�`!����"7�[�O�g ��NN2U�Y􆥺4�+ʗ��w��y[(�F�h��Vv����jжܡ�.��ub��nA�j�a�F�Ŧ�}y65^QD�_t87zk�O��v���i�mV�����rM)$n�����O8�˰�� ٤��N���[������U��s��Z���M�q�fܞx���'\��-8ދ��	@}!V����=��ˤ��:�Ft�S��?�j���8D�DQUV7�B5���|�E?Uȏ&��ZR���)KeKƝ"t��ak���[�@�aik��`����`3y��:5�J�
��A �H���V��u��g�<��v?�M�g��d�'N�.+Xk�g���x׊hId���j�1U�I�x[���2�+kX�բ2��ͬ�x��O;���!Fo���h����{O��/�K�cF=������P^��AG�W$A��`J�9����"��!�v��%�� 82��__��|�cj6H������H�TcX��|+�������-U�}G�w/�^��~�G6`�4W����ML䦗\v�j�	|t�C|�X��`5#\�=,�N]ɇ�,�6�{���f�`w��| -r�H�Z jV��x��Ψ~�#K���"W]�]������ų ��I.��G� �U����\�+�����0���8;�����"|����Q�:1��(�[@A;{RtN=��6��I��t�N�-π�_̝�h�u�/�D��kR���(�ji�6m���f�C�F����U�O�E��?R7,��Z�r��]#ѥʢ/���^哨^}�K!�9夜��Z�,�(y���n�總6��z����dzd8�-�W�+>qr��CY!T(��^��,��5�����,�Fv�d�-=εk����h�����D����O�B�����P$-��/Lne�4�U����p6=��@�
�k���e��O����g�߸fr��(_m?F�{��\k����qwxٛh}�(�:�N�a������^ז������\���t��d���nL�f"�"��Dj�vhd�CZ����`V=�;�����R-V�#	��Pe��՚� ��=�qap,�${�pǉk��V.�!����w������1V��U�=�^D��Pl��R���0�	�.�k���~Z0�t���#|s�b�o�{e��E�V��9U y1�3M�~�
�V�%V�k����(R2�*����#��79�Y�y��צ��"�z|{3S-_r��A��r���_���Z"�m1;�����uܖ���y$�.{��M��y�`BȪ]��]t��J����%�I7���I���@��=j�u�Ȑ^- |�t����M]7�P\1K��K����m(7QXN�|�>��y#��Z?C��V	p�xmD�����ب��$�;A$`��jH�H�#)����8W��yt_NN��cPd�˕$�3,K��*fK*Wx���m���HW'0�6��ɫ�!a/�v�`�E�|��2M{`�}���)Gp��|��xv`u�ԧ�*�J>G�	,��5m�@�U���#E	�7��M��r�ycK��n�|�
�/�E1�;�Y
�^$����-��������Uhr�����I�
�E�e�����)��(�ᓀ��(`�^e_��B�_�v�\��G �e	�]?%*�8�X'@�zg"���e�^ ��&4T�����.����nKJ\�2�J%�D�lEo]��p�i�*��b�!-/ꈏ^Bµ�����}���R�C���5�DF�I��)dvԿ���rʁ����G�U��9���cۡ��y��'�F;�t�px
����9����>�y��c��2�1����uh��gUa�D����k����s�~ZC�V�ۀ��?2c��}���ݿ��΀�ٹƘ�+�����(�g1FXu'Jj͛[���EHeFy�G��]��|{J���x�J5�%ָy��s<��Y*��pLq�'�a=~qI�8�ʁe���R0 �14\��h���]G�	���Ǜ�M�B��A$&]�(���bw��@���`"�����5���cI��ˀ|(؁�Ll5'�	�O`��XB0����pH!1T��"d�`�NI�n�/�
�E�X8��|����زFkO��EE*>�AnI���mK��x��e��mÌP����-��g|�
�����^U��B����p/H�0���-�ﺡ�sݶ��ҵ��$6_�I�=�^�~!��5ְ%��Ҵ�#�z�����:|^x����f�Y}���gXy�V���h�AF��c���зiY�;��n��I���>���lǧ֢]�ʝ�V8�H/��X���E��TF\�<�]�4������Ձ�*�W��*t�u!�_몔���x/d�%'h=�s?���;�=Wϔ�:��4Wl ����h��]g#�;����㰍��=	��k�`j6Do��.�+�61�f�j[�b�n=�Ay��{G�R����VE���u�F{a��k�U}t^�n��6g�-�c�l�����N���\��ۀa��Esi<{-�l�t�Γ�NL��dMtn�Y�ػ����"��?*��7��W������~�[���"�~n���=�,������]Ԇ�"K���z���)_-�5^���7�]�-b��r�V�5���Y�1\��w�Vf!�C&t.,c/�1������c���8w���E�u���y�Z$&m�o��Yz@~��<""��x�p����Sap����F��v�`ݡ�g�f�f�`M�}�Mm�'�QB�ܒ�s���ZXl:���4�J�V��y�Ps"ć���efUa��*��x�/�!�ߍ��6�����x#��Q���g�3�0�w(��� ������� 	N2�#p�=��ߡq�59j�S���<���}OEf���$2�����,�fyHO�t�Z�<{v�!���F8\�ʮ���R���_$�*�Mw>��uV�����qE.�_���n�0aRK[.��v�����HxJ���D�'��q�q��ҕ� )y��K��YE�Q x�o�)�����~a�Jop���	{�RVL��;����8�����.��u,U�w�Nl��_�\�$�ᵡ���u��t\17�3���o���|E����#�Ն
}Y��������*�4�܈D��Z�r�9��T�����&����m�]V��F{;5��L��ĤGv�l�1wq����j��̠3yD��F�l`���ɤ e�>9��-���߽�a
�ܝ���t~kC���XJ,Q0W7Ӂ%�����XW~4�Cl;�t�j60{:ˆ�2۳�9TI5zgT�=ZVj��\�2,L������{��na�9�M��~�|?V�O�T{�`�sw�B�l�x)���#ޘ<���U$[Y{������P�_[�[`xM��
�u�^����8�0�Y��m��Q�K�����MDZ�t/�%;�g^ ��%�[���"ӕ������!;]ԕ%�0k��n�( ��$�*�5��A�G:���]g��������Q�������y�`M_��ף'����	�R�g�Kߟ���)�P�U��ڎ�sMp�C[FU4%P��X�p׆L����OJa��|%SՋ�{��?���=}��qo ��⯂[t��iatջ�Ň���ғ����!���;��oK�@:�w��|�"I�b�{���A�~��+��?>��&��s�~z�{� �Q^��|�8���t��)E7�g$�`��Q��ɠ�O&�Al�N�i#���B���#�\<��b3����i���6MH'���'��m�1V�a����.(jy3\G��?7�h�	WJ�2~Z�(���#��uv���^U��!�O��B�Ц�oI/����e?u����p����Q�AI�#���7�F��"��=�� k!���$� fxE�Ni��-�j��KEY�$Xu��Sw�b#8��cA�:a��P{2�E��h�9�=��]�}ܫ]�La�đ�o�E�(��� ?��#n((ܜ~4xp��&�$�Q�%�o�z�e��5�G�*s���<��T��v������2nO�68�'��a�.� ����/<M��;�#��{�2t͉0���V�r��Q���W�K|���}��@u�J t