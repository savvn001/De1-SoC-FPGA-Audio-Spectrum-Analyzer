��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��YlU8�U-d����	�Ug�}�6՝��{�f�C�%����p�kE����\��b�Ad�t_�r��KM�X��cZ����i�-=���]�����������
�h_P�I�e���钠��4���d��{��u20�l!O��Jw�����gV�e�F�[+|t��Z����aa*�rk~��;�:�M[�6��T,~��N���zm":oϝB�l�����Ŕ��1��0y��RΚP�pə o�<�D2_�*N^�t���D�j�O��cG�H8IZ�R_èM�:.�C}EA=M�S����6tvdxך������Z��T��k�k��\�۹��ܞ� !�Z���b�ٳ�����e��H�^�^����9�Ӷb�?���\�ح��h^�u��֏���v%Ș���rP~�_�_���d%sxre4��s8[�^��~vb�cĕ��7�L����c��s��G��k��/�ZxG�pF3e�{�@��b��RQv8e�ӷ��<]�I0��~*���	��d�I������<k��YmH�m+AE�����ے�	S�_4>:�2U��R&G�um��_d�	-�b�J��Y&
�xMo>��(��e%��%���Y����QNfX��I�ڷ>�H������^�\��e��Ы��Œٳz<g�s����H(ӄ��,�\*��<7Ul���m_�J٣b�d��G8�i��K�R-E�p�@q��8�V�s�*��2�����M�2�M$'��x7�.Y�~M�IL�N���$P����|S�d���B�c�.�#D�<� W�����`��`�z[+*-B�[�*��b�H΁ګ�-���KC^q��;q!ӥ1Z�\l��N�0h�.Zt�_n=ۮk- Z�!���&�0��d�ӱ�r�x�LEZ�mχ�'D�lYKx��7���CaHwZ����78�u��ؓ�\�!��<�Cp�L���t����Aʔ����;�n���;�iz%�s���)�cI/tp��߾in}hwie!� ��1���F�K��w�z�0ա�H6��$N�B�Pş�30v�E'���AD��n�i���r�����:8�R�[��F�Ƃ[�AV���S\��u�z�A��;�-��lb�J��׫GQ��gQ܈��,�'lT���*[��Y�Ş�ރ��>��&�s����K}9�/�D������Sa2����
�Z0EatxF�jX0��t�C@�bߣ�|7�GH'�����PGP�g�����Hئ����X�K`+N!a����_�E3������ �@W����a�6r�qQ��� ځ���]C�
֑�>��-<���w��K�x�X�+�f���t�1B �U�p�ѷ�E���V�B�PV���7����B��q6�3`+� �А��'u?p6w���u<�5���DC�/k�gZ�B���b�s�|��j7/c�RJ�d]���,N5��%��Im�O��#��ֳ�V���]O�8%C[��?��x]O�v��,v[��c�R9��n�3݄�\4|Z&׀��)�^8˕G�3M$Վj�Z�H8)��Pp�����v���͜�R��W�qx�3��qohl["��N����Ƚ��͐���F�Ջ�u�ʁ���Uo��	u��_����S�<�����e����d�٣3�p��0t�5!GK�N�b����z�1��jԧ�S�@"5�s2����n�d0be���Fd�}u2�˖I$2@�9���*<�<��ېyZ]��N)�$,z�a���ʉNc�#���Ì���j(a#N8��]��A�U]�ϯ�Nak� .&�ppa����N�!`$ww9�f)Xf�ݑ�\OW܉@	OI��nA[cG�(�<,��n��F&8�DR�S#�"��A���U 2[�����X@�qI�� 2\��2�54Ww��x~P�ݢ��Ҭ֕�H5�
���7�S�Wjp�؉��|,����Ѭ�?�c���|j>T��F�5����M�J�w0C�g���C�`~�j&�/�H�����I��k<r��KIbT�G�]�O�E�g��U�+oٿ�����x�Z�RnW;G"����n���⬴1�*�7�e�@,��L����N$/G�yrg�5|��鷰YgLt~{��s�2z���-UH@8�)��1,|\S�񹻣T��J?6�����6����R?�l��>�1Y�=lx
X��� ���Ԙ�����{��uJRZ���ō�0ۧ�I��`eL����������W��Fg���HD����P���7�/�#�`��ܸZu�'lA��>�y�Êy���'����mg��/*�n?�1l=5rqq�n���豆&k�Uq�̬�@{��NO�b�0�d�wh-�d6�}k���޿k�A�π�p�B9�����n��?���9���)gU�]�����-�?�.�Te��Y�=�X�`�m��Z�K���$��gu��4'������3[^�|�e��b�0��a�HߩFq�Z���P:
��'R�x����f0�Yn�ƂZ�Hz��>cf.y�7���9�����|f.bӂݝ&ɨB�dk��ݎ�����U-o{Y�Cu�����*t�e���(�`ҝ�PY�ڑ�p*���❊�� ����6L[D�aCa�-&w�ꡤ7��,	�'�[x"��
B}]M=6B��ے���7ԗ����j��-���%޴>���l��P�Y5�61,����Z�:Y�J@�R*j����H���q�6a[�-%�$��W�M�^,9�d�-��[}T�;��tU^9� �o��,E��6t�K\j����T=�����}׊�T!R��蹖��Y����,}���K��y+��e��Wra/�����2�`���&��E%���bg>4�����7BE<�q�k�2&҇"�M�F��
�����R���i1Hږc;Z3XJ�D�5^ 0�FH3ܑ�2�mz��\	c��^�dh�O����U$�zn�0U�ϸ��Y�kn����Aݳ$�E�U/���Bto�Da;�
F�nԦ���2iFK�Z�JF�p���C�3�n��(f�* ʉ�ʾ�7I��r�R�E���{f����L�nn�N��2�H(�*���&T|v����*H�E#v&|=��q�݅�O�zy�4+F<�5�{jG�{�����T)�
�JBo�;P�%�Ń�5)�A�����wG)fPn����ݮ� ���Q�k���RJ�N�JH���|�O�W����!U�]W"�] X�`0dKu���}\�,ߖƷ�>��d�� T(�ܺ�F��tBZ���bR^Q�	L�g�)H�#ӭ���?b�e�Z����04��"�� Ա�7���� p`cFt�f�	�&yAՅdw'�Y;�!6��:����C֨�8��j�L�M�.x0	�
��V�(85������W�L�sl�C�o��ڀ�7!n��z�o��lc����=ٺ����qa�L8�# S��P��c�/i���$��%W>�K�8����
)���?F#{_�?!�|���?�s�����\6�b����sXG�_K���Ԗ�S��(�>��G,�( D��$��v�J��l<.\8]��@@0/�|���U�|%��)�S6w�yͩkis/�'���p/�� �B?ο��� e[9�G�;l�b0i��+u�ig��!��_�Z��b6��6^A�Ȫpw �\��\����{]+A[U:H�Z?��.�������v���a�`��-e@tͲ@ү�t��#f;�A�����K��+���8i;�.17W���=��_��U_uGSd��K�K�P�P��-����Gal���I�z�o���P��g�Y�I����uU��M���]��A:,{�G�va���� ��)�J�w������Ί �����ɚ�%�q��A'[pnG�6V)�U��{( ������$��9c'|L��[ *����lz@�����$�C�k�����:�[�!~b/e����\������	���`��׋��H��Q�o���Q���D��H��`�_���lg�<S'7��(��&[��C���c�|:���C���� ����� P�@�eַ|��mġ󼖿�6��z�S���|<���9� �|�s�����<|e��K�l\#�7#7�� �E��]�#eV'�;�m������%h�f�"U'��0ˍPk�nS/� י���^�C	V&���Dŧ�T�qkn����w`�B�ŏ��}k������|��1���}�0��B�
���Cڙ���RR�chX��sԎÝ���EW�_�R���A*e�X�W��m�L��xL�#�C!5�_(Ʉ��~3��u���cw���Ao3��%W[�@��<%MVe��Ҩr,�k��C\ ������1����� 0�.�k2l0!T
�QaY�}	 �Ѱ#����B�H��a�����	ӦV�2GY�bc�6^�lӓX9�:����HcLqْ���f��][/m��o�-�ϗo�&E ��Y�yR8Z���kKpd�����Z���G��L1����	J|�Ψ2;���R��'#�A�D�#��4�_���'j��8t\|�k��0�]�N�@��eϋ(5��d�8�G���kE�~3���/}յ�F�N�����K�h�����au�����3�U`�:���7�-����{���-`oK�V��Q�gOXp���*dҗ���x����_�%���v��ys��ə�aܛf��ěZ�SU$m�b9���L�3?�u:բ���i�Mhd=�[#:��Mg���*��S���iE�/�L�%�aT����W����x��&<n֕f�~`+���pX�Y�<M�Jf�Z�T�����In^�(�&#yq5֓��f�	%����2�o'>;��ì����8��a�3T���3t���O)b�h�rQ�����I�x5]@���ҏp*Vn��K�b����I>�TzI�'ʎ�G/��1��Լ�����X�R�RPp
��:�}��:<�z�}-�!��^�{-���u?���H�6'n'�f�
�&�a�d(���]a/� r���d�F#g��͹Ӕ"�ϐ���'��_��J<?ꔜH��
�i�7��Z��jWSS�xo��>U�\��@Q(ouI��l����y��,@�h!�Q9�Qie�a � �L���CG��q~ִ#;Х�N���!]�i?�� !�+	h���qE4�Bz�H���q\�?P#\�����_nǶa;~�)��b@�����<��~����d�T�ΰ��<��I>��Q�ߘ�9)h��3��*��x�gO����X
C���
�6�i��w2�6�U&��ك�c�Ob�VI*]�Zi}y@Z���JQ�i)1\%���q�p�H� ya�u�F*�?)�I�I]��y����	����c5�kw��?��^����Q+t'�ȴ�y��HM9��dU��+��C�Eu�v�mf��*�3�|?x�����N�PI+�U]��?�0�����1\���ZL���u$��N�U؉w�?�� 	��a��� ��7�z��S�>�/j��~5���/�d/�*�#s�}\���k�iw�J�= �Į�E~CĦrg��-$
��Y��Zv�r$[)�ޘ�B���\�<J%�TsU��E٬4FO�鱶J�����4T^	F�Eh�A-��H$�ć�-n�����x�ٮ@5-���'_FɆc_u�����S �;}�Ĥ�a�.݀�M�.���s]����)<�D�Z�t� �7�]Y/�A�i��d��#TH�Mr�y����D�j?P �X�ӓ�D1�q%���O�T�Og�0C�q��\)o/2zة�������ݶ�/�r���p�y+fO}�g�4����I"��1�)�N=ՖT�����'7
��4�|AbR���,� �G��tU�R��ɬ�_�9��d�us5���M%���c5�=�b+��Rj.#i�e����J�+Ǳ0|C�c���6b��pT%������7},�or�?�o"yn6p��}�q�q��Ԃ y�5��v9�>�}�߭��h��P˓����n��I' ��h��9��Tf.�JV��ߺ(�YD�� �-���� ��P��f�]F�s��逆���c8n �������rO޴�s�U#}+�!o?�ƛ����u��?}qm�q#�40;l2���MFN�Q�m[��ا���~����������)yAi5ϜM;� /����w�2bw�i�1�A^�
�I�2Xw�p�*�����HV�_ۢ�\���oU*�X��q���z?v ��D�����D��B��o�7dw�yf�'1�I�\<���}���d5Y�>��ӯp��D-���2}�q\�}�(/��m�B	�*t։�G׸�e��hͿ����w�w�d��<$��,�e�"��(:�.
p�\�8&�)��{|�t?�.�r�L1�Z�Էդ��Q1d��+���i@2�4Φ���>��H{�?M�E���^��ou��H�l�}�N3Ѣ3���S}���[����z�^1��'g������<�n���WY�Z;�BB��p�o.����u� uď9&;6	
"�z%�j�z�����p⧒|�Gڵ�#ubG�9A���ϻo ��3�q^2h'Z
ߵ�]�f#`�&�y�ö��^(���$����eL Q���I�M���gҩ�H��[o����$xJ>^�N�Ť;����aZ�F5pji���'�P��u��,����^��D��(���;H_I(�X?��	���;����v����`�Cy����Kb���X1��������[m>��x^$4����'[�o���K�y��=%7��<���]@1S��'�FϚh;�FQx�z��8g���y�&L��0������{<e�+ S�e@���X5��}}��J��q�(Y_˜���ΰ64�_��~@��qXOgNmv����d�X�e�Z����b�B��w28���t�X���/J�/<�y��}�O��W�:)d���^Qb���G�_��BR�ڗ�� 4�7���7����htv�Su��\�W���\��#�"K$��)����(�+Z{��n��9�1Q��fO�zO�
����d�ՙ�\�:n�%�%gG�8��s���Ŕ�Z�5��}>5��0��{|���+��� zeh�^�>�S~��!M)t���$��,L7�T`���s�zhF�EnU���9��Ö5�m�(Xȁ���l���c�kP��b����p+mkR	��M�h�M�����#�a��x0Ex�A�B���N>Wi5�&vQ$p��<��sfb�
q9��D=M�D�!8��ٌgpL�zh�jL�"�<�K�0��Ғ��]uS%}�Gx��?�S��Q�O8_)RG��9��3e8��h������?V���k�g+t=�|��k�E�U�TF�4�i�]X��R"����H�W��l��+"�pX1/��� ���j�����Q�1 g����Ղǫ����qS�^Ir]�����>�Y���V��X�~�=seH�Lj��@g��>�H���­-Q�Y��#���a߻����h��3D�k�H�� ��=�*p�1�����܏i]Fa4�<��J{o@�W��:��w�d��l�,�i%��4r�2LЗLj�ܦ7q!��E�d����� �[*B5�M&�?Ј��R�*{?#I���}�xm�쉽�I�m�8O`�%2K.fȳu%�˙�~_׏��;�^O
�I(�mm
bzS�/j�L�Gc;���t6�_��5l5D���?s�hmc��T�vgw�գoޅ�Z�|*n����Fa��X�ݿ���mgt�҂v�y��Jܬ���J��]'wKYQ��_�̬zv��ڣ�D������P�W1�v����:��eM��e��/��!�oA�� b��������q~�^�����SY�_�0{����A�؉�Dy��_�Cܔ�c2EF���3�ii�{���7�>u#��YsKK*�R"q~��y��^��,=/$���g6`6�o�����t���9�ydM-�+U��ys��[
�#khHn��c�t�mE�^,=t �Ÿ�}@��C�W�� ��!�'�_��o�y�^"�V�^����嚛)b�3��Ss�`�)�~�%�-�Hb?_�j�*C��c5�I%=�Ԙӱ������a%I˓[x��~=P��B:�y�4O��1�,V�}���
w�ĩ���-��q�"��gμ����}mq��N���uxnIJ>���`��e������`+$R���Ɗ7h�:7Lj9B��|���#S+���#PB���&Oܟ��W��|�Rā�
Q�P��p�D�Ir�mŦ��9��*�6�@�M��Z8���g�m=ͼݎ\kf�L�ŝ,nQ�u�9�8����[�P�h��  ��/��
zmeN����V�)l���-f�J�OQ9-�^��&�o��r��k�����hl���NZ�;�=`�����y�$��Z
��[36Ĵ��Ӄ��B���w������Խ�|�Ę�}v���p�F_��~-�kѨ5!;3�ҢmQTpَ������a�E��*r��E�la���Ͽ��|{�>6�̇@,�"���78Re~�+���!�PH �?�{μ����u���v/�[[���S��Qδ�z�@��B�

�M��2�����1�2��$8�����$��@Te��s�����]�6A����~�����]#xr+��!����z�7�\�+u���R�YR�<˺�u֔��OшԄ%9'�8g˿�[�eRvk�p8����Ps�"���{�-e4�/�41_�aI�]ǿ�)��5 H�̩Mt���0���04X8���g���E�<�N�Zh�UL�:�,�`����゛���pȌK�oFJ�>rjA`0���ֵ����P��\
c�F�4���84�O�.y����=�-� �ƅ�Gi�����u���`�м�,`�n��J$H����-]�w�15�~k0�sL�h5��O��r%�0d�����4�S2�3�����p]��y*p���OC�}�w�+�������~��|~�۾ò�����,݊8���5$���q�0��d+B���������T_z%=�U�ߘ��`�1��X�yl�됎��3���=n�p}�U���M$�k�Z<�ஸ�`� �\j�T��K�o�3\7v/�a)��EB�e��]|�ĳ_B1�*_�R����'QFr��̒��?��Ӆ����ұ�������b��v�Qwѯ�"�p�	e���E=%���zgy��q�0a	��&����i&g�Vg9+T��Nn1�-�t���o*�H���T3%*Ln��2q��B����{�-��/s�HH��7fôd��̣��V��@Ӝ������u֬�+�4��k�ڄ[1F�jvK
���G�#�p�X0�t��H%�"jq��*���Q�y�'�Ig�� �k��v����"%l�G=�%c�A:�ߛ\�ǡ����6~�`,K�O�Q2���2��%~����^�����dg:.T��h�UfLggHc����o��E\ƃ;���		��=�:���@D,���i����@J@��c(e���cM3{�5�|��s%�%���ǡ�m"5#��2Y�}�(e���xE��|F��*�QE�����^=Gb�s���E�cHiy�O���y�!�8$��Pk�W�U�cN�̲�Sh4�uB
}4Je��U��3j�9ϼ�7c �5,���y��>�q�D�Y]��aF�-+N�n����,F jEW1�x�IPu����b�U��(�C
���
�V�V�SÝ���-�hy�T�>�/�$����g2�SE)���|���^�����������sMB�?�Q>��u�M225��.�u��u,��È�l�"������G��ݲ�[U�����Tެ��w ��� �;oW�{y;�y�"3U�-X�v&��E� �X�ݜ������=��l,���	g�E�V60qN 5��� O�9�=�Ew�/g��o�
?�����M��?̙{��g�g���}���y��z�h6���9�3I&��E�Y��M��/7�
e�>�:��k�ݘ;A?��y��'�u0Ja��A8�u���5�Kw�!�Xi�V����;��aЩڋbA�N��7V��M���`3�>��2���i��R�,/�p
��D��C�o���R����D��n���me��V����ћ�
�Yd�4�c.\�4�ɪ�^.b�`@�/�����T��ЬI�D3DxD� G�-�����]=��$����b�U��]�Um:�O6?J��rS+����ј�-��lh�\]_3�?��+�-!r�ᨏ����T7M��T�i���UO�ʮ��ݝP���>��da-��u���g�V��|�<]X�9�#��V�0~�����)4�
|-m~#<�X?�l੐��Z��,EM<���m����Pd?'؏N�,uf$�,|���{��6�/�~3�.e�(�A
�Tg��*�u�������:�K��WK��͕��?�u����67�̥�vlN�6+�[�������h|\��&�Z��k�=���5j�m�� �x�Rv-�[�9X�ɣrP&?ߍ(���Ih�{�fGͫ�uJ�JQIdb�Mi�s�MkB�Ч�v_�V�=����E����Pχ�jL���MB��z�K�wUx��R�XT��c�k�
�<�l|��G*��e���`,)��t�f��g$I�Sn�\�(���nO=f��M����dQ�L�"eԒž�1�JT�Q����Y�r�ԫ:������+ע4_��^Ϻ� ��qJ��Ṛ�E���v��8��H����X+����R"B,�$΁K� ��V,5�r�w�+u�1n,^�C��L�˜#J��̖̏N�~��"��f}W.�e��~Z\��n���4�ζ�����d�Qw���|����7�Ϥ��拙n�W����J褿��#brm�5-�$#�V��',��B.�F]����M-��:�L���Ϫ�p@ff��Qy�"��{Z�+F�&����f�ы�&���"D����F��&O�j3*�i='�ހ����)�XJǰ�ZrzWł���ҕX̂ff}ij��X����?\��Q#�Ss����/�a�+Kﺂ��ё��Fbʭ�m�jt3|h��(�m�XO%	�	Y9���"���"�`_���*#�\qgA�A8'$i.ٳN��{6��O�J�<`���[���U�į�N��aS��>�]�#m(ŚԵ��Ot�����eW5|�,nӅ�L������~k\0ݘk�Qe�����z{�Z�-�}�%��2I�I=ێu_&�c��dȸ=��S��B� �U�~�0��p,�i'�N��[��@��|w�p�,��� :��������"�X�h�iC���S����w�)���9<��z�Vy��B��ӌ�"=���v�	��3���_Q)��rd�k��X�����J���x'��b��7(�Ka�Ɍ����=�,.�΅^]�-os�=�lf��� ��[�����]�t���l���%O�!�U�����Z������\���ٗf&7���"����gy!��B�%:��)\Mj2�w��.�+�sRwT�⼝\D�H�����TfZ�34���U��_>z���P9+(;q*f����M�a���#�`��3Z,����X;�m��ȣ�٤S�4�ٜ&[*n�*�4z)׏��$䠡�%U�u�%˽&�2��/���T���*��6C#B2v3^��4�CK�%�g�YH٘'0�Nc��EI=C�,��llK"zE��5p$��s�CK��4'� ��Vk�[90�t֟��E�ޛ��{�����?��0���K6<�������ݟ�ؙ�ۯ33�XM/�˨���Il��i�S���i������r�S�J�Z��ZF��cSM��$C�R�����j.���m�L����Ug��3�=�����~�}8���"T0�;Pش�' d�k�k�a���2�v�"�;\u%x}k$��;a�������b�+:���#��^S��,W�RJY�!čJ�'H�w���@t"�
�U�C�Ax��T~�����mn�xy��y�յ��i�Q,�|vʪLp3j&���*����$��ؠ�G��qn{��{���)���S}�Y�����a�+��h��^jr�O ^���ɱ�-HpIs�8B���&J��\�p\�B(&�6Z2�Uк�)>��c�����NK��Mٽ'���˹b� G`F�;%` ]�����ػ^�E͝Ǵ���7a�pY�܋�M6uL/�<�֛�^���f\A��Oc
tdq?|�"eaR�i�lU�`�9lcfst�# IQx��'�� ��k�c/�ajν~��9T�����)aM[_3Y;`fÈ��`o�Hz��߹���׻��|�F@i*L�j��S�~�>��.���C�4��<Ց��] �+��Q��s4���{`���)���c�(�ꬳUO��Q��[�.5�*���~���5krDQ�7i�5�T_%= $�'����n�=i��tcw#a���['� [v��"\y穀h��D�V
��/��w,+�,ҧ��|�d�K��>�SR�W�������Yj%�����\��8�
gQ��U p����������U�g@�����R��$9C�YW_=|G[�$�^��[���$�<�;����XX6q9�+�1��f/g�2��(�d6���
�8C�͇t;��"~���D����ZP��[�f
?�o)ʌ�bW��m9�2��{p�ٞ)�_� Hcz�G���׌���=a�z*�x�F,jf�n��f�F*��l�hd�!�o���M#F%��$cMAct7o0�X���`��j1Pq��3b�W�uNS�v�:��1��H���eگ��ˡ~�NuQ�!ܽ�����g�7��Z�V���|�Er=���*no�uļfnU��@��/[�$�.���CL$?{�B�:�z�=n_��d��^[�K��å���C�x �<���&h	�0�d��GΉټ�GkB�E{�~���D�8�J +��څoQk�.��x`�������Y���g�1�I<��7�q����5�PH�����^=�M'#�k3�O�Pv�LӝlL�����\Mh�L�Ú_����Ԕ�/ӕ"M�o`N�	i�T	��kR��7�*�fDx3���@cn�f��{,�o-��&��x���*\�8�z+h�f� ���EI�M��b"B\d��(k-E�8Nk{��vk6P,y�0=��`�0����e$�)�����zr��q-p�0
H��><����g�׾W��` _��oi���rlc}�q��U���?�����&��\��Ń7-M�2LW],�<v���6<��G,_�����rV��,Z��I̙�ʻ)&�gZِ�7���f}�|���$�k��򄽐Џ�?G7���a	?3(?�M��a��,�#^�k�{'ص�Ҽ�ؖ'_v�S�1�(1s�O��ef���܃��	rh���Ӏ�m�:Ts�)����!��C
	 �xh؏[�-B~sh�ꉆ8�N��"�g��PT�B�c8,��b�10�w�T��I����~�����>��ƐjW�,_ц��C�f�5��e�E�9�#����O�������3�q\����dU�yG�tu��,�M���z�`�]@(`d(J���+I���"jIf�F�P����Nئ����F��h���V<l%Ilsݍ]���/�1�Y/˱b�E,���!���YO �؋���E�Г����
Gi��MM���Y���۞�zu�⋷ە������l�M��\^��P�ɡ5a�V�D����V!������p��i��SG|"�< F��6��"N�r��̊s���Fʆڻ%LT�q��n�ݞ[*S6*����$b�J����b�j�+vXkY(�Kp�P�H�޺cv��ݜ�+�����Dp�{����z��K�U����?A[^�_����D��0���/�8�6�7���X�����1=yNG~Nę��\�O4)\;� |!,���+R�3��d�",����Gì[�K�m�8h�̃��jS�A���.�a^2.� �
�v���Ç������r���Z[J�&޷���4�u���-���W8jmB�"ڟΧ^��߷+��V�d;��{�vm�1GF[8���zy7�x�GIU0R f��Io���B�����Z�OW�f�3碰{�(��4T2\�����\���"�}�P��ч/��\�����5�����G)� ��R����� �$�ɘ��uER׶�FK��{�=�nx�k�oi.@��@q�AG�.!�V4�6�P$W�K�^�-9w�۟�$���Tl��&�Lj=.�U��Xa%8`��A:�Cc�y�:yl"�v3���WK�P�X������0�>��,Grz�V��'�&B)w��eZ=�bn�ecHb���|�m�����;6��*���R��H�����x,�9�}�Y�lޝ\���K8J����Yy��Ϻ4n�}6{D�[�nT+P�P��?�<)�����~��vX����c0���?'�U��l�
�J��a���,[����0z �dz�.$���x̼	ϰlW:���fK#���������V�럙K�ݷ�7Z$ +d��D�#�n�s��#
4�.��6����vw�pM�U��-C��ՠ�"��5�u���!'��]+�ž�$[`�2���M�?9��莂�P-�!����4��U/C+ �6>���O%O	���H4ߊ�Ȋ�AC��W�i���E_�@Vy��؆[�����$�ƃ��:Z�ۀO#���H^.$'*������"��n4�D�!+���ƌM����:;�q'@.$;t�N�$���e3ƺV{u���K�����/����ץ�R�zh7��讋�w�8?9[����{������b���YZ:��]���@�������ٲC.A=�2.�7Wx���k�.-)���(�B�u�:�@TG��A��̎��*����[�Y?9B�d�ob�qD�ZDa5�n+�	�ݶ�g�]�w�>it#�T����cڑ�#��oN�T��[a���<hX���i�Z���m@q�L�G��D�DIi�u�[J�Lc��Y_���\^�#)J-�+��?]Z��2�Y*g��?b{����O�J6,�gSA�\�U�٩m��WVx�|����e�am��I�L|����~r(_���O��Ȕ�5��0^���ZH�⯟�}�\1{C�JFnE"=�bDq�M���jȝ�������aEC_��[��hK&��Q�~�S�S: Y���&���l�u(�#N�oU��e����
�А��%�i��AZ!������
��3��sx��;d}�ț��D`�2S+E\ƴ��'29�G�#���]���x�` }f���#VX��a)F��ݼz�zF�<��5��U�f����ء�ڻ�HMЊRU��i��e��[�I�]Ʊ/�^T������̫�Tm���WK@�����zbS��&�stcΝs�]������y�#�j�h�%m?�9��,����ϓ��KF�q���M7��5%	m�	2�ܣ��B���|�V����a��-�T2�]9p�Jy��6�}VB3}�B4-+�x�����'W�~�*a5��f�H��/�mm��m���(�kv��ɤ�@]�+$�#.��a�An���hy�Kf�q�8�?Մ��v#�q���"J{�.�c?�]�D�W71�g@���^�}`��Ћ�]�e���wվ��w�)���Y��d1�0%I�i7O�"=�5
센yK3��^��EM-mh)����|-v��=�^���y�bg�ٯf/3�'���mH6²L�GXEJ-�N�޲�9 �Y�}1A��ʝht��FTh��	�c��C_��ۆt����1���M_ ��S�H�Ι�7�-���o �\s	���7z/(����������<$m�@2�Ή��Bn��p؋k9Ki�U'z��1���` zq!ސ#��vZ�aP����)���Zr�f��W	�|���r�������!�r�0�ng�6�(�w�B`�e橥��4P�OtQQ�K��J��Y7u���!�d�d���Sk���o\�N��,�B^eLH'�#���wD%'	��������$�aq"�A8�gI�������]G3(\E��#Ve�"rUT���cM	KHG����={>��_��d$%�A�F�$��F��^ �������Ϋ!��bC]S�
�|F�{��>��jj/�%^S��_&�]Ō�E��+ �"a4��B��6��8.�o�!3���V`}@S����9�?<8̮3�yz傠q3���LR�q�r���T�̆��Q}s���.d���$������R��j���>|E��}�2&���F��q���ͮ������if�E��,s�wkw���Xq961Ѳ�M�V@'�!���X�ȫ&Z�n��6LF~�A��j��s�~Y��W���Y|�$��5�\��F�3`�1�� bO��jp���h$M��1[�_ ~ ���n��;5����/!�Z@JFnv��ޡ�ߡ?7�Ki�ʣ���O��oG|��v�#(/�`G�ͥ�M��!.�4.L�X�T��kE���=o��T9G�_&�~
�5�Bs�2���[��~��ʿ�!�p�Ab �g~�DC�Z��2��?|i����=�Xp�~�����O�����^�"�����ӣ��p �ݾ�2��V�	=q�`J��Z�T9�"&��(0�	�����#�a�?�(#D�Jx�tY�=�ЧD�f�����x��RMuٸ�$�����m�I]q�G1<t*��$��W �A�p�
� �l(Җz6���3i�oq=���}��I�<�<wAZ����AV��?)$���V����+2�g�m�$ȴ8�����tN!LPڶJ�	���t�`	�Z�!�L�8'���l�x��s��B#�`%Ӫ�j���B;j����(���-�"�p\
 U���y2V�xS��|1A�Z(��"��kc
pCM��@c��8k���]@�ܐ��9�Oj�X�[#r B ځ'��G�6�ւi{���_K���\O\��#I�-)�2���+��\�#��đ�xI��>x�R.���[�?�-��+^��5O}�4�i=9Qo��Ԑ�B=�< �ؑ谒S7�]�������BK�1�Pv50p��o�B�B����
� ���Oʹ_��\WX��
�C����u1�fX$YWm�Wv�OD��),x�F�I�Ge;Ry�q�M�+�0��sc,�Tj� ;��l'E��*o���ke�!�Β�8�����s�O^�z@ק�2P�}fL��F򰹏�u�<���+݋�I�N���eWU���e]��r�54Z���*�?��%�M�"�lP�D��!{//LCQ9�j�s1݀�
�u�N9)h�����L�މ�-�3���8��%x�n�������@IN�5oI�5z���X�lŘ۟hMR���Cawm.my���NN��`���6�	�2�@�We�L�[��W�H�|�k��@��n
P���%�Ɖ�����?"`݇����5�N9��7(�<	~�_�,!'.?<���Ђhx�X�ɐ�Mp�!�"�XW�-)xh0GOrI����e)�;w�#�|z5��!}��؀*������V+kYr�$|��f�s8<�n��I�xdnG�W&2֥�f�ۃ��]�2d<N
ChR�����+A�斲��� n��9�AC����%V�"��D�+x;sS7��5��n��ԓ�s����ݸ��mȵa��\b;�Q�6�E��_�ԁ�ޱy�v�g �J���������y�Ԫ3��w9iy�`���A9��D����� dG���D��p��~w����U���k^����K��\���!�Fc�ǪE�lo�T��{�:F4�~�K��l�{�]6'Sg�ȓp�����3p���j����7X6�>o��!e�n>��c&M4eο��cA5�Q�N�S���^]�|8�S������q�z��	�N��P/�����������?�,�I�e��!=����8�S�^4x��yղ>fBja����h����Ӿa�?f�|�K��H1���<,�$b�0���5�	�|ќE��tOE�	�����K+4��5�A�9Z�V
R�pP��\�k��n�g��2�.΄{u�{�@w;֑��k�l\���]y#��ߟ�t �L.%��2o�4^^1�b"��C�'Ɋ�8N?�)ok#�Dݪ�:���޻���s��&+^���O^���V�fN��a>�� ;����2��]PiP��M���{��HK�s�9�foa�9@ �U��Vu˚���RPz�E���Y��؞>׉�++G9ބ�>����j�7�|[{$*��+l��/��>�"q�˥����U�9��]O��/#��^Z��N;9�t��~�yZ�e��{p��˦��=ٮ8�]�<�:���hU�N�^s�ў`����y�'��HF��FSTB�������@S֏4��]^`5�`��a��\��Qh���@�E
��%�J��0�cەlT�	�Cs��H�������}�C})7'��R%�{����=g����D�>�YG)�n�L�<4��?}��C0,N�c4�v�ߥ���E�����y-��X�!#4�n��&���	P!�|E��l���V��:��KK �|)�r�P["*��o�
�J{5磌*��3��m��揭/rB##+������s�7��ȝ\XڛE�[USLĖY�7�ߎ��V��0S��i#PgZ����o�p����hH- )�-+��QJ{��������KWu�i*K�r�a��3��ɥ�������������D�]�w����6���?���G��y��1[\�i�%�h�2{�݊mt�w�(�p����ϳ$R;E�;|�݄~8�v�7+���	��sap�M� l8�=��-Jby����x�Z�ŜH)��[��m�F��h��]Hs����ks-����S7E��i���nå�nxxI�\���0������6DB�VA����d^+��WB'��DZ�ޮ����!�8��W{p�яK����I�0y֫16
c-#���I~@
� ����7���K��˵C�.�ԩ�?��a)[��i���������m,�X#��T|��'!C�Н[ޖ��I����j���k��~��$�x���fFT��1(L{`�M�&τ�>�$ɮ��<�NN:�̿��+-C�D�m�ީ��ӳ�c�#2'0Rat�:.�Vj�9<p�d
�U��'SyH��rO��(j�u �����g��
��+��W=��lX[������3�p895
a��"� W�M��j�t�9��LRF/Hn��@,������D�-" �U���b3�/7v��]�as�I8��o9MQ1T�����I�p�Ζh�U_���wx�%����$�����(�[u���+6�|1M�GGC���!�B���?�E-���֊����{�ք����_#�N�~T�1+I(Iϰ�X	E���,<��� �U�I� z�?����i(D6�aAq��L����5�2�������V�m9'�����TG�%�W;�8Ar׺q�����~o��7&3�I�SP5���|T+ݛfv�.hD���7��,�J��q��Q-�N�H:�x�l�i<���)Ӹ�����@���'������G�
��ע�Mwn���&x�3d?�8l���6wjm)*ƅ(�R���<����黌���)�9�6�
^�T>#r�'��&�������cy� �\�O("�&�"hϴ.z����
��:[w��Յᭁm-I�*�4�Ҕv&��gҁ~��kqL��m]�,45���nWC !�D0�0ݳA�ڰ�5[v,w�i�}HvB��>R:?��P�8�����C�U��_G�r�z>�0շ�Q�9G�}�@Վt�p���t����S�.h�,�lL6�U6�=�PZ���(6|!�=ߟ�'�����|�����@KwE��IY�����t�{�:�8���-ɿ�ƨތ� Z��~^2�Rw��㽊J`��t���K`�H��Jˁ$9�/�_܋�/��G��O�*����<�f�(�\�y��?�ok�����l�-�!�ϐ-�t��Q�r%�e�-���=��7��ǩr?������zÖ�l���n�@.�2�䋫��Bꟓ��=�o&�� ��|��?��u$��T�H�7��؋��:aS��;55�5�|C�Q�ޡ����ܐ�Z�U�6�H�-�TR`�&@��d����8��7B?Ik|�\�1�`�:-ŚS^f����c��J�J�V���F�6�Fm$vj��ƿ��N�-�FD���|����'b@)�5�9q�>�jˊƎXݱ]DZ�>I���?���:\� �� ~�T66 X �̚jʽq�'s�Q0�v�x#&k�_[��ʎ�N'�H����4X<!�4�V�a�4����׉A�@��x��� �mة%�ȣ'��&��e�y���\]�q$��g�z�i���K :��y}�-���cEf�
�g�y�L!xr��5�v���G�Ӯj��X�x��7?١�������D����ୀ�>��mW�3}����Ja#����II|�[���0��3���4�dBI #?�6��\�"o*��g^��-©���.k5��ʉ>Q۪��&+�0W�LDu�fzξ�����Ռ�Ό�_֝��/�$p��V�,���%�ث4U�]4��@E��K"�=�~/��J�[N�
^Ht�!�[1Q�J�3��$�:x�]�5�um���ݸ���H��?�wb3�R�0'1��� '5�ũ,�
�0��u��x`Ɖ�6х!����ޏ)\7��ʳQ�~��\��>�T ̡r���L��!�_,��u���t�������Gw��h��#�6�b]7�4�Vv
ei�5�y�G�]AU�dX6x�C"5�����k����]@�Ǽ"c
�.4���n���cYg�i�ԫ�����Z��Y�)�)[̈́�XIas�3�WK��m�`j/�n���vnd?��=x.<��&�U��7���#nL� ވZ:z�F�x0n����%#5��̬���oo�H����b���O��]��{��qo�x�Vt7IU��i�z4�-4��].u-RnZJ��ƣI�^A���򯢸O4�3���U���`*�ܽ)<`�z�9^�I뛼��x�,f�[`(pO�P�`v��*�}b�F��W� �����CH���V<�Xc)�^1-���Ǡ�a_�����iʎU�[�>���+Y�i���G����x�Q���ψ�����8�~���l��5��w����B7��t�+G\���-p��х�'@(��ǙԺ0���]�(��λ��qP�{JZ&����~��S�8��Rx��%{c����������m6�������#�㎞���ϫ��s\#_��mx 5��C�u�;h=�d.6\{7[ ��w���e��6{���3N��Q�r��0<�S���=Hߠ&��5/����e�������%����v��V��-�Y1�#Y��QF��,��x&&���X؟��ZF�(i�b��1S�I�𽸫>�Gry�n��sg��u�~��?��LD%���CT�BGަ�5C]㒺�'����S�������#)��B�j'�����r� �9�{�A�Zǐp�n��&.%��?��y���w�;���J>�,��x!��|�N[��e��������wp8���c�7��j��[�� 8�L�Il
�24r`�3)߻@.�ղڏ'�����@�@�U$¶)h���B��+�6�4dt���/�j.ԹJk���;*;��w���V̝�{�V�:�e�mo\���}��kǊLc�6�،��mvt:�����E[�Ez6|�R���]���NJ����Z�̌�a�>�`0
q� ֔ۜ����_��c���5�r�[[H6G�,����"�L�咴���m ʺ`�(X/�K^�t��Yw�k9��{=O�Y,{E��t��}�`ؠ��ͳ��+��L���
f�(��G0�W�qd�wyw)���r��(�)T1�t�[�?5*�2I~M��JP��ƁT�aϳ���r�ؔV9&�̢�)5 �,�
�vY6�������������Yx��ծ���<���J�\�9�٤���m���a�W	��e�xJ�{�"��ҫ44an�ٸ4NBn���Nl��5�u�?�e#�\9g& ��X��ʙ�3笚�ڙ�P�-���v%����D�=+�JU��b�CLo⦽�:t�Ĕg���m6�����Y�kzf��N�R~L���B��T���G�gtU�aN`�4:Al�=�u u}��>"��S���OH�澿#��9�����6=�/���k�Ց��\Ʈ��k��V����"$!��2$/{��oZ�-�r�B��o�x~�[o��OԆu��R����TeD@�Z�jM����E/<�S���M�̔��/�=���T�#�W��
%jJ͏��UZ�`w����<V��g�3NG؏��#K��HH�����r�ՕdԱ�L��и�Ш�?ս%�gs���5��^C�g�9������`̖nO p1W�L~n
XN�h�?D����<�8�Ҏw��p�9��>�+�g��?Z�p+�̫��Eh������y����f���]<�:�{	>
4�|B1�XuG�#_�"����O�׭�ƃ��M�B��]6��8*)�r���DV�� Me���T��ńC.�R1=�'�̡�9^��oE��f��*�'u�D/����g�X&�{E5��m[ٶȂ�Q*}�I�H$�b f`̆�e Ĩ�d;�)#I�_�����Y� ��d�z�siM>5� L/!o�)��%P�9QB�1���y����B\ő�
�`X�o\ox,??|�|�)h�T������(��P$:�-���wB)���4s�}�ն���a;.�z��aم(q|�S�M��~����P\ ��ԝ,6.{P�ZF>�Ż�]���Y�OUk�S���qF ��J.�M|^#�k�s������T�3Ѱ��W���3�� ��	��%A	�.��������R��+mw�}rrnG&7o�������J@eˤ�A��MO?�"�K�y��؈��,0�wy�) t��N��r�~��� @��o�s;W�t*������a��S�(˕X{�{��� k��?_.,y�6�:�*���q.��v��<E��������P{rҁ���(�W����?!��;�酬=�	`�0�Sy� \E�N��ݜ��`ϙGX�(�2a2��pjȳXͪ���XNb�1��v������k�?$ ��辔�5~�M8�
��,y�:I��wF�PZj���i��	c��B���f�},YjAĝ�b�s+�CK�n��f�S/�E�n_ي=YbO{:�U��� N�E3�	���#����˿z`��`f��L=�Xq
cJ��OD
rt4}�	�[�>k"�w5Z�7?#�~ �폺b���f�a�,:��u�j�^��L8���-�\�:����&��j���9>n=B���$��|�|�Ӱ�I;*@�Y�ӥ�Pή�iBè��۟�_��b�-�@���z��g�)��4!����^;����j��*h�Z��קA�<�|� �H#��
�=�m.R{2��ͅ��,��z��Y�y�2����/�v�o��{�^.~@CE�D[
��3
"���/jA�
@�&�o~i�����~,ϙqf������@Fa�_5�� �I��z���^,n��X�6
p���[��6iT,���t��cwr�J��&z�D�8�����9�v(3�]V�F:��k�ڹ5\!;��$��8��������ue�n�@uzx�W�3��tF��U��OF�T�;[l�������5%�\�ˆ�g�;1Bf��;)� �4-�C�Z���ƕg�|9� �X�9������wO��,B�%�	�$7�Ϧ!i)'�:n�"�������;۠�A��2初F�,Zr��8k
��^��xԸ-H�\�$S��r��=h�[�w��3�އ��z�[��&$�7n`�'����m��&$�&�hN��㿽���º1VRoQ�s
�h���g���$f�t��݈���/�_X'e� �������r��ơq�L#��Ձ�)J1B)hsG�TY�;5x�s��+��50T�Yn�����!�[�c���@���;���p#�����x��[T�l�ڢ�j��0�Q!��	��x�'�	$�*5b
}.vE���[���L� XK���\O81�͛ʲ���_7s���%SʷUco�'���g,O1�6��6�
�9#Z�%�jJ�]�*���jG��CJ���O�_\��R� �6�ة��u{�4�*��lP���֌L)�{j�`��0���4j�@ա���>W��Â����	$%:D�1��$-T����衩��S�vZJ������u�I�ʺ�ԣԬa���$ӿ���U8�5{��#��X$�iy1x�e�8�*��1c�͕���{�S[=Der驟2(҃�Q�pr#:Έ��ER��=�+c�ûQ|��`Ma;�ɀ����[d<��t��mW�3�`� A,�[��}y�7w���l~9�j4(�v�XV^����6��_WI�����D�������1�̧�`��xv�IӢC���eK�m@8'hu��]�?&�ߘ��F��V�h���@��ԅW�k�黟�8�+�l���0������-Fft��|�wW�b��`Tә�"��ܣM�N��^x�a3�B�E�`�ҪݙU2x���6J\����}r!�r�c=�����/�"�_R���!���K�k�k��� �<'� �.�{5�GK�CLO��H�$V-��n�Qg�J�#�a�B�3[ǣ�5�Y�V�`ߚ�% A4�!'t[S-t�4ߑ5�]l�fӝ�F������N�d�,P�&��%��eXaW䗌)��q�e�m����(R߯��IH/KXm������������9����[�B�m��aF��縻��Y��X_i�؆��!,Q���n�ƀ���{zj�ex�o:U����p��zN�񒊯��w�mVD�=<�k��W�N�\G|5��̓�҃p!�����g
Eی��V��5��[>���
O���o�����ԑ ��g#j���[K��
�1$�{�@@��J�QYPDq	H�X[U��^RS��0\�:a���WT$���/c:�ފ8��ۢ�a���Ћr��n�z��Xh�,�"y��C9��w����9zO��Rb��\ƄE}�H K��*���6ÈR����)ڐ���F+���bͧIv�'K!�MB�e-!��Q�\0%^K+���h��}S�)}�I�Q��
aN�m����ۛw��O��\�m����'�����˫� �t��ų��ٝ@W@��-
4,c$��k��?���)J����C��_�x�:��*K�5�t\i��݃�7,��ds�uxw~ᝪH�`��P�1�=���7��V%r�J�A��հZInQ�Y���������Sk�[�O1��EKز0�PF�V[:P��x���F��RE��[��:����4�ht��#�Rs�ՀS?�#�g
�+���$�!^"P�D���Ԁ�[��x���l��������g\=C#�^��2�$�'m�b?i�9�\c�B0�ɚ53���%u7�׻�پ���?.
�.��$��	�@�����ܳ�����6ق^f�- �d���:(�4M¸
+m�hi(�@϶�u{�ZfnA���cWvC],�˚B��4��1?����=4=͌����ȡ�Cp2��c�d���P�}�� rDJ��6�s	i^����R~��ӄ�����%�,^���T�8��V�c�m�t	?��'����'˹���7��r�&���B�r�C兠�F��S��Ө�`f2���V�v�E��:�|� �+� O'b[�Ɗ)p�z�.�:GΘ�?�,��4h�//zO9��i5�����`RI�p:d5$>�����E(����N
pj_
Upv�A�0r�����<���ox�6�;֯��ut=�j�y�M.�����&��!-�m�����@֥ �f?�+Q|�d�	�h�Z��j��Bݳ/t�5\*b�G&d�� ݖ9�r�|�C#�mE�����*S{������2R�v��fFN��=�\�B��<O翮1�9�)p����#�l�Q�KsA�R����:o�ٝ��k�{R�]�گESH�~cuZ7����hhN��Y��ex��0�H����E��4�p~��F�hh���W��ycԤ�x[�R��Uة�I�n?H��'͡�r���	;�|k�S��K��!���/cŉ�R%ak�;g���OFrP���=I9v�k����c��w]�l���ˆ����[�����J����`��o�x
Q X/�����(��c`��.W�f�6��8.����ԑf�������A�0ڔ��['��Gz�M�m��r#;�6��-�׼�����Nĺ9F�������}
k؞U��� ثy� k�����;�w �	Z�����n��-L�\���z�c����:n�#��6JZc��[�~�1�I��y�s�>R��M�_���k�E�W{�He�s�3Qo?8"�4!b�����J����	��00l��
d���Ʌf�ٲ�d=!m7SaW9�1�y�aӺ���'jCi�)Қ�@"9:�_�Z'La���&�"{e�*����V�N!�!����L�9�D�LW�!6F4���_���a��f�.�߰���I7�Γ���rU��';�̲�te�!�
~�"~ꀃ}�Ee��n�������U�ҍ����ޭK`B9Q���G�&��u��::KJ���예��2�7gw5Y��z_3��%˘�� ����6JL�xT���4=��K	���{�gذ?���/��\�=~����Q���J��%�ۥ.�����B��K4�h�)sK�@Y�Z���
��~��,�_#A ��"��yo�1C����A6�hmD�'ç�4O������sX��#숋[��P�;�W�s!k�:�2a�B���ޣ���x��o'��MJ
�1��8��-�o^�0��I!��땯vA}G��y�уz!>! �ǌ4�u%�y����%&a���������a'����5��݊<�0<b��\P�Z�5�h�/x�>���
�]�0i� ��5��+{v��L�-c߫nV^���FBrGdL�� ��e0/�ۦ�&��+��2�ej۵��qX<��]4@Y�x��:.���5�w���s��Ӽ�X;f�iF�RY		�QN�5�1&	N/
�1��m���b��H���Iv8H�]ZXQB-��q���L:�I-��D�v4� !b�v�J�o�)�&�K#�O�7�F�9g@^ޤ��ޥ�ˎ�t"������lڣ�\�zw�f�Fz2O&����I�y/80JH�c����l&K+2�������yƑ�^��r�T� �ǈ��C�7���mw�>�&�*��S�덭�L��B�ο�U���A�˦���D�q�;�A�K����	��~ U4�11睧���c��oUa@Hޫ�0[h?q��m򚷄�N��s�A�-�^���F���[8����TH�]ə��G,��ՠ�4L���3� ]+������Ył�ĩp.W$.qV�d !L�懩�!m�=Ɏ���'�A�S���nª "���NM�Ӛz������n�w�Q�u�A�VM�C�5ԑ|@}bM�+��I�M�C�������Z����[������g���V�jNC��Qv�J�0�8�F�-
vZ��I���J$�P؋{�0�P(	��d�G��Z\8�!)d >���ߏ�g}IP�K���rJ�����9Z��8���+��gU�<.y.o����d�޳4GK����[V'����.�P����6d����1n'G8zȥ��8��ԭ@�����_Q�G[t����@ns([�K4'��[�Q�j[�V�AM*�ψ�7�|�y�:��+�ؘ�K�b%���K�D76�:�b��K���oT_���tC���گ8TZ�_5xp=��`���t�RcL�Ƌ>����藬a�;ypC<��5�k���Y�K�-�$ث'�Q|Ѵ�z���$�8�ː��ɳ�Ɲ��p���\u�P%8�3�V��#?|w�a���SǬ�����Z$^ۦ��Z̿��LPTh~�"I�WM�v���b��̃)�Ս��S���p~��C�e�8_S�ƙi���r�P�ˣj�Y�>��u.ݳn��n������ǘ R}���A������.����k�O��ΈK�7�Y.��?��b�u��9!W�,����6<�����A��3�i\��#�S�΅�f79aVT'Pq�/�䯝`�����W�C޼�<�i�|�Ѣ_��+z���oR �?�9������Xܙ���l,t���	)�g�cY�~_��/r�Ԭ�n��
O�s��Z� �bժ�i�������{y7J� u<�Ϝ��$ϖ�T�mه}H@�����J�Zvc�j�s�و"Jz8�%A���p8������۷�����n��[<��~�G(.�(��b	��-�ʋ��Ы��Q���2��`�xP:����2房W�Qzi�<��펙P���j�h��i07�i�������.�Cq\n��e���C�(V�f�(v�������.qձ��@��Xچ���m��U���ߒ'�g�uW�i^�����L���moOsg!M���dm\��)g|a1���������̌j��2���X��dj9j�}���01��ʇ�jTyV�ՃS�;�k��2�<�k��T@
Tڶf���	�%��������+�D $�P�V�a�<��je�@g�g�,�ݱ`D�1�&���GK��z+O�I5B���j����֬�+��z���d�A�c}m+w\�܂�d.T�|���@P��א�[TI��B+���� �ts���l�Y�|>c3�;��t$��K�EFΑ- g``ĞG�(�ُ���m��$h�Ox��%Azv�Q����!�m����gv �����sj3|�$h8��j���G�؛#�Ӷc�I�އq�X��m�`���Š�����y`���o`D]��(Y�*�+�yj���=����T�Q5?�_``)Qh�Y�Hk��O�䫪�#
|u�� m��n��Vӽ� "��1��;�)\�G>�v������}t�Ε��VW��I7�֝v����8�܅J"��V/�R�J��	�&I%)�+�G��P��$�[P�����=�x�޼���T$
ǁ�9J�%1F�GMLB³�'����(�z�$W ��5�0�/P,�n���)SR�:Y7���B③�] ��7'��r��E����u�n��E@�
.�l�mr1g)���U�>^�6.Lp�3l@�F�QA�e(ʥ�zmآ i�`�鈐qN�@u󙙹ޭ_-؈p�d�CQ�ы�_��ӡW�0�Ù��o���d�JÜ�#r6�>�<���?Z����%���Ş�!m�p�P������E�u]Of���b\A"$ ~�M�����1*��-�j��iRW��q�p�=q��=Q�Bm���kc�qGhQ�D����3�|�i���DC���ik���(�]�ƕ�H��k"ų�~~p%�ʕ6�I�t�?D�d��,Xs]N�6��0V�J����}�S|@�t;��� Q�3��V+�9��Jc��J�p$�ک\��tA���v����)ui���3k�����%� ��Rặ��C�x��h�����M9+���y��.�|�;�#��w�����r5#\F�.��w,@ ��%�C��Orߣ� �A�/��v�qt�6�1�#� Cȉ;|��&N%)ݢ�/�PTj)�*Bdf�B�V��l�j�"Cqb}ϝ1��@T(��v� �K��>m?
趴#� ��i�<��/{I�,�ƻ���q���'��Α?Y�H���t���҃}�)I)��{)��H�&��4�"��#g�{(�`!^�<���x��u%/o��tU Z�M��Q��<�������=�0f�:�x&Mji{�W�ei��t��c	T
���a����!���H_Y�ԛr���c�����z�6�ݘ.&E��N�D>����[�ز�U�*e��Do3H����Z,��������D̨N�<hժ!��F}��8l�^3��\� ��/�Ƽ1$��(O�w4�~�t�H3CU���/�zPu5�'��O9�3^��!�n�����*3 ���a+L�p�Kd�R=��_MH��$���5fje�n�\h�Sn�����(��Mğ��՟����:����bӣ)�	57@� �ؔo�����!)d-_�I�VыD�����o����FWh�����lsW�l������nt�'#�L?簝�Ϳ�a����6�_�U�j�z%c(;A�,qe�V��Ci���d��rW���N;4�c1
_}�+v�cx�6o�x�\c�kaʍ�*o��K�����N��%蠔�Keq6����rV8�:��M�x�5A>d��
�n���^��!2�34���J�I���?(�5�Vw��2�0����47��f�lw<
���P2��o<9��x_�-��*$kح"1!�(�� ��oȚ���+j��,�`����7��V,������w��.�R���C^�`a����j]#߱��PnN3���$iH�!�a����[��z�,V!�ȝs ,�[kb�G+���Dv��lA���V1�/���H
J4����p�@��hH�1��8D��S�:�M���[�b�\��0�	�>̷�a�Q��,�ܒ,p�Vӱ=�`5�#�E�8�V`l����2�| c�M���<siM8�e"'�p�z��_9�o_5z�`^�C�j&|��h��;�^�v����RGO�Tv��ٹ�P���-3$����Aj
{����MS�^����s��z�A�Ӱ�^e���J"t�,�l7u�DP�[.h�x��c�U�v�m��C���QH+́���@7�E2��ǥ�r�VC91��@X�N��H�ֽh�|]�®?b�jUMK�Cn��@�	:�����ʹf�%cam'v��g�9�Y<�+}�ޟ�xA�ƚ�Ҋ."�g�zrɁXWo�5#Q^�sї,a��V��c���廊����x���ҝ�<Ug릤"gwL�k �	SimL-��d�RsftقEAf��m����
��/���2L��h��F m �Pq��G�XH!VXi�� ~�c]f��_-i��/u/�i��Pb��pSeNP�X�Dw���ʨ���g���j?iu3��=���^d!D<�DsH���@��l��HoRnQl���Y���KL�xU��tv�޶�x��r�C�T� "%�-�h��}���_g�7��ӾGS"aj}�-�<?i�7�e	<���/�< �0�I�CP�K��̒~�{�8z�:�V��F�V����FM��e���]�*�M�b���U�#�9������X�p!�M[��׵�Q��U�,Y�0-�4�J�@���^�o1�ZQ#������Eޭ
$$�R�����\\�~Kb��(b���~Z�%+��q��=�:����
z���{l@]	� o
Z�IKAs\v��j}3SWIt�?^kz^�V���&��Q��������#��� �Y :�矣�*��� ����\ҷ���w���~y��LPAu�?/cu��1}sk>��w�.\U,��9[}�B�- A/�Z�jɭ�*�45��?H��qY�%�oJ�'�&a[Ÿ��۔q�������{<V9�P�z���j�<�R�k��5�g)p��8x�U�g���Ӥ�LLC?�2��J���� g��\h�]3�eS�y�NY�u�FуkaA�ar�_��t�����!����~(�j">Sqk��h��ẋJ�?B���p�L��1�X�w��/#���nk'������U,7��`�`��L�t;�.�^�� �[����pˈIJ�2�F��,f|IC0�^����;8��č�%�0=��y4) �P6�K:�A 'RL���	�v�}j�Ip(���I��` 0�hª'NbC-ꎇ]T�H7�����5 �!s_d�?��+����JCV��0����� 	�R{e��k5JK��}`�Q���f��Yw�IM���ȴ)W\ι=)5���Wz�NS�wg^�	��΃�F;�1O�9�t�|4�w����k�g~����ˑՆ����s�U��J��V�k��!U.d�,��=�LV�'ʟ�?�#u��~c�@Qw�>Y���m��&����B�zfw��%T�.�1�YI�����3^����*�R����Wrp����h�$�")��o&�Ve��k��c���dc�9��s/��K�����%WN�r�uk_?h�Ӂ��ÿ�9��w�2��!��=Q�<���d�P$�rAe�$���i��,���.���a:�p}�C���c�-����fق!}ݬ�y�,�f.[�ن�9���$�;�"�/Q�Mj(T9!}�^���m���P�N�
.�ӛ��o�ވ�g��A���)bU���o��Lž����%��帪.�L5,`X��ߦI�H/\���o\CEo�|noY�(-.�����Ӗ���+$Q���nT���آ%�H�	Y���e.������y8��0�*��|ඬ������+D�:1�����2�S:n��Jpi���q�3 (��Y2-�d@c\)p�"����+U�ܪ����i(�)��|�F�!���4�d��h?e��ܰi���j���|e9CyW��Y��N ��+���f7Y]�r�B��^�^����Hn�	 � �l��.L�ЪG �j��l�:���c�����P�4��Fzǈ��`�Vr�탅�L�'�0)zV��.��4�̂��{�� �ɋcT#�V@�)ف�5L�p�g�@���&C-��|[{٘�R�R�YƏM��ckyd.j�2K80G��r:E��>:t\�x�&��Ί���C��\iQ���ڻ�[�2��nItIN�m��9ah�#���:���x�$ΛX'�M0BD��aǌ�1O"u=��JC�;1N�J�&ʳ��>=�)�oJ#�R��Y�Y�%��Rx��m��Y�p@�y�t)Tu�c�:���[{�6�X�_�iO1��.�5	
_��~�g��٨Ϫ��tM�ŭj�R/Z��c��n��6E쐑� 	�A""s��=�,�o���IPd���/|*�
��s%9�^ׄ9�HC�-4�k�Q���������!1���;�WVM��^�YI�dn���o4���$���!���R�za({a0¶�935�'Y��+�B�xo�r��L� ���b`	9�8��oM$�0�v���oH��B��O��4�n o|hH��gUeاU�r?��2����A��`�[1P�lL�٘6�\�a�hPvq��#Qn%�d�ʱ^F9'�-�p��w8>y&��7L3�|��M�c/Kܜ��ɔ�{.����5�H�u��H�k���Z�Ks�E/y-#�B���Ý�\�������n�1}� �uǙ��t�߷�f~�8�!C&F�7���=]��u/�PT޳\$$/�	����8iɋ
��,a��4m�8B_{�T���it�FTi%�[�
v���g�����Ł#wY�+!�G���oЕ��<CM C��
|�����*��3.P���s���m�v���S��%��0���K�F���������L?��%��H%1��������j���~��v���\�Sa= ���"=��%�?�P5��Jv���y�0�Ì&���c����[��Q�W�óc���|3pL�����e��]Mq/�
q�(�8�LT}��8���.��2ߢ^He0���:It�b�^y%���=#�Ry贯h{%�1%r�s"G�_EFO)����@)�ҝ���`��Q����\��(�ȯ�ĸ��|�y�/i"N�m]+�7k�8���d�'7Mы!5 ��Uw��Ew��F})�s�b�x{
&v��^���w${r/b���`�l��۶�8U�����B1uv@U��������w9W�}e�����~�0���"CԨ�����>�X}�9���s,��;���(�F���}� 3@��LMw��(�(MN�~ѧ�,�/���4\{T�sE)EA��o!a�
�V�WE����]3\(��r����P��C��#��m�!��)���Cs���N&�d����6�$��;����`y�,gS�?����b(��9�
w~B���tP��v�,7�&Zg|�7{+,���i L_���-��7>P?"R(��y�w�Rxwq"�VQJ�ϡ�:�k�"��φZkh�L�0�+�x�@����R��~��)t�#
@�h�c�Xp���,�A�3�O�y8kU���� ^�Y�YǶ�3�L�M0>� v�5�;=B�5�����l�>sXÅ��'�G��c� ����-#2�D�)���Q�,\|;^����C��M�m~5��<�&�s�j�M;lLʈ��T>�t<���@�Ҙ1�wT�In)u1Ç���I.'4�C�YU�K�P��Z��$V�'��"�f�HTqȈN>O��I.�d~�����"���w	-g@''{�5��%�ܫg�`N���+3��������֦�Q�[�+n��e���w-����	6���ֺ���c�|M||r4�݌H8n�yC���h���W�P��Rv�ԁ$ЮX�Q��+lc����|�N�\��!?���oC�T���G��@A��;HG����t�z*Sg)�L�a���0_�}��K�� ����^���kgP'چ��nǀ|�<W���+�v����4%��iPHRdm�+6�׏h�<A�:�Շ�1~�&ν�%;� ^�G����\B��)%7�%�+��B�h��ո������R&��۱CzIz+i��[C�{Y���8�7�g��d6z�=ɘ����R��0
AJ�F`E��
5�*r3��%왴��?l~(*�E<	�am�s����"��ǎbj3bx癩t�cvl�J8x�}���f8����9�(�-�7.2S0J`���)S.NGO��aߩ��l�/��<��>o���3-�f��%Փ,�E*�bb$o��tj ���S�,�˚b_N�څQ� �7�#�!�w�y��V��n?|1htP#~�7o0u=@mKA�m�2z�8�Z�ȱ���υ�u1ì�i�q�Uo�?�k���h�/<&b�h<��;�Ȑ@��&W�ӅށVK�<ӿ���:�0�۪0Yқ�ŗ䟾"�� Wc�&�a=�E����C�=ty^Op�H�%�����-��j@�rЉ���u �p����_������ޕ��$S�Qҵ��~�'��-ǎ����8�f�,�E"�#����\YD�<u��	�$�[�[�또���W��S���,�_���������Ŏx~ӣ��+]��Y>���ow�  Q����<���kXs?�竩	��4�D���Dϓ��	C�F//��d�^e� $���gf��Z��cP��ps�_��XJ��b����|�Y�*��s�Q���$O�r�[m�"\��?����AQ�h���G�J��ҁk[�V6�^�2��&�Q|�0�,���W3*�Lf�+w��$?/ᥠ�;���E�j�{�D�$d��#,AGBٙhӬ`yo��k�5M}�|}T���P�l�9$3�Eލ���j��	`zH�,�kFs��;8�$W�h$k��I�0cHH/��ô�%p�#%����.����E2��s�-'>��9�]���U�)����9�`q�Q�~��x_.x��@��d���Q]F��*/L'q�����7w�4;^���iu4ep�6�z&Ib�P�ၐ�-|힇����u
?ĴV~
��u�9ԃ�W&D̬��O��[k�Q,���Mr���[{��*vT�9Wj��P��*�� 9u`�z��;��%�y���;�����np,�n�8��<d�.�zno5��IR������1V�ڱ��p�(��߉Z�X�������X�3Kv�L��:���M��#��-�B���;�}AHfvk�OԲb�g󡧯^EϷ�f��C�{��NWO��f��Q��G�Gm��N�@��H�ڑ_��D�\��ҒzŃ,�{N�_��U�,ݟ����d�F�!r'�O�u���ݪ����!Fk��=�]��z<N�]�a�����G6�P҅i���
�Ɖ����|j�9֥sD"�������v�-e�|͋[|[�D�x�H#��Ca�Jj@� ^�8�uB>���`�(s����W�r9�����'qo>��;��w��~�ga�����#����폮'�'�ږdcwy�nQP���ڡC0*݁�Q~(����#e'��`u�"�����n��f��Q����+���t��%�u���+�՜��<MGY�u������RrJoc�`Ј�E�"��A?��|P�7_�PϜY�����pD6( 䟒Z3�Y�Y��;��R���ɗU�ƻ�N:v�ҍ�#ih���o��v��� �<������0	��*IotY\f�t��b�"4'�z��\t��<)��*�.�rU�u�J���K���=��I
����n�s�X�>���.eT�4�yuU[�eU���=(P�J�E_�KH%�qS�Dtg���s�A4x%FInx�;e�ڛ�ss'�yAwA\����r؁�B�n��kۖ�����'�8��>�$}�h=ه>o5�aaD�m��%C��0��B�`Ƽ{#?����rg��^&l�o^ *_nC�<9���2^;7U7�,�%+pl�r�M��=B�r��,�	&`��w8�&�K���F5﨓Jܭ]B�u4N�
Fș�_���ư#�B̔��6߈���3M�Ӿy�5�`��8~�ڭfs4�e����sޟk�I�a�X�
QȒ�t�=X��^�2l̽*����t�{/��}�����>^�Nڡ� �K��0>"CS?�B�M��ڞ��x�te���
��$�sdj~�-��4K�y+�cjմsJǂ�C	�=A�l���`\���V�5�ڶZ�t2�;cb�jz?ۗm�+h�����#bQ�iR��Φ�A¡~��	<�Lb�HMJ�!���ä'����t��y�q�xd�GZB�8#+�N�;����״e���
�����:`h����)��we�6$p�����#��x�^0�Bz;�2D_��e&:�S��1�C�*}�³����-K�7�BZV� ����%N��|1���7�	2�oV� �)�V�=�3b����@��Q%��s`���"z�Z�%`]?��<���v?y�����5֫�4���-�O�hd^i�� �|���j/�_m��� CQ�5����R4�&�ΚD�6��<��t�e�.d��-�Ǯ�#���^���B����e����d[\�|9>4����W��:;�)w��Pǈ'���/9aCJ*��F�xh�V'h���,�d|@���6<��۠s�yBc2�FZ�H�iY'G.bRi*Ƚ�����|*�l��yU������� }��f*��*z@���Ӝ{��Y	�@�E��f�۝��[C�\_퟊w��?����͎O*{d����Y�C|����`�n�b�mw��5��Q6z����y3��e���L��p#)����oR������R���Mts�ҾC���StI�Y�!=w�n)��FU�|��J��#���*+/!���|0��Dk�F��̹�Ё�:(��3.y^����+(;͂��r$գ��a���ǐ�u���Gy2d�Mr���>y.��Y8��.,:@���o�Ukb�V�6��M�*/͵��_Z1�L�oJv��
��" �P.�"�0�'/i�X辫{f�J��\�+��N��I��$TP�E��S�h���;�pu=��"{8I<�T����N��77����,������%봼'uxD�$��-̦S��o!ϰ�_BK-ri5����_$#�R�^�T���.o��������d�ŅӾ2�0��vͰ(�������Q �P��6��F��}h�<f6o��o����hy����
�4X���B�ZEC���k��fs��4�)�gͨ���8?Yλa�{��o�{q�v��3	���j��V�ʤ�����\:�u����ֶ$\lB��WC:��p�G��x��꘎˅���-?�`?(�)��ꂛ����2k!ư��W�>�-T2_ҚP���~`�U#�d~��u��E�&�����Lh�WX֊D�E[$��,��0O�VD%���Qs���G떿��v���� w*������P%���(t	n�����r%u���d9����?HR�~���N��R֣��t���OL��z�r&�g�M32߷�T�.s�x��к���$3�KW��ⅾF��M1� ��4[���
X.��D@q�<��:��7���U�"c�i���W3���E�M�oq!Yʈ�:>Aύ�P[�n�w��BQ�jh��dt�D���i�[���&�Zu�2�O�X��}W�4��]Wk��8�#�Zw��Dg��z9�R�>(:���,�C$c���
tB+�aVU�>Ы�����'a��{3�.�A��Y% /�;Fe�dh
��,�'Ð�����7f�h���T	l3��JOG@"��sB;�Nl2T�\�<����z��Y�%2Sy�E�0�b�Г���N��!�ʮ03iMιn��-Vt�a	Y�F~���OY%T�(�Pc�����0ud��˟��}k�~诌�Վ:�Q]����yѥ�y�gb�ջʙ���MM��o��+¸����;/K��h�ѯ��䝊Ŗx��w�.L�Q�_������0���tr�:R0���E���_����Ŋj�6����K���e
Ƽ�Š3���)���y�M!���X��#�[���pN�gO�㝨�)i����2��  ��#w�"�M/�)lq��l|��a�p�i;�}�E!#�@:/�C&�.B��/,Y"��K ���r���8�/t&�Y�>!�#����L�\������,�n�V"�b��RS��j�=).��]_����9@��]�X��aP���kx	���� �rR�?o����x+�P����-�z����?8�G���0��������g'�mBщ�b%q�k������/:&o�ø\�%z�'s�����_�T��6@�C�B�6�9`�J�͉�`��1�ht�)��7͆~A"
)��r�@�SIn` ��LΗGH�u6��!�bR��˩�c��>2��a��?H�(eM^*X ./��Q|��c�����2���C��.I��)�DbH�ϧ����G�/o��}|��D�N[��q����?���>�8���YyQ`�E�-�[��9��q\�A����#xD�JQ�Rϝ���[�x�5����>���jzn˸,��&�@�����SP @�"�t��g�j�}�/�@���4�	�-���k��$�"�3�Y;A]u�|��.�� 2A]%�y�k��׳��@vХyY�b��@�?���/p�qIQ?$׼�8Ur� ��*|����]U�vO˝,m�MPP�T��a%��y9h`&Q�u�0qQ�� �X�-�7��a}APʣ��`ҫ�����서�vn��Ǉ�_�����-�������X�娬�0�c"&8�9=}"&�0cE��|��h>uD�H��p�h9��6�x��)��];���m�q~��4/�M``�h��۫���`�����&CC���n,���-�++���L�l��É�P�=�� Dn�F�A��7��K�u����S�e*�P�ʋ#�%�Q���0Ik��c,|�ܾ�wK���;��m��;WhH���'v�L��n��'�}�p%č��us��(^q+��q�ر��U.��YO�k�:��kx�� 5���؏��[�~`uY�/\Eq�`��KN����`sL�<��%ǐliN9��Zz������T���`���߮>��$R�9���f�'A<�m���(���O	gDh6*��܇3,����/�9��ꮳ3<6g9�2S�c��w�?���ǥ����)e��o�;��T��>�#���Fh�Mr��d9r�s�m��F��n����o�P�,O�w߿V"��#��������7�bz��4��-�`}��1�&;��c4�8�ъٷ}��
IL��T���琪���E���R����'E��*��(�7*G���af+��תhH�k�P 3�3܃�Ԣ	Ӻ�N�VO�M^��RJ{(z(�E�҆+F� �9DGh�3=j�)�[����#J�L�BZ!�f�-��NI��֪e�/����YR�3�ܗ
�LO�x|�jt�D����\�qD��M��u�������Ѭ���D��h�/e=G�wdqv�r"Qb����~�
�LJJ���������2�ӣO�!��
�%%�V��z�Z.*g��<�U�Y�6��X�T�!��4
��6�$F���t��/����X�-2U���Ȁ{~C�_�ɣ�z���l��*����ƴ7��ys&kh�Vj��xwbDm�)`�&�im�u,x�؅�WWe�iH�ך�ҫy�2�����<�8�b��,O�֩�m,��'�V�������\b��1i&(k�x���s���!�M�(|2��)��!�銑��z����5�x2��q��ɵ�+n���%�ܙ	h�w��Z�g��6&��_PE�',6�S���g:<�W��i�z=�,AH�	Y��e1HPm�짟��r˓v�l-�P���+v(h3�n%u�F=�l&(n߭�$}�̨m }�]�(D�֯�f���e���m�aAp����R�{��SI��$<��N�(�
���tQ�!:Fp��5�!!�>Mtln�nU����u��Q�n�S�mu�t��o��Fe�jy�Ŕ�ru�z
b�$���U����7�`�˺B�$���ʱF!tɹm�]�KM�)�`��b�ٞX������\M����-�T��I�Ni�7	�ӑ�ͥ�'�ot�6y��@��f����]%�;i+�z]���$��zٛ��������{`�Ӽ��3��	[5�R�P��؍�T��X�^[w n5�2�07`"�]�k?��t���ua������;��a �R7i�8�QE<�wK0K��g��h�C�q�~@�8AD����8=��^�/���0�n��bCy�]�ߋu�<����{9��P{W�k���U'|�
��Hˬ�S��WS�Ӯ��hu�pj���?�k�e:�:g���7yr�zH�nl�s;ovpGto�>��T�?V_��O�.�Z\��޾�W�o�i���k�AI�b�9G�&��\Lg������!ܩb_�3i� x �`9e0����.�ܑP��!��S
čvȷO�CW�EF��	Nw�I:i��!ɔZ�r��P�=G��2%�KW�E��/-]��F��?~^���5�����@�kA�
E{��K�Dt��ER�}C2��!VV�N��0��ox�HCw�h�?d�b�����KL����(������l[��n<復�n��ʧ�fiB��HT�J@z��m�k�]�8B�����f�rXc���J��t�*�x����}V�����m��ǌ�j�W�i��	.�-�����:�t�*��C�I���g�gKw�(�/�/��ѡ�4 �6k�C=Q{ʐ>v&ZhD����A	$:-vP(�1��W���o5��M�Z�ML<��1>ϴ<�9s���pl=���e噾=n�QA�][t?�����F�=){-�|fV��9]�?��o��{�ū��*���$gu|ėW_�v������^���O���~m��Fz�v=e�l�39"��|r)��v�Ҁ�{�Yp�ˈ�Aг��������kdd�[�wkP�2�����&i�j���]�_�>]׃�z1HKp��oI�?kU�v���"�dW�hK WE���S�� ��k,ƨX����-R�͑�fܞ���y�
,�ҫ�J��v�ʶW�l��	��}�&���TȸL�,��⊴-G��[O@���(�*ӏ@8ix��GJ��c���*y�Kk�5>�����S�҄��rRH���#�����`>���I{_��X݈u���$�E�����W1����=*L�l�C� �<(�0LQ)��V��c��6yY+b����d�	`�0�\z�i\�b%���u���>�\�m������q\E��e�T�Ε��0
�w��U�~�[��"w�|�m��y������}��+T����ȷ����,��7c&_a�.�:�ve� ����2 �&��V>W��1�>�ë�nzI���k�k�������Ä���tU��.��C�b
������)�ƱI�j '��|m����b�k����˹J̉i��
��}��/ ��=�NW��O���j0����oCR��aL��-d`"��D�5ۜ9�U��[�QJ"ٿȉS��V-�P+?gL	�K�Ԯ�x����T��l�`�94��5M�xw�%qՍa�0b�Gkj��E�s�����'J�:g��5<�"R��n�?�p��8��{���m�Ͽ�X����XDlV@@rAN��+ȣow#m#�t�{�Z^�_�j2פ�]��������ܝd�bR3F��YE+��*_�~�Ś淞�� <�Lw�����f?+[0�(�3<g��B,b[,��z��7�'�"ˍ
ң��=���3�6�x^4��HGt4����a�l�Y|���e��" ,��c L�v�Uk�K����e�˥5΁�d�pkZ��D��[ܻ��c�ƃ�$�3�ls��� ���4CA�Cz�D�QX8��Z��:5�.K�E�E��)nw���c@��Ƹ�}�I]��+��H�3!��������_�p'��[x���^c���M�R�B<����"P�G�`�&"�Ĵ&[a6��j�H�2\,]����EaT��`/�O�0��$�|�~99��q�<��hk\y��L�/W����K�v��iQ�'�?�L�.�����]�%�7�8�Ir�w�yf"��a�w7�f�G��E��gI<��ܽ�)֢���p�8��bD�����;v^~�4�!���@��as���yX�"��z'���=~o��C�7k��3�ŋ*N�
�Yy7!E�,́n�����Z��v��$Az\f_}QN
����E��~Rb�]�G� gC�|?!9�>��|����ޏ��j������t��pl���ⁱXDtpaWeiI ������
��YՎ57z���y��a��~�鑘�T�^�H�k�@�����!�B/���/��;��L	�^N+�؊H�-:C=U��6~��|���n��vۨx�h����wɹm�z�Y��̬~���`iT[��~F��T$��==c�i2 \>�*`!2k����L��6G�����u������d�8���%q��w��8�cbKg���p]Pӵ��0ZJ��5j�����J�1A7�e�������7ԝkO�4�"�uS�*�UG�/V�N?�]9�=�p�-lR��κ�3D3N2PW�������fp��+�}����N�?�Y��܎Մ���Z� ac�n9�ܮ GNZv ��ݾ 	� �<o�@Y�0߻�0�,����( cd4vN�S����BC>�N
袸8?�r�}&P�Y����Y�ȱ�2`�˗-���FH���M��T��rV>
L�t�[���a~�j0C໼���������P�!��;�;��I�i�g�*��T���D�k���\8���� T;��c���HЍ�i����[y="
�~[�G�m��_9�@�3yh��l��~��/ѾԢZ\���k�����`�q0D��� L�V�{q���ᐒy��`��M�b�n`Pvu��MU����vb�P���#�F�F���!���z`�_f�Mc�	s݆uN4&��\Y�@�vG�q�����Tm�s��Slj�+�t�G�_�Hnm��CS3�٠��D
�M�%�g,��x��\���[(73��SyH�}(hI�^��Bj%g��'����8�D&n��������3��BQϖ����PW$�<	ա]��|ԳsO���u1�`p,Ns�n憄[!0��l�G$�b���l�����>d�J_+�	�fdЕ�u&e[��\�-���lµ������/�N&�&�y�:Q:k;�s�[�<CɓX��@���]r�!�!j
�!	�C#f�[�0鉠�����>ܥ�"���W`��zË��*�c-
��<��kG��N	�-��c���rP���_�c������d��>�������i�p�~�c��d{� ~��^�XU⟍H�k-u��1���݄��^�G8A�9��������i���9��%�ی/�
����s��Q�D���	�Z�v�QP��=��i��b��jʨ����r��$��#�Wr~�K���[�X2|UK?��kdȋ뻺{�(D��wx|��ġ�٪��=�J<d.5$�?�o���T�˯k�3�4�3Y�h*�gA�6�G� �]�4E����Y��.��w�b���;Xŧ4��(�[��j�:~�ZY��"��_�A�����FԄ�E/��RZŝu�ǹ��7�SE�Lf�S���ȭ�e��W�U����� ��W� b0����V��i��6�2x}���7�E�L�0���_b7�)}�L�/Q�u֠0h���g���̶�������=��]֑ڗ>��)]��rՌ�����~ߊ����[�x*��#	��}��XN���֕}����M]�NU�9X�XE����@�ؖP;���*��4��x�|�n&_�zh�ժ��c����b���5�tN%�
��~�BH(6���IŇ3��(���8W[Q���2���+���MB�݋3g ����lv��ΐI
�����|��� "7^Rf�#���A�(�e�g�X��L_'�	
�m�y�0�&��C^��Д�pKZq-WO���Jn���������B�>��<ե�a���^�D��ɭd]�(�w��a��WAs��]��s����[�����D'�F��}/(��vNx?�cb&[`g���Ï<�0�o��jD�n��u�x�C�P�>�鯽�҆1��^3@{��$�#���z´e4��񰑟x��
�%=��`R'�w�ި�����^���g��ia�l�q2��4r���j����Lk�_
d�����w2�+ؚ&뎶��*ܐe��J�nJn8�9j4���OI�њe֦�slb���=�g�L��1zJK��@����y|KT���4WAd� �S��%����*#}-��-�{j��R��y�C��V�y����e)��qn�8�Xz��I�*T@����Z�]#�͟���� BZ8��
�p�����`�]e�N���Wp�0٥ز��1��"�
���<W��,����L��Kv;�3Ԋ��=RW��H���ڛY���oi7�7��X
�6��޾�cluk����lgk�y�o��+r3��oS�j���ý�%b��` EE�Ӓ$!&�-x5����	ʖ�B�X-�������y%:�i�x�;�NS��͘j����?���|q�Ɛ�	ʴbF��'Yh�^!���j����z�r�(�z��<1t�ц��O�	�=�����~���P�I���q�:�=lK�vz���W(�&��L&�����M��լ�	-�u`r	�Z�O�<�١`��@<�՞���l���������>'��Q?��0�Z�E�Cݘ�R�N˫e��\�<[\����s)� '���Ł5wyi�o�6�a�Dܴ���^�v�cA.ۛ&�'R�S[�/���>@��
>ô�Oy>��d�~�\i]����7vH�#j7��J�)��W�����>�o�����RI��0�*��DG��G�K]�>#�����f}��&b�aW�,K(�� �Ԭ00��ՑMk`��&qZs��P�݇F���?p����"ہE����fi���57<���]:���P���T^������������ii�~������1�V>Ab/}!νZ� (�F�)�� �v��٦Z��d��9�t��0,r�CjV0�b\�Uf�h�t�-L�}�$���%?�%� ~�&]OMm7�P�bO{���[1��q�M����8W�6��[�RX���&ްx�����?W��q�D	Ol<��ܼy��i��� K�:�ќ;"ǋ�`�#:x�)E��N�D������RIi�v4��}�xگ�#�u�&����(���f-��go��RՊ1�wU?�=�S��(r���y�r5����"2\����\�l�4nF�W+������K�t���������dJ���&!�"���+�v�E�Tj��|�5�'&ȞE�%��%o�FcmW.s�_��R7� �����?�:�V��oEy������K���`����ۆ$`���F\΢׽��5�I�f���k�2@�ku�_oRk���f�QuCJ_+za5=��%IZ�����X�aD�#ã�e��֋����n���ٷ��<����zK�[���d��A��S��3����nϛ�b�C6�OQ�k�a�Fn�N:�"�{��N�q��ժ(�k��M�[Z���mn�xq���=��f�5������+/��t��r�1��* m�>1�u.V8mۡ��ɑ�Ua{���$�]��ɾݫ	k�tP%ų�Y&_H5ہQ)�w�dy<�" ��Mu�P�B�&�aL'k�����)|3]xW`gw�\��	��aO��n=`l��a��fl<7�1Ç�,�Sw���*�1̓~9���H/3ۦ�����i��D��c�z0��}�HѪsq�:��Z���N�;�8�R�οB��$f]~%�u�g�|�x�pVC��vJ� �1 뒣�������Ԧ�	껅"��7p<�F��@E��=���b����D�/r�HF��O��Ć��V'�#���t�^�맨�}�W'9�{l�߈<���>�d��1ǂ+��y8�tT)���a���ݭ��P�-yɁ���lS�M�p?�ćq���bP��o寜K�^����Ā�!X��C2�#`�$K��5�<��t`mC�Q^ub	�.�m�E ���>n���6%�3�o��i}ѹGdE�
I�������S����;�ؑ��$���o�8L�p��?&M�w�B��m�1��=���)�5�
;j#߮S��;���3{$A������LC��|�|w�i� �#%�ڄ�'���M��q�����Z�ަUqg�����rN�
�L�B:�u���#�*��<֣I�����'���$��0�����5�/�S/�^��׌^�Y0"��D�}����h#������_��U�������A�uҌ,�+�$��0;���l�z��3���z\�^���^��m����?��fŘx���$�o�������+����(�ϸC��U1��}ȩ�����V�mØ�g���S�Q�a�uo��^���w��"�ȡ�m�A�A�ڌ��[�k�I���l-���<-(��;����#�^��2�&�~��+!�yO��>~#JZ�<�3I���ݶ�$6.8�ct�g`25�t�\�T��ZF*��I�#���s~>���a-g�P�Đ+{���y�5y!�E�M�ڴ�S~��}w��ʞ0Eq�+���������}�� و ����?�$��XwK��p�����TG�/d[����'1߇%[Zs�N]�*Ct�axh  ����1#�X�@1��J臣.���^���(�QV8���p{T�V�N�w�š�8�R�~�����㯦�Ы�/%��h&�<|h��B��O���WMy���Koi�Q�F�l�00n2<9��}�ģ�x��p��wXG��|�	:k	��F�R�h�����G���ag�E�VU��L\���B	?�1x����Ŵ��CT�4�j��:b��6vg&}��k��*^���:��6`U~좄��_��D,~�O���pJNoY�����'�([�����7ktJߑDk���Q& Z{x�c�0Ͳ�'����*Ь	�ƥB,�Z��{z�e�۫����ϡvhof��ُ\�#c�DCD_f��x2�S��NJn6���x�Q���P|����FZS���w�A��A#�3��,/}�kp����d(�TAJ�o�:�����S�Z_/��o�:������&��m�ޡ�,*���:s�H��0|d�������2F�C��u��pu��zc��'��~�W>�͵��k��	��R���[e6�g�0�����,U8����e7�V~t&d�o�g����k��;�.	�k^k��
_�>��h�.�������:��a�++{��
'\������n�ǟ��Q�)���o��4�>NM��_4�I=r�+u��^AM�Exv�T�[Y��� le������]���y�Us�(�|�6j"�ݢ�$LU`F����am%��
�g�NdI�����@��3�>��'L5I�¡�W��J�5d��V�Y�O����K�M�h��jL��}?����{����2����9:{��_���[��W����ދ�iz��N���t��yu�-���y�8��~q6U��)`:d�`z�?�T�h��L����Cz]}﯏�ँ�K	y�
幬��#�Q���*$-�3y��w������F�_����p��(�cc^q�b1_B�
X��I&��Y%1��Q�!�A���wQux~�+Ǆ\��˃��cWV��ɉ�Г�;�?q�O��cʸ��5�D(�k�����>�E���˃��;���/���Y�<���*@D�6�J�X�[��L��?9���[:���ĥf�����m��\!�Ž&B2�
�%�!�9�a��l�@TnȠ�y�ud��u�OdOI3U�s6�I���Z V��~�hE�|�M9q.[�����X��-o���"�5�l������J-֠i� +�Th�Ɗ�O@<�j	��������uR�$�F,��fVY9QH�钏B��������Pe�iBTb:$�(O\P��;�H�?��rBN�a��A�]`S�����b+D�l�B*�7�)t{E��hiY�i����o�A�"�_��]�3���`{P�c����8;c2CQ'��C4��#hr��e{�(�}1R��)�?Hty�A7j�LiP)��r��Mk��� �3|��w4�e�$�i^t�+S���qM�q)���#��E*� �!��N(��
�d��בȑ<���̃�,��q�9��)V\���ӱ ��R��?���Q�R��J6��c���f�mUQ5�s#����	�IV�-	��O��t)*�uX��Q	�m����R� �h�����'�\���������������������ƅ�|Q�������	K~���7�U��Ս���B�
���$9���Ə͹��@w_�)~��ŭ�/Ǜ�-�N��!	�Q���WK{tJs�n,����~u�
}�(���jv�q�z/�ʩL1U�w20ye{�,F�0��&�U��׺���x�T����@>lY&L�t�6�����K���U=��:1��k��g�y�Y[���*j�ɧ^�<\4�U�Zo�����a��q����A<�l��jx���C��Ow7i�w9-spݙ�o����O�X���e�7�գ���4�B�#���*�O������n�y�'C�Bu������� +���k���e+mW��WI4kq�֯s��gЛ�f
�7 ��i�#Y����Z?�Ya	�/��ع(̇�S���n���jj�$�N�������Q���ER�AC�uE���
z�u��Qw8�-�(�Q���*u��$6��4�;uUf���ێ��!8�i���+ۢy����)�B���.��K;р|Q�;D�m2��r�tP��u��M��3�C�̖�?���_���ϭ鿊�݋�B�P�ˇ�����N��	���f<���Q<��i����K���%�;��N5�H�["�5\�l7�ŴeU,{	�.w�t�A}#D�M�Brv�xX���E*�~s���RP�z���T��աG����a{��^3�����:����!�2Ծ�E1Ӌ�P��,/�_�\w�c���sE��lL��7mt~����)#�q��q��{%H~{{a@'6p!�:8��.���BO�.`�Yn���t�x֧�@����xX�������Ԓ��H��y�?�{�,DW���t��\���G�W�N�(�y�2j�n���Es1�j�V3QHy���R�X�o+�'t���&�(��t�#%�5�'�i�a��uȎC� �-Yw1���q+�P��O�1y������~
~���V�Ǝ�)���Ԅ`"X��d�5h�a�t?rQ�zn���X����zs{+�벊G��=��Pp-�;���绞�T�[��ʕs��!�X�FS"�]�wM} ��rc8Ư������[����m11���n�0�1��d#��G:/6}(���4�7�K_�)Lŧ�藭�Z�U��/@_$��Mw0���^P`�4�0��Ӡ?�y����;Ќ��9
�8���~���+�L��@>7��ġ�������`�<��h����#.�0r/uz��,eF�e�j��w��=k�m������(������6�)�����8����R��I�39����T>�.-����wT�-f$�t/mDY}�P��}f� �2�kib,�i�WL�I�ʍ���l
�߹C�����̪�d��ʵ���JC�f��Ӑ�V5����!A�d��C�Z�ϧ�K�蠹:��v�{z�?�9'�5�d���nG����RF����=��r+2��ْ�x"���E�Q��'Lwt�`��������~Y��6/5�:����e��A˘����Sꌗ�é��嚖���[�S�f�	����t��&E�y�U�[�h�)6Q*�ݢ�M�Q���7g���c���\�A����/�.6p꺎���wنKpZe�4�4�Һ�C[��,��Ye��Q���ɲ�s�Bt	��}N�:��F�V�Zؗ���['TS?٦����'{�k��"n�:�{���O�^�G1s�b�96ԁ�0-��9��jŔ����&�@Q�Y�	Xh;�nV�ׯ����s���O����j/������z��
�����(�����������"PW?h�X�h#
ؐI6Xq�%}[S2��^�04.��[ڏ�?�@#��)KVGtx2uּ�9���Cl%4�9+'����������	�:�'�ΑA�ߖ�����ۨdY�jiN* �.�ܟ� 	�5�D�2�Ƴ�xĴ��#+���yf��{�
NV��4�9/>�������܎Ќ�=vϥ R%��%�����C���<�\/M�M&P	]�~���r~1�b��+�Ar�����~��1���6cHL���1,�eg>�n�Go��JE�g��v��y89���}��I��HY�Kµt��+�N\i����,|�����Qi0�m�J�%՘�c�����]/y�v���]G�}��:V��V��ʉz�!*GWA�:�j�t������Lg��Ҽ�|����g�˥�-t�<!]o����<�{����sKl�?�.����� V�g����z��|8E����SW���]���?�� ΆB���C�0�39�87G��[J���3N���z�D"G���<~��>}P
-y���0����LS�P��t�^	�+��F9�p�{��Mi�4���h�S�n!���fm�ژ�0���Q��J
n��l�f�$������j۹wO��^���
��9;--�ѦB�%0?��l����!�
EC>�8|g�����1+4|��w����
�	�i Ut偃=R�C��'�5�73�a�\��=�ZYx��n;�s���=��|I�+[�f����AI��_ۥqI�ٲ�S�P����R�b�R2ұ+Y�vݝ���
�&����L�s�ș�a��H6%n�g��Ô����9���.��V��~8�4hLh��%'�lǟ�	��$ʌ!#�	���%���:�D�/�f��9��F�Un2�A2����8�h@ �C��nf{��tV���r�a/�I�{]�sh5��(�jmcKc���a����C��K���5�~�:�@��a��E�j����Jż�E.C�<���d6)�ޱ9�9���˘��\��Қy=-8q?<cm>�"i��ݦ��a�T�\����B�(���	����St�%g�%�`�'�J_�Ra��g�0��ňy+��6�A=-�B#ɒ�+��J�F�Q!�!�v##0�c��ȿ���� �k��>�MXU��r<�O�`����������ڲy]R�x4��=V]a��4Me��h���"���M��`���5d����5hľe�H��>��&\"�9�E��[>�;�VX�p�~��C��%ĸ�h�ֆ�v]�2���kU�uQ�|���RB��7���J�J�Q�鴅6����~4�Ff<�d%�j-�`�w�bo��H?U�Q��XF�6��:	GНQ�)������T�y�#����g���t?��؜�jwx�m���&�h�m�s�UXw3/:�a��(�t�ŵ_r�����T�^�����"�mJ [�W�QP���.���<��A��|"YZ�4.�9���K=��n|�m��UAu[tZ`�{�׃_�G��Q�o+�=��*T(�1Ӓ5�-/������8u���ɆXM��؉���
��{�������(�X٥��� �bE�Y�9L�Af�$��;L/f�n,�_��K�U�2�]���4��u���IB&����Tm8�o!�u��=�y�E`?JJA��)a]�eŠg�����E�����c��u�)�,6W����l����Q>��_�?���n8ըs"�*��̬�S�F��$���Q��h�M.�\����5OL$´��<�jr5/u�~Q���>h�JS�s!G��6�QHq��
f��"(�;uZX#����/`Y%�����=�������EL��+�s�U����y?���R��~�c�>w��e)��"j�e�*[<�@�)���
�D�.v��~y0Q{r��Q�L=FlU�N|��������`jse�yt��o�(s@kԐ������ͮ];�o"�eh�3��"$�uO�*q0�2i�Ov�4*���0��?I	ߪ�\\�H!Xž�I'�`�p�������*#K;9�Ƣ*���J����kIJ�wf��r:��b?3?��!�fF):�}�k��m����Ol����P��7���/T6�h�')\=�EZ4��@^�d�8�� ��2\RN;>�#���A� �H�__����3<��^5�"�{��t&�`�2��Z� Qg�zFH�-�hS�MY���S)�oB>��9m�&Ɖ��C�jC�2jS0��/�שT�f��V+��Y,*y+k�3�*Y�������إ�����f 
��-��	ϲ��fr$
=J���S2@LF���ߪ�c�=͊r�;��&�;�x�ϗM*Y�g�PJ���7�/����
�ë��&����jv.��bƷL�$��5g���F�?��<���=4 ����^��C&�jV�r�غ�HtN�_^|��D�;�/�h�I�i~�/vl���{p %�:�a��bb��s*�Q���:��_���dϪue�4�T��i��e�/�%)�?�揠�$���NHuJ�Eg�������ߩ@������~Y�cu�:MkFK�z��j]Vǥv��^���ݔ��AO���%�2$䄜���;�;�7�%lE��+�Br����cɕ5h�R�8.}�U�A�B�)�:��1z*�^ӣ�!�BqW�4ADX�l6I(dR9<*:W�e��}��7���fm�ćKP���6�(ڷ���f�Kd�JQݛRc�ro��5��QBV���	�.ie�1���W6�9PQ�|���v����೜����"�A@YI̱��7�u�C��A�`�'a/q|
��n^	0��$w��3|�xps;ԟ�r�?b��s��(����3����kr-X��x�2�鬿�Rb���~{4�.(#0 �O�<�Q�R��C�#+m;��%ՀtH�^���l�~a!�^�ai�u�Ty�f����8O������5�񄔥c�;|�nb=�V8M�#���	�B��w]0h��⵫�&�K��JX�����S�f5���%��ޥ즷A�ά���j���O��|��r���GJo{i�e�Κ��>LQ(E�`�u3n�MG����!�F���G(�/;�5ZR�1J��A��K���O�s�����g����\?d���XK��<9x'aMU����H�Ɲ�
�\�w���'�pM���t��0����8���e#b�N�h'�/s����󇇬���cP	^��M���8�W*�uŪW�!x_|Ee8�qy^Wp�k��rv�o��?==M�H����W�Le���?wgM�y�N��<��ه�T���xg�&� �>��� �+���82d�I��)������0�Y�Z�<�.���NSx�1�a&���*'u��Lb^��-GY&=l��;2���Ǆ��czR`�/HNɑ\��Y6�r�هz<�XX��rֈ\nvs>�H#���|NP�n�����VtF�qV;ؤ�.6�&�Y����͖��%����L�b�l�`4UӴ5�L���O�����/�3y�鲟{'��~g�0|�W"C������vj�l�$1B��<,�=�S��O_�Hew<�/p~w����J?�G~>�#����K��L���}01���D�y���������
z��]$Q��#fY�
r6|�YҨC�	������T�wrJ�͢�̙�l�hy�I���5>-�9#�Ҕ�+�uTZ���,'����ӆy��bL���"�v\�W�K_�1���^�P��@�Ie�{�8�xF03uo�pOvF�x�y�
�4��=�����Rc$G�!3E�j����?�C����b���"��7w��X��u	���60�e���4�-������74�������c4�|���=�8>�E��哗�������=L��IX�~6�]��6]���g[/-�;L�gl���+-��X�TԟGz9&��J�|F��*��nǶ�|�Kܙ�2S}��y��s�L%dlB�tT�\���B��L����x��P6��*�� �
�	0 |%Z��c|��?��3�����3���7�IΚD�~�1���3���ӑV�q��w��;���{8��ESG�۹�U��� Ԁ��5)�p�ʲ(�՜�;�IZ���[2WWy@�8؄~�ǜrE�ϗ<���=%(]#Ao��>����t�E+�����.�8a�.͖������i��Ik�|,@�eE~*�t>�[T,ƹ%����i<,���}��;n�S��3ǵ�1l`�
�f��\'�~��)&+��@��nsd�F��#DM[�!��Qf����g�t��������mv$�a�2��_��p!K�K��k�@C�G��v��,g��k�g�ADH�J@H���ϋ��T�ӭ������=@ϸ�2|i��M̟2�Q��0ʫp��t�o&|^�MR~�?*�����I
P
	R���fr$�0Wk�����M
!ń����(Eؚi�24l���zt�I�UF���z��a���]�s���}_�8�+���I �#m��H���}\h&[�=�.�F%����/��U?�9���.]$��k�c�O�خ�fkg<c��&'m-$E)�q(��TV.������}*��'O1F2ӛ�3�J�?˧X�;]A��¨�����(�Gx���*�!����b;6�k�f���q�ށ� ����\Аpk�G��"�=�v�딢�n)aH���q�����[���.�|��
�' ]+\��#t�#J
��(N�rI�����s��C��) ���[���<�tؾ�����L^ ���6.�HK��r����	�)��E:	'���K��n�:
�4,9ڸ�g��I����2�aT�~/�\3DJ0Qo���A��~�.�%�ɳI�U�"�`��D@x��UzV�ѻ��m	�Q��l\#y�=]��;9�t��ך
)�c6]�F�e>Oj\x4��M�fR�ylzf�W{�>l#�.6-}�{�A�k97g�7� J�LG	]�6��6�.�S��b?��G��1�e��XUQm"��Rjm7�����f��^��,*D��ˠNmPS�Fއ�^�?��|�l WS>���wDw�QQ]����flp����D�`�I�ΤA�#�I&Ϯ����d��9[8UT�A����A��n)z��e_X���q�5%D�Բ�:�9�E�KD��7�b��	
�-�I4����6�s��+�e�\�Qi���t7����)�i1���&�apB��u ��tjGS��DCdt���/>�UO<�	�|�v����:F��0g������^/?���L9*�n`C��g�=D���v�_�z�u��
��8�'p-�y<K��Cׂj�.���R�q��@�;*���C�%���B�>�4;�8�~}"����+�K�vp���Re���1�.6,hވ��F�NN�_/O\0h�]�Ёg��>d��G�O�"3e�@��8i	W���W�M���`NZ��s���M�*t����X��<^�I�8}���Ř���Ȇ ܏��uX��)u�2�T�o�I�X���:�;2�6]z;nL�F�+z����fPd�1do�*��_W�lp^�g���^�r*&�<�7`=ǦBqT!ե'ta����ڶ�2+�\Ӧ$� F��� �C�B{�;kd�ЭrzV�T�[C ��Eڃ��~j��B���J���1q�qHz�^E�n����?��qUw0���8�2���uP�T J�^�������0��󡅽t���H6�kv��~}�|d"D|�:R����c�����mw��{~ɸR#}���.�.]���X����=��\od��P��D9�A�U�o���/` �[@5��~GA������@:,�2뤢Q�b'��J�����{�y��2��Ⴀ��خoMv!gx�����S��	�+�rBxN���9�@��<��=-�=l��%������5IXT��xI&햆�(�/$��w�}��P��8���tԂ�fEL,pE�Ȳ=��z��7�K�,<�3����_����jr%���ڧ5�Ť��԰Ӆֵ��\6��عBʡ��b���c��T`̵d�}z%b����V��U*�cRJYV��|Τm:�D3tmG�6O ]-Up �}9*�b�������Br��Fs��^b���>�Yp����4D]9�r���P.�p�-�3g�O�%$�� �*h^#�dJ�P���x)��G�?s�w�W���:f����v��*���<|�
Oo�-�J����}�|޴�9��۵z�5���E��kŖ�0�m�-�ri2��%�g���aM"��$��=��Ok a�)���1���Ā����3�g�D���]h�0&��گ�Z|����-K� ��i� ���s�]��ȫl����;�� J��������)��
/��u���)� ѕf6������r�<�� ��D�!��/�o��O����8n�����4kSI��{q����z=� G�N�F����Gp�BҞ|39Ce��NWVi@ʧ���	���SS��a(H��=ޯ[��2�)���&�W���kE�=ߠ�2�(o;^�}0��&r:�[۔Oʞ�'�wL���u3���-j%�-m9YL2��&�Tߟ6�[�u�vUڃ��+_�D8�(d�K��.�l�ys��dEk��~lfț��(%[��u���-h�J��rlL7�˨�Z��vcG���b�D>��e=��J��I���Ei&u�I��_��Σ�������
/���;;���:�yq
z��ٳy^R$jZ�!���Fv�k
��;]���oX����K0��ւ�`�*���CL��t�v=o�E ���G�\bF��Y�>U�n��1�%�E���f��y�ʮ��e�.�AK)�:��j`<3hLb���d�$Sqמ)�/f���'�ZP��47�I���}N��l�ѐ}��A�̶f�����%�r�t�aEp���e7i��d��&f�C�PC8dU�F}���ATU�uWT|Chɂ曯m��4��KA�>b�hB�#�����8�{�r����4�b����|���􁕋ej�<�?�*ߒF��(�C*5�m���T�V��$Mv�2�:±`����01vu��MVͥ9��O�Ս� �F�a*M��٩\���_v�|GȊ���>765�D��*/�#�t��g,i��m�)�l��	Q;9��+	�75��*�х��,��3?b�cAk�u�V矛'�2��t1�,?��֫
}�~�(K@~b��(6�X�LD�䫃�~��,L�	�[�o�'}#�%���ᵐ�\�*��X�ޞn�w�%���t�=i���v����<y1m���Ȓ�Cv�P8
.����v�D�	"[�,S�l��r%W�	�a�2#��p�;ª8�W�ޛ�Ta��ƭ�&���(���������ё�S;��,�: cӚ�G�K�T�����v��.��!H �4�?h^�F��a{9�2Gg�9Ts�<P�T`�f�����e�toVEf���N���<�z�%�2�_��O7-�$����T3��"������ܡ�1ĵ;�u��=9b4��$����a�;�kr��$�U��E�n���ltS�M2�n����CI�=칤թ���G]n���-y�>�"�fy���P���L˥��w� ���Qw�$�׈���C����FZ��:���@�T�1�,�eYݕi�_�u�u�M���tR��lv��!�>�G
;mmG�����=ƮT�B�����?MH�oH4l�4�?��`�q�ض�[�V��c$��8o"��yU�'���rG �*��w�%vò��޿8	�s
�b�wp9�`�{6�=Be�eQzūk��űi���Q�+�D�
Z�5r`n�j��-~���ҋi\�B��V8z���\[t�6y��A�b���͎�n�t��b٬Ok��d(^GN�z���̮�վ��]6��:�8�1�����y��
�j-��r��B��?��K'��Q���#�F����=��%��0��rW�LS�$�W$��s{j�{�|�=0�6T:Xr�!��E̼e�x'�C�\J�a�J+�7l�N��f��7����c�)�I��i��j�>�t�~�aY\)#D���
ѱ�YA�D����I<=.�^L��)@
�6TL�A��^�����v�~�ŉE?�r�"�b$���~-[I��蘒�dj6�`�lz�E�8��܊�Kd�R�4<|l-׵@�ڎL�I7��M?+��ϙ�rgWyU��OC<��N�6�d&�_M�_U#�t�fa���""�6#���x��IF� �(��Z��F{cD S����f��%��֮+jçUIs�%(���Xb�o^h�>Ph ,�q���x�8.B��N)��,�}��$z��bɋS��#ߺdɚ	2_�!�x��fC���g��&)ߦ3a�����%LՏ{7P(kf٪��@�I`�C8�]��L�>PO*�����τ�$fp�$+��-��ŕ�uq����T��^�Lohf7�"���xz����+�Z�Өo���S�^S��o&IA�O��3�"�žYO��4�D+�\�Ǘp,���듍+Ur������|�!+��T�T@��5�6:i`:�'x��4�V!-���j4�VF"��F�3ZC�|�|IXFi�94#w>�.�xd@V��B�Zl'Ee��>��m�����5(�f9�@�|�t/����A�^�B�8�txV���5u�y��Hj׷�@`��<�7U��Ly����#��?�
M�8��{����s�Vʟ�g�f�Z�����Ȫ�����3/������$��2a2Fc����n�{��֏�|w�謏ݢ���)��+����f���Y;
�;�Ϲ�A��n~��Y�S��Yں�M�j'o_���a�=-���~6���9N�)�5� ��O#D���@n`�c�<��+M��#����(�׈�ӏ�8|��u��u����vqC��?�j�c0��}���N3�y�t;@H2�����	��	��!m���Ow	yٮF����>�G����(m��дz�B☺{�I!������!.����H�8�dZ�`c9�[ GC��!��P�O`��D�ᅹHկl���7���I�@1�|T��b!o����t̘�M�P��E��jU��.=r�;+�}N��'Mq.j=���S�fN�v�^*\n�@��jM���I-�Q!�Ҕo��/��� ��ԅ�kp���E�T��B�*�)QE�� Oѵ{�x������A���3� }�b�V��Ƹ���F��	NL����Y�Sk�����=� �:a־D9�w�DV5v}�l����u�D}K_�*p����K ��/��U)�Mˡ�	P���2��a��/��F�o!������~*�����y��� N�$m���SѢ�K燘������Z���.�=��0ڶ����m{��Q������%7�4��L�A�� l���"I��C9`��E#��'It�
�S�ǲI�>y�5
Izp'I-�����G��j�E��x��]t�Ã:���T�|�!��R��Z�َ��9}Eo� ?��k\q�y����6���~�@���Y�'j�h��^��j!������w�|x���JacR��Fp(+b,��c)�%���p~��N�<7���r!�7��~I���<�F�C��Y�\0:�Թ�mK�4�-��2'@��0u�4$�Y-s>U<W�0�1�wO��`���,2���Zo![QX.w�A����]�x|y>���o;Ŝ��~x$�]�v3o��~T�&����_XG�R:����'�<��0�(�t�/U����������)���Wh�3���(���`u�N��W+��^�uI�[ef��R�]ǆ����f��񄑇ZL#tz��6`�&85�^�]3��K
c�K���1�^�m���BE�<�,���\���N\;��x�jW���h#�(��dݰY�Ap����}�����2͞���={�eʰj�9&���X�8k܋��=���j���>��f�qo�xW�f�?XSX2_�0h�礻^2I	}/���RC|[i�ۭZE���d?:q��V�F�A�(�ˇ�f;�u�����:��gN�pGA�K�I=k�����`�Zfo��xr��	�-2���P���v6��<3T,��T�W;�Ɂ^=��h�����lBXՍ!���/�h �	�_��[k��t�~�O����X��Ҁ	) L�����������F
���N��	GO���t��:�.1���3t���gk���"�=���Ɛ��zaao��O\����,����OU,
P��hD����c���yKH�k w���U�ZV��fUQ~
M��t�f���U�\)vA���h��CnL�$|r��X���s�k�Ƶi�K�{�0n�7F��6>zǗ�YjfBvW�!�9H4hZ�>RϮ��������Ƿ��,�FG(��`�;�9\��p�j���OVX�����9��d��� �����kR�J�m����@
��y�$ \�{��KC�!Gd������`�0V1A���0�g[T�%�f#�Pj'v�A¹��N���{.JA�:&��C�d=P,��ڼ�����o�v>����"����4�0��������^<���0Y��M;xo����k.=B�ǒ<=k�v�}y�;C�	�49i�����a�T�����#7%�+�M��*�W�$�z��(\ea��7B��~~�A�_Y��הA��p�h�b? � ��<{i�m�W��-�Y�*��5�Qu�Q�����6ǤT��.m�x,�o�_�	Su	�~���
����K���|���^�9^lbe��A����*{uo��x=S ��@�����3�l�z�1�ei�NsgL�ϣ2�K�)�}����]���Y�m{���Rً	����d`�"�	�^��q��x��R����0Q4RUq�9M�Mo�?����TE�4�H��%tm"C�}����6�iJ��� >~�z3�/Tvҋ�h���L���og p�I�9qVy��d;��1e���S���L �}:����:lJ�KR�8O⎰2�k���R���p�vB[�6~�o�ڏ?|iqܲt�r
8�T�nYO�\$\ؿ�Ɉ@O�r��|��|�>-"G��Y�
z^8v4K���������h3f)_�6��RRќc��=��wlnYcQ���Y�RB��RR�t�*�F���p���8���귌Y��t�d���$z�ya�iH)�`~�,)��NN�W_�������+$����M��z��ژ��[�*��p�肥S�s��qBs}�O���Kz�h�X�U"K��b���:{��E��������rk3a��+��x�ƁzP��>��FaԹ�؆

T���7p0�
T��޵$d 蹁 �Z�a֌47r�QL<��'��F(�I4�ka0���L�r�=�t#��5+������pRv~�x>���������`P=�&6���R��	LxѸ7n���8�	�lԶ�X~[i��9����1�y�'s!�/�Y���/g�\C��(�k�����QU�;�8Y���Ee�E��O�р�>��cS���%��օD�j�/�=x�n1��ѓ���a���Q���4�	`&uo&Ai�$���h4^K'��(q�$Ӫ$X\v��"�#�aN&��~�;�q�����I�&�{g��ȗ��`|� ̎����n}�X�U%�y�B��2����<���4Kh��-��?���������:3��C�R��� vI�݌w�mJ��Ib�,4P]�X�?�� ec9%��K�)�Vo�iX߆�3a�5C׈�`��t�<T�y,����7�3��b���R����2�KD��'|�M�\ɕ����_��4��1f�ͅ2�= .v)jP�NQ����2�<��X�B	����*s���Q`�]�l�	/��vMO�c���q̀�(�va#w��z\v�>��X1b!�neW�R 9ƣ�(@'7�ARv�)A�$H�9��j>�8U͚	8vܫ��d��M���f�
�50:G��fHB��"��P��r����m.��`��8A�s,Lrj�t���H$�)P���2/��g)ꄏ⬅0 <�Ԛ�`$��c��b����Ep����%W"��%�r!?Q����!)@�߭���Qj���G(\�7�F��g$Q]��:+2����q�Mo��7�ƅl|8TY�����0��F�q�2�W�ڕ�I��Z����)Q�+k`��+
�y��G�~4춭� ���޹lґ�K�8��Z+�_��?�˛E���gp
D��wВ"���R�y%�"I̷�A-�߼���O�<1i��0���D� �$Ӿ���R����i<ʤV����W�'�g�ˠd�ۥ�D!/k9C`�9�d��q.�tV��UÖ���6hR�bFf�	2e_��Mg�5>�d
iS��xn�{�Z��Kf8,��3�L.��8�lK�}��j�D�,/W'6l��g�]Z6�?��$ʖ�(�Y����>��jn��6?��ט>S��a�
��R��S�|>�;<�$w�>FgK��T�KV)k��d�祐���Q����c>��\A�eB�כ_��(��GM� ��Hو��p�� ��'��L��s���E)t��-?Q<LÈ�RY|���	�O��a5����R�#�M���5ǜ2j@@5x*[e�!������j��2�W|l���5�'�d�
�"p%/c_��z��:�����ɚ|g��ε�w�>C��Ao`�r�7�	�o?[,��o#��z?,wB5"�����.5��g9U%���3�+�q�o�?.�}�V.w'�t6������TI8~� �[�}�X�g{���gaZ�����#���9K�ˎ������ P��XU|��W1S` 8�D5<\?P�z����n5E �=�̪�-���k {e.��E>��?@T�)�2)p-�F`Ѡ�6+k\uC��q�z���'��&9�*�r%12�\��F�Ӑ��*�o����}.��V�cP�lb�����B��r37H�غ&,`d����xv�6 �Y�w̉,��ФN}�@����i���.�U�C��<�8/0F�W���:����%��_w����Ê���[�2	�H�6���A���G�@x�Q�a{�/��!�ST�ú3�A�
v��c���b�jo����d�*��f�!)y��7/��f}�Z��mK	8�D/k��&�`���4����O�M*��I}�����&+60ϵ2줹�o�gVsU���@��I�p�v]QF�֬���}@�Hzt���-��R�)E���g�6d)��<�+����z���Q��'J�k2�a��o���^�5���y���IV ��(檉#�u�LT�E[$P���k̳�e�%���lH�oMw���g���=��f�y:dP\� %L�fK�N]� Tr��P�[;���	1��E壾$R���u��@�H��Bw�4��T׸�+�PY �=�b�������_,Q��2�1,�6�e�8 ��،>��]b��_VQdX�m�Ó��?��KY;˦s�'F�G�����T��\ˮ��$�����_^&����(�$eR�i���SJ������|����8�Rd��Uݫka�2���ґů��T�2�
q��6�/��{7�:%�m��N��Y��g�a����)nԆ%��}GB�0�")���:��=2��$,�Jxi�a��y��R�.��X���Z��z�hB�S8�쨭�m�ؑ�جQ�H��=4�"qK�/�9��2$��5e�'y�}W���Eɬ�V�H�~�LS�:`����c��}��3�������Y`ثj	"��Y���At�i$�����x�(X :	2ikX�!)��E(H)2'ƞ'`}�S����e�¬�U���E����v��WN�˥�,�۱(�RZck��0nףr�E�y*�4
G�k-�C���b�В��53fgl���x	k�ވ���<�r�?1Ļ��PC#�<�Г�(�
��|V�z9M����Ŀ�H$������	���zc�zB:3Q�v����|ȣ%P��na�i���������9�'W ��/�'���i �d�&�÷z�b��H^�=��dBl�-���Bu��\���E�<��ӚT?�0����rx�~<`�j(�7m��m^o�&�%��9�;i���=�){�j�^�Dߟ��'*ّ<C��9��[ �B~<��T/�|B�*���z�m�Gj��e�� iL�@���e�CÛ&��x!=Z-Xw�Y1Hz=S�=��6tAA�"�����y��L�3e�}��K���ц��-3'�9V/�� �I�َ�U���
"��0��.\va=��̍K*>�p!o��\�H]-n�̾6[�1J{F�%�1��$Џ�E�e.����l�/�!�0ݝ��������6�ل^�����O�^��MKv�@|ySɣGq��<���@e>Wc-q�Q�/����9wS�OZ7Yi��D�m���>��z#��z/���B��|+k��m�Տ�_��d��J 7d�i�TU�L��vo�o���Q�-�t���#۴T�>�f��U�쇡n��6��P�Xa�Y15�EI��W�C{P\�s�<(�����!K���o�}�308&4;�����[��gb6��#�C�Gb�Bvy�4�Ќ�+�1ɂ��:����<��1�!���׌ӗϲG�l�2R����L��0�tQ�k���}e3@����H���#�O�	Ő�F��k$�iw,o�B���$4,~���w#�҈�"�&�:�뎝. ���|p�����ۤ1ԗ�(Ȁ"�W[$��i�����r# �r� qA�1���i$ɨ��<���w9�!�|��UBOի����3fk[%���],�23ه<����U�!2-ܡ���iO*��^R�dǟܛ�5W�s�%W2	p���u����s�a�r�F�*#EXg�"{���/V�kQ� ��u�K���D���k�Oi��O��R'F�|�����.�U�rJE==�Ɣ�����.IP����zHY1�K�H�c���ßħ�SL�u��#����6�p�`3������|� ��!QY�'�d��-�s�߹�����X�D�/��e(� �=�@+�a�Ø1P����6V��O�Uy	�J͗H��BC��6!�1��7�?��Fie��p��Jr�B԰��kW�p�K���0�4����:v���.��j�Yy�p���z�[ 0!�&�r�_���p��NeTqFL��N:���XkD!S�{�[T�x�Q�χ��*�����p�'� P�'����*�DY��I�hLe�4�Lv�El7�L;�2��U����}j6���|gEz��O����N��*���/������)_r������>���@�h�m��Z��8ހrro|DH��	( �]�u�����!|�_��0��L�8��<��7t�P`?���<�":�A��H{9����L�8�]q�ڬ���ٻpR��TW���JB��M�>�<�[41c�^�A��߬��b�᮳�`}f��^�Jr��8?�9�"ԫ� :���&9wB��RMK�h	�h�4���8.�f\ �[?j�p�V
��'���n������wˮ��/�x����oG�0[� ��x�;{Ԇ{���-��v�<Ti�h����A��O2�-��Tf��=�s	�?*���[��s�.&�Y��1�p��hu7y��w��Ɗ#S�MZ=\6���r`7�V�`f6B"ڜB�v���~;�T���6=ގ�tf�uw��)Z�]���Y���B�����)�q��%C$#<�W	n'���
�P��x�:�o�=�j7}^�'W}<0�Ayb��;(V4���"N��7�=�2$�B�s���O�Y?jӾ����;�1v	1g��85�)�v��J0��h�p�A>���x�5��l�r�]F/�Xj��A���ӲRq�(k�ʰr��RI�a��� �.Q��k(���^�!ڪއ!��2�c��\}N�����Y<p@[���$��k�cF���4L��,�K	��Txz��䶜��T�@�C���>a��!��v��TG�mw	o2vJp}�X.q����AR�Gs#߰OQހ�H�;ߋ�c�z�#�vTo6�Ϻ���m����;��[H�i��+��%|~��W��({��1��2A%bqד����h��$���H�҅�O�4��˛�A�ѲΪ�B��/x��֊&��RV���m�Oz�)ǌ�w2��_G)�9p1����r-��Y����h���ҙ��+����3� 5�R�����-����@����4O����A=PS{�3U�s�.a�(����~�P�0��m��V�![ǁ]�I���U�����\�Ԋ}���#��Y>/���t�-�
S��}��;G)�����@��(9�qr����Pn�o�Z��]f�^�<
"�d� P���T�3nP����am�-�
��06@mh�5 ��!�{��N����)���eı^��)p�.�p!�y����@�H�� ��䉪��(D�ib[G�?%�l�
1za����
߱Q��y�D�8B�Ia�4k���
��o�	'�>�	��P�Pn )?��~qg�)��2�}��!s_Q|͆�7{�c��ڄ���3[����vM���qy�9`9{q�����T�%ֲLzl ��1����oR���dl"Έ��y��/���0BU��+�M$e%VL��� �3[��1�O��[H�y�$���.���ʅ�1��X���&A(�n��oU�Ov
�׏������w�!��nh�0;qGs��s��Ap�t������FW"3�:���H��l�p�A�-�s�#ZԱ�*ң`�*��M���T����O�Wy�Vӻs�q�"ޖ��oh����W�/8����I+��j�ƅ>cCא�Fd��
φe��_A���X��3�sXP�}����ͅ�׉Sc���s淂j{�7�S��"�P%�]A���l��v���O��^U���y�׻%��T�TYl߲P�L���̸wV� �m�����Fab3�}�]B:{\�"�x�mdk��ION֔�hD�9`�X�����K��T�}ՄJc��n�{)�ᮮ� �ҁ��~7���[�;�dX���ʧ��R#��?`V�S�w�'��V�C�縖��\�&Li���F"Ȓ�oZ�TU�����>DN�#�W2�Gq;�Id	�Q��a�-D�P��I�3=��b�=#ԋ@��p���F�+��n����4�5p��pѬT�Um���_������_)��j����P�N!���d@����1�o�^!�g��ET&R�A��nˮ�)�6;1� ��7������e[ 寀]��38��A^=�p08��^�N;�E.e>g��>��A�p��(e���eNp��^����E���oC��i������e�6{"U���wM�
5�Y	�	'-8V�EE�3�����{���9�hqQ�Fl��W­��Ҕ}c�~�]S��|e!*i^JݙB{e�d��m/��ӌ#�7YR&l3By�צeL�c����&���!��a����Lj�@J"��E�d�1�+�Mry�=�Y�R��+JCz��MyQ����qp+-����2?�YyI��(g���K�e�P���,��3�W^H�빭ؑ#_҈�7�H9�ZW1n(;:#���,��7_ ��@~Fo�¥�}�n��@ OC���К��H|=�H��+�r�ɴ+�ү�	ģ;FD�\w/�8�E���x�iW��p�Lv�o�j]�SF�5�?F�I�&	�����F��LJGs�r�"l�rd�B[3d#�_�$�W��������h�,�K8����I�@�(Gv��?�3��;T���?r+�H�EX�����-K��h�w�se�1� <���t�ﮙ�T�����´���im��_a��g��u��pK��Q*���Ti�"���;���s鋆�";�o�m�S�Yt��A����B��7�ŉ�]���41ًlh�r5]e����	�!���=���_�����j��kotQ�9L�����ɦj���H�>�_�,>����yL��.f.F����P>g�<f:�صCY@2ۂB���4����ƀ������X��.�K��Y���
 2m�u�� �n��̧ l�8OА=�<��`��u��Pq%�UU���>��;����f���D��0��F%JR�'XC"p�H�f����r�n�Z1w���-�&�sz%��E�j�͐���w��}^�?`p�c�T?'xg-=(3O\z� T;p�iV�M&D����
��(w�u�h��*��c��ς�k�����v\��t3�NW��L+)8;<i;).'�י�oX��W�+y��K�i:��7���:Aa���7nƏ��Y�)
��B��9!���
�������${2
�gD2�C,OJ���V�P�^�ث>-�N҉6<���3���a���ZI>��@T�������8���l1'_�,`�-�X����U���T���jTR�#���' ^$R�JS��lɺ�g�4�}hvvs�U�{|O���
�'I���+��Vr�B,'�.�? g�f�[2��r)h m\�a[c�z	����!�g�x�!2XL�(�����^/*F�qF�4��]�M=R��Y��QnE�a�cQB�?Λf���hN��O$�%Ÿ �aL���j�t�\�V��Ț���E �J�Y��9��P/X�j��=P�T�`��f�g&?������ҡk$�H�J|�D���능������y�9�4�,/CH�3K"�`p9U�RG	>�t`���a�[0]cH�6S��ˑk�7o:���jD�ҼF�g�˵*�K{�����n+�F�>��vƤi��!�Nv1x�}8���-��GH���R�X�☴�ތ�LJ�f����������'IK�DEE�98�a�D�	�Df>w�����>��lik����Ә�%��A�yB�ٳ�=��IN�ۨ���v�W�h�YW�$n��{��)�5Ƿ��jNj��Iڃ[�sol7S�&���GJW(/V�T��3a��`)�N@���ln����[X90ӽ�?A�X���k��8`����'� �������iEܲ�̩m�3�TS�t�n<�2RN�
�w�����#����/���Ԏ�1ϫӽӁ2�<.<�$�|т6�+��@�A?��,�ۈ�?�Z�ђO�=��wZ���BD�8Hߜ�[7�q�W�#�T�|J! gBРP�rΡ����i�-�'����x/l�������Os+`R>����)�z൞��Я쯒�n�:�ǀ�-���VL��0RY�Ԇ������8�l
0y��/<%�#�U�}}����:��)W5��ԥ�� �bv+�E��d{�/����0Q�m�e�\X�[��ה�����z�͖pM(,�4�\ �L5(�1�C§LU��� �r�ہ&��lq��y��Y"�v/�����P ��ɡ����C4D2���BD�0B�[GH/�Œ�s�h�@oMm(�'���
��Lxtc1I�4�y�_��Cw^� ���H7vpEQ3�P���{�_�&D�=�E[�P�|�L���e�{ �=�&(�����o��4�B%BSH���h�E�-����w��a���0q|&��(�kD��H��L\�#}��'<WMr��>��~�h$ ������u����e;��)��"��5pD��(��[�nA�+�(�ͥ���J:la��7Ii�U��OK״s���:|��.Þ��X��3���&,%�	�H`�lS��ћ6.T쌑X�#@ã}z_���c��$�t�bT����N�1٩���U3�e��>ؗ��X`Q�S�a:av��6�F�͵�;�^��~��c�j?�װG�X!�bf����?;ZQ��-nו�i(*��7�'�oN�?��?p~�P��u(�U���&�8��Bp� P�|�4䉡[�:�ۈtj���9y�%=dA����vI��� ��eh�<IoE�7TJ�9v��V��׿X6k!:���N��Z�>f��r<C�tCw9��7s�@�)m�0*u����=�m`�ښO��0q��ߩ7�ĉzv�P�4����
L}�ʀ.��K�"��?\-q���g��ͦ'�\�O@`T!U׹�O��1�x���9�G0�:xK:�=��Z�[�r��U�v=����$=8A$���N�	����0�`�Z(K��Ym���5ǝ�$҄�bL���|P/��=����^rop�?�'�:��T�S��U�{�x���v�)��k��}��q}�C/�	�|3����}�76��z���ֿF iF��缓�=��\ߖ�b��]���qyS�{��:�#,o�&Cիۭ��b9P>�'�C��e��ULv׌wI1���C&�Њ�,�ը��zR)T��(1Rks���6�i�-tӒL��i'���V@v����D�~�>��� -�h(8��*3�����d��8�1�r�;���@5RB��}���h -��jK���:�\R�8v_9��xd �&��p��*�v��cw��)���r����_T��勻p�"��F)SX���,)Qk&fS@�=F�B���$Ȏi�.6�j��Nn��C��A�d֖��O��*7��͈���4֛}j>,K�u�BE�2Q+\&���2�d鐆��qc�w�\��Whr?�m!G���_��UWtR�(���ew��aHl��g_b���gTlX8
�SE�w���
��'=��L��\X��=hi�ZS4�]�ڀ>����_t� t
�/mq�h�
�EyŅ%�$rx���ʩ��{)p@[G��bo�~��a(�Z�5����X/Q�m,ԄO1�F���޹ ]o(I�F�}̹sՇ�� mF�r\�N�{���EZ�X��zOZ1�n���iu�ƒ.9��ŕ�,�X�4�"�1:�@ҩp�C����a�W�����q{ӴQn�][v�n��r0'υ��J	k`eh��r	z����ƣ޷�W����f��P����ս���~���_�s"D�&���kFM�nr��y�ěW��_DW&,�X�_�R_z�5�)4�*�%~$�Cr���*]b���ث��Օ)�Ѿ�}	I���mx)�7�l�����_~*���:��]Y�p�ad!V�^�)���P���K��jW����x�{�5Zt�e|�Ȑ,P�Ez�P��=�]؃��UHÕU��u�pn��R�FO*=�������aE������SX�h[�0����{����NԢ�fAҘ/���;�;������PwZCn�]�oI����_�ƒL+l��/���c3L�8=�;�wv�"8�����?׾_�V����M���?r�#����D������t�]q�I>_�y��G���Y��[���_�t��L8�_��Y���o$���|1�dZ��_�n)3�;%�4������D�D�`-�N,�^����:_-!ț�m��S0Lv�\�&Z��r�A�}/q��j/v�S�.E��0�%��[�j�����f�|�߅��O���q<AWw՞e�3��V��a�n��}B�7�`$b����pDg�vD=�V�+u�
Y�QtJ;jO}�8̞/���~��#�2��-��
?LF�$H\�lFL�]\����N����H���;U���up��h�!\r�,/2���jt��Y%�����@{>WB�[�P���ZD��q��Zs�M�"����~�:l�Ƚ�֡��5�ݖz�nlp��Rh�鹀������'/�2z$l�аױ&1���`����Y�.�r����牒������G7{us����Z�9�>��
^i8�#������0�6��,�YF��Ǻ|>ʢo���t��6�*:�[T�ʶA��1^s�X�=�#���`���R��7���V{T)��	�BC�εwo���'J|����Q�����b'�Hf^C'�fv7� �j���rv�v�M��~W4�N^G����T�Iĉ���fR��ӓ0�	N���H�����)nD@�l@"S�(mP�eb(Fe��C�E���Y��%C)�,��6=�SBIuW�����	w�"W�3[#|EB1��tLŬ*��T�2��uT䅚9�a���8%�xG5�<.(���?��i��hHt%�{���9��d_���T}�ǿH	� �8[�N��<�f5`�� ���X��|�������.�(d����"��s��Wa89�W�����6�5 [L��io�\`�TSac+xL�7��y�jq�Rz��I�H�[v$��K�ϲ`�]f�-���H s��[�Y�����{w�rW��t~�c�����'v����H=T���ν�e,G�5�yRB�CZ:� ?% 6k�Y3�߫��~����a�J��hŨ��[�|��ma�^����9�×14"���A%��kf�i��M��sp���?Y��č��(b$l����f��۸���z��Ӆxv~';}骱���k���pp\;F"֠�;UP��4��^e��:䐤~���usҒ�&��:~�&O!���8�ż���Z������reǮI�� 7��R��Z����Z�OI�n"�^Y�螶�,M�#�L�:@�C���> ���f�+�M��a�8�1DQ���(%��+�3͈_q{Ԯն�"��W*��ܝy%�e|/E�=#J��E���������U����ޣ���[W|k���E�b�9��;�U_��ˁ���e�zj��mRwh/��"����A��>֐W7��9���
A�-ί�I�M�9����es���!w�{X2�?��GͶv2(՗���kr6~*�Ƴ��F�m�=�^( �=��/	�)���^�W�"L�x^$,<��W���JYC�x��b�	�Ch� ��]���W�\#o�ۘ���#{`ǁpL j��/-r^� _��ޯ�J�W�#�0gNk�f��4��̅��>4}����D�dMj�q�f����~,\ ��������Y����>"�����}P3���>���X�!�������c�1�(m`	���K����|v�}��Mi�xno�$�l��\=���dOn�Yg�C�F��P�u'Uv���-&x^���x-IM��B�VݽqO�у�q.���]�|�"��p�"Y�����D��k��b�*�g�
 vw��S��EB(;�4I�vϣ���pu>��' ݱ/3�qS�#�˯A��T��N�Y�k�w[�����:Б����6��k��Ԅ��ee6H��|�}�y����@B�"px"O޲�l�h;�U�W���ދ��/D9;��m�	),�_�͘��"�d�R8��i?�WG���(����x�����R��ݨhz��������Ϭj	0o��-5$�����`����a_
U���y�Q�V5yI9�ZW��/k�4���k���N�����
�!���g5������Hf��V��5@%���|n1�:�L��Zqb�	_=��.;�4r�藌���	
�+F����
�L�x~�b��f֐�\W}�zo�O�����$��E5�!���{c�����d�*w��x��sW�$meW�v=,VV�8�yw����`�Y��ɷ�X��щ	�Z~�J���rY.����D�}�a�d�b�������ozr�ӧ4ݚlLO�_p�U[r�G%|T3IK��"I�b�VsS,yO>�ѣ��n�7�B��\�rH.ͭGIz�pNf�+!�n�G����z�3K:P�L�� I��I�`a���;���ٺ���c^@�%�����\��$�W� 
��7�y��}��ڙA�jd����`|*&M�Q=�V�'�����m�U>=���4�ܧ=S@�Ul�K#�x��X�]��!��ߒ�x�i���m�EHͥ�L,�2&��;;Y��C�w嘬�>X�Zі�e���4,�R�������|�Oh�R=^V 2�&
�=D�=G%��e<����6'1dWL�s
�9Y�����c_Y<0�Vz"Y��Ln�bV(f�,�D/��&�o�X�G�'�s��E�����{8<�7�`�MQ�����,h����ҞG�`�*"0؂��-�XO�^���'Qk\�o!�����>R�����ﾡq���k�U�i'hK�e$Ǜb�:�A��w��������Vu�e�I�&GF�r�^4��~�l�/�A���ђ�z a��8��L@\��w�����~�)*��Y!�Bu��>��6���E���tq�W8��W|c0_���'��8���bNZ��Τ<x�2)�7�d[�C%7`�ꕵg�k�L�,�,�S��s>'߾���񔴠�?6�4Y�L�u>ԟ�(�P����Ӣ��7^�ԌG�b
ݔ��̲�ʦ��"8	%�AY��l�5���hQR�f2�l.&�(�`?6s �Q�J�!�����00�e�e��a�ʷ�Q<R ���؋7�A�lT�	�*9%�kT����rD �5 \zP@�K�˅�^�+���|�P��!�/��y��Cuq{4�7������ऌ>��ˑ�lޗ��4ǳ��t�-�b�HF{�}�\�:<t��������@O�߻j��2e��(3��~b?�������/���/сW�hޗ��1&6'��FL�~��wY�+��P$qI���4R�F牗6	�L�K�R�Ma#z{
/C�%F��f�U�-�JF�R�w����! 5>g�8�Y�$e_����rbi�X-���_Ū�;(���������s�+�S���tBX�/����}�JL6!�2*�g��͠^Ɋb�"��qD)/�泩�����m�yU ���ZR�ds��L�iS��?(H��Ɲ���p����s�J�{�ʼc(e���](�[ۖ�6��M�訫��X�Hv�CkJ��_O8@�@�[��,��-�}�0�!3���[� 6��{{�~�B.[f��G�#7�/�J��Eٻ���HK�X��s素�z�˃�r�!y��c��t;j*������.O����2Ŕ$UW�B+����ٚXn֔�#@}��L� ��T�Mާ��i�(I�k�=l��<��O�Ӑ�ao�Ѕ�GX�p<�[q�>�y���h�g1];�B���PK��ZIH;��)NjySH&9SB�h9���Vه�	������������}>u����H[)A	(�$)��Y�*��c�'��"�5*�3鷭=,�Bŝ���5N�D�4��P���y�^�i�+UL���b̴B����'����u<bm�JU�xq���I�J����ӱ�W������/��M	��� 75m�z�q�2����.!��/׹�^���6�1ˀ<ʣ8�4��6�VXo_�#F(w'W����h�.�kz׹"D)V��z"W����I�pZJҨ���L�M��4������I_��i���j�ai0�fE���Y�@��M���Fr���j�	:����_�=?�A��YeP�ok���2�
��Q���9�͢rD��B)�s���MIX$���5
�~�B��x9�5V�nm����H��/�'�C�g���
������h�~G��/�$�g�+�FA��dt|�8XXԝ�h�xEd�$��]�4(�A�!Q�f� 	^M�B(U�K����'I)_ۓ�2q���A*�vߵ���|��(�	x1>٘rA�W���8�#�R�k��m�m�?RD��A�ů5��{_V�>u��D~�&#u(�:D
/A����
��8>������1��L_ņ;�~��@����ڡ�}�H����XuXXY~���>���j�|:��]�J) &uY:���/��m�I}���Gj!YhgY�Z�`j�99
�>���+��O�F2��ߎ0����F�c(�h.����Z���pW���
C����ğ�qU��6(WJG���V�D�VP�j�޼~�A.�4`�AZs��$'�TKX�䐒Gh��]�;��2� ��؊����8�rr�>r���_Q7>�v�]���������H��d��l�M-
��szx¤�@���� W�O$�K�U!C(Y3f~�B�7̑�����D���hT�Q]
����>r[�����;Jb�8�C���/�i� e��w/�Nr��) ��e��M���'�����������Ue��1�	e��N�rPeߚ�ۃ�^>� �!Ĥ������V���A�O s>�:k"�����)���K�sf��ǈ�^�K����UCh]�xM_�L�b^�!،�XXJ������� ��Gv
��6�#�먴�
)���t�Hvq3Ub��@������k�⮽9���AVKr���\��΂Q�^+GGI9�ǂR�4�����Iճf�u�8���Wb�ߙ[�8�[u����2?ݬ�N1�,�Y$3}����~��{�&ǍT���E�s
^c����l��c�mF��K�Z�w,���v�9TG�+�F����H���0��� aZ¶)r��ߥ�`治�U� �A���ye�?��1��8�)�M0,�3��47^~54�
8�I���8����WR�\��כ����2�u�IF�\>���l�iH��K)��̣A
�*Ch �����g463#׹�w�p�'W��p��>ݧ'Uy(e���#j��:ON��#�%�l����xt��� �8F����q�^K������tg&�y6��^�S)jo�j��)�t �;i���~�B5_1�z9�}X<sE\/�a��p���t:�_h�~���Y���D4;SQ ��>�*qug�@���ɔ73L�W�j���t�J�xOx��Ҩ�p̓�[��#ٙ�3y��aS�ǧ���v�՗\�ڀ��>g�<<��mX����p ֦+׭ϒZ�7�Lc���ft����GnG}�Ҏ"�WD	{ [�{h��ϚB�K2o��t��">�Y*�6��z~9�����	{5K�5R% ¡�"�~���I0���dG���20�1�@����3��^⸴�9?�Z��T�= w������>�8�y��2�F"�f.� sXtϦ���b�TV��lZN˟u[��p�3�[���u�<o���'���'�1z�������/.�QVPZޣ�0��GE�(��,LJ�ѿqd``/,���Y�#��:z�<X(��9�[��P�*����������q�����s���⏁�nռ�1�������'v��UD�̢u�/n��+b�r���F	�*����7�g�B���9|h$��do���91�����b�E��mGjd�2;0��a��cZ�����
(1c�'v��?�_�O��|���MQB�ߛa��N ��T�#��#��z��'�S�v[z���:��Pb^���@`�u&�?��c8����b�i]���F�[b��F�g��Vl��Fs���_ �k��0��������D+7е�Q�ij���U�&<?�Snx�c�C�]��э��߻H/#�%N��G���X2|�ǅ[��.*�:Q,����,�J7.4�"I�0�������Z�e����N���|�2�~o�,�i1;����j�D�����J֞G2:��f,�h����%�.���a��z� �j�ڟ�[(���&�����Id��g��ԫ���n]�0|�����Hq�Ub�Ӣ<Xd����9k��=���D��ˊ��*>]��}��܀+0�>�0@W���7pzY*�)��=@�.����1d����#*V$S O�ah�'��k�g�^�n5����k��?KE;t�����Y/5�U��P]��X�9�����ۈ�*��p�\�h��1+a`�e�W��K.��m�k�F�h�����_�kC�������玳:�&��r ^���t��/a&=Բ(Ǹ�t|����4��9�ed`!mB���y���hj��Q����ZwZ�� +P��-/C$�����6�CԨ�9!��.��\i�L�z��tC�7m�"�DzH�áeM����P��w��z��Ą�-+�;�1K�M�T�����k��ٜ�NG���W���77RN�XVZ�o������w�C&w �!�c���a��t<�?�S�?�Z�]L����5U)E�C1�C�-�(�$��P��Zߗ.Ń �&�n��U�]�b����cc��:�:T�	����[�S������Զ��E�n�^\��y����8w.�,mn�}�tm��1�^V��/;�LN���a��'��l�Ӓ��j?V�0��"�w�,�dj.HV�hZ�ȏaR��6�Ð��6U?u�x�`��S����v�|<鞘zf�~��4����K(����4�{�����>�W
���v�Z��S��|4e��_��Uc	�H�%���&�Z�R�������W�������>�z����!(0Gx<y�"ֵ˫��uW���kv�����v�g��f4�MB��!���Y@wU{��4�04C���M�@��y��N�_�;�_�;�~&=��n��4�0�	�_��"x�d@��R��
�]��dϷY뵋Ɠ����s�b�-c�2��,烑v���i����g�9UK����khd��e�8D��R�|d�o"�L�"�25j��D+�"�ʄ���&j;�T��EPh�Όmk
��D���::㣵��NԞ��j�_-c���>�� �D�O�aq�Ce�,�O�9�F�������5�#�n{����dϛ38�D��p�F4�q	�"�=�S��֒۱ס��"'���:GZ��LiI�)���0�]6P�NЦ�N�-��ŗi����N1�)c�%�;��Ȍ���,�7�/Dtd\���fP�rl�͓w	t"~AE����	z�
��\�����7�J�a�	���Y ?ѽg�\�<U �s����pT���YXЉXt��FXR(iX;�����^6�1,�Z�zLܨ��(�g��3yG܁M�-f���Ϗ55�?,Jc����q�*{O�@�1�� Z_<U��p���ކ��1�����J=[VV��G ����i����1p����1�or��-;����ņ5��� {`�4��}q����IJBj�9���A`.v��q=Χ�e�6��+(~u%}���DQߗ�� )��m%l����FӎLwϴ|��T,]Q&t����(�Cײ5VB�,}�_K��Y�?YX2c�}z���%�h@�<]�κ�C
����B?F��G�N�B+1���8|��`WlX�?s���C7�Y�Wu�]ሗ�N~�!i���U���8 �˳':�t��X�S�=�M�/eی-Z��#��{N�@Y� ?s;w�F���h�}��M�媣]H��τ~o`5k�������#Z�-��9����~�L�o�o���.H�b��h`��_ҕ�.�9��ýK�����݂�D$е�p�a����h�#Q=�!>f��Qa�~D�9�A�L��|�\����*�mY����x`��\�W�>Q�ʬ�T��4�3��123N�A/�}�;�Q���lZs)O��=�Y6��$�r�t��7"��NC��4�&��m�W�3�@16p�L`��*"]\(5={��&,��Ǜ�˧��Xg�Ώ9/r���`��L@��[L����/��	�L�f�.Uz�Y�@DQ3c��h�&ۿt�(�����uoKd���c`�{��7�UcI��c��ِ�!�6������5Uy��� ���i�X�8@��rX��vVo�u����������$
�e}�l���p��Q������o���8Wd�����c���f�|���/aR���/m�p�I����k5�QQ4)��'��/�[��ڵ�h���wD�.���۹�w���a��y]�5��p[0/��Gҗ �?��>Br�΢�ƿ}�Ԁ�4j�:
��5$W�3�/7lp��IWa�t�w�<J�v�Px���X$�~�!��,/LS@Efȡ� U�h�:�彩��h��i��nn�j�w�kma��Zw�y~
TS�>>���w}������;�n���\_hwE ��sOb?����5c5#X�]���X�.䶻9 {j/Z�M^R���7у�%�T� AK +�*�=����uc>�D�
h�9&V��Q������{�$M?���5����w�G��zZ��hvVL(I7�eQ���懫~ivEq��@u���.����O�Z;)�\\|���Y�}���O�V�'p��dýf�n�N������z���}!���$-����_�/��$U?�ʢt��s6g&JE���Uo��������rp��ٰ"��";h͞�:W�%�{א(��c0ɇ���r>~�/�`� �\