-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bn29/J+Txduhle8E+NQqk3zo6iymGjmjoGF+5qbsCzV46+IjrvKNEYUb+c+sPnr8Mot9iMyMIcrp
BTO+jTlCg0EHXyHwrSfrwwWCaaMfbUyFLtP44jJA2zsSBZeJUnUhPHceskJi9eCB6yhoMQTlUA+Y
GRJf0L+5AnhdbL6ur19xlKW2jkHWnSsD3uxlr4jAN0qUOXoTQQRDJmNmbQTSxmce3Sr8uR8vrYja
SBsgRyV80I7Ter04i2Xd4j1YTtpNYBossO2nL+XDzWc2ufzTACSJJPo6HdmOxvV/tidYGmqWgWof
UBwcGvRgLgv55B4l+NWkFJzoGR257+aKheiAaw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
Y8ZZMzomedst19QcTvT5jDNKj/GpsD5ZcnonuHKca9UMq+Zlq7u+Vy/bDShqcV48LRRj+gESGCuW
3N7e+b9kP3C0n5HMfEJC9fMtoKCWtL80f83s5jhAMoqI07Tw7Ir+HlDHzu3h/We9ZqPdMnPn/ggN
cvUDcXoOpUHFL4Jh8LSBAEBK+zbQkDORezEmGjCVUAO87eA+s3GItZ2JnGxPEH2DleqOiqp54zyA
p7cB6KrwSTSrlvW/TuKpWyij71bsJ3quNI2DCJjggY/Jzp5jutt54tyT/IQf9XZOqeVY6j+4RPql
tPNY10QIrMw30i+VyEiBH01j8X/+WvZjwAxN+yX+3ZHjv9e28PFhlCponnCfEALjSZhITiZzwPOw
Q1NP0dWeiJLtRDZadnK3GftySlJkt1OhAKM6AWkA+QNVQulDKiEYy99pNRnlNGtJarnUyoVa5HH4
Yc1hc0P62T36y3K74SX5K6Gw9wUE2sATa1pS+TLOwyvXKQ/6zAKy3J64gfiYRO9wC8+GscqVZra4
UyZKBb8khrlS9O7uX54IJxPy8sVFW45xgBCuYLoQuiY+fDiO9ZI+/2y7lgHmg/utVKki2ZQPHmyL
g9X04m3MuzHhwATyG/R/67N8R6e6eLd/pkwXQvOBTlGRS7n4JH79MC6IZ7iHnzi/8K9jceMUtDu7
YMqgkHaSBzu61UqQAa+iJscUIRYrb0qEgpt2uMSiaNpoPH2bDou5/s9AbqhD0rtnituDm/Eecynx
pN5LiyOTfPMHNijbYusNWjgfbzYvkc7ogV081wMnA5f7c39GvJuPN+vY6Y0I26Uo+vIkRLQDIcdq
fK2NrzkWUdtUGLx8/FrYWqw8IDqcKIVHZTbwusRklnVeoyXlIt1koMJDLl/jvImREAEY/umC9dGK
2pXklxWPoEVQIeDcS9m1bsJcjflA7A8jWjsBbhoHhIMpNmgZxaot/loRuD9GmMS7aATMlqvMkhPf
7IMIJ7S5Hr84YphdnADlZU0HNw9WC7MdFRY3FlKl6346ovJQAzsn+uLCOmXEq0i+sC8aGFzpHHYj
vO2YyRvKW/42LBjdjtrRCZQ2J6wV+byH6OcT+p16pJ266sSmY2LOsHcEwuA9IlZwYnMUKkGA00BU
c0MMFmi0SXgufxObvmphyAC+WP2YvSuL2PeO4YQzoXBG9QKFfRgynjAarJhiOmHs/GvimQpA6T13
E9+mg9ckfhgtC5KnNaS9FWSB4wdX+gbtvzF60it72PxVMFuXjqbVu7efFSUgsvyQnrPAyhcxRCNr
opbSPdS72Mj5RZXcktZBT4xfuIlwVHlZTNN52JbwBG653rCFZmBEgfjrti+WZJ9asSKEpe2X94iN
JDB9sMW1rNLY/SO+ywt1HE4oMjM1Sul3sePdLcImcUdNl6Wui6D5a3yVnaAesuMzMs4pywm9GcTU
pYB8/q6bUcsqEi9ZbGDiDFidC2qUpnUzZAHlMg8Hp5iCrQjTd8cpfsR82sH/SDw2/gIxxIPUDOeO
hcJLu0d6xstxXLlSQcj8Xc7EvVH3uYAOYEg9OfwvayxG7sTwcLboTsV9Q5KjxxHvVxj5nsIHvqnG
fU4Bbga3Uo77EIzBSB/WMTd9vAieVDSLlFJ6Rn+ojb9cSIOHuwpo909IRWRYUXcS4RXSn2bzugiT
57VajSqrlAeiOZTz1X4/refVgx3emw9AEzJgad/WDD7ETHPntjYotysZbUa5lZSS9eP9YRySty1A
hMgCE2TcUVyzrKxzZ5+W+rlrwkKLC6ulBkZ42XS0cr/D2M2qEWS5LFc0XYivw4k+lGNUZqBCwCUr
hrNIT6k9SK2xFpOgmA97o6dp5Fc6MttxbdWJmsmxoIXZ4ArCH5V7RENx5GIxDUhZuwbIyjaxYHaO
NpM2RIu2VhzQfaDsU7wKaPdb/hLJ/5k4Rt9VYCVoR0fUjp9sJGsco+lfRmGwFWpP6Uh+X04LAi40
yZ1uAsRKuwxxkIIYKVHb46sCV6ltmlELuRIp2femf4VMPDbprWZ1LBI0L1LUrxBixuqJVbPR0YNn
zyOVe10SZrwXXHNaLOc2njzbVWuqjWVMKxjp8msOwhQUzfnOhuDNc0+97VwFD+UlC13KdS1bWXmh
I9CACcPlu2k5JQNw7p8fCS0Ma+DaQPpJLK4Z5mlcmTvLxl22c7ReI1oR/gOUokuQCcJoN54e+bv5
UsEjsJZyzpP403AW8QRo5ScrXTdVTn3PhlQTetFKM5bK3lkFtHG3PPFrlG99CkbcB6/W4LT5BLur
IzfX+8x3o/SC7cNOtd35MPXBqoBm+PTutUKYsVZEdSaGj5VM8eVVNquLkWrRb6yVnevETWwxqqvD
cK+LwSYWZbAPLS7GbdA/l3T0ymoGCV0Z+GJKEcf8SegC2kdAUdqWtrBFdc3lIz1GAcEmI73YW0BA
4f2z9rc5SBUjYZ/zM5OxMTxTV3Kvsr5W3uZ5j5yR2kqpcV05ATvKnLwlbk9xAdcOUbGfYcPoQ4Kb
CgRZ4V++hfBCpz41z6jMvwzIu9KiDhPFjvTYUAHz6svBT/oXG3qYYWEd3syOOXi6aoKU1n95YMrE
a2SUMPTBXJ3hdQnNs81zLKz3C5psdjhoypblCybvYfLWmyis3zt4uknhBlMQ/8+ZzdI4TpM82ALy
4Gk5MtFk1x7RyjscTHAq3Gz1cwJJLzCinHhQZ1Sasc/UgVqEMsoIcoqK14llUjvH/tjCXwXHLV9y
0/Ml/teOYSgWpJRzmMnd9LBvoK2mogcJP2FOh1z3ORU8pJmgnNjPPnaRA5TBoBcSo6kEZ7+DmIRG
svqnjNdWCfK0LarfUjkMql7toW/XW2tqC00PWhLjQMn6igt5EfVEvDe7FtjtHTCEfbqk70dZ1axQ
PwIKjMObO8cJW7DapDipVD6Ib/9giw3/FWr8iHg/rrDNR/ejUPouE0M7pdYJ5RiVV6NhAub2KIq7
ySwz/lu4T/7WbJ+esKL/hZG8cYiZe7UPELsP01LV2BB+qp3SztWtAo+t3m98BemsHMy9ONxn9xCi
/nMeueqW8yidzUq4bvBVzI8JNJ8OihliRurdJ8HJEM60bPS3bXAn16cmEpmAQ1rizjtm/i1T3UMh
Hx8tCm6aOZQNq0ifCS26zOvYKkM0pBEI9kszfgkgfYduKvPwCWPu3FXsnBwvniI3q7BX9bJf7NAD
WKfnmVSYspc5LiE4u8mvk/ugRisnywCEFodnGumY6tiqfAQ77GtL+wrCQleDoRkZrS6ycf3mhW8J
xNSEbKQZzog8G2fWungGDPNj1/dM7gavA3I4BBO3T3yelm38hxS46qIHRax/aE3DVmOffYw72yKa
pglUyQayAJ8Tm3/0EWWh1YIZxFisLMQbWuxZOoWVUkAkPtEzJRa6jm/q/34oDxlvAklbaOCAc8Bu
chq0oLtJIlyLZwfna2KSHdJjT4TkO2CL4vgn6pycO4TNrV5zG92dBc64Tj7KqsCiUfAHnhJo2I3/
fAVsReuWkKyFx58Qg4mjVhlZO8U5QzDDCmxAr9/qRDeljrds8dn96KNKqqjQttYSDjIjGAftw9fp
wO/1IKePQvPGTLFjqvVKV+bebR0is3dWy7RVTnlMmGd0CHonkIvCNGTCIDbJhjjElreOq/aioJc0
TSUZd+sFLp6kI2latfmGOEJwlhRW5tSsZaxp1svzuvu4qDS+gNKIotzZpTW1ldkQIR9FPfRPu3cq
oMcvTVBkFP9WDjZsFwNqqtrJyJXgRZFrUjq5i0zc3tMieG/lsL+cRzepIu9eo0CBttMNkzQPWwso
0SU3Z8T2BclmSze81kY6zPqv5+IT1CI5diRVZ217IcP8y5DwZIdcvsVmauq7EBS/KkbIfhV6QZYw
2iYDptfj9AXBefEQDEwSKf8xsCYBKJKo0t3wNqqoaEWpQLN44h3fkMOPZp4BeDrbMEo2wiP8j78/
JPiPhHzGL3mEdu3gOOn7Zb/5ZXtrcH/g9gwWBt6dWJqy8emSPzBhPQU6Qeoxpc2EZ0QeiOH+to+D
qt7Z6/mMoVg2s88ilMwsYeIb61JQO+89pgrpUSu9urcKqZ7l2XU7rPq39Febo8mrzfQvi/zZaVF1
iinhH/NRK8CWUnRxkFz5fEuNrF1wScFGNIpV2uLQeDrKMKH9whOdGS5Fjz8RBxDDVVsufpPXm9OV
pdgb/zG03lfeIjkrTomrJoW73m0t3wvzuMQ1yvSnRf5x93ly8gh9pzWwTjINPZvKRLwpX6kZY+rC
bq6EpXothDE1mr22Uu7zBhnIEOskwvKHaeMz7YNfmvdJ9R07YRaf8P0d/rOgWOcyCOu3l+hncgAQ
BCEzdN1qfSc0BImGHDX5RlDXdYoa1natwXl+DtV9KpwiWzlWdIsJqOnA8PU1Mj6Lc1YDXc1o8gti
g07gi/hkIqvImolccL5QSU444sVP5fa22xEvQ2dHHDEJuTjTe74zn9a743aoYERG+fP9qrtDOtyd
YLYSfPY/qlRP5aryd8gKF17GHGhIL5aq/NoAu5w89Ku7wrGNk/C0XrhCy3d4wufLvgKE0V6jc97T
g+qLnejqGQcgTwQMP0NooGROOaHNRDvw3I/VMBl5AskukQEc/Q7kD1CtzxOldkICgIkLEhwPknRh
7fVldpOqD7Os/wboMWOMiZ3/wDzQRArqzj3v2wdjJaCWX1SNWHihZmUg/BOMMVjf4ArQYMPpTfDd
AajX90tJCCkoIl+w2i+xFzpO6267IWU/LlL/zO1F7/EsMy4N7ZMmrAil3KmXg5/jUt0w7rFRy+eR
pak2+XA7NJOllMOxvZhPStHmTGsM5QJTcRHwSuEd/X4GXJ4PUb3SUXJZIbC3dTbU+D7vny08xI+0
JyevBxxC8xTiysqDbXD/WyRxFwltYl7AW/8ytZ6h7k6cd+OdQFpdbyhprHdFiQ2OlQbEREWUvbS8
fU6DweOyUpDs1WjmT6S6HZYLi9JU25NZohWfASCvI10pb5HPopYnTePh28O2Q72Bb+MQd1ClMl1+
4ppyfniAbzGh2HomS+ptJBgMnz+jsgqWLhzom2GrzYMpRhhtpJ65t5f/MsEcwiWAsn7m5+0SS+kp
kvQ6SPuvER58k6xsm0DMRg1oBNmGxKGyOra5Qrnnd/VfZGobniRoc0HGruXbksdCjurdd0HBRGVk
Y/99t2d+qYPABfUKDl5KDw3u5v4U0lUfaZSf1q6Osr0FU/V4Z7n6clp8Dfd3h1OvR+GyRWEzrmv2
hYeLf40KQkEMx6zWxyzQ5z7jIx9koaVm5Aw4IEvGPYRFaufIDi+WpxWX5CPyM5oAUl2A/4wRTXKZ
Rxq692HjEApOXBC1wTFlc5q0lmVv+WUln67DlD6CKpCBDpRV7qpno6mZO+qmTyHkJw0cMvY/xl8B
uiPjdth4oycpS2kTLhAixcBiuGUdNgua/CB+f7nXyODe7QmUylt2czTYn8QVrqj34HgBqLZVLZ34
jSBVQjD+QsMDTUoImX9kE1064nzvo/N9kUEfmqy6S50T5DWsvGptP4Os4KVryB17FltD6Jfdfc7T
i0FSeHnr0MPztcxNoRqc978iKTb5OFT0ldu6Y3cjl5wfJWm88QNyAwK3VfgRF+SyFiIOPG9PPD41
JY/SJumEGYDZn9l4aSNiIncm0REKYMsjw9DZAiYAjx4IZ6PcgG+cVOST+uNUhHAOG0vJHiDDxyN5
+CVj+hxqQ7uUeDU6CFlo174q8dz6Ml9Feoz7fKH9Kdp16/qPsg8YQv2K1/6PT3t01Vvpehu4IezR
VyBumL4IoU/J+F0ZDmBViVNWjXZKUXxQj4gZB13+n54j+IydswMmzWxh0Mn1htXvJbtPA3DC7fBe
BxZBho0it1wVK3CQ0vOCOsNUZEMiM/rQkSuA3W0c5LVsYtjMNBy0TlXIinNPYCJsnRx1srsPkw/Z
CMeftyfhiFezl/l8/FkYk/tljsWm0Byw/LFfLuzVjwT0XOsA/kV6cdVhE73ZGgm//4ivy5q77iII
lbDlg7+4btFm/rjozYZqcExjnEUXYp2hcOqF+39se0VqFkWjD6xz3sfxElzl3h6K3exzklQdwpUL
TxZB/yeVsb87+kwXSL+Mc3X31f4YdvwkiBYBvtlHWY1qn1pBu2LOH2HD1jdsMoQax0B8pT3tYpKB
G+QCI3IUg8qz2m+RM7GhgrAZDlN0iaeW97sybBypyUgbA10/+46uVvKRYRzAq46XdtRjq1Hiy3KD
PK5bTWFqq1F+XCgNjWI7gHmxZDxtQOrdM3KLHXhuhEMP3DjNbyn/ZzkcGkxnmWC3yfbmqnkELRVb
/npgILRGKLZ7PjjCcjgBvUIDlBg1+jaAuYSayOcFkMCI5t1QXZlHWJlj8lphdP1E8VFlRkAd36WF
dAItOs0zSk59oqjj7YCuc82QdPS2OrxuyxiS3K78Po8JITAT6ndhKptFuSazSEDnYZ04vkI2/75s
N6o5k/aTDhdewrBOsOJwy7tNuOydnJ5X0gope7ICdyFJ+IP0hQcOlXl1hxR27/0u33mbBcmYTmoY
rFXm3LFh3NaRHtPTgvr/Dnt7W8HrSZsumo/0Lq7CJVGwRPpBciyOjVVGDD5pmlXuw1UuRk3UVJdx
FUzyF/cXnL1MU/YKP4CCNRBo89zJf3er/quaQd4S3L0FYqdS5gbi8gj1hKzcdMTEBPsJnH8I0PN2
dlAM9ySvlk82nw3+g55Zr/q7lqqvaFzrkrmv0O4E2ss21AvJ+LMVjitRs0YBuiWj9DeW14ImGFVL
BJG2mVdmJIFHvAlmBXb2O9CVIC1RYTDn6306z+QTmhmSf37XhBlGNfRqi04/wtR9RplQ930+9t2R
8OwVlL1fKjHThcHfMzl/tQ+XUUeAjxSmqUUUQySUqizP4kznouUKYux/ddVcXSAygXZOE9hEdc8V
8waKDg+DkGex2F+G7Jgbmv+3bL2tqm9OI8JV1D70l3LKeFE7NsT613ntNCVTZPSvEOFT3u2uHi45
F91Ne/JKXaA9JjxsE7OhNAz3ilBp9AnLpqSg4KXtirx8fg9blTQMSSPjOiuzViToZxXB+mrnw4/I
gje0S9TkIjU+AXj8939eWJ6Kp1JHnJDTpDJfNQJIPPsBDW0kMPu7U1JnwWx89GRyydKp31ldBoB6
5n//osu3D/21GuhyrHTRLRkOn0ximRDX6FFWuIoBniyRHKPXxOdSYgr/diI3jnobeFq/RyhKXauX
c9RsAKgumDi9V2PNQcKAbWeC4bmrymEbp2efMpANTwKji3YIli+H+ewHP1tlIUhogBMwAKcqON/I
qZiJ//WOxqxqqiyiJ5zJzmWvTBdSM/kfnlMcn1CiEXYT05AAysVNLkQFWFJcrNtzMjvsg1JuwkVn
a/lcDgPW6RymYs/dbUp1C2wE+hI6euI2Bw07l1b+gkiUlW3WLUDQWUYK+X2Pdh08FPfQrmgAVZYV
Dr0YcRjo+7dvSaiUsm0wPuHAnv0MlJBdOc62a6QmMf/c7+8kv/QVLtHOgCTCVkwxOPEdpDP5wKo3
Fcl32rW5NrRp/ws3AQsAIQ3ruS6vx/Pz3YaXQ3VWi94DowhIxPgNspfPumYMFy+ptujSoPnC97bt
mfCArVEGHP3YH/4KWJO8Y73YTQJE9AS/Jp5oEAOswP+LOrYu7gAIfCMU1NRV+Q0mXSUcNqAaHpuC
N8M+Je3R5kf64YyErrReIGAmRlDvNJiglcCtPXwYRTY+SbSP9Wz0vFxhAURel/xADTkhhpnUwQYb
N7YjPZBul41AvsyhOmczE3V042SNJ+pWpcQEu+166/+PFJvlV1SeozVBJVH+8G6310uU5vEyRI5/
1HIZaYqbRKhNmRi+dmVNgUfA+GovjcJP/91fZsCr0ghRmUKDs9Q1HLDg2UCPf4uY0M6HojHkCf4R
u2qCjZmv3Mz1V0i/xxczhmo395g5QoqRiZchfbpeTpHEABl4pld/lsRyejZTTv+VRW7N9YfL6xKh
UWnLXjzdKkxebgzWK7tFRhaoIIOqxb2TN0mH/4NUE+6Om9oYsVxZQNhI6T3fbsKAIURHJjFYd7Kz
UQFJBG8lCHUCeMqJcOZ1evBHltJkqLPfKcgMKoIo6SmIOBk5z1LaOdPq88/z5KsdU5y7j7EdggES
wEAgvOC5SrFf1+zJ4RyjM3WWN8wmNgzb0Y7BJSd3OaIzDjsEr63yX1mHzUHnVQF29hDwThUf4Gxw
srGyEo5sWwsGdSbomaEQtkMuluioEDtvYjbZxlIB4jR+iuCj/jiSys6kufq95HyIhufqpUPPxr/+
XEuicMePPIW6Ys+UREWsjyiPA7mp287kAZ44ktXyk2jf4329F7OfKdSirpq0MOso+0Ral8WI3cj/
cwdNbN2T8bWGRmUeA/ITcON78X4nh+rFwEzgX6A99VOwWpB3e0kqCuSXqb7xoLe+uszHtwxKcU78
zkmGoiN7MwIf4WqtEHGwUwkij/t9hBDLFpbp/I2qrhgnETovez1kfdur52/HgBGJrvEOmB5DEei0
E07/B93/xxYaqS7pgjF4Un0lZgdN+kEF/mkviUut4QHVM+8NYXh5N3g/MNqOX/egmaQkpPKzuJ7o
PHBRZCG06XkMQg9q7Ky6PMA30/XOlpsRzTiVFu21S9rAsvhg77Z3M1nQio3EV/Rg8x145BYKnG30
JDSam+dOa4e/TIl8s5L4/75F4F4W86VxOP209+EWkSty8edxTcgzoLF5mMmNNBNvwEpBw+b1klKn
tW22oICW3taWaYP2UFBsFG/pth1VdQUDl7wGIoJk1BjI+H9jDSp3zLFud6oKcYxhiMoMSrnVbRah
e1RHylkMabyNDy4l3lbCNQiV5ZwweGX+ggRViVvIKGDSQEkrArw0vN61/LqiorvpUbZKWKIGvrsv
sVGM9mXA+0DxQJYXz4ixTY2S61YWKS+ye5zP0uo5fWQuAhHY9AGbxr+aSUUPQDPA174E+nPUK+Pt
jdTbc0AHOO0GhrknKomH+KYRuUHnRoUkINfIko8P7FiNPl8XGL62YWJDr4Y11CU1YmX0X9fYUPar
F7HKdNbCMAX0P6XBKykr/mrb7FKYYLPWQOhs+fssiEKlWjVh0vBtyZMMheNzCq3OHQtSER7i+RH1
V2J/17p3ZOUY4Ta7ShzlD1CpIhYmfg/Me1SLE6x7TTr6UGNq6MKk57opo25XufnkYcrBhYMj/v9t
V1lLzJGXqam1rquGRT1iTB0pprBV9cDwTaK1chInzPBqwR7i9ljy8hvJFbwK8mFD79IMQQ34Frq1
O6aq/5M3/7axthTw8N496iWi1k3Up0e2vN77Y9MySgFTyGOStfi5pPQ9/tBs1qQz4aIhElrUBQLH
oeajiAIVV10YNFz8EPkSFYcGHP/uWD1pfxIGOg1ZqAwuap/KS5q/wo0+BbSvb5JihJw8Q3tdpoCh
FIV7aMJ4KSeNRFWFuWR4NKujUXk48yWpYLBlA/r1ZXDlVk6AzUBtajS2Wb0aOwK/M/hkyKdzecJy
p5FBAmjBt+Ymfk88G2eVAa+IKpj4qTwVWiT8TEHZVel216pCYiep5vD2/JdcHEF+udc/OjYwdus9
y6iVbNSSHQuaDQgi+fre4Kis6ME0InD1REiyKscZlzG2+Kr2bUg80S9a5+SYvk5UDXSHa7oX373g
vgrNNvigS8Pb+u5drqBB/0U5yS7YGWvsz5yMdnFfmWeytUu38EXhTLiFp0iG+QkQTBLIBhyj4my4
BQhT7CMB7UD4RrhotVjZ+56GWwMvogyiBOr2oT3YXWawI3ltuufOrxYDCWs34t7NrzDpma4sYwo1
E8YrI56oXeXPmz1zMC66qPXWt3AkXqzJ5F1m/RYJb8vbJS3pW6Jao77l3ZptIJo5qEBgI7Yvc6Fh
EoA5+3J5yvvEaUO+JcZNvbYLGzh+95I+6Du2Y6Qndbv3O8ne65wCZjDm7wUKmEMxYKh5iNVGwcQf
2VE+bI1cYrCLWGcfaSLBpwBCoptkh8FNRg+TGpxqYfjoOONh72NR850mRf/5o8WM6B0p+FjivhbT
fF2z38XDqJwZWzFjPEFMhYVVwAMSyc7AAdzI/yYxh2LT2WcTbshijV+NGwE7q+/g40KmPXWuAQBQ
/tc992nHj/8MDLZ/3k6yQWWG67/c6THlPv8i1rRrDocGAmYOPu7QJ4GfvzkziiqJ5+WXrhYhTFvL
5CKDGvzkdivzs+g7rGSqKEv1ojYD6Vi7EMf0g9RMxwwQ82QKhXTX2S7jfiPAdHBX0N8W1gXqGMsw
68f3HMQs0ehtZ6D8Xwad5yI93Mm06FbjGVJHHyerK2Pzh7xlnbt+olY5zrPoGFTGDVPOwZiyXZCV
PMJCzgjxVxcoNkXBo4POzkkGO3j/jFOpk9ldX3HZqUS/mRy600dcaArRrCewjNpYkGbu+qXPMW1b
J5O4ECyVgC0cb7Qx0vED9rJknhdprG4kdo6BadPGSwGi8p2F1a0KQTyJIQ2rBUpWksy05f0r+1lY
fP2yK/jyHBq+JWCBgj7tviOAk0himSEUHyDxtIzYWJJgUpxc35Elu9kVrI6CtSvL5iANIVzsTvtl
sPbwNIRpgek9wOjlqR2dKE4n6C37JInzS4ZOHXkB7S8Kv1mQ6A0wBOdo6RnAnSwIJGALJvs1P38Q
LubjR4wvRLU+BV9ZJcR1vnekAg8ByZfnzxokVmeymvkYPV5uOsNmjq7YEwB5NzxDRC5ugQNdfm+E
T1bTTO3AOfpa2AenqrXmcw5TwNHZpkPsXfJNeqKFtYBVlnlTQILmIdXfmgg/t/GYyyIJef9Jtr44
hyDCBaEPRxA89WWXyyfiD8p3N5m1KXXL6XbRl5E/IoMlskxlb8PkYVFGl/AIHfohhxZ31bZ7mIjs
Hj4vZdq6sDq9SqFDozehZ+3hbzRS+tfUyF+rIj13nO261O3yd+fw7Fw2AtNyLpXxYumdb1HSs+sD
IyMGjJUYJ3PqK5qDr4IexFT6cLsJyQOqyzSZcc2oxpjtI4jH20XVAOP55uzMTRVyqJA6NgpGp/9z
yl9KInZp9VB5cM6BQbC5t/SocGHLSTZXbXxunSC3S6s92nMj2t6xi6egNTEuA8MNNMY/DpmV2U3m
e9OaujgFsTAszalUO15ogsT75MiuEgF8EoR20TQ6Cw/udZwquyljNHNPlTyFpTptpX36FRN5GtHJ
y4nC4smLvzf771FizRr/dWJvTE2l/l6xveQ7gRzKVovDQ4nhjLZohzPRfjxekHLk3OgrZsP/Dr27
AIycix7M9XZyFBx9ecpI5GnwOzDKwsKV3UXgJnkONxoeQ66B+HYnU7Y+xlVJdKz0X9RNspkzaEfx
F+x+ObGtGejuxOg1dXGIBDPQKtaxILjRwPzJkGeIF/VPUso0iejNXTTN7pTm7JujLbGAoJTSHRF1
n6LS5g1Nwxzlc+OkfiyksSWjQ/G27Lh31Fm3JDoJ0pwkQk2qjOR35lS1715R/QTWY3u0wChU0mol
+qBvMlTquI/Kf0nrO+OSAh+hPhvEagATZYT13vIrgYKU7gYMP8J9l0jbU1sq6JQHWubEtnGrHUOj
Tv+yHLUyn2pNnup3+uQ7yVYoCJJdyUA0gqHWYz4sRbUOQx3KoU8RS7P7z31G9+g+EcAqYnZGj4or
raZY+LfkwVswvg0sk/7bYPBkrvbdsMm9ESUSOVpOEflZ5lo3cCW2TxhjSjS8VuybvPMZuoq1zMik
AlHBx1AW2/L8QZ9dWErz5UoWZhJtFTPvbqOyVcCGdkGDiscvcdeFWBllYkIu8rM/Of4qczfu2Qxo
b6dlIev0/0O92D+aHHece6cvyyLXgpSx1uHA52s8a9SfHjwIDD4Ik78g7Hb4zG6w+L9vdGOVxeX5
57AdX7AdIJCtUSlBovUCiQ45ABsSpZarET1PR7F6do5/Xj2ZW/zL8Ndlg4sEup+Jy66tN6u5K/qp
GMljAKp50pc+OOUeoTaAvoW/VYovG0UevUOb8V56hz3+zzxadgxKow3ryzWaLgxMLFWYxEykR7Uz
AQWQGEn1U8Xb0KWNMMYpnWUP9qkJd6AztKrSkgDoyli8mrTummx5/UqVdcwf6TuPedineq0kmYXZ
8Ry1jxfBViG/Xy2e3FN6kxmBNbbimE1Fspe6yglDJ8EUWZnxYdSY0tGLl+DY4IkDLl/r6PGlbyTP
hhPHpjVUOAzZ+3/S66lJ/IrETpqUCWZEJLfKQ9pUSQZgC1FvXF9NsLChinhv2DM3yisqQDp+G7Fl
LVNAqQQD9U83JWUkgibssTm5q/FCMH63nxOTzrchOMMh6pFNieVE2rMe8IjCd6yOKdOMC6qSUOBO
GS5mbQX7lxoESJKtgn6MO0YZVO0UtfwPo9FDESxtyV+L1r/ahV7clPUDPDACRcFuBIIQFoBtMoD9
55WgBaKAo6t/mXwbqLjX/8cr9tdRqP7B0fi5SP5nT7FXizhoOOoxe29ZV21iE6FqLK0gt5CZfJ7C
wDJO29EK1T1qkRFffg2JWeAVQtFB6+2h3aIFbhvJ2t+ITj2KbwXVEHAoMGMvGDE6NnOOqCMpQhwc
+n57Uwu29IUb/yGxB8TKoRIqDrZeGN9Z/mSG2Wg7hFLYJY/ukeheF877MwQrIw2Lw3fusnw5H4vY
3alyeGjNb7vXlDAU7BbBdf4vvTH2T/FFPA8a+s8twU2NXCRBkSIFI7LEfetLNnWFCi+vaKwQ51UW
6LZ1SiHWMecNHsSok16+jRpnZLnfmzS4ov4s7EgTBrQTRE5uaJ+xZlxsa82dgRFJtwm2rm9rtlnm
kMTkWCcV4moHB9xKYga4Cn5dfXdXXJZpoVyZ3RHBWHi4Stf14nwcW1fhfcPTBJuveq2h0QaSIrAH
SH00afFsdufOFDUquN52zhWAd7C8RTpE9iemY0A1iEkGnTsS3sfp+FTX0z4BoAwIVMxg5zp3SNjC
rS+CNaB25I8cJ1f7B7cMcaUpRxM4gxpGeCzj0kpz32sWogN6WCpIshdP7RERUz3dKlM7EAxuA9pH
ceRqRSLAG8Z2fCBvf7eA9yeYSBQ/l7U8SL2ey/6U93LLjwAF79waQqL/G0XY58m+kWHOiWs/807e
FZ4Qlyl/KdopWRLfk/F5sNBCYU2vYvAg8M/QFD/dBQKPHlkx8m3HEJbrk0y0QLQGpfEkayVF5PCY
xa0xMclM+92cviVyc3cgPmNqAVSyhaYrAJhvD5iFVFJCcH8f6bmaUsZQ7UYybpdZ6JVUd5JSMWWG
5TksqmtAQLJjRu5asOCi4QHVutREBoy5KIbNPwkot9cjJSy1ZIQy8SpiGRREevRD5yj+Id0kHb0n
ZM6+WGobVA4uD99M0eBR/OxZUyhiaKdbs93Lp38GJ8nkCS83ZuNtvBDeqY2FSmRvVpakBxIWs/gU
3mw+Ow6yj0SKFN9jBuD59YAndu7S9bZLjfXc25rf7e4uPhvhR095ilf9p8vlWp43a3M77A6AdQSo
0MaYrvgtwWmy8Nfnu3iuysQCn+QQCMdnOeyErfrI4af39PXSFWvsw2gQmASMq8rAmgZnSwXNJ/b8
Y6Ev7mFyNcF2alFB4764kurYxFRQXUZn+G5O9RImvRu6NUPn38oIozsfY7kC3wNi+A2DPOyGzK3O
TZJAHRmESKvc+WM/1G4XEVaH3DC/75SyUeIUwuGCQgSCkO7ilQ5twwc0yeG6pp1Xv87rCYkDY5ql
kxDbWrdPRrpWUP7ClgHeLAGRh+K+CjPCVq9XeH4P9Nqfz+jQxKYqS8ufdd+cqXXsJabsmwZg6471
xCeUuk4CEDpzEm/E9yN2Ir4rMjFOC40Vpm3A+Svw0Npkxog/CcAQmGMNZ8EWiurCPTubdGpb0/4d
HoGFBxieUhzgjEHfFaPokGdbTVWAAv+gwhkTIgGl/9vAcyA42+3pjqsDkqUYfO05buyiSUDEizu+
2fX7kt0Kl5jrAMyxqvbFzGbDMfV2AMDgSs7JIa9jhWP/Qc/qzq9ryYjUrCq6DMFYLqY7pqpFPyGB
+ikpwoI3ouP8vY9x4Kc4RvWzl6p/MurKNF7Vpcg0nGODgqe8wVisbdCPoQmfyaQEACftISjUt3Jh
2xADVC4/ff2UewRlDSxnkTPCYiWOBN+lCeYKK8+fHwMx01rbGMggD/Q8YAgSl+hyDp7FndsEfrDV
FXkzD43DmkkLc0N0HvdQ8FYc9UHaRKImVMBKUx8BfyiOOcebGAPLvNc19iTIWzB9gxmGa2Fknqqv
0S3ID0eolXMhjSOZGnT8Kbf0kF19Q1so/S6G/fr1dIE2ZoOf5711JyYtzjm97BbxO6nmC0yhoJIz
Wkx/KS5yfw0i18/4dMowTuH/yj5zt1UNHHOhjsXRLfe9H00AUcN7gFijwaCNz1fWdurWJn2J3TuV
V8/QKECf1i7QiuYYl1eK1IZ6YwXtedLFUCKyudNdgGw80ppOiHidcV9XaS0PQNYSE9pt8HcfJXJn
HbRhxeWrlfMBmir27PkFuwiHaishGAXD7qdLnLPEybCnIoWk7Ovo7QZ/0T8fT79Q+fNAEAVgb3DW
5IsTvKKXv41XyYnB/nVemR5LGo0NAaK8UCRmteOP/PzGwZq32gfI2OZhF0vLtH0WNLyUMP7tGAor
mogv89s6NzFeyhivUcRQH4oCwGlOH/jbX8/Z1agEIx7tgW3O5HjcU+u8KOERkTOrHwx/UmwsGnU6
u2H5glcXcJvcRWusuey/6Weg324utiHOwm9+gZmmgwYyG6gG5D+SH0sZuv2GkfmvhYOuiusjoGyg
KU+3anqh2pSQ9eZMdSKeBDtjEMF3fkQ2YsHUh8K+79YIOsutK5AGhk7VZrYmiS12wmqtno7uOlQM
ruab30OqCfnxnYcZ6HlsHHkynykRZn9AxF8PwugiRTFS9IAVN0A583KiT+f4qiKF4N8PbJUMHttt
0OzSNhhF5XpzSG3PEL1JF5WBXC453+CmpaGC/eqWntsy5TZbRrTpbXsBCmk0TrrYZey/oRZhgAAO
XTKxzK8n/7xuWNhyMut/t3wlHm/0nLsTwRlF2VgwgGd/K+uH8CN2YzomoLC/2OL20EkWhXQUvpDZ
ze4JQ50SInRxR8AIDHgepqoL/K+inffkHbUvBpXo/CFifHXEk6sGfORB2ETiVMXFKc6ejyATfPZG
AeHCgnBpAWp3SyWcEnJJ7hL/XBHiJkKYJMzw4aZgnAZOYrwhk7aWEI/vNY/g/cCEGLBRXA6qPnxc
q+J4RJjD/KdRutEMlym7goZWJLFoOtGPuPqJudjLVQmEAj1X6dqItIXNcwIlB2w0l5ANW3WI9CR6
CdwdXoqkA6KeKKZp5LhyOIR3UY7XspVdTP4NzSD2j7ozrravfW1w3JgE37lp52/FqRFJwn9TnEwH
UdzCRBRuUK05hEpAB6qvC4zCAWtAberU4sAuOeg5oJhDxuPs8EA1TqzkQ0qHb1G2QTlPWhaMbuR+
Mf0B3Fx0rpacbypxwsfHvaTBRO7aoY/cDZs72rod8WBd0zqGSmrMIfOg95oFJwLhuYSWGEHnKNXx
SbNls4nKuAGpzxY/S7Dr2VA7YgQ3JOQKvKxJoGLZRl7YqDjX3OUaXPbn30yhvxdALWsXQI8znkNZ
MFxP3+AzfuXEHa68ReP9llkp4k+DqYVgTr7CDTANx2I89hwOs0hugeZjhsEyjIkAhSYxxQj2pWck
nd/JvvXRBtJfsYjmOdeMgR/hp2+ZabRxP4Sok4fUZY1kB/OxMDIyHAhOcToZ7fjrA9+GPZtJnrDr
EhPMOQJVZJkPf9CAotz2JiwmNIZNfeUc1fso1RyeE2K+JboBfet7RpcALt/eU7gij9P4z1qInzLl
rAJVGG/Bl8jP7c9gLKtNpxNnRqMLZU4+aYrOB//luKy/G4kOQpDisyRg5euwa9591mRq0GtVyoXA
H++SWzlxIXRrFUhNcYq8r7i2NTw70l9I+nxGPEauan4rG4EoYfKH90w2/2X65OR4Zfp34TSx0sBL
eAzVld8z3rV/5gDTpaCJp01lvC6KomyLBscJY3dLVFHoMpJHt4Lm1NUhyJnBOapzyxsuOSXJCWip
uGyzfenVq18ibCpZn8+XpOYsdYRti9UvPsmkNe76C8Cg3rePE0RmlCNoUyEdqlUcKBX6MVZ2/6JK
MX04wlr/xMr+NC0BFHHOp32sXwDJOUIqG0X7qfZC8Ndm4HZRzKIBiH9pYKGcvdwxOw5bJYHx5QU0
Kfi9Eykl8do4soTtjaVPht3iGSG/s+Xd69j11ysAcGfO+315Uvgwpyp1E0IvNDlkbYMcGCrhKKmp
UbQhDD5c6lEXBo5u52F9J6W1TwpDisvOd5uIZLk0KuIXx9GhCtDGYImxpDT8mVd8GV6LrY3yidaL
Cg0zKs3cVVo+7osg5Hw1Bd4MZqqncVrZuBq9firayHpItUZfsYPsNbnfLoVCpRVvrm/Rx/8Qagcv
1032+Xr+IbnQfNnSxGRM2pwWt66hrFZbrc4hLIM85jvN7ufyQtH4mLCI4qafSMKbk4UvLi56e0np
jkzHgeOYhJDyd0mKniifcfzGCGgdwpeEeZkFIJHwkCKBIJl6b52YlOgCZHsIp1xj1QCUJNpD8Xll
/DSLd877egMYtvU6zhEpOuwQtsS69eI5QlNbQGweYY1UeQmUr+4+L2hFqbRADpj9989RrkCkrm2P
zR14s2kQgRe4eXABd8Cc5QvvBlHp+1S1BFQsMyKSU/vYdQ+5sEYq9nhtWzCEXiqckw6xvrxX1x7o
K1PPxY921g3TGj4urQNOYN662HLS/fJJFj1miF0RGurCDVNLfqAFotj356OkqmrvAYVGTF5TTy19
OWELzyXtsM33NqJE59IaPhuTmIWXhlhZaZx6RPF/pqCGnoEogSLb+lk1nk+YMjKSgJ0WI6C4iBZG
SQTBPJsUTUeg71+BjjdC/mLKBHKOfcLrBycSM5BOqUHQmKQxVU31tdfqSJ+aormoMRIHvMxeRqHx
Il5RFgPTWg7KLbePo/C71SUHv2L7N7qszGwx2AcxxqSr3BMT4mTaZMFpbrpcdp9nPAYXrSibA5aH
3Yld/diWm8KOIXrLmzlqqh4ooGeykCuINn0JujE7C5gEi19b5zb0kAXJyfiNc9jeVFNRmc+HHrJj
aeTBuXj0y9dvdSPM6RDXlOxWrGPR3t+NF1pYECNgwjQyyCVPiaMoKCTH5uf8xKpnTys3Eh04AnZz
9L97V9DEUJyRkijh/dNx6fVxtlw2/GUOuePqGNZFiA6scHIpYQ7ZMQOhk7/19iFB5JgKN1YX0JRV
0RzGorY20qO0tEaQQNY2XR8C+YuOEQDSYbMReLVJK4vWZnhOxRgHDJg0urR2q7y22e8UdPakv8Rp
nLEv5PtI/ILyFZAlxErJt70N3J3ucD4vXbyjtuwUITIJlhSVaJhYZgtI9xanQtvLatYzflbcyPuH
SCGBEUYHpbzE6pghAd7m6S0uQpYEdBnnXDGcmnAsBBprN71NypX6CuS6Md70xgMszkuxxOhkvGuF
btsuWrK165RIgh9ucOIv1cxTtREbuCWeXoyB1sKiB0IBFpyKmsE/PEMTzJtWGexNpEHKFbGaAbh2
WuUuM5OzNoDsB8CUBznFCd+l4n9NFLwx+/SqvcTC8RIGUayvN0EC4G97MfYdQpclFiASlV+VCylz
DfoJFUda+Uvr2t/3SALF/CPrf8c9APr7Ma3l8usXiBFJPxJfoTBw2/4RuwYpkuh6CpSgEVSYdOB+
s+ccstvVscPL8CPFy2efqyTzaS+eJiWNmPb6Zf44mMcx5iEMlByBluzjOtZ578/YDWN5CrQhG4lG
uHB8UxoSU9dNLC/QeX2NauxWsVT6DxgQF3KP/yj2f0+XQUEZRe1k4VBIgvM2YWkCMqu/cHSUOIQ9
c+AY6J8ztq6q6hP5PlYHvkZ0Em12pXRkibSWutJSMaiVKKBtJwDiMbhqnIP9N8n40u1UYpovFntY
kDBF0UlfqCQjmUEDxqQV/cwtoJMWm0RPkRWJmwX4Z7uxYfrCMWsOF0uiwVutEO8oORobvvLYulel
ZT/ul51/kLLUuBo6csDtgoYtAQtKB8J/p71V5hvt45RILd0Ihw+y2/Jtcv48IfkRKKNrIf9WzZZ/
Kih1h2B8s6qrepBHi7GVpmuzNgbAghxMl4ePwvL1GCMI0boBafEdVWnRQ8CZm4z3gx1npuIOTB/c
ztUk5DfcPCohK8wgS+FPXPSRayPlowLDPSM/HqYH9yv7yicewCt6+aea9nrqorwjnOwsSeiy9Qt5
iNcONR1TMIh07hFVjfLFcyNkQRQcifCseIxT8YEeCXx0mZFKLJXiesw12CyPDz4OPne0O/JzwLZS
KoS43wvpWo+eIb9Wc0lYF6Yl/BNizbf8oFmsJMjKEE4h3WKGLpFtKGKLrcPJphBVLbejZ64QMTuf
EPU20b0CQhKJYLQQ/LsrRKezDKUsUohhKA14RHFDBvjNeqHd9f1jzCh1QtsP0+LwDcXJ5uG2Q5yJ
EC4ftpltUkrpT7ozP7PCDjA1P1TSg6jyTNjm2ucPL/eWjDO3Gz0jfMlDYd2yhgeDVk9X2RUPB9G+
PZidprCSl44n87LCf6RPBv/Wz6BKojilPPl4Mx7Oz+IdLIyx3Kv5PVLxseFO1kDxgOlN2qhPoXw8
KwP0B5I6fr+qJdrXGd4sB44IWFxFNFhTd7AHR+MGNuNb0ZvOYqxwlOGcY7rkhqKsN+Y9GaUOdM0L
o5ZKLZ7GiYDPPnU15ZT7qBNfWBN2XnYqTi6LwiW86DuA/UfHdwI9tALZdoduWx0WcRrY3wblpirN
tmDt4G3Zlop22h5JqXR5+C6hb1UyYdP80RY/MxYvB6daUflyv8rj6O03T3h8pXYzG311N8BmFudh
Q/jUWLeljj7UjgVqMA6lZFD1LoiHovWT2gZOknlgO9WXxc0HB68p7Mxi6tlzXHjaCzcvPLKVdmtT
VOZSd/Fm0H+r6YpJgwLenlLLfV3uc9OQ0mTGdAVcpP3BulGb/VNYEHmti3QtGZZOdkAHSX3odQhh
8F2WVvKGq9Y9Ywn7CH16snXcZd0vdii9W1BxKcXiiFyAjW8OIpfH9bzPumBbonJFbQ0mHWCJFMJH
h3b8O0NVm95uoiucP6gCfAPj+ox0mUaXbJhjC4faaaQW+qtDixdMUf5H5ykONqLkBtkVc7DXhyKD
3IXZsuGirj1Y9SbVnxgdw4eiGS8PMhlmRfPplXmIUt7QrWsHQiVfqH0n3Se45U7iOeVngUjji79a
GwV/Dyp04kT1xfuxxG7Dx004bRBSoFd96I6hC5lva25fkcI3bllgftaQtPtjIOysRRwp5EOSd9x3
/UFHbbI4fS4oZadBMorw/Eq/X1pVp9TS5Fpr0lPMHiEjxIznWTBsASv5Cmgi65xguLdFv47TVwvq
zKA5D8juYSiCS6YrK5TIvaK6gnG6iSW0oVZENucyQv1Vdtwkv7H0PAwLw422eEDAW6d42F2gqHDw
9A3oM9bVyGQEZlU5CT/cE2jujRtEeSVnZ0WrKKPKMgot46vc08zbSpBM/qBhqLkU8qLJhYNMMDTZ
QbrNW4RVBHWwwx2vyZ0HsJN11jc8UMiHlCNwCObeKeNxE65jn+mnYusj4ffbN8RbO1fI08BX5Vx+
h6xFHaPCMqRLmNzREk9JfArGNcwsnjUv/HwUfaMji3xjsdv2P34cXWWaF7TcCeG/BID/a2e3Z3Os
CxRMGTsFJxrtFldlOXrm9UpbeYNkj3Pr5+7U0MCzK9ZEGX2d14uqV2tWO4JAPn9pApYXiofZqX8Z
23V6ELN4rHlL4zzcw/6Mn1XFDvEOu/iGg10q4ArUPspn+iDgu+Qfyt+XWxK2T8NKE/vtYpOhREKy
6Ei/NRFIJICClqlf0vgQihPXkRz3pZuxQagEyIo0S9DCaEwST2w2RQuySHCHBq7eXUbsy/iJcr2f
OjdzwbJtQ0Ctmjaodagnk9ZUAnF1pgg8vgowbrrVkOxoKVs4ixx9K5R2nuoBeZ8eXgTGYHH+h2Fq
5iWThCM4slB/vk6KIyV/9SrPx3kJA78GRthhohbk4sYDykZs0wkc2rWVB5yBoFCoXHIBq+Zii0mY
vysan4DcVUoedPirrE+LuyI7+iBTBaZ9atxTPMUrwfPuA/8NuVd7nupvDelWkUDH1KMpGdZQ9msF
NgdU/8nlqfJSaT69io6vEQbDFDrsMQLnQz6+BfwN0dBZ+s9w5knuY62j/z00T7n/MbbYiK5YlZM0
hj0d42DWEA7t5DNvd/n+/eATftt5VtBrPZCFkMKzZgtUWGnlUOJotcOTqX09mtykEO3LxtG4Ve5y
SZHSJhaKmjz+pMowyDDxOuouuMLN5McbfRSPYiRTltmqs1ZIu0csmxu16z8v5LDDWfPINjBlraNl
kYX6WuH1vttrTL8KrH5g5cvNL+HpX2LHTE80IO9y7LdBjRK62VmnJnBiwZ46L3mnVsDLp15s1wvJ
PyTj3EvEqDWyRrMWmm9ZOGz7/RynvtgFXsssp9+hRJzVLaYPEAlDYEiTQt1za7FzODv6r5tuv0ds
PFJLXtM+gR97ENjI+GnymzETljiC0JPRVzrFmR5feEJ44HNz2D6zceWnIjOJZRWj+5qHl4RBFR77
1uVhDCKRkuheqLuQkltsaGKZvKt8gWiaONEPzGZ948scoxS18lBn3I0lSNLL57asov9SsBDC9SUh
bntzRgTivWzJRZagJ0mDFrZWmtbYa78LCqDbSAyIOJJiR0KnPsKcAHxC/dUwog/Km0CqZVaB6IZw
mJRyJMFAqwe8dDplL6kHAITZN8Nfa8euoMWOjj5bva/9Eay3J3Ku0JwzlESYNS4t78f/OW39zu1H
WUoEMuhVn6R4YyyTgZE7QI3gyunkv9trUh9c358ZSl7iIHuofsgjUTMrka7o+5vLdAB65YFYdUrM
NrEBnCSmtNIO5lNHvFMvNE87EBPsIHJZsESEWeAFiLu7H5LwTUZv0WAOhiQ5KqlbyfY1gW/k//FM
Tc/Vr9khVF6vx8L+AWvc7tw+T3FD5Yk8BdUZVGlO+PVcKI7lOSj+qqygmm2PzT21Q4kgG1nqdP6j
ID7SPVHn5M92FnFFHIJJ33tB1cc00NyOqmhPRH3Ptqnr10Smere4I66ZzibjQE6reu1SIyjBVHta
4x/f3BBTvwh+sI+/U0/e5HWnnjW9887VhNfpBzvRZqSBclKzS2Lruq911HE3G65zZZULNE6iGKzo
FJ6ItOQTPIupILFNaKzyy9nzPW58YdR+a/ZvnK8wSbi9bPAE8j3unSvGam2fEq/ep6NKylPQGxMc
7ZYErDM30AjYYR4ZcRZl896FyEj7u+ST7EZ89c5CbNSjJS/jyBZJ9ZiAf1yr2wqBuit54lU2IdS6
lfh/U9Djw3zJRKVaM2QyZn4VIiZU9I9rJCsRK0FeMUPB3yP7iaj5spAQuKEAmT9qBW9CAhvTlsus
vzm4KKOvE0RfJsUysUKF0QwvuBD9/l7RYtnEj2RRiX/gLv3oMiCaL6lt8U+goNpT2/jF+CEETecB
2YICiUIGtLYg1Vga0pjCszed6exwy1H+06nLx4mET7erkQAyb/bonCtNPqXp4v13e9qHWawyGzPu
D5jR4XvLqvCMEcFEUFGajABo3YGUofWlEI33xGYwmPp0B7CVjM0PF1mf29Tbn0oilq3EbSt+lM5k
9D2U3OkxTHtqzdQmeFgDE3fdQjLa6Jdx0Pet7VdvXFoseftalq59GbZoMOF6ZNFLBJB0M06kVEz+
ByT2lKZ79cnlXOUC/TiN/Zs2rIM2hcCGTKrO1Gwkw344NLIynazklCtXuT2p7fiCGqbdNV47yd2d
YgxMMrNnXR30AVEFZIU2T7qR3ZZa7wnuJW22au2L388FxKhLOwS4d8HPt6dYfsa1jGxJapN07je5
okmmI9mVkwgL0UFRENz7Gt/gVNmAyL/uHfZ4KUBk+2GgNsxQSW2THwNB/VpS4WZnTNWy0bTU7zLY
QxQ+FEn9HCUQ8lD522pVFd2tSXTAjwtJHh0qfBLLLqw1v/wWSRLqjhzt1agKaukd7b/c7jeodAYh
SgG3t3WAt0AH12yRaDd9Zd2wEfanxNnLpFkYepvZVDPCOsYB33umV9dpawDPCaw0tHrWQLCUosUy
qV7cxAaIAnIL2qXaQrvMPim/Y3ZUuGQdi8OvyQ/o74TXzmWc78yH9xe4lqbR+d/bmbL7Qn9LjQ7x
xtFM+oNMCc7dhc7DLbBUTZI4LEpEoeng/atknh9OHRqfHRsZXSOnFYXEsEsxHvs/ov2kKIIZ1tOO
68eEZBuSA+WohB0xlwwJ7vISiYYa+31f9AvYoVHkBBRHaljr/XvjqELsSaaSArg+ykp5QityqcCW
LhC4pG8yx71dFWCX7+7kiOfKnSs2i0tAtNWUzjriV0OeESgjY3tMT8P3xx1lk8TIjKCD+ztHpS54
40UX35CxHXx52TwgnTmePhZZKOT5zyKad/QJLhi5x3Cxpu3SABjeyYZC8qa1egk5QUYYulHcEwpU
HALvj/3D/0vlTHSAHdA+ZfeO05PoLqrLpO8j2yyK7RY03IyMbtz4nJyvORXcPZugimijM9a4veoh
ndD0932AF8VvFWe6ztGl/TIzeN3Y8qwidhvNBUG65IAFETohBnkNzJzZ/noaL4qhL/sxHxB+8H1H
zx/CLabKi346kpVcQJsFynbVkBmMOl6i7C2UO+zZBfJOyBHtxNS1k+arQjww01AK+RrMRX0+g/Xk
J8mc7URL5T6D/SJTDFoim/7SivxK3o4xjyqHHHFaFD8D17lKivQh8QM2xm8nIHoONaREWQ65Umxo
AD9O6Gfwe+HTNJK6zihA5oMET6rUef3xeaoqmsiFrVcyeIjD1kwdUjdlje6TKMgnl0gGTBARMCN/
rXI493HL7CrmduiWs0isA74WnD0peq4tk/a7zz/Q/EcSfjbBQg285RHWTfUdJfO3MoO0jqfRNFMv
e7NJb2BZQjaZ+/wteMivgll4a6vhaYHMIFYJR+0athPoZUl2010ZcfBmwC5spRPT2mx39gXBFiuc
PbSo+/PkLXtf0hqLe1FDTy3gKDxXMBVpUPttMHv1wYnlaP8yLbGDHu4CxKl/ZTR7WCcxI+akpPMY
Rr+NB2bcpNMsFoCzaH/kQVqIPxnPx1jpoU3dnBDq19cNBLqHuwxW4C90O1F8lkbo5xurujo6s/dh
0HhmyrM6M/xLO/cq2u7pzaFyYbBJHW7aLX92biHzhPAa5vFFRbAlWx57FGPhNg+OC8t3IPWmxu1u
8p/T+sM9fsPpUonDGEowTauIQa9QELjALh5jh5Jlj7Kzek3+E2Nnvpv2T0sr+479+vqXrjFxLM13
xqBeKudvbJOZDDDl9r/oXZ6c9u/3tFoMEy8y9AUkNUApnTqxt1FWP0NjPZAsiIcVdfySlRAy6hyA
Gow105+7qOKACZXPJ2IF9YHl+7tClI0ki80W1Z969r1T4P7xjjF/CLVv+Z+KDMvARKwRIaPaVHOy
e2mbR57ReAIPVnql32qlNoQogY6BiycqUMm8ZYaEzTrKoTQQlSoAKjh8wW/ffH4Q72v23HSf/mRF
jEfk3d7StDEDXsUx6zpk2dtU+fP4wuyaVvKoNuwe0+ehXE8kkRV6gF7PfLyIFuPivRDyWre1E1Ad
1xz6/ODdoy86bFJd8beKUPaQ8VJwvJZttMopKZfz2o6fJbsDrmEpFAWBJC/CNiqxBh3/UTNJF5xj
g/IhcZejWnAaPJTwfXprO60/HigTwP5h4Uh5fe6mIxrAFmxeDrvPHhTVdZcDyxeqnEA4wxslWxjV
fBsEpKXIejzN8wqpg4s/TahKivKx8L6WUiu+BJyz/AvAvtlNhU4rA46g00HVTheY7Wzx7OXtDg6W
et0XpRsvc7XwT5l3BvnGFW6QVEjgAwBINELc/AWrKDmKfLbmeqW4p2U0uoysNUgQNAiFsixDBn6U
LOgJZaw+NnX/WpOjH6pomVsDTkGh44tYMyUZ1zw5CZa3xTM7HBGtHtMQUYbblIUYvowvzDwIrEEA
3LcqTTCp1sRxPsBKM3b2uwwYBtoBmtrLz5OO719kcxHtwceu4iMNBCewP8EB4HDbr32/Yk2nEZLL
dTpmKU0CYljPKGPPOKKYPRraVUSfCd4mRAxXqdc76KU9Vo6pyyWbMF5HXwiW0BYtsSIgncQTpFOC
phTe1g85Fzb0aTcfoTQMwL0Dp3HQU9l7lzN5MTNINX42bt5I3LUJlx2Hx4H77iktwVYtnzN+RjWV
NAPA1MYoGRGZPSWcXSI66+Fox4r9F+gRZF/Gl15SQ2cfeMXtGN3NsATqgt4gjmv4WSJcBfcSBBhn
vDb6xmBLUJlF3jktVxrIx64/moQYg5BUQ1drc0k+HpRCvkmOLpSsQw3XW1Yb1qh5HMQ67escf94J
7rscp3Ax2hlzVi+4NuFEiIEtpq+XGRW1glQY6EBpSm09NjPjH1W7wb6c6dziVoC73/rahaMY0svt
dOvQ9/IA0hDy6LOS6y1eDgTRvr7Ad/j/rMq2VPmPOhYdT8+FskrMAG18MWlrobE7lb3zhdNQYkA8
iSAkZqp1waObbSzgvcHY47WS6SvhYXg00tEKbhFH5oqqNMTW4EGEJSGjOvpQEzKDZQ22o54k+/AM
AI/9mcU/x3nLaA05TCWJRtFZGBA2OeKhQPRTROihCt/z+jMREHddd5hCYkg+802ALXmtd1wG1ij5
MlG8t0XXi/4CJBPlVt+JvX1MOsNBK6npbdKLOMukRFlJQJzs3dLeXNagSBMWcYJUF/CWOLPks/bx
L41TRYdLE4ydIdH1nWFo1kR8yc87I+Z5JnD4/ZrnM4QRWN7YLW8IEcC0JkkpZ90coCQ5tT5sZXlI
l2oKNjE2HRL/A0/sjpBud5nJyMJ2JC6v/fcm0/w5IPcaFOpIcXlIdgjWH9MKzSas4X2tJJdoB3Sf
ipltH4DhwkpzbZIdWln+Ok1BFcwPejYMdQoOjwjdmjB3Y2w2UATLbyeQK5xx3NtfFc4BfjJ//+I5
XmsmU/QWkOr1YkrW1pkKhakkuX6tclOppTA24wu0CB/iao8NP06g7DVPHE0cTzQn38CZucuV6QD4
ptIav40/ftUw+69E9EMGSaZWacowiKOv2kvVs+phmEkwrGcPR6qnzVvJ6OJbblNSDZLYKLejVQd5
qVinaCXyp0y8804NMyx9/tFYm20VYScEcr+P0+crhHoc15Kuks00EQKBRpPtyN1INDhc/FMW8wki
G4L9gmQC0uHStNxtkxvb13FPqFS/IxHNZhDEWbYEx/J5EjEK8kzl4O5gnPcyUSV/pl90TGiTdRGp
U/cle889lfi4h1ea7URliQ+t9b/uSbyUGoYaMufEUNsn3Fr8iY5YFkdVWlwa/H8XDF89j+x4o5/p
YLcNcJKvVdhXuRqa+23dOoF9EKSfb2SGg7MH69HE1at/5Ca+t6pktlw4+UHAvEslb5EbdfrBk7c2
rOPCd3fKozuXZpRja+ylpRRqagduepTuumAyUPOM605rkQhhCkT5BCiYkRGkuuZNL6yNKPQbHheH
VkrFC/YoJgDr9urcR5WyVfAUAcrwVGzp7wvQOEAiNc1gr69TpRR4hjYTZkH6oz81/ATjfZWTj/X9
hkJbB0fhk60K7Y7hdjyh5eq5KAI4kK12hc6RLbiuAb+Wen95393OGk7Ek1kNnrxKg2OtnLMeb7ls
gGe83h5FqwDeUjy9xJ6U3x1KPoFRtnrOerw6nZzDpY13T1/D/N6rP0wy/RsNClND2G8eg0Q9repK
+zI5vTaQ6Is6XXJ8i00sbzj+ZBRvSzD881d2m+x7hhaY7Tq9KgFVca0h4Cv77R65am8GEK/EVWPa
nYZMYbXh6/KNowNxfhSD8rg0SWnp1x2GVjnJOCKDpkdrXy++SywDR8Qe606/DFn6IU0MVyhQiLj1
7lwfCzfh2xYF3pHyDEWmlFa+wvJ6jBjtPusG4qP9qzR3E76pvvTUKanLfMfe+UbRlZ28hHUxtVUE
RPpYLio9RvS36miXt0yMIWpeQJTSWZtkGUgpXwquDl/wFs6XWeXlYp/UkD0xgfU13NnG6iZ3aAfm
auqssQTE6a1xe5jLYlokCQxGqPI0EI7d297lx5XI/p6MAIoxaso8GFP2vIPzSZ3TkoLT1ykWueIx
usgYZAHrBo03Zmx2WNtLoAJY/Xn0Ltp0HCP+P+TLOj1mfn/I6tlyIDZuc4rKn1I8qdX4uZ93HAJA
Tcgckbu8kBv6MvNaEX141Xriyo0PXy/JjPiNqGDIKVwj1bZ/FvLWrKsq5PKaNVq7LHD9f182yxeU
t0m8lSeEdxJzhzbPcWf86iUQ2VAVdyt6KV7pwjnsOXw5FgCjoGq0fK1Midxfi/2no9ETj52uiwdL
kmqtof2Mm5gR7/N9i6mTQdetLgF/0VFZ1dLg7hqpZoxRS1f3d3AP6nRzn2QdaTNUClwPw+jZ8HKu
5tk+gI/7GOITzLvvNt29kHZdCoILRg8dy9z3wtQX/QZprL7rbuTMeiggfZb+oQ+RPJoQyslMSf+Q
1aIDblXz43fumX9arYVQO4Kn5y1UcYr9VekhWzkDwZEReWpaFBwhFChPUiXSfPnw4SLkqLLs0faM
oH4oZfk69jB4Jl1S/D+80AhIJTFWSKh0uUz6I8PnrF6TKCpL0NKG3r1Y4f/Ssqj7YOdFCZl7T1u5
Sa3AbX28LKfpSjipTXYvam/OLzz2ZSmoJsUSJlGXs8iwPsGij/1vDm0or9zNas4EbS6qJl4pQGmo
MQ/cibuwDCpFlcr1vr3umqIX+lTH1xsoPZ5KQwm3593k7MakEgcBj0VJ5ScNQOkMbDO35C2MdU5Z
CpCeIydr/FADdgVQO+QJCnhZG/+0bg/tAEd06XyemubwO3kiTcohXGSA1eCHfEpSdpNSIl+f0our
mhYGgfcG8P3acEpoS0zNp46QB5Onijlldi/BB2OiVzQRTPrjphGVhJy6iMO7wPfEOmI7uwA+kGVP
9hKGt4yRLiOnioKAhhZMPQu1pxpgNDfay71Sw0tzu1tkhWGa7NhPjw89q8CADUo0YXQ8ChA1E7Kc
9u86TvQvLW4jwTLha0O/UjfUAcVcG/wF9n8OCBD9KAYGiF3Nb7WwJKum0n2lwDJ/ExUdPuJyP+D5
hY+KwOgdHP/dBPc0MZXIQ0NFU+jV3kyW8yLu8HoI04soF2jFOItLylFlKxX2BwTuTCd2ivROUsxk
JkFG4G4NdREDvbgyHoTG5gUcMd9Ruh4H7IbD28MqaXL9l0V2oMt5XGDd8VMrC0yu5peZdOkNZqFK
+EERW3bWjdX6AyBtA/7VbO0qxf/EkXJvgaBPHJFLxx8Gzlw3KoABcguJL/5V6EmipVw/M6H+syB5
Gp1LDqgjdutTvzz9Q0a/8fjSKufeOIWPMZXimGYEwdEaXLpxr46jHPFungAELBI3MCwPVOPvNg0Z
tVzrZEsYw/Rjy87Aheax2dxXETVNFGrNQuujU2MUkL1csPgZz8EmYae0/r25gW7DL19t9BHjGWEP
Dy23H9nXA7ELIJAHxOC6WsAgAFX6KkMNLQIyn9zynD7xprPqQyDWtIeUxPfb6Bobto6tWOff2eZp
rW/It79CgN7HWjpN4bHgLWsWyBg4gkM0nAlDT/47e8f7Xda+mWQaMZiyhkHdWLl2GxrY1lvzM/OX
j0VWwsZDSiV1txHdIfY7YdIRD8Xew7TwnK3ESb1IqbYt5VhYgzfLoZsyVGkGLpxysmXr0AAFU9C6
8I6WKrhPy1GDb0VM6p3Ot0FhXM03CHx0c4tn2vi700HYkRgFUhpvTFWX0pFSjeCvZRpKe1enLK+X
PfSmRt/wTs0/6oj7Sn22dNaKK7EIob42FJ+xw7xDbSO3jM/L6v4snlyYjnkUk1rV2NRklxZSdPYo
7x4c9JWo8fUUrNObLdRYusfI3DGZtfMlJsloP2YgKkNyGxOGqiBKHseMruj1RKkpYWTGRCFLlwX+
83Fw4tmzk3ZTV4TUE6ybFnXbV3mbFHGUwUnkw79FsDjkqHdApe6O3WTQo+m8WQt91cG80E3+Gd7p
uKIeWZb3aGS9LVuBsYEL0MPty6dUM0DQpO0t3FrAQKjlqyjstWiZSATMpUcJKskteH7Vm9VipRRp
V2G55sQdWevaXHHIegXLe49YKTJqJxrJKAufp2q3koj5EbaQ/e3bCdujQWq5ImMzCUgtT4tDcPbH
sMuv0E28E2nhiloyxm9Eif39LC0N/ytlD5Wy0kuefROQ4ulp3rHXmxzfDnDce+JHp75bofxMXrEh
oSSPOusy2ncoRh7bWeHu30Bpq4D1DmeudgDbbETGWLelIDkx9MI6+jQZeyMLB01NM6jdFuZJGsi+
jF2T6EPTf2sZTqpH2XrwJhRpmJAtHcit/WI4ZMcFpmsdaG9jYmfhpcOagpjN47EYJ4dLAaSTPMk/
fY8wMFi5L8EmWTTpGx7dU8JeBhP3sV8MutPIl+EqZt2vGwzULh97iOM0arRu2RPWY7xnOZUAq6FG
lXfy1ryNpMnT4nHMDovyUlJYrb0AlBcr3XlalIu8HPQ8U1FuIumgapGU1vwmdTNAot23FMS+0IWL
Xgm4KNzC+njpjf1AGfYog6eagbclDTqGIpqkN6HalNbw/5FhyEVNqvH7U+X2SmK7rG9SGS9/Dm35
pW/EmFep+g/flQdoikcTtcPTeV6ZWKBy1CLhe9yvcST9S0QQUTHab0KExMFtaIRams7iwFcH8B+a
/bZAnbCWv7OHF8QRyytmkeNFYd/3/JhkxPm+tLBad+QN0T8loruthCbEMBkCzLzYZwva3x07W60W
0lLBalsdn3e35y+dCQcR80SbYN9woFxAoI+xPFfF678sEKl8DaKJcQzgxDVf02B4QnB35JoTxTNl
Wow6YPtV8OaRocMn1O4NgcehXjXKVBbsom5usLcW/03A9//vFkX6viMMyiy9WBj/HEssvbed2rv7
zPkm7bATeJh1ZsU7MWMpnd1TEXxJ9oVAWdAz90zX8K3NJ8lWMMunfmKHbiwjI0Kuh3j8R1RKZrN7
WhtWlBAJNPPK56IaN1sHNjXZUsh+knhOdCfbPwR8ISLAGZA7eYeUm9VvzaJxoZ6eyRif99hJ93ZB
2u2z7o8sM4cnJTZT3933wc7T4VtAeldtTgS6D6xmRQLnRrWnr7Jf1X3fgP2ayi6uQ+mt47km+XVZ
/goakE3aJ04CY9CIwmoTEiL98sR05wQeKJLjZi8wa4oa3sKaQ9Wxy0JIkmmHuEhjUyLsqpxgpomi
AfJTGCyFsubgprGwJTE9IiVdgw19B8QIf+ska5W17gab7A0NdI2Gf2iGdCYuxO0Xjpv5N8slw3NT
0lJZc0MvDL3SojMECpixEiCuhU7ERRONVTMD5rxXzMHuISbGG3JO9Rwcj3NWRz6ZM8lyc5MVusbg
7ndvQx0WshXPqitYjbo4OOLoRCXkH8Bn3+uYRkZ7XuaGzyGe3gaQRH1+P4INtq4NjB5FjQN79wX4
d6trbu1S7UYstEjxhIj6ck28R+0OhS49HlN7C/WordwtS9ZBmai/roOesve6rtB+RQRcClTFGiKd
59/ME7Ot7MPwsrR8V8WNn/bV9v5A+i1Dy05WC9c96H59/l3knIX+Ryvvw/eqXblmhvh2WQzAfZWO
2ZzBhS6O6ygFmXAbDa5IHXsCN/K5vOT3RFCmztPsRLSncSw5kro24Yx6SOJ3U17uNUMRIKiUK2g1
nUQxHndk001yYsN0RLYeDSK4Eh8fcIOnnUeFH1URO0yPeSaLKto2C/WGabGJBdqAb6OqPbDlad+8
lbG+R+I4Zi97PRcwr5zbsbvqfBpphMF1XwqzCtDI12xpnMjDnq2ZsuSHN9Cv/Pwb/UFqtcvS0EYq
KdavrGZ0swYF6734eLimu7qQ1G32gLtnVdpBXx8h0/xQzDg7IeF8KQHYJw7aZyWPKlR0ybIO9Iey
jHDPSj5CTA+AptvLaMm2cRxeOLq3mdVpJTX0jj+2c8HgCv/EB/gpyTUeI3tj5T86Gy643lIs6Cbn
X8nz05t7pVzsEnRXCfnRlL0KYk3GEMNHDU3Fp+R60z8cdnrVDuqta0JopZcL09+o8Km7zIMeyjXL
Q/s9BHgaJodUMYFI5g2spji6WMi3NQ0rdbT00fGjNhNGgPXscGgIWdnEXjjvbptAoi12iBBziY2M
H6uGgcrFBCv5l2HfIl9qji1uyELMOsTmQiRMc/TyeAdcT6OSAPXp6hcSy4h5Pv6+YyW2VKc2wjT/
ALay1lIAik7ye9+gY4uGMZlnE9f9d+SE4TV1knnaa/vs4fWwpu8ftJ6FvvabksnzPvrit4dHUPYJ
mVaVw+6C9KxHf8YMwB7QN5QPm7RcCWtsEdDRTb/uFrE3vSN02h5bh7UV2SRagn4KMrQtJO1BFv3w
xaHkYCUqoem45T1ZZp6A9Y0ELCbnYOiKOElJj35rUgOX2UI3IrK4PzqHMRS/YqJxmPLhzxV9Ine8
b43r9mgehW9933wyDKKRlWnerIB1jpROAlFefaj3Klmo4JvVYWWw1PvMpnwuK5WwbUOsvovJitlj
wR5BHPAbEMSmfvT+sWjk+7DsE06OToIld7rRIOFqhE62cCs0e81vsvKCMze4FmeJtJnZq6CrUtkv
9xVbbHEWp8sSXQ9qxr6ZqRifLB7Co6BSNmUFzoxVfBLvSsBOsJTOYkCYVcwpYjnQGLLpWReT8ngO
3rGcDAznjD4kHhfykMclHjOqu8/odT7rG5NujA3wVmw9RcZ8KsxISK54TP5S2+wIDzaOCiHllUcE
nEsIOD5Zg0Ixq0ObnK/qdmyEDwcjibHEbQWyM5Du7iPAdHFR2aXI9+KtULnaui62MOEP402GtRzO
lqHb60kTPi6XUhIIbBj15+43+7es+PMNnDxZVKGi0ArJZTGdu2md03MRaRRbBSVdFFVeEo5GdyYM
p3QdSERQ+9zg9YYcpOnu1CtEiO9zWIR9cJRMPq8Jiu+1YaMz4nJIPP43cxZ3fkEWlww+W1/76bRK
ei/IeMair1WrpFa16SnBdMcwoBzyoImtjRo8F5f8KZ83xPH87VRp+m5yLzjoARMhRM2NuVoi46Vz
IYFwNppqHij1MXybDLlSJJsbctjVrTEnS9OIipUkf5Q2tOG0WnpJC2Duqt38JZPff/hlzJ9SfR99
Sg2t/QCNxCoNDnKdYJsPF7w7cQU9HaFHcOJGcv/TBlje/6Sf9GEFVlXDlcy5nptx9Xlx4Rv9/W07
yymp3rvgUF/VL0Tozwy3MFhF7JMKEHDCMvVz8wDqj8EBtdUOpFhNuaqycKtHXOEw3lvHXZe7SLpx
qUbOovsan0hrGlCZy230IeAv/TaPZDx/GyuSkAGMQIpm/2DS8GXlVFlok1OG8TXRdpAMfe1i/Lxy
bH9fFS5ZyKJXgX8NyWy2ZQu6wACE+U39vc3nk9hZ7kk/UhZI0t3tsnQYIvuWFvB0f4H7DkrTlJR/
Cqkh2O8QpXUm0Vmk+B86WmTFX5KZqyb+y4bWsuYCQBOI7F3HqHcXLgxIYgr/ATYQYv7AXGsP0+e3
Y7UFzaAf+X0xIMp2v+IYuaYA1PYavkAquMIK8c/tuHzXOLbbKWcPK8XfxDH0cgFUBtWs/iTX0UKb
3/5qgmaZB5pWPRSxy0n9DfW9qnIbNS6NQd8f08FTVaSPTtb57yg+ofC0nlJ5IDzN9gUbXqchrP8+
FBCB5TwiuBseMhKCf8gsIn3AfBncBvaG7Vu6ykEDiJB4vMLrjoV3gLv6UihvqcA/ktaSkc4ewSLp
ThDCL2+hNwX4swY7i7RQVgagQgCzXXHhdw+cwI4+iR3WdjvjTsNp23PXjThKBd75PbofjPF51HvC
XOul6tZEVrPm70zV4dgL6znmQnbKKcT2okCL+HxZy3ZRNBPinSQFn5r379ziYsMkIsmGLqNazBHP
AmlLpPa+NN3V0eTWkPugC7OvT8IY9ZdcUfAc9Y0VA7M7a5ibv9wq+81Ygj+RkHjpGvU62pON9239
YEqVji/AAzHLSk0X8i3rsPCxrZSsDp2+1k759C5GsJiAnzFYR0N/DxNfDRQ6n8+EUIRAVDbxeFsq
L+scEQR78bPO5XgV7ydcQKX0RhX0di7A9x8ya66f8SphMlJ4bTaWr+lzgPFGqacAWVq2gaWKDwsY
7OhyXGiDJv2Vc7dvwNsovTPy66ZGkAHzmQKiLBXf74Dl4g1lrAq0QL6koFp5W0IqQW1c9OcM/f9X
lK0ZFJwhzkm3FDNiAZo+JNtYHuVpXc3jSQy8e/6YR5tYUKZOwQGVNY4c54ftiNN+YYv5sh3qblwa
0LE0423F8vwiQR1PJje8uiQkCCSPDgaxjFP9k9cO567Aj5yl1LGXK4EKEkxbgyrpcGuCLlXj9r1g
hQ8pqd2A8yRetPFWWphgqxB39l35T6U69w650SJYfMRFhleD4dJlxJ1yuh3jG07H0bNRno8PjHM8
/SDtL7XgBy8g5Tq4/Bp3Ko12mAvM3Ztws1lpAfva0t8SLNF3gVWLC5XdJ+lfJDo+Vmsr4N4REak7
R4DlHtjxfqpnZnQC81/ivGPdtyVd3mfvJ/tav/VVgZnoNK5hNjbSXP85Xq9a0RwR8Zb9GpyKnRvr
gNf5WgXOsjWeU14vVwufV2zVRLDQGOLGkgcGhXY648GNKggqm0SMnLfVvD/d1/zMKYgG42PfEF5N
PFhXgAwq2MU/Ka2kS6AkutlOw407cQtPcUugv4FdE2L5HBqruHPCaq6XLvT2pxnCkKYVNgciaIsI
ge79iYt75EqZze9RSC4qHrjMGCcJvY2Lg+dpKR9m4MDnM9LCsenMWh0K3NTAv8FeWV+9O04cVmyy
guZMV0hfF67+CDiElla/+zMCOFTNad1wdhHfCg6W7F63sZJp5b1ghHaWqU2WS+to6DXzf77QLlAm
PNSQ0x5oGK74NHyGFluFEU5sABY1gNoYRiTSLKIxNcTNjYrkPxzlTTt+c+gCeabsAUjZd48afBVd
h/dKFpIpxa/nn2BYbH/qnD1uEDvZS4dxA4XsXNC78yoTwXNmxrs/vgng+HZ1lUb+r9SWgV0Dv9Rs
QulZ9nL++he1aIfD1BqBI96Yi1jM3RFiTpQtq+p3Cj9MONrXl7NNmfU0b4tif6C32wxuq0yld2+W
FHebfK3UzXCX2O1mQjY9E+vo/Q9wPLQ9LAzLE94X4BDrc8z5oaYSN6n2v5hDJFloVdKSlLF0vax1
gVK/Tsbx5KxvBP6tmkecZbrKBpqL/wQwq6KugyH+lfvocYOnSRJPVciNYLFQhoY03oo3cwIcP5xc
IkDYZVMdF23h6soUExBk6Fo1bEpW2yCqV5AQhtfAqjuWR0HRLwBRlD1kLbRBcJXsYJ6ox0KP7zAX
rJMBx94G/aeJsbI8WbnKvu216p7im+i/VTe7t3Bv2LOTmem+KPMi86Q/wmn1k2i/hSFa7xdSgxFu
2Z6mq1uFCf5Z9TZCPmdEYJA9qSCi4D+ZZ6Jf7lQARsGB2mDpIG3e25O+wYBAXJ9Zr35KeQDdWn8O
qog/KpBfObg0pdmfd85NFmqjECEtolij+knOqwJ9/G4MiV8Allq8zG38RGI7mVdJOUhApxn+TU5A
1z9jX0O60aECIPGK0bbexFQIdI/isjdQzHJ3iLf1YsRcHA4/EcD9b2In8YET0k5GRajxelpEKqRg
R9SxykvYEFTrQDlnzKrlkPI58r92IJY/aYCSbQxtfvhyudhgOqJGW3OH4w1INdA1aqiooTvAQQPU
bnG86XevrAFZ6Gjh0fH5Ma0u9JJTHf1uNmtGcEhlxZUIDx2yC9httiYQIv0n1e2UWjeHRodpBjEw
RJ6hfDk13HTMLy/10LMnKqJZQLL/nWZFZpHdXJG4zzLs03Qvnezhw1R2hmmdXj+/iocpcZFayoTO
/FwMLy0V+PjYc9EUZd+ZT3PwkkQxfD8eE0BMKFeoeIfQj717v24tRLhEGbduc3W4aavEch6tD1p8
Umu4T2GQBYIirgVcS2qpZUR/ljwYhj7AyfaNeS/AaOzIZrkOYDHPmfBHPmyP2HETNLoex6edGmtG
UQOSNolFgGajkE5sEk5pW5NkMdZhO7/QILk7iPTZKqw0yIkzelt79GAeAnp+yJmvfddg80Stmenx
ujhex+qtXELrQFfflaTjE90X6gMgMf7SGlH9a5eQJQ3y7CkH8QASil9+hbMB+7mb/s5T0SydXRKI
Xu9yApD/jmFFJaY+rT8Vv7q2fXiBlTNRw/VUrk+PJ71F0pQAFv7n+qenUMU/bQNQRg4lKQtj1dI7
42Le2F5HWVLMs0lF9TaoiTxjxeX3+Q6BoOsNrtzFb2+wRVc3P3m1+S3obxCFMqStkJQ3kGs0nCKn
TYB3lZSsNrMhUA1D6j5TkCWJ2+Ym8R/eOum3GV30GitFoob34Neg8PRQC8RHXQ2Vfd6GU64J5lY3
hjjh5JHMasjrAXFkC4ZdxIFNwI/qY8UX72ZXedf8FPlaBYVsAsMJ+5KCK994zr84X2r62DdJcSmv
Z4Zu2l3KN0elzdvtZHgrixbzvG5CIXTKe6E3iUs6+NQRlQNbJPKcczTAdpHQYNig+PAnaVu7qRYE
hKB0ZTBF8AtvkcG3jOgBsWhHvtG/3j+XGXwfXyq+KDtRBX5A5eVj3sapGz2ZLKFl07ab5IDjxrCf
WuLQ98LNYmqF7xURzR2TGA2KgrO01dbWNJKxquPylk9z41Sf4+qcFq9av7WS8ViNUTiKpOPeOunZ
LtDeXeTWpntFZQB//RISB7MZkf4l3HSKWd/3I5LxvJGtT5UMSImzhHSUvfKTXu27KqIDU2OYVQXC
VtHD8ve7BGpyDp0fCAG21zc1JnYautrrI7zNaC8pOy3pAdos1VPQidEdfkhP/XcAjpFBNQH8ZAPW
0254OpXKsXm9ftWWwsP5J0C307kq0juHHOzbYWRBrJuQ5CBLtB4n+KWOX9ZQOH5AgZDgFea+vhmr
wY9+fngQu5dUWNmFyPZjkj95nlqS3SOuoDBywcjZ+UYnb0RjR3VShdPX6ggClhq7sAwe/5qDa0v4
abbCLMPsN2KMlYkGXFtKqa+9tKJA6bJaAkApHKIkZ4l1n1R6Sd0j5XZ/WC8RGWBAJMk6tbNRbJPS
Gd0blpDFYSdQ756YUQcxo+Z4q1574S45kE5xiLh/aRf05HR39pZtKM2N9+z2sZAuPPd7W/RFkh4K
nMbd7qax1shY1KF/0aDKSfapqAkaWkWQ0e3KfITF31U8MfkzPMUqyxT4uR2QiCDN24d7weVZYeVe
2BqJbSDCoa5tajwf+3zOAjiM78TsaCNh0fZ5eMJaNoffWHIxHMAYi8tSnft4E5f+qxz5LaKInz9j
PyuBU0gt0J4zUGeB/TZtvfJ9UDS0m3fVMs6+VRB0TGiv/5z/lVLT1viXUrVG5SfuMDt7Q0zfd4Vp
mcCGki43YkhdbnNyYVLxR1hPeEn9YmieTgAySGfzySN/D04bVOXqaEpP08o9RaVdwa46UKZ38U6E
6ZFjmXhg31+mLr9yDXIsFJXY4f7NtKM/3Lt0pOkf+8kXp+XGDYdp7rwlDjQlmOzXQevMurldW6NI
vlR5Mhgr/kVsv/g2w0lJUF1HpOyKCiARB46hBuAIwCcC6xF4MUsfIGoaPQGCOQCKmYj42+kDEvmM
msvDHa6M/sKJgAfly8afIyakMl1PrL8X4m5YitL6V+c8VUbA7EJABdxVDhfGVfeahSP5Y2Xrgfga
Ebzpz7YQ649lnoP8rektISVU82hEqre/zdBeenuVRyhBvSFabDN3R7El2ANa0+92tE9ZMRxD/kZ9
29mvF56T4Oa1xFAqD91tUnQD/ClkSaaFgoA7S6j7lG21JS0RivbqSOFCx8QgVWN33Pn2NYwpSGxo
Fpg2RTXhTrJ2TIpiRHkyVzmA4ZAJKtx7lByEmcCA1ApcPn2w2BCspHwNuhEnxrpf4EVWlTNcypNA
6fFTCBs3UJCtdqKmkyakWhE11gOEmXVKR35Cys3QueksbkJA/PCGpevZzbAKD6NnDBig4rn0Yooc
qpdqtR3p8ZZnUEgGHCOhnxDUnkaGBcfQ3Hukd7iYH2DEVvLLzmsTLGU3n+AQ6k6aplr5ahxOhJO7
/fmYMk31oIYS2g7JbeO8sJ59H/4pKdLfJ0H8+tFr2FwXXV+UBBijkvNzUx5NFgGV1sLvJ1SZInCb
s1Zxa8m5YsAPua/gQwcFJyM7zwo0OSgr9sct7xkU2VzSWBXioHBNWcATu9f4HJE4WUt4YYWnIzRq
4agjIDZXG9q6pD4RRsaD2/4UL0zPMOjrztthjiVkM3wrRcuIrRsIGFo1mLhXLUqrj/2IlKIr6xKW
c7wPkUGPVs72fPG+oAiCFS0INvhshCHSZ1ER0xFklo5DK2rGFngsRIN59TFdL583c5G7GVj/FJb+
yFC/UXlW4QOw6UiofR0H0S18FUdH3l8pVMNxiKTigi1HEvpOl7kvMUObsAPnVWukO6MNFtykzcLx
e14YASmFeOiTOL9QrzgrwfYoOfcSf+KWIz/7RCHS+AuauION90v+p3Pq1ROg6VOnjoFAWm16UhxX
rB0jhpredHr/eA2VmYEiE2XctELNZPR08arPX+rXDrjHmFPTkbyNjKXajx96jpV62bnFmcawwWkf
MTikWfAG2pC0HOQT5/2KDeVkmgKR9gcKUIMEaFQxVQ3i+4zje7RHIv8ScgwnsiSTIczfJmTQwgP7
Rdcl6lX6gZx4aL4Ane2VQyavFMPkl6erqqo127RO8CGRcqt8z90VhElY3jophn8wIIL8MZKV1ABu
6fqKQJb/D3RYIk1U0ExNio8qlOOueEkvi9Ura9jFKGRxTBKAHYp/CW5vB4FDcMzaYIwc/nCYDqRJ
I+99MPb0H8Jht8XzIwjkCELZV4rNj5YwSyjS+HHvjqSxM4zDvy6ztV4VpGqOGmJR9wY3BYhnpMx2
QLBr3wp43gtglP6PWx4d4oIOJircrNILJ0nMbWMbaiViP1a3vo3QBNKd5Tk8PozLtXbQN+q4bH4q
j3R/9XENsR2z0meCIiN51oByyZ56mVUh1kwygd+b8gWfF+0vU01BYqQIKkPLT6224Zv+hlRu5kdZ
zcQrJp2oKCjJAK6nrafKPwH79pmlfS63IDPQB/mzkT8CeofXOGGvkD3pLAHe77e8aCXq005w0VTF
5ZRQ34OHA0EWg3akXsUTYMCgYJPBiqWO4LAzQ9lhVIb4Bx5foe9Hbps4agI+KnRDEIm39fTjmJCx
HZuGtvFEScMOlyK0ifhiR0kQtHwaHodPaGXoi6qGGVx5xcQHil6Yrp/hhvw99bzuyCvDqix4/cB8
r5VorGY6ECYYOnTxHZf3EqTJsi+0/fehVfg3XILertXDhIOnUf7knKkEy2MdBq/PrVqKkjVKqdlK
n8Ji4DG5yT2Fu/KUZdcRTaQz8V3diSt+n8MiixJmW9X3cifIupN1hxVC2oi+oqGxY6h0FTYOo2f7
5uYwGoQGKLEjFptu60iKaMXRtmwJaED6Zrl37aPmIma3FUFa1yBaTGnwfg/I81itpdLVhOeuRLVk
zvSPMH2NPJVTiIlEAwZEpqwAq4zuHZd7wbPX7RjIysYsXgdW3oniG1xkY7nLnY6L9+AzBXd8ZJFw
7FlBEyOb3+9mOG2CuFLYEt4sm8YHhldVZ/Z3gpQqBV+FzgBLTIj49e1lcPNYbr7Ymm/ZQqVVIrvA
5Zy28EhX+y3OLN5qOOy7rk/heYC7y3bmSFgiqLXnzU8TOIw0G321auBHD8LnxH27ksQYt8CqllW/
km3VfnXrPNA8cBH8i4zynFwCfKK73OOK4bawdK3LHijZ5frz+ITnOO40dPeaaXsvSQRWGbegatJ7
c2yCjMd8l0ad48AF1etphHeSuHcmcLUH9JuuFpNa/qP2Oy4G0v/qAPBZuLzz2RNX+A2Qzf1IXPmg
4+ZjlGERl4F23sJwwMJjUxL47A/jKuLUwNJjfPHNVrsJAtRWmKWg/FItwFFXYQMwTMVUWJ7NDILA
E+TPyuNN8bj+2CMuCNXNuEazdbBfb3OgI1/JWt4F783giFOMXaX9OVRJ8ehxEbfQqy07WYYF3E5P
+Et/13Q6iKKJKxyFO++Wc1WAhk7OGB8nRYGjpypetsU3XNKv6YX3ZeK9ekODMsIsByIKkpKNyN9G
Iny7StPNO7lQvXfV7H7rDkRl2iitqjavXtgEJVAvGwm0rH/ioYcIfJQE5p8kvwjUan7KHtYaIR5f
APyNt91YQDDdWXX5n+B0y/2xu6jbWQQQ5zPBnDINrkNam/APEEoUw3XCo7yP6MPTmzOQFBpI8pZY
p5hR678AYzZ65H5PhcxNs3iDSQOgbeq1DM+Irbn+6v99wi8ZQFuuVxoWLBnWuWxIe49Ykk470d1v
iJZ/1ib93bdjvn4kqY77ngwEgPBOfSQBgREyFw3s8P5Z3qJo7HbQQ2ugBfIO3MDPTv+d4iRIK3QZ
zXIFvPZOkXhcrAiln++KHKarQur2YVxhchWY/kD+bY/qnC+of57iSlo9gUV8zzOgYehdYz3kzPeb
D7ZtN2Aj362YKZ0jEIt7jFuIGMMBoZITFPAWvUGywVmH0rGhv4/YWA64ObC4CkK1s+L2331KXEXP
S1wazjE4e2cA1ue40hhPKmyzcnO301PtrB3tZLgOW3hUGSae0z5OOyUj3r2zb949ttUp5sl+9kSN
A762knraawnp/CR8QOje7jtngamtcG8DAvNvpdqLxrxd+vAj0jEB04eigEVD/4pdY89EHzXj++Ua
H50VtaUNg9PHFP4yn2vg5FskBCNxBdAJ+EQl/sGWXz2WzD5um+P7vPE5kiEo2xxzAcYlp/V8QJQX
L7tbTunCAoDFWGZSDNh5/GupKTookukDCy8mkJ3ZFyeYLD5NhYOU+ELUOThum2jPKEDLWwDp05jm
gLrtUMlDiuRKlPaQIuc9qSoPtA2mJkxna0hB407pw/T4aEKO00u5d2eywbMVLz0Ii6kHUcdNV+d4
kdzEiJTQ1MPmhzEAR4YVfq893BKqHgc99E0JFqnoYcwpYYQSfPUAxndTzuuK30vfNmBq+YJZvdwk
KnjQzDaTh3HpV164mXjOiKl9ZGrvMF2r6iE4l9VG6LhHFWg4PL/oMSG0oxmzMz/D0tzMZVOVYBg8
z1woGZObWvUR9iWWplDClpALCNIyXCQEHqSwImX+V8OYg8GkSX3W44wSmeu6m/3+3bocjodOEmno
mIf1vNvUCyqOXEjvBrYpPTCtRE8bqSdAypzTMWD0nmq7GvKoFjvGSjyB7cPvXUG+8XRP+GYacanR
MANT7GBEgTWn+u9fLze4mC0XR8DCRT9ysKGGvFhQ4zQAwGfqvNihDnmLQHZWMNGfYkg3NSv5J5RN
vbdBSnYkyyp7pHVClmAeSKPajjWeq2p8XHlCT4I77dx0hulKnBAfJ5vWZAutkZfVxFRwr6aaupGF
1cycSffNJNk2MrY2xiFwXaAfUJknwQIN8lXE/mMKmCZAbXy37T172u/9ChMGEFLJ9oyAIlkkT0xG
XAp9rsYFomG4yzXsxQbClbsaE30ZBZr+P2anWRdpt4lEoqoHqriP5Pnx22oEMoIA6U4NuDHEhzZD
qKR5p6VSi8m28cvVqsqq3eHDdDHZdlasbkl18no3klG7xKQnUnRas2I6GR3QsStrQuj5zN8Oige3
5Gi7XENdne64RhQNlnRt4FYNDZGyislNIZCr+ML6lFTEKHRTXS9Fay6kstyprn2s/NJFh5XuGnKf
sTipa0xLiwXJVBjY9AHWxmsF4YW91QnHxNU0Wc6MR5EOXnfx7fAC/YVqLaGYZZ4beeOL6VSyOLwj
73peAjX3U8Spg/jnkkrz6YeFbJyItWwQ3ns3qEEeD4oMPsXmxJ48uUOmPxqtxgDhVqR12lsKFNjk
epBdvLOF7HeW+Un+3Q1L6G5ZJT5SV9q1Yqvhe9EZ1zhXCWC5cR2aWaOZRj1usz9ydRfYi1asqOZx
bt60HELoo4rNGyolYPJokWv4hHphVrcZS+uWGnt4xZd2RGe5KILq0hzjipEw8fcGZODbjHFCK9nH
wViVVdwcwS6MDAXQuPU68PLYlnLCIWRG5fgrgDhe/GGyWFNHyIab/bitJtLuGOGVldYsdr/J4fui
oOYFy2UlNvEyoOP53KMcn/I7TJHsm14Q09UsSVYNNt1973dkOK+j/i/06mA7bZ0vj66yBAwqL+Wg
z/hGcaEg4pUGyWttXQeegT/STitdXCiqJIb0V/rrgvHuV8tLskwAkYvoEpT2HLf1j5NFM8BbYq4+
qGozRgiCbpdZNhTnukgJLIcp1AWmEtC9cZbYOkCWpMz2GBn0Kbp6m6FOLGts7RvHQ/N53VEGNU0l
KmBPDyFoIR7l5F6RLBEPKTj1288ZsNRpPxff0mqm1Jq5KjD5z8FOi5UPRIbMZBF1q9kmg5/QhazO
Rm+DIVtrHqro3Vf3AvCE3b6W0IvKpvbGKM03y76qRLtUlYW9TMk14/v5rY/c4jq/EbKDOmH/pHHm
WO+PuKl/F462ZA2u7Wtj74wfK7EsF4laZQ3n3LVBI/o1E34/ALBTsrVzO8WYk7CHp+aFd3NP6iM1
uC7btpbo1d6FQqkOjmjq5aV7jHmztWR4sQCkOZ++27L9fz7KCHAZg4yomxS0EJYw+jWsYb2OKRus
wQ0ZYNuxBGYV1VPCSfJFribl4cojekH1aLYcd2VCUZK77HxnzAgNBRaNZ3SsKdKMFlMXgjJuTaYp
P1IOyQpwfKeB3P+deohzdpkhLe19s8XoxnPPDHxxI0UihKQP+bOxRrhpzy2Ea6cord1oRE+NWvDv
KHucaXL1w1Y11mcb1wEnvfKa1SmE8sSa5M6qkq5Qh6HxeKd2iv80MXZSTbhW3QxIp3mJRglxbRrc
mHaGgVCfh0oessNaqMykMn9y0f7AKCfa42QuKqaeuzlwUydja4oYWejPEhhLFUh0g6SoqjPiWmAR
Vda9tzTGrzDDlyqKuRtWiVRDRzw+9F/mtFYAxqzF7/tryQ9Y4raZMykZa6hLInJtWJXhzd2Sc6Yx
xziu+x7h+Ba8BDZcJrML80MMxbL6HZ/8LHVXP0fzU9X00ViC2dffX5HKYRSZd1hhA0lCAlQDmTZL
kT1J9XKyaFUe0nLjmjsf6rHndxNUOgNI8gFOxYqrgbtM/wrLri5fv15fD6mhV5L51YAX4OSWt0ij
tfGR8KtO26h3eD5kVixX+sL7/zhY2ffTFn/aXb/T+2ICo+Aw1KiRYLb11NbtS2q5riMhlxwZ8bTt
Jts4+Cs58vC5CQZpASiUHkggjqeXuWtvnOaXUspbYD3I7suH4Diz8k/UlgQPfnqP1qsqedu5kWjj
hfhEljoUXih87YHoBPf1Pc+ejG79j0iwwWBl1FftbJtuUQfhtRHfJPv7qtXRSdQGB7p/8gowdRWS
wL5GjBJy/IIUDXpDsieaemLHS67sjlA6lVsJSO+jrOUTNR3tBm/KCiKB3kdP3nN7tLF84epQYsxx
banpPpOg48zUgbkQx+PObaRm+eXYFUXqrghCqZVRd3N66fptQgm4KHjnxND9LYovir+/tfCq8ETZ
QwcSuQ16d+Q1NMO3PChecP7DN8/0OQC+SnMiYojl7VgycUDkxofWghdtbwCq7sWj643FAR/R7pPZ
oKm0KfB10UNnKCLi5t4Bs4ZgBRsTwRPznsCzZUwxziLVhhW+fm92IIY3WgFdqLtpPq+ik+YJXEw3
Sog4L0kpMUmJktvQbS/W4p6fcqGzygkHGaa6xWHijvaImRKeGPimwRnk3QMgN+/KW/bDxeCPXcsK
lQwHePNd8dKqVqvdEtiySskIv7DPNXqh2zM9JGuW1qIKL+aDX9RTU15jiysGET9jPhRom3/X5cM7
G3+nVRizOwDycshz0qyXN0R5UfZapXl+iKmDt4UazhidSAsev9RdAt2B1YMYDzr7i6vITtUbPX+R
9zXEdTLkgbxA9rN40+yAWgDzK3GuoSzy7OBABuic07QNeghape4gOt6b3PCwp6lJtwqj5Idc7Z55
JBJIaIXTAbBfMlJ3AFvMHJJUE7OUgtZNyankvYh0fWDAgJvVtJH+jxlri9XnwB4N63bZ4yYNnen9
NTApH52kEXuPFNa7ZuCyPcvkROVqkahKM40DpoGofXhFqjEGspHwVIG2US/cN0j0eaJvETZdtVaf
6D+dlmRBUORiKR+SKPhNghRusiv1YJWUl3M/INa1oIMOhENE8KtZLDJdbtmYSPbU1/Ym2c8sYTbC
foWbGUu5+HKGSV9/sQEfnCsNLl3jFJNp8wN2bM4q76DLt6DXT7bkpt4NP4a7gc0LInnKnHbAx7zb
U3sHfoWT9rXPEsvWaLZQIIEUqPUwVimDyYasxoGqBAyww/jdm4/sFSfX9o6UCVf/3b1D12hUH/af
0hfJFs9bik0iSVwNi598d4W3R/GOjb+BouQJJD9qus1LWYJrxxk8Yc+RGiqtsr9+N//DHMJ299AQ
/nrIM26CKJstW/vNuAWmghHjvXQ65P7dHCws3MYy2tbistjJ8cR87PW4dX6BDrj8py2yJFd6e2G7
1mfVi62+bEecfK7Mk1SU0wJJch+17fW8ecY/1SEc64U8ldMIqgloDeHCMnwSaIWS+iiEjO1uwOW3
YWFRNn612xrLdeP3H1S0QEiXZRpYzjRpaFeWaM3oztNgggqxatrjzWICM532LPV7ON1kaqGU5BUG
u28HaMM/WkpdWSUbzoaFJI+a+PAaq2ypyEl+rEQQLxAwBTLTVnFovw0sWlrwdnZWFhJP5MRx41FB
qTMwYZEI5LTzPtoSkUHIkMKndjIbi+jQBQJeX0ElYm721dYH2+2fFc1KA3omi6nIoTPAmlhQvUmN
sjw1NJoGOxTcOhTCTE/mK+AhCYruiNd3guWn1UnkL6V3wE3jNOngV9mXaFdhqqRnWOuRkfItlk42
oe2jHrTn/s0sDApAPKo6Apv7/bP0N9jHK4hTbV8fIMo2rs6z9YVTOw7KiHZPOP8RzIwrRuk4WYKl
xEPgrvm2EXAMemHu0AmefI0loaKw1bR1cfYKmU0wSEJeEmsCEsX4Iay19ePd6x8AlAZIDXA3siai
mySkvtXkqxn6ajxTMkKWwQF7dyo+abgF3ybghTkrlk+e99jkF+nrQ9mqmWtQrmhXli/5uHey39NB
GxE0ksXBJtbVxrtqoZ6QY9c8pJdO9yPmbnOPwOtPiCVvs5fYpAzEWrK5PjF2ppdA0sZtnCK4B3M3
Mvmj1B6uIyhbUOfSDoGRKZXMuBaqnFj3qib9W20RPJuACbnAb23iyIeEO8IRg0xxoT7XsCWMDew9
anogitvOt1Sji27n0bnH9fIh+7mBliwane+7BYFAEKztp1B5JriumfQaEuImpCDPwtVp/jA+I3aZ
mkADK372gDySC5yaiIpATmr1aZp+XIHeS+QQmKgKEnBJycWXZcA8YZHBWnSOdIUtHop1v+tjySSw
DL1kOQOF7Gf/YCUS8lTCau7i8jScaxNxVsOImSeqFU8yLFtOzA+Irx7z+jeHCvrDmpZD3lVj9ZVM
ofBNdVpmkeLOG1YU2GRsXGjxN5q8/o/MNFiEMpap/eNWPFhsc5mEy0sNhlqXEagZvjxsUcHOMrDY
AczFMQ18YjBwg9e7Gh+8QaZXIjrchMr3L7CBBQJYnQP8TezDRzQa1bXd2VSFmH4LvJ7gMOjaTqsM
bt9bTL/kQD/8TB2zoIM3ukB5xaHV5ncShPIG5PnvINH+pg/sfq9u7YwDGr6Tm2qU78WJ3s+dw8Dn
rRlOLUVA0eWCjdjORr5l6BRPdl1AA6UdTz4yRPy90SuKmO/ybjfJArZffijZVHjmNHyJSXv2ZD63
iCViNsnCSbaQtaFerczENQ+pRK9Hbl51O5eCIOQt8Hxw1Pc816nWR1Kq3FgRQInso+nVgrfAARJ5
Q1z6rQ2kr/IjyVtqt59XVgE292Km2yPx9LRkUf0G8S6OYalm7UvONRQCB7jHAHMJGnVhu0Ql/mha
geTjBw0ZmQ+Dh03WBASSj+3a0SDHzLPa5CkKv75LnIcMhU2tBQgL44udVRO/a8V8/I755V/gC92E
QYhOKprfPc6ltv1I1Y6fhal+hEBE3mnUczuMODWpfzaoi1yOuGXTixGqKlvCIRmq8hRRgfgrm3Dw
bb06+7mEVN6yKERulZgymDZVccqcvUoal0tx6wdjEj1VsrujGutEcRTAlF96nbn1LkwJGZ8CkJHq
qcY3CCK3ARF4hHyLoZ+KlmLAPhBq+AXePRASzq5bjoH4dXJiSm1Oy8i+OP0sPap0mgo4mgSv665A
ho+RaN+PhFH5y0Dp2pbVFXmZoKwjvdqoiKoQo/EpYsQlNovr7sgWgISaX/xB2d1jubRb18RmeDQJ
Z79hprvkyy8HFreyztfXbtQ+oG7QtXCfnPowPdn/WCuu/8vHg6aDYjVc+VYfXMyUOjU0AkGQDv24
s52xO0tL/XocMz9QL+J40vzGUOwm/kXjY1b4eE7GxteihrBuvcVtHPJAh/YUPum11r9Ird+BaPrp
evk/jV7Bu99zRIz3egANqxprnweM7xY+xiqqheDW9EOkzakLtqFIqk7QJD0iAc83h513eikPA4xr
MYTDW/mJYrG7myCP3gGswLEgCuYvl1wWAX+cMFLOYKw6lNKae/xzBoIVMcG+WRw1J1Or+sk7fcMB
JACPweIP7m2p6HtN6KAUlkmMWVqIxYLSZseuSqwBNjH4DVPQt4+QE+KuO/ULb/55BpeM6sz55E6s
Cn7wFlNmEhaceHA9ewr4pBafO6ZScS3y3g3hWXQbBmeBcauT9qdkmg5ZhAEeRKfy/3XJDRvXznuh
j872Uyl1Vw+hqOxPlpv0/cDeqVl2kl3FEXF10Jb5F61g95zV69TSYdq9Cfg439kyfgq+hEWwvNNa
EUGi2oCG+6v3Lo/7V/edcPxIR+65JuWigi0cjAaaNq1RAJcRbNNzbFlXV6LA6fKBm2kcLqTMgjiW
GYm6KKJ1v9PVvmc/0Dl/e8iZRjFLSRNKN85EDQqi5uuIZ69gGcY/+MBqwMQJzfyvbCNNruloIaQH
0ftfZThThgg7I+VeWgQXMXPjmAkVf8NlVtCEGIeZJtLxfq1Xd12zfHnIWBlZgySk83BTBafFhHpT
pli/7aMtThMtcjeW729klCJl3hQuU5TyNW+gYjWFX4uYSmelIvII9TXYSgz4Ag1TqHAHvt9AQaGQ
FYuzjGsY63ZMzKtjewJJ8CvVYtWrPXX+F74cE5mQXo2oJAG3vzx3znwbzNtVQeND41WbK7SZr9GJ
f+CndF6tR/7xYaeqyVBVqMxLkmlDkM7IbAZQQEb7MjkndA6wXX3lxpmA3bwUWkHzA+PYwl/eFqvp
fO1BR+z+feyZrErMrQvFLocfboagsCE0g4uXJg+2MeXc3Fa+3mAvtjJLG6/FlYof05UbeQqiqxzx
x1ZQV2jynJ5WrTsBu4swUVLM1/pOMONzsGduFQFVGkRG6TELnhnNH6XTG7locwPnRluN1ojjBekB
m6Z6GRrpQznwKSaxumE7Sqw8jRbbQtpRoMxPo/0ZhpyZLaZp/vwS8tZ98xOyaMD8x4YQOdkTqBEp
ho3sQfkyNiQoQaE7Ho4/XMIM3xs01BhHMZ+BzxAAZ5BTU3vpm9G3v4gwJjtz3lovKO4Uk7kKhIHl
AevJ1jN6sVYRK6ZUhGx+N6bRTna9zBrEfoI1p2LTJr1mJGPAqzKJuQAl8VPuYHKsY+DgtvpgNVH+
UMKzXbDqUdvVjDjijCO2XPhuXgdkADLUAJ8qqiVQ4qM7x7SVAsI1LKMIO+9LzvH6dOfkQ579EhV5
npi3b8dMhKEfA6C1Tw8ZQNs8fD1Vurd01Fn7WaKP34zavbJWxQ+oMQ4r8ap3G5I/uKeIz6jsfIMg
32uDmsjQT3cRaqpRXfpa2IfStcC8p/rky68fnGYh/wDIawjM3DW3HhhtiNFw97vou1Nl/t7u9fgR
1Q8AzARcvirxmww2nVZHxb4GiPT8d+tDOZbQv6JZxubih6t8YrUhvw09ghXJ5LA89E14L+upnHO6
irDH5mDBUjsbYPR80XEnBOTKgvZoSF6xQy4IdtS+8x/pM7coFXWE2/71JJeTjP246mTT5TesNov2
eXOQznSK5R/iNzq3bVxzJGQgTaIWuVN3Uk2MS14JRfubqeGPj2rObkeCjfNtkHtgbFaN27e7J/Wx
JfT8zBBxGfmZb9EUW+8WxdVnIAQY5XAD9VINIrNaZkcKFtw/L3KpK+82Sv9llzSMfe6MZ+FLaU8N
qABrgpOn1MJAeDroltVGdtdZzu/yKyqZpKgDMBp9iGlpq/ZTk9cvaeKIzgtc/j39Ankkr0RpmUgL
idjGYwRnXqUD3TQznS68W7fS4naGSNfI5HFHZlLo+byEDyvWbkNYsa9Xgabit7JfajFyUjtARk4P
Tun6Q6dlIySR7/2FgP8KGwAJJIklxi5eODk4v+fzMJ63ddMXoY6iPOqZJ1oGEae2pO+11CS76TeM
xrfw5Ecy5+Fw7HdMqNL1Sf36ajawyRhHzX8762TppN5whBzxS8YbX2FO3DUbiVf8b3kVrzrYKSqp
rAZ8QedxbJBbfbmwcxKIjMm6rQQ4VP5D31yAz2LlBIYG5DeqhTvZe8xZGR4hHEhPnK9ECRdc/u5N
XTob+TYU3MQ0Vn2DvL/UyrxFIKRM0KiUtvXeIpYSDZNdFxlWPmVBO31JuA6pGnT9KSzWwWSoCU/f
bkn7sMRjPebVdW/Mf4P3zfnFP71Crn2zk5JAiGEiEaQ3XXhl57y9YTaE4L7sJte9J9/X4FqLmueJ
U1BJRiOsdOKs7qicxG2gbgZJP1ivUR0/Z9nF/iT6tINI6gmreG10x9+r7bIOWV5M+YmDkup69etB
ecryLmEy/LVczIAv59L04txcDibT9TSGsdY2UN9EZVQyW0FadYjW5dtZpeIsqHADfZblgl6L78dC
9wsNVV2Eye74wYoUuldY2OzwtCivQ+NtewWhV+OUuse8dxo41wDHYoRfwcqUut0yqgKSUKnzEb/b
YzZYHEfByIZlrFysotSPONaPhcDHelXfNZyTGat2bJvr0cwvmBO1HygQwY84U5G6K0t75Gly8l8a
fz0WGFrnDsWn0PzJ9NKZcS+y3uPv7u7nToGSjCeLQ76mzGmgIjtsqpa51dNyV3SYOZ+8gz2V88Ft
tXG9VAiCVrdUxWiKWf8+6GrVsXI6eKrcvUnD2FWc7oKDbqQfqFOL1Ci0GF3QdEHUt2uBFrj/a2Bm
UIaHhoJdpVooyjkFMJGrtxwoemEEIiZKKi5Q4o8VRXILbBw6IZgu77WOpimlNMI0gPSkhynWem84
IhMEredVeC4wb6wNOHC6Pyr3HJydUvUZIg/ZUL+4McrhEYf7a5nCDm96hunervhVxufhz/fX9lQV
8b/zrbEyHIfvwtwfqYQOOdfUb13Ys7HEY3MkOEIsYleMue42RyXZetHBQyF0aHYwXAi3AuORe14c
XM0YVjRsPm4tesiEf2vdrt4nQbleNkzYzs0eHokWw3B3+rFKw+wbp3+gHx+A6YqDy/zzA9t+yvYq
/0hqLsadAhCF1VWQisFpqs7UNymP3UCe5JLPOSLLkIwykXh2tXKH1jiCiRcYNFMMERSoPZKC3+EJ
+9QwR3rDsv+YmGQMl0WCfXqodIrY6cbTFh9IuTddKNU8X2vz04kB4XY+xaxzNKKvT5Gx6mB1kGF0
UzVOex3Gz/Z4fQi8zUy4OphogYVeKezoCBfT4ewF3qbkCnb4hwscSSOtxQRD+hiuHkg9hI6OMzM1
M6gbdMWF9GJ51z1r9lgE1oiECEr8goyT5nJKF14IRDGJrokVXjkSkoUgHD0g5FCdzA1AjUSwaKyI
Cs8oRqWe56Gx9VlSEr2CE1jKVdSfNnHJ74HxZYR09zMwMuA5TKxnNBZvJNy4NMa2vlzKLAxdE9hM
5ujuLzdm0UtnM+bku2mBaUyNF3Vw6M48QLq65RRs660jRaP0++NgsiH55d+N45jacLP22qy5sT/A
gHkvuKgGQuosfuhzyWHZdL4xUMLbTIHeMtZiE+3YforLedX027WbVDy8qekkk0JXQRvyFBksNNW+
UHHdQymu6ISflSAA4DB3zFcTlhGOY4pE4tkVdjx6SQSaPqp5MHYIPL++qjTpYEOEd4UBaDKCfixb
eqf8p8tNL7uYgaV8+cMqmao7TLBwmi6CqOKV/W7WclxLDorJiuJhKXpNnTMAUCtbZGsNt39wG18I
UJYasxDpyFb9PzrN50P+s189KFgOeB4ZGF9mHbyG8WxTiQ4Ju4f/YnqKnz25poN19Ih2MtEXLkjC
Ftz5D6a4H3+n4cPzs81bg9/LG5aKVFZwW8WKcwvnrAm7H4qFaKT4Guaq5EPBGoA/8xqib2DgRTUa
7F1kMOUX3ZEuE3x/APJdIpct75FA3IRXmHCP2RXV/zRijKeTLub1zsGgebAcrlR5EM8dgZG0/rko
LBXPTl6XUVkBrquJy78Cdp3LIFfp0XrC8sw9M2TgFB3/NioskoUuyiqRqO+ypqcydrK+msMovOom
mSPMFH4y+jdZ2JcJIpJLXlCe6N0u8UDcnCrItP5vjxztdxW+XAj8vYMj3yQc9h/y88rSOoom4319
qscugMv9HTEI/t/nX9IFN33CvF/Ky233MdYcYfstlAbnlsy9vs1KL07JfyDiJa2ZGNY37dczdUH1
o3vrtHT+15p1TEBwZVY7LMFC2jKKadW7RkQM6UNFN56E0WnMzJtK11myfMvVthdo/O7LPml4y/W1
RgQAx/KMMk4A3mioZgz1AfsWDn2/1K8b5LvxWTRaBA/KjG6+5Syw/Avbf/95Ph8s73w/OIQFNvqU
vZT4MB7btOxQygfveqLKPwGwpiCJE3jQ9fJiTzCX+0zdwx9UEZfkVbrGGqRZI24qrdsv2GaH5FaS
OirsYRacMcolhFRv9zucyoBCWLHRQsk+nhVjussGpvufZsFB5LHzacrsnyD2PgMi+1jEAJWr5vAW
ev3VVNlSRnWx4pAuckzSjWNI8C6rxqU7E/IUjy3Scgmo1WREf8f3boORnU4WCibQYP1YbZqwkmRT
HZuvPCaMilRcLTZ969hC8UhNMVvF3xwuFTcqGnOhUXxiaLuRGtQUsr+0E1/ZxamCJXyFIZJkNU8F
iKusGXhOSJxGE+VNxBdKPYbtRcNIpzwoCj+cZjmZB1JOyho7hIP/ltdch4ORmu67a5AnTNDKAE7b
uU77fKWJnqJmx/JWbcA1WRUfVCSI9643mh6c8GigsiqETBv9m/91i9mDOADpy2WckaVmHqWorqzC
oa5b92mFJ26eBKBwxxgh4vi81V7xu64TervHolA8qDjFXGetiIsJEzNKERk/RNqbF51UscRg+Sk2
dBEycUr9GxzpoiFg6IUvh5r2TIZB0iKns71A12tZRdNPTjkOIWZYsYyYTJ91ya3vCE4R0cBgNbtz
rgt5I920DMrwS833r1hho/i69HkAWZs6tihXMU1fccY8/9/0Zg8JXtj4gpdzgUaMIBZgwf6p9HOq
NHYVoCaM5hsHqAhibmL6VEJ1/G5hTKf+CkktEsbMx+QiICHM3ww6FPO1WgiIKnyVb8OjTwDtdSaw
jWGs3EyJY4CLC31Cfr1ePwQEBZDQgd41hh7eUJpCNm6w9kLB4ldZN4yjQfFudxnUHQNUE1jqG8DS
wS7hKoKNfSHXSn1tS15FbjqgjMZ76tu8cZ+BknRxg+kXh80hLfULSFYg9x/4TsKnV47j0wjYwTCa
OvcPhXU90ihV/WwFj8t1RqoRhARh99FeFNfLVsiOafO9k62kzjVBDIHkfV3FVQ7Ubnl7NJYLSwxV
fVHselADNnLlQEqi9ojo1YJH5jWjL64BeVViL2rUY5Lk4sdcMEXIWWCtcQErXMH/oSmAT4Lr9CDl
KtTf9oHgWvy6QNfGY7WvRNzjbBOUNvzmUbctq4BFrFzcC6hdsXn8OFbY60yhnA+/a5qdP4bu6Ie/
J4vfBfhfldGnF6xXu9avs08svuzRffuzolsu9tZ96Ip7i0R44aG3I7DTi3RmP3f6gjy6bR0D8rOT
wN0XreTd5NtJ1boagP7BG3GxJxvjOOIdQ6QTnW/3BLTgJm/zF8vAqmpjj1ZMp5TqCfq4QfdYIOc5
wdGrWI8QyvPXOVoyFBSEypsEs/dx9vg7HNV4KLvKVrVY+iqNGa/AQ1fDV1Mn0y7ozKGo7fMksLHj
0Xw5wDPDrjbIlcyqGOJ69NUlrAY/pvVEYQQhGXgGhkHBSl5OqwYniG0Tr+YS66oYDq5C2VznlgyK
H1L4DvZn1Un4VntuRU1c80ZxE2WFST1wdXXZmD1TzuOr16OhNFtG1N33M4jhjG48b96eeCGcmETe
9UpH1o/7feCcZN148udxpnExwltyziXNAbioZgSt0e8vb4lrsCKWG7+CFQOa+EtrjqOZl389T7Aw
J02RgFKSEyMi9J0GOY1xo6drvzjXzFAZAidOl75F83hUAsgeol06PW27CsCx1ekbUdfmDUD/AgSq
27LMR1KwU2oqPCRdbzsRr0ogY20ktc4dU+Gcp1x5nIMDtsRk8/yu9XMyUxAq9kekD0AB7LhnN0p+
3ZURFr6qZ3e8d91qnkXXK9renAtxubDUB3NRR7jYfmWm5JgC/8JSoAUPb3mwTqra/r0p7wljhBaU
gALabq6dxlGDfQa9OU3DIcOK39skcouVlBEEmMCSKc15Rzf/W3AabQuibDNGtzIcyIv1WRRPR6uc
rNjRc2QA7l1B/p/f94i9f5v/0TxkSiiIeej6Dc8C+Kwl3ZxrpgHSbRwXVc4euckq9j8gG5dMTV7S
7kWhme9quADUAtnvGyx+q1GLH95AxCOJmP5WH3GEbOe9+cLfE4gJkXkLGdgZVi0aFfraP9BUPfje
2K7Yl4qMawLa22pDXkZLA64lcjp4D4umwy9xnUbb5qB5Tw+INTsN+82lDNIi0kXosCHV9dSwbOZP
QEF+Txm+tPcFVgY2FPDVW91o3vycnfADC/uTOyHO/lIgFPbxgzsUB3WlRwdGdDEmE45nIxjRa+bb
1DE6qMt7okPoMGFNNj4xlFyfOP5kEMJu1gV6F/PO/kCZz0Oj/60kvudhHIEPyodQoD4UdbLPE/Jp
nv/drAYmqxxnBirk60+mov9ix5kkmhqi9ac+dHNzpr8QBnsBtkyBmn9cmAP1HWtrTPKjKGE/uZpC
Qfrh5TcpgtP24G1QHjA1zso2XfVAy5GJsSMnZNFBrqoIHLSIeDHeOkOtzL/gCH+cbouYD0dqsMkk
D8+8aYDQ+qnDM6gBDwF/hfdMs8vhmLRaTeuWOKh4+YqsFYTFdtmm49tk/4pwbum6sUHyUo9pEtt9
tXHMWNM+ZoiB8ew5WxTqzWfTG0IK+A16yZ5UFvGilI+XnDWmf2WiWhqxdjN4gNKVftBAYN2sl3Z2
Audk0BCrMiPzhMgu47WCzwb3QRorLSBEqWqt3FYfIpAHBd1BrdTT+TG5rrw37fKfOcYxsEbqaMkc
+P+q7X7TfcQNMqNqc2C1RCwA7O9NcP1C/z0NQukamoYbtqPWvTacpZF9XhykPlPpbsisiosm2Lpf
opLTAewJrY8n6dq1J4XjfeW+OPwTNAWJH7rMmq8t5mKbQJA1qjwcHkEeiou/ifnowlWqoqLp7jM0
GT7wVmP1HovtmXIYbpVz3239St8e6AuZHCmbBsB7DB28HeYDn+tCFdw8C+BmdfiUDTluopm+uhFZ
aOmNG9Gl9DqUjKhARY1LeBX/oKS67iXj14IDptDXoF2J4No2VofTogeocHQDKd1gRIwltIV7VWGX
agtCcLdKjC84FvQr5gjN85VPJtYtJJ1njGx4IhBg2vp0/dTGTih3DvzUqDDzNeidWdszQQBpTii9
vFwTMk38I2J7OmVeFgBU8F2s1ZeVSW7ngHWx9vhWRiHjztOgUmi3gsRNmqF3TA7ThUucDWITMfvq
q+PnOT7WmWTFSE099fqlJAC7iPXmSkdXUolS7JsUvJOEXiEePEi3swGtGUd0d+rpOjK0g0gYEo69
IcT4FpbC8Cr1IZne0hkIEOuwnzF3ndybM1exl2gbC+zZFl3WWWW/qAQr3Z0se+m1/QA78U9qmQPE
W65/Y956L2htF0LIglXv2xu/vobgrOAt0KV+6z3aaIExOFZlJopiTcTwnYbqDRCYrBT6P/j97sON
LMCHOs/OoLO2/Gxk3OKfVx7SOztvVXHcFOGzuBxjGx31E2THFqk8HnuJSXTA49xyeAZMx0Zncgjp
bro/CJWiuMtMoxkNClc2+QIrSY6BzLKO53LAo5F4l0NAJzppqNltPaSUtx9MeMfB1ri1bBozg4sL
UdmVWV1GjPWBLxTLm2GzbD8I7qxpJTvIMqbrFf0zDTpgFDiUkEdp0B4WQy91wndM9Vfw79G/irbl
Rgru2jf2Zb9gk4guN2bkqLMZrSHp07MVmFrZlfnOFfNnShZQjkHcIsUSajWpx/t1CjoPguPR8fsu
lCT9JzhCWVjbkqMOT93PBmW7wfUCVJO2nW7sIFy/aTgMjXcj8HcUwQmSLahIclKfScA8a4BID2GX
LTQCuJ9AXcGqwop4H+mo8u+qqa7MBQnjru4Zf4kTATa6hh/IGaO0dbV0a3zHEpguiqv+if7zL8rj
LAucBQLuH1xaKx5hWzQdbO015aJco7svPbRMxpOllQhCUBYti162wCsYZjI89Wu0tBlC2xBiSCq+
sJ2Sda+wYNULmNbkPvxISaAg3NRBKPGTSfmZT+JVOPNSoUUbVfdh/0rKI6nOguyiso9yue7BkbW0
a5jHcveihWMHyCAurM+wqoEYGgEf/iT6qN2eGYq8VuxPS4rAUfw4bN9J0mDCrGWPgbWLCJPa8lUU
eg6lRLKoSgKqaLjOE5AzXQf2wtbvON47VCUemedIuXukcZwNwD0WGyPnVBTKn/a9LjA0Dezm71he
OG2TxjO+O0mq84+YEjdnPMpwLuSyYEO7mPOhSKbSEKyt9i69uJMd5XbxiKRmDeV5OZMFZFUUeZ/M
pe2RYF2dNQ6wk+/sUkLW4PV+kS42Wln1v1kSJF9jXk2ZdRH1WwIz7Vqfmy/lj4JtfqUpJgGFuT1H
pG20iR/83qbPsMg1sCwlHpkEfJkuIP5F7cCPXUBK2mZ0yPQreGbGsLYmBf7O9jckulIECeMiOMTd
o+/Pnmw8zWm3WDUAXArlnWqw6Z0OR4Z2MJEH+taa1Cn+DMZIjqEJYV9K4++vILjuII4WludeRqja
Lb4JtbiaFNsS/Cq7JGSKRRKpKpqNRgkmuh82EAfXqHt0CbKCn8eZvQhrMXkrifbr58f51uOYQqTv
lCvdJFaUCefqZWnF2hru/9MjjMu+m0zayc96EdHSbcvQsY3uUEQNsWwzN2PVUGmvtICCaCPISahn
dpf0vIJj9J4LbuzDKlhVVYxYDT4RB2qtUF3xv8Zk7fHuVfyPhM1yKnvbuFm/QxQeHohcMmK2hIZJ
pCx+bghdK5+EqgobE2FXTp4CR4G24p8v0Rn10gMBY/XjrFOqQOMxLTH0Xy05iZOUL6nsLwXjhXA2
1TlfXnBI8HnjEo6jgFkb4yu4a9clj/4BHGeqTw/u/0DsRGNQ7ZMz
`protect end_protected
