��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}��,d�)q�n'a�s�0~��N��C{�OƪR�)��K����Ņ������6+��˗5���#
��	�Wl�x��LZ���=K�r�bH�����[r�u���b������9׋8� �$&W�JU�+~ T�~���M6(���W*��FC�:�6Ɇ��]\7����,x�&w�gx�}�&��&֎Ղ�6���L��t�pA�4z؇�}��T�ny����M���;��$�ͤ���Z03T@��@n�=a�C��B<"����-S�uI&�>�z� \��T�'�xO��?+R���i��n�T��� �xLV���f'�&��h?� �8sഽZ17�i�����	��8��)K���B�w��Z�#V���/�{b�Z���*�uc�(g��w �R�3d�,n�8+!zI���w �̽ ��I�M@c�Y�\b��U�[��?��������4�u���z֩����;f�:��S�89�֙�lJ�h��.zU^<�x��_��i�i���#	o/�ʛ����.�n8e�+�����]�'�n�)�bp��G1&>d#L��?+�ی�z�-����n��>�^���;�!A�R(�Yz'���/`����`P���ߚ�	��$�C��Ԗ�Y�}�:*�Zd��B��-�B���wf����ş��0�)�Up�y�؊z��9���^�J�Y�:�e->_U��]�\����3�U0�k���̇�������!d�žY+ �SN��B��^f�	"~V�>&�?�$�Bku���glYHDd�T���3	�t���8��?9I�niin�I�k8<%�sؒ4�r�L�_�v�<�"��Nd&��+⎙��2�.�h���5vL H"�\�u�5�>�T*Ħ��џ�u>g6c�x妺��f�=��La�)�O�)9����]��0ms�g�xH��DhH)orM	����V!�I��N(p������&��8wP�5
�Zd.n�}�k5��>ⴁh��X0 ��y|F06V|fox\i�U��>��T�������tn�i²E�� #�k��т�8���kV�y|����z`��A����Ê,����Øl�I�Qݺ|�����7{k@�|Ǚ@S]�p�6��Mu	1E�MQx������(�o��m�o�R�Qw�(�p�2���Eic�7��������nY�G+��:[�+���'������_��$��;���<gb�2��-���Ŝ��+����'�M�ܑ�����LӀJ�phxc�Mpj������g��<X�>���W�Y��`G��`����>�`b�B53N5�K�36��]� �S��Z��C�z�鴴&����)g�]�J��k9�"�.R�>�t�:��R^�TT�����&$�Ʌ����^�6<��^/���N
�^�Wl1{(��0�N2G$5$���'�{�?.�g¯oCU˭��/#��r���	 jMZ���S�9 ֗[O KD[�?�d��M�kk+���a�j���=L���tU6g2��=���ziܲ$"�����$��ȓ��3�pȂ6���|��Ê��I��xM��G���E��g�[� »�Pz���>�6à�o~sԉ�������}�����
r��:������}�t5N]!�m�~�v��He�	 b��5�B=v������%�;
كw�ւ���^��'����et�_��pD��]�9&������S���Y��=��r�I�5���T�:f
�!�3�e�|��.�.5���<_�+<�{,�fN�/^f�P�������Y*���Um��tvQv$��Zpx,%�9���QG+L�*Pw�a��
�p��Њ���kttHim�(8e�I"�ˏ�H�zHU?Q@[�n�����j��5�?~W�#y�$}���z&����v��9iC³�>��V�9�0^]b�����U��p���{�_��Q�͘p��N�h�3�eECu�g��r�I�q�|}5�L�%o�j�s����"�#��H�?��2�6,�ƨ�)S��ֆ�Z�w����5�@4{���]s�a���Ɛ>�?��]�D�Sh�� �T��v��u4��ϵm����r-n�ɝ{	�_�:��5&0�I�\�{:��=>�)�9�1��Is�n!�4�W9^͏.����$�PA��?C=������WF.|�:� 龢ڊ\��UG���j$Ny�V�T�NPğ9���&\#f�vYɟʁ�^I �U����9_� ���.֑"&J7�51��\��P�}�
��,S��a�P_R^"]�x`T��k� r�+��X0���W\�"&��*�fY��X+�DC���)K+�4OX\���lk�O$��t'�g��
؋���~K.�P�1閤}�D"�f6�D�,��UHſ_%x��*#X���W��U�$��s>���P��)����D\�Z��
D��ͪEm|��g�~|�K{5��߄�a�e��@�[#<(XrsBK�K�-3A�G�Γ��p���F���Ǹ(���Cgܭ�/ڎ�R<E��:���L��r��r��xHA��xZp��Y��Y��zB
MX{�̛$6.0���Kqa��6Q`߳��D� �<�E��5_��N$���v�E6"U��.�_M����;6��5&{k���1z��i���|��D|�ĪQWK�?e�;`��6���]�z�U�U�ZY��~��u6�@��� ��ʙJ
^b⭩C���;��>��H^�
ԍ�!O-����0F�ʝ��G:�f^}X?�!�{�\�"�j,Q�X�����C������*�H��2w��G�$r����N�<�{�]8����	���l��*fm��;� k�J8\_ ���:��T6�9���씞��~���������,�|���Y��&�ne�s$S�I�d*�I%��$�1�-?!��LO��V^5_4�JgBo���@+��h��}��\�5|\:�8#���D\����@������z,��܅(KP�;�Q�fY˻1Z�5H@�� �lz�뫘�{}�V��0퉐��/+'S<+�Qʣ����LOuf8�`;�{.T�;�"��Z�<H��fZ�rYn�ۻѕ�4+��pa%�=�*A�3�ɲ��O�,�3Lːq�m4�z9"s�J��@�g���h#w]QR8Ejk��~IUu>��nb���
���3�`c�\ހl���)=�&U�����\t>�}Xp�M��tin�&X���W4|�i$.)@ }R5�ϕ���g6v�]/b� hbe0����C������i���
;�G48�V>P9 `e���jK�N���}�W#�C\[u�搢)�3l�mS~�9�m�oR�����&'�4l�h��#�e=���B-/&��_@����f%Q�@���胆��˴A^��.q�G��:|M֛���9����OyT���h9���ܿ�#k1�ݑ{�J����'����a�{��
L�܅����_Tu�O��*j�S��&���ySB��j8����ޡ/%(����
 g����YkV���%���yx����!�m| ��t��z
��-�,G����`�ח#S�)$�pp��J��nXA��Ǌ+m�M�����Ί��SQ��68�7Sϣ���Ya5J�
�{K�BX�V������ΣOo�ȹ�z�C>�%�&�|=����(�f�Z�E c��}@�0eKzx���x�U#c?��_E�
��4L�e~�1��>F���2>��`VM^i�MH��L�ĩ�|�<�����6N��յ�J�����t��=���V�p�P���mS=(7OڴR�m�!@E���d]�$��B�1$�"i�~WS�N��v�I²Jk]�o9�T�)��*Q$�'�娛Op��u���Ǹ{X�a�JVĂ>v�A�i7��5'K�*9RFE�wv����;��6c��=#3W�B��M�o.+k�G����I��^a��vK1�*d�ӯp��uy���	��4xM�w�_/�>+�H��,9�0��P'�=V�|ݏiJ�]w�����hچIŚ/k�ы���ܽ\��)��	t$�����W<Ȣ:���~ىI�,q�<����r�������үs]wy&�=�^��\�y�:���!ٙ ~AԠ2smR6���|J	0 E^���w�oY�\��H0cG����K�f�t���+�ro���dq �-���æ��#�x]��oљEyV���l[�w�=�y��	��:/�����!;|�� ��f��6rf"�#��wS�2���� �Hݤ� Kɗ
4$��b�2��"ܬi�5���ȗPb��%Q����#��k�J��B�-�e_�b�^Y�ɩt���������T�f��Gy����F�����y������69��d�����<��B��2*V���!"�*_C��,���S<���p<b׍����wA�)��j��X���U���b޽��,�τS��Z�Y��Z�>�0P�f3�E����,��@�Q����p���ǆj��G���7���Rf�כl	�� ��x�7��oɩȝ�x@�1Uؽy�[횄 8�I)�\9$�4�� �h'�3�r\锆�w풥9bq�-s�Z?����]f;�����Om��1��Cf%E�1"8����
3n66�R�����@3Rͻ�W���p��e�ox����eq
���|���z*�z�4�?�O���t6`/Eڬ#%ӱ�P���so^D~���&���&V�O�w��0팟v$�����I�AI��띔�YmT�bD��Ǘ֛��l�Rg��QǦ�/x��ZhZ��z���4X�]���k"��,%���a��%n��^Ig��WGk�+��ღnU��;_��#?�_6/Y�O���y��2K�7F���۶�;������90���1#/�?��\���a�{���2u�}���@�zgax�]wڶP(����'�.:�F۩]]%�2�V�8�r����dZ�l���@]�+��-������)�<Q�quybNE�<|,n�R{���	,�r#���b�tc|�~S�p����P�N%�>A@�rF��.K�l���WReI(U<��C�ǲ��,���2
�K��G�
����F����
��;'o���<��4�D�K���p��hI[r*�ˊ��m�����ކR^�Q�P���6(dd�!���3���!@3MIQ�R�4��Fc.M�;�5G���^���孿�p.	���L�ԇ>dX6�`왙�i�5��)���`!%v�>�C+t�3�oG�����G@늀-lmG��z��-�$����v9����p�Y{��s��+�q򥁼3�d��Z�\��.�)7���'n
��'S(5kZ3�>����i�֕�ʹ��$�x4,��.��곾z�du}��A��֟��sJJ;Oѻ��~H��)�1_,q��Ɉo]~����v���3��1c+X��梱�����q��^b��P�B�c�����4|��OM�f��L�a	Ǔ�2�)�{fEO+��h���X*HA"]�Ü:Ά�W��V3ַ�s�FG����3վe���$�*�����cm�uу�\�ztv%��a�d��g[y��^� ��풇o�Y�z8E��ȟ��g����to7צ!�n��=��VY��i�6���qd��(���b���;� �f� d�j�&��l��ԣd� 
��}G$p�+�$��t��n�d�t���v#3�	f W����0S6Н�Q���
�}U�_�sc����P�G=�D��n@���7!x�SQ#4�W
�ی�o�T��LB��|T�1���FXbz��� �@��Z���VrYJ���3�_+U�\������v�ֵ՝�T�����H?�UK0�p8�����SB)�,��U��Վ��sxהĳ��K5o��L��@�eD�⠭�]��=GZ��#A\B��+��B�Ћ��"���~@^Q`��
n�P&:I����#�^���Y�Fl���&�;�г�W����t�?�� ȶ��ϱ�돱Ե>�m������������º�z��.VHԌ��׿�_6=�C#�F�ۦx�(h K]��SN�ND�xۍ&U���7��E�$���`#�LlI����zt�I�(��g RU�>�7f����D |&Ve�(�<�;\�e{���A�Ж��]�[8�")�� �cM���#��h������셿��#.ir2¬������ϒ���r�U�g��y��V�a�.�������&�*g���2F�
�T�d5u����/��4O�C�����C�|�=[
r�+w��w.��>�v�T�� ���
��� !2.�e9�@��Rn����xͲu��˄��1I���
�Z"�OP��|țlZNm��.��r W$���kR��>��ǀĄHG��E\&��E����y���Eu��+Fk��9{��6��1����1%$�F5�s#n-�A�\���kݤ�� �M_9��Ijeˡ^╲��\a`�j�f;������d:6Y/g:��l�>i] �4��F2�3��V�6�7�]� ��朷ƭ� 0x���?s�'o��L u�OC�d�������i���ئ��s�Z|�O�����>eXUV0X���������������ة���Tg6�*U���8�:��o4�.S���eH���|~�����-r��B�:>���!�%`�i5�����~F���6��V���C9�`[�����M@�	E��F,pf%��Z=O��iB*����{�a���Q�k#BQ7r�cr-p�MX�Ý�^�!A�T2�1#7[z&��XL��u]���'B���+J��@=(�u�����!- ��.N�V��<0wʟs��S�&-��t�N����"�g}S�A�WES�t's �^�o�R\�*<�|z��K��Liܟ�>%b��q�$��}��sv��>}a��w�z��Z|(���C�S�p��P��T�8k�
����^#lv�/��U�A-QF��{�3�Cܴ�٪'%[U��RC��|���X �hT��������[f2���?G�i}%��-��ǰ|g�0'��MU��ű
7,����k4]�z���	�H�/#�ZܷZ$��q��R ��i� ��"ɄCJ)�*�ʧ-�h�
�.��_��%��K��Z���0�F�l� JF�
	1���Ý�W\��g'Ss��҃|�(~��5���v�����A*t3l���e}�X�:f�������������`���O,�"��{��0��ӝ�,�a+#�˼*�%Qf:�аv�|j���@�Y�#�f\�[�W���A�y��ct������ŪReD�r|����):��Q�;��/�^#8�3���
U[*<j��UaH�h? =���V��e����н��c�f���k����F���N�S��z���"�K3i�ZI�F�A��x=�<7?}�y��2�m�{:�S*��� ��Ae%��f_���-�۴'h�;�6�,Vw����J�	Կ�Ŧ&-�a��_��`��Pt@���G��C���j�fW�%i��8#��K]?��H���?�`]�Q�r�^��x�봶}�����ռ�g̳O��t>3�����p��$�E��W�l�,���(x��. ��.&��1%X�Ђ���]�<O������T����ù�����d���@���]�Caͭ�C��m����D��9�KΧ����C�거>�
��l]��f��t:����%Ƥn��W=��P����d.��B�h�@�����;wy�9G��\Xh��+ߜ�ӂ���T�s����;,��J&up,�䎊>i�����Hme����!X&)����l��3�+�Pw��l�f*�@���*��|N�68^x��"�� !8�������PK���;Xˡ�ά�"��*U��<�@���=Z��Y��??Ό(��f��v�/k��bW�	R`�� ��}}K�}��{�w}?���tlh)lS�(�x����9>�n�h�!��Nد"u�R�|��� �w��4ſ�� �yN%�&�t�M����$ ɽ[y�i4�*�P~����~'j��܃1������F1Ʌ9���Z�5�PÒ�J��k�V=�E#s�TDl�6Y�K��f�im��� X̗*��`R�+�Ό� ��r�DHn�~�A���р>B��c�j��'<�0�{_�������k�H;m�(7L"��b�d1��R(NI~m�za(�1П#��[�*[��᣶>���brh�:���^�C}$�����aHJG=�d׳6��<*���}�N3l�݊��px:��� h���{�bwA��g�vO."z	��I�-L�������P��U�8�I�5�����7��.�#֋��MB���3� �n�6�W�㲘����^���>#R��o9�V�e>���ka�}��a~�i�|�9M#H:�^�7�a���J����g+р߇��F4�q���Ŭ�m���Cu��M���d	���(��_-Q�@��ϗr�
 Z
��q	�)N<�������N�Vq������N$���V��Ѣ��,�=Ȃz�?L�����Y��� �� K�=s�x-L%��8ez��?_��AI�1c2�����Q��l�