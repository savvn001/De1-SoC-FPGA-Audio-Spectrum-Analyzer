��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl�-ҕ�J��6p��p�SP���+b(*��ʴ/~�vJ�v�)��ʑxv"���(D��f��@ u��D/c��|%j�.�:��@̟�d�%�I���/�
*_0���i��nt�$����
	9~�Q��_�A��O	���^3��1��?�[�A��:���j���j/�X��7�Myik����d���Kf=D�/p���)��0�C�/-�qb�����i�	#J�p��\8}�U���]؅ª_���n���H�o~��3ӢK��	�uB��{�䁀��Ɛ�m�w�_�Q+�GE"�xJ�8���Ä����U�"?Mk��zs�x����N�``����ޚb�#���?°K��Գ>	��FJ2�w�Q�{�ڴbT����s
C1|�{<�*�-g����9�Y��o+xqyB' �j�a,��=��W�p�)�	;�քg��B>��l��'�`ɀ��4&T��^3��HO����k�n�?���?�VLh�"Ξ̻)s�ѱԓ�h��/A"p��)ɮ$1��wd������h�^���)Zag��p{~G���oV�)��0�"�����7�=���Z���)��ҝ�Vu��.�W�u��/�+֚H�Â4	J�ag[ҵ$M����$�U���s���8~���̪���Ǜr7s�"��/��S�=!.~%�sg|�x�K�Xg��j�����iKfk����ᖲuc&K/*3��ܨ�s����O6�9�QF�	�67���sYz���+�����m0�U��h�Pv�c�,��UYmT�ٸ�"�=��iX4Ȳ�OfUf�FrJ�j����^�\}`�Y�t>���@�gc��.�8:��P̫��_	$9�08!���X�C
6�:H���r��O��o���Ȧ$��E]V@�<��
S��|�2.3%�F�� �Mz�t�Q'��L�f�P�QWN^��)�Y�'�|z �����ţ�!_��*�� 7��ف�����Q/�8Y��L�CUjK���YCGicV�M�I+�o���|Cf�H��*��/�5W݋��b���B���g�]&:��G�_���_ڈNV��k���ė�MP�!L�$f35I�%�N]J?�)mk(�q2��C���' ��(jl�98b`:-�4a@w���ZD�����i�rs�0���:l8xt�gn��T ��eA���3��v�"���n��]s�蒚��s�w���GY�4xú����}�|����~�W���Z����S'>=�^r�{���X{!�����4&�)U�[���w���5�T8�%J���hQ���${�vUԟ���H��e��ưi�s�p���AH���?���3�����
����TzQ���j��?>�O�嚻�LjG.��� )���ѷ��{�i��ޗ�D��i��{����W)m����)��=�M�v~��_�����nb,�{̙h���~�?��_T�$������X	�*' {�9�ە=��i
V&�R�[�&K�v8q�s��S��0g��ĕO,I��=�w�a�]�����TY�k�x(�f(�6���RMKue���7R�?:[���GT;���~M+���t�Tm��Э��[�i	jk�C޾�I�Ϡ�#����D��^���jZ���e�N��4u��p�{�0%k�@)	��"�#"W0���%*kr�=hw�փ�M?8]0���iOɁ��O��ƙ4�-�V.:D�$@����S\�� �����΅�w��"��k�Jd$oʎv]�
Q�֨߼Oə��K�s��������hGwOŢ������ֆ�*�Wӗ,d� �]�*�U�2D��e�B��������ׂ�6����M�>0̥������s��Q��ܵ��� �*�.���F��2�c�M[}����Qnl#����S���c�+*x�FÏ7����D	���&|�B���HG�����R*������H�\�v�aZ��^9]�*h�X	NT�`���u���)tv���u/�����ˑ���2ф;�(y��H��m��n6?N@��b?�I`:���wZ��!&�����I`�ٻ��Q@u�5�V����O=:��SP��ə7����I�"��WR���NH�?�u�ɜ���h�l�ZE���@�!�RGp�5��'��qn#2�5:!u�(S1R��c@y+(3C�4�*�F�916�9/v�������`�p@�o:��2V�'�Oe�Q��ٰ�$�#��Mڱ��;JG~�k|��p��.�H;���V�n��y���0�q�48�ͣzV�5�j���yl�yC���ҀϑY���ӓ�GjǱӱV��R����|�p�%F��#((�G�{;rO����Yq���s�W�M��k��^�������9�
���~�_2*}3".�rς�Qc�{}@���=Y��Ld�逬�����1��|�_���N#���]�g��q%V��<�>m<�M�J�9G�,V�-�\Y�j�9����귈p�/����_�\Eu�n���:e�n!��,�Y�m�[��/ը#�I�"-g��b��5Eww�DPbq��Ⱦ9�ح�~i4Bm�);Xk�2�Z[N�vM�2�HP�!��Ft�6� %�w=-v�\rd��kIT��!���M+����;Q�V��ǘ���Gj�a6���!jO�ָ�Z�%�n����=�x��3_h�s���E��XI皎��zh�����n�A��8
>N�ӗI==K��+װf���Ԁ�?�y��
�<�ϔEhg
�O�D�[���9�1�޴�@���(\(�pCv��>��k��P����� �����b�e���"GB�~JܲkjEf�<c���x�H��3���UPK����`}R`C]o�5*ͭԪ�?|��3��"����o�*#^�D5l�1q��4�)���X��	gAn�k�w��0A�kP㊱B��֕j]ɤ��Xy:S2�r4�o�
� �U|jo
l�-����rE4�U� ����]?ܺ��0Z�P�v�>�F����MrQ
޾u�!q��lPa֒�[���a�|R�����W�AU4TPB��0Zp�Dt��z�ۣG%fސ�c�v-+��[���-n�h<r^cE{9��u%zP�iP�#aY�Y�^�Ag��Ů�rɳ�����Ĥ�����X/�F��*0H˭�o�s��PƼ���;��D��OAګ}Z�FMB��զ��vl�h��ً+i�%���G�9����A����Z��rc���w>Z%bI���$b�ciǭ�=b��_���ʔ��I�|���*���5~G�"
�Sj�f��3W���ղ)����D���+� b.U��ľ:��H�@z"�=���}7u`��}�""�S<�qM�\#���Q�%�Ц�ט��7
�㗄�	jWG���o�p�҅�e���2�9.:k��!��V/��	���T'�M�(lv+�gӀrc�9�:>J�%���J E<#V��`�i�NM3�!��`K@֑�"|~,i���"Zhx�nş�J,'`D��4�}�3f_�ϖ=��e��$,��Q�/�	ݪE5�Ţ��Кk�ͅQM��ۧ;î��@�8]-��3Ai�!_Go@��I�����K[�){`�J)f/ޗt@�o�.r#=���Ti-+P���������N�7@n�{Y͚?n�d��nֻ��)�N�����K*�:Ȕ��/"E�'���L��>��k�!�Ư)�Dׄ�lCA��޾��a.���#��yy��խ�7g;-S{�y��؛�{/����j�,7��@'7$����<��Z�A6��%�4���AE��#��gW�;)�~��Xl��_��� �������"�3���)RG�; �AAP�+&�it�q&}̍xlʁ�O���x�C����d�mIS@�j'�,�LC�9�ڼ�T�w!���Ҽ��F�FQ5�^��1q���%�Ԭ�~�s�8��t F����A�ә���̢=��ٜ�X�����%�4Z�)�R��a�eoRH���'��w���|�;��h��	MvC&�ҡr]~PЂJ!�ݻ��q�tt�j6ܦ�?���!)�=9/+S�9�!h;�ķ�ᥳ�{�Jd:����4��jݓ�'\����}�Q1�ד�<ƒ!��""��(�����p�@��wWZ�H�;��f�EX��῞�T��p�Q~_�D���v���4Ӭ�H�����{�s` �:C�nR�@��փ/�$�4�VB�:"$����sOZ���t]�K�$��>�jF2�#��"��zi���߱j����hb�`�O���+{a�]R���j&��A�f����XQԽ���-��g!���)x������l� %�o��U���K!��I�>�Q�����R�H���ֵ�Û2[��ok��Np�"=�a�.{��|�9�4�e`@�FZ��;��nD�v��X���E��=�tIa��0~�t�&���O
��D����a��&m`
�s!�"��,�ͺzd�-��fS��4��$z�I�fpa�w�u�"U!zԙ0+�����\{�<��t���gvG�hpI�{�r���*�x'gi#��Ss�c��F�0q����&ةa���j#Rc��a�"Qx<�K �O���Ԝ��D _SP
�F���O�7,��������4���}�=H	2���j`��ZEG����� >c���	�V����4 ����C!a!�Jr<p6ݓQ�H�5�#&f�տF@���$%�(\ؗ+MyF�����Gj@S���>�g�z�3�&�1��j���c>%� 5�H6�����|�����Nݷj�س��t�5OY�)�Q�"�eR�S¦�����Q�|�6����%5�a���T��1!V��K�* Z�s�M8���ol��
����mooD9�J˂臛���|����� J���=tW�����nH��T�I�[�@����F��)�,Q��P%�w�9�l�[��0��ҴK.�f���V=�28o�x%O�Jf��/�@G+�#
�*���",��ؘ�%�ק����H2�+?YW�e#�,��
x���Zsa��A6)�c��h��<�s �>��&�A�\M��Q�[δ�c�JZ,���;}�Ss/^�|�Ä���))e0��r��8:��X���p7�5��f�z�����qw?>췸0B�9�rWQi�!G:�b�U ���H���	� �"֚y2���1�5(���=2h�x W-��uK�O��P#z1 �$� �nl�P4���Q��*���1P���>�7Q���"�I`��sz�R똈)���#|G����_p�S00b(.��?�plUP�o�`+��L�l��N���gl&O�ºU�r q���Kn]�}埥ӈ|z�#K|��+�J��*�ӥ�TP��fZ�7�z��S���	�yϵ {�x����&$��0k_�.�l5o�7��;Eu~����6��b�su#j�kFo�H��O�L\���7��"%�J[�;�k�����a���I�Ux�F`����]4�f��㹩Jd��i��Â���:3��洮z ��m�0�?�c��h�6�xNq�#2]�e5{����R�8�U�M|�p��y*s��է8�b�t�yz��ti[�x���׹�����^
l[�2��s��ː�sH����d�4�2��p쀖!�оoo��!0���uƯ�5���9�3%�^��Q[	��[�r�Ȓ��L7��]'R���K��z�1[WX!(�3Y���i����w���}��6	���@��J�J]29�j�ƍd�)<���zt]2�K��2w�*_|�7�j����6K;�A�|uv�}�ٔ��pE7*�qu��J����=����d��{ڭ�T�\���]&�|v�<٣��U� =r'LX�(fӃ\�W��k�u��J)�>�pM����s|#@PM�2�$h33N6E1�dVZb`�,	�X|�?=�3�i�����P�~f���ɵ�S�ϊ�\���2nA=~ĲJ�3�U< �W�!�H⑙�Z(!�@�;o7�2�y5c�6h<!��O�����)�W3s���TM�1ہP�չ�����a�æ�-Hw>g����`+����y���;�?�.�����f�%5� �k!��e	��B��jǐ{;`���gYF7;q�����bi��<e	0�т!�]b�-�a\yh��	� ���\�qز>�DC���	�`.�i2�˙��>����YnK>���Z�r��e�P�29e4hD��wś�mDB���'D�����}JP~x��!��D����-�Ԋ������v���l� �j��M�zE�A��Yy�[y!�8��x_4�����R�sp��3�i^�C��sU<��� Ӈ��:r0`X3�-b�	�����#w�;[�w�(��iQQ���{��w�&�ǝ���&̳8���C��bw¤���6ADZqw�M�G�5]�$��ߌi{��}eܦ�U���F��5Ǧm�w� ��֯�o��Я�1
�Z�xs �h�/5<��z��8���irGN$^kKj߳����EQ��	qu�d��lt��艈J�C��1Vdcjꟑ7uyP���B4@Uo�&UL@��f�S�>��}�TϾ~�-�D2V�v&4\��q��jڀ1UX+�F\�R1$(]*��Z���I�<(t�����ѵ��0�{�y&k�l�����t#ƈ�9-e?2q|�h�RA�;�=�]�c5��"�{a'��џ�_IvI��7�1Bn*vO�>8Kk��hRQh����V�fH�8~Dq�
����r�w3�#�P}�L�`?-�����ź�"+�̈.���쌧�nH���}�����-��
�8��c��C������QUjl7E����^�e�W�g��'/����������>jGrL�����,h$_���4~�k���!��+�G����3&��[9{����+��%L��� ���'6��Lϣ���1�b�%�Gv�)���z�T��"t�c0��DDEA��֑ݘ4C�+O�*�1ȼ������]�=+���')?�ýY��
^p��x�*0e=N�)i�o�'~N�!�AAchMp��z�c.�����_N^$�p�o�!���=�J��6&Ȓ:�9��g{M�"�x�gz
�8�5?���S�&�U|$�FXH�� �����sZ�z{��~l�~F�;�ޏa�4H���>2LBty��ꀂ�.� �;Ϯ��n�4�\A�|Lk	�_] �����0U�>2�4B�J�<���s�9$v��M��`��sJ�C�;�f���*�탤�.�3��0%��і�S��w: �;��\Sp\�C4	8�Ζ|���#GA%��D��	fʱ�:�|�G;d�*��~Q(������r�eI���c��ž�AY��{�O%�hl�H��ľ���PI��
�*[���i�����U9��4��D�oK�����=)�6��x���|�k���ˎ�}�^@��r�g4b���u��r��M��âh[^��?�V�I���X�<��]�GG}��4���#�� Ŷ#b���%g��nԼho�2^�^\�|?�M�ë;)1A-��ʨ�,/x!�*h4LA7%�����/�J/���/S"3�e�C��y��`��
#������މx��2mNu ����&/�E�.P�!�;���!gU.Bf�Kn��Z�"�6ޅ���I9��6\�CV�[���a�S�\�3�zt���B�
��Ok����ƌw �N��|T�\쪅�X6�Z� ���sf�~�;��9�����-xG��3WR��<lԀ�z������4���< =�	����[��3�Z) �ʔ1���3e!U�P=\x֬J�OK}� ���9�5�E+�V;����<��K1�ԫ�׾j�Bd2}�	��#�x�C��6*e�p�FDq�KH�FB����
(}��x�O����l@j߰���=x�����z��[�n�`|��SN���0��Ӯ�(.����xc��Ѫ�H�jxLx�丞�����Ǯ4ޜ4����c2uZR�T@�%�z%���Ȑ�3��d!��N�6�^�S$KE�wҽo�H��+���(Ro��I�gi�QG�4�2,J���!�z,���i6_�v��kSm����f%��Dw�,uЋ�h4!FK_�/���h��⢧�a���Q%_�1�E�c�3��fWb�°6�U?�zw������7Nv���T�����V�����+�^�L��4Qwv�!�Q�jAMv~�T��vs�� =k�\�f���>��F�Ei�I)���'��-q����mkx��"���F'�1��?�'�����EI���q�Ӕ��'�
���(�&.�W�Ǜ΍9�(c8�m5�����b`L-�;�����%Q�L��Ŏ���5.�\~h9Ū�!��D^�z"Ɏ�-u�KS?e�=�&���ou��>p��g�N�Ā�K�����.���q�����S��ȷ~i�'Cʝ\[��(�U~�+2v�2�Zٻ�1�/�y*'�UX�$,�Φ�����|�0���h׵.����n�_ez��Ͻ���R�Z)`�L �2�6����#b����!���B�>i�o�|	)�tg�TS�n�����@V�b@%4���<P�L����?��]��G����/�����y}£W}��\h8��A6R�H��T�O���(�߼>��ϳb���51���R[İ�^Zq9�v��@kfw ��>��I�nvU�T�|�zN���-�s�<����`�j#�����7?��*~�#d	���I�I8;a�n��O���`��N�G�QA#op]ux��F�3 ��-�rp>(����Ҳ�/a��z˜V��M���V��̚��G"�}O���S�Jt���ѭ1��R֣pW;S��6P��~*%e�c��1-�E��<��D�f�q�'6$�Q�t���0m�|N��`�:��`� �ei��Ow	�K�_h�/E��7��]�?u����z�"~ X�^qF��x�����u(z �)+K={��p��a_��{g�҈Qe���~��`Q�/���.P���{:���1.�bs�W{,E"��P������+iv>�L��q�����5`�~XM�0�)$�g �@oK�z!�WT',�����D��9O�y�i��7)��I㷶��9�U�3�!�g�rI�b�6�ֺ��O{opG	�Jz19R��5^p��Ѵ]tƱPѬ�܍ �5�^_��d��1;G�jz�{���� k ������m�\�p��ʰ`����� ����5���,ı�k�o�!��Ip�5S@�HМ�(�Xa��D��,K�@�V��n�9Jx6�0��/�,د����rz�F��2sNSrR�vA�	�FP�4�<"��O��K�ls���O{5L�(R^��;ӟh�H�(��M͹XrBUW��l7u��E��Ţ/��I�eL`�#m@q܅��나�l�\��}��q�u�m���ZW�D��#ˢ��3��l#�>n�x�毰��l��B��~W���ȊE=K	���)�}I� ;U�?t���g߈�7K��%>m�skN'I*Z�ۼ3#F�ڂXuЧ�2��s�[𿾌�a"�ʚ����/����߿�0܁�ݪ�TCB+"�<���{?_��-�����ĤVsv0υ�+>$*���}��T�u���A�W���v�F�X��fz6 z�N9�}0 F��E�7�r��)v���p2Q�0��|�%��cx
�Ū������ˈD��2�v2����)]��u�ם`�%x�"]̈j�o�N��Q�f��h0��T��)iX�e�=�;��>��q�4R�Ï�� ?��
����ؿ�w_��|�c���ݛ:f>ִ������V��r�;ˑ��C�p7�J�����79�Wr��bU�a�mʢfX��ኑϳ�D_;�M�� Ҕ�(�J�7Ȼ�����J���ˌ�MB������0����v!�I�;7tDKM6l]K�[�0��6�]��^b����F�����3xS��/��+���
�«�N��6b��R���B�T�K!�=0s/ڌ �S�j���bp5`{�t�Ѹ pY,^�J��t��G�\q�,��r� yz�˜��>���c����&��p�l��ȏ�x7�\�c�U&)�Թma��h�� >������_�x��B2��F�������4&�����K�@Ё�����N�镹Of�������ޞ-�LB��[�0#������z�0������i�Gh^z�{��O���Ҟ8�80����Ś���;JU��d�7��`o��\8zb^?�OT���ؾ���Y���B�3sS�M�H �3�lZ�`�����1<ᄽ	�u�D�A��s�A��˸�:����U7Ѻ 6<��f]4���ߩ���OsD7��O3RR���-�}��~6<a[�_�_�< ���.��Xt4h�N�������::h�sR~vbȆ�9�N�Ŷ6�-�觉��ǴŌ�&G�_'w��I3GDad��Xq�ݨ�)�4^O��Mk�� jE�D�Z�wN^���W)����=p)���f�l�9���q%���Q�	k	��Y�e�M�&2S��M}�f���B�2�os�;&����9BK!A؈D����$*#�}�q�����2�4E��m�"!I2܍��]�����5s~@��G�0�ʽ�1�uK˼Cz��QDHb`�1���Dr�9��S�z�U���h�`�~ڻd&�La�%�]��o�(?d�k��'m^20Z�b��vGVjbgM���F1�}0 �Ѫ�Yrwr��C8:i�QL�0�������Ȍ���e�9=fȾ�@xbQe��>��|4lag��rk�zN'J��kSǈqly�k�8�l-���J�6��r�gU^��uQ�AYb�[�I��D5���OH��d>��Qh��46��.;���l`�n^&>u,�_$�I��S�S>�J-�|f�jtn�,8Ha�p�nY��cUG�mE�!ixЙX�j��7u�x_�����J~X�Ɩ�Pr��:���ܗ+/�Oק�&��H�A=r⌲��@NP��h��
�����Fa���욢N���~g4\����v�}(ˏ��	9�Ú��4Up����K����zv�*���f��ОE�~�s	]��O<zS��߭�^Y�%�]+}*}�G�~E�&����x��v�`�x�'�)@��:�ǈ�+gNf_��81���'�*��PW�N=�A<;d��̄���e��>�%�>�5�5��fX�8
r�
@nE��ER����/0��BzVN���!?�O��RX:&~����C N�t��!8AX��g�o��;w�R�c�}H�#��
������,>)v��DnD�ޮ[�4�:<w�% �~���]'܌�l�I\�`O�J�4��=*̅��� �Ћ��6�1�h�ξʚ�V"�qJX*�,��;���=H��/��Ծׇu�@3��Nyb��L$����(<�M�{q
 ,���
�#���3�ݩ]#Is��/|�U��=�G���1Iw��T�^�����6ɠsooTL��T/o������$[
ն՜V���a� X^��}��(����&���}!��5s�ﯻ��F�_N�������>��h�Q^���H�[�Ԙ�!����B���g�|8�G��ك\�����.��H�r�h�K˒ڹ�%m�a�$x�i�P�S'�8��@�ur5�	qyl�Ъ�bq������C���[P����U ��Dm�z��{�B�����;��yM�f�Ȑ Pf���n.�Xd��Q%7���'�?��dR��(`I�$��$�姌����Rk7B{ʒ��?%��f�ot�|��j�M����0���DA��-�ކ� %n��<Z9��y�Ҙ�uGQZZ�wI� ���wT�����L����;I��������	��8m�x���O��6���v9+04]24A(���4L�#u=h�T64x�c�\�.�d�S�3o>����y����:�#4� j̓���:*��J�w�;��A�����Jy��Z��f���Vi)7O�k!<��^Ɋp~��߿���9n��7y�ѡc	o9s�d\T|5���'��)�f�T^�~#��!{��fX��\�	1:��i��+.C.���<2|���~�&oq�C*���F��C�s�8��V(X�ɼ&��D���S��[�TrH�*�\��[˘�lu�WV����suU��Z�	_͟�=c0�L��d�y;4�0{�\#�b��֢���ec6�=z]��gt�0�Gk�[h���ΣM���Y��l"x�w'�s�V67���fl� 2ᯢ.���+5�Wrj��1#�@Z�m+A���@�0��'XM"C�jG�����ecZ��w|9FSǉ3o�Z*���_s��!zٹ$���7Z�oT.xNWz�������q�x1��6��GZ���JT毿��P
%%�[&��נfrR���A����>�a���h4���S���M���� �B*9H��:��ڳ��Ct��G2�%�)�7�~�1A3����QC��w�+��K���PO�F.��ձ�a���`h��kt�mA�>Q��sG�v0�K������-&%��"�b�C��v�i�˾�U���,a�.�"�A� �uꢉ��K�E�g��:{���� )�H 
�y�����OΙ�H��2�����Q�0cX����N� ��m�� ����${����D}?�82H���@�t���<7�h��X���g?��!�Z���'��(I�ηg.Gm,�D��.��w��.ZBDҳ,��U����>��C�hŗ�{?��S*?�n�F�G\��c/m!!0��ޕ<���5A�Qz�##��H�Q���=L�筌��T��P?�z��/z�!��޵����f���1c-krs{hz6����>H����ʄܮ���l��l�k�W���]����c������z�6P,~�~5_����X���fr�/�����P���R��D�t�BA�t+����v�>C��o����A�Gu�'YG�hwpv�2�r�Q��dОK�}
���s���5"z�V6E�΍�Y�qA2��v�X�'+�
�GMP����jt��6�v���iVw�4'��x��7n��K?v:���^{�!#�ڱZ��0����|�`������$��� rz �`�H�S��u�?2���f�Y������B�x��}[,�����T}��W�^����F�oZ��s���A�,ᕶ�4a�Lʡ�2�@>uQ�w�'�;�^���� p���X'
�����YoC�n�3��!�P�,��ܝ\(��[�����zN	,������[����Mi����@'�&���'��=嶾فh� ��F��f�]:��F��k�!���o�b�?yJ���,�+'c��]�<�ut�ƒ8���Kf�)C�*����Pt���W=@�y���ɘȖr贱[ͬvZ� �Jt�j�*�LT�o7�
����0������a^J���@��@����a$[S���}��%�7��t�3���Vpe��ޤ�<<Z�,�Y�rN����wpr�K�4Y]5�}Z� ���0�|эb,��/�?�ݩ�:5M�v�3���Tuc���U8j�~hK�n�ŋ�d�p�"T��9j!��\Ψ�������^ˊ�/6塱0m���.�'3�j�'@#b�(i��Ɉ�V��.��,�R&$A���5?5��ت����r�^8�XD���2*�{���Ci��OF���mD��D�E���옋f��@C1��}�٬��L"�m򛩧�!�Y$�>Y��0n�q��1T�k����]�nm�����$I�}�٠��BU7H������_Y�C3V����,{��~Cn1�E��?�j��ƺ6���:�;fg��q�^ԁ&GF�����uD���l�$�7�$ug�![x�^{��w�.b��6�^m˸!����Hk܉��2ENdF��3{�2i���.�(ht���@ f'�%��XQ\�+�{�C(D��I[�`^0�U+���>dT��;���tv�`��� ��-�4э��j�дn;Toɓ��/2I����v��*�����qZ���-�M�9$DU` ���[���s��Hbftc��m=�z���yv�~��f���C;������A�OR�K���jt.�% ���-8�
&�A�ǳq��P�nᎻB�� �rUi��'Ķ�Z�����lN���6@&�&<䞒orǴ���փK�G�����X��`�J"���Q�g��r�W=�����yP^��89h y}b%��U�DFP�b)\L��3fU�t�W��B�|�`'`2�XݺOG�X��V�� �z·h�"x�PlҚ
ES}�����5F���7h���0з^qC�_=/�hb��|O^�����.W�j�\0�	L�鎓pA�v;s<3�Ƽ���']A��4��'9ǟ~�A, ��2T���R�ܨ
Y^��=�s��=�GN�![�G��R���jxY�e����&�~��h��A�-xuo�t_���/a��-U9�d�D�Mg�5�|�����+�ԃ���/����i���/ë3�\��������w\t�!��$�
���+����Ю��oK�bL�cY��UӗYUڴ�EG@Sޭ��D�I�W�,'j�����3���+� ǰ�?1���` k	z!_�Bp�ݔZ*6����:-H�֑��Ng���R�hG�����d���m%F˘��$t	��g�v�D����'�Ҍ/��iq�0ۂG,_� ��W��&\}� {�LLԙ�=w��>#W��������>>��8�!i�"OBf�glT��֗t����񨪜�,�E]u�
�<��l�������r�p(��g ���(e��{��3�t���[5���G���=�N���FaX�%���菨m�:;��[��.���x�2�C��@�o.x�q��x���g�w��ZfTN��eb�N^`�]���2{`:�OϪ���w���X�K�nS6�Ғ��w��<C'��̷ms��R�;��!���}@��œi{h�q�G�s�N�
�X�H�v�C�jܫzW榦1S�)��tH� �l����2��f��VvL���c���cފq)�~@
�^��
�C${<��Ml�U�K`���$$/��Dx�]�7W&��ҹ=��Q�Ϡ@A�vK��&�]k��$�P���풋�����Ec�a u����gC)��3}�bj�-dW�"�)�ĸf5U�u����tB���X�_������uW�Es��oj�y�h	�p�]P�h&)$�V��]�f2�NR~ �<~�� �i�����k��#�b�t=+���>��$Pp�j=	�]$��0/�jE�G��6Μ��� �J�|i%F ��7}�����K��J���m�\Eq���,�qGH-}�tIOZ�+[`Z�h��
�H �7đ�zy���^�/���N����c���~�D��߮*0S����N�x��D5�p���O��	r��v��\M��z��[2?��^#Qm�K�n���m����Yʋ�w�m���?Q�R�x	"R��C��E�eҖ�:�P."EԄ@�tZ,+E*��#��� n&l�7��S��A�>@NM%�]���q��+3�D�{�r0�{�"�sg�4�+��������C~�F�lr8�?{B���j�Ĥbmk����d��=�� �"�W���kgsdd_��*���+��n�JLqʪoݽC���<�Fj/̹��s
d�Ӟ0<�����=:h�P�ѷ��p��Զ^�u1���h\JT?��h�m��s�d�0�ɗ<�8<�ƭ%7T��Ќ��6�o��B�]_|��oV��t�-@�ayB\�U�X�:P0�2����$�j��s��`id
1N9\vs:Uyƕd}�h�����	���������"��'�oY���.�O�0�����z�u��[)�	���!�<Yj� A¸iZ,:�(��F'؆���έ�ݚWL)�Y2�p��+6�jֿ�V���a����F�1�"~j�u���|A7�b�&ro�A����Q�]k@#��-�W��&�kd�b��[��R5����^9�~�($�����@3�7��t�i%�[Җ������/3�l��;2�R�@e4�2c��h���&{���_��3-�j���j�1}�<�2�0�Q.��I����Z�8���V_�4���gy[�=�:%_D��˰`���2��s���������+3�f�=h�j���?���(��d�t���(\��*,t�6�����o�`�X��1�Wj����Y��t�$?T僟�F�a�^�<������lʘ\��*���9��]�`��U�'n�M{���)p���V��h:f.,�El��)���P̮�Xr����6h��}����W���Fˍp�/�{Vg����6Ș��|O���+�1M<�����?/�ޗ��h�8 Gc@�F����gl����O;{Wj���9ԏ7ʷ�0V�T���H�3-��{����s¹���7��f3?��?��v�7�o����J5�H] N��Fs�5���k�%�Y]�f�t=�R)�U�O6������1��/$P����s�*������r����;���վ]W�=����-��z�)��j-�xT�lKO�ThaP H�W���`m�È`+�oÙ.����-���=�P�4��?p�����_��ś�2����IRuEw����p���1^�ے��)�� ������3�u�ÐP@(^\�"S<�u�@4~M�3o����'�Z��v?s���`���<�(�&��s\^���57*,��(��7��v�(��?X�_F0�`�-���M|�Z�fM��2�j��MW�m�J��Zr�p 	��Dֈ�GK��m^�i	mAv�,|U[�+G�%f���A�F�۵�	�������(zQ�C�ЖSޒ�c�dЎ����?��5���|�i4:?6mzo�`���x�E���n�r�.a�#_\�͌:�O�q���wk em�?�]��9���kR� yJi���2��F[������{`�5],�[6 '<��LQ$��6��jF)$]RM��M4@Pa����]��:�j�*B�~�Uf˝�l��B��Zc��BNx�8!2>��d��q.jڶT%��d�^Խ�Y����d�
��
��\;q���؛�I��<��u%~�!X���~v@�r1F��V:�^���@;D���ڀz3��~O����u6�Uo���62sd&�l�,�<T3 ��+언���է�����S�3�.��a�e�%�,'�F�I���\@<�u*�^�Dؼ1��Idsѝ\�;Vf����A$��8��KC���G�:���V��o8~@��	 �ގ���R��a[6�?�'5��:@����$ڞ�;�ӐI)����N���w�(%�����	����,ZS��-EպCG���mi �ٖ2H��C%Z%_rE2�!��[m�y(�������D5���#��v7���Ja�V��5x'>������D��u<q�{���aZ�mx^n�(���z���[�ٙ3q8�y��h�*�g�t�Hne���yu�����`y����	�~�����Y7X�h��9M$���2��kbx/&��]��ē�"����S[r�H�R��R#z�2½��Bu��f��\��'<�)#�c�e�7{����$lO�({�(g�=�=�/����?Z:8`�h��̷ �{�8�4?��l��+����Mi��}r8[CHj�~����"�����6:�{C��Ԟɨ��6-���}@�t���������o�A�q�ܟ$�o���]�Sq� F�����,1`E��Ȥ��*�Q���[V�型��9�É�aj d$�8V�b�����Ѩ!c�������x�f��M�J�o������ {X��'�d_�E�������__��u�8ٳg$�\�[�Q$�i�#���b���?�u��0Fݲa���F��K ao#�`�++}�8���\u�!Ks%��W/��q�'�gv6 Y�Zc¢����nv2��L���f�����P��{�X�(;^�B�z�*ˀFY0��$�9�j��"��&���O(�����hCT<Jedz�}����Ax=ϩ)�N|�٥I����o����7�A�N ���45�����w�$����{���O
�~:~&T�P��J���V^O�����6�w��D;��Z����5<;e�i]٫|@5���i{�F^?�_k����Q���yo]a(s�Cf���8_:	��Ӱ_F�{��C�*c�U��hk�^U���6�%��}N-.��]K�U@�睗��Y��"�lBʓ >"���vr���.����]��k{[SJB���.L�=~�C�ͯ6U��j��!��%���cO�f���I���Û��