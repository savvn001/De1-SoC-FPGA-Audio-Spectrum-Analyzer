-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BG4RMR+LrAuUd8zd2eVJ0ITjDG9Dm2eLN3K29pR58E6HoGYuvQx1Lb07ryIu2B2PaAREzcvyLfIR
Zyv8iyJrn+6zznmXKvXRp85I6x5z1uWARKuokwpbtr4KvdUIeOXstjGNiGYe1VJq/Y+rPOMsPoyj
wPC5SXOKuyDff+vUVeR+J+Bu+/DSn/fVxoNDkLSDk5FfF3S3JwARMOfFaAG4zoQ+8ZMN4rOJTMNw
1xvj/TVQjF5XcWQl/0uwVHU0ZFWPyJgr7pjo7kM2F3u+WoJJHzr/Ca8HpC/0/3Rv3/gEUQORia3Y
+jhOtkBzY6U6uMkQd0CfiI90CsaiD4c6I2eQvA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
/hvD7YD2pN5lhaNuNrWcCBuGIVi0nluJHF2Lw/gijIzX5uxkcd6U0qOMsbH6C9LoFlDxw5166pdq
VkxDszjHWHCv4CTg7NVITZnVXTvVn0/DUywL8aaG4c5PacZVsHEvbAkk5nECUq4y6bz1JNUcoNpm
+Ys3i1fPFDy/wVeSkujkIPx8J1LkkMh3m/bNkEt7xl1vEQ/B0RPQjt1RERKsC/lcr2SxsuOaKReU
E28Gf4S6KnhcOl837PnYYxGwTXIrtqkqrzydhdEKKlYpnEUQ5eiQppiZy7gm9o8fM+7D7UjDoNYa
XcU7HxniqY8B14SF9onzZkMwK+zrpEtbirWU0TOzByESbfRLP+CH81jiiIU8cUpdz1wTQkyMdZEI
Du86uddm1x+9DRE57jfcYSrohLw24Li5NkVsZf/e77K3AAFcEq/VSCZqZn6P3hD30WBKdlo69YaJ
7gZeIZUAU/AZvxug5w/+jGkbG3Xh/YYMDYwtbMRRiRUs2eftDggTduA97ogCN1IiSYdGN+JxInkf
2K5CtFkG9O98paVNL1vsUzKu5/kVWpuRhNjxYdJaGIiR0lwCLLpxv+gT82006UwLUi7XTYZAICpS
mA9kx4zc6zADccNi5rv0oEVEj6D8EFdjGFFnbC2T1PuXMikWWAUHcSJqweL0pxArjR+R/fPsEihf
qC7eUhXMKkavsR41iJIAkzRDm5iekFcrTf36bxv1v5docAbbzKUyRsZtlHahxSgIAzPTNgO6PSGI
04HNDGNZBF6/Glih1ZaVjbWly6SOY2FCXfeAvl9X1q3TQdAPJG2I3N7sP5XD/JJ6r3Q+MmGz8j3C
h6tloy+WjgJZ/dlneCV3AOTojVS6GSEcu8x1DCzSEvzLLxri01GHo3hy8s9zodzbWMQggNMvfHpG
xNn0QxETAfefLaNaxJclKjV0bfdcnN720xJjz3RpBPA9PFuWYaqQ+ULEPt/bci5BTIXm5wHHbdkd
hU9QweBR0dwkPGQQ/dY487GKOxIgBxKLecg1K7SdJU3heo8nS/T7/yDGYcQ3rYEDWvVlcVZrRkcv
jKEGzj1uH8XyLl506ZnRo+nmHxzNYUcNzjc2Lq8RbOH60mEUsQm1Yz4FgCUjQP9JA8QDZZCPnDfF
zZlFABH4KFYx+WgN6RMuE8xuI6tAtB8aMLBbeegIN6/1w7dvlVJK43L2Wh2lGrP/0fQUt3BOE7VV
IXDQg+sJMUjw1qjmlRtYjhEvWV3zEVqaMTYoyMjaP3gWbeSSkaHKmAMowEOGHMIUUKmOa3J62h/A
dm5rWMs21Ly8xmzbWeFJB3YIujA8XDT0hChNBgWwkEvPZTWxMrPwCROPIr5tVUxs2kP9gLEM/Njj
KdZAzYWzmT9J4VfFcBafvp+LGpZmrV/aQ3qDXQyyRLBCvtZPT+kfURUiczCHxXaVkoz4xMOeOt5x
MeECgK7p5cpg3veSOS0mcgI4r4h1vpPsJLCWK7Vu7/1kY9Gg75OBz4HlUPyqD/jNN5kQvapJJia5
0vp4pdtHwsy6dpNQO/6nwfzYysWkW6RawNsXi7YkiJUPzo2ru60OBCB4bvpQ7xehJBq2i/AP+T4t
Xwv4NyH/3R6P6CONIwGocqzs+tKlVIkYi8RKLukEQ3BdCF4GrleBSbq70n6id3Fy9Ll/KIMecMZg
a0nDhbg4XynO/jeMe2goA5Es5zlH7kliGrSbNRG6THoQGUogRxuZj9L9/IdWDto6RBg/HhdRDhBt
n/bLPgbYY2SFOoxWUSoONZa9MnGGDMmJOFzOyzbqZskz+pWyP3vIgEd3D1OLLVXirxYmWVnk3I+/
5BUaxVSB62rG7ptVSXPrsNkDWnf2V77ztIl7JKhRme1E9DqXsNo7asq3gqFqO6dycW/4Qh8fqZkl
sKH5BeeA4L4aByU5teLl4zPbHtuX8+Y1UMV4c2qeKVh9rZmkE3mZxnM7JKEwBEjNLiGPF00cuz6+
nzR92B7hlVAegwSaCDT+3oWPfxVLCI1mURMsjWB2YuI8dXUeKHA0cvkWpxh1dvTFzEt+yZkhOhj2
6zwFGX3aspKkrniwnrcLOwCrE/Ox9EG+yDUCVyZr6P5sZQ3h24gYnhuTLY6eErF+hUERbBDhffUk
7nmEfQfgcPswJA7awl8GU1zxutIl/mjw75WGmbs9mNp8927kKd5+7NCcY0ZvoVFFRyRisFpJE+DZ
/ttGBMJoCRooDWES4kkG/gJSEa/Z87oMAlJHbsogdDyi5VNM5Kup0E9QZ10zNXV6nXeBPy/REaZz
rIe7tp8UvFlAGjp66TdUavuEX41P0ebZbloRSqrNgrNvxpCMOvr9GMNDGNUruXv+q+FtIJSyFMP2
RQpELAVoa4qSodtO4bvd69F3q6sZgrRQ5+9tWsB0XKar8DcVLMRQJPhaCUwStOEaOZGuzkBtYlK2
vUMK3TvzLbXIdpoVbqaqflqRpUK3qOlFaSFkQ6PPDDuu94Kd2ubSpy4MnBK/Nf/uh+0Qm/7F4is9
Hu/NjYgQglHBs5fpx6NAhh/QAabAQFTrVTnD3kBeZakcHB0vCHbrXyNBJIQwZSrpl01emkzewvEm
1HAZAuUI60HueX2quOuSLxezoA0qnknPZXQSu8DrX3uAZCgrLTKbeDJqj3so+sco4VhrZ8ypJhBI
emhNDuCblC6Gq6bfKRAGEqsq4XQXy10QUkWW3o88ONY+VnI2oR0OJY39aOMf9WBMAU8qlSEgt3nu
CbeMyOLIR8c7nxYVUzfy+Lhk174vlusQoLMJaAgcpizZmI29541MwADGKgcMIzZh5yWWLlCjnKRF
qHgEXNyrvQ2MBlFFp/YOe6vnjajbuH/Jv54c8hA6bgm/wquBqwYje8T6MiRaryERX4NsBKDgFGGs
/bnorV+jw9552AMl24YGdNZfobPkTTIu1gro19oHmJLOAgJjSIrHG7Is78UGGoyqY0l/eIt9gCES
4Jz0iefYSCoMeX4z0Env/9iPU2E1Qo0YAWM2je1ZCUWVG8nekIZimIPcYiw0RmyUFgI49ciuKPVy
4hRMzXDZFnYBm/699HBp7i2CAnbgvyvqQaTotoT6jA7bni82j063Vgn8jmX8umV/rsgfPgq7bt+s
yzcuwVg5kSnVnxFH6dGZiX8pmqXZyjYxmOC6uRIx5l7mpTCzG19ZRN3EIjUQNE7ZMOrEwggzq9UT
ZEGGzBEnsCXQnvyfGE+B5stnnkvj5GNGNSrxg6I53Oo8OE/+JldrChXk3Omcnfe05+Uua3CutSj/
KpsPR8FGUzHJLKPXaxdePBScCrKbYlCvSxrlX4cfgR0Qr+KI+ebYhX9qXmtmf445w6KqpZ/F6dLA
4Oi6Sre224+nzY67ItkgsbX6qEyREfAnf748xoBwpdLEBDxpPNAJdGjLLA8rPIKsJD1Pp3p3ybFo
zj0N+TVE6F4B7KEvva9eZ/xppWH+59b+D37lRTlGYG4IUsb1KgKYyd4r9AgsRfAaZYbFw7ajmmiC
ZHVFAXrHlfFrehlSreLET+Z+ozzijQnG07cjNSdxr0sODFFm98siIcUbQ1UeU5+y/PtfCgxmle3j
a/n9xayCjH04TNwGzBPcXucC1GTaG3rx+yLZt+Zin9UMA1qVyINqMudrZmVoK1cSsyeYHJPCEmZg
d7sCJVlqNFjRpS8gq4HvYBaxBOVG797gEQzv6BAd3lERyYaVK6lSZfV7dh/+IMZdMvHO2RiOE9A4
jIHd+u/u8AwqaEo+9mEDSIRqImSYfESwsLwjwY/pdrgZ5PX9ELKzNBF+FaIz0JWA+53VT2zUFq8G
3AYJvIRXlEBLjSVaEPEiPr1eW5YQDRCSWzxmzkQ45GwyxekIyEg9BwUH/PR+6kH0L4NtDXi6kTtl
U/Q42/NuwTgPtstKVsZF9FMrCt3Ub101r3MQHZhjYrPy0AzNEKU7ibGGrDOe/5N4yYn3XAp+3cYY
eeOre7eRjtRhRy4hKdhXI6ae8Fxo9GtPjyuJjYrZVpeUi729h6I2TEEgynUTsLIsZu+K6JkytVNn
CQJ05TVXnpVMLPrMOvP/XI1ym/asdLyQEdFHB655cX62n+OWVVyuCES2iohhneaGHEj+yKobYUWK
eKoUqF1g0uAtCFL7Gk7RyQ49wyZVo0oUnHDBMoBCKamBX6AjValbbDIt2QiptdoQbItbOXORwKgV
tiwjFp9Pu7E3LC3sQSbxaRGyrtG4fSB8tySAKxyeQVw3iG0kh1Zwq161WJd9Bz213C7uuSi992Vp
dtoXUMpsCL0N6xwLXqjfS4+Q7RoAR1Lee0z6aNTCwWuaOt+ZlfSuJN+DSShx5KR7xqpNxOQUb07y
uR6EfC+zoAJK8YoLUfg/XbQOD+nNlQ0HP9RmNm2CUyOW0AoXpzi0slojf4KYkH6osF70MQhLu+4Y
ukCr9q7OC0AZ8BzR82ELFNBdR7vr4YLXl0e7jfU5kYJTTsZHysj2BFsJ28Lyw7hkt5wF3Vd7gyWk
Zd/xUq8JRaE3SrNa38SjNpyZiLZiMl3oAtbFEXVDj665W5/9G8kd4umJmweTFSgD8GgT4tb/s9Vm
HL68zggTqNlbB+7O4Gtn4aZFZsZExwOl9KV7LZPtChSoLiADlImnfAplnNTSbRdzZFl0NlrgVeMK
uCHXTYjJ/k+thoN8RBJjZBieSFN8/rpvYQ9eLFwBvjzeZ7nm3t/dpiFyGmWS8MuKQaRXvvdjQv6T
9K9MBvkGJ0Vr/8/VbBbgluR99XDPrFoG7f2H4ruAcXBPQVN4Be/720F+FoG7Utb1NHiUXUhJwHOS
+KoU49yaNxGV14uzyd8CsfeW5fGmVpwTuH+0Btcln7vaaYI+xvzLbAsD3ACM6jlcfdg2VH9lQjVQ
bRUwXOGokSB1SSYOXvOor4GbWPqztnXRpzSlMSfM74o0DYNNpaCTezlYBPpZzcnj0Ze1vMpkfony
VhMFhZhOlER9Tmwo/4U8A8lS0MMSu/2quZwFH8WnEccAmKDWASxMKXWpSnU0TkK1TgUHRuVu0n1A
Cz54senDkDeGR+CfhajO8OAADmSALP7MimaRaTHoOf09p460mgFp/Fmb5hUewg/6wuT/Lq42eJ69
RhJnL6LYWz5HnQ4Dtzu7SBJ4l0o58OZUD86sJcFmXw/O+GYELUOVMdPFEJzBLr1+xaxvwJCB+Zd5
p77THO9MSTQMMF9NdnYZy4D8pJB+JlUnE2QFUIf0nU1HJXIBCxwrWq6w3bKr1YROCEGXdyLCSDGc
bzbCvgutCDcl0+oCzNOzsacUdGZCKdLgsV/ZMUH2irY4yL8n9KfA4dJ4HMhhNu/37hmKExit41Kb
pl4Dg1diIPj6cnKjaHqg9+esyYTpehzVHua0tJ+AyO/tb5DwVhjnxuxNfoaczZcKaacX20ytB+vP
1MSAgcTJ9nSYD5zVHmFBjW4WNEKAFLfxSuj/z5cBaZbbITgDHQGn1QuhnMiLz5CCOEbQNguoJKpr
Um3YmI4FEiRRdOBsZlr7v6WdiDj70OYkT7AgOI9K48C6Jd4MwwfBcKzbSYORs6HxLkXIZgH2Ngq5
2lK2GpE9/DAWT1w+uKW9L8i44byBDPr5S/xVws6+Um0SWON/H3sXylHrzmgn/DkMapf2YzkuEW0k
vEfMcW478XeEGy708fS0u1d2/WzbaIQtwpjFO92/f91u6+dVhrLPWD1UqdethCPghE6TKJKHsuTe
1UwwFFr4c8d5cV9xclbYFrsX5b/l2ZiWFSeUEjWtMqzz1nOfn+7hr1Yq2UlTuR1k1dvJOROvF8lB
HrJ0Xrn3HNTY01Vz9mWC6pzmjq39/9+gEQYjETUhxnTjyoOn4HL4pgsrQzor4Rux+R3s5MWMlm23
JJj71Mu8i5x7/PiayJTrip3RdxFa3qYQHD9undZ9pqqSuxiqW3JrCiqsqir8YL2LFZ9kgkzaxWdL
MgfpgUcB8VCEbCjIMFDLV+1YwUspUuAflh8JGcLisFW5XIGiH71Hus2nqMD65o/j3a9SBEE+8yR/
S3qmd+QomeNT8FSQXgUWtm+1tVnAMPV0H4ZUoz2rnQho+yHqQCWhlYWER9sQIcHkqKKs67bv+/c3
buD3/srokGzf98xRWzifrmisn6wCkUFrgBvpHm9FQxTtvDysr/QF1cO5wXNncImSFNQb4yVjKTpN
Em+NE9qUnVXuFsuIvLKMCTHdGK8Dih9O5Ih0oLxa+Zesw4F2UxDsVLl0t1RSaZFRBCfKlnfxE+V0
RALIvdyu6TlnGOpUgXT+9rs/c9x9fHAevQz9lP10LM6EOTrcnqml8nuSKgei7j261O8kDYK97MtQ
4iDnqm4cLdt/WwE1mTuJ+397mH1/Lwcgm4xR/Wj0Z6G3earG8wAScokWISNSGpJcySDEAJk8NLNx
Wk5NaFT3xhVSUjF77u0M8039gjt8Yw7iLM2ii8jQfDDDnFwtcVDlHMHg1zCKvH5u/Gb9Sc9xm/wY
4Pj0c3pP3HT0ICQyePaGN8sKJsIKrm/jusYGCI/ND3Y368PaZf/WPUGzh1WkKw+vCSQQUSQaCjvY
Dx/ZrdYKkTnD8toAh0ENF4sYXR9xof5hL6Br60wn1iIUNuNVOZeTatB+B3FdNNeICtnlA9yKvj61
x7y1v2TodBL6moQjVkzb8LHTxucoy7zzcstI7iZTbOZRkc2/8DS9i59/i52JQV1nYvEP8Eora8op
7hQhgffYjbQGwDKEjWJ0ZgrAZKYnBO1rw2Ih95jt1D0GcGj2j7stRs6FXymC7+xpnBwotpn/UYbU
7U55kv4iqbSZCHSXLhVrh1kRxkNlbhv0n7J1lRFi7j5KtHJuEqt+tO2+ye0Rmto5zUihtlC7Ur2l
ClGANaMfFr7NbSMROby/FLEgbuy+ts4jPbknu/jsFGLHdGk923uofWrBwi6mvJE9lh+nY6vtOFZr
yx8IIS5xU48v0mGIRS2jv2oL6Hv+14ruUZfRMemRxOM1g14IGt47h/7xUdY3PRGDdAIssBof8iE6
9P1uOXwivPd/QCnrzwoW5OqGfSd7s4X0LaQp3LC1uj/Vsyd8cctqaCkm94T1VD8LFp96WPLXRDGL
jj3f4wgxqzYqhzVfutZvB5IJGMMCSwjh3xq/LIXkgHZ3wejRA9ypfYV2fuOiPepVmvX2p/fGya8B
8lQOskk/B9ZlYxg0XGfYjTwVBR3u9f2ZvFjhw5IPs4andTMbw8dnRdsDbAB2QZ+o9GwnkvCL/K9B
+rFI7CXDxeF1dWEYMSp0cClpTMsDe1YWPYKM2+6yTTQLP8JJLYBc6y5d8EnqLNrpA4jKM9mn/YBW
Pg19mkn8S1h158P96veBE8eb1yOIaRjK5h0Q5LtBt23TPZS+OzcTbwJLUDAljqH1XGE7RRuwcrEn
mjYq7zrh8+Eg7vK/CX7lN8L/O7Xj8MGOzCqPqJ07Ox5jwmjqxNqRLcYL/V8ygb2tp4BqiUTVMslG
7FCfAnRmPkIEL+G3pT6ge8j58gdc76ep5GXduNujw9JwlB/C9Bs/8RqXcs2YrAq1USNj2cxddPoh
IsJfaLhbBgXJ++qFq5IkQfsfX6mN81m+wmamThnBYH5iULqen1mdXhh/RRFdX7D1pr1mbPDrcTU5
uPWFvooBUQMtShOpDsrdzlgjbLdn8nj0yzzTae5Z6Cs7c9mRuKP4dvVlMg0E0DYbr1oXtAfln6J6
cFfP0rTH3sD1yJ+hA7maqKXJ1Pm9X6Awa+zCdOBlKmNrEZfON/i9HiXZy9i9aQyKrKrTymRkAagX
Z2DkTCKi0uCEa0BSfODhnLgkygVWAUQmGPQHno2NBTLUlg4DdswZlYwSsrSIh2/TWlo5v2I1pmcu
Qi+e+XzIa/vuwusjLCd3sRynpN2LnkgDTRkcEaQWWTXqf/6dz9XLW2EPJ8fJC1zjKyraXhrMLh+N
/ZxS6mpug1S+OwNtzqvh2eVXEy4kAyU9ugUl01h/VuTs/RJwA45NJhC8DywLE7yT0abKunXBFAFF
1bQ9xoy9vIQE65BsUjTSQifoUiMFkt9d3yIxH7yuHxeDpLZLB4LzkbAm19n4ipvt6pj8oR/Ww9ZG
segNk6NyUBkfOmhacekfM5EnVLwzh+hL18b15J97Q3dJPJ7hGeAq/ypPVAa76lzn6yI3iG5EO8L1
nb2Un55wdTiFDCAQI48h2ytdcKBTX16FDeUF7Nf1zg/raWm7yXunSLtp3fwxNb9nqQMNfFZJgG3A
4V5dIKoBlMFOwqGG+tAvSKNm9WFDdVBENZ7rLfpUvfd+TI0u/KPH/ScX1NX9HPqi0ZI10pA5QZVd
cNHSy/14k2QDDZMJHx9S7nAwo7n91skvJzkrOhFj8lcar6AhasJo64fjcNrFQvWGC/EDcg6GU5vG
dkylrhcf1DQC3BmCy6O619U3VZlajmborFpe39wzVDACdZdO3CVWZPUJzh3Vwu1hL0ar6Lz/M0MW
7VyvnNat/1a4b1sPZ4IWdJilBlE9xun3wz+C8OlxCrCEnuqdD2slVRVxaxSZ1940vOqgJannRzWV
YnY1O8YzpjPXlxERr1+sCU19Nj3yBN3pzwesndBcLKXm8Yx22Csq3OIdDwhdNnhJj97gG60KqTNL
x4gT2vsePowDUrP9ypN1zQ6thomPZGDSemQvF1AhEN46BNVzZ/jnNLW/nnp1TvMtcjzL6IP3HoJD
UU8YkwvPCjaw8/m1P9oW1xuj34rZIv9vTGn1EwazVo6OSuPfFVn52kzGGHRzeZ9vJeJmFXO5t5T2
kOcHUirMbd0rSanSmEyimgLJGFo2lpdAoiml6Y3wtK/mB6227qJ9XSVvsY6rDNwKzGMJ3W+m5AX4
rta56riKWB/SLyXq9WhfG2TA/9E9S4Ykg8wKs4RExqMKiZR7IPYFCVPGG5+gPoqSNmxR1iCl5RpY
chu+b4iIIjDDupg1YnNJZLiMnaS+E/jlKtHxsGtrmVw6tWuRdRuYyF4jLfYLPB2H+TG3/dX/eV8j
jbmHW6ikEDPTPbNxv6VaVlkosp/bU2mgrby/V6JgQ7XuD45ozuMeChzUGvRmPjb+hEwqBrXHeyP8
ARTwXdviBo9CTKWCyeLmstZjTF+AC2uvGjJM9weh43R/Y1xVsKKymLGurKGvNDcIspEZ29t5CNOT
2rHqc+eo2IVvOS6QJFtbJrww9k2WuV0YHLTt9X2PKdH5UIER7GNJjtZOYJunEN2uZfwdGD8s2BZV
yb9bYiD96zU7t0GuOaXMnKBynSaIdj4jcdWLsSAfrMcbJMVThtg229C8OaNMI9UVL7Dt32QQiXRd
NXrrRe3osT6Yrmz4HG+JNK7mbiDz87GSQca0rlhDLzhYzJE0AFhfQbj//LtIkqANK9nsHzXE76kg
EI4pD7eJwNpuk5Y00icm9x9JMioUbxKT4VaKRMJCZaaqi8UibFqhNCA7NiY3eg7hNcxnMAgg5Qhe
ChPR+OtorvGFcssh4yiMbNrdFakz9brvHOBxOMhPTWu6bDx8r9fYUG2brZg0BWn0vitamqjWBSOo
bG1AImqA1VcA/YDNaB3wGMR5Pm5ACgNJBa9zgXxU/VNCkQNB8EG3CjEpwbrv3pBfVf3D6hItHxUC
4lfWSxJMwMkjrpi1k9POrG+FMa1xE9Q47Zm7kO7/L2qCWt1W9XIF3xrp7/t7LDDOQQu0Bnuj4rxt
ZXlEYuKkK3OhRvZGKRCKlXkpgLfzzN88tNarkUIiOz+eXqr90wqycsK9d1wU0iT3mJ4wHFThdibl
Mxu8gLNMQNCG/kffMyBXmPjljs24Zd2ywPV8VPrW8r5EL3tzUpo0MdI4IVxA/gUfssHQzlZ0MT+M
4JBgIBCJuTp0QP6QqiSewFJ1HH0UvjhXtmbif9OotNRd8dvoCYNVO9SoLX5wd8lxx+cbCUQL1jtT
mhcFq9jWXnnHef2goI22wXxAcXf7IoJCjt5wRKCV7FsEYOhE6v+kB2Rael8WcaDQFIdSucfu/0Np
2cTeUkDDi7Jw9ggWyXIwBqWb+Ac8FNe3gnnV1Z8w4HBD9Rj90ut1e2IfFuNRtCEMl9mzHdwT3dz3
NVeoxQaJlwr1MMfIht1RgZQeUGsNam/7yO89vTWkO4pWrfnTUIndKlCH1N+KiyhK11GBVcnqpJjH
SIO43bPWlFq/nKM12Md6R4lQIobwcOxiZ+XP6muh7XcsRsAddIqhwK1+cnY9gV26AUu0B0YXn5NS
t54VKvubp+c5yYLhMbi0hlbAnGYsPu95ii9KH9dupj6LIok3fDcg5S+XMTyJrYEjZI8il97ESSJ1
bE+Lq8tSARqikeDl3XwMECfidF3Tku2iOPubWAqdl3p8vZ55ZN3MUA1EauK+PNnCc5hbZDB0oanN
4Aryws+7fyAmqqfnZsJF9BtClrdfAplXsWvTZQb/VfoDGNvRK+2T1SR5yTHiKvrvzt4Or2Vh68mD
PiJJOOQdyPTG1C2Rx/woAqe2bY3gt7rgTCKbLzdqyDJb6NRSQnl59k4YNrLepoApNhPKIePk/RzW
ggTA0lWwHbfc6AyCDsi4hVJybrIWonIZe01HxhqYU3qcCE3Q0+wEbf4h8+tVMDIx1j05oU9rvdli
K9PiJ/BLC4UfgIb8ScIxhLBW5KkmmQHSr4h4ueIBtLmYs3z2Zg6W9fwdjFiHAHR5ixzCcssnShcE
m2BBpBAKdEAOSqSpITsDLKjhCCQiS46Qs5sXTVC9eYHhZMZCmVHIvkYbrKQxNLvvuA4xoFpb4D8S
xivTo+Nc/N5+JfNMfIfyCX27GNP2JbeWGXgyJOHiHIItkYEajgNbC9y1l2GZGgsOZ4EL+6BsKOEJ
UHFoc4xuyfr4nuZ/3JiYei8tzwRa2cxXdr1uX0DWfVjcmQU1pP7mNlgz0PBL4BQ1SCRDkCVmNVwu
1Xlux93qzO7atGbX8MgcVC2UyFD/k/8ypA0oOvUg8sj0mlYks8yW9tGXQoRgGbuMh5dLmRQHdOpV
tg5w3SwF7GDwwTywxAYu/O5XJAj45gK6A+LxQ6g+ivE5/JvTXKQYRx8TLWMprptpLFV/heiYouIX
effDq6YaKvPlfY+6XPLqDsSJ69c/AQYC3nWlY/UNK5eK+WjuzjvCv1xliXaxyWWptKkSO1nTUWN5
4Y8YuIG0KF1xsXVyVwjjqixqL+bnwnrnejx3V1gpbO2EA1BGn4lHdjP9hPOu/NgZb8X0CaFVUbX6
2n9iUw2He4upd05yAOjqtQ9aczL277TkmrhEUHaotd1XrYVShYkinSYVXFfV9/I5q39hMN/e8CVM
7ibLHpthQwjW/BbIf5k4QNu7qgcCTpqAfpGFZVVdObCiFzyDz/L+pOrWt2OLcknAwq+RSqDuRbOY
HrFMhC3gnvfBInoYQiogNQJ0Eddmnaz3PC8gc/4PJKHlVPFoTpsWPTXZyEPLEKfSjZjlTAltbzr5
RQBgH4rtmkN4yZKon4t5oAzfgamk+bVjcR3wA8LgFuz6+P1VflQq9alnlM30wBQTZtyod0OJnFh8
chjMWNuJhmDxPkYO9RWKIBkHKfel3UTK0ROISPVMSfiLEhzMvtP/XOcBopBW1+y5l8vXl1BlHcRT
F8NeOtWNxhhlinE62QxXNSBLIzJL6us+OSvWx/QP66dh3enoiLTjraGZxr9/Hhfsg4iTOPmZJCzv
NdBcFJ0YueXlJD5fka4aPTrkLT0NS3Q3RE9U8L47hhA3zi3tTg0uN4Cnomelw/kBaAeicjS7m91Y
IeSXEFoMo+B/GvrHRSOBLDQTGVBuijnAsl6iXrE+LzbASJu3DbY3cr22w2h7GAB9WT5IbQbP8fQY
uVw/1Ywj+jtRYeXXjgcOQSCxjXUYAUfaPI0A0peP50oIOTWVTGjkY8mjZar6v1M2uDWE67XJg+d9
9ZQf0DxQ7qLIwuUxR6Nho1DnhBG+TXURl0bDe5KGpSk0ewNYyK13k/wiB4b6byTRrE4/qUYjJzas
xunXIkDJGV0l4hZ8eUz12YxYPGK6QYQNZ2vUR7BGmamfjr6gqFSMm/te+qDQw6oGc9hQM2SdHy+p
kL1kc7mMitXcfhaSzc4e2w7v7Z0zbv3gVo9wI+97/ald2FLgNmom1toiPZ0nsT/eE9RlaBgZ2zmZ
ZNXTXM0lH+U9wsmydPGVEqPKE1NlFyGeLGS0kMLseD2Wg5DyjQnUayqSfVeX7j3F3oj/BiEMeA7c
n/gKs/T4RQhGMPLi7WaXyzBYgu/WOlJ4pjTYhDLxxsX/CBDBIG0Ywkj+ONL5fo8liRO0+8BDWC51
56Ph8Q7Kn7CCZfPI8mi9IWaYWTculeaZlh27vgPLRjyUCcDhvfnSAbsHf3B8ZOGpKzN2RN92HE6z
/eU+mfjjjsTudqDAwoL30cjvX1ehSij4CLWkfBv6J+ECFE1t/Dwn1p/py1lm9+G/fI7jYsdE195f
vrOjrzGZKJxLXYTzVIOhQvP+HGEspRgdE+JuKIezhwl1MBr5k313Y1icMkN8auXd7fL8I3HlrkRJ
YGEXQXZiXB1vNm6Hb1PsZSaABZ8pRqnxDKeOc2GQSDPGuPN5LKnqjp2zaXkwmnY27LB+ADb/Zhr5
b6d5zAqnDfRLSdrovmUqerKI6iYjdiWQZJaStCgzsI16z9H5/V+6aD9oml2UVwsJYWnAzqfuGyYu
GYkWWLqOVAWj7cbITlZ2sOCl/D2O3G2oVnEfjXiX5cCzvb168s/DVuUnbsq4no0l2bIFRqH8lC/I
U7jQ/CgchyR6CnlJizSHqBd9UXS9DEciEKnaGbUwbm1Rb6c9OUHwEJ7hyRloeZJhm7QCGqMwBsoh
TAfpSJ6noX7pM/2tNd4KIs+eu4CKqn2dYUXstFFdmYjylKXwV6oybOJ1FtTkAsaOcPjTkCoiwsHD
1f2d0fTxFp60mFth/ucPjaBYM39lJ7NAt+HiNyockR5TQr3h7cb9KmU9ZpuTSOKAqFZTFMdnsxUp
+dfwXSqPQ3dWvDcuBf1Xmv3N05Pmce+n2jtp00+/P6Ysn8+OaZpctxcYkkuBbxfTwhSadATZL2hK
a9SnKdvoSuL8pJiH7yQCW8seFET2co4Q/3HOLVtbw2W6+SPhr0pIXgjsROaATuUqRM9lTIDH9XsJ
zBEqPkYmFNZHJWwb6ouVdi7Sx4DbdzsAQIx/CzD7OHNccsIyhFSlA1mon57GgvBqPHSkehScOeiY
XrlLNAjDuCysI0uWaQt3xtmC6AekQuCn7YS4i7mGWQSa9G394g+O03Sb3T16hZJ74RDX5OXRgPXr
IW9JE7OOBsQHCAS9dFUn7OGUMgqn5kRxW1ejSBeAHDrH/XQVwZdGQPRXHFW4IelXS1CP037l1K79
ZIQT/GjFQ5IEWQMGbB+K3rqKj7M9zBsj1nnypzJEniGikBCxfb/cfhhV/CHur/IyyNU2K2C4erkc
XWOkXGGxlWEo7jRmaxzuk2oiZn3t8WLRdON+VaREzQgup+7bxJ3vwPLIqYTSm/bF2OR0kTDgnjw+
tYTAgH1WCw8Tl4BGN0400PVomQ6GDGgQQQt47ceLISw1vD4xOl1Pk3HG01LZCEXfdTlPAjUjBOFn
45pg5SsSD0eeCR4rrviAlgm4bz83w/wMtv3ducgqZJ1AxbqWe+EZxepnUqDPeR9/s+/sbrsMGZwb
fWUIWlj/XUMsDQwFGBoF42cRztcl3L/iK6MGkkL4XnD6jfEYlFmtZ3CNVgbJetjsSXrq2aWPYAJR
IEvfjXSP3Slx78J3AVsFL85HcJ+pzfCNQ7g/3Kff+M9+LfcoxOE3eEC7scoIaEGzdv9/YRrcKof7
LOJYMc/el+NJ7qklwczJRyxV20I+qHZsWxMwcoiuwEoeZrGGbUjgxK2+Mhut0lObtynzwuQrQFwy
3U2Lsmg68rK5iwLZgAdQ5qXDRqMZhMuJpUXW148pCc12SQzc7cgHZ2Pu8WWlHnQwGCKqS0FvDyNR
mPoEhvIBfPdnUia1YFX6rKpl2ahNB09PsLiM5N4nArK99Bxo4DAGVYfFx3ihpZTdkQyWcapRIJty
vg8ttFVQgnc5o0vn2riCArkeiHFwzGzjA4qHCP4SFjXpGDffS07B3kvYBF8se/e6hIJcovvN/eQd
V4YrYqQ7kbXRcP7qnvGhQAXMITFwDpjyH5k+oIhrrvJbIu0acEiQobV/XsrypkKhwxFVtbUenPGl
2vP+XN57b4bSWC+V4ByWtiumJBv9HZ0wMiX4J4lC+1Owi7CEbLHdFgUe42mh9LKxrR1Q/EFshdCX
uUVlcVHF8+6JPrWox9qFbfaRIYvenDzicVHoFYNqrGeSz2+/EWU3MrgXsquryLGvOofQufEWcfm9
JIcGAOatNahkAEAUgOtaS1vcLTkeV2uE1RfihvyW/daNSbmCsjEn1YDD6g74lwcNmP8MDEUw1G5g
t1vz5nbWFJ9wvgGvLqFNzUNxDfNPCrsVqUuHteQ+ybZorjslfopQZYlddpv+BsYHfzRswLsncwJh
fQvSr2GYGc949s85m0KAJ4iPcy+47wyQ5rYBQ9hBrbQ3g5o3X/DHWqxao6A4SaZtRnTXkazkqqGq
mNmRgSkDpYq2rfg4dLyYmiN8Zmbjs8rcDN4N+hzNzuLdzKmzdObamMwpJUi8MnW/EiAPWQ9Q3Tou
pEJgXR3AfXeJS+9ITFNVnpE4DgxVMrHAybRUF2tbRaFEYrfoYTSHuUyUCXN9SWNPos02D6Ycco3R
Mz7D1Fd/Gc3zOdNRrXnhSgtDakHvStY1y5FEmOyfzFQ9lW2527tYFeWdRIm43vfZb/SKnQPnRKo/
V9vpTr5zBP7TnSwx2jK8t55InhaTSC11W+H4nMVTaGr20I+4efInJ+abop0qCqdAPGGmd/iFr0cb
yLySEyt0uzs4xAnaSAu8fMs+MlnrtFVoATiqDl+HmXH2LBfNxUmBCnqcIrYMq2/A63aNQC7iuEz+
TBqRsbfhkr1o5I52DnOe67iTPYKTQrligjnXaddyW0ImAq25Jyz/jezbs4hnQ78iNQuI108uzr5o
PI+jQ8+BbIyFnWNDTx3xmNWYLigR6wQ8N++wdop0oPVCVIkST0onUsshvHbGyJV1hiKAcTtGe9PX
DGpxB5MpKvFK0cDDlIGbaNeAlru4HD1TVHj0Gq9ilU4DkOQz4joHqGgWP9SLGDoEB0lYhLHykLdK
rqs2zARCtL4KzUYylBuSLX+XsoGghpB7YMcDpOc0i9TSBLhhfvbWpzd5T+9vLI/vmU8VJihFww9y
XuwTSBIMLqGUETfW2oEQDgR7cj2TNXrAYE7B1z4Y1wbWdyUFUH7lSS4HNWyvqKAqMcg0/iWniKIB
VRkwWH9y9wpzb6WKy4iLQO+c/xVI84vQC6t3hwYMuBd9O+aa6LQTnivnI7ZUaL2SMcD1w3EUqaWs
LV/vP620JkChD+8/sgyiWMklIH6s0BPr1g5FGuI5f84/UpZ8nBUVrFOugrS8WP8ii5xaLTJzHSOS
C4KXT1AaTvDEes/BahUD6H9Z7oy6CC58zU7nfezu/u3ldl4zzsPDFNgMDp9ht9X/Ha0nWHHeeycH
lyxwJO3EI1LXNOrVcEW8j76v8KYxmRcOqAPZOWdN7uh9IgEc0XBuGNRUYrB1ruUiBclZRMBRKBp1
WdJCk72RzHxcEr0b/5xYUMxTwlB15kkEYfzhFPMVRfLXTD4XXGMLa+Yp2EOlhciuozZFC4ZD6Z5y
lzDfU5DfCQ0M51YWvCBDFjY82MJGsEoh18L/294M5nZ6c6eUh9pchF1aFLWRzWPj6MMJu4dHJye1
k93Zl1/0jFy8+1jj4gcGsvmWRBipQHutnO2xVBL/FGY+X9PNj6lnOW6nWb7cm8pe/VLOWL/DiWLa
0d+Qn/UlBC+AzIaRNIm/L6g/pChrDr5V+YOgah6GZ/qT0b3P4MuUxZIHYPwap6I2kAOHv/uwIHV0
e1GRa/IcqIcS20tvnQ1Wm73xB8TFtfoK9m46GzRPQ795dZST3skfXyNPR1bEOnbCn6PXKqh9YflQ
xnSF65jULGmrp/BOVBFAkaBcJb4y6qqd+x8Mt2VgF93ZRxFEJYwfy3qKBpCeYaIo/HUDE1muPN9e
Errztk7Mdz3jSDS5cAolZKtrT0xauKD9o40gGD5OrnemekC2fH6JVGaBvHMksjTMxpgaciiUzRR+
YwZbRpe10kRbdee0aEvwLY5eCCc/XUecLxunugnnNUyvirYAd5/EoGELMTgx2eWM3O3had1wxy6k
uan0ilJ+PN3REdw7NAr+Mwh6GjWEA8cmhZDg2JQQROJj03PiOGcMhkl1FtviTV4dXEpE+cEkSCnN
XKjDiD4JuMpwMpHO0lzSkWV/FW9GssK/fyfjdjx/PVBg4ThN+ySmQOHNFHr46uNl/xH1oEUeiJXv
XUbTORcOWGy+isSJzKjLIlEy/R87tJ8bavbLQtUtvyZuNa3gALDMEOW92VOo3ZQiDw2B9B5E/FMe
/aDW0YKip85pTY8GOrxhRA1awHqc0pszxRw1SNlsyZI2wPNt/tOXOl6qFHDE3fvWzPjoN8TdHCZF
Ck31lx86VxSeBDC6Um8ZfR1bWzLmMPIAcn4pIbqXIlWPG4Sg0OAgHRSQbz0aPtnEwF8fHrxIjKog
9fWqEqUNvzB4WJE5BMeb7dWhLC2cWL6GNB1tVCvuUV0hyyr/sm/oE1i87smkRcn6RmWNUoPyN0sh
qaCzfqxcsexbk1tTytazODsh2JRN1A8uLt2p/DAqbHWzFq4evUutjtlrQ+7Mjzfirtr7uMPi6yry
tMdnlN5gIayMBnHyWLojEbeCCP/XVL9IsPJ34Z8reJJljUMmHB5jksVVzUYw8Px4aBC6wzO6wfPc
6/JFPtvMB17ETC6Pjp9u4dghYkZQ3hzAwZ0UEnTPFOw9iqHl+tiZB5gVgUe4ieEcABEudfePxrU5
jlk3f6xM3DxYIdmxjvRccfRWHxIrCmkij5Iw0RRbU9a9HNNC9HS7qjAY+l3K+zZ6pzfTqZblgoNY
Z89uKSt1izn8sWVai8zvBfRMT9zWk1O9YnRgEls3NJwpYjS3E+ickK5bG+ARbSgY9NcOA+iUfjN+
JHCX6cg7QYGoW3xqmLocplznQsslgFJTCDi8AQX8rBd19pSHnSKmsFFVPRxVLXIvMeFrQA42DMDD
SCsl1e9Ii0H+GVDYo8oOmaAA4oie67R0nDjCWBhInGLpLnSmACuprB0GzfHI4NDzICwXf97h5vLn
Y5stLu7jJbG+wy7gYskZk6E53PDvn3k/OmUXp7oivJOdntBWmD8u8Uty81/L8My469leC0WxAyXb
xLIwTY03+GYWJs/Uy/q+E1Kb2I46/Xr53ESKzq4icIPktx783RFUV9ycGNwwXejIYYEPJKmPXtAF
HILs14oVs9iI68Y9aao5pVoLKXdzJPMyCyJS4Hml8AraDC5x5tAodD2zoay0QkirXuj2ZcBFdIeK
z+6ZT/a7sA6bnnHEvLw55ECjsEUfTeE2i8XSjK07+2dOwo3T3ShBxXDbOx9aG7j2VGrbmph5htMv
poubgL1ZVcLQG8ek/HMr8vH3VIzuPE+zQb0eJqYWs7P/377wZO6ZlM1olgvA20DpGxjQBiB2p/FG
Lqz1m7cNL5MUS/p6+Q36AUVXxyA23Q6Sz0sIe5KswiCL+fNY0xgtljV75VwLAXkeN+z9xbMTfqcg
xRc6tMzSKHsMsx2Shuox+FKKtO9HOdfO2HvFGh+G6EW22jNcvFzWp6HMDY5fLaMDw26GI/3/CuXP
vjUCss6dnLhUc/2J/v9abi+dMniTOivNoSwYMKfV/w+oqUwRTpRABbucqqPeiWy2QSFpV27K38Ku
FJQKqy1H8uW7V1724iEVWtwzzgNYWSK6NYcpFjgw/mQSG72LB7s5Z++A/qfAClUApM7a/UhTtiFM
PbfSP+d52F5SN9GMMVZ/qlCoI+LZRV77FDigTU4Vv9z6iW7b0e1IHHOY76ryuw+1XNzEYuVUFbcq
XlgOitKDQDvjhyYPUCilulEW1z9fnFYHvH5m4SQwM7BHGdm7YHbbkAiMCbS4pNJhdmbmJ9wS/Cnu
kDySzm+XevRMq8oT/s+4T919Okelx1JfxEw6GPz9RuMVBZq++BJ4mQxMpBvqz88jL8NdNAItdVPo
/0vxsKKOUSsQ8ExnnkHV9SFFElI336rHQyMBEwgOXcsuKo3q1xzUHsKmKrMM/hVS/PtqSnQIck/H
QU5sUpDpwYYLqKgHuhcZirJlkvc7xTElWLu3k1dboOEbgueXp0T687cW7lJMxGOzeL3C8pQkMlra
UVMqj2k2nQ0IzuBi7lJhUCkj1hHLO6KSoRSe7S0Kti/PGV9yjSfhEwHMzj2cSnf3ocAyaqoP7AAJ
UbAiQtTJEL5s8DPyGwoQglr/SdxuQALUfNHQJWeDIipcGBvbOMoHMxHZNlh4CtDn/48YPWvhzkGq
BC7ppXugkIrAQhRmisHY6mf7dDDTdxT2Uw2sTuAzVplTDacFo7rtsjY5tlMLgFCQ6A+gy4lM0nHE
5nBL9E3JRtu5c1zuahqYNTuGbifJCkbS8682Kex1ioUBy40MFkIImcZ9mqInY/svrHmQMEatbdGl
qCrOhUyxuo3CYIsGWfLjxn5NCmnatvalvYkUq1YXVfEHN39E9BVg8LAuuGQ+V9gfI7VpMaFVPDuk
fW7O86nknOLiw0Yv0U4qR4CnqTMNsI7qU3Wqm/a4y4WTCYE5vMOcHW5iddhwjz0Fq2dDlSoUJXk/
11fOKwA21d5UYRN2BYSR9q+sqTYja9g8hpTKEbLmglscl57TnPJbeuKCnKEE1zI55F3VHdSgI1ny
34auY6oeOiJiJ8ZiZRbsSgqqa1kfdi+d+uh7pN9R1mlT9Uik5Y2mhc9GMu5rCWS+nY9Sg6qBpoAV
NewaG7id1aBFdUyMD0isyLCSY6UfOimFVjcDYRbwsZGNMj7yK3ksH2SNCoNRHfzZ7mYBvOxdizTj
efDNQLEIIw7O74Esf172gEDbJ2EYI3FOQmI67hOx/iFsrHasgvhSFsTjxJ3MmLS+2T5QNJ0UU0Q5
+VZXTJVXyw4Uji9k+qSuoVPmqGR1+158jdYqDK2bOBbkGrb+3tisxRxMRjVaY2Z/2pHtg+aEHRtR
W4zbcaHliPr3ZfDoynM3Ftf8Fph1oIhsonZzduMNDcOcrgSK1Iphd9sz2P1W7oOOYfKw1AF6gQnZ
vda6fXjBSca+F5PZ9NqSWRMcel1KSM7BcHSn2vkOmjcmsWCQSqGxPPk/Pg8oqicXl3RMIR8n206P
6dAFHs5pe8Urwbd6oIQVLUmeEpqzMBLt29+qqntHxyqDrNueuUKHII+zsyUpuWwUjlQ2CFeMauem
HN8zLcKf1YNC0heeYMWPGlWWlRQIa9GI/TQdEeljsW8zr9kyDI0EC2wCRTN799YqIf+sdV3sFwJp
iQtzQBJFc8hfPrIyzeXRiIaqcJuA6KE6gOrQGUp81d0ktEnE/lq/fsrUbsvbfXvwcuAf9gY/0bIt
fSYQFEyEnXiiM1o4gwFQ/YXoFReAH+hu/4z+QtUQBVHrScn56rFcCHb3iuhM5x7eRkXZU0lRgtpu
YQI9bmEOJ0c4ZX2A1iKOQ5sPdTflRVqH0QpOsf+mZH3MxAMKTd8RjoDst5LTrFr1bVmUAXNDF20q
cNlLpc3HyJR2h8wDhS+HJetUaijUm9p5Gq8ZRZtt/2NrRDaFgk7pmuBscmUQT4zFd2kzoJv+ZkKs
mLXe299URm9TUEetgJDL6+h3Vs6jPqZiSjJm6cObrQ/yVlEsy3kf8UnmGT+hUQzGmSff9dGqJmtv
x0nJ11cLLjT/v4JeKr0NkPhgwJ+VlwgS0vZcVNYaoN3t3mAh5iBTQQRdZHCt0lqsyfXWela5gk8c
a7vWMGz6wNASdEplj2GANwKDXKid2tMK8doA5kXY7RzElfrR9nW7gMov6fM7jrjefTjbmvpm0aqe
oRplfk+WN4J2zDA4qRRC8OMD9ovMLnOPLUgK89urx3iyU3R+IWjx1/H2BB/PnKjtAAERpP6Riwpa
YHunSXGDWfvSd5wSpoSRgn6Lrp33gnp2ysPTqRKd9bQg2zrof/9ZnZRMtZn546KzO9l4d2bnqKsM
wLuQLM5knTVlkUinTfyKEewx/++aMhXGuObZ6CagOt0aZv41eKnVbHxWgkQl530BlN8M3kow8XAx
p0SXQGQTBS7bO7kwGJ6TBHHudJjekRCA4j1LAZ4iTbf6Ix+mA4NN8E/Z2j1+Rg5/8TIctyfrfRlE
ZcAOFNSmx1tQ+q5HqvumVerqfd+vaf8MKxnzjDcolOwjMS4PT0DjZCZGqmDQKloIhprEAxXyZL6z
AZcjx6+xcrr75oImG2gsQigDTrF3/6K6lZK9ZCmDeC4BY7NLxTeJPbTLkEdz2FSU6OG1lb5g/YEc
9+NFlXMlzUHp1yH+0BcRdAmE/2QBFutHAMyddLBSEVJxzPa5PuBVhKGhA1UFL2lwyDdPJuZWJGLd
qmTTwGelt72j3WAdHTJwyVxwHxESL1/CNphequivpn56GkZgQmlMLdqLIW+/w8yfd7ILL3pS4QVG
fG3y4x2yBT0yCsP6Stf0DtFmrRrDfdRoS3tMJSDIWV356TXBXd2144DqoKohpKnDvvSg056ydnC8
7vzmoyN/GEVuoTRMwgsYBBzHMHJ2w4RZJTXzSfP2kt+r24gSOCKmVlIde7dxSCT8zalkWwMbPukw
s9puAErLMzhUsVzAcU68G08L3N0NVn0qZYhbllu3Ha21Vd6ih8IYHZ8Gqtxqd1LyHMs8zHDw3fMe
ZYfqyiGhEelaoxXhysMVXflUqzcYVXxZhx9vM6XxxXKFBVSeC1MBIX8y5exMLMnYNY5YoFiwGdGU
uhG0VqxnlUEqh0/HOIQAwf2Ey8YHodfwWn3gqG6s4aopKkK5yEHXHuLzFQ+pG4QwTEtlhRaBzL+b
GUgXR8FDQshbhi4if5O/dTds1Vsu+XHk7+wsMH5srD82b68Wkdpf/5lhVZC6EsnvU0kk0Hgu82ra
l2+YokIMVSXMrYCJYlRmrD2gZn4eBXHSpjCFdEdABx73aWnJMGS9Z3NaB2JzAURk8oSU5KhLQ1rA
UI/eVmG4G3lRBbXifmarYm7fjaEfLKEhkiTPKHEQqMbaA7kQexaU6NY+M7RTXc1WK6JYVgnHk5hL
xYcnkdKCft1x1lcEIfAcpZOHp1pk62+CuAqd1SrmNDffiHjB57CbSKkXnnee2oeRjBrSYgcKZsy/
IXjb/0kG+nyTYuzdYG2VaxrV776lSQtCcpq0VOu46Dcih3MZDfFwa+zVFsdbT7y/sIDXdHVkRIT8
Yy/NPb7/vGR5nE0Lcy78gNM1za0QdQtlLKfAAG+HO3YvskWkgs92TeJyZquXiR24w2FvnORSwj2X
ZyuBk4TKjyYHZnnoUcTjDf1E9/4OST19dk6hvZYjYD+YoEtdTrSVR5lpVc5FCVCr1M4frgHposGM
aFslPgSMbxGJyBGT1vSCm6PLsn4QKF4wk2g4DVZ3ObNzlt62biyhuJTg+MKzAvxIiYA+uFJ/woYr
rM9SOukrLYreiR0uRl3FOsZVr4OgbubUwUuzRQsKzhT8XSpDVZq8VqAgsvJ/X5B48M02lTOw5fuc
6c02hXDWJ6NFALVQzuKkOU+AjnjgUn9LyVlwhHPdJrM50KYeJD99ewS9Z9/4CmaGhXsJUSgcOAgp
3eGiwubLqjqOgu6HUamhK6c41A0gxMQjuzJH1zczM48o6VdqMqBvBOANwQUczxx2ihhvq+cG9zLN
MvFC4fJT13ZdyjTY0tss/wcq9elfmRyh6pmmAN0I5y7AWBhfV0x1pQ4QUQ+kkSc8agPecO+HYK+5
PYz6jqsKji3OEJd0BoDECB4YdUMKoPzzXhjHK9DISmAvCP1bcelQRviM3q8VcCtVkkg9Rpl7sDWK
yi6lzBha55s5rKimtQABXM80E/gOft6fgzqcpoQz27rCq4EcMWEA37A6VFubatLeGNSxfyzCMBhn
82fymYtSCWkoE1SZ3RnIifGbYrSl0hZUaK/1+dYk92l7usWSzhDdWl3LRhykUwDlP+oaY+6jk74D
tpsbHoYBhFTwFECwTyH6BuQtaY55ZDXeg1DCz6WLUwJjkMA5O3lFm1jU/tF6qctatG6aWURfdiXn
tOG61iiM+lsg5cTCaPlPJ4A4AbO8esqsSh1SOpapoEMhP+dbv7DJJBoFyK3Yo3KPPTr55eakptyB
8hFgOkihP96+sgSnsPWZypFePdW/XXdSOQSFGsgov2MnSBLF2395A4fCoYDekk0ixkwfKUyN7ixE
bRDcg3b9NNbRduLoM5AaHkGs32yMg2bmZFOAvQfjVJDAgGoHtdLyF43X7sMB3nQuJFkFyltt7AOI
wvKJ3m3xZiJJHrTKs1VGO0H6GA8+9di8L5z8j/epZZBV+SII5BbGTUyEstA8wkTMrGZJMQtpmyAI
FVCpoNf1A+NNvQcmICtCBG74hL+Fg3HSb0lNGFpIYELoBO/1Zly8IfuXst59Q1V+dv3Ex8QLkOF0
WKsims2FzCYywrVLhB5v9v7pFoIYj1kqfxD8gTj6Ne9gkynByj7ODzIBGE8DS4wzQoZzN9fGsZsM
UxsCBFWfvXiumEWOhTDyBucfJ2DWG4kFvFoUAZTAt3ZMYhZvGgr3e/28V7X2JfbFN+JZX2FPfLm4
3/LJJ331gnJrQmRpRxnBETIcrvjtOIVsY1Q4CjED0qOXP/S3nDwkvHKTQ20wODdda27/mk1SjCWg
JmftZE/EwKixTRZe6PJWv0yeQwdEd9ngCrPNeY9EhgKtdhSf+myBSNqKkip5INRaf8G7WBSBgDmx
fVKkJImWuHd9yp1aq+E/+FMavmGqZRWhbfHFpt4KexIhfa8ORcYDhl/p0ewuAeWrGO5AK+WbDoC7
m8fox56lvacRC5jPjx+bZm1DMi3I+PTUIqG1O1dzq+OjsmsFzJpdrlhnMZghCSX+Y2eBcwAXDrur
HlQVsR2EpvKMV3gzjOhDiyeJSOGc23GODzXHsjylj5kQ36pivqeX92VZH6srdvRO2a0nVTK+jcPK
HXikXbNdRW4c0Ct2e1NrNhWgXvo8tYI6B67GWdhvf3d6LeZP/9xeeerX2SO9j9BOaQOvBhNljcrs
eMIDZAihuLMQMNlkG9caQt7Z+oqAJ21OE+KpcQsJYgry2Uk3sdv5mOL6q35zp4alXbhp2Bxld524
WPXC1HY7SJc2zQTFtDi2zplMWlWzmbqTj7cC1bxroi7Qwns7bmABbHtXln7iAh+qcdWSiT9ocm3Q
LCNhpCc49mQDLdMlwsLdkoI+UK/nrSe1fbXLttxGV1MExirIz+DO3rp9ypikGfRHfjBdq8TFr8J0
Al5FB91YIK3SmdcIByrdY9XlGft6Zh8U4C5tOdgMakp3zSmCt98fowszaEwo6NKxB+RW2ZnOq1V8
kn3N9giQegt12WLFB/pvnuIpbd+SnSmFKvfc4QRRWbBE4enMqu4UasaSZtKMUqkaHLF/8DIFNZUQ
wyHo85XwT8+3NKgOKslKuKyDBA1ngOZfmvQLBskcRve+NJIo19mBZcRjcNlkFuCEg0idLIZjXAzU
GU3xDvcPMQZicc51UoWGOcaqHoVltSaA9OTim5TJwFMiE+U1khMAvaEVEQKVdSfdaYA2osQRxy7I
O4t/sINOHnKawHPufZnJuz1Z6xjvLr9/ihVFaMrJbDG3nFjMHl4oxZqYy5SN2Z3VEn0/sqowd95P
28vSGcXxYpnPViionj9hXWfJaAVuaHvG7gy+UGwwX8uZH7k75avbHPTOoJqtpJJj+cfXmeA9ZEIW
qID0V3vk1S5N/UdgEIJjZV1hxxWpBCTzXGJoYWbKTX3NNOIwgAeiD407G+9PmFveUqoXEkxTEeZz
honiNMO6e4FDPRXMm0dQFe6ViQQJLH27P5pOUA/0M6J7eZ/XQdR89hITZ8db2+JMYicfoLD6cZBK
HL7GOytCkpJ+Cc9/4RcAdDtItk/pQtClwQS4f9be71ORhZyNLWlslgZjb6HXBL5uujVoW2cGbtWA
5kYchnAvnjQtKehx0NWOT7cllvJTEk06G68r/sPaakJpYcTPEGeU63kS33IJMjYQHoGQyZAlus/6
dNfP5rLocTS9bHc1nSoGk96MPVu6SWfscrz3tI9sobY8VLF7xaLq0Zl5KOwyZn3JA1u2e87yRY/p
i1tiuR+6yJq9cqfHO8f0/EtNYeYIMsXEvTfGfnnqJC+6Z790kCydCcdRd2ktmYMuOJqaevNKNWLK
CG7s2oAwZnnUCnlpIoTFByP+F0gXsTgwbavqVMT6cXsbR0TPYId+Q2vTwr4S6hRHaXAWol28Y94b
uh27eyfKT1J1vgVjRUC4T4v0XOV61rtM+m3C/tfBXMTgL24HqPteO9A2pZLUSicUzQMiwh4UMR5F
4bcI5D7dT32r7yXNxBQ3vjzBuPTznSO4RVd9Pw0HcLvyv1paO+qv58Bu3bcNtK0Yk2w3Q1Cf72HZ
r0dqz+JNx55bH+fpbG5EQxN33xV6HCg4vuySLqw05PwA/XbhcdaGPfL9+YsVayhw7iUggrkWW5mw
wTfV1V3HlWgqgE20MM5PQX9VH9hzlmO87kPXrks23wIOyTG+k43RT2mv2DnqYTEMidam521K2GWy
6bojM1JwCIw23DE1KjZ1uzfSYMEIcIdX5C/DgMcE4aa5Hb99qvbPz+U+XVTeSS9837ZauAdmyxho
bzLK6X3wfYQijf/ZytOLJk/A3FeAwgy8g8NIscEc1Iu5F4SW2o4O6GItLbdTPvlKokg9zqv97eY9
etAyk0IFXo44Rzi+7DTbBk6uQjZUIE6jnmrEC2gOd6dCKGXnyYnlM82Ekb+qVVT5tIhGbp9hSqEK
oSG6u+fhe2vWW2B6mK164YTYvL2svQ1AsIJQA+44LvEg8xGWSHPO4WdWUSVMgtvIgv1DfF5S2MEW
rF8D/hdvSz1lwKQzu+HTaUnqT4+lb0VObzHOsp9roYklhN4E1jjn2ipllmF7FLxFEPyr0EV2lnvt
FzK4bsjHVO1hwA5y/m9QRdGicYoZ3maSJEHsG9wG+2VtzHsessZoYsLWbiNBE0bwsNxL74wNNZFR
O9Pk7A36peApQkA3OxII3QgO7ozhNyiA7/mcYqAxQqjouAmk8hUeHrDTA6AyfgtbtDnJ8BANF6ll
zC2QfZ2jS/z9KKZAVjE/QFFOkl2eFMghMIPOj0q7SzT/BC1oexal4wkbKjl2Ok7Dr/ZcGjf+c3/3
5mo3ZY5HjDi6FUHNwqUjz86K2xke53zqRK2lTZowaOGUY/Rbmoy4uvQ2Fb23zW3DKOusMZNx8nbj
w5ZuXarN36eyLPPsQJZBHNQqcV8FCz8DTbrvsbhvH8PfNlNKMp0dX29ztJIFP5Kazk/rhDLZ1Gq0
aDspE1/wbnJPK1Imnneuy41i9VADrVZ/Nw6xd/uucBYGwPCi+Ujpe7tKh92KzPt0XzYSnbZIhsiv
E3CK5SLtLQoJABmL4v/7ZvI0bYA8cUIa8Ezio4nbWY1ehKMVi53I42XGMwU3vhH1cXsI0yobtG/L
g2y8nTWkfWYqLqcRQIcjRqnwp08vm1xKGzFXGsyymU/p2ku5jqLxtdBz3e90AS6s9EPfdXI6s5Yn
lMCZvOVuzP0+bLQOYoxsE1/crqMg97wng1/xuLAqynyCkYvQx1WfbPnLEn0JOPk3SQDgl4/0gg2j
YAuDr1t620ASoREjnYGAdM+SfluTLXZDByt2Kpa2u18OapYhn8hJ1m4WkxvP/qiLgCZl3k17ROpN
vNR0zUM0vDfeFXWoog7nkhEVNmpEuJi000e75WZD1fxpKXOzCMdChE86mwaUk9gJ3uoRl5a/Tgpe
+9EUdyWG9iS+PJCGcaB8nIGCUCfFA2ppad5cDPws2VjZ+AWmcVAl5H2Cw9Kg/36x04Co+9xVZpT0
h/1dqT2yZBPZLP5cbkpnZub5/ydqC1v/g3Jtv6civo6WU5oMHWIJVFlgWXUE9UJcfdKOazDUFMWx
LhvpoOYJyfc3tRmhoBcWqXbWHDlJhuuu7RvVuudK2abatzbeYMeamVW5Mk1SPCZsMNzG1VrzrGty
8Hfbg2RRdEfquqpEziMVJ6kp6FkCBBSM9AIiZVP7TssmK0eEPq6kaphTbKGgyNx0ydcZ+ZUnOAuq
+peUmkuExB0tW4fDSDt2LsNvI5fXnwLsvzw5RkjmwAepY54Lwpvejq9nUOKvduTH35yLhqVDPgWe
ion7B3o+2RxTVEYEVEkyIfglhUd6YKhph6LQr0fVLfUZUi213S9Z7YFg1PQsJgOD5UdDXXivvbHt
Nynns9pbV+cTlrhJv/VS2ATA071JbGopnepeyC0bNRXJ7Eb9OfCUS6tPLhMOT+QEhmfbwMPIH3+M
iHAYxfIU7mlVF39mh4vziDbAoVRSaFh5FZ/NJtDkfsdrHNXyhD/oVateNaFjVasmn0qkZw017oS3
8tZpICl+06VL5GwjfwSlgYKK09Dp7m6jaYTunAhTkK2A7yV/BcyEsq6aLMmlgbyI42xNph+XiBpQ
WkiLrHCAoVx/Yy3RiH4Cn2tsx+WeRtydKcHzTjulKxxal6uSEMF+IiIKpyfj6hbaL8eP9r9E5Huz
0UXxz1W0vZNPrmLw8/m2T/T5kK60R0yq+4i8anMyTQ0T410hrtQevqLpNSQnL40RSqhZshwsuNpJ
pbUWl2nwoumT6UpJUBb4Uumjf0BBG95Sbqk+6zGAi5xrOekIFh5dKgYuIz1CZg8jeiDyxPpBSebR
qoYkseN9OVaKNirA6d3fCLc46t1jADJe+ILXTkKYIlob/Ka14NpLaO84txGPjMKIAfn4Gc/Iy8F8
zdk8NZx8Ks3jCj6k3Pw+5Q/Yn+gahCiCbXHpARI2tV46LGY0+2YrIMupE9hbXR1txBZglqfnxkD0
fqgKVLPAaZsqvkRMsiB84qECZynN3UcBZErGQNGSUFiFyjpFjZ8dFmuYbpCRUaWGl5tzkdFEL7lh
JSmMQBnape+/pZZE3iBIweCWuBO/35NNGY5HgGpOaU6jgCKm76Tt6YsQeOhPOhMg9rOWn3EDo/tE
XfX/hLECu0VP0tzxZ081UXFju/NN4R18JeHyynIEjcwKx0cke7Qxyc2n5qaEO/n6cLiiKwckT/ZY
gzW+fkIdQvCRD7mURhnn73xzEZoaYPtqztUKktU3PAv44GgjQJmXGD6Y2puuQwV8TN3gK00gPiW6
eBL4AKLi2KA3vgv49sRpHdoJQG3ObvKyFHt9CsbhlpQjx58m0N2e1n/Qiz1sKQzMgd5e9Q09g+lj
Ydmpx5+rzfGlY9q4xUYy/Ji3sxpf45ePmsic8gZAQmmUBJBxiahaAHTjCV2zeIOQYsCHT/1/0IwD
xffQF9mVxKZwF/h5JnELq33gSaUxca8yS/2FCgsAenP+NNre8dqGkjRna0hWfXfuQh7K99iAwRPs
BIyY7p0m5si8QE7q6Q8EMgJWKw5bS9ILpS5C26fzVBUWRm0yAUlJmU6BqQU/9yYC8XVorwU+jsuy
5dwv+Mgx8wr+ocuMOiTjOqps0sU61aVWiIqgvDbtI4emuUDoLfq2z8TEbwT/yF9GbBfNyjZnLus7
G8FtBGD0OFdyfd0uALQZrCdTL2Pl/Cz9iNM/y1aeXY5IAEMFDEwR8xzShIilvP+K81NL2u1bp26J
atv21jgTUspkejXljs/eXU24efCGLzaRRZiHlR/adhK7U4TtVxXxVxPY2Sj6iEaB7KywAgEWCVOC
/Yn+nkzivAn3HagpEWUJxMbtfTZNPrweYloxmkm9j55l3/iqu5vZTrKdhTAiTMCRp9t7D5ERY46E
nWi8dJgAfr8X2fL1vs0ou/WtgYzdoi8Mxor7kJA5VsISsRy5zkeePv5Aw7/Y9XqGOhNRSc8SMvHQ
QpHRLJgrEuSAcdbZ9etYoWwUsfws39b+wpiJ+QX4qwabPxhasOxDR0gAlkrBWdvnhjwGl8QpQDmw
g+Cx09Sr34U3yDepy8Q1PM2sTkthSTRLIO3VZqvV4pMRCEkdRUNRc0Tr7UV3/DKbM4g8pWan5+YY
U1fXbhpUyO6xNReHqAL7leNlXCtM7AtpaF6QpUWJCCMmDd5CBQIQJOkZ/d1Wsu5zRJtixPxWlpgM
jq9K7iAEafNZ6xlrvLF8tJYK1Uefj0Tz1RHbT1635PRv+Z1G6+P0q8wCUBCoaMKCUD5HWQQ+scZX
ua8tNPWl1dTxJgpyZZHSW/KFEQupCWaA3ty7LCecYyOOpw6cdTmDQNT4PhcwCQwCG15F46wY2QW5
Wr/racJXKYMFtXIldj7SZisypjYgRx2rtncnuj5d9zblkwxxux4GKkbJSU5NmEVo/TZh7svEorlu
J/k30WUTOWRhPxbW8fj7RI56YY/aINuQ1Ix4EKgXFutvp8acmwiyKYJTT79acgNPrk/ZkOY7kjdF
U8UfpE1yKGEpPdvYt7w5dEG7N75ZbULlOGv8UHaOaDA+eb/4ffHEQaXpiJLC14Bt3x9fEdjr06+U
GYXfU8hpCcUWMmuq52V1aANVoJ+RC4yvNpLygaRKA0OTJ4rKHs7NgeVE8Kg7iEHe7CtG/qr3XJ/9
OrP/m/SUxywMjdbirt/3Kp0+0hv2jC3DAEOxVYjLOAYw6tETTixwxTG7ZPnFmucdFSNoCclmMusS
jVhO+5gDZhaYht8HGQXR2/GW0owdkwTre/yiezzO5U0EmX5NUoohxTfOg4UY1wOYgGAPr8mtzOSD
VFWqitGR8m91zxlNcta+96Wa+IoINWELp3/gL1hKHIxbhfvwj31W4HWNC+QuQ7SJEJjl1xot3/wP
ZVORhVd3exKSEDxNECd9vrpSMrj2Daq5+gYbWKwBwC25jRX9LLseYYkGlqN5Tpb9DbF00XJ/Boba
h6utWN7kBSq98jQIKZT7U5imZ/xzY7bXAM9zwRa26wQ1YJJ74W1AN6CqkO3KupJekuDY++7ZgY0z
ZE/0Yxz94nWclHIt1j84m0OuzAkk8UJ70hEmV/XQzs+Bdgi3lcshUFfZDMJ4mC1dpyoEgzgfGOku
YKd4TOQUaHIryl11BTfmWK7kPwtgLyMpwx+oxgAuKgQ5n+VdnRSDjK1wTo9UX9VjKzKaLkCpkYBz
1Bgl1ykDpHAyenpCfT6w8dUnzc4iRf9xRSCf5DkTCKhlfIRrg/4XHVjhjrZKdOE6w/N4cfY2kruf
u2VVlw+JLWxxG0V1bFeBUfFY1qmbcL+iqZigfVMLMIvZkGHEl1Vjc8XnGN+I6LFEKkMFGMNDip81
XkAuTChMlqdHFHNXD2UsoQe+jA0g0gwqCTJ0WHrETrQq90zSHARf4LRgL1D+qQdLOBh3Y1p2uvCa
jFgjF2LQXr5ib3Xgt9qrSmEA1jrMKzl5VXyhYJyK9gtNZfHLkNFrUAKor3n99efmNur5ArWdfx8r
H6+aHbEbt2ALnsJRo3Xrv6rV77wAmgTIlLjYlPiELmFhb2wyPxlvnIrC/XHg8C1C9vC39GY0OSbd
N5mDawp/Pytfo6SMZLNwtzhstWJ2e9EPw4/d7GcAT7i3rBwAspjbNLesXiTBtIVSUPaD46xxMoO9
JmMs/1j8L1ubEuzh3MeasB0PQKIgmIuS6f/bTPkxtAIVAAP9hz6WKL7xBmaMGnInfYj8lQGGrBl2
sjLgn8CSzhn1zPQ3anVKYRiegjACwYFxwPEgI6susOKq6oiC7+uLCwimggC5D9TOeYZ23vtJYzOU
n0kGTrawMfpd28F75SPk85qmIq6jGe+TB3C8PolXS0V13fl3RB9sutKoJ//CO3bOLKkpK798/yfg
59MwDwvXfCPjypm/kawXFrE88XtVMvtUVCeRKWsDZ2fMg6+9w2nUc5V2Ubnpd0ojmNJE+NNwbghG
L5jpFxRfglQB2pqDxckuY31rwFqZD9pd8Aek1jhrqcdUmYVFA+SfeKHc+8McnWLZTY4CvLtpKWcw
VhYhd2QkfwxpSMIQCJdfaEG55qMObYW5qsRQU19k4Gbj6NNxlHvho2d+j+AG8+in1DMDHBxizhWy
SxIiB9gCteIKxltLrRvZsE1Hj2o2lYYtDVadot3qS/NNHzQuUIgZ3c9wqyv/Fh2XJ2j7zDCZdr9w
w1FplGpAlDjoB55lfPN9kzOoFJ1p6zhiXPN4e/7VV6FHCQ2HFBMK7Fs1kbXAbkqJ4O5QsJLQTure
iQH8fJYeI78qdXEFbeMYNBm9cq9tAoLSyKy7OMqOCgENh4I7loBwHztUUWJzEcvXWWWHlSUUZBOF
IeEljJsiykD54ZQSwKgltfht3uxgsc5S3OtfktkZ9DcmoTIcwikO5oRf2VZhltzcJFi/etjuy6Rx
lcAa7P28zFJwpTPv6XgopzMp9WdopbMZtsyUiQfOH7ZlH/XRtfnFyxfbxb9mwwR0elVzVTRnyHp3
YOzU6Sr1UoW1RJJb6KkL6W2PrpNWyQ51Kx+XaI6GfRQQyuzpXwlC3fg0+L32aNGBoWRStSJ4YHqr
fpWTts/+2t49JJpPviD72WygPy50A2Hby/5GZoQ6y3pe3hhp7nSNldWrT3HonJKlrBWN26mlsWrD
NJbwseuhv8zApJuTb7BxG8aYSGYrWK8tunN63+6FutUwP8/Qvu5ZX+zKnpfYH+LA72vlrPP8LBCR
EmkzAXaY2jruzMJBsF7IHvl4K5SPa94xHkzZv/oorMj3CiQo1etEU+wUh4BiLayq91sw+LYGTj7j
gw8nwwIlu8aee1UUPba0O5PYIywSgiAKkyCLop88gKzgrR7fxTxnFrlIeYMU0HuWvDcwlanueY3r
KYDeEBEX0FbZ38A4hjg8bDzuOGZ5n4tj7DqL5d3HbATPMum/F9dpXwZ5sEGn1j5UglocwYYaiQTq
JAlQ3buxfrhIAJj4jLkzVOKHHulodcsor8susGB5x+dsfSuoeZbF/r9z24HxaN7jnv9OrXyIi4qA
fVcDaL41AKVhKryQUCYUHEA3gy9W2xglyYq7BNVowO+gytIb5uPJxSXDufhsKzxKcXfp+10DpgsI
1Deqy7JGyHN4JpNYnDIuMEc7HsL+uX6EP6tR+uJcZavMyWu2n7eUc3sOR5IDeJsWlX0MJYGTDHfh
TGHqBhH5OME/C4tIQPMOdOaE2jBh6BeeNDSLsbRyxv5gBeoeHlWwdReBTyp+JhekqJGoU2oZmsWb
Jd7npvve7M9/aFCkDKzKI06UfmkgLkzQI5zCgv2e0TyvWKAOnEZcfeeFugpHS7COphbNBh4p6Q1j
/VcKJv3mxBhtv8GXv7Vze7pjTy+vu7D1QMN2LmIBK4oBnIYypDzpc5vs8g+VSO4AWnh1qYUHj1Bo
anZVuJFNxKYR47A0/1SMGwvmOfN0Zan/pxloIFCKVdJop5LK4M1u1K5D4mfbEAa3qZgfYK2OUi80
T/tZ2Eay5RW2ifgjKA4YGwBsu5+ygyB+sSn3yjRAj40yBi//m+7pVFbMU0X1zxtyNTMhdzMUjvIe
qM4FTVsCbGR+FVZOwCt8NdyxchKqTa4dIwgrKWvrOcYxnZmCISDplFIh5LdaA7MB4OkocjlaMGte
3xBilBxARQu566oEM49rl6pQQHE06Aw9gygR2aIw2jN472SFi/GDKsc1JqnGybG0At8g+EJW4Tkq
5IzSdLEpO4JM9txDt8UXsvcFvmIaAwaO1eJZe/Nfg9YHsQfLXRKRsXYdjtsJwmgTRB5OET85OfcI
2vnWgcntGipHq7pXLbRVP/EPIi9lTIqustNPatdMf/FvOidA91B8GUHmIV0YlzSFWCKIQ68oUhQD
lhRslxtSz7M26l2L1/Gv2D679CPbfSW/HXpFwnGgNEwtrP9V54pwU5lvDrWh1eLjmVkjts2p4IU6
gG1wVY1alSWE1JhDCEZZMtfvA6BrWKbwyNHpFzV11Lgc9HWSzCjow7qA2osfOznpWo9jE8/4Vx3o
oYwqI4b79H/GTFy1iUPCtP3IB60BkwLsqS2fPmCJalkRcoPLL8YwRQLr8Sd10snD0qtRJph3FQvf
UbWRSF/4pPMyulmrxGnLJ2x8ILX5NXD7tXnt7ylH/ZsW5vShXpcS68OHtktj2gAsdDcOMkMVBEJM
SsxXj8hraeiO3EuIwCVJs+Mffxv1V5TPEclP+rVdPRqseDFFRpWV/9NpT4t+TVa1YTlrdiE2+/A+
sV77/OTq7ielpr7lEHzSZxKJvi0tXgXqOcII6c6S4HiRL2zx6q+QK+YSQRtffO+E1+Va7/VedreR
AQNXWGhWupouvCYF/Uh9/tSEXlPUqHHN1ne1u75MNnvrurXFSV034OxG/NadB5/+DK1tMEO985R0
gA/GBe3FYMyTQvZ42S8iIjfLx2r3XD6ixc/pqE+FrMMx3B/LZRxlocvuMoJlPMoGKzxLoCANO0ue
AcgZXSbe7KlGShbwJxKXpmKocs4fc7zQfTEtz/vka6LUnRvD9M7jU/xb1Ij21ykYX7BqMHF3EBYQ
BiloRhePwKfV/f3R3sYIPycoXN7iRkT9zlOABF2P3gIQ/ikA13Poq4kXs9J2b6MRMj9FkTrnORO6
Nl1og/HlPc6CqKpLUUvY1AQ1Oo8fVufQ/Uo8Yjig8IJYUsaaTuNpI8Hc4fsqnfrEK5jm8+I098N7
vQ0elpIdmsuaNtENSghlCA7YzQi586orSM1dj2imlV7hsXnN0qfpK05ht0Jz+HFdMD4T5cL9uL1Q
yANLAIAtwA969mhitUxv1aLMeUnm5D9JY2I8ADrMWiwkhjld0z0UAlxTy8miJS7YWGlWZMRgr0HA
glu/gLI/vKrIFXstIBIe/QpkUDZ01BjpxlBjazGKhJoXFtBUGQDaAxTJJ5gNYT+9xcehR7EH2g/9
YfU3yGV5MXj270XfDG6ymyN7/w6gc5C3mObSn3seZh72wLt2yJIZJzDgE9veGQYaXcrxL6tceeDI
4kqxe3YBu1vU2LcWCDoe9K1pr5VULprVRiBsMGH+AbuCpi14qCJEOtK8eNBw+RFPegYjaCL7B68M
GppsTZ11o70hD2zy/gQzgmV/rezr0Vw94Y05EhsV8mi6Mi9nUVrsdhmpDKRgGstOqES7xY+rsd0F
dCgw1Jx3JHHftn8XckagLEoDkJHCXQ8Z0zJx65pioWkPsgo8yZOKX6VbqNizDmP2UHFBFv6AO0JG
6BRMbqHwuQBAaiI7mJrML9suuuBqVwpz4FmlDz+8Me6DQxE51Oy+nZZ1jdlEP6VjdzgBOLas9ouw
SBBIqWq6QLS5DDay75vPrZokvN1fEli9/W5QwSxn5d2j+xT+mtKn7C6/mvXi6/dIjz6BCuh1uwwS
IwTGhFfUgO3V9WeiuXxRiUYFZI6LezPGYPR9HdmltxNCzxA+IXke++sTHsGYDWDHyPdzXFq8TNxR
S3BAWa2CC1Rvm/gzt8wivaRAOSTJbIVp6Utv8nxFx/jIfrT1c0tV5uDmviV58dqFw7qVR7Hhf90U
yRJBM52FqStrFpC7q/PM9xyOCxi5ME5Sf7NZQzqhiLubIExuJ8w3lARznObWBm+EHTdSY4THcv7z
oC1Q+IYWVY3pvHQGXDMDc/e0I7QRALK67knXcQd9Mb6lEamfLKKbCT2fmj1r/NkmrIU7Ho6NADoe
t0sTS7zNK1nT95wprmP8mm0UuSUmbt5rZOGDqNy4uGqSs9nJUV64Gm2nzibJuFAkO9o680keUKwW
AOo/jjlMHBomDghh/Zi2Q1b+JM/BNt6EviRIexbc0Ok9vA96RKa6cFZoyzx+s4w6EayCxbxIrRq9
p4taXBVqAP3gCB/t/CLbRbuBbtv5vS/IhHL1e8VANkuGygxDnGSnJaRFQnsjwMAYm3OOSJ+zprSv
CzLU5v5FR/QmfTna+wCunMf8cY1S/B9PJ4sm1YI+a8+C2mg/Vv6QOoFsQAnFj5hblibfBK6Gth+s
eSP17mU7T+dod3iifemCU0MsvPZBQECbzDWhgCNm4lmTvAJsXMJRq4F6jnyNveqXiXY9O57xUWs4
Z10Jhb/4j9vzhrNnokF8HbQR5iX1+yo7vsVfM8HAEvcouBR0vxS1/ZQt08fE8ritk9ta6NgsEtKa
eN9zBxW12DcAFyTS2xMlnQdIsTsirDn1YMJYB6CQkGBOQdGZE946DbKRyGkTZvXOxEfk4hLdAMJz
gf3skmEwuQVHEpGkBgxId+0EC/AVHObLIw9wBFJSJ4m3EpmfCsPeK1rtLfdwf7oPnUDy1yuLbc/p
N2yo5bfjK51ShUXSaKWrWCXplVvdr7weAfbponM5LBKompRYM3DGPs1DMkg/hJbh/sHr9lUzJMsk
HBFpkCiFnbRv1ICvFSIIJ0O28N9/GNpEww4Q8xrsChsRJWa7Ca0whFgOvb613VIVO+e4xmAergop
GOP3o1Rlw7QDhrGI42A8N5ZFi4Y2W9omqt6vONc7bP1ZPJXW97E6YZRLSij6Pp9OW4ymSFkaJycY
kVQm1AEFuHdrtI9O9eEz2YtS5O8rAglR8PJP355JCyRTrjE35dnjV86rVGU44Zr0deDQBGTIwk7s
32Wc22m40NBZHcs2bMkJSpehhIov9m7SCwILIr9M0OwUuHEix/jGujyISYGHCbKxItZWr2KkYqS8
21WEDDUNC0X0TGXRT6hhqtrClmhxnV92h+FABpT1fLQGjrp1cZLn7KFijd/LL9Kt5B5WCRsdAkpF
Y3ynD/YOjBds0tNkDbXZylWEuWx5UyhJSAw53y5gnJJIaF49Nv1Y4ahAnObZRhgGJWCL6/ZgQiMh
f59R5wImRxsAFnm32UEsInhq+e/jno0aXCY43/tbWYK8GmleNUPAOxMFTzY88Uepg97T3NZ0VsQ7
I38tqLjPYHNQFByUCKteLsioteNlWY55+f9m+EuIkEEraJ3BPHKw6GbV7sIP/OjdbrXdgpesGEYR
7C/K/0vCi5yiegbqDLNn3n4Tql/eWKGKK2HNbOGGj7+kbEFt5QWHzHm44Zj8GlCksdCnhUMR8FN0
i6BkY1vBjoHR0Nz4eBdOKp1VQNtrP8H9B/vTTbZhabJTRxgWFNiCFpEH7v5K7kzugGUnANE/Rva7
wZ3VOo2+gnGRT7aZCeGdY79DYYwRTjdB9I0T6jcAg3R6fKWoC4+WABmRdm43RC8BduHATJ4j08yo
Nwsk6EU6OQMrxS7NIplLL1/UN0INTty544m1iumj5HG/dH59XwOfgK+ijwfP4HWL7KjstLNH+2Lx
bNP4PBSv0glbesMgNGWh8tmLqmthFDI0Kq/HAJ9tEj0oam+jNQHyWd5WjQJbBSHqp/vHkXXAa+1c
ToAS5iJBv6wXK/8tiT0Hfm5bWt7D4vlO5rgoq6ImOE8utZKM70v4k0B2XvpyhKUkuO/PWtjogl2+
YT70E5GD7gdc8LogNeHlltIFSP2OofNvcdO3oejLunXqBTRC6BdKtOEO4OuIj9E9dtG8OhaUDVUx
9Fu/OkpwpCCw7VQ8GQN1zQD0AgewevoU+HKnoCeHmxfUtUaqsK7FKCGw+ndyel6JCBoXvS9XqaHB
RPrguI7ig0mn356AoA4QH7i36OSXVQ+RsUZ5lrAGdAWlHy179vhMKaLsrDJj9mWOjA18Y1ufrsOZ
u15WRo36rrp55fIUWAlYSICKrsYFPybJxpPbKqAJxlWE6ZFHgeqEQv2Yr48YyTEl+7L4Ho6lbT4k
gXhWTr8/J23ZftzyyIAjj24BtrMIM3acNMu+asnwUmCWykdsPm3AFcK87Iqz9mz7j3bNeDAuM1cG
Nr1BbWG71Ir0sTx9HqJzaD+ARhDnRTPDRODCkWR9yjJucLaK5FAgwS5bhmiuhkW8Dv3t0iSteCPo
GFkYdWjAoM3UuFKhl6oOp7NAOn8UPGbmbK4iD4GczATnxuvST1md6KRIKZMSGRc6Hj/Jh/VCp6FZ
MXz0Z5CxisR6+QOuSEadvy8qT6l5iMfut3AXU4F3dFx/MpRb3nSYkwP1XuiYrH6gFkLilsLLhHfQ
6NQZNBSZKMIh4vKPcyeUuAugo1GqDd91Om0IElGOj3C7PsAmVYEar8TkU2znmHxM8jcQqSBUPxwn
mdX7emvn5XSliMdYUnCiQ3M+3DnAgLkH0DuZlZ3xzTGJpKOYSz26RnW6/h/xw1i/ysc6Fwm8UbtY
8eoJigfZwB80YyDK/pTU2rmsMrC8vGuX42NirxZM1ts3++bTl7RSgUob64bVUM++6SoOkfKJEUnz
jvJFHsJpQK3izpak34cweNPv7FNMBgutKEpc0f6qtxrNxSgz35TbPS0kXzJn/D54WLN/rqevq4iu
PM/ZXx9NfXQqn/OzaB0j6tXwLmCZhAkoPxQj1G+x+ZIpWsSfSCbIMlHf7G8Z9hGqy2r2OgBs6gbX
iWbpdbovKlJLYeMpYFcdHMxnNQdyTDCnTlBaBjTWLF9bo7vq5800GgzLUXQOPR567DuIUJWyaQ9F
Pu73+/yXi5AosNpxZWa4SB5OhgisvX398tPmz+j3DBI0YzQIIPdhahOqePSuCOr+Hfb+RxWRDG9C
Yo6RGIYgSd0/PfhFrN6yk4vhMeqgMpfx/uaBcGQ8GFeHCZlM9iRloN2K04jdlxEdUSiloUYkdGrH
NZJQpdDXet7WN4ClAgjpk2Z+jbtzOiEktXln2nWdrf+FHA+fejBxIBjRR4uYkzZXN/rE3VOGzeb9
KIsiAGLXKU9Cf+Fd/rJmk6i9LS/KAgjtCakxhkyAYj3i8wckpeMVBCILwdknWjaf0RoC5GVkQFdK
8RnNdA0hAkVaEiposq3bK9JxpW/jXLgF4kFbcXchCgMbNcZBlZDSsEZDSrb7lWFkrcGKPqUsmVRg
8n+kX71SGEo93dVf0IRfon3u9wRKCpJnVeChOv0zGJm996BYRxnqSD7DBFyxiXUrnDD0rfFumgZR
a5WkUZ6n3LA0kbMwztYKs68gFVvJx0cYnYC2n2rjK0ApEL+czM4SldKhf3kUp5nFO3WnsGMWhKNf
YBaDZQCWFfjZwC2ZRvjKh9jvWe85S7Z3sKBP0mYh8MSMbrVqJTrIhFhdSyJrUJN4pN+aWyd20X04
iIOjpiJuuS7jrfCv422qC/anYkEylMgenAYt2GLJ3542igW+EFPb+F+fu4MsPEe/L9rAJMiIGkdw
ifEjyGJ+XOXczQVweO2lobq+Cy7ApujDKgFq3czAR2kqUjFQplAnH9ydSfI1HS1q3nQCyOwNsoHl
mcu89d/gNc2uaZy22y8QbdCx6TTyfzxhXEAkrdbwu/Yn8UzX2qg8XqNFew1brrnlWDinSOigveqg
2sw00eCok2ZDzDsgrgZVpusJ4wSShTsDlir0hckWVu6z02Q6v9AOfORrIbzDPbo14UztLCtK707u
GOHsxNQW7RTiRpfY/MMWI1yeqFUm73zaS+B5u1B1mzWk64uQm+/h2Mcte6Ex96ATRiajpn+96Xgl
fyZ69CFEHpx7Tx4DuudeadkqbxKRtMP8YejnBcNJ4umvQHfnUgUncL38Jjo5ZBBcEHhYwr1GqK1E
Q54RBEVQqnpMLrQX9Jgb0Trr7JKHNQVy9PtXwqeZ924LMx7AGlKeaj88Fsl3+nn37dIq7UrJnLQp
Pu9NFtfXTVCm7kuRAksAufsyurwuT+/RKpmKFRGMVo5gc8yktBPyJHwZP/nd738a2oc1oDPaW3tZ
blEohnfCgRlXQetjDDetiMAAufmo8H3xf8INeE1vs14kkUDtX26uYyTGJDHsEi6kkAuKJbecdpjx
WCc1fGaRHSwhBRjNIQzM72SJ5+cZ9mHyIBgAdXE3lXTRqoEPrLq3YAuAHuMUgzqXI+BlGc54LJ37
Y+p72zHAY5wO+qVHK2i/frZb3txytsK4/Lftym7MHwfXuXFUgYA4xaIK+6/cMXomIR94f+eXL6nm
gVMqRee5newo47rxqh2RP0aeVgppkgGR/TCnFD5A3YVIMxhjN6bx+9Xvjg/RPVeZ2HqK72TsirYP
9BAmP03bDAxpad71GI5sh6hDZOtC8I2pJ1nNfAlyoXHbRj9F+A2NVClVH3WLY24H0CVw9VHroRBr
+1Xk3WlM5/tSxSr1xlhIk5PVdE1n+zog1X6wKxFrzW7wXiqD9iHyWBDdtLFGjn5aOqlZcHeHZVxR
aFiXOSruv0dO0FaX9ftjQbKE3uXYEVQktB2MoBc75ToV3hJbwavK9ZOXl8PwKy1nVEC9UcDS2+wd
jcGL5W7fxqrrByFouJ4Dr4CfS9haTi/kjhv4R/jpw/8oiqguGYIdkQAexCnHE+lygI/Eq0z/thn8
+kLmZ33JTIF9VovZgDZtxxPYzo2uv9zZW2vagOVAUNf8JRv6tsSJnClt+lACyh/EqA7HkhIQDrfz
uTsCRZaCmwFi0uXtB3e4NXkl4AiKomAEV8Fm1EtV+7k2Et6YAwIdorGQOfMF68CWxz6Q/6kFoGym
99Ipykwe7Gv4keQIFu7/rjlh8hSDxTiNbM8CFyHiOYauX9QGK3EzPu2UCD1VZ0iLIQrxh2wm0Lng
yz+hlq7v6hQc9fRXIwyPIKdZVkAYfM3qc5Qw6he0RLU9aoe/lj44HZtE4r7kzFsLOX41oO/2Du5V
MTsbMsVYJKJZE6ccVXudrHHAxNQUE0YMYz4SpulD1kDjMXjjUIxqgcCyi9+NRcPa8LitGv+IKo+E
BiscOIkD1Yf0iT+54uVgjSYL3a3KyPp5b+fDa4s8IkCCpg8ommJKNjrfX5G+HE6r89s+yV95W7FK
jhfeso6TDkmcJ6K119BLT2iA/ZdGtXKEAEXupn5gZHcIZXdpBwXhWVBdyjLcxioDXh36CuhqroH4
ibYoqh2JHCr09QxdDF3ime+IS0fG1ezKBaxI3eZSxsDbxhH7n0C9UOKAoIAl7afTpw2NSMDii03C
nbltmA7bQO2HOJjXKomrTcJS0htfAr1qShZXNeoT+3cDjozM7XatAM2jLUg14Pkvf5e8TS37NUAS
pvgmgZ6EUszaqL5IWJ+mm5rAEDgA3H7HMLDLz/ZB8EZY5gD6QxY6sbCa1CuYB4ISnGb/ymoCjI0l
ILX6JyPdJbqjTlz8mvrCE1rl5k+HME0C4RA19xZ3U3BmxZdgFS02qWsczhqCGlISxq3jsnamaDFY
fiD+gwX7tW8i3dHYe1KwYKM8OUTup54vmVrrXeJO6flp3eNECRFvY9W5skD5bb8nvBIFnCf79bfK
uOSPSMbqIm2ve6nypshDH8jEUxb7UlWqBtcPxFd4McJMey2cCS31af1VNkndj2OtaYHQNsD+N0RO
Bhl+MAqvzSWLwtLk4EkFQbUsQ0VKYbj8cXbM/YB7fBEasr4u6Vrpg7djGl2zDSzCvD7u31nAfgUE
FAEEYr1X6O0p3Ynkau9uGWomvPhfOyfZMZydx2Q768SUBQoxCQHPfPAF0e11J6ghMWRhag4IEbhc
DYuzr8HlJBO+xymWGUJxWKIwshFj8uhFs+nzX/1C5MYbjQ61AMcgjeHDcwrZXKWaK9wHP+n0vVS7
LS368jw/sz9lRR8dJnXe4XGqogtqtl+FsPL2Ur9/mi+2w5o50qRgeIyu8sK2e6ofeWGec+dv1VDM
USV5121+1AzchjqFUKWLN3wjPdjtajrYoZdgyCpRAuy+lMNfvGCExaLZNhoeZ0zPl1gWD8s6oAfG
ckytjE5jMQ5UGCgB/jPvGRLDL+pPbXcnekqIUs3jethQD5otxPwicUDGkCu+a/ZMn1pmZUpAS2fD
qKFB4Qwm0dkixeBr5HvH7bNkri6kW8tw/BVf2B5OMuegqur92iQ5f74YeT7XIV+5Q5Nv79G+fEAP
IFxZfF7wi+jp/4G7dgG/OYRbQCccO8hzaDXGc17fKB1z/i+Ru7NJG/8l2sGBgYx/u2gobebzOK4f
xfpeqCQWk/G1UlnPaVOe/JmDIZkLiVgZpjen6kTnihMBJGhpcUg2N0/sxZC6eD5u2YWKmPEkioOE
Fkc11KsDodMrVfSz2BKj9MOY1NKJGQTditvJFvog4x2Qe3YcjqKyM281ONl4Pa0eFc1eXPcKxjPM
Y2g5YaYVzcB7wtSnOuUDIvtQ7T3C6Mk1zHASSqRi3DFydh5I9DqrnVZC5GFToAjtc11Fbh/lYeBC
2MJlGerxYCX01g3b6MRPz/arqxFt2jsKfJ9jnpL2yj02ACYNN4hVlpj8DMKKVVBHWPzdHfPZggTt
QRpymCIASTEn+fvZ1B3Vpe4MXDpidQ9QpX5HpgdDuCqGWbFm4rPzkFUcXmUkFDO5zSM6Uq9yv48R
oz8hSkvRwiX0It93PeqqeS3yg6z3HJ9SzEVgdPV8iyat/WLcVM0xPSfIc6HMRFcPW0R30e0pfLmi
xCIpnpwPlyNSmkc+wuQVdhSGJnD2QqHBrvGaQh1VI5C8InPw7570SrQNm8Ckjzz7uhmjz+QP37Ef
+1a95Regut2oAK/UnTGtaIzIuuyGSDI7WvPse/BA49+b0BFZfqq67vr/UIRTyQOi7TFR5dzhascH
/MNh4gcnu0Hfov3ztdPfxTIZSl8TgIRbXzQixcmFXFHaTeJ264a5LzCj5aK0LazvBmbd67Kq38Jz
dclvOqD7PPyRXd6H7n9EwuzsKIwBjQJtIWfnkl1WtD8qiyW9Jb8LLAKMkj/rD7dEk6kbhQx7z4Xb
+/ZtFBhRaFhKQNtwiZvj/iGbIbavTwytUYY5OPdguy7oz+p6SNsTPwFXKmlGUgtlc1SXi/Q0Yl2j
PgopPV1stW3AsU20gaGyEKCARCi2Jofixp4SKmK5GjH6P0sL1wHLC28HtLFo8rQbXdQTPr7RQ0/X
gwCQcXQhEfQileuKnR7bTPTKdCPxAFMj4264jbRl63nrItf6pki51TiwyR0P+5eOFFnPKjGpm0C8
7vvIj6RSTgp8I6lqSemQgdQJQdJpWWGD4uTm19Z1r1pimg2C+Yar9uN81qVCO2HOzsbz+XAb2LZr
V3FxvPB+E+VTuWmuGzET9ElWeg7bpjam+PK+/0qg+BKe/huTaab6jMImeNOwPFZXZDmk1hqFWBmR
V2jo0VzLseYI7UlhivMTr0TNFv/pxGiLc/pA3qDXpdx5/0DyVmHHFr/IVGw3f8E+LDCw1yqsPAm8
frXlLlfVRoKOe42PXCRoI5wyM8lEhyHVKHf3RZXzDNIZFtNJRSsbiP3Oiz/tQmlYFeUURidkkYfN
ctc3J3ppZ5Bn9ohAEbv+GEiW6HjUdifaXoFKyoW/gjAPnzjq+33YI1LE8Kzqm4MBqB+A/79Qfn4s
6UIfJtZieGdzLfCXehou95ISwsLZd/8h8rKrZS0G+q+Ae9kfFGN0AF1lJyOrkbjFp9M/cUvgD8nh
OiY5We/kZd3HQdsuW7ScodBlC9wXFxHL/u0NGbiHIVzjAUj7S9vLxbhKqqrb3UcA8WDcX48O1djb
J5zWfW7FE8w6C8CcSr3xeS+DFtecVaRTbIWeNH9J+RTHdD3h/5oFv+MNHMOgESHxEz7Zvsh8DY9L
dpRTYoBKb2QaeR4hkIxR5312My/KYPyFQ3Bdwf6XwbQkkYl6R3uExxXrPFlD/Q3qZaVfUoBicZnW
788vweSdP1ojeBuL+5JiLLd3N5lRwlzf3VtENV4GF/m2xBNZ9gCFQiJF/DimiYwc/FrvDCqVIoh5
++V7sB/BAYsnt2RsVtIMIWzn1b2Fb6GAk9N/Lc9XHhWgLNhsbkxwqkIrsMp5z8p8g+vJnjaJ6n35
f1oA1cByz4tFCQkNUqwxB8cktmr0d2pyMAB/EuH4Er44F7Xar8jioaHleeUl5ES9No3xr6C5SOaU
YKss46dmxRJgP49DwCFXwgh1AYu9MFKP3xgdart0LRKcpfnZhEoT0TzQYHcJDVfRTftskwNO4Me/
Xvm5wDn1dyFpU5UL2AIHDPX5Whx17MNV3kGQeHyN0y2y9DtMWBS1JXeqBlT1zOnoGgYFaT0xn1pc
ajshjQBf9e9bmABkRqNYiu/kKlEbmSG9mmG32y5BaOeQI4/rlMpQtVaibDSUySQGB+pD49UTaQwK
VjMES87rTOoslhsQe+QWHinSzDaUTTI6wKT61oGik/BnJwV7j0FrOW9msxKsn4pKKhr50k9fMYt5
AsjIKt9Y6rV6lAwMjSVseZJ/er3ju4mUhGzbW6aNt5Dez0qrXmcDlENND0jub5mindnP62jOaTWO
Q9q96hJcn5uac9186Z9HRt7vAbR/dw8DkkJQf7YBNwe69oprVB3joKB5+DGARfVNFcCngabx0Ffi
OCM6TlJt2PkYoiGJ3aCSmeuYN13CnpoWJNf4RRApKyScSmG+2Huf+aoJhwHuQaGI6HtKuYGLLFzX
/OPpZISSrVMMe0DU57KMDvis3b08doqOTm3aJxpPG4E39OR1pT9FB47CCG16nh3wIPXvHfOoWVlc
Gg5K8x4J5Ri9Ng942YrdKA7DfKV679+pFCHptVgB8FtYnTp+vPv+/6ZB4sfGjTqR2RS9vzbNQFBh
6Wa+GxQWnhXVB+dVDt7w8U6DBJRRm4GFfO/Xnn/NIyMFTXN/Ynh+YPeJmNpL8tfnUFgF539/ILYI
OsBulGqPxqOT5i1yTtEQqVLWrzbz1DqTRl5P2c5IQIXbyORYZ9tB0QARYWdieBGe/jI3eVdGMBzy
YtPsmy9nMCndAv/kBB0KdmoaQHTDyCKo6EAumwFrdbkPzLR5zaA2zdS8mohaNfvAnvssctGDJthN
uTKdbTvtBoyb0Hi/oQraYqV7SzFWaQIQ/I4D9VXiRcLQiXtAQpSeK401qr0qBBrWCDToRVY1lQIV
eYgoDbZqVz+AmFjgshHswx62ls18nXMUflAIaq2KdSqvD2II09bFKKw7DwSXw/+17uzbQF8faubD
ccohluGH9d9MXVCCMSla3S6po93aduyOzKr+ERABU5pNm+3ZES79NOvQjo9BazGLjKbLg9cIDnpz
7/ID7VshvmKFr8msKysMKCzDbKCkaejEyBNpt5Dcr3Lc0ySk2OKJPwOholMWCCObPcx3K0LbSLs0
wMtN3JrIWyAc/WoSjEitAGFO2OlHTFEapSxOLRqa+o6nl9SGOwAS1N9tjq/lZfILgezC197OPWKi
C/aSipIuaFZ+5jYzYNJrTBWwFkJl6P+sDCodSd4usiZzInZmuO3RCF5IhVnpzeYzPGVpwfFN+bmq
vBNa+owGLIw2aW5Ry9qHGaOnyq2EkZW+bwCh0Y1eCXsvb27u8xZadt97TaXoRf80xUIOT5SEUhgW
uMNqLXLhPyqoItT47+EIn1Wge7FBmM2UoYYwdUBL5pJq7ZPbJtla3ov1ZHJZoqkPoXZudWba2BeR
urhoO1/z/TFeXrydfQs3wL98+jkACF4bjhoI47WCf/SoRe7dkTKN7FmXsLHrdywZvSBLnlVJop1g
HleioVRYGLzzqBinlBLNpsfj+nRopA3k8QMdRh3FsQQP1D/qpvRMA/kWMjc1aBC8+C1URNPWNuRl
SnkIXRroWByaUsxpLKm+IAcYiEsNNiHfa/tcQynB+az+rAz1dbJZMN3srP4iXKcbXsNTIIfzzIhM
afU32j7U/XxbXKoqRSjYAgksYhgml5NjlFXOMHD18+LJ3uHcz8Qjuz4rstSlFMM/tUSnFtREinu3
plD1jOX8FH08RNyUIu1Zp++0k1HKQmbhd3ybxIIFj8EtBOAWBdx21WCqyLgkO4R4pBQIHTcRHIRG
Fq5rrASarafyXZubMjfBEZ7TUv0R5agEoouCogrSzpkCNGdl3hX8MsDl71eGjW7KGwg+JuxYg5lY
q+Zq1K0tjhpmSxkwe+DMJn2c1QfOEOpun2XJOZOexOtFVg88/GpOpAO0TEMPCY/o3DCKG7+cX0Ii
eRfclBOJisQB7VR+/JmWa5rDRzSxnuLrW5lCb+M/SyOQ9Qd0h95zPdjFxPjU88tbLhJ+ZA+sseX2
8aCzC/VxcSg8YVgCq0GhkJS5VQ0upZI1WxMaD54JL+9Y4ynaKmMDAML0Rd9at9fjFu39xpayN9L5
L0iONib/xahSSvWlDU4L19Yn+eQoFd77qQL/w8l1dCRtjXcDMQWQO/HBtOLEytz7cvCrTz0en4Xv
LMBCNX5wKRfs3uMhIN73dVIKR8TdC/VBYCZ+7FYfB9E0cMZb6RayoHWWkIyrGrK8o8cokgqDAQ3s
LiFTL6jTX1kHghAl7rRf+rD8F48IqEgxNE3PFhoT0/79gVxJGoZ8Ev9qhWhldCT3rLcB0DQv2fkI
P47MWzmUrhhqsduR/YEiJpSGv6zEE6avBZoSm/J5lnCp5i9OY4VSRDmgoN2iZ/ar8y8CjbX8QotP
CbLYY95qzU4A14C3/uEUC181YdwF5qWOecx7wdLNQqmRijACWVk/Aq+aNkOShfaE7DCuaOhgKJUR
WUzvRB7EIZgf3T8zXzsWCegAqHJay3ySl7/VIsQrQ2gA3lQi8ti2QY3KXc0r+ovvCtUT36lXzSyS
nN3rv7czkw8Jag/Ffc3ksha5XyNNY2e4qUu7p1adZoMV346lzRhnCLnSpMAHzseorcswPsHH97S6
uYPyr02Gw70c0xW+P5Fms74p8/mzu2ebVqUpnGlFNq+H/+EPTxiIhvolHIcyUZWakx4AFVfigyyp
0Dt4MJBwVqfNDvEtDTs4JXoq/73s9COi4s1g/8YAVX9wxCHPED15EMmqG5L5KbGLgeI68kJk50Bb
WQFCXUEU9mRymwADxStJzFtg0NwvCtuBfJxvCCT2QtY+xdRJplGIC9aS2XP+oXljFA03VzpTouib
cTxaWuVRbOwUC5xbe37Bj5vSw7kqHWrR6yJ5fhg3Mw+WEDycJov4uJj4SjEMSK978xzKjKfQVv9n
eZmm5Wpkvex4RV2cQ/4Ir90HJCR6tb1nW4miCtllQ3exTIK1Mqylk8Xq1/TG0WqfF6FOozL8jJsB
p/3a/QatRqgzVXVTrWw1suHDSdyzUyM0+AC0EGRRBNgHAPF6cYK+6Lt9KWuuFH7I5HclKogRKROH
oxAWtBzjdojPx3WDoj2HOePe+r8/Vmy34Sy1rfgyE/p5XO9FYx2OP2lqIXPLG5KfkyTpA4N9dVvA
bWPohXScidF0OmUUiWCwcguEc+wiFXc+3BB/245am3YhaRiCQ7m6eJVmghy4JaVehD3EH0Wz7xlX
QvnHpYBjHx+v8m2hsNACzVjK9LgLWAIRdMaLlXXLb9bqGf4O+32cg5UyblT3UxpiE1mpRX58b+82
as8xpGe0llw4VcJWaA4/XMAY6Np7qaNzZuNMpS/6gQ6PCOYp2DKvlKTMT7rGgnGt7f91eUMqFIvI
tG5tCkH/fERdVJf8xHblzUj9n+t6DN3kAdg4aU0L8LiSPOUWo/OO5IYDa3kQUhr551QZRQlOAlla
nGyxqg2xDdj4DrkuKbBteO+uIDCJXq/Mc1Hwm6s056UFu8ApNQN3Tt2ueE5wCgdXbWmu1nfr1NcX
QWYxPsyhs1bmyikVurZ1UY75qOH2tBr3/52ALu9rK/1+XbyAY8eAKXgIgk6xcYcvMUtYIpUCaUJ0
yHxNTecic9RXuilnbNLFS3K820jLk/vtkZd1ZUgk5wWDSwTJnJr6Hbzk6EzO/vy7mhgB4YGh57yY
ly2TxZI0xcrOPC/vTggXD0TXWrE909CkdDjz7ya5b8Vm49VlfmMfsl01tP4WLIHQIjQqeDUFpu/b
oV3D2829HaFuwGdsxXkDEaic5htKUJOKVyl8pIw5fRqeNHqA801StJfPy73GLEFnICL9/8TVvZp/
TOELIlkWUgCYbgxZIrvUGEwJqwbEOe8lyszv+1mOvYNl7p9kjmntS7cOugKV4akbxiYGOTMfCAut
AvCCEa/Vcj6U/1cQEiIkmI7UJCe1tmDAiHz5sS6jbg8rJTsuk/+cDWsPIXIYJv09OTgZfHjF7DH0
HuTa991jVfoOFsq3HR4McCY3pZrfN9Y+YftRUlQ/MF5sy7PgPPzdGyNlT9cmCGI6qF1ee6lJh5Nw
c0UZZWn7Jtjbed5ShTTwy+ojdhREVbtQczz7K2svLDBBgabHj0tpt62dr9cvkr8yoxAlRMDy1lKQ
VsbmgY3urPoW3oj69FL3usXF/VHsA/k1sTlgBwyFpGFp4WA8X/chVI+CJextok8aRR3fNqwLSBI6
hax5ZNqD+FHdU9QQiuJ6+RfhMCMQDXc6Q6T8JXeg8sxxFCl5Z4Wbg9JUeW8b50uzZK8OkRMcsz9v
tw5pi+5DgFARRAXDS4QIxgl87uu7i8pCTGpeNNLaSgsOhdB96U3+b97gW5vKjyjw3i/XLiRftLrg
s9NsbFCkl570m/554kpCxFJHFdPH2PhMP3Gy7Vgz3EzW0etWldOKEYCsd7uBaTfDdg7DwY01gF1b
eV7dadZmeAgl/5iXSJcqfIyXkMjl2AuFyYOcvccRA2jfulWBAo7hl7NG8akNQzK5q8BqLanyRZkD
xRpUOxGiz0kVuV0OSUFwnUDMkCwYDMPdPB6NrXev9m8Oqjrod/IC3eSt1AXgu2CkZClOyENULy1G
e4812Qyk+HbAdieJf4HvsbpaiA//EeuRwqN6P29J8TNe5/NvePK7wzjS+0lhihZQDmBq2W0XBvbF
K2eDGSCEF/gkzoBanmmgJnZZe3v1AXDKwWpecax3J1Aj4nAKuRsx1ECEmWpmShTiM9qJzCcL6GcC
wD2Nivr2LHsgySjRBwbzEJ2qctrr2GOE9B4Lo4m+VmK65ddlSWCpgEymBKghSMVgFX2lp0WFW6Z3
ks96AEeDbRuKjK65vbZ6v6BQAtqCW/l5BYmPxNGUt804XOdjhtoMDPuxBHi5FejPrIXfIEfsjbUA
kjSRbwEL8bT5BNTgVrm1GjvIiDTLlMXm+2prpaPqILctPHgwsVAls+z5VRQShPxAuchUKSboZ0SC
bzKrVu3TJi2bYmxdxpNK7lpUkH2WPUbGsguXbaSef+PS2sY89IRAE2e0YhdH6tnynx9MCSLPtCbR
mxoOnHEhraoZq/htTvXGjRSRaScIG5rFyhQ+HeytcL+nNu8hvaFbf8K/YzF1fiGl8lnx6JaknTTl
z159o0kZ3H6F3xtp1IiMuUt318PsxqBCx9HitxyzeVVA0t79/VoMxS0ShJjCYNO858Vj3zQp4f53
zIovGXtDtsTFNYB14ghgwQq2vMiO8xbmVida4Y3kbNeu5eXNUNyfqpE/aLsvai2U8NRZjMIXcXXN
+T0NYIiG3pz+RowQe8vgAcOJQpw+3j6g68W5NRqnrwla2aqPxqi971lGkE2jKtMGia15+yOmEpZC
/oSN4jcRioakIMScRWYrHrQvPSgkrsXaZOElS06a2zykEY59G2hTe+OUHpQtYXeaZdGZuedsZK0W
tWJ1dkFRlJm4v+8kPrpFVYh0AXT+kbSm1ZJmjvYttnLRm3x1Nvg1L3+8e5e+006iBiudka9oPTEw
QFxvb3ix/nc/weLgmb7qE2LEiN4z26PugXBfV9DSodcyc/i8rt3DsqdDzBVvtsxFvh/UjNqRXsta
LMX6iCxT/SpLTPNrciilnbWZp4EBx+LatpeHW4AlMOjVbVGQol1SahbbTO36TULl4PlMOyFP4dkY
7dSvgPOPTtF5BG6BB/SPVitgGjsVgFyD5677/xEmBzKLZ81x2uvaAkFXzO0EP0gOQJI2Swu+tBNT
qSYEBki06O5rl2FlwnUy0ezz8Y05uBALXu6fejGf/abATZ7/hzHwA6ZQbHexmY1QCvQYVS3vUVL0
VTZ8hHA3YiyjXEMrahK8faofoXFl8DhGkYT+/BNLX0sNinyTozcZ1ZbNjnAn3xvgQM2reH+pJ7Sc
1Yf4kfkNIUZF5B1aKTIAZfX1KIo1Vnect7VCPqwuwktdiL9r1aB4Zpxl4FCAkoBruWNfUga09g/1
36mvOmzyq4yOIm7jaHdD8QYnyiFpKd2HqyQJ3r8vtw5NmuGk1/kGq980Z7tzg22uRf1N2OhQ8gLy
Dsh2nvHpW5MGg4QHJph3xtoGBuyNPASQDQYVLU+/zWr4JnQ6XEGavIpVB9DcB8yAsjJtxVFdWyap
0/HIuHMVTMbuQR7SFRlZ+h/ZWi2XwYefTeIj/DEszdOJ0MPrFsvusTJSVjX7NI6Jxqt/NYQYjuTj
BWIchqhelx/7/dF2s9YRTg2K10VKl6EHmUYT4EaTdskFrdTmWkIUZwc61E33zfwiZYqVvvyVxkUK
gM2qJwCCVu77F6QSXLGf1ghUl0gkIkdqy4i1VCklWqaNaMgc+JnzSEryhBYaJNFsl+i5I3on0pcw
UxMvI/gsp8VwWtGJOA27EAoqG+xELJ5YjmMbiZ8AmKcnKoxppxcElry7v4BJOOXOVDdI3OdWdQDV
16LRpi6NjN4xPiYW4j4WWTfqMPgfIBdi2qL0DkLT5/knNujmGS8kvQ+8c/yBz82z8CnfmPGu3Wg9
aAnPj5Hnv0S2H1r1Vos1vA1wQXg9Ne6ELBYmoBE4mgc/25KHZJuD/3ptwb1XYQ/o8JdRXC/ZuJJK
XJf1++DdLvf8UCleZEQVgT31JtTZ+MTMZaVf22+b5R4+xpHnBNktoy/ux9Jignt3ZiCp+7xX19rh
FptQkxoqklF4P3a2Gac2jydN1oEPTWEq7JSO0yKOzavdFbydSpZMW1MVdtks16it06tPgPWBSq2f
4LFNgpGxRLy7hUapEce8kRZ9b8UJty/8vC3OyxzKYyu00BooEGYnKa1MkkkeDRD2RztHQbX0zcKj
OknlnIkOkQjTpJG4FoFxjIxjS+v1en8KgE4b6XufCnbTvrX6tJQbTMETh51a+7Gaa82EjnUOvTfT
27/vHq//w3W38x99fkR6rdemiF2gNHor9SMEIDYLH1gWr7KGhL40hP/DPIyLbi0d3S6KsXkwul7l
iCVkjSRJd2cLzm4O6Bxmrr6VA4u75SqQwX7S9Hhb9xHYvEqJtwb6uQDUafuWClDD3+hto4hCFCqG
aC7xUKsF7oqX6EUJF6fENgbXmj/leTKPAsnn1uz/UlvH4RnZzlGQhS6XaYyQWOjQkVFEEEipb6Ia
QbPoC/HNdK/R+Rkhc/JxKArK0OWXS3Fm6ullT1U2Y6f1J5RJ+Z9gc/noyZY9owqnvvQIg7T5j7Ec
xj7UNyo6H4aspv/EyWu2Aoja7D5QuN9/UA5jCYThGU1tndoRbtfjLXfpRGLjMf0MvWTamYhYa7mY
UyMXmvgCorKyO40zToeyXA2SRPlJMdw7D1b8YuG3c97Hb+Xd1/VjbXyL+EgNLcZs+QNuBlS3FNVi
eUTy9KE5E0auntnbzQ3UHvFLTnIJ6Yu09AanvBu6+LNAnQSvk+4uYsMorzUkmmFefPorhlBitK8f
omQvBab5Axb97oP1U8WG6vqABIp2mvuUXQwOp2ZS0odg5ZmnOX3M/AudjgyobYyorP1NN0LiRHzw
laEyLDLAO1eHs5gO9FU83Zg8+1lg2eBCP5sHNVP6VgAtYtHm+3EZeVfA3Xt868abRwD4SYffXK+6
gV4jelxVNVAY8XfV8hyK+lZTl9ziLWGa+UItKsbXjK9IsZYa1L4N57KfJTt1r/6HQF0g2mAvJR71
i8SA20IvFopYc+EhJAJQW9Rjxu7Eo+AGms/DXYLMb6ZmFU7FugqYl1jAHCOR39N/1RtZtT/UHUaD
R+n4G4wogXZi+66GyqAYIDLxc4arNBic9Cp5wjM+AXrjAmcx4GSRm9NtVSvwcO5DQkfGryMg7dR0
1M1wXGv/aKlVuBwFzXzl7pt38tPIswZE2EGk9wKJ88XwekpffXAF+UoUVJSw8RoEvUI9TOqH3t/T
MT3b7kgcTwvmK5LGym/sTvE1rZ8wQDKlkgSS519DlONq9kDvYnVpkzA8wXfNEnYgCtzKIinpD2LL
VG5t/GyQmEJk3Ykm+p3RMniYhbZWw+5LRa62tsINhyBeOo+HSuoY0kMQ4ai1u51QFSRF9jiixnMt
MXfC6hfn7BLwPxFTOD1RsbtCXwSCGIkzzTbgKJl4YkRcVKH76gL9THWgDIl77gPGslHkoO3ATtYg
Wee0dy6kMLKtQiJrjlhlespZmN9oJoSOTPeDzPmodTiGJBqdssMZ+t+oiotTVCLlauqmbKKfxCO/
hSFr1ldmVbzbWR2xkqVF3ShVTtQa8ENTNrBBtJho0waEDPLRchKagw5327NJo70xhacnlEYckmQl
oHcH0F6QT9nhJiEJ2t85JX3XM1p+1EQOrJqGWx6jw7GSV7TgYUxWiG8yYWXOQ6XcukUM4TeRFUDW
+dDVUBSYDiIHTbuQW/vQxcJBTqijMzXAhpJyuRTItL4NkqOgbVoNd3iP00MXgvLEOZQeo5ZtdhBi
Nca/7N5gCkap/4neEzBDRfqCFE+pow/LK7MbI+tMgtPYRfW+qqAxnZRyu0DHF9LUEUPQ95nJJdnH
vhc+M+I8WoQ5onvcFA50auhRehpjzAVwYCaV5CaAH9fIfs6thCN6GROGSbfaYolhdh1pbtNAZ4A5
X3mkDjq6vhf8PCPeF1R35lFBCzFwGoNbDb9en//Ul+GekHFiSwm1KvdonhyA2vVrZEr8GyXfu8xm
PAWIcylFRjFgFo7ReQSTt/QhVOoC19oeaHcPfc/Y3/UUdjPXk2Orj6u72vdNgLvc5zDDTEvdhdPr
+gLV5w3MGMAZELh722AcuNX7qAHAUB8d6ZrflvIAFIIz8mEwkp60O9Q37FARA31Mt+EV6q2f0+Ln
fS1ejLBQhpWqmbPdatwG7Wf6b4l7MUIGX4QyrlztPqEyA2dvLwQ/kJ+WEzV3tKUkyrnOwj0NUyK2
JBYTuj9FzjSH1LD6K99VXCPWm0MO2U+bM3IR5AEcZweWIxZsrP2Jtuy2zlz2MR1fE7RdM12MYuFW
3pNgK6oil9bREXAma2dOf7AT+Nobt94/K0xOeMm5Pfb5yufqWks+R4spotYfoR3aFk/XBglddwlI
RBKOT7tkXJLIKxvYrRU37YL6b/VanLnA7roY9jQ934YoEp0D6Ikr/a/Kf1Rjc3u3NO6exubJfWEv
YffsJRDALatZa8j87f33+u+VOsDy+cDqVmMv941mYAb19DNJBotoqjr5XTocga6iY/+tLjbrzNZc
Vh0KfT21IqELa/NbFExvfahZFoeMchRViJaGb1QSxYd3ulFBoBtfV9s8aMBQQFztjj+zIObLScMO
T9tb13/6SIprBVxHVwmfyMxnmx4LC+KlfuGz/63KNZPcxF/mzglzfgi8Ieu0NqbNo9LpKfEjAjD/
DxaMd3HYYxX/z3HhSzfaHeIwhhqpFPhhwloXMP776za5LWzJtMEl3LQzEij7XVy50mzmvK3pTJqI
Vl24boJkmglOS7vn44b0eaarJQfLZ1EoAAEuj/s55MWF5HmXH87nFGkyfy768PqnlL8KfUGHuXBU
2qK9OELL45kQrUoYcaghDQwLhIA7507/39VmiYMbqjFpBAS0YdoeSjm3vwiOQYDHyht2RHQ8uJ79
OO+0f87gk21+cMhv8eZEKZgi6+WEwlg2t2LHF+oqkuHZAEAZIHIk40DBdYXyPJs5YwvUSwWaxP/E
jckKXOesLOF0NIPF6KLXoUDepNMKBc193x87DUVhEAFuAhu77qxlwMMXWxdTHhXq5u6ZVKvh3VoV
ozg8jwI36YNicZka6OAK+C1Kzh+UPTYWMFJVxyx/YMUkMCefkC38npzpYx6mFPPpl/lYmZwNjzFa
hyl5O0Ykc5XgRHe/l0lgsFuhcQREbZ46euJrtfT0JimDDk7FHq/MhL+rtKUcWRCv+wrtJhWnDFsg
gMn6fvY+2JrGUElm74nZWvnWdWv3s/ApoFcYJua95OIbsYHt7EP3R47Dye47V1ytNtrmpEUdf+sN
5Ad2zIPR+XJwUpgERlPHrWGPnVnJlNlsbNYtKWPWONuwHWkfaGi4GEF7wVA4YhPaO0B/eJiR/peN
72idUHkmR8FR+6yUsBJwZ7A+OV/2NQOR/H57Nt/2mpFZdTMG3qOD+T+7pXDdc9f0Nnull6S1Gj4t
vH37vwq7FdEOt21T+0R1bJwJiBYuAB5dwZSuhaWbHeyYFCgnqW3GeCWWxHnegWT1IUS2nPpAkw7X
vPe/q+70RGSbvGMRQcagKBdg89f/YVzzeYZOuS0nhJ/ZKbKj4fPOtHaZhaIaprTRzIrTKW9JWjxZ
SegdzcPXc/fZnJcz3CEPF/JzeybsEPHPh7o2oaA4WtCD73aH9YD1EM4taEaYmTNvI68EuMQbMhPw
g6NkYKwCzhY/f/DtlKOjVySP3SKPW+ts5bWiMtQ1p5n59vjRmw2ZyQdP81DeesR7YdbW0HB07JLJ
y4isin27ssfdVTVLGq9siqiAX3DgCm7UhVUnBg4nquzpmzs73jbwhURU6NpkPHZt9WjJ26gUs4op
0d+dP4N3FydYBpUG9/03e6cO9bY/PQX0gx7xr+3gaf6JkusJhjIRO02lBrF41srdHmhiO7L428gH
FSdcF24xsowM+jo+N9b1Tuua3LxaN37NlDH0iGNIfMMCMWUZkGZzM0W0oF/OM9H7NsTuhrRDsbAc
3hokB0lf43sjo1cqPgV5QP3Fh+0kYmLBre063IQHSDhNL+u2oG5ts8Psc7XpX5r8qW6X77EwDewn
foiaNmlCKCWNo7xko80P4+lOxwZm3Y2SDm073220Roq8yyWdsSiyGbB8cJH2+uKvns/zmHt5SnWj
agmcX/bfEvlEdZ5LbRdawtOm6uabU9u7MguQYGEjKpBPYum1Pl9/9Abb1z80Y2pGMpEyU+5k9ZMy
WgdCD55xvNYYzVVxpfwFstX2IsGlzUuKqeHksbFDG9tGpM7Sz/1Io6nGNvXSEXaLwr7kQoyQMXtF
xF7C23Z9FcmNFcpDt4i3dyrQ28j1EaJ7ig7oMy4yxMDZ2EwQ6fNpH0tukRIRrNWvCNKHkoMKm6/v
GevVUhr3HBTtTkN3RtWSksyLpqqEK8CPrrXzxqF79mu66zcDquIadE8hHtAJE8ChsDlsxVe+Pu9Z
nCpmUgQkCSwpSECHVxFSsNZ1fBfdxhXqINweLYhuCUV14eWRbnXQnbH9jvTHHhyZwHZKi7xKy8rU
DK5q6xm3EdVnc0PoXaf7fDB4JYuHAM75EOH5v/RLwCc2brTWd06fiAbRaQX2B+woajERHHDI6WmA
oj69USeCUtK+5WUzQfflWnxwMoTM1Dd2Nd51Bmkuez4d8Rcus/Yq8kBtJ0AVnUWFPV5Q1hkjpXXi
Dh5tRwtFqVqJ2VwKFIPzuzClJrbRjBfv9dfccfJLh/ACLtQCdgmLdiCZQhD2qV8GLlag4xQXOB/P
gfYQXZ3rbPJXcXsdsNvDa8ODdAAeEIdb39zXWNs/gbBWsg0xc4Tk+WmK9VvCCScYPqCxJxCilts3
usRSM0ImV/SPZRA7jbBQKoMcgW2ks1ISmGJABd5vsxuQ/NY4QNZJy2WRKAeBUoL+kZ4h4y/cNutC
r5XZYHoLm5vlP9DYxMxKFlKgKbpLV0LB9GLOs0Q+auWG0w/hpLB61txZ4qTijnD4OU9mWAgwIth4
q22HGY0RbArnXRD6LWW3VpKfL0c66ZNv9JDCq2ge5ervDS4//cDNl+oNxpjFgsmOYgT34FeZDTBs
abdD2io0KDYxvwgAcUnyTkp1W62B9X/O1BWKvxMM3tp7BxrtqpSzYMqZ36qx/7FgMnEw0oWllY2L
qGw95SnUDiI+UiZkNxOpCLGVev7PsFfa8wguEeujD5k7ZDj52cf3oi7qHjnItECH6h/Sh9b9fW32
sZzqY+gwnkHkEjIMiscDOk5mVvtyaTVDjdbc+JB6llOmV96PQhXM2v9Pz+XhLJurX+3giFymFo4H
PZxh8dmeTB8lV58bdd5o7XPRsgSdzlkaZxCkTUzedHIVH1etw8pB8WDDoL6d5cNik1tsY1yFe4SF
JmTJUnHy6cYQG//BAWek+2++18bu4OWw/GiCT6EnvfHReeakgpp0mDJEw5WDkQvom9FMeesxkqZ5
KJLpKg37cvz4ahMeC/IEYhYOwyqpUTsNqlBQMOPTFmpR/wO3f+XogJFkYL1RqDOgNEu6/dyQ2sNo
EIRf6Uy7peRHQBl2Op2NTrxAzLBCtBnMbkgDQ0LnJ/KBJtJoYWitxqgwcYy1PCEwhNOa9hAbgEKo
WuYzl2n+QoaItM9OmxWbC6a+ICRny32HrW8N1qX1WUML7UgG+MrmU0fxVPDWzEdmvyn2FqXEfZXv
TRLbfT/RUi8l1uNU9dUyJMmS+Vg8P/eXybDbyhi+dlR+n0UGQYj+BaYB8DuyFz+1LVHZ0hzLnkk9
2aWYXJhGsQoWEWK7K3c9b9susR60N7mZvAb/Q8CUojGqMJpJ+yBwJc2M4cmH9dESHrSASpNurfve
nbxJHzdCmk7jHz9FfIDX5D5jE5L3S+giInuoLlDtxFSL3JqxuSb5NoHV9AjE32kgS3FmP84PSp/M
KodO9MrdsdNn7uD42TzqpSUx7ecv5W24HXmDpNkhgKCTvDuN58Odu6K9qouZWXz0d9iO5FWa9feF
jZbVqGbXPYeLFosNDVlaVb4RMZmBJ9L2QJSIhl42L/eQGfOPN0jwyFTRyoUBM7yfa73aaVjPIPqu
jvxSO8hdHAa3Gv85gRSrP4GQYzyE90BrDu9F2og419OoPbwmF8vZiGSj2pY7nnVwKd4ZyxMCe6bE
nbOQDLpevA1kE1UqQRVzT9tYrd2FNyVMONYqes4CBffrNkM4M6z4psWF6Fo89XEggMhgrHWwLhkA
pwkyTKex0J5xlqLodk1CS/VKEsnPoARGQA6mXp5uToY3OlL9tRSO/qmGjfj3ItQSYPHn3z2clJLZ
nZfMm3LCQFUrBd90RYfmTUpdugTFJ7lk0R091TVv4+MEJQJFvWNSNVcg3pkUERPTWfOuHBCv4pZ2
jesaZ9CYy0uRGA2kJ6yWvXXBrIBiTOSw+3evKpcuSsA1NB/6ab7nGbnCQchGLF0JPwObFP3gYSt9
aSXuKujNpGhVb0JxcEFl07zIUfpOhruWE7FUCjAivrYpK4XsMEQ8ZiDgwZmWUoioktFcKWyC9Fcj
QWQVDvxWU/tHGNdhEBcxP74Ul7KTpViEq9F9KpeQDzsYu2mABQUav3MY9KMlfVodjDbz/CLBNaEl
W7kCVsRk89u463ylZ+XSYPAmyAhAy1T+DJObYNTvCMWfAjU4uAFLYd7GvkxWPvtR3L8fecydTicZ
cFbo+pBzgln2bl+8AKP9KKLeBWgVPKQveu+MwEnPuJUI+AHK6hoyy7ZINEjNO8M8Ugvy5iH/JTEt
D78fGufzUz9u+jBOQlVAHRhMZKwE17P8yKzL7yF4GxHpc2WWrNfzR6z9YKVRriQmVgpuFaS2GpHO
gKBoW+y0CWWcjfTU7PDZJRbzhfjLRN7pydTMnt47877/UWqeVhean/NcqVn46Nobs6vHJtKElAsn
y3NkCorAkhvg+rJvDW1OLjibvQ3XkQ/r/YH4YQtmtb/l/6SeaBMUXS8TABZBgz+2yJDk5bdUjVaR
8ITLHG3adu3JxuD8RSZ8CM/nZLJ/QwBRLAjeh9t8jJb15um8si/iZoXk1iUrMwWbjEC4djxyAlfw
2PeAZnWDB1Oh9jfKAmJ4VEJwndhk/CEnWzFGT0RQzzKJEq25HQ0wbZfiwvhrBGlWxkJu56u0HAmD
VKiChNd6WEORmbR2gRKm5QR1sQl+mT2OilAw7XMbfFLW2wNDaLU4wrLyxIT0Vp7QlMT9xqV9c8qO
L3dbr9/k0yJAAoV71XdgmaSx7suNAu8Gfe9IqsdFQA496DB6TY4wODgS9scrHxBK/4jq30VuIsEo
7+Ialm4tnO3NzWys+s4A4rYl2GCdAIfz2D/yoPedOuQyYyvu4G4N7/FLn5aBUoubBwsmOS0d93db
igVaMyHL33F+c3jBnzHD/EVY+Oul9Y55DHeCgbRLpUKxsRoud/3LyR+IbwO2+Wqx8JNiPSHaPX+l
lktUTr+OmNNeSOO70DWz6rtnLIHfHIxHKaTYOHE4Ojj0SbJjrQdTm2wSYMgO5SG46kRLMYYTEwvy
c/wzDN8YWNB4sDqOBGJ+moGd1+ekZhZMb7D9rAQwVlVSU93RtQ0Za1Bbb0lDqyQpacQinWLJl932
U7nraiouZusNHR8ClTlalLhCOsK7oICF+2EJPlGvRLWYcr9MOCawqHNbqMpC0VbKgqnH91+sFqzt
LjGVPlgGYwXpY46Skpc+MS/Fdba4PUVwdu8+MjoSY+3s/0ZPymDK2t1FdIrD4DMwncwQmFeUrjPt
rh5Yc8G0ejawP3qQY/LSciHaRvwofQTvzfgRWWKDc2h7KjTMq4US2H1HHG/vEwGLb6jEaNfxC655
H8mGA0RB1yDd/stBqh5Xs7KE8eXiIRK6Z2C8d8RNKrroz/K1IYT8Q79wbnKk5m4hKMtyTXskoiQl
jjvQ6+Tp70/5mvaHr6KSt2zd7tUStfkBDs1AJA/YrJU+GL0su6cP05Somewi9haxhCyDP1FI+uhP
7iY5cKC6+OZQaUlMLcn97yKsQrFnWBnlGWk1QX9dcOw43p4IDYo9Wg7CYdexC1RMf8K3p6V46c6N
IBK7mQnmAa7K5OjecrYMWqdRtTWn0VvWox+VM7UDI0dSmFtWwBU8A2qU/WYd09xF5iIdwnoKHi+R
egHkBGDy/YgPrxFGye1sRvfyHs22j5Ff0eWNn+ZqmZE/yHRn/RVdUso773ngWtoKSk77vvGJ0R9H
MLzqIBlbh0jD3AVk4aXXeSS1d5fejb3C98jpfIkMUWelr4bPJEy781vU3EsAXE5QVGrLv/CRVA56
VfwVjErHOvzAWHNQv5BSBOvfXHYbxOcQLphtp9OtKM8lcxFt+PxIGVhi3Ncm+/bt4XW1Of1MPjUk
cW8nASBbc0PHK6aJpY0LvqtyzZgbgRe0NDpLiqxN2uUpwcQf+pOCxvKm7Rhs21pLcG1KbBlv9BMu
a07wLBqzRGk5uNN5VQNNaHEU8YYupruIYO213UMvjYKTKyNsBUXZT1EhDGomSGbvyF7LJGjjBsmQ
61IX7xPJzxA0H3LyBjRZ/szmkPcF4EWWR59Lvwb8d1tRN/VlSF1l23SFpUjEK4VQQ4cSKQbx9mdK
alW5BQdNq1WWMsA3MWTZiZsE4mC1a7WpqQ8PtoT5797qJZ3hspcMtJF5sj2FQbSEKq56mSezTrqc
cdHkHN/JMpjXzq47dpW9wJ+L+2rJnNeqgmv4VFeUuPkwy63A6NxWSn2ytINJj+KoKSs4gCgthUFX
6H6duooP+YmH7rucYzIHgvQRqSN6CGHUG7RgXx5M9yCruKKkRqAnb4G9StHAPdGEAXTXRW8ZaAvP
PMP4TWK7ek3ALfdNnApdn8RL8H177cXF+g3+iT4BdepkV/Uq/KKJbln2GlLacFkE9EcKAQrw3PGn
+dDEtxUUvGDi5POHd4GeBnRDp2eVNB4M7E4IHXVWc0+7XiCF1YoezRv8tIACYwjRQRNbMxzXqhbS
aj6m43cgfQXcJGAlSRWNj/NwbelFm/55+FO+OeW6r/JeGBiAJGL0DcW+v8BBinZE3fXB09oAYHaU
GS2nvTTd5tO3g1V6W+mhndzI4KNK8T0vRiXJ3cSdNFTWk6MgpYlnACO3E5ge0lLteS9fhI0MvrKY
iywAfisaFwojjQptRXY4E9K3avA3hIYC+gK7MzJXeofyvhMrYuNN5/J6+X2raVhxVXAQggSN/a1w
MiV8WnY+oQDUp5zWJnYKZzv/MKMphHbxFexh64rEGqetj9f7VuQaSnCKEuvA2ABVrxpxJ6JwtSlj
tUU08Aqrw5BisTFdokKaq3UyY0Z95QXlXimpSj1qc0SNwXfcmFktswG3qLCh0zzOKB/5bT/blcjN
tEvSU6vfcrxcACO7vad9XxNqplQ7q4sZT+f72mMQ2IfNigvBdlruWviLhun0PU5+UV5T4TX+PIVO
rZQ3hoIPKkKOV9EJseR3KKjzDAAeYdOZUUNj3SVd9t0ajwcYJjLkVjvDmYqPr29O2LGeHgM96ni4
3OhudkSgQC5hHfu9PycIJzSZzKv9ELuEvXfVeWNEblQfRKjEMVmfeaOlLGn+/8Cqt4QMT7gUrwx8
bQAhLx5R00zU2m4uL9tnvok3fjt1wMxsDZCJCrXiYddWZXI2XU9SGWk4jt/5QWddFi0xEZlhc0s1
AOjiEd5DV8nEm4/2BhbucKr15UFzZBAXKfEJB6xh20wAnTAAWt5erIcTDRXQ/KLuZdmC3Ut32px9
t6Ba641hwEPU2G8RVp0gO6cYmpWT0ikBlPN3D2tjGfl8Bpy4BxKLwK1dR3ytHmZqZXhS72oupsyS
oBCzaVVAS3+JGCpM3iU3asgdbYJLUNgTjqPDGcxP6olyzIJm0wmnR+nLcXUKqeD5BBsKR/UsQMEM
1EuGjUXUMYjxbeav7xMmFNXCZ+wBeKrvme+h5poiaUz/Ax9qFGF8c8gGsTh4WTB2XlQqrjjaiOzY
CcfJQlO58N71rjcOk8S0oacv+CcS+0iXfPWiFibQCPOv6Z2QoxqpwvaDZTfc4IOLAL6kb7EmEVuM
X0ALVtqZT8iyMSDDMk9lL3xDcQa1hxt3WIhdd54+NF8hpEWxihTZTJHWQOrD04zO/nW+vhlp1lRd
7Da6iRY9gq1SpAPyY7IGWi+pGydlpcRgpe4KSiyjeXqzbouqZCBGNRYzagsPAjfs5H+/nt7oerlJ
19QFgzP3LdkAhzyQv4UTnmzvs6ze8vTay8ituoC5Cfjo14Tk/d6CRStRCKp3wPopr5m0/qlpUo3h
yNh3kx4FvFmtTriQPtOMHG4CLh8Qz+7mEqLLqg+zKUugEBeNcT+DNa1vkfCO1K8rH9l5kRAvuwOt
dAxPKdVrLRaJCNoxHPt3U0axfZ4BHHhAwwRuRon2gXtunriaHUa5W9SjxgrRefvxz9G+M2SKP8u3
Uz5YK/pZdr0TAobLbVa29k4f5fEglmVIdijke/Ba04FWSEPiWxboKXij2EQk//hWBfFZCUdHAiAE
CzvpSOy7pjk52MCmbYkDEos3kTy6DLVwDvKfKxkvxaNANCX7W5TmWF5y0nP3A1NJiWDz6ECErqx9
C0WJK6iR1nqKs4ZCVmTA/6TKGHl5cgpXON3GlAfUc/xZdfxUNk9Kz4xGaF4C9ovRb2FGM48XuM32
nboIEl006gG7OokoQ4EwWzFUDAW840f9L1Y+UxdYKJ0V+pzV2ej2dom2qdXEh7JpeDp+2oneYnwS
JEvuhOrfs6ArQQM/r4XpjTPYDNLu2YeICb6mIR+f969SoBWizeoT8O2TtTDxHGyNr45a9wKRcUD2
SihB8w+ledAu/jNfB/tC3kmsnfW31OXPfnC6YMBWaQnSC8blnmVNuzR7w0SMIFd80WoeZy9LeFzg
8xMG8hLLr4hpfqfoFJJRC2to92aLXyW9A+8lRY9BlwCTFleLpfP032uwPncOUlPntcmZDq4YjF7C
BI/oK/rXbFKz/1cDu9WChEfAT9fMmZNhZxgkBTNDtvcWx/kqqVgQ6bsaqhgD1Z6lVotWmbs2s14O
VorWfBuRQRlWHjFe8xXhdmjhHAorcL2x/GnBlZmIrFLPZA2+MsccAeVa5y/IMgAgYYqmK1td40aN
Akm+fhj4wh5vcXu4RXEQHogxc9FcslNxOQe5quKMO26911L9+oXuFMLdvh5h94z3a8lmIfUxEHt2
FEFRdx1JMFOx8zEA6RqWwrypL6HiCGhqcO6qzq/dSGcCWAv6KOJXkJtyxpUCYGuV7T8Zo/yxWLg8
MvzR8YMOHAFwaJG3UmfGN1B64jBeuzeQRx4yY6+doPoSO75/8drUacnHRR/WbToYOo25K5QhKUan
A/qoMHeGUGVsqS9uQrrNW9KYX4oQUJSXh0AkAF1oed4TEu0bqyLpbcZKet/E86xSAEap2JLc+dP4
ZiKD0audxgSznUDutmt9zbC72d2OAHj5hk6q0oT60mTrkJs1hilT5pCDM0jnhA1fmrscDTPIhKZV
2rLSfLUxeJL1xmXpMv83pAU0iTlxOvdiwKCcmwoeU6hHrm4OqeM2GwZDwJvs0bTUS2bo/J1SV9vW
zPhttATeJMGVrcg0bc4pDJ5m3IRQaE5aWit+cZaPuhgRIFOG48uLkRl+SWxuXIy7cbCIE4t9l+Bw
lo8orB5m7A+qHXD4M8j5zZDXS3lvgDBAW47Ik6+KjTfF9M3zBRZXHNe3mpiyUeFN665uTLQFcbrV
TibnYFAr2QYi9yJdQ1Shq9+BkOX5Z6mJPEmIfdRg56mrgghRPBZORQFu/3JihYB4vDddy2MzftF4
i0WwyhRpf5LA2fVdR4DiHqmk07UbiytmXfp11qLakGrNnHisK0I0STRMJk1appxCy4X1GeKDW6i6
cBMcT5DEWW2qk19elX9I7A1iZyafPQZi3K6xu1zFaPDGhSiD0Ckd2IwQn8noRQSGyODHaglpSj0p
wnhhwcFrn33dcB72eAwXX68txlRH+NNN58babFIm2Wk/s2ldgDKpDExqus3VPC3LiaLclO9mjjPY
bxtVeaTiJRTjrcm9BR2NLj765piMEznlHegmHR18ZvQ0l0VIfN7NpbWEzOP9ja1dHG1PcOP0kRNG
aquhbW8tfruMMzBttv/QWHog7Jwh/C+yag7wVIIqUgyagxyT8E0eZBk9DEWYXajn9bUBmAPrpV/b
qIZnGlvINAblB8Y2SZhNP47RkMP+kDTAMryJPFEL3gFlluViA9ubqQ1xYNAR7akFpxTJv7rF0Jbe
TTP38P2RA55GY7hoy6UOREuRcL3w8fizh7T3n1wo1EgoumqaoSP0Dq2n0JsE1OtDvtilPfZNN1pH
oHhMz+PaUxTPAh5srzgnpDp+cTQlTOXL/cPHGF71Aq44BQUEu0BTjtwYCWd00z2U8Xn1iIDlaehd
JApIBaGbImBdYsuBtsGyX3QVf0a0Td86hu8lF5LarXqHy8VSSr9dG96K904v2AnR8yNpjVXXPj/+
F98BpUC01HDb/UpSY0n0/unhDOMxHsrM+p18wYq68qdkRr0Ax9JnDfijAb7rvl8QwSNMCmo2tRxi
jRFqEmIubvvN5iCRsPTtwc3+GFnNXq+qmCn1uAS0EmC4IyEGDGGN/DRnRAm/pC/EbPIh5JfWBIsg
nIh0XO3S0vfm2Mc6ORvay1AEv4O6jMRRQyUHLhqAO0M53nkRAtH8qaCJ94JeAPLoNDdqaPWVjKQ3
qGY98wxwL+mst4Fsy2cNp7NaUIsyNaaqFCVjWa8jvQrNw8R5q02Uj0ALXU8nIeGBtnFya8mi7lj1
DskCF+HWxL4xOrkis2CZ/q/9+Pe3HmkYpy5lhqd80P8B77q4wO9qnQh6I6AHdFfYzNykuj6v9hoW
JTY8Q7EWvytANTyCBYjAelkSsc14i0UtMERn/VbtpF5689VzhYNaydw/pu3LmH1lk2INcHxhcPKG
1P/Q16qy4sb6Cv/3Ktvxlz28gORNEGFlYEMFZuCNztHBfVlC9T/W7iT/YXgCRMMoC10UnXT91VJy
8ZAAc5yCh7s2vSgf4aJRVk6BFfFgXkUCBIbZP+arH/3v8IW9OV+Yc01/X1UrC5+oSXMU3Slujrhp
kiWFT/Byd3qaplLqrcvZriA5R+Z9DGHnGOj9ryYk0hJtu6/JqmEm8tkOlU49IuCZnbXroql77TJf
qFY3PX/Gv4sG9yiyNJsDcDyGVGEuqoJ0vLZNDAQlfJ3R/N2oi0jOt+mY9shpz9Alg9h76qKLGWF+
X8Me8OqHUEYcVjD2a7sXnpIIHeO2c9+xl2RtT+jm73N+GznfDgo8Bh/b9dH7mR0n+WSKAcQ/qNIx
joalwSAfvFeyqtmoIdNrR3t0Oof4sarxUS7f7LrnhXl79c1cF3d7gknugXKu4s1FvVKGc+kDKFam
I4iwO74f/l0EWbGWIZ7H9Epa2SUPGLCojyJa9UR+iYJxyvwpXcojjL4ztX0U2fyitqOu6KXJikLP
8ErKYa0vSBAAoNGTrT+Js0kMSbV8LiV6G0m15Hk4EvyUQ+7vLPgZL4ngXjHiqznnCXoAt49WPL2J
txlsvdXhuWytmHurb1nNx0Kq4XR4sPCE0+L0lPq58p29T5BZTcnDKxZiQ0Jad4HlhGCyMpGWXPeA
hRzjSe5wJnTnDS1OFTo/n2LPOLkeqJvhqsb+aRI1Y+G/iXdytWmz5FrBZ6vDXY05ReMuIAHslegh
4AdVw253YtXrnekVZfAJrz4cASyOR6Ggnaowxpk810gZ4s6qGfilGULan86VGnEqJ2zTIz1sXjcf
IqKjAtokheU83W1wJfFcJrE/MmpFlMwZx7+dolU3UuUEmYYlSGBlE5Rlv4ovUj3EOrxsbiPglwo1
s65JAdQNaJJyB6jfgYoY+qUyFW+PhAF4N91gJdVrTL8gQhovr9LEWJ++28O0ABZqQD8DBXBFAy4t
DCvebe6aGNtMBfj8XoPAhvLbfjPBCktvbxGVxn5huVBi8iUURfrUbh2quX6LoHa3r9JCjduwq9nD
SHxrHP5tATSs6+cY4iqRU7eoxrw1Sikj9zLX5/OnvGpc6MYmWVOJRBsfVNehSkjyevPJCBAtG6Ba
ZdxntpoqBf30kk7Pr/LbTPE5e9dfCcBmO4KSfS2AqpLNMZXOjSjhVnRb52qNZ3b2uwrMRzUDRlyu
HNDV5n9BmPCGltXwc8nX61PszuUcSMXvalx/FU/6uTVQDfDgkbJF4kf0i+8LOYaK2x3pZkMooRJ1
3Rz8adaVpJ8BOc9o/N98fAJ8q5V/gy+B6iVXrEQSK4sy3J+3hyoQCWBNLp2YGagRZQT88EtV+/3F
2HKsjNZI2FNKXrd2W1UrRitPkfFsucllcDO6FMalcWC7Hcqkjpfmcgy9NQqDRPWDv0CybE2zxjBL
dVh5MDACZXGxqT4sQ3q7G9QG8XlYlEg3S4KghSI6d8P59zwe1euo6cayQqSK0Zzt8MbVzDFkNxsG
ABx0F4+N6fBKyFV1msJh3XCUl9smb1qxdI00Pcnoq2URAPQWJATcwlAPHvkDCFJD+lAedSEz2pZX
b5cCwIqxqpCABrbRgmEF0WiUdu0gUuMbTRZQazkDVgIZycMZ87C18CC+CDJaESdrL2dC2JHq9IHo
dMbToB2hMJud4x3HMcz9Aznqk7I22n6sXfrsA/y/rrdXw3PCro7vZdDJ5ReiGTsqW+/Sexdjw4WA
fGMTK9iPnksat0QAAL8Zv7KA8tuQ3R0RAP/6vMiT+BwJICcFgC4zRBwJeiJpUxOcANL5I8SxXShj
VW7lQ7vVRa7nU4CD9BvLD/Ha6VgERbNMheXYFEclFPuE4wfJDno6MBNnxD2xwe29j4Er/lenxk1A
RzRNvMJIJevl4S8IKLGqEfg+Gg5M5MFPfb3IUPMLQnZyHdt4gwKtdlX5ixky4tAf6PJCUtLaHs0B
Esl65exowOttHm0EmqbgNowNHCPBsMxPUbcqFNxYBvo7NhupK+91MZtHBaHvuUxgtr521mV88ZcS
J8uSR/uOTBHXrvK7KLkp8srA9A1BGavEZQKdI7q2W6mzky2LBS7cIsL7OKLvKW9bluzIQRmysVqb
5OJI2WoRdXIX7w7NRxBcyqqjp5cGeCUz/YmjF1YN7/D/5TE8Er+Xtzw3He8qCfDV96BfkIb6N587
QyyWPV0iSyQDp9VvDxAWWX5PPKG3Yh6Fq8ax8GmDscbu8SWuQHwz68s1ZFEwT4UnGFFo1eQyn8zP
qgjgJSzCbGCG0ozJnaq1Fmq9THVrJEr+hjb/DBXSZgfCuybM9klfeJRnw/n0gGOTbJpzF2k7mCGc
CQr0Kr/r1COqdzm6dd85upIbRPeg4LPoR7TMxqND/33rkIy0Kl1RwW/JvVkH/wtO2fLF5Lm1Jnql
l4qhW7UGJi2Moi5G3hNeKhlezyuDSEKcPhYm+Jpndbf7q9auW1YahLXjmLrTpnXHnoPgYoqNITU6
UZOtD24j+m07uiwWV4rCHEAruzplNbE0dmrx/HZvctsBIBPHW6Y7hAlR1lrm0X/NWAgh4UsujYo7
KM3tUb16A9mpW/xVOQTIjjOCOn8BXjkoSE4+VqRF6KjEzqO/cMpN4Clsa+KP+bIcxEdc2HXEUGMC
dhny95ekUMUV7uZSgHaluGf+gJVDQwY0d7rTZ4d3FQ4MBhjpkrySEwicmsbTZ4KiKjzs8mmfLU3A
4HPgAvPSLgmypjVsVJLGYOPNdoIvRNsYP6Zx3Ln/OPwlK5wxxcAiyuVuKEiHpaCJI35aIhQYieHO
GmVngz/dDogrZQz7osBlmh9mTxVCPucZV1TN6vappcLaFDJwFKf6oLhKt01zDwbs2zjxBKCINIkx
8aQNIcx2cQdOTR7VPP0nERKmTImtKQPw0EHFCpckfyxK32T0KsfXi3R+qBUIFXVUWSZM1TLIXKog
ryOjFfvo1CKGpFjKGtWdr89mP4SGaLUXHz8km9wCyFs1F9Svh69hyhkzjRJ4NdSHjp3Cigp4ZjvR
819FJEjHHayGcX8HjhHPB2npIikkVCJ5YGkKScfrgcNqgsIVpyoUnc93DmThgkTiJEHsQWZTtGPW
jxE2JgX1D8/tOQizqbYMZnj/KrJrP1pKye26f/ZfQOts78cqTikHrbDj1G6klJZEtVV8DdhiBiZU
omBNS+cDQLThblW3FEs+XX/tmwQ/coMT7vR5c6emH/ASFZQv18Gi8EFnUN1onNusDztu/NabDtXl
V6xd6YcqDBlpZkX8s2kpn6OtHvhh6SNEdggKwc/7/WuN7Ju/58opec96h9ZyBldI47M7m1jCMfHA
YYDoONBJa+UDJGCkQ3dp1BDzcseKSUJcaTjZkOrHoe/s5GObnGJAVqtsEBtPwpMZvgny6Rox1LNX
WhYZ8ExpU8g08ibdaXoe/r1t1lvtluFKu8ewQygXh32qr5AhwlqIFogiekTyFkdfNaz2ntbG8kk+
o2Y8Z7nIf/K189nyVNtnW5sBmFOgUELRaY5rE/fj82SvY0LZjPVryeyRPz370vqg7/w0NDzKyo9Q
+U7LPhWrFHlXN4Zy7QmS6yYs0EQn2rRg77HKl7Z/SkJDsveWPcctx6jC/y7sxkAFjEWgQjz9gcQT
FRdI8nmbhSpjlDriiRirh6DklDzuRY/mXdhwIC+pNU4rAEVZnGXef6ivrxsx5/a+7qNYchehGDZD
QSdUHzZPQ+Z4VLXVdtIGsmu637Yb0fZgBYq05EGNtIlby5/ESL6V/rgBquHYxQYxfWhxAqPwIwJB
LGo+Iz40BYopsEI0pDEgQu4lO3nLLh3a91XyH1gsMLcWOIE/Fu+AGjPFpwNbAxSj+xpDn8AnUSmh
+0YFjjwAYrf3JBg+N/gxQ+GRxHTUnHcr+9bA8R35CZ0I6XQBf1bD5nVTDlNyFax+Zn3z8gbmp8tY
peZvmz04zfe4CFdK6T6KGz9dXHfMFU0est/MLi3sflieg4gncCSuwRa82RED6cTw134rEYBIZctW
qksRRT9n0edNoWrduKUq4qHlUJFmX0rEOQX64EPzG9z2jTN9h1B0TCVjdHAKQfCrRu9s6tqdKOKF
Px03OW5NXnakb9h3Qp+YuX9I5z5upwUBicRR5TvFoQpt0E0opGJViAjjs/dK7hBYjB1CLpg++VA7
aEUrJVhAABayHvOcFaQe6dC/t+aaMZj5L+Y6tH4ph4HefIcZBYpLVReCsIwfmPbym7bfZWHkImqI
br73rrYEzH7o3qg3XeAvz7kYIzRmGWKJaIn3SqN5OgQ0CoD7DCvw/byfxrW7YTOKK5jGuIezGn/F
jyINf3ZUrb/5IW1fJ30+NZ5X+CHS5xRqRYtB3PTbeOxAWqkmRlRE9dVuD7jurs/SGW/XzQVwg4fa
BkpirLZ+py8LSQUBrK40fa0iHjhDJL4JftO6m8fSCooSI5ZakD2N0/o/ykr34rEeTYoyG+gRIwkG
okIgsKUar1VxLgursVQuQm9gUF1n3VV0jB83peWlRRq4+tfYYdGfjaVGjwkCklw1s02hdzPxaG8v
SuHA/45/h7HmbH35iPuqPc3/gkZAc2i689aqa3t/oxABIGKdQ1c1sGFfuzF5dNfNBQ2qqIgrQ78e
d5mGaVq31AQ+roi6RbhjhUGZyrpOf8J/GJgjLbRFeADjgQ57VHvP8OESoKmBFBAI67HsEtCdJJLF
mFnQ+2pzNBR9VFhWZ5Xsoqu0zyYhbJXvUpqq+ylgaL96QD4MhCPHNmK8iOvittde+C9Ng3XTapn3
1SYoe8OVISRUjtZKlv/FNyJC2HNaS/W06WA0Vdf/g0Lk3CTrqJbWZWXN4TaIPTdVhzxXuBgG3OWa
quoReBIhBOnTW6VV/xz5V3xJXpguDjgeKzAQcfOLdcm9tlFT9tCw3F7VyLG0OTpvfFUBddVBpkNm
0s4c73dJiYqD9sov2wZlfq9Fyd6CRwJKdFBE3XtGW0PJl6gGVfS8qXS+AhjTm8PT09ZuIjJXQapX
z2xScSiRdrxEuESSgmqQWK3TwxHJUsWD66eeZhV1M68lYK0pnQ8mIebr7Uf0C8wKF0OJLPZSwy35
66bsrTomxtCbIg1MD+baVDhfTTYRVk9kWE6+bDcHskaUz0HqkczvaXcu1wOjqIkjJd2nhUoVP+yE
yYEloabNGRhJFN2HcQ3LuwpteiXP/OxAqNxzhVZAe/TyWLtCCOT/UNWgfYqThiR9g858n94STzm6
J0aXdDrkq6NeuLV85g4h8ibprXP4NrKv1GuxutiL6t6GmQQhxB+wwy9ee+FWG2HDQq27rnTvVwnu
2J1RBwqAqbeESKCAj0+L9XGMnxG6NoAiQY6GN+p+NvUbHrOMGMzDQbJ5eKltPFiMt0Eh/jcz8AO4
Q/fhnlTcNyqsq4XDGq9HdMHHKCsrktLjWhodRI+75q874bds+X8aaD4JtPb9aP3Pwt81KNpHO6zw
8lziiKJOVKj09UFhk+fGOV1nUwo+2w/bscalZkX7yX30p883vqz2VQsb/GnDIN8KZyr5DGcKRft6
gbomS/bpVOVfhzdWzuQVMlaf+RyaJ5hs+/5Mgmm6gFYkapjIH+aiwAASWdUirj8Ox92HPFuKnJF9
Z5HYWzusOez0U1Pteo/+BUC2ENsgAljV9WZEqBdbT6b/WJoPtdtlT/wHqY0n6YoRqHKr4Bpy2jI2
yT57fs23o1P8wxP9eOD1BX/3wrC5OYkeAf9KrVS91ff65IAYNH9NuIc3GSPs088qdQaA4Hdpfj1R
N4Yk6XaU+NWlqr+Z+XTweGlsztVNaPLK731bIEfmtzZtIjIcJbcBpJpQVKFEHLylQ+BT4LcAZQLF
dAYJirjY5ujBGTD0BEA2Y21WKw4mKnrJsoTE6fQo6qRqBCSeKb8roCxTtb4sxhrFRclqZlnE76mb
mI6wXtRufkBvvDm4Pz6O6ZCXLU3tVImBowDrKFbzkhK0TwSjs5WmXoiM54B65INpWHPf7G/qv2n1
/AKHicEz3Ubd7d2MaaArEmGVh8Ob2gnNyGMe6lJxqR9EdIaPHdJyzOc+EyqU+I/iQ2jcanpiD0bu
8/+M7hYdYZE8L7swzpFUuWA6UdOfGccGsHrPhjaOGwl0qs5bkBhge781XoS996hYAGETZEmJWckn
U1oOnN82iGgjqDssYZ6agE44qJgbJUnxGCmkzA7zJAaTfMw4R411rx+V/qBA+yF5uP/2BxMBBdMu
2BXtdCuJ9bfTS92oOgv2AfZ4jnVUrATfJ15XAb8pvloIVwsS7QtpQxrPqbVCzxffXxLzF4GtU8EO
LxlRsABQxCvjEBDP9HitZX1txf6k3kQ+mr+/hC93MKKkfVxfahvHrlDM/d6jIPohRopdZ1w2mzHl
XiH5YpOIxNMwe2irW4h+KEh3O9yLA2yXNpQQ25nr7avfpi1I5IvP074LWDuLIbJJeXOVo9yWjhgE
UNebECWG2CVHBRo3mKo+CWfpfqSHtaDGcGhHCpOWMjwrr5oBIfRl2vGgNG/O0veRUNMZ34QPSIJM
VgkhKMQUUEmhBt07E4mnkrPgNCDskRMrjFgLKZzMoj0c279COjaz4BLZA9ojGa83pzeTjmpCqgUB
6vvbObYB5VLItcPzRew7I/grbtWn/XxlKWTjBxgI54mGG2IQZSWYc5Or3Ab9f7wjEm4HbJQBPlWZ
IrzV+ka4uuFKXgFoA7jfoH02K1GVAkLqduMHpmBxM3E4vNP/6Jp05nAwk2Jbj7fzXqXDjwiZUKJ9
Z52iF8RUsbm/m8CuQQOKorvjlg8jdhoKOuFA68k2yJsv/DoxK1g/xI75sCUK8Ug4a31O1tfosxIO
45v9+5/vaKRVZOKPnAgDfewB4ScwNNABeoiKMoNK15sB2sV7dzaljxtVvtCw/YJKxOTsl2aNZBWr
3gYlbsWQHq+6rOIuK35Stf0MqfROPaogZ1HeKaFNx5tXCnrj8NaNIgpcphAMx7ASP2vDmVUwxhur
EhotSQNF3WNQPI277nkXym+Wxz3t/9M0QL0PWSTZopR+SGKJiYPYPPi+zxMtr0BtXA83PlACIvf/
YXdcB0WU8D474jbil/t1Dyv+LlAvneTQMl+BFVo7bloGrjlmston+guIGOhAW48MVWJr+K8gWeef
A/kY2hRgbXnJT6SpLNsRtleStk0Jn1aEiMah1CGWqnkfn68h2co8fGrWCjW6gsnh0HEjBTVaMcfP
n4pUTineFUqE9Hlg/kNrcemcFalH8InRo/InrCsjd6vK+Tfg040oFmkby/ub0+sPN6R7mX2BJYAc
DW2rcpilXabnuhCHXZ3bVMMpR+NHJXzjF8KJVMiSzRm1e0wZiB4jCbD+y1MO9iNuZTsXDVXmZrr/
T4ZrbErCRqtAcpFSQkl5ITQttdABJRBkil0GJoYDj+lzOgBfOmG1cK3UJNBtgXNx9HUgO8uchjcf
Tl7NXsRvh9xb4X3uKWhS73cjGi4OQAiAhVXkGlNdiaalacsF0OGeDFavi2rAHhz1F4/i+0JJICdL
AhxlIz92PGDOGQwGWf4DlE1ZUclt6Xzb6zz7jII0aY2d5N/GSjgZ2DcA9GnvRDhARle4PE16Ph/0
of9MJB8bqc61+gCeFWwUY4q7KJ/qmfDTmpHOmJM04TH+to7hizmOXL8ZLYyEYX1mqXSKYbfCRPSl
9K/JgIY0JTJ+KCauEbWzyDYe5kh81+qeyHzgxcHAOZSR+PddA8GCaPBd/ccOlFaXFe/CudwW1B3a
haMna6+ZDqmO+1PZzWrlDor/8v3K//fv54EFqi8UAgZpijhVol91gIb6Lra8FZscs3/kJr6Rxedp
4W9rsL4HJJFwiyRMe2mOQaA7PWvEPVTmM+Cr7Up4Rm8yDRGumipKoXxoVkxt0tw+tvukK4gsiRK9
zJJr2kzK63c71ep16ZJ4jmcs2Z578x1bQzKQq5T0RPVM5dBDuBY9dHBoDZkCCJa87ez+twTWCuWN
JTrodzCljxGS/Rj8xY3SIkwjIuS9JVLG5QUl3eReZR6F1OLCZu56s9gd936iCtInJRpKpcHLu8tS
AVN9SjvPBwpPMOz+O2YWL0W+UtYGTnpfsH+iOg6yl+2dq8vLimZiWqBsFnTcIl23TyV2+Tzp1LE3
JO04KWvhBUmMVPAyZbaXRf/4kHcGZuLjYFM0vEU4XQZx/rGHNIs/dVMW/ZKIc5qQLfVVhO2w3cf5
tOf0LdCEJXoO279KGPrUUuYWq9HijNW2zKYbtt63pO1Lsmzn+eIqTFLvKETC6fjldhz30YrRahvT
Z+B5P6wZfZWlVINgLr+UTr+VYvrKdcqGkD+Pns2yeWIl0lzS00FeN9dQzM4tTQlMfEwsZIigK2hh
obz+WmS9fPujowwv9qJMRckPcwGB6rSm814Fmwwsu82zOXzhQMaF1Bv9/SjHmzac2WUXnUwCjP4U
sbRlYNDKiaIab2NV2MDTvCxVKlg6TL1Rlyj20zEqS5kKv7IwO1iPcv057UlncvwVUfxHhCRXRy1f
Rykf5o3Qf71CgEV+yyitg2UHQMDJ3v+eDr9ZAHs02qVnuL6qVU1DKLRViBP7rtMQb/wPCpddcIpL
QW9GpdsOiQ/vKjcXOip3jH31Wu3ds/Bb7JUgTrqMtcUpg2HOI78rdXwCUQbff/NE9n1zH528r6mG
JqrLthTPs3QrRrfRGjaO940zfEvO2NuN84cCm1rbl0/G8S54o6zbkQKq6nJcFUhZ1ZOc1htLfRk3
Xz7jjDns8aWw+zkGr0/UrXJJAl/en5QIlm0W5l9w2+T5Xzu6cTe4uV++WsOiqus06FmBprSNToQK
RluTF9LKmTGjtPlm4jfvamslwWfdlq8kb9GcObjmLfxP8/ei/YcEzHJnAmnBjqb33APxM6pupUar
EXwhb1YTHWLXF2xZyHAlGt1N7e8/nLRUHiQ7n6FvUA8kA2gScKyEMudWJ7y+yRDUHTJ2IMiv27by
ZFME3bYW3e1ZEHXogxiSaGOmzJFSW9kHT6oL7yZ3FToV9Rzjt2+6iyrWIKrstM7KsJ2DBvm1nR+g
JgIFslKy0RRDJvcFyf9noCcXJVENQbofgSa+xhnsRXiwWCan1miGVYCHgDwHrwXsPEC6waDFh0kS
ogYtxhsY3EMqlX7kyrsxbNRnvhfAswfElKcq83jS2Sco5vtwG2WMAz9fA1+tu/E5qnPpK2SIfaaO
QDnSzNSYbXF9/gsYY7sC2P1VMoM9Rsqu3Jk763o78rmFC7mmU9r+J3elo6oPDFNS9F7CudWglMma
/DHWVWHStzoK+odZ7NoYZpH/GrorSadg6cTSmEBhDwvM+orneb9nP6PSU8aR/9CNNSLWZ95y9hvI
60Fb6ldw7tiMp3LkGvxx3hGjBdd09DMSYhjS8PeG3he02OU98YEBgtDF6oT9R2npe5No64mjm4Zq
/8QC+1KT58kEQO2nDTze8oRuTsc1ro/YL1yss41w1dbYFjoyJ0nlEgEGPgoVW2LAaVStKO7KYTOa
imOX/e7d7YcAegOo4gGM/jIVskLRLBsAfX2TxJmlXmSnWf7BadTcjGmvkvIwezv22g7GpCdlDwsh
nVl5KJ7qSVxMj2kI57BmoBcgzeK6PT9vEJQVhBy+qlyY4uVjXBvlWpbV/I4mvDj+w1FgSS9khlza
UQZjNd5yvS0eQllGoNaYEuabdq0EozytmQjqlBXStTUgtBXL4jDOPJb9K5nc2SMnk4NZx5N3j/4r
V6uaVYw7bvP2FmpQd2sCEHTXQ8kDjxd9J3td/Vi8KETtrEY5cnRZiRJntFnK3VRfkUdgidGOMDZz
zBx/hiVUgv8f/zFOVcC8N8jK+w9JEEw4eBRNfV2n4b1wO5tBysnZC5S+260b08RAFI+dg/NY2rFP
alrd5CHSf3v3OoX7hqWSy/uZfdLA6FIBSfqNeF6uslOqMFWSUqhKrymPLL1TgXN/ntFod9fW58aV
PETyhCrKZTneBJYcGu7cOG3aC8Z/O74TF9urN0C4FvKWDMh+6KzwN0xTAakUqBDD62FYkQrv5Wz/
QIy6jivwHRa+cIUm1sY5Ww2IGOPP0Eg4e4v64tvUYQpG3S1XiHf2Sw1bbAeaYJ80ZKm0Jp6Ibge+
+47NWjGkp1fyc2oRnc080te5yLiMgtjAMpSMvkG0EXp+uScFWPaL2WY7eUfisRc2Zh6jY8Tutl5H
ibxrAFQ8vgFl9oK4At+3rF4geZvF9ybX8diZnzRlASvYJS2pd2zDWzIqcLYSViSSAgguTAbKda63
o9JbXaZlI4eoNHDQ9k3cW7RBVTIXHP+Muxi6bMJNsYICZr2zplID6RifS2/NEfvXQfa8l+xZ/vCv
mlTpbpTqdwpSqX7kvSOwczzULEFCJgcpht5AC5HcSgDYcVCrntheJtWvY8ePFK2IkYT0izgS2rEL
YBcuCGXbtsKm68tgqD7eP8rwq/8N1dH6DoNwy7hc2py4j2KPu8kee+mCEgL9TSvU6snOjg+Q9fy9
VKQ9L1CHF9Kw0F5cnOky5svN84MQ29Jp/O3Jb5Aed8ilNXbsMj3ZYrejQkjjofuGPuLtUkPCYQg1
27hlUlSFM9bFod+kD5U0Xi8zDRMok/jX/iz6O+d7cFNLnnmlAABBd0Rp8kYg37whdBxuvBxwRzFk
M2xw09kCreY7f4nG2wNdmuGDlT9OC4YWU46eWTiC1gjX4PDO8Ey4Ekmf/mLQ5n+VlKISRi5D/L7R
XA4K0RLJK0rQB8kk/gFRpm+LOeLKpZny0Kl/nqHdik9/lPBftqJD7ZKJMI7JwMtfFofPNS0rtV13
m7NvfvgL15PUchhFL5GueRlc4yHkOG5PjnN8+Wv3unTLlGR0zd/A+cCDocSP7a7KxHp6I4fcEGeN
AK3Pe0So8HfQ+/UuwUXPq6KO5NL5Py4+fI+QtMzy8az5lQSAlgubw+I3dpSxnRhgyp8qqb8OKiw0
1TISOTN4g46T/HCnuQQBudBuB42j7uycWMcbvkAR33tf2wcqS8OTD5HzQlegsVcxTYOaZatqzp8Z
w0DIVlZ0QtkPkM1/aICLsYTOuP6CqzTeOcPVAEbsAVAgt2C3+o+/QOe2XhFuWtyrn49C2FtZ28yE
svibr7aE8LM8o4gAjZmie1fGy326BXpboPTl3c3ZFuU7iMw/NHY5YA5sceHOMY++hfpYcVnX3AXS
2Q9D1HegMGypAXx8gsiF0ksl6qnPsXeUrxTWYYVzajNQGQNkVLuwwQnlPlEttn6YcXExDUTOSEAV
yk5VldoT3IZM6J36Qc6OJjy7Hslvu5Tt0a9c+J31R3l6PbERagWRo0NjhdI3D4cz0lUnMoP2f9V5
a+IUhWXcmO+gtiIS61SzovDkSfV1U05E22zNXQf/+o7QhH/Ofk334PqB2NXSBCBn4Lgm/zAS5dHi
+HIKqMRvKDE4KpgOiNshMisIK/u20ZbxpMJ+bwRD+9WoHg3davafxljVJDewPblq1zm1kHJvW4MI
jZAbvK8zlEwzI8Y8Aprh9U1haiKR73BMc04ZHb51VF8KTe4w0/VOM3O09DjTfpdzC8N4d5xIDz48
rEL/baRAJ2Tt08s3zC5ah4BOXIpLoxcL0jp/u75dGsnwgeCJKXeKBBbMdvaYDXBbbkW65G1krtiJ
ibH4RaW1/4S+mo0+yzjUuktklohQ0QAr43keRQ2Owc/NtVh1XMdVwTTMgnafOMeoE/s/BR6vmfWD
9WGYK+pf1PNL5g24ZsgsmJ4RQs2Cqi1DiN/wWpJOIKm+m70YtneXsk3Br2Fz2ud4hpzzFlftA4xc
OAjOb8JM12bdsMI30gRXtNFMZ9VO09X2IdAZyux4BvVQNdN4+gUg8SRMlGLFa91dtlG2Gu6s0e9i
QIm/cp+6Fng2udD2wVC9TTp3zfuY6fh/pLRGg8ui9Z+tkcUCi4GwTwsNRgnS1egxhX4se5Onz0td
+PJkCdXHDaogwW2eyXXt2iJmGlhLstSb0WPfi6wU+YYSjOgTO99SxFRRFg3oq9LncoTzSUYJxb+O
OCcukowBKQssP/P9djV5k2iPZPUJZGLdgJ0Hgraff1otEcnSeVgKHghbwsU0ArOyFcVzWEWtlbj7
z7PFCGikmjdCTYdrAhdbrYBGxttduFEs85+XI2lPQL970+3eSxjaZtQnRS0P38mc36IVDbJVySK9
rPfGdj5dxemk6GhgIxD7lyNI/0VKgVHqGwXKByD1pkNdogVXHZo90SEYdgUdpbNznqS+0fqzNy/u
TYwJritOPzMRTCng2xaaaObboEHoQm6VSK5dRGt0ciqLjIk3AndfB+T4D/Vi/uVxvWiRwLAHuMO2
1UFILwE2XFr2N6QQyVrUGnEk/qqkeBzcH88673EtYodTjqYZaBIDrI3ianRdhhfqBgHo4RAvPpHl
ULq8dwcg9I7EX8ViksbltVwTkEzY+ymNQ51d8ye+F9lAQcEtPJrnT1EQUuYX8qY+z4EBvflJDlBo
gDTpHs4nmyKpjbIRsC85wG6/gpTloK5xs6AodHBQne8QRJBsx4qrRZSVtPLknJLCBBeIQY1qcYWt
kzM/dLOTXehon8yehMj2WRWJcncEk6x0z5NvztVQskNyc66ZOBEkaabEXuhPjxc3nwpQQYBvBG0M
iclUdcQdetObeP3WVgKUqRKoHT9IP7VlfJ3Ao+6iRJ5OM/b4UBKM2Qt3Cy8xNIH+7ffBvTjbDlxs
4Jo+uxZP3z8JIMdQiVfVA4JmhJlJEhajn8X1pmE7hq1Ki0NQDp/8Vt5hTiVbrlAglh+fCn5ReUoa
BA/hS0MSNfQcnJtA68FPMy1vZFmgF2xPEuJQLWjuvNOAWtrt5LUSN3EfiyJFfGQ7nPqVtgHbshW/
XiTuYLcNnlY4RVazr4omBiIdzEw71OjQrL19hX+p/RqwMBPmTXd+RWRf+Jh50e47csxcP92WSTtd
WDT9IkBFnGYQep/eR6kycOMMPcsscYaRzMG4ckPjfAGGS3ePR35Iwx6dgJyyewzE/I3/T6fXC65Z
AKh6z+B4f6BUgLWfv0WYkSWltEEhsYSUnkkxjuJJWMYPI03hvsNCRM20ns5vBL9XrE7TqsWKsxPe
5J/Fzmie8DYTF+mcBho9juDui2tywdE32HXjw0oIF3C/JIzpCUtmjTwGTTcp6B2E2Vjf0uaisyty
uE4rW3ZSFBQr1+Id3vVT2ZDWT0S1fEJLHlAdoN38RZNysjrGOPpiGzTtvNjxnH+RQWXz51RhatOG
n7SdnUrsT5ATzmiN0rGDQcae5nsxmq7qBbQpJhYQJsDpTTqz8ErLZH3QX6rbdc1OPHFBAMc6c6yU
lQ8a1ZU4TM9SKntWKD0uARTD2f98sYKALfEBT89JcQ7BAx7bw82d3xgxu3RC5DvTd2T+vDQsU070
wq/EFUrIjYb61xI6UaWEQ7WaUu5o3OdPpBXcwfBaJZ+H0YGibK41T7ASgAOCjl0DaS96DmfjVwzO
g67mLDL9QXjPfhzw5RFzAwkvhGMyBSLzHBvmHIb3RIIm+d3VuiYCyEycMLGwFnqdVCuqR1C7yiH/
p8C9QUp/HfULhivlmfLOf3w92HPbb6g1nQimzSp/K9S3AmcTtudO9tCM+L3I7ZauCIbWh5FtW2Pl
Bfj3fDFtoyFNF9sbf1c9p6ozRne5V6anbdfKL/f4EHLqhnKwIZfsZiUW7Y2wSQM20EGfS+rbfpbZ
0aHpzh5bhN1G0jiUP45ogTaAkNW2BSKUF6EUZpjELhXF+p5hAJGZbXKRTimwaisaNEwZfn3TXm13
O4YyLCxjx4j3Xvfg8crDaXemn6x2jVYffxvqkDa4Ir89m9ALYalzOKYxVYAyKfWTicPrfEojf226
tPpGpt3wIi+dio097b5zVtDIU17eCobYtd29+SNEGfehtnRa2RNXVdibDokBhjIip6L842wqSAJh
io6nqPlvAzQeiQO2/MzWMRbhwLCagtkrvl/KfI8xttqVgm63wXFCsk8RardrR+Aw96E5GcbIQPLw
FI9LB+2GXQX01HhcEfB8FWG6pD/sao9sWdyeXhPExRNzQeRYvu7MLOTYYPPUMlbYClWnCtjLqYr1
LObAr5Hq5WykIgt/Tdu06Pdp3TelrqQ2HTE1m+FIzAoeukO044qlmcp9cbvO89zJqVe4E5fX3g7K
yC4k+qyvIo8L5ooZM1XPbCJORDQ1i6LTk/mfturf71OfRKDtoEfoDs2I5+MsQFRfasRs1LC34N9v
R9pp4mgPYA9Z52d/xd5lssYZWkSw4THTlyMbAuIK4+qJqiSIQ1caeJggSdVw23RFl3z7YkJs6ioz
lv0M25vwakqdlvtDnl3IORjOgcSJRKXSVrEpKIVdsL4Xnvslr202xs0NinEoEVLdOvIdO/lo6QA/
uycPDWkE1bWqytpN4/NePmMoT3NE3JaRgUfIooNBtZx5SV7sTvATEMSFkBeaAHKR9BrowLF0OqjM
jCiLVJQS5PwXC1FHV5rreX0kH1KAcaX6GJR0Q77qm89oqunJ+A7w6ZHxbNeiSfpO8X/1Cy36G7Pm
C2Fwr11S2y6TpzRzhvNciLj6Sh/9J+cQLa+G2z0sd+nxv3zoLU4M/ylg9nLMfpaXFfZeKM2MdaCv
fGb7yd40+bzaBnlTgA6WkqJ4MtlfZUJJKnDk/HkYdjEHcxGtpBnEgXjMc7DiqQzmdv0BtOSGWSPO
iC4uB5j0ELfRCRiWmCiCMDSf5eMxAyTspho/K4V4yGfgixosJPQnCu9AGQlbQq8pE5IoU5PWUYvs
a2rDob+x05wKUhhT5wU9SuLQ1NwlSyayyMBbkWScUFYoz7MDyphWQawIgah1YprUE5fXxh/vJq6y
Qe7jsbqKXtZUq/9gjLE2m4/4ozrYvrfrLDcNmMUrp8eUNlMi+IAkQT8a0SAyO8aA8XJhokyOblCA
RWmOcQSNoIpBTcGIoCUUxIZy+8lmqwRVc/LRWwHt9XBAmxSGwtBSujqQngEDtesFJNNE/CpM7Wfa
onlHjJNHuqxa69+KU91HXZ2uXGW1iWQ6xKMTVpC+dIE80qDXnFLoeqqomskx3TUy80bEwdE3oNxi
V3a0/hepiqabP5RVoqRFMpvenLBDYNhePV/kywHUkjadygdG4Hg35LrGwRhRwkO9wimkwm3d7IQF
8w9SPVSsEj73usnp4d89yLNvb0UCnoWLj7P0Na3ZACg1PrzFZTAlpFvng589HOOIkZU8HbZ6RxcN
sRVfyT3xocu/x6t1f7tL+MV3tXpgXfjcB7wxw8Ge5gbw8UcbsNCfy7wm10rYl57KziDCJILKWitJ
0QWBtGp0cwgho9h8JvWVASp6qrG0FFAk6YPLp46pDHeFoK4KNA45uC8skcHz7Q7CB28IccdQV/IC
xtT7q6mGOiHt7XHQmhY08I+kqD9wE3elnkQJQCpC7b9zvU059oH9bJlVvnMBwI//Tq8GZq/fvgWx
ivPZeSW3oiYnetAj4hGF3U4avEOi4P0SyhKP59tXOBOsqsfXkq136Q6baq85HRcqgJhzdj/gZyyv
hiLOzTOhQzuATrq4Omi1O9HyMRpapYINFY/lt26Mr5lWEh2LJu67z2+GI08n+VgOm+79snM6vKR9
PIYTiaUqqBVsKLH1ZR/F0KSTRqZJ8Ik+8KJL0V4JnrsfvHgGfr8fJLtZOL9by7Aqq/cbVzq37SFd
9ViooUXa84Thr1CrMsRWFWzWB3XkeX6SFu+ho0yu3zyM4gW6EO52r7LkSglNI9cxCB8ozFpz+jpV
iWrnHUqw59xIcdyla6H6qkkofZCmRUnWTI3Ho0vFtuXu+nnu9VdKdveunwPoQlt/Zhp+TK48UKtc
ZcFiDwjhvU91cfqmba6qS5bXG0El70dDTonZiTePu/VBNWBQijU9D6U/Mp7g/iQTMNfpk8VY8q4t
AKuG7IzmNEX82sDwH4nFdcxIqZhK9Oe62GgaJY1diADLESd0lJzY0iaE+bWLshElPk+Uguw0IP6E
6qQG1qtif45ONdemkcYP4NwcRddZzk6J3fNHAyWsoJNfAasR/jP8u/Y1IneclFZ4KFFkX6XkHhVm
pEZioljlaUgLnaAZeyhZwMwTqZFpZdbQv7Z9P0Te5ysy9NIU+Y9R1ZLtcvSKiHekOE38OLzmN6kF
jo7Ynj5nF7wRSq4L9dqo4YnTqW2XKfdgGMPiy/Wd07JfWdn1ck4M1xJuJRzZFJ8rogi3XKEdPsLQ
ZDO4CKEQ6rcCf6v0XA6Zcy3hSqYn2cQ4w3uBIUVUdbRm/vX4Xa9+Y47663SyVFZcCQeGZQUOQgJD
rhNpuQWFbOeohhAQWmVy4p8Yu+ZB47qMd41L7By+CpPyXLa+xNHzQeJNw5kpy6uOWrkLbuAz5Xla
j7+XIsBGMgLokW/AU2Ytol/PP0iAK75uTAn9sCy3Hysuc8yPfp+DnJFty7ZmJn/+SkLPXaQvnytD
zwaJFHMBa8+o8FhdhWfNfRUVbcDHO241fGeNzKAGxj/Pdw8ot6I51jYLtclbXSh/Noo45TMsJ7Wi
eMuGiw3pBaGJBhT6s3x0ZxTTzQKzkLVTBt/Rycs+yE6zo7vlVMN1h6gkAnhs2046VTm4ZijMPljb
a2L1JaLqSqQloaonBmafxh8t6OZCO4XbOB/lWZin+/WdJRR+hZoOH7jDDyXo23cyNTGakAkfPlxD
REl4TOHT0770EyOohIb3XYT7TM5ExdmXxUgGmy1ZDxzGovz8+TQdEWpzNUX5N5gkr2GBqrns5ipf
2OmjrER7N4PB83dW6hFCd4zZh0cP4y2cQFk1mfA922IRPehN2Bncjnscpwn0vLPWHHMRsM6XdG2i
GPewQYaCVQQYAQXo8qibAuXk5jk25VrqP9PynCR8h1jOh4AsnSxTXksjUMrKKVSOQeajLaWiMSUY
EEvJdwW+tscD9BKCZPgASPV2GtO+dgMvXd+rRkpiGqgYWmKgcjV0//mF3RYLz7Yoooe+nDcrZLII
OJuK6OS7dYfnKjIaFLhr4uixjU04mw1EyUNGUPgNq4Unx6d2NgFzmAjfJu3gH1a7KxgaCf1mKKLe
iCHMGDbZXEX3RxBfBjJuiag6i31+6pCZB/5ITQVCebMAeBgNuHbCV5pqBdXHkuIQdrXVLlZZe7w/
qjNYGTq7cIHlgbH/n/WPLxWlATWPmbqBg0qNlDW5ut0b6pOAW/Ws21ymNkIN5F7NhAKNkgLfnZQF
Fhqa0+QjYAZvUSi92sPdtjsXh0LAP2oYA/a5JOq0T1Qjw7Wn3JaHSSO8hgzxY95bujOfJGr0iZVZ
bzPecNlWU+ATKCq/oGA/eoGZ/WdRHHVPOW2fGW1r7gWavk6jdQr3ZANpPA2Uh1B7YuLxZzh5kGcE
8AESbEVooJgot22Qb1dJ6z7NzNt5KZciDbG3kzNkfAkKY79ah9pHoNFw+OzviZ6l0EyKY0yBr1uo
A7r4qm03pz8+APXk1GNqLWcr7eFp9TYh62g21H7IQ0Q5u81PJbYJz6arkKJt1Ta3hrohtVcQo1xi
0a+rrZ48Sbg9k4V2/FiVCr4HOdlDU3ZIFYz2rubgTRUdxZo3Y2wXyvESfYSNPWSTdYj+/gRzIJou
+/09SYPs5Eu9GHvkiw+wEns+uUN343M2i4PB/rdUJAVPyztrKaRor7ns75JSrnsXyiy/t3du9Qiu
NH2/wkmV9xCc+erAxYnd+0tfjlrQ1Zh1B5/LHHnqFejJPqLGizmvY6L/hYd1L0AraZupqmMS3lKD
AzIvcPL9whrNc6D9V1CkG15wXZv1v5eOEX3SdBNxz0VrxiLHcSj+aItUE9mpcnsS2sUPpWYYl9AP
4B5tTHGB5H1Kz/KHxmBMZ+JPpYuzJgMnSj3D1COv5ntnVnz3CAOb3XQCMoovuHnmL6PlLBQR0erF
NuyjNE1gi3NXkT9PmD8QhHKKmKVo5TGfmiOue+f5XQOs1MaqdGF7vfJeqw5r3cTNhGQoq0c5DHTG
94LzyEiITnyIYbC3FdMYM/FcCJOQpkj8+7gK7ZPXKBL+5RAaLoeIYvnhbg+EmjxX1xQ2zY8DviSU
4MxKsGiYxD6XSeWhvh7/4utmG5j5cfQ0gmTD40s5m9InXqYdnmRBnkWyseeOknGGunO91Db3K1xs
yA5F5uyl8n3XfIjJyWve/kqLdCfYLrcMWGUEXsS1dEodWmYRUxGtXQ3xak2syjxqSJkYyGE9pNBT
Ta3QDDKKRRFYssse9heSo7NT/lY01UCgT0bfTeNDEx9+IMTa2KMit5Qv7ICc6Sh/h+Wo7LzxzPI0
JddJa8uAY7czW9wwKfDYKiJjQf2y0X1odLGtxjBTAHVxKq99YA2TrBdpqfQVqeic8lwMlupR2SVy
ahLROlSO+SBbS0GpGDblwWrrGsYsT8aFllNZ6050IJZ6EO7dH7HYcj/w6NIaZxsunNsNPsBbJzX1
VTsMJRvsMk5oSBgPtJ6hIs6DzVycHgJLc2N7zA0vdSkvbBy16xvBwD98q0D5Tz69314/0PgTHxiU
qEyhSRzRGZ3WEWKDDzhquiRxZ6nJ5gHEmWmktg9j6Szcf7Bts9+40DWCUB5T/e7m93/SzBnrvToc
IzQ3yfzm107aTodWqPYJpDG64lF6vFSTNMPCoSP35gT6x+4YCgP7IlRH8BJ6//V+v/J0LWioqFFI
G86ie6b8PogdezVquDOyB2x4R+2IIQ0Ne1sLNOY1+8QFkz34ENyO9DSqWTZHtP26DYh2RUFRYhCA
fmlTdApEJeWb3hjw6q3qPLz8s2Cf80GFnK+ETRNnuppsgbFpuC1mDzU3jzJ+Kjpft81Cn5J9U3xQ
tjcDQLhLSCdKB+42bOQLCcCMTE6IwNVhmaZkKWoTmLEPa+v7P4eS33K+1PrfMIGNjX/mACvqyZU9
sW5OrLvDTIRkyNgC8z9RVPt24/OWPfmPP/DQlfRMOEwc4HKH6m2C20iEQvy4FrcEBxhI9Esou9sT
BlDWDoPbaJRITEiTb1vtOzNtFCZI0RSKY0+9jr5wxQ3mLeB7v/c8NWXWDDA8pFDYdt65mFfprW01
rAfZ+XydbGkpMjFqB022AP6p9oPgTPLkuUvFylmHpyUop5tTDX8IWW/J01buee66rrN0uiBSlgxA
h7Bv/A/Oy00VjxnB3FR/qpbp71ufexjck9MXMCNQ7jViAxodU2DFmnW3Ra7IhQ+RGbVtuXMP4xYO
lJPFi7hDJ0Zm2o8lxXqYxzZFvek2kQ+SHZooqhs/oENpGvO6H15lQGkBBe61k7CU6qT6qzplEekb
q0o6DFpZIMFK6zshNp/jEHsbNKq5ibZMxcg/AgJ6IoIh6SHngumXAEXPm8Ydjuki4NW+FOUe/2Ss
qJKYkCmtl7SMPS5toLst/wqUNxHxTWU3WBIoXWJONVY8+1xdIFU48MOEcqFFQD6OQ29zAFC0eiqN
whQTUGh/auDtgWbAtyDRSKCTVjObsprThMn/ErpIarJXaYzMCD3vezObvkQAP3U7D8WDH8l3UgLR
VXXfrqZztZYZfzyQDrCYgmeZ8O3Po7gvO5pLYH0wBqRnBfLZIminn8YYvAvk2gMjzaw0toqM2qjl
q17MaXB5A7MTqFnbLpLGkt/H+4s3a3uc4HQN+Wul/efZvelS/P1kt1spki/jOvT6wRHbtd3Vqr4H
paBDdGkN5x68c/XIs4NDFmu2jYq7Ikx9V40QUG9+SKojNrilPVc80N1mLmJyrkTFQqqCOgAVi8w8
S55UE8W6+6ae/jULTruzfBVuteMmiGNzv8Y0Inx5aVEiXWcOxxlXf4i0WM1w22+2px7gbpKgjUPe
geeKr6dmZQ9xJZQTTSnbByzyFgZU3jU8VHNeoRb6VuW90rd8AS2NrJ0Sb6n+rOBwarZhJtUJa2OY
80P3zbsRs31em9fuKBel9m4QElCJ4KnTWmO+/SxmvNlcqDxaw9uwdT7CdQCPkVF18RwNtcLoG4eF
fbZGDHYgvtgWeA3fo6xRa2Ffo9/dD3l56Esvl36mMkl87spn/7sowRHZq0rmhy+h4ykcIDzeiLbf
wFhf1lLo2d/2fco2OXUtQrAjlP//EtqdeK+iiYXER1jgY7S7//bfK4VhRmgYq13VYpGllx3tUsHp
GFllSe7zn9s1JQfzdylktA/QDXBj2ZjQSmYehNAK8suLYbCUQqvaFfapTcL58Pt30Dc0vdhJkGWN
Z12Cdp4qfa0yqqK7PXUKW8u9sufhftZMYaXlFj5iWRvF3wkcT9bUSrbQb8ET/N6iCXofOKTpHOCc
pza6OwDr2UEWm0hSvKSwWRfGxZEvrZOlwCmc3NLKNivk4D7rr3f4EPcVrfkj0R5mPMby4+5YfqGn
GJscNaPwLHnPyhXMBSbzDLkSCwM8ghJNUe9SNV3mnfllysR+kDRaWazeTFYhzOjmBkKTe+ppylgQ
UkcPbI0svjvZpT7K27wQwsSpWlrkohC1vLkVopmm+SB4RsIJnxHk/6XqzAr32R1iS8i2B8ftJkRp
ICbZ4us40bs6FtgWiPDm8aocOoA96paFKJ6yNNxVf1NdK9zsAXQ47U5so6/bzHbm1g3UpXoWdjIh
S4X98tRN+TipUcoocJVo9hw1iSCfIQm0tIT49oLTL7AvwK3pkTjsOK/EY9VgEmyjY9wFKmrRZqwi
QQ0m+VBMuyhvNKamL+f0LH6SQ+hObiCpFV2Q8yf/c3ddttkoadJfzoEFjbYjsncU33T8+FKiPGeg
CilcaUEq7qTIUPXFb83mahoYEFbyXMCtOyNWdGBnTlHFz5ZJ+fgytGtNM5NaSIK6Hfc9kVvznM9/
L0YbXaPO8TVKspA+0VoQP0wxGxqOM/WNzMCycVlimlKIfRyyrbGuSwaB8o0WvArGookaCCNiYGDx
4tk/Vcd9h3m+izJuhnFaehbBqz8g+KOui12U+rOvwYxq/weB1qwEXOqhYtHpR5EtUI1HfqPwjgA5
8/z4kiBHnTqHpL1anL49FfEAHiEVGgETgVckE3D723amrA+iy+jG0AXtIf0it1iEHw30N4iUQrCP
ssJMG+1ETig78NL9x5vZVGWbunMYgbsjx2+chQj7P1wYJimajByXPMMUNLLOUtmKKTR01cwzKkNl
zW2X05xhL00JyRUeAZP1C7S+6Bn8dXnUCIR9W7xh5ETeNulgKw6K0kjrkG2wAytH6eJGd8CwFq0V
znBKFs768lC7wpy74tBNiqfw3Z6DXq0hAd3JM8qUl9bDJeHrfAJYS7zdqDSmRy1vOpn4k57M+5Ib
97k+GRxZP+JJviNsu9LaE5pg1bIWxgdq7wSJZsh83+6yoDKWv5l2TVMO2DshfyznDBiksUGmLCcD
nlvUS6BTH8Uz4k+lK+aseyYmV5bTkSXGa9OlCFeNB55sKjHLDHezoFrDkc9eaeIGF7mBko4wYzaT
jVQEoRKnuNpdSoqH3rwBayTK8DdDFB2V4w7tiAd6+daQXlTlgqbyS6ssTIa8rh0jgS3MqCPDbr/K
Xvlmp8kDNK64lYDgDv+ywuRj1axdpBdbPxzmdmtV0tpfaxF7nYwruuK9y8wmuYnuy9HK0wLrkonp
RmLgoo/L75kvyRUdlngABd5dBS95Gu8H0RF9Ej+ESmI+XOaNR6LeL96VfZUT3EOZopRyeVAeDn+B
tXT33HJ/hH9VLI26NB5QyO/d9FeDold1vCi/bJBXU+sVHpRFTEar7YiI293cOpqpauRYWcfsnrg5
zYquy9FkMmp4Kx+tTDz+XUdz/7RKIm46ETwuF9lGq+fdSkQrjx1jlcQx9qyjZ6wy/2wYYZG/1VCq
RD4GFxQHftGUuIph277/8OEJeJKDv37iQPzyZaEyXHi26fu9IN0fLadz74GSwXU6ssE/le6LP24t
d+ysH5MMfudLh8b8u1YeK61nDFksJ11GWa83ZVLAQUcLUCaA6MpG5sAOdx49/qpeN7oU5fR3qQ+J
Cm3RA7jR3bx1Gbaly3kxoBpaCpVh0x8bdm+9iZZba1YqiEFrADOEqYZydxhOxMZRNzNLZpsj/4Rj
pr86a7D2/dWC+GFxemjy50H+1HjiEmDEYuCcMs8xas7TIKOIRLQMsifAtqE2KgINAfIPX1BqufJ4
ruao0krXRve3yAlWw2PPeMzXdeWVjv+Wc2NmXiCIITvFUbGJ1hv2A6CYNTvliCSB9IvMGF6xv0Sf
+GgM5pHvmxCjnSM/hbUczjzN8XsMX6/e6c8oyQGYgTiUbEJ5PB5LuWAjCetV+Ojqp6e/L8ijnh8r
RMqTLUwXP5u7zVkVYKVbn3YXawwyiRQwZeNiuIzpkF6BPq6vIIEm9xlaiouvb6sy0OIQ1odkIyCz
xa9i9ox8RGXE/ctBVq1HIVToH9XbJZuAmhiv5dK/xVE2AT9+p8H6TzDNrJ1sAg/MUFAevK6c2o7i
ySdlbj68q7q2P3UDblP5yAjQ+clw9Oc3HT8cIUfHv9beMz8DCiwTkAyTiZDr0vVK2WLw3XXFYZit
BFQGMYf0h/+HmfR8rTnAZM46rCxA+JqZx8iurVVUkHutnpp5gwJjXcmy/J9mwZlGq27+sh+HAKt8
8m8hDhRCG0e0OvsoIngeV03UxYEaKkVHyFpjhFdoZDiSUa6ps2JbaY3Tn9Tr//r2jmTR3UXyOOUG
Alunyh83zmDpKNfUXgJdOQhecCGW7DuL9sSQMM5+Bss3D2spFunwA+C6gkF/2Yf26kZQ8JEioCAq
b1Aox/kAMriF+HEfMBidFDLMmh7HzZ8x3EGS6UaUbD2naeFpkAeFZziULWBsuVQJHymmA4X5d53o
85OinS2lfbA1eXB5vrZbjfd6v5EaTBDsfv/7fgyUB+CDIniTj526gVJObApNvGO1RKnxhHt5BiHs
lvlCFd2sB2lysMLkle2ql73nFgK4Ny1FbB2SMFFcpMmqXjf0u0/3th8rkY3ydTA46Cd7YSYgbWjP
DofXOu+3zx8bXm9vIsC8JpO3HoWtS74KPndDNZEeLpGbBcqdzCofstnIjrUo0BvDD0hAKIWCb7MR
OpZW+UoWYjqtwyxwQB+3B8SW/ZnK0L07UXqgtFbLzbuc3F/Y7p0jM/FyADXcRB8qjMqZIP5soQrS
3AnQ/rmgg9Wjc/u6Ek70wNy6+O39+DEQPkJ5Oi/zVigs2D4rpFoj/2ZKe6iybxElrukKeYAC8Qna
k/efIFVoU0zsAzY3+gXLuNP5KDH9XUOypidOlOSdtdiH8oYoiW3d747AOXxRPsb0wG9hHTkpbTNU
/tZeeazTAdq+VDiYzekGx4IgZzDhALik+I9RICVqmUlbzxLDrNTrRc70asTEIkL1RilD7tK2C4Y8
Rl0G31XL7kE8saRO2nmB7UQsqTaGvGgIRBn9WSTMvp37dWYO5Tk+FKumLpPchF4YeN4EGkVCGH3s
5meemq7QRfbBBi9uShYQDMpHJNii2I/CzXJ9EzhJDpylyZfyWnySFpf4gOhZ8N4e/EVyi83gLu+/
Nd7qAFjyD2QCsP1zIiipwciHNwMTuzTdPkEVWPSOwF8vI/kFThyoSMunnMLrN+RZE02q6Rtodiuq
7L4fzrQchM6EGQOFt/CDtM98mJEzg7KEFxgiSgpdWsuIBAFevZkb2TU+bWf9Adswknuwac1VUMvt
f53XXXP5dwUPsl+A3tRuqv0bRpNbraFia6FrpVgiTLs2VgK7FlMH2i/O4zYrNMc4aSXSinm3KXnV
z1vAzmvzLGfPFuti8lrgSxaSACUasBEa+ULadGShAaeTbnh4JV2/WBkgviakaN/kf3T4BNwiXU5+
sI+YJfoKDvQbIGDmFh2HvXuar7L0o1I0goZTNC+1KeKSyh7P2m5jwC2m/5BO11uOJc/xecxF/5fG
kZ6vYn1tAHJ0772ZgAB3oiE2SsOMRfePVqBSn+iCiZcDoVQ8exG2aFNPiDHRTMT69FYq1m/l7Mjc
LawYdgDRumK6yxj877Gvtm5covcOw+4o6WxyZbDUQILOtWsrfeEE/XOqUeK5RPO07xoOrRiFEeXv
+gZQUoqLteNqbmu3xn0zj/zPj/OLwS4Slf98pVSWECzPPYmG8sKnnA6Ty8exbfSgtv1tRrIbi+k/
GGIRA6QScodMIeV8CAJugoqhY8bX4Gw1W4NvwdOAUwnlZPwoaAcpjQ8Rj5xeuNFY73CTLSDp8x+b
r+ox0U6s568FM7AnIGvvWt/JtZKnJgU/RBFR72rcRjv4MspWw36+0DA8epWgot/6U1Y+cZe/2nUO
HZmA1DKUtLqHG5A2FI/0q3OlNmXL+8/G9sBGg57psE3LBCjFlfN0ZiJk9hUFgccN69qzZKaW072z
G7BtrDw33aYs7eiqmh1QiKTh9GvgTG/2gRkAsqgqchmsRO/MU3bsMBdJc3WyR8/fa9I2JLMlE5kY
DfiJykn1DA83jaTKggP2oQSutr5fA+gjJbPw2m7Bo2RhFeXAHzxDTyukFdVmrzLyY5OMlWejwYta
ISGklY7f8UWwvUhx2iBIihUbvdVg/UvpSkqhQusxkal8vgUpcC5/qPY4CteaiAmJMuET59xRBDoU
L+zjmmxPYWv1A8TAC5bQJ+j+djBoVjxputh59WoqsOamjDLPCaZfmCqVtHwgOWjdYgSR212Tbxrq
ji203yDNB3AarkRtmRgC380PGvh6vtSsgiNxpsR+rUZh3wXBwSU/OLDXkwCUtLqvC4T3CNBp4gle
j7rAqLW+aV1C3wbEDu8olalqunCegAfpmP8xbrvuA+j+i/0/6aa8Wl4lPmkVEw5OeWWeXlv0E0PP
giEmPLQ2H5rEH7DM/r5DoUGiI8JBRo6dw6JoieeL8o7OlwD0C8fHir25T+BVil6hHqv3CyQyLcJl
Qn4l8l2GROLWng7v1CFOGD/B0jMkw7o6t/HaqXFihQ9rYzYJSX0QfQ54gsKJ83joVyiEJaF3KAj4
RBAcIpZit3DG5GH5+zedk2o4udXQRXDUghFiI0ep/Bn6Z/b0/++xX7sW4zG3HSjTtPKKvH9le/Ga
6ZjvEAfMV6UD39ZZidbjdRMjJKwP+qcTIXYKM6/yuvj++t1DN8GSH780KQ90oQ7kaoAcZGqOGqiT
vJw6kcRDB0CeXS1G7TQBLj6QsabHNjqKOxoDOw/K/Z2n2g4npopfXMpJRur7jouTu858FsNud0Tq
GR99fqF6bZnFzl1T6XyYTKv5I7CO1qTudjT5ujK4pPtZemhqxx6D/hT1WWpgd7zxoSjUdlXGDgPC
qO/zVBNV69Mti/RaYThXsGBvd9Svnx0Fyj+43VAVUvPuYeGNBLUyuuezHkIutYkTZ6xfNh8WO+DK
rjR1L27kCpRS53ZQpuChUMaY/lMpDtPBZRw02pmVsUUL17jXbMAhy06jmGboSQjqajkOIRo3HmDp
IduuqLCB94JxJqblPmQP0sQgrhjOOJ0wOwsR2xIOF9Zq7oZut2sQWQpVHeMD17iJOTi8QHmURgcQ
kuGE6U/1rqdg/9dAK82/oXYfRA78byOJ51eOcYRpcCrFtoZeT6cFSemSBT/pnvS0IYoBExs3vRl/
HjifdBoLzM79Wlay7HDHEG8qsde/OHK0PfFwzP2R9LgYT34sJQM3Y7jQG/71kmYaY/J6ZgkPdS1P
MBZjcbBLjGha1pv06dHBu1aM4E0ni1zmsnuez3eP0Z9Mx0VtiQSnbjtpQoECxhpNmrG+9QgGzJOn
KnaW8HClNi+GQA7s0vWEd9sOwokdBbEDhYRmhEhqtHZGTvnfuUnf1Bnj174PBPfEcFOIVAF4Lgc5
JWZs+xUMnq5CvKbY60krk+720gX8afcNzdYknJ9n/DWCnpbQFQ/GjmoTXxDv4GC12ObZ9lwBWTac
p4HT58Jr28EA6gdO7JkV+RxNoQDZQLHFGJWg27r3UPtB1R8MH/HC0NbfEM3AY6dgOHfOT4VlgWFb
jb1kjUEQficOyi06Fgo0Rn8PWxxwXSK4OCgaeyyPhJaXauWXlzxYQADDWfxBQnuZC5nS53XSA+m6
5Yih+QOHoSjmyMrOYYVzJRkqO4Ilpn3QTbhPMz5AtKDNmOHLzovlFmC2xIBAq2dAVLLC4NOfC5s7
/kOU5RLiiaJ8MLjvNnyMRaYjWHI64CsRUp7K+TuqRAlelEGUnErATlt9dDx7vQYpUZCJ6qO/BON/
Jj5LBmNtBxSLRM4KZ7Sk1HJVYpo3vGDy+2f1RkrrB9mGSZiSctZA9/s6qNX8vVCFt+WJp4p975r8
MWzDb9KknKGqB9d3NABDUXGxYVA+M0vrPHIjtyKJtFmZxUK51F6Xkq9in3bFq8mH7UX4R7XvKtOx
oqVl69osPMHaCdopRaAnTtbo/g24kbQevY8j1jJsazj8CisL4j4s0mog946UGa7yezEg2aNSnH13
xqJhCx6Cwy3NzlvlNFvkbI+8vX3FYvnjnU1vyPz5/B+RTZ/OnNmECgkRD3WVoA3eB1Nvk/Gqcb4N
JeOCtLv5cJ9CqiFZr6rFiol9QC9QHdq9tD5L3dH06Jw17D0EZ73zyeW/bww/WpjpW7mFlt3kAQlb
sW5EWUrMwtKaG+F1F2UStbmP4wTThNR4caJbC1jhoFAFPO2OTcZHgQBsArwhnjPoxpvxyuJUHTIN
8r+hz135kxVXPk2Xrv/AhMQF7VsIUV8TPcNrw0KRv0wLjRpdghyegr9y3k5scRFXXPoG5IWWLPDi
5zYvceLIG11m3+/ASYsPO4I73coq0SIBLcCJT1Y4l6hWCton4esxzK1KgukkYJW9l58dtWS+aAMr
A5tNoga9JJ4XVJoJmTYw2+R5foZaxOxt9uvFKm7EwtaqvN7cYXUtRILUXM5NtZgrQTPjLEGYKuJX
KNgXgn390qtXCrgMCtI02XSjbmzbyZSYkAm9nNdVerm+BExjEoiKokSHPb0kuHISSQ1hjm8jw8B8
6x3L2S1JGfQd/XmoY8hvUcgcMw2lOvnpHj0sxE25QlCufBS8zf1fTr8XNe0AD8YazNVSUCHmaink
GyTebwQC1Dv898ZCtT8XA0sPpstqq8kE710geVmuQZHeKx4ieFV0tBcjKdcBM9/i9y8JQxfP2NC6
9ECY7dFjqdG6qX5imMo+HlXxjNtX35gFglQP858nCDlAYQ6lHjyZqQrMyAsWiQWFHHn9P3YoQI6Q
bSiZdanK+r0V4OlTHBAgWhj7ui7e41DEJXEeDleTw/VXka8/xEtESL0ZEISe9qs2H2jDJw9ye7MY
sWZmbaTcQJqjVIohiPY3PW0AqoeR6hIOMAycsy3sQ3MXwiZbm2eo8aOF3IDGDPs/wazpMHMFmsrU
Xhr6Hi+JQdcDi814Cw2vsMSri84qg5+JdZDAeYu71qbIKCbYXDJuiARbInYWpAFofev+AWtbZfIa
nKRXHkLd8J3E6hZIL2mv91iw2qDkAMW/hIO3tEITHE9yQ0hDziUi8GNdWTG3ycJVM9HWxlHagXth
sXj6sTEw2jy+IwmNQsYCV67BDPh6bIcrC7IXmEpTx3fLs576xYjyU7k9EtcZvvKLuy90XgZMTeLy
MINE6w+Z5NCKLUeivUEZpVWPZrV17UEpUiGo+rh7nqFUt2BU/bln7t6bpenlNXmVlzEXj5AkYBnH
jNnHsnLxtXVM4EVPTrGFLQLSAAoP9+kBjxROaAZPBWDSWuKXNswUBn7nxNQLGO2Dd3a1qTA04Exl
5M/Rk8P8X39AdIysqyRmG4Z3Rg/fQZn5vlwcWOPLoMYRw3LtA/PCNX7DuD/MWPjkhcrA09MjJVtX
xvNjLvjxYEB/xrfdUWsU+jb1N9U7QpauAUvefb/0NCnCd3Rpi9NVmJ4kDIg+EdB1gYY6P6cCRdhF
BfGrmhL8sY+M2ARhVH8S0GXeH3/V9+hYA/yN4wxdHLJG/SMpZwussFl36h/vwi6r+D5eSu5pZZnU
40mL/tFR51Jw5fIc4KSU0VTjWjqadNA32SsnXnYnKhpOJyNTmhptyiDCjB5WdA1adq9movxH1Vkg
w3hnT9eFyZ1r3rhQUQI3J0XfPIVgSZEO3B8E8SxQlPAFJEjcp3WibI73lg/jQ1JCLdQw2UKySRMr
Sj6G3wy1TgOC2VqnikFRljgIYiGS20A7OHPKwMIwmTkcyVaeH3l5raBdyu4wKm0IFGZ+sh/y2LJp
dVWh4RC41puqG9r8UcnLrOo2oJvIkmNHeeLsqb4QImoRU9KqJOBSMJGDQutRVbZYHDv3mSKVj+no
LSrNc4vyE6TbM94sudnCWX0j9vREuQQy87I14xqMmy4Dd/NNy7sFlQAlMaPsfGTJ71gcSzm1CV7f
l6C9iQ72BmkRUqN2pcPPuSD02se7si8jmqHsJAgTi3tssRetqQy2t/b70GqqHQiD7rjlum2VNR1p
QH5cQlVscDUDsCpIop+m9QWCS/Qs1vEXSHDYT5AFyibYpyv0gp03bTTo0sTEy7jhNFk3DYB4i/hS
xOye9auOT7NvLClt+0UkqrextpE5a+HOJgurYnOjpDdtDvJ3JYIUZljN7Rl/YHpclTinTrN5cAmD
lVQsF0jvyYAI+kD7CAQTUkWJh3Jripz2l85CRarlBfhCGDpqdwrOvtMITaJSoAHkYjwLll0dZ9cq
XaUp8oH2dr7RK7HfUCTNxMvTE6SArmIOPO493rlFsUDf9JrSY06Tlxu8AMEhFqsA0b0vtBEWDOud
Cx9mWKVvrbpiFu5yP3tvyUMytcrruRoRHT2DxjeP8yklf/HJXSKlxsjaIYdm4eT0cvaqyl9DKlb2
V6gncMXqfDz6ypc9tHfqVE+yHCniHEDSxeUI3jwgKD+n/kP1UNEXI0nW2yTJL1RqTuYV+3wgiO3c
Y5XU6RDglQechEeqWVbbrPFmMJ6GWGQdQrrao/kmAAnWJdZMd46FMu9rVjnubs98uoq41sOSYYlK
DQ/j4AfTj45eA/ERbKJEUIwp2yYdTnMCHoSlXb/3d1JRhb++Wi+pD2/4qn33ceGqLQlLx5qLL129
qQzIylT7mOo8kpihzlgpjcbxzoTurZILZN8Ub41IYdbPWDcReNj8SylZGqRYRa2CY9QlGF530d9D
ZSqzdUcsf5KcTyj8gCPpvxZdqeE/2VLnDDl6dgi/do4ybsjv+KKEUC5AGfkojfrx3QfhE+hO77Kc
or04O/SXFWECHKbita3ZuIW31B4XTM8SStnyuUvahEibBfu9s6B1okWhG7b5sr8z3pBOuK1lFtrD
pEm3XisxASBLyiISZQGukKG+DRF0gwOpxyfusNQU1GFSsQ3ylKlY/RcuHDqHTL3PxII07xtMJFTw
rayuChmj8+Bhgu5oUoOA19QbCHI6zA/qKahjIuG/Js11QO931yLCBQ45IJnTO5jXqwrx+vobcfx2
aUMbBAoSmpdNE7eBzEJ9a3jJ6EeAxw68lcNFTIikJH89ocuMKk6e9pAhjJ2bNDaJqxFFuw8qTZqD
7E6NLbSGxhaUjb6iD7Rk4BMMic8qqMig6sagUW5CZMMHR3rDZbfXWrDJwlvBOaFf/ThXluFxe1Em
2GvMoT2JkBuQft/QJV8gUha2uUysMm+8E+s+uhBKqe7i5bGUKkDoUAjYLMK5tD1dGeejI7xRxclw
s4cN2WA7BNd5AveViYP3DD+g9gGcq0EeNrGpxCLKb8RC1UzlTBTV+wpiOf42jYPghDljQ1nZLkCP
1kpZeZGWGZXW6pSulc+UVCLI3FbfKiatni8lf+6VDeeVZQUwoPjgP75OtJz22x4v9HyiB74jbMsB
1ezuXuoMtSnZSswU/QV0Gik6NALnkAJabEMxq3MV/zMe6s/05poPqxElvY8o0GUdFpDSA6GVavSC
qveHKz1RRQfGWroJ5JMsPUO1iYbTRFNvi1jgjTcolv18aBMXnNWjz7IxTBWN/Y0/hxdEyQCFqpgy
KoB0MGQSIzUrC4MIzNWb7eCGgUI8IV4C/NRgYuUk4y4dUuCGFHcb3jpZWi8Qd9wosQrkU2G1ZytH
JGRU0PuVVACscIgt4O4BFGIsKz+qX50aFDVrCnj2cZ2x7Fr+p75wdawHsUVVrqCkQQF1QrCDJLTw
i7H5wD5naZ64PzqGsyKlSjfqivVvNi4c3OvssTmD1w4WH1MlEVpvRatQN3gN/473dAjPi9B9rmlV
JU1LQFQQy416ZiNfGI5GixNdYtvPLFrgd88xLa5UmHvewztks3DoHb+sx4kRcVkAFp6qlmgLqhPH
AICkmrZI8aMEcauAJiCdyIa+xRyJcqwTdRRYe34PzD3S0Szhk4p1J/KpJ643tNknzIkZtqhWIE46
LIwsT4Mvdeo5HBzDxc9CunN1REDaA6rxICH8+Hwp8zrAKZKLxLakiwipdJX3ES4G00UxNRysidbd
nMMYDwQ/aN466jEPWn3+u9ttjrLmSMTbFA554+/tZx9/aY/LbrgvZl7qwQHYFWdWQvQ5Sz+MHPvv
TaPpWRf/YlRawCBuQAgtc7PXSavubImHBK+GJ870VG30UYiKeEJu1vRc/nRLg19D+t/R8E9aW/s0
ktN6Gwwj8PIXp2YfnME079Nc67qmr/xlVBxe28xL5HG/B+WEEyYqkub2HOPEbTHn2UY92MepXf74
sc2pPHKfIdSpFVsNioBmELK9DCy6UCGEQzhb47KOmq6wCD+F0jbMs+IdCkfNqEDmd+cKwshUDbvm
hau7fil+rVV4yYv83P24N+SWWBwY39DZg2BCs9N+b7OWlh7120LTAfn3TQ4NKGoNrcf9xhPSKHV1
HhJ9CHgDAQCnJFhwLmsiytUb68LNUm4Yekkv1GbM+XnOi1t4zvlYeF0t3JhLCuRei05fVPrCWKlc
qiV1k62/CyUg0pdH9L+Pigtk7Od9hqy7oUAQlQa0ytF8dvspSDnagZx7byiXAV7TtZA03n0PXiq4
dmbiX78iSbE47sEFuwf+X2iWIf4wIeDdQxaKP8cXvtJDNqmWja0L03qTr+ymViALx9wh8psQunmw
yl9S/0m+Aui7m0ZKJmf1uurClCh9qP5f8uj70/CUtBBwNXZhvPVtgYgiTqDetCdsIqxx8Zfesg4N
SKRGDYbcU1KYcIEKDV4l35dHQKjuLbvhegdaGXeiZnO7E4Btf3E7cLPoZQMFz3JE8a9Q//hJWJvx
ZuZFihxheSgWya8LRQd4rDl/pVhd7CznhDE4O/Iz3ldqjG8bWjYlgLQXYYZvBksPD98ptvhUro/b
gt98l1WAjZZuBSA5JSrZx7Xu/0ALGczDhTNgN4tZar3hgINB4wJvibibYYLR9sXD6lzfLRDUwXMB
WZ4fGsgSy2BSbopLGHUeI/ZDvbUWZpn4xZCEZwRcTpI0ZjxJVm+YuSGDOsSyFVXjnXrmQ2Qg8Pxw
TW9UhmFy4rwHtXEkMoeBhVfWQHey6oT9y05HURECrlvgqwCmWNbiJoSHpJh0KcdEYV0IHYBbTuxB
KopIAvnqxtzzBVqr0YO6enFqHllXm0Hy3OliQLKtrbwNwmMk0KYukq/RMq4e33cNpmcp/tBSdClp
gCXRH21wltHPr1G1EFLO0XpO+OyVguIpAO8DJAGQLUHszTjKQgjX0VzGZNYjkktNx8QM6nYwPTjK
5ZTHpI7RjVttSNQ6PwbcnFTTwLjYfvkILDAeBI+U5JQUJXjAydaSYXWmZ/kAP4FtnN6KgEGZe6i0
o1Rh3mm9ZXHUyvNyrxG60T9SY33mwRqM7JjTReFxfs/B2GEsecOYwZsGVkigzVzGCIHRoUV/ZMXE
rYWcPxV3Q+7bkg+Mz2isp4NuKQpkkEZ/kd/LQOebHjudKO/w8M/qsKmCVsHzTHpwEaCuPNurTEdE
P10tr2uM2a88qcw6GPTAM+U/O5HaCNRjYeuT8I801I9reA1/vEmzDy8D1Bv45Y06eG6PBrB9QIOD
dHbD2flvofKn9liM9aL+j1rfsPdF7Qfz4dEXd2NiW3CdbV/f/55cLPyXfkQpy0Id+a0ZQ14TLAGz
eY2IxA7hFMhUiZb7ua9KS4v6AIl5Cm7HiSfC/BtGqBwu2W1a5Xk9jmDR4yiapLOqOPdGnFFwF1GY
F9X/ugirsAY5bTEfYswOAro8goWa4JGc8x4ODBBNSdAK9dM0c+h7XLsPk90FbInklNrYiBtIZOWV
GuLZgLUkk4GOyZ8bn+JvwReEqI1ET+CKuKcLuCMlfdUDu53/iCdrnkHzQ/3k74ZS2jH3RBzARbf/
6sQPbrd7n1tz22aAKPuXTRM3OT2g5IC16KuIBk0DuWhsp93hto8x++YI9B7uN3iEtQqDlYb6XVzC
n4xTu4FXk7xphd9aGP3rAoUwt6DPJMaXKTp0JJvD9Wi8q8s3U1/Hl0YuHoQnJgWj1n8715k1CGWm
hOg/zTa2IDwtD9ml4h77QMaNJvTLNdSPORv7o5a2f3psexQWlVjg9BLnmhpwyHdr5eyNunSe8BCT
FNvcs6QxD1KPclkuwm4cgquBSVIa+87M4MTFJw+kGX0dECpF7PN7kE4ZlYRJqI27kdbxUTEnXXzB
wWunrKoZXj1kmg0unQqqpjJDLbeN2Ey39n8s8nOplh5S7j3zmlqc4QneXzwH3PVlucoLz9If6kUw
YPCvYt4CESOzv5oohAtvEM3B+YzVQ5wCfnDgzPULw42x0i9VYnO6JFVd6FR2EbKuntkXLr4UHdSY
ot5N87UjWY+RoClfF4acgeTMhrr8cXDPWsWHFNzw2WPoPQVLM0vbz0PS19Wnv7de3vuGGTeO+m3D
LKuuqrsHo9buBedOrWWSrsh5nUKb6a9TbVGzsayxAOeVMPcldl3b1uFMoiOImYp3+Lthr7GEd6jW
ymmDvqPg3Ud9ERorZWp56dDe/o5OlrPWtAIzCBIkB3kYcL8qrAAA3eaCysMRqIIZqbYmFzbU0mdI
/Sb3HHqeMci4wB/FOcj8c0nWuaw0hg24i0CT07Vbd/yyThWQI8qeBzFO5KUtWHmwo7r/ePnBjhzA
xJ6WpBuGd7KWO99kYZK7hwlhX8rbT1ejdCLmuLXhojtfOQMzCTisMoxK6ILEQYZCzsCtDJKhkVAn
AuRNlzzfRHDy0lB048wYY+pPPxYDxL+JGbu5NC7qWxCrI0vCZWxtV3OB20NfDnBsug5nU6WVBsea
j8xaacT158RVat35xFZcnAVPtsn31z3ypJa0vBmLkILJHcHC0qwQyiSt7v6pU5ZTJLSyomydS8NY
jangyTxUYELhK2JadoXQLQ5QqiKdz/WSUZRI/SUWZUaQPMCSu6izAzjKKqp0h3NmoIQnjY4aOWyH
/MlbZXBpYYwr1NlD34FdzZeEYWqnjiDHgerMxTsTfnOm4Y8f8UIpP24pX7DY464HxRP1noymhrQZ
zHDaRFbFaJx/n5NWxg27itG6xSYQUNGiYlhkhR0c/ubLfSoK00yIKoDRziq4NE6tCtbDEijtRVV/
u5/ocwKaomq3U0QmV5NzbQyodm2GcHucdnNNohL8aShuNRUBRjDx/yBSCTZXRSSqPCnKwKHEHbCq
BUuE6+1MFyE0ydnhJCxFIRJkiIB9r77oqFvrEYNPQ9BGPHScAEsMhvWy94L4cCBrzj9smV5rNZxe
3RifevsghV2IRdcNWgEFqKcOrqvf1yPYYQsF74Adyzh00OqPbLNMGSy4WFNNKi2p0kbaIUpqd9Y7
9fw6ESGIOdRzudQXSdDv0Gp52OmCJUUQS/lAV9FfeUjdltA17JccJHqLGYfhY/+6t2AKgTScKctE
OavsN/WE7SjYhl42JALnvvTFzcO0S4942BgJAE45I0BmKWy7ZPlYHE4eILOHXw8Q9PXdfZFMVYOD
leV7z8pfF13D32sBM2SJ147eBJY2e/ai5quutH8QiKQSule+VxxXKQZRCQDpi8X77JntG0BdaR8F
sl2TmNA1t2qYmj67ZptmN3tWU6jKiPBSNYxcYkP8Fjlmpc1jdcFhXMeeegeH1nAQEOxLChSref3x
wKiYFi0jn/HQtS6ZVndqlY1lNv8m8Pk4FuUVP60WSJwrMPHabALd5fVO9YctB6DDdkqE3agjtf3e
ApKFTsjLdIwQmKkIJpQPirj6PYuFTaKYRXqaLmvoQRmmSBpXX3wtZnoHpEwtVN0mgR2LhJ8alQEs
6WCxlFXxESYss137KhsDAnrbGXKzcKajXWtm2+MkKSqPI5Jxx5Som3Dijdr3w0877HfB7OYYYNa3
6YYP1cf920uRT+gJbi5htaIJM3DOAnb32QFD8CETYOm56HzmsOotssg300Waz4IvU4OA9Ye0VVRA
/SbJJ/Ol38mq0Ts02chzgNjsVMOPYKa0kSWy0ZWeEcST5E4GMjYd9hi9xE3LM9z6v9pN7b+VRjS8
ezHDkJ/ekpaB4wK2cr6ewXDMiF4Mc8s97rNyFJ3TBnTt7To/SlD0iQtJSWmSmECGW9ErveHXE8MK
/MNp2J13KBzJ0IvXfRDHKr/WmENxROG6k+X9sov8Zcidu+VnV1UABz3FVVqlSvnO+Y21NnM9+qu+
u/Q2DGbhP7CFu0K4Y0ctp5iB6Hy0sbCRvUkjRVvo+xwmBbKQ649xfSgKojIHi2X40KTO+vmL/QNg
jJLpw6wDDYnEeZnVM9WzlNtHuRWmOH4Ajjc+YaGnxKFsSlP+GgvElp1QNNaVJ4wm9iw1qqQt/e+u
sHce1vX8P57qO1YbyWGU5FgljRMjeyqWGHOyZim8vz4K4ryIB1oIivg4xO57LKKXZ/LRKXOq4Kyh
zZGhNY+OTuaVbl3MJFecTYx9EfsisN8FpXQ3N8MLt6LG04P/T1YoDKP/uiiPjh5+AMTeId23ow02
L9f8qGNpfA8pis3EwY8OnFULgZWO4Cyi/ZS+B2qWm6Mh2XYRestXjSUnAOsIWjtwAEPRjGEnkGT2
FwJB2ZOsRsLscUo+CSQR6XyMRdwAajkgUO+LWaWgk6/TFC2mIbPWvDjjokxx/R5PRuTVE8rFa1AH
bcEtnPws59dgDZYH5DvMh7PliSFy3vq4PVTT/t7QVLDEdLXWN3IlCwnu0noFLVfF64DPCJtfyq56
L4RFu+6LwV/7AGL76XrDlxdS7y3Aix5Zh6Pa7ZCmBt8NPb3lFKtGJuQGyIdvtnvTknDYBy0lU3uB
6C5GpY1Zg3P6Vym32JegEM0OfDQxeO/Xj6dbm4wbDUTm2jXLEsjOwrKz3EpcqZgKmrMdz1c76sda
iu7Aes/f57mP1YruLfdjdwubJxYJfzTtv0F3Bf5RLfjUC7yjuEH3SOuDfeN4tnauU/7hkPEmKobn
dWTUs/XXi/dcRq4tSqS1W6JiPJRQCTY9j3RsHGNMUQ3eg7zRcerCOtI8eNdB5hYv0+9wtU+lPidi
Pkg/Nap/7Ic/G3aMT8nW+D/ti8T4R83hoo23xn/S39gfquJQyRJfLdE23rRgvp4DDuo6chzPKXb2
LXrI5fdf7qMJXX78H4fOj7RbGgkZmdpJDQYysTjQ0mWy+1JsilFrk2RA0+JpzknhB73LggjBKtR8
yVaHehd3d2AEkA5V1lXuIlMsvHWCdQh5aNQyzYXCMIrKag18XFQFY/uKFhF47AXWRFZ7u+t8BJFs
iLuXFWuVA5vnYxRMTFg0D/ARYG1JVOWgnmXmPDb+FLKvYCPH9cNhXms1UzM7GAX7hi2HaKHW243F
rnKDAh9FJVmk4x2Pi51F+CCdbjkT4iFXMdLjGVh8HNOFGZ/qE1Tv95cRCcfsxznck0cdGeBhVguk
K6Qsub77po8c5Sen+PKU8MBVaoSqeeFYousSEPMpkgTyHMjNUsF5pFZRYwx9UqdoT4LRPRoFXu56
PEVXIblroa6kTwOrHgVbcEHG2vOlkhI+vIL70rNrV5UTjG2SSFoF7DR4y8+mUEJBNSbTjlGndwHW
STv8vuSeVhHQtN30tFQBxb0ADx41d0IG1HlCNhDuGIt+IMLNSsuKdK6JJAVQccU/XiOz9K3m0Mem
LfUjnbKgBloc3CvFeOCe0/O9IqgSPuuzaBS4HaNPEM/8MKa/jjDVTPS403SeCEsktEj9nvUJsacZ
TZ3XOElyYP83QzwSYAT47+kP2tTvdGavNBVJdBuLaGo79SKWbuX8VeFJEm7j9LoMpij5EFbwhqio
IyakHsFboHfCYCrtcXbB0BgYf9BBEp8RJNpLltFLS36aBkWc4E8q5VJ/13LblY+omFRjgfRDIO5e
KZ3yzkf4GMGTANGkHh6tFjBpuYya5xd8JYO5bA8drK8X/dhHb8S4eYLN1aUu3kXEtpXx/1dS7lrb
SZkjvfcKp970TueL3727FwKne1KqakcW9hNoEt9vJilYG143l84CO/09cYEQyh+CXbNJaw+rNtbz
bU5RQVeFzgzkXV75G+22t5tjSOk7PPOfox9KcHSh1rxilaVUOMDEw3pH+uNpccJbAuY7muQSERPn
uj7OjScDTIAtamZRTpMNXdrv/N2vsodlERTvWYdZ0evr8MaoA+K1tzE3O1eNMuOjBp8vcrkrREsK
IEkFGYrG9LlCo5aH6CjV51hDM8bp1h7uGYJSU6kjq9drH8ggQoRy5t1/ob34P53Od9pbxeN92plc
cqGo4iBguniBbCuU4SfF07tt6NYcrjVwkuSkWA//tIv6LyiowbiriBOyCV2JD/0R+LYSCDHd3MeA
tokpJMvKvjPQFgDCaR8eQi2MILypMMrZp+tKX92cDIZeu6SXqPrNJMGpVhhpphCiLLX0hgW23laL
aRpL61GMq6Pwy5rmcjYseH+ZaVNTmt5itZiVG6C2E8knXUeGueO2lbPev12lk/lhJdRLVQVioOba
0wZhhIKq6U92maFRIbQ8BBgVsVj0k2jiIjTtsT3C1odcI0KS4T0oFUvldkSZ0JyUNPOOc9T/Z36u
aLz31EdLwCT9kINMI9zYrQ+EGotmvQtTkmkNpEMt8QVTJpMo70pluAIxOwJ4N78o00Fr5T8hrcJO
FTqPNUn5/S+UZsKEDVKcsYG19PIef4WQrzQVWqqzCwirTF5UCoGcQ3IlMhvozCCMYcAlAXZcUdCT
O4FGFmkrENacvZ+yVV0LgXgYOq9pfxjmaWOde/rwX9oXNiFTymBRJ67fOkrqCLWPgVfUQrKGQV4U
t1shIQ3LI4OZi84htm2bbhhjmpg2onRkfYM/HjBPWfIVPyYPIZdCByBdcEC76AcZt7UVgfeH9y+3
X2QUURHmXkCqxNn7Qb9offcscOJoo25LOfslY0L2NmZlMWVkt4gC2Pi/0qt8T7bbl3t4Mw1CwcWH
dBcXnQ62dfxBFbwyv2YY5drs7VNdWMZT9mYMNL4UUZhBNGZR150fF5kntINd65thknpcVlc2+DqW
9fM6WCb1JPWzdIi50YIzINOIui+a8vGEctxPNpNeuBh31Sp7GvY76z8rC2cOwWLYBj3g39PuA2/D
LgXWj2aoQ6A809f12SQAaG4/J1yffTg8dXSEP+JwxpJrU1dokI48ZRN8I/1fGqCvxFG27qDmtNk1
K3EYeYp2z/fEqjLGVBxsOdwl74NKgjZP2RTr41p875194x1AYuxRDniDBinRdyijo8pDkQdmBTxi
3A9bP9nJEtHdQu0ytF1wInzjGkmDHaAjw12Exga0ZrZdY4QS/PxjURSS1+l25EnEX/5eSytkRLUE
+MVRvPnj9y/KWTeHTFOqcKiwgsubdxhNb8pnKD4YNeAo6f9iO1J6CgMi/Sr11C1VCleQRHkgkTTN
+9vTQjMGc3jN+ATR7iaLhFjp0ogEHS1RLtfeGg/SfrFD/fYDPAv2JYTWxeXq2YX7IKoqq0asuwNx
0NJ0mpwvorQtqEGLBpn6FjAcaZJy+J0is1o6/8vpc3XeEvqpzX2VvqF+wdFiw9awuwfvmqOACdS+
FbJYn4RLS550zjFGqf8zzehGXIBWH8KCRTX2rXRN5tCufY6V1whEt3s2AQ5APn7wHvPqH33mXXu2
gQb9cqu0NkTLThxnZOPAtpajBc7BVZy1zzOyN04XjVuhKO4bSVngqnSjMVl2TXbDotFTzsLz/DNj
BdQF0ROEwsoOFAeQrzlkpLb83aWxjaX3Dq9Gv2SykXaDwIQ89Hxbs13/GwoeeWO+HSfcq8QpZmme
AWSr0B3uiLgRr7nxQM6qyh37r0ID6OUlGeYiblovqKQ9hoObxbaXbViOovmEfz+qogeh2LcxlOgI
Qwtd62T5rWunDFwlsAYItTZeQQ4G1NAcI1BiWtUuTiBGTRq7f6tgMx1qIv9+kgP5DDhTNS6luMEp
c8EMAVTdArn5J6xeNmGgNm8WiNGbsxs3r+l0D0ssO5SrYHDR4RztHmkKtHgUAZmOrfcoPBs7uLiO
gNGoCwTrQ3IaArloyzvLPgOdShQdLzNeTNmT9M8ODig+nwluHGvM1QcvCo9e+O4P6ixieavA13Wm
fg2YfQMqrxKRJgs9uFX2sKXtkFRslfFe5e4jTgfIu50gvudSNC5CVc3TDAo8GqkQF2Pwk6hZmZ0g
Wu4NH74daOitdcD7hjK09P263X2sicYYz0BlMY11sSBjPAUdOL+KR8t/dNZDdCjeUohLf+eRD68K
L9lTheVNcE8+7fC7X5SpgBBXNrVwgLFKe8SIG4UlhP+2nn8G+qGl5jva5oD/vZm/wEHzXkU0GskE
PlSc9qKRyJmySgU2zNFchTK0FpAi84lqGjBy8eGEM47hnJ1ho+IxNqJFFHq5vFzaXhOSeroYLKjZ
wqdlB5LfbF9zkX53IXCJHaSmvjZrycu5Nd7ypHE95UwaWsQUuwFUm0oL8mnWaiNcDPJex3L9Jtd4
6cNhcfzcm5qFhMZ84K5+tMLTS8vi+jAb4ESVNTWvaYriJtBLL1FLIDQt7HBsGamHADGaP40YFy4e
Xb9OqgjdZLxR83mh9PVDveL+xczNSn02r0Vc8ZjMzZtQL+7hbn6YxUFjzpPAQz6xdB57+Ew8x33V
KW3atjNZG4Jo9Bg2+sowVmbq9QoMWcTkk3fVArCVXr7y2oJ2pkwOMGB3LeUKDLIwz1dcM+MAPdVz
JHT+z6N0vpmDqdyPC6G6pTwzYaCY/UUVvjfKkOJBhX8tXpdOy6gNbCn7A/xz4COIiI2Xph1d8umF
IABKNjmongVk71pYzYORw9tmIOp7oLQtDwOPs2BUyE/+Kp0V1PQCWGvoDPCUtX6S2VMpT4NP4uTs
RBI1EzQfy7dcZRDHqfAbjbyRMhB2pr4bSNVW654vNvsCrKfqyIjDouWv378+VKfdxNolkwFNrjGY
Lk8QtLhXQDE3byGOL4g9Mf7bo00Jb94P/qEgnyQliv3iHMCSxjssHE2X1l8qB1e5IGhupLcNI3vl
qBgFy1pxaXJ630n2HhXFWts8yEQ59M5tFZ1JikuzCaEBt8TLpvjKZa3LXaNEDehKVGQ5/q4YiO8W
KcqvY3QcxbC5PaEXeTDi0jzrfGczlW1n3M+lfKxjpWRl3/8GenMQ0jCwHYPIi19Ecdbyg4hchMIc
/y4yx3jaDQcF0NTzmfdVAwvXu7ruLS4oeZb2xvOgmAi8y/Rh78Gs6eiYYSWuti/JlvKrzuPAUwnr
NsYwoUHduwRlG3GkSrJvyAVpOaQN0P2Ub0q1qk/JHbsaynQVzZlcleL+qPO6Bb7AnmhJ+ckYcpJr
4KEP78FIquH+mSgd0Wwj3SsCfwUtMS/JnDevH6ajwSOUlSOsM2V78NbhkJCtM0rcqZGvTY4Vcxej
/evEUqcUDWyDjytCfXo6Fwj1oR6b8abVzIwC8Eg0PulXyB7k6KPCSvhA9hSEm38jkofYCT8jw+ih
ou2RPL5C9u57Z+p843XCiP75iHApO634xji1BM1neLdWNAraq8+KbHQ013x7PS39We+jzA3Zkl57
1KT5BKvcHFc4V6pJqkATdB4CIxUMFdfYevLI3iqirvIEuBdNrOr/mZDfYaAknMAehy6dcldaGgjm
ecmnvj1+9SegsoRyB89WOWHSfgqgLuyHpazkRc8jO139GrU6Tb1di6qejtxzoDXmdvTe5At6W71a
omKGNvliv2IoqEBeLxZRQNqlkKGgiYM7g0IgFadSLP7iznjWlwsGdiJbYQKehTR6MvETn/TK6NmQ
PssYBi0v0ZgsSuGsMG8ZyQiYW04//p+rRuzIzywdJk5NNzNLxU4F5Df+jwpGtCtzPbQe+4RLvrAw
2dKMv+sZbYanvCJFBsa5bZa4EfMosFccNLj7R9cdnEVXqLIIxCsz0jSuLtsx9ADc4WBEsPOwxr4y
F/HDiFaAayk2Lo+8P2qsD3gSUDgJUYBAA2JYoMdo3GugTSmqH/Q4Ago6lbNKAFdgeEdwCy1gvxMf
zF99abKKY+EmhRSO9l93ltXNc9XHiJ+RA5iWrmKsSywc6bLnA40g7W6yoHzDBYMBrDRmrJSourvs
ei3Q8RTINRt1fsHj1nIB2JY0Pq71us0CjiHKKbQ2xyutX4kfdUyHpQIB3sRbfNjazx1545i2i/oD
ewVA7aoh8zSVOddf3omkMDJVeIQYejyvfpVrHuUf8pl1YUDQXfVuxJogfONkbXs0+wiyN9shKPm/
ef+17px5Hk4enlHqGOway/O2XoqpvXWsSIJmMmUm6jToVFVQklBMTYLAIWH/CBRzZTx/UAoz1jxO
WINb5xtZ/ROzlHdcy2HExwRKgW2S27O7KDDBwFZcpin8DGsU5Vkxg7VNJQkSrfleV17rzrL/ieUj
HKV4cmWenBehC65ngKIQFXoQ5aZ3iATYfJmhIgyyA5pViLtx9fmwI5Gc3WPCzMAw/Vf8Hlxb8ZkX
MNpfz0Ro5arm0WeXD55b9DjopmU+UGIqXlZ+WbzE7xeeusAg3nLihY/xVR+J4TmT3dftUuajDNqH
OZ8dJxqyPwvqVwnJI7QRZlJ9hWMrwGZZLHYEq5Fr7PM0FWJWg7+E199h3bIoLtrJmtADQUtsQCJq
em2OW1MQXGBUy7SDuvulqOSAU6yxI5UxkGLHDrZIq3dm1RsvkR8n7wElnFsdnwPjpYu0sLn4eokE
HOSjnLVtfe5qqh3pAvq2PKjVnIjFneXkRaOPG2hxK2aLdb3xUJ36DXmQ8X4UFO+NskjmrQ/duxxa
oYpXcaZG9Tm4cF+V1UZ/qn/seXHm1L+7YWa1njUmUH3GCuBwKE4z2/ln0TThAzuax3YybSFWKM9W
4w1I96qZDvtKfRbvLLNYgFKMLnhD3btoAwxyARy2NFwYqT7KEzrY+kDw8oRjj1bpbs1uGqqnyk7A
idw0CbBuLXaCZ6GRRxQcA5JfQ+EDc22vzJ8TuBjK5zIYAV6pJ7LBCq//BoQ7qzuBk3OK0OVCYkUz
IvDdQaB0mKaStuflp1FmrIIRcV5LuFD/UNv8MowCzR0TgJ2Op8xW/C75+pFhlygWbD9RZ/lv6Bq4
rAb5x+iY1oQGXf9JFjt8cRTEjqLcKcD9Vp4yUAdb0r7PGHzMLbY4PbKmkSfL3WE6VSqHZ5D5URoE
gQd1GYmOEEw27/rw9f4CBdzoCf2Lot/0O4AJwXZ9uDfi4otZyk6orhkJrmfLXsRxPkgzSFLeI0zj
91dI432Dg9U+/iU1bJEJ6fs9OdC0h0NZLJGjpDt0fbewhet/okM1WNnmpQtEZT3ZDP0ie/vtw2ts
bG6lrUm3kltyT1RZuThEgL/I0ftFKHH6UMjiXZ9NRyr+UO7/qb2bGVB3VsYJGRktbgT+5o3RBmpn
rdeA1n73mKCfb9bZnWwjmfY9qcyYRlsQF67UOEtcekjNN3n4UmduuUNKORln4zrxqYVcVeSxwZH2
Fvoyde9Fzr3VnfSr/RxEBOaH8teA6mBEHaiQY3BL6/oTFpIxuWZBWi+mV55pubcqMB08+fwb8Vel
ZBUlTyEV+HNtdUbVGfy5GjOWlujKwaTPup+QlRiumnKpJiUt3shNiNhx5m2fKnY4VdaW7zZjkjuB
2ua0Son8buxhBTpdDCX+1SP1JU4KmfcEZ16Ak26YySesm4i8prCOmshTMisXws3kiyjGUIfuqrgr
zEd7tCOm2vzkcG+738O6oXZEN3EGj+vlf3lKXr77FeX2gKFziPWCbGbuXzjs96wjmbZdb2Jifiqf
b9RXjwY9cgcizTMXaZdThl9Nu9LjiKTkpSU/KRIm3x4m2bH7a9iQlE5BemPlPlyAguOZ5HKChgPJ
eAZ0lsAtzpWi3lmItP6aQiqoF8YF8GQpgLvN+HA1EFA1nup2SIJrl8hn4ovay7rEk9xSz0y3XRBN
jvNAyauW17+gAgU7B3m6eUREVGAxWoyfl3cii51BqeCRnGlM69vgNiz8YiqKII521zRQNAuOMK0e
yqCe6+WNbd3VmxlgIr9F6bXYracFDWibsA5UED2Gc0Sciy2OTIwL2eeyIB825n7v++0uSMuz2cy8
xul5nogACr4EmP8EX8cBAVFzMZCcZzTj0HS0qzUNfnK5gW2EGt3bEtJ+aGujCiZXhIIs8NcSRQBL
MK1e71+V12mvZ/UFdOmebh7mY+TpqRZlRLsqVsmfgnZqwbPu5aAkXFdgRbTUsQxh1VKSABmouNSa
/Kh0RXIZ33r55DS9nruI+C5NRjKJ2bXGPPe2TQ+z7k6ViWXsq03Uj9WAbcOqyKS0ms8ImyY4Vjk0
U6UR2h7hX3+ii5wCMoDwaxqRUf8bQbkG/Cc/dDcEV+kK2flA5chLMl8X3VlP/eSwMW01kzR7LMJc
n7xFOL61GWpor6zaQOoLSvSOlq+meqlu+pEy+i26kAKfC9gbW9loCkZt2NTWDqlciSJUF39FkTcj
Vo/iducf4PI04nKpVkzgQMczO9pgIOL4+zjzbWo9sDGW17aZCSI6MzgTV2/5zGhwsTPIcBokitlk
kMTIxEqM+nbBKVpKQv19geyslB/Uc/QMZZR1dNTqxtz+0bbUXpahgcU9TaqRUaf8qxwL95XqmC6c
EgwgvOFjlK6x9Y435oFKQmDTg4pgQ+q2zHQemRqYKtbIvvzoUVQ+iS9p4xXHWeMpxAv7kg6tFpmi
sSDnnT++0HduSDs8Hr7O8ADonLkVwwdATdIcd46Y0u6zZ4pbAPvDuf+Bq6bOEGJhiU27CrUzrNS6
VKT0/LkEukW/GubrZHDtOuV/OLTASeQraGqQFYFKWhiCL5TWT/HkWOV2tf5GVdRTWjtrpvRtVIZR
H2GhGv467o9ZWWD3ttapedBw9VxPb/EXXE8Il9CvbHqLIGd+7CHnYQNorMFi/JAkXC++9Gd0Idz+
R/+Acba/2em/v548UnbED5aSko4jFUX+OP/MAzx0lSkxwVgIRr3M+Bl4TVZMgOHY/amEwZVtcEYn
O93pUJMqmV+Vw5wWVcSWTuM05bHFiwom8pHzJSM5z3fqg82L5JwPZ9Wt0PRvYA9QWU6VwwzfA6kc
4VUhV2df4+IusE2+LZaXd3J/orohZflfC4LpftIO+gO6ALhQGtc00Dijk4Uk2MqnHEO8Gl+9lSEQ
2Xz+y7CWn7jQwNgpT6l4k4gebHnaRenL4yQLuocZew3CIWhCHgwElor8ka0IndbLss1RWqYHsclo
7svl2WQZJX5mQKvwWFj85jm7zq/j9PAyirmrL6Tlc1kwtePbI7XB6CDO6aeWCT3TpJVLRbcfafYV
d+lIgBLGI+NHKgaspLtckhfrXz0b66gymMvAPuuBYeWBJE6AsgfZkcRAj90IuA8yvB975XHNX1FX
ExNDJMXAtobBtd+Waq0EXIz0TwtkXH3uXTFC3GSno5StBPWwihj6BFEhTR1h58ZZKaOnHK2HWqIK
tj4e6ZeriOslOGTum1kb2U5AXvHwPjyczz71VJ6SC6EHe0WRd/iPJze+mLXGPfxYfvq15wFWYNU4
couzyMgyvXEQJZAsIew0o1os84AltzzXWrapPcEAqPGjUJaOuTy167uKP2DsURKciapMxSAMmb9C
PAu8BCZr6lE7qg5OddhDKEvvU6tHjFTLzFri54vEFV7R/yAisfDlV9U+5k1qMixrY9yawJfketXH
t1tmoCnnHLI+KRQOh6k31g8UDu9v7pazH1mV6g2zP8FekzKRPnxGowJNHhAYcDIkFLrVTFsLhmAM
o9RcGa+kqa4Md7t0Bv8avujHvQbPB2rbyZ0AtualU2Ii/Czrn/XB62ES0/Ww02obY1aOP6WjzHel
Ge+luw/ojcPEqdTrDG0DNIIFaR4csDGX69ysbIigNkCmg+HXGqvF9zG/Ap0hpZb3gp1sTc7AA9Ei
NOoJJmdhytd56j1+uSrGMxvdG66vnPYl0hjmaaWZzIEjFHQA2aGCVdjoneyRRaIMuzxarHiwrm+T
XoHvY9RO2SpmD7RaYbPnCGTmQH8aYxry6VtIHNFZOUOhKe1uenOMTBq9SE6Lgc3WoHLFk7d3jxK3
EHkOVS9dY1sWSJ46remZjFTq4mAlJvQM8GYYIlQM3lQiJofIHetAZm0fnK70YkEFPFyjSwAYafIW
XsZt3eaRXzyI5u+6l/jTY0uwaxoxNjgHifMjd54TXdFyuGxz8n7WZjozEO7rA7WwcrtpH5ErNR9S
sqahlqRqETHHlxsakJuXNRgpblTntqbJRYjI/M6+8eiGtK85Jwlw74AbhuGvCN0M+SybWw6U7Sgp
jY8q+WA2Mc1WGWKHAjqhbeaAjFTAE1d7I4LPmxAts4G0GApOfkyP9nHljF41Zd8Vbp74HPuHIL4X
oEiqdWLr+ZTIMH1bUM39rKgvW4CE8ibY3DFNctVa6jBe4SOo4aaGRZO9mJlQUMSq1vZdY90XtJPi
ihNs9CYwG1t0EZVnwUW9CjCjh2T0dC774HVUUYyD2EjJP3s1A/GdsF/mBw1FNmKkaV3Opn1lckVN
itb/XcrdqJFtYBbYzPdLKBCrnvKcPOX3+oVfZpcht1zouvHU4kIdsKD1Pajm2TScolrsX+gZTuZ+
w0+ZO98JEFqjLjpU+vIYkoSa1P/BZyaZIDibYw8AiFQX8/LSKcR9Kdd8sRjWufZ1sn6VH5NG5tye
v+ZDzCihZ/ySbBDnpvIZiNcBx0rYgaDH0TlkKweNPY26cUPOwuQuLmrwwTyHhXEVvGt2zHTmh/CD
cuNP7gCB/bzbnu99ozCPzoJH4bBF+pORay1C+LmXRaOMcrzlElr0Gg/xiZdfLK7QTobDVHs2BMX0
2REmc1wwWnK3IkFMRhSnJ7KRJ+6OVkuy2xHV47ObAd7AE0NnayZjOHZiTE1+1s8o0OytTCVoghJE
As586soRLMwGEW4tzop0UH+for/HZHcRjNfT1R6Hr6slpjwGDyFg6yGZjYMbpWSwon2H5B31bK38
f2HiaCPu3FLLl241PqFiXkwIGCug05q0F6p50oVW36E9t1F3xuGZTuuwhdMDIb3d4HD9sskvh+/6
8EEtlwZoMkd7jJ6kKWTJSWecE8gnaCZABIrNaoS72wChUEwKyuExZztViUOwhzjVKY6nSTLQz++c
Q1EB8XTCBMrFDHpoQX/xkEn8T8n0U2vQes3b/xQ2ClxC2VxTLbKD8iQiBlwukGUKqEivOWFAR58C
48k/Z4RIuVEXOChB48qNByG4Jz2b+68jM9pWyeQGQK8doPp7Dw9WfzNdYVsVIO5g8DJHLRSJYhmI
6aU/9r678n331SVLhu9oKQKB9ihyT6O3pvKLYqXV9oULbLintHfRaBhcl0CLiBkseUWgzKtUazXY
2/IHoOwyCoDTkz8Icm8H6khe7HmFOIghQXcUFxtxn1zRyCF+zJivWYr6UCdtD9+OgqSOl28C9K5y
bCX5Q6ki+xWShWZ689grU8NwEyMmiM5qHqmn6VWRpBjIyHvtye+OjoC7Kvlpvk77XJ5fKZU/tM8s
fm09gqAJVURciOmplbhatXIYuHGnwp1nSLa5K4w+Lk6WnZCXc65vkYA2sZZqw9mh+boSwsbgDQis
U06tW2SSssmQ7EVHuxgvw0T25FZ9J/7xt1g5fLd7y/IDdfFySQdOauwhYDyT/Sor2ZsX2ugDB2U1
Txhgwe7yPjTImVDkiuI9NNtZWEL8xcBgP9YZ3Lc/D7oIKJ1zLLiuaCeS3P9XpdQFOsG8TtfSCHgi
4Y1eymnxzIlyCzQ7XPuhbj0UKcN5uPxwO7l58hvueFmMSbB7D2wF/bihNHcvZrNiWipendP/rVze
mBEojhaWSv57Bsw30yrfbxaYnRfbK7zT10UKLNeWGj1/l0YnzramXq+1529UAWVCu6y0Ltc/tCb4
f3FV4wSxZ/JkL3jt3yVEasKRE4Gqfl+D09XgLKMzTW+gD3itFCAaM5zqZjEJUz0tfwFkx6zhXPV8
Hb8wiO/wd3c50VggRH32hK6BRunWLG4G3ivU486Af1zBKvAMWaain49u5P6oaJzQHYM+wzpXVWHE
iq3+AO2MHFsb4fxSA5Sujtj5Wy0dHNPZsh7lFt9F6P+j0uRPRC8HVw4A//T4YCtgtL9/NyqtKtO3
yldKFwA5Q2wx5pJ0Sn7p5DaeZa8XofbYDzei0dZaQ8Btxaa6FPdUoOE9/RKQDcmiv96YNXOFd3eI
nLrECRW1BPWBI4ISZ0cSEH28CeK96Z/xWyDvMYxyIbe+teFupiZefgj8/8sO+yVwXhLHw5kxSbpC
6+gUoSeMPrTPpNzm8rNeYoHckPfSbIQMS2k1j3LCWr9w91n6dued9mtY3zyMSy7dtrfQH8VJ6VYW
Qgw2V7c0B/hg0j/TTPDgGbyLVBu4mMevzzWv+sAscs8Azy05B2RUyqg1Imn5TnRz5w1qN1M1qcE2
YEdWAnXt6+BLv4wJQrvqmnAzRHy18AKIUOWe3Kr/55WWBALMjGzPbQvVYmkzdDsxITw/kaJrdses
RiK0f0Fdpd2diQ0IcJlH7gie9mETEtmTbBbI9CvERdrkty2T4S0KBeVWhi5oerL1JPTp1aQLha2N
tmymFIWOFt3KuKYb5DPsso2ZOQdw2L/Qtevep8m/gyCyOAMLsAJS3psmyTDyTCAjYKWKAouFVX8F
4/qUyCH+dc9PAyoRLZCPvISUMwF+uNvS/xtSZyCUHPpKsIq0PaIep66lcvM6giUbgs5jqIVtpiPs
BPXuEX7d8Jwcfsj7fcp1sEC6Tg/c86sSdV6WFatkPELrWYHme7jFxZMQURPEtIaqus69uBpERxjF
hVO6BitJlJflm29+F18ulH16KB7ujBtM404eaCxIxSMsS+/60/jOQ9zEY+57hjxmM+UBKCHjKZN1
l4lUsTudBN10Qp/wWuCFOL4qAn4YHUqxCVDMXhuFc+jIC6vTkq19CX9GYd4atlM+tKrsyYxO/Yu5
k8+eNg73xlLkfY3bIe3bHvrTlZUefdRjjC0KIM7LJlMRom7F10dXuA73Qi945sha22zTsde6rxai
fLbKvIM/sN3JpCpiwXXYwdnl6kCKQRgjLAMfCHVYWGPukltYRXyE2QRGOTVstpitldQAIlv0cI4U
Aph2OyaMpDZN0UhWTBdFqsg5Lobn05lMJqSSKw/z9g0xpUlM7Re5CCsQLBgD3W4wKi0RzvgAd/4p
cwe5lM/1BzuC4ykDfoFdmWhVlx2eWa0SVwZHfAxL5DWXTdwZqtXbCZnurG51vGt16GX/Igqw3jp3
Bk4OaCn43zpGD+zzHaARrrtHnsyNO4rLvWJW6xaqOUQEDDSCS+gnCEAq23TrN8citWsDiCevSCJP
mmCPHi54TnmcC9kSPPqytoU7G6qNFkU3PNp3suq/vFzHgov11Ic9RFKSHMGd6PwJcGR1jvmo8vk9
PF2ELEG63CySh5Pr4oLyC0P94zOmEAJLlc2d3csTwdedVi8p9Fq1pqdwZr8lpzW9Gp13lRlQzX7C
dOKr/SwUOXNKQT9O0yst30TpWCPpc9JMgCJDY3jCPG0D0d20Uf2Ygh3hDzsA6W3lINCXVrwth7Z6
OvnDNz405oerWf5ul1CqrNfLPeqT2pCrSWjOsJkpNX3umyMP3lY8EJDqE6jeZfDAGZGB573zHo+V
dgzXUo5E5T/faUhyzoeg42l5BCp50b/HPuQ2N7KlMuNzio52jBpPAUY+Bk7u0sTpP8JZtAyJgeDQ
UeLaPgW6lwzpA8OyZcJklyi6G6C6fW4PjLltn4Qf18dC/w0LsAcEzVlUUp22ZtqEGqTOxEMEjc6j
7aY4N99y/+4Cg6aKJsiacLFJ27P899s6SKMZMnTyRGIV931KaP9oIVzfuqPpRcnKVd+SSdKZUTKm
bFhdXUlomPpsFQMWJg/MoiWzzOgdJPopDYBbPT/5UwgYeUKZVd+ksTYAqInRjIKtjjY6M4iI1w0m
6ccCd+7vUKev5cHHa/MZf6oXxmtL7XJ8MLlCpvKQKABZFOjF4Lis8tKn+Yaw1OYWb4KuMkF1b2pW
tfzvorAGDcWffLw/2WSEDjnJrWmB641jEZl24UrO2/h3EqBujVDWdCKCMal0CUBUQMpBLsqv++9Q
+vlq0zvPQG/ybcEdzf4KSH39zhfJwYrre08juCI01u6XDwKF5R01W6aI3sVnLG0wV2oIKoXzI83I
xZygRB9oRNZG3Md38Pdsqq4Oh/gkxfoumVzO3J3cDEjdM+PeH4jwt1oTtrUI76WZmNyHi2V4OnuI
oF8Fkvp05UQQsmJi28HcV+GvkVaDrFBtu6eKlkW3DZpYy5ZQkDRNypo0D7vKmPEFtLnwa1BuiiwX
17yBMYQY+vMfkYNJCIl21xVijYI4Eybp+j7StRhXGtSAUNO5N35nmhzmJBhjL1wA3MbM3JjxsXe+
3f/I87wdLEAtHOk4g0P8vS2KLWEVL/9BjgRPrSE71RCSNgfeK1XoBYjlITeAuOxpALD+wuYx5PPw
qW3kdYH3OTZTONLHNOyvZmQqhEqXBoP+ZSQQ200+44HZbQwvZnmEY7n+E19Rkq6msqUUM3nxHx16
tbJzKrE7hmMffhBRT5Hxo82fHJDXe6zhsfak4j1mXmL9ceeEgwn2JXdT5eZqbXeZyJZpTI+SdzSN
Db5a2/qAjKWQxX6XHHU6nBiiArztQYGDmkX8D0+q4ccy+IxFeiw/vfmikAr7bD34zzGW9bBMXFPs
UAz17RDTDGgcKPQ5igvmmbJnBZOqmXbNtfTwL7u017qp4oRlEwhAAOvFiIWRKTBg1ylVWz27Z2s2
YoWmrEcme8bosLmRaO1vDa+Jw0hW4h3LS2SBRuz7ymBOup2w6F3iq8fm3dfmmnnJj5zP//7Quky1
S55NZzYon7Vz+LUwZT5gpUIyN9fF0baNkGxkxtK+vuL6jfYZay/7YRnKWuK26qQd6M0Y7SHv98ta
iONPpvRJoK4KAPjmqq3iqC13tjGGw5Va8TN/fEAUXsi6EVJZHzQcPFPhZrRwQIFKBN1+pev17UMH
96ntEQ54LVP8u4AmhZg3km22mKpuezdVGaO8uaBBjeqAw0hjQ1qVZ7500Oj9N0bGdtQpB3qpZbht
b6JjO+b90/47Vf4qZdZ8Dg/MkhznY+9sWFBhJ27R+nXE9XLtyQiSC6/k/Ia8Vr3/aMzd2xR2m2ew
d1knAGKvTDW673NGMfAN0w1pL7a1Zl0T+eWSaQTODZgzmlc9dtIiZzUJbYot+P9gtiENWyeUNRs3
7eNN6sh2x4Nuhcuce+QKLOgccnoyjuThYn9CaYQvNv8jFPwLI+k5xZNHlpqUBfCaiRtaAdzqC4En
gYJpC+92aplq63OXAxATHQCbUeZB9rb458iTRJYeWa41frKZTsivXWxqNp7/BtKwY+YeF9BLze5c
sXtUzUQl+9WuznTHate7WbsToEjO3adkMIDlQGIprhO1Ws1JapBA3fs23iJuCRSSgAMgR3a5earJ
iIpIswk28E7E9qwjIV3HR/OUbTNiPdfDC1+L2qj2OSHS+srFfQra+dM8jtlqDeFQQPglJ/7T06UD
GoFZscfszJa8Wr8lqymBsDmNfirWrD9xuFz+uYuRypzo6kZNWiJoAJ5E6V3JbCSzLYWnUGtVZY7R
6oDPB8mtX17ErQqveO0rtmDIsEynXfQjFtttjkKUniB/p0AuUUb0RjeVNdZT8mbppGLgFE6l4XYz
3+EYWh0pgo7h2ILRDD0PvPyCZE1xlZV6TVPi8Q9ZIbOS9vH1XEoKzBtw7IVrkYjlSwDRSnSqwGIL
G2aD36Cju+zq4aUxkNkDD1rCIuFTMK8zNDgZrDt7dKm1Rj5FgMintwcFnUBSlCYFKQ/Sx/aSMEUl
+qeDBbNqiyzS+wwU6XeixARhIpJpuLD144NDL5PvLyzTP8dQtcqFoQFRYPY1+rBhstzFmZt91ylo
Tm4gcgB9yucGkjShXEaM13HercTkaPPB3O6SLs4lvshdc7t6orrWY4YSTsTb8kime6/a3HGQ1wwA
FfXS1Y7necasWYv/WDl8wXzmTO6cm9oHfpDQ4wY7cVaQr7QyH/t1255AzOSz8AZ9OUxKESIW2BYv
/eor+nafaSwzkpQDs2imvrYhAqwNuujuNBFkOD5AtzvWNYabB6yxX4cSol5ICkl7IUO19+x2Kacj
A1YJBGmnLj3H5lFYKloTzN8aSqbnkHqMcjmNTYhp4dxxj6HXiMTq4LhGzF/ITG1XJwou0Oqmzi+9
uh+ezYxrhl40Oy5VOOKQfsC6uDkc/AlLSMxrGLAyu7cDmRQCq4vObeAx/dC9cjqkkRbgargj+EGg
jWFCW6tLXzAa49hAbi/R1UPQCaDeJKrLztX4bnwssKU8Si43y+WPKjdVmkK5tiuIUSqNufHhFh84
23BpndB+BuV0AZgx68ymkHmZ+Z1lhPj8/7sqFb8BHufLZRZNopV1ltNhqAJuXGIDkUwYXqaA+iFw
FTzrs8h8xl2X1VVpzj2JSHUUmZsBnw1mz17iwxsykSnKBxaNLu9xO+o+Z737quct8lVxUgaiLHhz
6gAxJTMiWd/4GUJGQVUPvqNgWeIIeo9rgVzFdmkL6vkNWzpu1cynCUvVkdQ4NO2fNvve0nnPIOb7
kTyLpMjCja3yCCtVSgKf8m6zafzwCCvCZ9JGFv5bVNnShYcz/+NiNYiO0EJCVYieyYUOL+32A8OR
WddiIohxwI+0I2WmT25+eVLoKPGXWXBKLYPJNAmg9hr5gMsY7KVRVoHXgOfIOam6brEtR3vgP1He
FbSdw5czmlGH4AlSP17tQjMcapNddBUZJJ9jEYa5JpkBQY8ObXxc+TveNuOs6IDR6SODSpWRz2GU
le09y97RtISBzhyVrbXDbmqF0A3ld0wdheF7x/T7jP367ibfXevzhae6KWV9/lAXJPo+FfEwvBSr
8d23FSrmiqVKln0n0vZCsLlKkyr4HBdMYq6E8lT/JqRYAUUiyVEG7pc/1XCbyT2oF+mR5QBAQjIR
UrJSPHOwNeOvkVrYV/jAA0dFurIOxQgXigKCciKp058e8E/29BAKPcJ+GKpMIO1DI3hW12eSE/2d
bMoGHOrdaB9FqxuwxOyxrou/DhA6sXF7hGt1LZNsD9E/haIF0YdUsHANN3/0gTOtIr/VNBIJQF3t
usuYSld4sDNzvXTr/0Wgz5jDh43yA7YfRGdoGKP5W4UlAk21PEW0zKfcG4NAkwOlUK2nHluX6BlE
nwznJkiF5VaXtCXFZF7kOktH11cXWJoOP0jkFfwyf9G8DwUhuHBmpBmmn9A08L7+33yz/4uTjCKr
ZLRs9OMShXIX3eTTsR0fdqdCr3B3KI/Fh4P/ygSNbthqc5Kb7BnG39EitvfkuovwXw2TzQPZ4/p4
AWappVCNPRk0pgpyrzvfOudcyb/n7ADOjgMSOz24invUVMPQyTVOmyDcJmlRrEs+K1qS3FXpghEl
0cgwIArOkK31FNfYrjgucl10e8SzBYAuQ1YxyEus8N7jnTJE9J1ZUUskS+GiJw3oygsEtUGeO8lR
6Qe5LtP5vqwlO9jy46DzI9vmvgNeZsZOTn4DPFtl4VK2+EgKDQGJBF63FtpPaaPZD9OfQBQZKA//
Zxaf2rmjBh9wvwLjEaqvvCV1yMKKE0W49Ar7t9e8URkDUz/iNw0rGa0lc3qfj0L9RUiijTjxvjfG
jkfRgUInU2XLM05ZgaQ2OcsA4DLYSmyvnjUFwuu8B5B8qpBcj7zhmdkcx2daHMJ9GL+BIpYGTCXE
B5im8TbavsVsLedp2O0ak6fTN3CobWzXOlJigJ7ZdmFTih9a59uT8CZ8lZX+HY6jP1v45RwoRdCq
3SodqEMgC3rteMBEUmloqcAfFoobrWy32TNmOMBinZOMkdTQ+ZLlQIcsqFniK/eogW//UFczncns
Yb/WlAs8uhe57JSEWcy8szkoXo56FHs/k5kPuUAaDWT+h1kf2/535wfeqRvgdzBpjet0dwAmEJQI
TtkyttJEXsrMwIoizkRoyaaIdqoM5WfS+WtAS7CT9zldclroZ5Go/Ii1jPdM7iLIjOWHoZ/9SfDu
tX+/WcTU8f5lXBwxlvsPwCP7V7kSrKfvmxhAXZAN4B5eY833RuH+GZTvMNxdv3asiXd1Lt4jJeF8
x/blRl64CRe44EgtDNv3c73i1SM5WJ0OT2mkyayjgxrURu8J3ILZUyf3qlxjrhkn9RPFYwkMdujG
fNHBXjANNnqkQWfpfAaIE2zbP0fizuQxHJtFq9epBJds1k9zqDxEhuwOZ2AnSeBEKoeWGYNA1+MX
zPNAz+LNdZyxhasEbjisV9dii2XDgLtEtsleUWdPmIL8v/RqB/T+KinR4moH+vEQy67MSxVUUvxl
TzM98ON/Jvg8ogYwAqyMfHq6SBEmlVx7WwXimv2nUbtl1m1ShKcAUlT+I7iqyRyYpwSYw1St+BPp
6MISqwo5E6iXVjn/+D4l8ruRQpf967Jpd/fvF/k7JEf2N12q42plwN3NVdMfDyniHLv5m2vc7h6b
+r7YjN+lnIavVwRFnGga/UP9Fc9chnVeEBspVaKzK/Gxa3Bj05VRAZGtVtdIUx9tdijv8Tno9xF0
bYtvtRUow5jgn0XxRIgs9WtpYDtj63pl9aGAK83x7z6eSX/gJuiUqeLQM9JmMKu4NaBPF+92rKO5
VZrWYlQddJjt7Q7HnWY/9kuxMsS5JBCpyFWiMFk2dYpoKA+awcq0rVtSzos4ZC8DKOWySZcIjfav
esliFq1r5fklDPnUUMR2jl9rGJ49fGnE5UYePiybe3uxwO4TCfSeCpib2fnGX1WXxf6KuTNp0Q72
8J9SrfS1hyH34j65riSnLT9WrEjBchyBzlTbwem2sJpJIUTE6R+5QTY9zjcpnym8wc0fsWZaye8B
b7oVWY95iQMw6xcoGACyXBGr14RYmr3Sj7hLaf4FVuO9U3Q8UFPt73XG+VIXYibfQ1Z6NwN6tOQn
ThJaHkD0GXMznJV4z1mcgrDqv4jQMn/yWEF4WRxpbMPinFYpg+/s+R2jL79AVo9tIlpNAfiiRo4E
ytVohdDtacggWu7eaIN0gpYAkm9j1OqW+tVCcjbQU+3ne4eLUXEtH0NlPVzRIBP/9acfEh52PQYn
K32SxjibwA2BZjZUi2mOdsQmwnK7RTDq3sQ/J/zHICtydAZH0IGWqGedp0jX0YYgDIiXVHRXoQ0f
L6n9MK3ecBRDTPn33xkiy4l/V3RMTJVvub+7ZBdsd6/RKl/qAOGq5kcz5G2UxVgHDVdRrSH7Jfr6
8g+8vGKnjhBwlqub4onpQ8pSb8qfFZ0+VNWifRCvir+DET2d2exi3zqDs8xpzplcS6VnKrjD5XnB
lKyIlIPgF2IUrixHxNNpRevq1JvunIBSuUXs/RBnpu2kdoarsD+O4GVwM/IeIhzriKbQS1LkMV9i
yAlMl00U1JcdeEgP5W75FDXsm+EKHcLnXwbzpjTFWbmg9uYPR+FofGQUUDrtJ972nqYOkUW02PZz
QBnnL8CjmOlrDJO1WE7MfkSRvZ3yWbERBsH13ksCXgmx2TtoMvbV8tNz+JDMYvjVxFZjLcm3OQHA
XKbRLfEYlFdMWxQRRniOUiYwj/hwT8GymMcgPOHUZFPoCz5rrVqrtMegrVggnLafTY1LXWdeXTan
uWcxnl9qVfu0d/nqViBCfIS2PKypx0/1BIOh5oyY/c8tw9an1XCrgBBkWdKuY9QOQzI6G18Hp0bS
+SAe0mUdK3sDRTWLiWmE43sNDukcEfyWy0tXxq2TtOzGCqUHolZAtPQD5qDlUNMlQu4jhM9wO7Da
bB0ED5qKMWwi8gRgLWE3o5sTEwRtnEMJdeaLyZMB7vq/vvC1CQDQmDAi/FGc1pdxcqn5GrDAIqpF
BmyfiT0XYqsf+fNrSkGkpMIjRmSJh6UjUUsIMspAuYOwTgztArI//f7Uf+LwxRxGOpAuMPcwmp+B
vMpc/fsBBNXa75ToMsAvINYqVKQ7uFp9WmorhrvfrJCaNNSFAlZbvjR8V8HV5zupGad2PNU7Q6ul
EB97aSInnOUDCxOLS5mU6EGQxIJUr1rPyFdovWA2fxQB5S9wctWwdlV43tT++n2T03i/eQrvIbxo
9Jk68eIJnOPf/RpYX3DOdqIzfkpjroCbibdIVcLwoN/dEvT/nPKix22GMTY0MJGk1wFVUd84F3pY
kMaCNcsrfPxxHBBzJCFyovzyKzIK9qNIww5YGkqScp6AKiLoSngjWGT9qeaJP7MywfCyEr6Nac5O
ZVlm4rTnrIckZF00desCi9j16fgpFGoicL+NFlTSzUU395I5XsAJjkynGhu2kCR8JNnaw5ZUJdRX
KRBxKflsY9UI9rpW1uUuQz6+Zmuk21CArK5NbAbVRfYfQZhZPaW73tC89GUSPmqEUfUVp0NcGffU
q/UJlKTZFzhliilCLfl5HUhnaHWqq7Qf6NyiJCDOzF7KlqwsBIYE9b1MmozItbRf2T98cHlEzfya
iqhRvvsVqiF9Q9rvrWpHLxHNetAk3L3madogSBDEEroSnnyDBliFvb5wrcP9asQWtcgo6Uw0kOEj
7TPe0oqb69hADVWF6aDhxPu+YTcUHeX3/OiUSVSbuZt06lb0zoBXCyUS3aNedEC5PMR9Hjt2g73L
0KQ8a3ZfIzgwvR99DKXi/alsu7yKO0Yk5+DI0sm+RksiGVse0L+lQSs4dL+XJjLOesXHDgFFA5Pi
BYceNVzkw6Ty0fX4s4HpMb67U1qEhaEGxFSryzZx4yTjKpCtPl9UrBb8Pq70YNd3nPhn5N7oyXtX
cD7cKDt4LGAd7ylSKJuccAzNsqDgC56D9Jdxm96alSkcnLVAaStuMzC0vcmhmG5xlpX3h9Q6V6Kp
UBNcY6s19DMJRj7MjuSCmgiq8/lgiEHNAiyQ6YvzKhGaZG+4JhQXd7BqtHG3UnB1BOhyJWuyO58+
uVhWRRU7usCF1neVSIX1Enao2AbRug/sxC0YpPxeAPaMl/npYg7Ep9kJ6kBhExNVKJufpxCKHr3j
ANCJI42Asik0miUYk5MLek9+q8Xr0Dhxt6pyREx8brWjp7KdzLc+DWlozG7fy5l/N+ipjat4o+uN
GjeAJi3SS0J6ukz7bufbClro7r9oUb+AowF4Q2zraVRZwGbmjzRBMhZo3ImlilVlBHIp82FcX+jl
tCYTRwDBPo6/eWNX/BRd7nSEvYlJVqxpmCt8ihx9JN0N40x0T0IwCQ1w5AXB9/Yn0S00+5b0q49/
7rGddsEh/l8SAbMYGFj4YkmjInEHlg6cw4uLuQqGyOlayUbduT/oNHmArpGuMraFJmOyzzEoA7hA
c/3ux+G2Sq7sd1eJYXMKQfCHGde2s53xu1S7+ij9FtQwOWFrPtfU+Y4amhUOpqTj5qlrQaN5IXZf
5TMi5ZK2O5Ig820+wanRy3OCO+Ci9CMkh2Q4++N4+YZVmQVZZjglv0ZGgadFKQ3VXaZtmCLF72OF
PkCSU1/BqgF16woEDC3kV/QrE2GTfkGo/e3kANWmAxUReuZAHb1fkPCHzvcPb/4PlFmhtqLlCwWe
bQ5C3gcYveVU0RaFtTCJ0Txy+i1P2sn3WJ7E6mVfRfppRvXhudKaD6w2ESnRmrlIqvmdK2BF7bAM
sNDU/4nPUBUtzhP/Cnpc7zQimiPi5VICBdJyJpJZCq8kxR+BR8F58bxQsblkZgVC4wlCZi0Q+jzZ
Y1HDhJPzDz2X79G5gbUdO2fVbGU9llDDDE9/lRY0NGONv0HsR/luS+sCD4AKc1FWyxNUanwWduOb
4r2+y0TvrKXTfFdqbSvMICeKnXhbbdYGqbublFK7w7cjjQyu3Mk8sK2nU+PAD1HkfUyHowLelTM6
gSi5mzYUtXZteQSkN/FPBXUXqgzaRuxkmPEa8ciMvR4ZQyg1PFfDcR5smWA7rMCHH4SNYDV8DJWQ
zUmyPN5H8RniF8rsnZ/D3CGPEU9GeEjsZZAe9qyH4z3+p29r5WYd6MuhSpPtXuoZdsNimQjm+kot
J+koba6QSiLQGTlco11hC2UC3uHY3yfht/BAGiJ8JAQFLc0DYjS8oe8x3ezVF+Hozxl93GofMxU4
TuOxpmXhd/YeOWXyNZSNn0ptQdZ+2diHwuavTDIlUmGdnbor6jgXSIcqNZY5fPi5SDWS4a9VYc00
IUBhmGrFEnkA1N6UnJcueDzUbLQ5yWQgsIZfLrMvF2o52c4ubO4Lv+xqFEX6iHAG2WJp3zaL0EhG
O8vqjOPUhH/KIUGKEiHW45uqmR8OTBbi8rPGWheTd2EZao8jrURCZq9ObVhMhBDGT3R5QiLSZ7BL
/A8ax4TaxJu7/OOX8m29VieTTFQ1eFGZwvEtk4ptBDLJ82tN0GEJl0Gj+v3GNiXEpf+YPZca99m5
kbp6HoQ3Zk0qb2VMciXeui62kPagTB6TXrYhlbQ6ccoxoCdlTvml3+Z/USFUoifA49m7G2eaEonv
2pTiYx9IsiiioHI1V1II3tg43C/zkQBSkiTVvGK7jfQ0LANhcKhekqsZ+9TMsiSEsZWrqGL4h1bq
pQItGzZLSCt1P5+EzWqehwRqoQOPOdLJQyZW4Qi7sT6ytAws7Zq5KWX7ZLWUpsK0yWwl7zzymj0q
rY3LCghnSGNHesgTiQYpp51tcmgL3Vhlk23I1UMRntv15zR9zoMnDyaquDjbcVaqa0ibGnUUfV/p
0L4X3hBK9KTMFYppv7YLbmIHNF9lAsH2oviLprmFiKemCuFWdQ+XatkEi1XgW71G4VNOSM8mXm5j
Zp1c0FoJtWrH2N64UueVP/331PV7SqevSIiiPOwHxTzpdZZtbgUPL/0+nVl/BP1c/9nDE78Q57Y2
EuWF9wvSfE3EewDdAiY4/XuFAcN5u36wjNfGxQlAs4oUEQa5eMcl2v91Uy8HZMuJ6srZ10pAglI1
YBv78zEhZorKF+wikK1DAZNpSJGQLj36HEqFEfGDjGGP5fx3SrsOkxMftBsYBK/hoNDNBewjZltP
Vu6zIHTszqK7h4/kAUhlxy2jrd9erzQNQRiCg6lyzjkkeYUvShvlFKKtgnOFC3yaMbVit9rGGa1m
eAjjQTn0NOpywv8fcXyuQfHSKod1TiolLC7eyuaCV/PWSOSBUyuNpH8tiaN66Cog0x46ggIiuL3e
5cncMfxf9+YwzZbChPy2R0gzlo2YlZekvmyUlNEcH9ifcAjdVkfQih2eufs++IXjy4322NNpbHI7
xw5J2onacV0r51ZsmltUlOY21n2N9SyGo1Q7LIUUJncbGIVlMD+Oh5MQKrzbUiqVaR03WP8wGnVl
G8eE5IevDRza3ZO8Xb7dQrTW+X7D2Fwx5jlK+shFiT7zJomO1XS7i/W+C73zSpiIhUAtFXWdhoXf
fxcDmQGg6e0VE/Y2qQZzgpPe0NTUMKTC+KkYQPncB5krPIeceMwtsUeE8MxpeemI9CkxAehpLNMI
zEXpGeXBEORmuyvWSa5+8qfFmeuEwRmki8dQwiGbOxB0aEjQ37+aFUrVxFaat7YJZ6bPQGK26Dvh
hWu+K1mBWoCEDwkvxZlw35/pYQgMqeUXA2tXDkkXAGhWsg1LzcAkQS1J2V7xvmyLnMBxtFj4ioak
T80uZpd4BFxLKj9Dtq6rnTsR0w+1IOhvz113BozAn/U6W6VtV73GQ55Cc3V9+mkVk1JVVbP1GCfy
ItlUbaqzC+NYl4w/cyv5Gb4Q7Ww4WrjvNrB6EK+JvFdZH8vgAsTmP31OY1cVPj2k4fp0Y0zZ2Iyf
eSI0ZxtslpuLvbuHigHKpL7JufWvBh0TOGGNo16hRqGBpWZs0JnZlZEmd22yLLYfyZHxV1+jsYn3
266PGFhLuwgaDt5blVTT8WHWxPcC2vptEyL7cpJnB+qFeDBH8rM2hQ9WqAxH8elkqOPy/yMszysA
e8hAuTm6h3SI5o0r2g0QdE/l3/mTA4IXQLzuU2dbvo25nJsnL/PUdOQYwwNJeZjUtpNAu5R5au+f
phtBWCuPST7Usdolq8n686Kfh0/5xQ9GWBwL65tD9MQX2X0plPhuzOZN5d2UuAWNFS+3Yb6iJTt7
LfCSP6Rp3AQBSArefnw6H1tzhybrS7f1rneSCiHBaMvzsTEJFUKdvKLm9teVuB8nZt1xIPAVKEFG
cIs/uhwK2UYCONclTNoY+M87nvvce7w/ZBi4wu2Jb1ogS+sJ+LG06KbU1tBR4a1kobnnal6JPa1O
rGlOIzXpaFUr/EKn/AlN4NztFc2xNyp+0SO9U8kSgzqpMQeC92XpE8UTF6DUdU/E4ROyRX6Cx90O
4pFmLJBAa7YhRIon1CGfTrDyzq2GkHbggaUHmVdOK0FYtcSvXvzrTyXRidAe6AMNsVyUO5uk7Vcm
tDRXhwrzCXgxR9AjOunNo5XXF9g0eTt73XWFONkm6rIr0v/7jl4B/tLd8ykDUS1UWSz/9YFriR+l
dm4cyZlSknZV0GapAZpqH3bQ0WAkKOBKpXOJoVWKpZqScDEQrv20ex68HG/7/2Ol3kqpHk71g1lo
NPviXp7pI3sScjLriW9SL+VFZCYDVKvZjYspW/NQywfNKcrpCB1q3PKdxnMXkp/av1do0l7fHHPf
flZu1dvXCf0fd2D4YSyR5O9IgroTY7fGJxP/+ghXJM+QqXO+6//e0OvcBZim4A2u+xcPbGA5Q6zO
InbKNCWwk9rADlXDRKqB35fSr0DUkBAvPWK5/V11r+nFBf7z/yMzMoynMjJeef/cmMVO7p5mCygp
Mztp+N6oiubFyK+eCRnVtCWDMPdGJX6+JZv1VEuH4Y5L9G9noN7ky2quTQujO0PpMStxkZES71Kk
JVRFBPf3HOTarkTxc1oNOmvhc6e3BcY3hJ3wzI26Jq6zUdRV2TaO22d2Lr1N71L/xxqnzEuIWy2g
UhXNwgXJe6pIbPRv2Vvf4HcHaII58kvu0MTWDlsp9+7Jgq9VkFXystT3LCirKpahsTomfTkI4jUY
stGcBtj1Ov6WcKJgLHhQuJL743uTQNHokZpFhfo43kBJ77fgW9W1pdeknXt6AofyfyDvfw60EE1Y
Y+p42hI5R0Zk0slglf8tw/9h5xma/MxImwA7ThEJ5VZympqVhnzrH+vJaunyNMmK5VrJ/hZ4rJ2c
vohI22c4bXQxdKsf/oNLAfs5yM8tNMiBcY3lg/GfLdgK6FikA9r/JjiZF7RiZ+1gk7xPMdsEWDHS
WDP4X6I7TYLpPUme6wUMPTpS+mEFh3lcZC1nwDF0lk2/ZlO6dPkl9P9zgHEKNcEEfh5kMp//mKTt
zSGqr/wonQowFoCxvyWE6pIyFj/82vuwOnYa+ADfvbYB9Wutp+fQUeItcjpQU9oxDde0e1tO7N88
3kJNCGwUkuiR+JWoD5WBJj1b1CQHfdTeyYKhxJGDziwAsehWbAvjJuJ37FjqC1QnBeaNt+lZfgcm
JDbblvLvy3KyJeooBhUDbpsUhPRloZS7MJs/kmHuAhd6UDmPavE6nkh9ubnWh/eCl58gkQNkUQnG
DCLqZey3Gj5aJwPo4avpue4uF1nWwW0c0FxDrshD2Ei8HEumQwI4a2ylS5Pm3TaRqqAShtu8vJwj
KTFcJo3TSJMZWYQBikDUoY0CeVUAcZSYyIsv3Cn6nx8GnZ7YmErBGqV8FThvWRI5EaQwRt2oexR+
VSwuKDxHcBubJJwktRYMslfjcZmZlyG9C/Od+Oi80+Jj2zaVtbLy4ty5W3eOBo0NoWzze+52XT/O
HhaKE+rzLH5n3uW9viTZYvBJeIlIrwplnHKdRcdeH8qoKDe6Wi1BA3I8w6vPUA/eFkmdwY2VGPs0
FWYAgihH+/6aR1pKbHrTmBXf+d8P8J8ebE4s49ZRopuItDgYoY7blgoNDXzfLyBWGNwM6rQGQuCQ
hO2EF9TeJl1PM3iaW7WLHGcWrOk65U7Ub3mrNbYxBwqnx9Azq0edx8AY/AaCAq+9Rf6Nb1YUXh4G
ImrZeof5Mc2xl0bdMGbNLfIq6lJDzWqkyC0e9POuRvv9Y5ArX6BlK3iJurY+Gyl8Es9anQ6tZAHe
xx6iT4ujTssdFrsEPK5D4+VLWmBfSko71q84GWyLSYA9GnQXCulIj5de9vNnhG7123fJwK2F7f7K
ytZugFWWmKAwmhccQeAUIaosNJZQrgFExTJ0p9qMy/0rD47u9QtBTTLJ3GQVuoeNnLTqxFwTKv5Q
eXtLJpaHV2ywQrV9VuY67dsL4QuI0BGT6W+2MRFTfpWbIH3TdJcXFl4u2UbNIp4Vv88MXxHn3//i
g5MkaWuCcKam7PoKB2nfD+LyoylJkLO5IWcaRdyOz/LDwdOWDYtNlPIZGn6k4Icfevua4DINKPHu
CtaoLUSvtMQ1mUBbDI/NjHrCGV3PMSQuv2M+cRCWFcOXyMys/e5Gwdf8YV45KH+LeszW+FI0AzF4
/vmZnpnYHWWgcHQgUHjpIhfNhT2cIkqiLzym9dQnXDUepmrHr0zUlLecErYK/7RAqY2oi0it3OMp
51UF3Xcb9tESljSNFhBgy2P1n6h+rvPBQLFtQivGsCiIcB06kqdHNLw8HBGmUCzS69A+F4S7UHTi
khzpyHGgSE3d8I4TbWbMBmkfi8mXSIOgGXXRajqM4UmyOk+bOU7K0Fadbdn9yLET+cjo2/x6Jkho
omNkz4QmDdtXVQ==
`protect end_protected
