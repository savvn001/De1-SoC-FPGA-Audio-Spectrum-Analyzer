��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	���$����u���>C�3�
**lc�@u�l��ZoH���7;�g�(��*�f�^c�9�����t���H7-O��U�ꣁ��H��q�[�Kߏ]+��l�Y�+)��/!��5{�;o��ӑ�,#������:m�@F޴nK���:ohGЯ{,��ޠ��I�ܷ�4�=��AV���a��YǗ��g������-S���%줩6��L�|"ӯY��{����$��ZdqJK�^l���?Qd|����b��:sw����r�c)B��i�����F��D�� f�m<:��&[��
r�B~���y�B,�W�X�F��~�<�]t�TW�>g6A�A��ŊZ�|<C�U�{�NVX�Տ2�0�(��n�
�M������ፉ/}����E��xM�'��g	��7~0W���]TS���s�J��F��Yh�	�Wݭ���.ľȴ6k�
�2%��5�>��'y ����\;�+�n�������Ov�[x�B8w�/��)�	����5)�ӷ�w�#�e�cX�CU�,C`X���X�;K~@ h�ꝍ'�z���.�05R�*��Z�_~�#�{J-`{
�K��JG��HxT����J[����m�{)
��.'^�`�t�5�{a��֤kM���Lګtڦ3<�W!8��
umyvio�����XU`��ht@B�{�ja��B���M_�{z1U��K���#�Ǖ̅��G��G�D�!:1E��pv���j6j�� �E����f@yws׵����xς�0�Nm��+iA(��M�V�����*�U��i��2ɏُvL��zq}�L����hei�\z���}�N���6P4��-q;���H���N�I��N�h��}�D}z�@�4��G�ŋ�qv�G�\J3�ky��7GYN�Z\�B0���7HtҪR$��p�<n�W��j���|�(�����N_=���w����LN�4Cτf��R:\tL��%��~.�^\���{^{��$o䳪�1sLS������x,j5������5�.�J���	�j����ٙ _�MK���@9��g�k��b6{q��By �zV�P$}�[6�i�����ue�V�U�  �ܤ���*j�4�]�"�X�n�ax�d�����8s��D/� #�nxd.�~�V�^��ʹ6$�Ҍ�>��!���:ƇYо{B����i�[�4���\85����� ,y�Q���9r9Tri�7�"�����G�?U%�Ws܉�Nzޫ��a2�~%�b}��7�_�	9���o�ў���I==.�;k�y%�q��䔸y(��}3�.r@[U*Vh�qiW�L�&��:(Kze��y��\	\�Ĵ=�:���*��)4��|�Ae�yh�e��pM�G����S��c�oO����Y.��t�l�ܪ�k�J;��9�_]&��y'�o�<���T�%Sj����V��boWcI��8�B���G_>bF�H����R& �v��^�qdS����פ-f�c[�x��kD9a�z�ETom�[�æ=I�����.�E�]�_��x�
;�����s�C�4/�Y2ic�0]߉![@"]	�N�]É�P�0��` z��A�S����Q�W�>��!RF�76��+��� 
5����^sk�`9U圧���2�	��ށ%���i��y�	(��� ��IW�?r�R���a�p��[��W��iӼ�I<�E�ub4C�p���uG�he:��B��Ex�i�f��]zGd�D*jUZj��t���hӁ铖���yV����W�������S=VEwIK����� ���x�^�oكb?��`�B`9e��^��a|T�$�e[ҫ5f�W�|��k·&���6FP���7����[�3�a>gaD?3®�����+�Y?����@r	�U�62q�tv��	� ��H8(�]'�Dd�E�\���m��ȅ����R<;0�.xw;!q���U9������ kL;��y�'*S\E��U���Z�V2\G��ʪ�u�O&~7,�Ĩ�I¨�ނ����֜�;O��r 2�G�̈́�=���X
�p5a�U�U���p�$��ĸ��sx�mwӥ���A펄+|�c���G��F�k+HC�z&Ft\9e�X�"7����������b��k��r����[c�N�����EB�Fj�A����P�"��b��9�~e�R�%I����V3�ȩ��˙y(�H&�n�^h�ET���D�}{=��&�e�+�6���6�e� .�����.׀�⁻�B�LM�d�s��Ɗݜ��=Z�3:�������0��D���**ێW�JS���ۋ��|n�n�Lan�Yڄ����vHS ���B���CŶ��&x�rK����/�Abn�:�<l����
�/�WQܭ��%d�����"0��E�����c�N�h�[e�S��p�X��$��
#�G����}*�[�w�4:��~?H���,W��r���56������:rHl��M)j�"Ǡ��]�<��&��gvud�+az
� ���T��he�HQ��_��ʊ�5Tn^�bU�8Z�±e\����6��v.��i�I�N�_m�B������x��܁���Ă4x^�;�VA����l�!����|N�R/����Tkb_'��M��}���@�(�
��ĦZ�ʑ@�J��8��>#�h,�g�ύ�
o���@�o��N��l#6>a��G�L�ͣkg��9b�rʦ��
����(��En�x���Y�^��5F���AtQ�-�8/������X@�1���-r�Th�X��0�������u]3��A��,NZf^�.o�]q��}�B}.��Xc��O��uM���C�������~&s�Q;G��|�Ť�-���	]')6�&b�@�Y�0Nk��)@_�>u��d4wLč�;3*�a�'5��^��k>��7�`�<�w?&�ΧdP
�z�鳪.Kbl�n"�~��x� ���_]����i���[���H�k1�/ƍ�g9��5�K�U�vwYd��\��ί�i�F�G����1=���@�}y?Ո��W38�2O1�"B02TY�FO3�~���lmz$��r�!�[��a *ĂFv���;e���)���rn�����V%t�:DD������1�\+�ݽI? �Zɏ�]�eUo ��c*��?�8���9�>N�Bs��>:��-�G�|ǖ��F��@�6g�f��S�X��b���c�;��L����J_�k��	��|��x%�|���s�&vyŰ�x������/pZ�3?V���@An�O�2���l�(U�
�#����q(Y���e+Q�2*2����&��=��e�ƌ�(
X�\?����<��Z��=H���b1�;B/���tq�0,��_��X���l;�(�G����X�M e7� R���-P ��p~ν%ŵ��m��[kdx��V����b3y��5��bRm-��1������M�u����6��4k��$`�n�%Yſ��^eJ����}��$�a2v��-s0��T��_o+\�VKB���L���_b�"I�\���^�y#r�$O/�6߆��8<�W�Zl�`�Ā�s��a��
m\,�YJU~���L��"/0f�DOӬ�6�3t���C�T|���m%�i�aT��������qK3�@���5=U�I�~*�+��g�4��EhW�V��f�+ٱ|}�������3����N�z�d���_:�+��RP����-��L��V�|�3j8����R@�a1��P����O��8�1��3pȞ!���Ԧ�8�Q:��^�4�]T���,��+��m_f3�N* �0D�����i4�3jGm;��K"��mB/[)E�7vG˚�/Q�h�z D�z��9q���	�.m�����SޭuXV�/n49{�q!��5L� �A��Y1"�A|\iQ������k��ԭ�p?��?�|rP,�M���Ʀm(U�xx(,²�s�9���z�r��j�x���h������]#N��O�=��$��u먬uo7)t�^N<X�d,���Xj�H�6h(Yd�X�% � �㸸�G��Ӆy��[�i�ds������&�-#?T�Wd�.�+��VZ�
 ��Ï�3M�\]��s|A��{	B'"m��|6*i�9?_�@ �`�ϣV�����sZ�TI�]Ԇ�e=�y0�c����Rؑ�7͕ݱ�(�(�Ƶ8O�l���O���I�𠆦�|,v3�2d�Y_^�m�F|��d��B� �X�JX�o��w<��+�h����m��ݐ?`뼧�Η�w<k������,��v�S]Bإ`�N�p��>i�"�)^�&���ml0>i��kϹ]�1m�c3�ڧS��#�&��?�[�F��Q�%YP��͡��'��m�WNc#I/�=Ij�+�����P���,dy(���@t���Y�Rң ��gA����tu�q�6�	�g*�"ܿW�ދb��$n�Pl.B
|V�6��	l�}ya/~!u0�O��#d�@ {����IB"oz�K�nGB��r��3�f�.�}�O#�BX�x%��f=}B���c�hg�=��ȸ��iD� �N��oډ��z�ث�vg��4ه����������)�}暍��-�1M�wc�Fw���Xz�2�J���>��H�"��'K���kY�������m,��(����[��4j���UN3�V����Li�x�"U�O�|k��t���g���@�|��Ѻn�\-2.��ݧf�uW��#�$&zMl���M	�T[�EƝZܲ\�3<ĳ��VP�|>YS�,�1�V�:9����H���hc/	h��m
���-�>�]��H=I��C�J�!1n���L���᲎@��w��V��v���\�pTN�/E_j�Ђ^���s��",y���y�i@��l����f�D�,1�{3�7J��]?D���\,��~�h.wӷ�6GUT�L#W7P|���#U5Fԉ;~��mY3�jN��(�/a�b�hΠm�2���r�W�Ȑ|���#�s�mv�`�nKz�p#�����<��»{&��A�P�;�
M �tv�ri�����u]�/�����۶l�D�x2��Rs�o����V������*�9����,���{WV��6�i5kX��{�#�vV��(��!�_1
�I�M�߅��pK��XD�m�_���4��6e:o3\]kCn�;[�sd���i$�!��e>�uƮ-F���23U��]���p��6���E=�"���(���%%4�X \㚢�*@��쥁���x�P5�|Ǌc%�ɀo�������~a.����봇��o\9�e@�	i�g�DV��6��	�!���p�dv��\�����l��Fa��X�Lg��uN-��d��Ӆ(P��yAE<i�����8ш�u���JI>e����)�5Ш�(��> ��{�T���a�҉�]w�٤��� "eӯ��,�]�g�ͯB��R�_����8����H=t����_nA��R%��y �B9A3�:}s{��Fq��#YU��;j�	���Q�	�"N6BP7ɚ)��Z0gY|�[�!���)@� �xQ��[Cq<`�]7y,��G��[#g~w���G�O _�ѬgT�1y�g3�l���
�x�������:aǊW,&�H�f���0����V6�i�Sa��B.h3�$�	�RL�0�����������*��? 9r�G-9$�ctK�Ϝ>��ofw_��&�i���NJzWm~sU��ׄ�D���@��hS�g�2�2�T:#Rc�ܛ]Bf�uJ&���<\��P��唡�S�R�'�%�x#�����%Z��M�3v��hI��Ͽ��5~š8@��k����`'�3�51��}  ��ET��q����I>#V&�/%��~l/&2i���3�D֭5P�a�'NoZ����Q@�YS��wO��׻dC��Q�q���:��X��8E�Dh��+'��a_t��^�ؾT%`T�=���GY��\(���9���ͣ���o�]��5W[�5L�}S�f��wd��N���Q�$|6�,�����;�T�~��Y�,=��k�ِb���UU���TW"J������2��+�W}���[+y��ݧ���IXZ�W��d�����3ޠd�=�m ���TW��'d � zl��Q���Y�㪱��S�MmPUi�G����y�^��ŴD�xc�g��|�@�g��+ �6v �1��h#��u&Uv�X��g]u֟��|{A���F���&��Q��RN�0��-��>)1	p�s��-ϦJ��a���z��'�����b�b�GH5�w�o 
��/�M�ǽ`�|ڞ ��eÇ���tګ�xM��[Ct��&c�n �=�R�;����p�UR��笘_���{�ә����p�N�*5B)�"X��q'7v7@���7sW�$V�m�W��!s�:D�}$�W8����Y�k�Od׿r���U����j��K�a~d�Y3�wa����|�,�^��3��f0h�Վ�F��d�{)�K��x�D/�W��X��K4��@{���vN=��$����[��	B�R��upS
B��z4�N�O�+�=�����`�6����Ccc�F��S�G�6n���C+�1��{=D��d�)�R:��T��sD�`�54�+(i�f�2^/����G�M	`��#^u�y�tM'=-F<#.W�;r�����#'h��=����]�v�D�ŵ��A�p�X�)XE:�M%s� #f,�=�%�����ml!"E}/Lpǂ�6�/Ugv��P�,V~̫)"�B׏�Z���j����:�V�/�V9����E*���:�B܋t��غ7n��ҵх`M̓r�HŬϡ�����	U�p�K	_Q�˚�{).�`=;�<�}��=�Y� l|YhC��C�����wm<$�B��`��-T���r�;6Hm斈2��������idM�l���qi�=����3a�
�O�Qr�ԋ�=��������R=q�p���.��(���l�b����V�>���͍j�&�������@�vυR�︣���f_uV�b�h���\�*���k�:Pa����#��<��D��,�d�P�m���
K���0��ma�Tk�@#����uc�9_1A�^M��E��t����i� ��X�7Ҭ7d1���c���xv�S!#�K!�KZ�(��A�����r��O�p[��x���ݟ�~]��x��ޯ�X��uBuq~��?/�0���r5��ɩ=C�%�z.4�Mg���]�A��Ʈ�Qeq�:�q�M�dٞFYa��dZqVu/}lE=D��]��K�e�� ��h�l<ڎK��E]�j�
ل��w�L�ۿ(�?M%۽�mt�M�W�N�-|��A�m"�&^ �`jl���'ψ�o@���Bt|O�=�|��;����E����a+�iv�$ķ}�7"�SuMt��U��$Ҍ��;�Zr�:�M04�)�P������zx���!����@�h@B#~)N����=s��Ě���V"�(�����,�p��0���j����ޖ��0y����ύ5e�F��}4B�Q3Ux'^�=1��YReA�ő�e�i��;FQI{*,������p�L�vYh�E�Rа�