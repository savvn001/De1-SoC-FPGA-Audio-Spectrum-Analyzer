-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
I5E4vECuthCc1/U2RXXEkXmdEE4LYNTUgYEgmfpj35aZVMAJ6v/9MphdQnShvi4w75XF7mg4zscb
wPu2fB6RUY+l/xAfJDzfPUwjKQ15YYm5wQ8ARJ/C3jE144OlbOtPA3v/FVjOVdCUFIpfdkQxBboA
kVlr5q+M17j6wa2ek9dLclagqVyXklLj6DK0uhLYH0AqH4ZCB1rUBl0wtrSitqKRgW6AIyKFLvDC
QLGIWRsMKe34mwmun6jXQp00pPH6VpAU1M08wZTpec9cM+1C0ZuJEjAubsqlCU6bBRGJe3lCg0o3
1S6528wIUaWc9EUaHMMu2UdhpOytvmxX+rlx0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
9qCulY8ULcxks/cC4KHwBy/9sBvLsRVGiMpYVY11SziTjViaQLiUOWPtFtyAlJVqtEOlWgXCTrnP
uzG0ufF+TNFbjFh1P13dOZInbfrvA7/kp5eF3y/00VCZsqfJwPMhh56f6DmiP9Y94t342YAh7SuS
JnQX87/nizzpuRMBoS0y1cjejY+8YMHZ9MYlWVM/bEbG7UQ5X9nMy3G8we/zeAJvbGbPZVGdzKyq
mE/JuzUXr93c7FbGvfFxqJ0uR9Kpf6hmSV7XzBcqkw/Uz5B8Z4gSGWX5GVE+lMj1puQPOjweXpNM
tGZnqus2xTaT/POiNvc67Yg+7DHJoIPrpWEqefat0Zgsmv0mKTns42oXNOs3KBaueTHVZhCzda6L
quxmoT8CkzAO5CY5S62/8MWy9Yp+wviHNzd21SvoL8TP3vgUbvezeqLQtj95ers0CXs5YorJZRfr
93wdltDtzfyFzh7b+PX76bZ2E24ROcpOb9JLqKUddbHixL+V5D8zxMGcjozOmroFYJ8vNbaqJ40n
0QlKmgQRtMOmtT4MfGgUnXZzTKwSAn66LKWVyLOsnu8agb4EVX88K2wWcCF1ej1dvIiX9UD2UocZ
zV60tmCetqo7OVeD1sagFiib+eJxb6uxwdqSwvEdhz4ZGD3cx2LUPqZ1mFe/jt5qS/o0myxlu7P8
BaGVxZxrqpVttgYH0qrtvcRMxjbN6ttwuvD8aWGGUOJtEtl0Jc3FJcyHUeSwpFsWHIb1ULbvQC+C
dErCuVrd/YeL9mkPyuyrTJbRvgCf4QgYgPKp0tb1HTxrUIufIZj8td59FGSSb1SaCSYCiXDwT3oH
wXXw4cAjS44gWoJSR/exaZ1W3CHaSQ4Zp59XvJjLRs0BqLXZ8O4y9jRNwiDExpjZkxlhu49zKLXE
tMm7R5n+XALjq81e1NUbANaOorVX48VPRrV+e5TY2XgBjFsO6dOXyVADL297Xtl7Y+06GHb6jejk
PUo4LwbAo5VewqEmfyb19OUM+XeRDjkW6rYJE5AuyU93M16IkD8NZYsve77dLRbrOtnrFKbbFYCE
xyyGf4lwQ1yVwQwx2Yks/W+Dtd1fTFqcGJyMibY0Ekduq5k9N+tRqCr2C628HcT+zmgqE1br0GAI
uThDV/IbLNRlUYguh6NziGm5w1aaZLGK6a5/gDyeyU9Ruc2rXtAOJBub9TYgBOvR7Vrd/EB5+YNF
7W3UG28s9DQnGaum0e4zRyIVnYC183ejGIUSi8X8lU+CwDUHVgj2IckQZTsHkoFzBtr94QF5UPMY
3b5c+SDgiA0FFwie3UzcqlBiCdrX8b3vH8dPx90s7rQND2S+t31Rtumfvke1YeqaRPEtFYQQdt43
1g8YdYPiCWvVqXiByabroZAPC59hmz6fmn7l5SWghCQQENvL40zooHTAj0+NnSHmXEvQ1NtyBO46
6j2mGDPyiYLfj2GHH5kWah7dhVwpQ0g6/Rr1P7ds4dhSipqpSQJRFYfl6G9iSq9wW/7guVr+CMrD
2XJxUikXi12gJILGU37d+glFz2RSEW0j3U19w9o2HUIyVmoBDxQSkAsqLIBu0ASZUihOVKnIzGTS
aMnijA8hLB7gBvInmyXiipCRwMkgc6c1/jVEDrzXMoodmwwLRhTma9hC18x/CdOzUUQAJH2fJC2K
hBs2Zrq9DpXIWNr7MH4atxroVM3Cyv9l7o2VpiOCnVN1sMbLvPGlaG79jzVXc2ryIWIKGcMFFPZd
yAi2ix8i7UORy6EN4I3/plQntOefB3G5pmghBLWzu9LsHVTly92HVBv11K5fqOPR8lCh46iOxkYa
RKqTVKkJSO7VRTExM57ROd8X4TY1FPtYREK127y4PzPJ7PJP5BLL620kNXyPs8VW89RZIeW5RRx1
KT5MsJhXa7buCMHdewcrBPYHwuhrDz7Zkz47JZuLWEQfF3Q2uHm68l7Jm14PgOSCnllpgZwaMCq1
/YHAeH1tsatQKjJ5etfezKO1BWdc31G9ProKmWBc1pJHuTQezjPJVaoTWiJIAlDjAyew9NakuCDj
d925v89U5OcxXFUOWzW5wCUeAdDsG3UgBXcT6q/gzBcoKTw6DG3a2zYWLvPrlvtKtAPufo1aztpu
JXN9uDup58f7X77Sn0oETR255E6d2TE+Bvu9tgApQSjdhWiteSt6LWostkUifjfDqJvAls5po7CV
k6+gNxXU4eymELHCPHaqRjbILa0adgFaXptpS+yVVwh/GBPT+Mv33Cr+65MO3LML/NmyZ+nzfTxK
9iXg3C8MiAuxtozLXtgnV9ec8C1ON9DnfG/GvTGbTVx0PiGRRCAu7lPIHTxVNv7Oo2enxtHvVeZO
Ngi4toACajhVqOioHMJm5TcCJLlx3cOVPPYvJ80jf/Qoyt5Wv7Pzrl/+Wc1KTMaP6wiGnSZbgXQe
bpUwvP6dKznSZIt1EMKcmttXD/zzJ+4IyVmy0pWdIrMCGJRulPxAVOLwpZB2LLH6VZgzbduRyxMV
zKF81Tr5AhxdoyiNi3O38jFssFPurHLuEqdj5TeroNKDSVwll4SV3bz++rCszZIsNW03Gk7GvIiJ
VN8OVlxNU9mfxnO/Yhrl6+jE9KpZf4YjCTxt5uUzy70kaV21Ml/HbxuBQIbgsz+hpwk1zxEE3rXo
VgalUH6zwZszsA9lYCelA57IdhTciN/KyWzoQ8Ob1zwqU31iNCIJQ3er0ICFQ2YxLJWO1Js8cnre
hkMvLSQcQhwrKDQoqO8xlEUQUGbpGT2vBkxByuSGSaxD3qskZnkshUK6HCfw65QIC1+G8ubAbsLj
L5NmcvqQQjltNTNn3UTlP3F9yvUlV8AQ+YcOoXknl2CDTYB5xftst8E1qNdZjmduhCwW86APgtrq
4tmRUaSEEbUtzhHkGVIONrONlAkAs4ywjLlB5l7frsuno2QjOdq4vlNWolFdFofLJySzUV4HkOc+
RLXLW6KvlTTqSRDxLvTbFaxmQTVRUllqAzRxEAeKN5QCdRgp36FfNvm9Bp/hjGHKZljz/jtZfwro
r0Y774B0sZz3vhMc5WGWv084+Ne1MC0/36Y6XDPwrOYRk9gvwFzOCfHewluJulwOswUNMjZwQ09F
MFyNQLAulIC2+7OPcdgdeG6zWI9Z3SoHsNNiDpcojql147xXxVPlduC2Hev1BZbepPD17ksNeTFw
Ms2KmSpbgIEaco0zrlWqjCUCc7dSpVz/RDurp0HPV967hqCowrU1loLUeaTysuIea0ykZyMOF+Uh
m0r5OaxJyJRe8VyTCqX1DY6buB18mUFgcf1YP7D8W/K1r8L86zo2Kqdm/1iUg/j+zuwbUiAfwZ/f
600ewQzIIJoDz735+03NjVa3j8L1iC/JrVCYciIsuRI5ovy2AMMY7UbgLzsAAVtEO4+uxR0I+vCm
RYgBYQ3yn0/QYNWdAFLhO+UyL9SNlUc8PxevXKn2otrYhSam3g8ZHJ/5XpMOKyTBih/GB46jL2Bw
FANrTi9H/x2giXHybjiux+07V91Z0rG4YFMOSyImUWl56YNYGc/Eo6iXIO2uPqf5ihhrM1bSBr7a
+A79NMRUakCmTT6/+LvxAUMGgc+bLLvIYisRhNmX/19jroErEQlN2WFXqDmMcIMx0HAiINyYeRs3
LRjf/82NqPWAryfDOoeFALDrDqH1DMcT/+L5NkFzTforLea2pdyqZaG5eSQ95mJqmkGFufmVcYUG
EeEbz9w2IFcjEj4f+SaqIbh19FobFhCl4dxhiE4grPtkkP1cSgLqRdPdiikwxOYPsPBzYIDXcyfD
rYoyqifkAncWynlwRBvWYtVx2u4WRbtlxQYlZXXFamwuGsr99R0faB+kpTOCTU5v2DY+cogm+t8f
5rihDKygi2RHng62hH2UbtVttBE4DNawc594Vj72XYAjezOjXhxcpG2HrZyf6KOpg3XEI6bL70vE
BCPyJMbVCU0BZKynPZriLaSEM8iFFFQyr4kbbLg8cVNIXG0iN+l89ez/zxXFJqGfZPF+cpFNllc+
TOrGJ0dQAckUZ+hk8+Ho6IlcaaRSOXp0qxTpHzBMdi7wmL/xk7FRVq/7VorofcQe8Oiq0PnDoqM0
Osnw0AUf5ykYt1N1YQdQlK68bjUP8nzGr2+F1+VFXEoMJsRbQdTjKOEsdv6QXFuGarEU7RLrcfh3
A87x3hVZ7sRVX5WldtVOkI+lYZNsz73aN9HrWYclIlSgMbMgpu2D5PH18uVew4I4Zy0Dz8z19R+8
0FYh091zkGPHdUq3X2CzHOFN0Xx7thQ6DISZ4ROJa+ktAKNcWxN3KB4cnyK/Y0mjf0Z9CzIDuEik
fGJuxFwncsi4BU0PTkXJLx+uaxpwHJm5OmW5rAtEBUOue23LjgWga954kHd91AmehEs3ikRgl0gk
zzm/B9NNeMMuqTlXhBX31lSv5twIn3cV/7lt6UxhZyfl3ufrtLGWPngQkqaRNpQttWdmMXv5gTuz
q9SpYmGKBNsQfkY5aridPVJOgbJQYk+ZOXK7hjUepN6quPzzZeRmwH3RjYN2jOoD7oghnYymjaH7
FmVlLVr31lAZu61zHXgr3eSaAX966Cu+f1kMb0Dt4+0lqsXJ/NUD+grG0odwYvApfBh/v3CWbVWe
uZTx60nF4dccQCjBRynq5uU4E2LAK/BFRs601lGixTrYcNd5A2LMmH+a4+uAZnOxFH3HWVULVWG7
B5pYRoknl5G8aHsQpKO0qmlMuZtT3NK6IfhRKGyqfXLsGbR+myhXwvE5Yh6pQ4k4G6zAtUrHbMbZ
M0lGnpJ8krEhGKswDSeuByljeHeJq6FMtMpmuq0zeH8iVF452DHvyCfHzHupiZZgmPGYEMajbAYJ
fSRdEm5GOkEMz44SwzsY629T+qNNNqT23K+m7P2j4je96gSVqH8q5ZP/akPVnc5fUGricnmXD37F
SsqoSIRRd87j1EqEfP984nK18otRO8iEyp3VOame0aeGiWQvy2u8nLUmWFa1Or0d8Ie1wn51iJo0
+ZcH79zfL/G6Sj9WxHceTyytOjqlM/C5NS7cAvbMNbCSl3Jc3bL6JFBBhKUWdgkKxjckgyiYtb/J
j8kjugDQuouOWLRc0Bs6BN5lazcgc5yEJ5dWBVLvemsMy6iz4NHelTaSv0c7WzTuYIfL6A6z3TvZ
iATXQxqEyXuG0UmFtgyWCECnf66DtbsJKkxthvGL+/6A8Ic9G56LMKAuu7HZRvsxzdsH7AJcF1VA
S8NUB80eXmwSzXJ+TPVspK8+qi9Vk5//LGL2NpjatBOO7YF5iAsJ3a7DwQXtqrNQ57/2bJdxZNVr
hV+aT7OdhY14rjV7WqqLkEmNyTqkXV3052Al2Z04nqP5cZnWR074K7TX/Fdl4xMHeMa6R9os/qev
wsPlnvAT2GuykGReklQaVz7WDHpOZXE9gdxQUb4yE2YKcTpVYpJ4ytyFnX86sgVehpbggy5wJybI
HzRhDpTdmjbWrGUSdvKTDNfODkDKHhRdq2C1E/cvP3vjTRd18gyrsLD9TOKQEhkDFnBmA+3+Z4zG
IAF0WWm+Nna9QRggigAngUIZtKCVlRfTbx+h5/z5EeDwD1DZ1FedRA+3bt+AoKhUbZLpb5H4+cwR
YYA80nMFXd8YLiVBGOj09j0gM1eLC18z686NE6cIZxdPp0JUHEw022tv87sLPiWiVK95YuupFXvL
1KQ4Wv5NFEicBtdPQDH0TeCa9FgenSGQwBYtffE8hHj2V7NFHGQJ2WUOg4PSdqJolqaJcjOSnnYO
X9OXGkdVV0+/ZlNKOwMVpZ8k7YHSOEv1YDpz8bpZgfZdEr/ekP1HhWWHqqpSfHLIYVs829mrPW5b
4Y2Kl94iK7UGU7N5jXyc4897vsU/pukkMfVDH76OFVue9MaswTv/vdNA+Xn6Tp6GGGikEUyrFwds
+zBUAx4Z8MhlD0U3run8FWWCT6FmRkLApjLjfp2LLYUZD5449mb1xNmJeIoK4Z53b6ES/VBB1j8n
7sPgejDh5GCozDqPoh8hYLFJQiGx9tyM/6a3hds9OIB4rXh0GMfnvvMZXy/NbfW0ErTHX/hn/zYt
xQ97YP1VYr+vdyzPOIQbUKCjdrI557jjNbBdzp216qet1rCiH4iiKITmYkujWl6FacGkddbEc76T
ajOEVUWKd0EiEElzlvJRJ+PvS7Z5KHoi11mVl3nZNa9ISL5zsEfMTPeTVSPrqX4TM0GLmWCbMELf
l3Hy58HqIgblO/Bk9hlOIF9n9qgO/LNrlra2tYN/soOyyGUUmBMZKoIAILr2v5hZszwnomm0hGJM
56ijnY/BInJZrs+tTPGFggLbS2BRy4vZloKX6nGDF2K+2XSlFZlJnuqzJu2p6poNIiS8NXE8GZyD
5WV+4Q6lavuDmc9Jf9Bl4UMgcwMrZZIzOjVS/RNF1eMMGB2nysKmnpUSpCQkGYmJjbp+L6grKGHx
eoEFfTiR1pJQbCmrmsEqYhb1yG/4zVXnyLMuLzbS/9mkswPhgtzr83WBQuamGGJmgO8mg/e5JpRm
qBTfBxgFcrruy1jMLrctgR2FUhc7s+VmEjL7FklTtqpIVm/r8EfuWOiFC1EGKrIlkxi4sLQKcN9E
dpCjUYxlKzm5j1J46XxiCaOKO92zQLu4cK6nHS55Vgw4sF4vyTJnujWDCcUGg++DvFSFbt2echrG
O/lq1Eeq7ugCuiW1WADt/btWt0zxWrFgiDtsmns/dDxL/jIz9Jqnb/kZnev98KiL3cXzITwbY0Rh
hqk8VwElnAckhahseIPWBqdlGv31WRKRg2nZOe1y1ZVfFcAk6d1g8BAN0+gZtOdHJ8q4Y5KZRk6O
nEKeamCDliPljEPAFTNmvd3n+mYjvec376FxEgNKPQ8DPKbO4kBITXygryv9qUvGAIx2z8U+4en0
ISvp0Sdun20IGwQuXRN5VKLOCQXeqhP0VPUYiOTp/Sy1i//Vkx5hTWqTv/ngn8tfpbU6e2FEE0Xg
RBtaaW43afq88FmPiiSLahJeuyrVaQXpnHxKXVHaI3dwJlxaVLe4VySNIunU2VSC8/WdPg==
`protect end_protected
