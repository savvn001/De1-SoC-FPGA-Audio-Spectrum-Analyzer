��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjH��mR�L�J8���`	774���%�<���/�0+�XP��1?��=bC���xk�J���7���[�P�8��h�_�$�[0�^�"��f�����"wd��`�{�ʛ�"F����8�U#�S�|{2�a�[v��RhE�Ý�;"9�9������<[Sh'�/8��%�(�A'���-���^����H[]�3$i�T}<�zo�+����8��������x�H��#ʕJ�@ҽ�ipP�r�G���w,�RS"*����SB6 )9X�Pr������ �[�d8כ��
Ng)�&c�RO�<�p�� n��V���Dm�G
>��8Vgk��~`̦��
I��^����Y\�\A�k'M��\/Py 
ҕ����uYH6�U4�f��Y�j�G�N�����8ǧ���De����ߟ��X,%(=� ��R��,i\�)�a�2S�@�������j�)����u�R��*4�I	0�ɴ-���Z��<�:ɧK�$N��kxӎ���\1�����U�G���M'�f�����"�by�����d�W�T6�;�Hl�W(\4��]n2�H[`��m�(�����pg(̪gv�����r�g;څ�c'e�%��\5KU�I����3[V�Ρ���ʸ�X��&�ɚ?}���1��=���c��&�@E���:���j&/d�3I��8.���!��%���|���j�������}ij=#!�/e�lR��{z���¯��J�h�����C�5��¦��Z���-��%�j)�"��Vas ��ȫJ6M/v:v!����?�*� M�d+���M��2�N�z��x��=i$�A�L�K�(��l@���=����+�ΐ�
"����F��-�#r�xc�!���m�`T O��1�j�`{��O�)��}\���r�-X�䴟��RY����m�ϥ�>�T.���x���yF@}9��m#��C�1��v9���\s������H�T�{��*.�X�~�*ٹ�|8]f=5�˽�@�,e��������y�4ߌ���LB嫼��Q��,Y+�c?�K��R!8U�?ߌ�}�Z�3�&'�~��ɖW�\�x޷����o��Z�H7W�"�6���j����M�����`L%.Z���̉��l !��,���h�ׄ}����r�q"�ܭ��3EhY�]�[D��������-�2�I��/�X�J��\̅��ٱ#�
�������n����$*#��� �'���H`}���X*�h\q�F�_o����XFr�������?lD�VN��u���D������ǟu��޵.T'���-?�t��-�M��tڎ�����?}u���)���	!�6$�5��p��k��IL�"ZuIb6����D�ᷲ�~�Q&{����@��ߥ����,��-S�83�h�;�?��O�Ox�F�g���^�ɥ{ۏAkF�(7u�V��r�Ъڬ�� ���a��ø��2Bs�S��o��W���x�a�X�9���WDf}��X�w%f�{����:��%��A��>�,�cl��>�����V��w��[��%'��Հ4d�H��xs�Zb�E�~���@������F���Zs�cj}��'�&QҧOy�_��k�mb=�c�D(
g��J����\�˓(���ކ����^�E��B7�)�L��qcWFd&-LA��'�e��]�5��;�\G9�����J�ִ��a�Z�+ZN\��T#}�k���O[�ILtU�SI�|���?�p�e���ш�fZw�5 @�&����8�%���]��f�@�ĺV��똧/<�'�O�v�mRXH���N�ׇ֊O7n�;7����PHF$�!}N�ց���i�V�[�ѽ7"�O�M}���/ "[:Ũvo������R�ϣ���]�8=7)�\(u�}TO��F�YH�_Gzg�
r��b_��t�vE�x߄x��k��g:iv5}��1�hn�cO�(�H��8�'%ӻ�&����!��[H��B:xMP'��SRw�N.v�����2p��
���L��\��p�l�?V�y�*�喑܊M�MQ��j�J�m���ڪ�O܅ub<nY[>����)���51:sUe�૝�{���8��3�J�[s�T��v"�0yQ��̢}	��il��T���gl�K.en|8�5�����D|vC���e�Fa	Gm��V����T+���I�-X�|����z�ai�ۯTV:?���R{j�,�T�fL:i����*��QH��$��\_j%�崗*g�أ���r9��K�j�jPײ8������1g��d�1����2!;v��y�$�oȽy�?BI����eb�4��/
g!�ݣ�;-�0[�n���>,�8O|�Pd�Ee^��RNci;�J+"�R�eH�����}&5߉�#Q�����B�a(�7�m�� ��X̹M	H�MuE���|9(_�vv]�mG��H�6��{�U,����-�Il	�E� �Ԋ	�C�2j�|��~u�w�cȋ�|�Pw� �X�	)VPy�]��a��Y����QT(���m�C����L9��	'p~A7�K���E
�k��L�7�ӲT7!/F�j]_��(�4�\~'8�݋p���b���H�>�l���n����ܿ���\]%0v�KI����@�f���<E��r��D����$��1��2?o�?n.�-�zZ1k.YA�r�3.}�r��Ċw�,��}�RX5"���
Tv\5�/�ω��6��\G��;�����2&O�
�9uO��Y[˪�*Ao<(.A!�1��^'���/fM�L�,��5r-��1�>�U�V)�e�E�X_�Vr�"�ݵo�V���m�h�p�2����Aɫ�,	��7��uy5K}ե>�	�l w\�	��Y� ?�u0(��Y�9�SdFh�l2�И��-�| �YeHFy��ܭpE���k"�/��E�z�����9�ؔ�Gi�����(؝j�~eU�bG��!b�����Uq���������V�R�8���˾v��I��������$�K��$�C�ݭP3!������Pz;��T�pd�eYc`1J����ȔN���\k� ��ït �����ؙ�cQ�J�T��ъ�oV�:�V�_���&fS6�@7���-vI�m C|ôįa�\�) �q�ǭ�U�؎�S�L�z�WV�i�z����cO��~`W ���/��-�Q{W3�;��_E0�E��p%&�M=��Z��}�Q���`YoY��ǵ����#���f��#%5&��~j2���
M�<�r���X��{��<�Щ>Ǻ
0�[lV����65�EH��MI��X�f�첛�
�\I�W�0OΧ�x���s���;� ��U��I���O��_\ۙ����<|0���<ª:��\s�-���03��:H�^O����DǛ��ykfk�>�� ���o��� Hl=���v������X�/h��7'���^�3��7O���ɦ�_��/��@h�v�f򪼐o�L}㻡��
f6����6D��}#֏�v�,>y%V�)���;���9I]D)8Y�}�P2�YF��wJFt�pn���6����y�a�EQc�����1�}(a�.�$���і闸�(E�G���߽�kR�ϓk���Q	����\�_�X�v��]�V,�U,��I!�Y�]��ur��2�ܕ��`�ő�R��aOҩ�J���1��:�4�/=��z�κ�Y`���꬯y��$�K��8��5t�h��b�]�+�d�|dX���Pϑ�-c
!<f
��&�;��r��=ǐ�6��M"�ӧ�@��7�O#���wg6�'�'�cM���S�lೱZ{�]�G29o=�2t���s��8h�Dd�>\�i��W��CJ�h�J��i�(��f��).ԆZ�= ̓�'Z�KѯV�9�u�v�9.��2�6 �X,C�w�e�����7d/��lM��Y|�pU)��`�4bW���q�+�}�D<A'+�]P����r}�E�p*z]3����l�,��Ҕ�LC(�=���\�a��|,����|ke������?bg�t�'|��]tw#�d���܃Q��6|����R�6a�p��J��~��9�%^38���u@�,W���s�R��Ŭ*�=u���1��Ox�����̞�w�(������E�?����H�ӈG�E�c�t>����׋��S�\w��B�%�� 6��kB�W��4���Q���6�C*Gq�[	���Q?���>hVV#OR8�-=25l.�Lo�AY:e�����M0M�z�ܤd� ���x#�$�w����|E9� �����c���ɴ2�8ѱv\�#�
�8�S��SZ���ң���5�d�P6-ӓ�cM?�r��0��o�LS���8�PD�Fx]'5J�a哀�-�D��Q���r�tf��|,0 M� ��d�A��t���}5�9�5:%�2�*�ܲZ�+}Z��Dv�g,�x��#!#nH�Ij��4�D5�����ǲI���;�J������6p��m�FB�@����|O�7`��C��7/Fy��G��H�&�3�(MV�:�f�C7���!��(uNQ�ڳ@��d�U��m]�ۅ]2rA2���`�D�T��+o=0��Tk��A�X���W��o�Ԥ���χ�v+wWt���c���W�f�]��?����R��7� �:׶R�.�kk�¢����=���+��J ׍��-=��?��Y:��˩�Uv�����s�hR���"��"�
����5�AU����ái��f��9�w��k{��&�)���,�|�l�_[��!pQ��A���	m>����٥-�l�t�"�/�%櫛ړ�n��	B.�3뾻D�������#=o%S%�+��cg��@{��bܜ��.⹏�#�����6Rﳇ�C�$����9G��G�jܶ�4]-o�����ޤ�̈-��d~g��0�%�{��н��f��+���'��w:�&8�W��MD�
�L���J�#F��`�șSݛ���m�c.ZY�NY�ۏ�{�q2�5���7r�b��M�.�ن�`�X����G'Gk�4��*mmNצN�y�D��P}�8$�ڐ܍�Mbj���/%�hR�,,�K����/;����%<n,��<�j�� f��~�6T���B�݋�Κ��&�Tm���,]zz�4F�����6����)GE�l�\�ej7�`�J.�$�F��[��	UX�i�"�ꃧ/>��IJ;�+fI���Nn_2�IpĥkFU�������FC2��wȟ��"�.�o��� E
^�'��|D����zl�9��R�8UW�meu�\_�λ^��U���e	�� �D4i#��ݡw9sF:�x�yD��JB �{�B�K�`'o���p �il���� �n�ۏ��o��7�h���h�
`�>13�{�K������,��3b���`�M��'��L��WT��z�_kֽ��}�1�.|�Q�2A;[�b�MRb��b4q������)����l��8k�;o�!�����>5<���&�ܪx$���Un�nQ��EZe�w$ّ���G�{wI5��	AÔ������J��w^u��R9��R��G�q�`����筋��}])/p���q]c�YV���s�w,��b���N�h�҇"֞�7�&�A O��r3K��+��6(���9C}�#%7s�a����Z�E�p����}Vo���q�"��7֭q�d�}p��;����tH��m ŀ.,s���-{���>,ׇP~l�� �{;YwfJ�I�siKӆ�<"չUe��5�"Ŷv�865-�_�-:��ad��� :E�Ƭ�+��X�[g��L����$�<C�TfW�6�6���6Tf��]��O�H�I �h�q�Z#�ɑ�4�>-۩�d�:��B30d�i JDc���/JS���T)����i���F35'�e��>��T��_���l�N���h��7]a���t%�1.2k�b����Y�jSU������[�@g6�{��ߕk��|�>)�w���(F��F� ���L��GiIoH�d���'��%x�^��W?o���E������m\`F�buyR=N����Ǚ�Z��D�\�߳�������词�ޞ�w
�|�x��9O>+\�QΤUW���E�v��4�̘�+ڶ�xL\
�m�e7Y���h�l����z ��%*�
U�E��:P�L����� ~�����E�b�!`A��� ��_n26�'���cjv�7lôq?9�}_��
�!�#��';!�6If��{��,� �U�e���J��v\��� �xH�)�[ �|e'=E���������h�8�w��W7ѕǪ늼��&�ۖ"���dP�q͙f�P���9ە݅�fV���*�4��9���4k �����7����"�x��hL���~l`fO�b14U��W/M�"����(���f�۶�@:4��	a�-�r�{�նP��Ք��a`8���>x�VPS[�X>h��͝dF�b��ht�< De
cr'�`��\�V��� ���Ms�2@|3m9�����_67��8��b�R�b0��� Z�r�p������_��*�w0�Y��Sfg�h] ������o�T�W�f���3�w�?�3���$M�Gvt����f�j��Ru��kS?�k ��x������&jI$�M�R����z��lp�{鸞���}��$���4孞G�<G͊��g+�$O�9ͼmH�x���
-pӿ�(`�0Wa@�YqH����R$�Kl�ƴ���Yr�����"��K5PoR�`�������j1n�Bfk���WS�!�S�K��Y�O+��'�Pv�wn?����r���ʟ.s�}K ����u텲�Z�%zm^jR��ݣ��[�r��lw��%�OZ��}����`�#��Pk�3�[���'�9��}/P*�����F����ƀ�=��v�b�Ǐ;�YV�;�����v�t��M�Ҭ.�~Cg�/z��7������ðI�������{�IW��#c�X�}����-���˾UPJr�&��&�^�j�p�:��t;�q�mڇ��_XҴ:C�)dni�g�ōi����.���H�6˞��AFk%]ڀ����}vҹ��Bʰ��a�����p�m�]V�3H��a\Sɗ�:�V��I�ƀ*���w����E��3��IXԄ�J*yX��D���� Z����W��j�H�i�/7���y&Oq���يĶ�t����n����8�a��}&2�����k�h�0��Bt6yM<�·J����6��y� ��?5���.�ұ"�۶�l�*�_�:kGҳ!�t4U?��y�m����1�r��K�S�"���$Q�3�0"A4��f�fi~��w��2�Y����.H�j�,����ə�{J8Ia\"!�:W;�����<��p��5��ı��� o�o��]�.b����������yU��$ϱ�~!���紁���?�)�w�GSn��ӯ������^J4 u
��Ǭa�g>��N/��k����wf���bK�+�?���,SI�	��>�t�`M�^�<���Rh%޾�4��w@<���M���3��O�����i� B〠�ǐ����(���ךK��;�������5��_$���X�������"�5��-�cÙ�����"�%�U�&�yݏ\S�E�
���M��Z@=��#q��6���폙;�[��0Pr�q[�M�Y��\�rܖ]ԴH$t
h�/�t;�/;��Ϙb���ި^�H�<��r�!w��^�y`p.�0my����,�|Am���ʅmu���{��;��������T�tR�:�f� ��SO��`�+&��n5
i������G{��\��v��v	�-�7�#ȶuHA%��L�bۊ����\���L�Oת���bp�6����+��b���q�N3@TC�B-��"��eaL��@�Y2����x��R^�'�&b����Z�t��ǀ7|9E�rf��9�&(S9�.��q{�ӹ��tՃt?N����t�X;�k�G쭳�#��qb�%oG��_H�>���wiŒ��;�eC8���'�Zj[��,1�W�'�LH�΂�W��؃�sF�;�����{Ԧ��60����V��xx�`�u&�s5�ס(�.����[���Dq�7�-�����@�D	�m��1�t8�m[:��Hv>�d� '=\�uG:��� E��i����5x����`����Z|s�s�k'�MEƜ�x<�<Ე��Ԯ&bB�QU��b)������d����nbW�b�\4[��L�-�39��'��f �x,2N�v���o�z�j`v�]�:F�բ� kyq���GT�'k�lܧ+ӆ���-����I�@���+[�w�~0R<��,��2�<�6]�W{'���x��y�4bڶI�f:%s�P6³�T�>eR���1����5B}a�{
�b�v��@<� S�W���r��>S���&����1��S��G6��Gd6�OC�dUd�|�,��Z��O��jc�;|-)��eC�����t�PS�WH��9 =�԰������V 7h�n���:�EIXdR����: ����̒���L��n]R�Tw��C1�5.\6>�`�3@�~oaZR�􅠍��R�B邒�4<S6�N�Vڨ�1��q�P�;�>��k�j��|�1+/gu#KyY�����Bt3��̄O���W#q��e*�IXȌ���Z�}��`��>0W��AΩ���4[�8V�\E�P?�YK�i8���:N0�Tǖ}��Z�@k0+��.a,ď.vv�P�BF���T=P{�������P)U��J��&m+rI��'�H���a�Ō���!�3�y��/R2��̣��`M���W����b/��j��F b%���#[�n����F��o���Ê�T�J��1̼5�c��0i�_�����~�P����(�V?Uױc~3�wk��]n#c!��HG!6ѳ�@+�@D�s��ஜ���V��F���8"n����q�J2p��V��V����۬�4Qe��8���pN��8��vep̕�����I[���Ҹ�$��ED�S��q���巈#F)�f�ϔб�@�ބ�	�KZ����̴��u�*5��%]�o7Cl�9���2j�2�ReK�k{�ǣ��<f ���L(kxf���eM��Ƕ����-%bX��wO;� 1َѹ|��/�0zd������Zs��kN�9m�k*	�-+�_���S�ԥ��׉m ���^;���_�8���D��أ*�I��97��n��6�>4�_���
P�����6%.b&D�}�K8��ԵQR�%�#
������}9�j���oV(�O0di�%[L����`D���B�3z��[��-��k��eg�J6ɑ^1�!
�Wm5G>�u"�6s��+��;���6*��~G��v��HC�t���A�Á���C�mG�b��{�%���QT���ڳ��|�h����:S+C!$��܌����%H�R��ZۙjvE�a ��g�O���c4s8G��C�J^$Ɲ�M��鐂���ְ�av�Q��Ŏ3�ѵ��6��	�g�~�es*��i�	S���Nع��#�D-����@h��C�!�z��0�Tƌ���d��M@�em�?�h):��v�� �J��="T�N��epnuW*N���<�p�E3�:y�7��y�=��϶1J�8p �1 �����쯐~I5z7o�4kFn��K��چ���ߥ:t_D����f��K��6<��X�6rإ��!<�xx�����&�`��`MC̷zU��q1��Z��!n���	��b6����0��о�E�L�*�,V��po�x=�m���/��-K�!�O6�0�h�����f�$'����zgy90v5���2rr��qX�T�`g��û��6����Fh^l=��&���������K���tw�b�j4ӥ<�b�ccБ6F�&J9�jþ�\�J����h宍߄W�{�Ag�����0�d�٦S�L�!:��q�)`��W\GWk�'Bf���?��@&d21I��D���HI8!���`�N�Bj)�	�����/ AMs�}&�N;ŰR��NuR˩�5b���_��`�=X����]~����'�sC)�e�Հ3���1i�]�Y3ܿw��ӝq����+��i#0����k�f>E��w��d�R��2��R��w�IL��\������#0)8�?��#¶��\*}|��$���B�'QM����q�O�/&T��h�at�D�|��#9�ᇸ�[����z8�Xr���J���M�? L���=�u����Hx��V:,F���V+�WMG��pY�p�uT�� �۷��#���c(A�����R��o�d�+H�&�CF�Ym���1F�Qi�D�,j�|7��WH��^b��~4���w%��9Sf:�6C2���Qj��6~X ���`�|��5?�B�M�����Q�]�Ҧ0�M�ʴ �/!��p�X`�e+��w�BZ�c�YU�6�#�J���NR�H��6��>�Q�XӋ~oiu�D2����mV㈗�]��~��鱜q���އ�d�\�p Z(^�O��t]�p����v�G_���+I��]��#���8w�wu����Z�Fj������HP,����}�>��5楹���S���T	A��V�D*�Oh�o��\|�e��P|܎W�=���z�z�(̂��"UeCE~�=�4S&x��0�<զT���q|L@o��j�u�È<��)�6� �0�~����LMv��3�.���,�U�HQ�B�&�(Xl�K��~�� �H�LA�6������ʩ�:T�>>�x���/�oA6(냗6��WP�;�4��mWW��ac�4z2����B�f�MhI�) Yv~���P/�@_�R�}j�7#��<��.:��}��%���sq��z�6��W+Ҡ�~� ����x�?I ;�����Z �� ��MeF1���翈y��U3�2�܁^u�nXw�4d~��
>1a>PZ��)N���6#r���	5�2���M�����ʲ��'�^1d�r�z��]�~fv�b��3�lHJ[T�W'��+�e:=�y�N�f@���%�l��b��,l��ag�p��^l-�C;�0��c���Ð^n܍NFs-ٙƕ�A6�7
�eL�J�iE*?�&�~�� �SJ~I���T} ՛�Y?��	\���T>�t���xl)�e6hA��7E�۝��n�vѰ�ug]�HQ�,��5�)���Xp��ϙ`?�B͚	�Gѣ� ������9Jq�|�J�
qIfq�f׭29տ@ҌѪ秨���3���A��9$��vG�N1��DY{i\(~�"җ`�O����O5 Ϊ�E^�ʽ��bh�Я(<r�0���h:ݲ�z<�{���Bv��ǳ��)����MC�0���CY�����Xv�<���j��(-�#=;�6�8�񡗀_ZH�|�b�H��M[�Z�L]AP]\�n*���c��F��[�ݿ<��cC�Q�\䨋��C��Ϛ%�Ha�Ѐ[@+�e o7}�쵉᠞�F 9�	��"�J�U��2X���~d��ء��m�)�u��v� �S�A�g�"y��_ٝ��1��<�3��Z$U��*i�N�`a\nP6�]/{d����&?7�X*��˛g��o��׆p����Gd+�D?\gQ�[@ԝ�!�=T�$>¼�DCu_N)�����)�{��K�DBnl0|f����s�Z��	�4�	k�f�a���|t:���n{s$ba��>I2�FT)Y|�g��fx���^r|s�U(��}�O���"ݐo�`g��G~7���)�h[x.Q�u��iH��M��|�{�!�=���s7��F^UO}��0�ܱ�:�)�C��һ�@�鵞S�!��P�r�d��=���;]�K
{WT1]�O�2|�:�)3���n�q�'�=�U�Gn� q �����8�2/�I1�Fi�x����|vÙ�/�5������r���ǎS�!�w�᧭�x,���-�?0�0j��e��+<T�g3/'��]��!��u�9��P���G�=�х������������+R�:;������,1"�P���k��Og)n	�q7Io�M��	�ρ�Z3?�+�%�$�V+�,���8�7]ބd��ɹ�
���F넰��N�AN�UI�&[����X0��������X*�k�el�G��WV8��<Sf��1ҪR�lQ�u˻\O��Ћ�)X���] ��El���8�j�W �T�D�����_�j�w��4?��AY~��)X���z	�{��F��I��'ͼ�Ro%���D*��t���x��d6h�q�����ٞlR���׎+��W6�����G�yT~����������^K�����i�����@�����@�U����?3����jڈ�ǲx&���L��:|��5��{9l���_[�(�5�2��7�\Ő`P,��v�v�(kpɞU�m���S��E3��8���U("���W�����$1\�R�t�K� րz-�X����VF�+�>��+��\�a������v]�6}:C�v_�	v`5����3`��>w�6�kyC��l�k���_]C7�5�B���צ�#��ي*;�'��9�����ҍ�y߭۾���ԳޜGA�,�4�&!�b�r�,� C!�	] ]�Zd]v~��N�d]�R�(�i{�w�?�p%�v�F|���g��	^6��=��n0�,�����~N3��S�� �h�4!�����`�q#R���O�q��n��ϓ�d�XAP����9����WF��Bf�"u���M�}1���y��_��*�Jg�m�w�P�lD���_U«غJBPO%<p��Y+o>�a��	�˸�O8�kФ4j�ѡd���j,f�_��ҹNin��)􉂗���A�N�v�Kb��ӄgY���^�Ufe0��Y���*}���#MqKa�ߧ~�	ԅ��
3�|9�Ƅ��Q��T�r�d�.��ɧ<���h|ީ�z�{M*�n��2�V�{(��������AK�\,̋[yU% N���<-�͐��V; ���o��c�+��|�[��<)"�Ɂ��2�tJA8��6�%F3
e�y$O45�*�SJW\�%ڨ����c��I4�=Y�� �Vg��A�俦^��lLa����S>���h~k��>W��7�3�fא�L����������ӏ�h9��[�nǒ?/��G��P����]>dUo��\��몳e"3r�W`�O�S�Ix���Vj״�V�'����I_���D7,7���麙N�r-�H|91�0	zF�=�ŲlY��/`S/�HS�"eN�-)�`<2��!ֽ��=����vF��������V��t� a�W��<6G���m��Ѧo=M�ў1v�K u�Taj�{���i������CtU�J{��VE�X�ߐ�6w�a{�9�E��G�؋T��C}:���cO�hA��\�QO���k&��:aYfW5�C�V��̹��J�V({��La�����-X
w|f~��m*Ɏ�D��4��_z���OpE���^5�(p_��UW;sB�F���I�����y����R�i ����/�h/9������X�\S��V�<8d���%���Lt�G {fq��O$G'��r�@kZ�@5(��Mt�,�݌X�N��8�ޫL�ܶ����Aa���^{�a�3G�P%�]`ݼB0 �:��K��;�o���̺���u>�>��Sr���bN3�6��J���:��J��[�$щ�Sv�6����F���2�4@-í��H����_� Y��w6	w �z>Ҍ 0R��눟��:,t�	אN�T��M&x���S���K!A�9$V-k�^[�ɼr�J%ߢ��~��o?]��@�k5�F!Լ��p�w�*q���x�s�{�N�qOז�T��'%?$��>[�#Ҭ�{[�������G���	&f1���k�"���2�q���Wx\�b�Β��aw��Y�+��O���ue�����d!���J6����Xyo���u��EC�k5bjiT�t��� ns~ۉ��-�e��^G�N��-�ڴ�
h�n��߸^�Ǧĩ;��6a
���o?�7EX}0�_(��%�����,*�1�D�RlsH?6���!P{�n�����hD�q����V�粮����ݯ�)2��&�[�Q'f>ۓ�#�b����^8������`�D�T~%���o9�XW$�q�˪�Iu�{F�C~O	g��~׺T<�@{�r��a���)
Ad���{����4V\�4̄D��iy�'Cfo`8=S��!�˒��ߤO�H������$�a>�ߜ9��Һ��8Q�-Ǭ�}�
�,d\= a�*�{����;am���P��zXd���D�+�$�j��N�?iA�q�/	{�*�1ef����G�#&AA���q���6�4qO�G�L��v�4�E�ˮ0K�B������i�L0ry$��zQ2�Д�f�wu&ˢB0uT�b/G�WU��ɭ���� ���Q!����uqIԬ��쏅�'og���^��s�l�Y;9��r��3�U�\��H��:��@����m��4#��[�9Dv�$�uY0��O��^?M�IJO*kU�2��{���:��`\Υ@WqNv��7�-3K�}l�Y�<4�x'�^���y�k�F�/T��lޅ�^:���hmT�����O�$g�QS�mSkA�tl��
:,{�EnC\4J�yL��q{�&c�h�s��Wa��Y#�aE^�R����-15�hܽ��Y�9�����(g�:�7�ج�3t�W:p�TK<��P�b��k0��'y��	~Xs��*[��ڷ��_1*��n���(0�ԛ�Q��%����{4��+��Jࡢ�����B�@e�4U�`]v��"��ߓ����%R%Mza��ǵ&�`*�13H�qwذ@<׬�\#`OaJ�j�Ŵ����}�*a���f�;8�t���Q&�WR��K���^��J8]��8�4FY3���:10�/�(Ҭ�oQ����U�r;�L��Zg��u/ź�c�ȼm$X0O�~U �iz�&U�0.�7+��_�<����=nS}Ǝ�����vo-��6`�yj�*�hB����ہ�\ˁ��UM��ml�ܥ���7�����?��ی��̎R��݅�ܞT��G���Z|=�	>��E��Kպ.�У�t��֕|�zN�H8)����ٮ��8�����)g�&���H�[8(4��m�:�j��+�Ab_��vҢs�s�J��B�!�Nsi�x������6�G8����oP�}h��S���E��<>�����_����p|ǀ9�\�P���n�DJ����!(;ׅ����� &?F�K	�+��VlC��DUv>	���0 �96ҽڴ��\��	��(̠\�I|�=$�O��Z$�o�ѹ�Y`�6��������b�����_�Յ�C�?b!~Q�!*:��_̚;��T��S�c��׎�]`@�em~JA��}_0�e�t@��\;��ݚ�WX3|��0������N"��^/䅴���!��s�wą��$R���r�m�i���q�ޙ$�sX��5��֙V��.Ȇ��l5�o���?��z��ʞ�-1�2���`���%2w4~�Q&5W"偠gsP�*9�eD��bչ�����B�}x��F�wQu�{<)���F����4�^Y�5��7q�na!4[(�yJ5�=HF!���7�ʞ|s�`��PRӭc��
ya����e�To�-��B��)���P�֓9���m�B�_ �j ���]��{���4��]�	zc�FH�� D�Y�x��ޛy��x���^Ls-�)�n�>�<��ՠ�&��paY���p$L[|/�yp;B�.�z0#v�#Sp#kn�X8��������u��9z�Y�4}uSu����B�Z^J�E`K����<�#�tF��o7��<����i�늧�_� �x�Oi%Q0�
�s�12��u1{�L|���q_��y
�>�OD�gn]�X���C<Hp��2�a�'s\BZ"�.�9�������tt�� �Q���"�=Cm�������న�C �Zk{�.fqvZ��K~�e5R���Lo�؜���1Ȏ?�X��V�4�:uW�4�Ș m��h߯�!���g�N��ɚ�K|�����k=�R�@Q��M�Pv��d]cpC��n΃;e�`A�=R�uDpk�Sr���0�X��NM�,�@��ho�
�����Q�L����=8_���@.�o�|U���k&\��(AD�\�2��(�b�$�N����7��;�0T��മ�Χ�E�����O"5)n��t�쏽kW�����[�#���Yq�jzq�_�T��LMi'(�T�ta��-:�n���qe?�c�x���ZDv?����2����Ʌmj����{'a�[j�
��v�]5��8��# �Ī�kzҫ�4�!d�ھ���mc�`<�zn3OU�آ��bg��hA?�?�&X�|7?�uBk�zu����J4P�(���)Z;�U�/�Ȉq�!���4��m��#��M�B2�]�AA��T�?�WmH.bt�3��T?@O�K����ZW�F�=Cy�mdW�V\����4�C�fw[EvM���(�1�Fvk@�z���a��$��//H�e2&{D�MMQy��o��]~u1i�}�;"Z�J+x,��ɞ��#>y4F#�T�bf_=5�|6�[E!᫤=�5ƋX ���N�;��v_�[�q�H�p>:���j�5��O�����E�u|��^�їxPU�y��}ז�V45�s�1
Lvar�������^D!�����+-�L�z:���ﲃ.t���a��k�7zZ6�� s��B����d:��]�Nbŋ��E�7��f�9��A���uL*$;Atbo}K]V�6�T­�y�
z*����jV��M�|˄��W�~V�2��#*7i8�eЏ'9ymG�gP��S�2�^���J���S�5������j{�jL�����\�0�$d<�Ý�������XYx��O ��o�wۥ:�ZŎ�xTP�f�;O���N��N�*��<��.��~QP�����1r%R��.�AxG|���8x8Ǩx�Jʦ~�f�o�ư��pCn ����tҰt9Y*��hW�����MO�pk>���X�h��	h���S^��A��]�e��6�@G��HS*�,�_�P�3�@�4&v�ɖ*	f�L���pY�&S����j����E�;(��ʾ ��ϕ��t�ύ�x��;��3l���Q���@`W�\�%�CI� _߬��� �Y�M�U���f�\-&_�g>�x�H�l�:�0�w���z�D�pb����E���m⸣��_��5j����[L��|E�{�-a\E�L *��	�zG�?@! �"����XJX�~�U�L�W�)��#$�5Ҕ���/��"��uiW�2�^C�����
��u�TI���#~Tx��ƃC�Ǯ=��(-7�ʹ�E����\:i?;k�~�����S?Fc��rD��I��4�Y�+�# ��C/L��Y�A� �����ˠҊ�%?[�0��~�hIC�s�/����:҅�T��;���f�B�,��E=$%4�Z���-���C���12Xy�6���+�m���ql�����P��f�B\KQEě�}O��W:5��,�1ǹ��?š�֌���kS\W���?G�dO ��-�e�wl��J-��qP?K"r�:|���i���$�eӓ�Q�,�GPgRVÏ�A�m}��_�k�'��밴�u�������jr�9��_�.@ҭ彇���̙V��rz>]�Uٙ��=?]�v0U���u&�^S�4��������0�
�u
r�fo�$K��Z��ũخ�D�*	�8�Jf�"(�a�����#�C��h�M���N���>�a	���j3�m�#.������*Q�0x����v��@\Y�U����I�k��AY�O1����V,��1>Z$�4
�!��A��m��I"��3!�)Ib������+�J����L,��F�V���8�߁1��'�(����rn+Q*���13�H�k
�uk�B����k�w�;�8_�DΗ1q�.�sM\��_"k�cn��:�7���PhC#�o�}���+k����v�Wd�}���K�(�>b�&���x��W���^�$�~lɏ2]/�I��o�@P���&>��<@u��|KOL�P �+�.c?a:q��)���C,}�Ķ<� s��q�J��/�Z	��:�����i۠�?�#�
"��<�)��9:�����u[���@�ܓE��5+-�M����o��נ� Q��zDý��^�R]����u�̨�k�ye]�앆�����5���'.����D/v�C	>֋��D��דgT�z8�T��X/�ך�ȍq��J )��QK�Wԃ@��pP�ºd�=�o�>���;+�
��0JX'�В��iE���z|��{ ��̛4���b�;�H�&2��Wڛnp���TgY=Z�d��1�bO�Ձw�2���X�-�9�'@�3�������u9,ﯶ�j�����.,�����b@�h�l=&����*N���.�*8ཏ�?gT�]%�Sm�ǑU*f�q7�8�`�����I��|�����䁡
����pI4��U�5�9k4,�\�:�k�|?�����-��	|��j��ڱ�r�-��NXL(o5�o�r��2p]���L��Ť��g\�I3��Ff��ͻ�	L��7�I�����y%z�ɕP���˺R7,A�p�o0��F��������ѯ�ə�YB
��Q��Ը�vjl�Z�S��qa�x6��E�Hg�P	T�끱�D��T,iS�BWR��T!*^������<�z��ooS����P�8ǟG�挩֫���w-���ۧͪA�O~#J�ca�̙A`������� Z�J 0Z��?����
���Ǌ�E�'�|��GP�4�v����6�F�~�7��`���㵂!�a�T&g6��qı�P�������}01�	�iV��Yd��r���_��7Až����@6WZH�"e��n=�
K��FS�e�n�H�QV;f"���W�<� =�~%a?��4�6�&B@?2�nU^��4�:��]�����{�<.&�@z4����AX\�lIX�
d�2�B�J�~�� 8bF�c�Xud?>lU!hRϤ�cpi�j������Մ��g�~�b�� �Y9AJy*�2H���K/a����_Q>��1nP����E�S����*Ӌ��G=8��%�)�Gp������[f�~���)�_�M/�g�N��T�ŧ\��B^���2���2���z�`�C�8O�s�@�ôK}٠�q`S]�\񁬺��<`��_&�Y������"�����=��Y��֓��cL�hG���?w��oa��S'X�^�am�A=�8�E-o)A���� �/+����=����6$p�����`�A���
��=94a��a�����1_G	)s�F�+�O�u�3�0=�LD�ߞtҌ�9My;��=�bv��Էt�XKk�&��W�~�CkeU�jRg�$(��XrĈ�"��]���TiB��9ǋ�}aMi+�"��PX�RZ
��� �Z$d9���9�m[�-,/�U�ڷ�g�l������oh�:thz�8����!X&��K.��R8/Ʌ�?z�T[$z�ȳ�5s��g�7ێ�E3�Ilȟ�4V#�i��Ю��T��{-���;g�ا�A|6M!�{��([�������
����9�+j�Z_�!t2�6<�*J��HM��=H�3���]�T��KDrpN([�s<�)q���J�5ƜjW_�qJ*��?2������-aDS>l7!^�b�H���;�I�	�'�zl�YHnn$����]��e��wن=��uAX��;s���ޔee����0 �q�s@7Eo�DA�_���{�B���=���&6��5��o�]�J^������m4u����X��"?T!��>��ވ���~��D��
/Þ�甒�-Z�t��ŵ� �`X�[��n��Y @$�!z���.�eӤ��
��63AV[ TnFސ�~�=yo�,�ȟ�?����,VG+r�鎫FkG=�>`?�������^�Xˡӏ/�w��<W�����O!	�a���[���/�xW��۰A�l�{���{	�?��^ѷF����!�Q
���+!I*2Ql���P���Λ�N�!�8�*��o�]�{���wh�d ηu�C�4<>�ц[�u|<����U�ly�Z3[�׭8�*}N���@ZדT]�6aŜk�lm5�4��n�bf��� =#�mC��m�ek ?:
���VЀ���?�8h�t6�Y�$���ӻ' ��S���0�&�xk���-:_��S��� ����q��e��@�*�3��#(k^��
{��x:�4�����D0]*������"sw��Dm0�H�x�� ����B�;"�+6�b��@�>A���^+�����x>O�g�@U)��oT�'���IO��
� �S�햻h~��)���q
�V���0nAGX�����|*�ķF��X�'Y�sgE�ʆ�ѡ��<���4Pߞr�@��M�#7z���vi>�����d]�|
���hc V�HM��O攳ml�+�D`��|�[���q���e?� �
,,���r��k��<�^)G:�-�U�O�UN����Ep3'��%Ǖ��0<�m�d�&�)���	Sk�q��6�\{�W��=�&.�ۡ�(4����7w*>��q*_¯8�{3��b�
������,|��k����&L������������aX��|O��@ o�U{��n_&3���ߖ��|#��B`���%��!�T�v�l)~'�:��x�1��)��jfB��~��4)�k���;
�L�D�Z��P��������J��r�a�-%pR
`�s����"�Ku����KS���4��g]����/+�O���c�
4Ϩ.�}���VX�"������p
o�鼼���`*�+��I;�7�z�~�"r���C6P>�j�'6֛�.'۩��*���?�k=97�v뺵!��Μ�e3!`�vw&��(����f='c���{�<P��CL:�.�v~��#y 05 �W��T�������s��xZ�)�c]���8���{���|]^aeۥMM��T�v�gp�� �3$qYK�ߝ� Y5o"�SR���oY&><ZNW���|�}�3��w�Ug;��=.��E(Vz�sk��=�T�MQud�q'����1�F�>�i.�c���R嗱8J�^-k ܙh�6be>�M}j	I H�-��8���4�6�91_0���*�����v����.r�!����	;Z�.G�7+D�\�,,sy0���.		䌸���7J�ɦ�	^P�b,�b���U��
��Ů%�=ĩ-*�稃
�8낌��OAu�"����{ݶ��+d"�\�nUIy�_M�rEl�w�ʿ;�@��W٥	Y���[P���?�� W�Z��$���*��i���M�Y\"B8��QQ�9b34g��sw�HL�ߡ�9[gI���IMZ4l�j��$�%s	.���~y1���Xі��v�:�t���𕆆Y�˹�b 3a"G�Dr����)5�bZxA�e��+�N�i�b���)βU7Kh���Rz?��W���Q��˄��S���24�!��{ �qIxIP����N��y,�T�c8ȳ��"��ׂ*�X����Ŧv��+Tp᏶gF}93���".�"��-c�^:���-���ru_}��z��d��9@.D8u!��#ҋ\����5��0��,HD��+4\�#�U���i#x��^��4&�޲���1W\�>}j��gX�w����8��Շ��9NN��s+�儘s�@|���*�>�<�_O2�jɔT���~{,�B�X��]�5z=�=�����'���h]~���3�x5}�(�N4�MXi�	�0��_�����ԉdpzO0���XԠ���M�E8�+�9�LP���_��%��+q�Z�{�����Z{��΃��"
c���џN#��r�wJ�Qp�y|��xeD�']g��Hj�n��h��W|L<�n�s�֏2\��>MI�"WR������`�Ϫ��4����Y�Y㎈U/s�<�z�uW`&B�?<8�]t�/��k�m�&b��˺&Aki퐑��@) B���A�����}���o��ޟ�98V�$1�R��`!�I֕x@���=)q�����M��%����W�K$��!�����0P|��[ xl7a�CsF��?8��ze��F7\<�_ aAm�ˌ�,Sx���W�bM��c�� D���S| ����)���|IEʀ�Zcz-�L�$��@	o�<�|e_�1||�����C�G
v��I�"�4s��À�0.�bU[��
��*4��j����VF�}���~ӑ=��~�FܓS�I�/�&�x����WōY}�'_�#�aՉK���e�+�;?�9f�b�-2Y^B���x��:L��J�W>��H��&>�)�K��ܯ�g��W�J,�����g�~�'��Ǜ���Q���f[����-i)�W��N$Wrx��r�ЎDդ=6�@��I��:�J+�In/{c��V�H6���Z�S_1@@�s>�����܀B���2eȽ��5��u6=�n�Z���V�e6�_޸����&~M9�$�Q�n�6�pd%���-f1�wF'���Y^�!�=�>jk�L���R廷��,��l� �aϿ��VҐ��b�%��~�rav����o�DHOk��mZ4���I�1�����/ƫ�s}�/�4�o�.4���9`qd��랒�6|�}S��4AD���1�p�1#��fAzY�^\1OI}91��]��w��A)xi:����	肃sy_��A�a7z��X"�T���4rA��Ѯ�+�"1y'\^������Lt��0d������~���j�B���(�J!��+nEu:�5��D�}�a���t7���:�ԬMu�$k��9�N�LN�;��~�?t���$d'f��^��h��= ��(�9�����+��A#�~}S�q��=�J�<@h( (:�Ul�,3B��&�xY�E*$>�J�P�ߣ�^ϖ�-j�� y��.��L+�Q#RpEH���oy�>w�σ����{)��g=��w۪�)��AX~��2H��D^5i�7�������V���7�	T\F�BI'�qB ������	u��W�Ԉ��룺s�7l��6��A��>%�7�m���@�?��.���t�`Q �T*���jܫ��%�~����}�rw��w�μ5����ˌ���wQ�v�}1��')<�MD9���n�?��{?I��&�5"#��6Ga�A�j��P���pw۞3�Tg0�t��\���=�8}G�ܥQk��=g�E0,� o�[�U��'��0E��39�3��x����2K��|0�!���5w���#��y1�|�QX'�໏hd���������i�ʖƔ����?4/���=k'TXdg��u4�k��ׄA7��BB���F�F}����I�/(Tm@I���	^���S稲��t�T��
�r�������Fe���uk�Ө��$w�CDl��:ɿ�@�D�c=�����'U�Sӹ���/�!�}���	QW���&#1�����nA�I�,*XҐ��؆�ҡP�M8ԣ�ZL'P/��OL� �Fjy�Wq�u���YӣR�ˢ̻̬V	���|��ApR��m��}�7��f�e	 ��S��M:���
թ��]�"�3��@���f�a*^0����^X�v�;���{X!���@i��N�9�`�@�e<\��w����s��@�
w��n�9t++�%p�����\[^Ƥ��-�"T��v��-��eՉ�8k.J#�oޫo��;�Q'���޻ޅ�jL,���D*+ݱ���j� ��s�H��iZ��B���<�IN
~�d���e��D���7�e���T���65[ޥ�Ռ1�ؖ��e(IC�T�A��2��(��v>f��
P3�.BDE���9�ôv����.��Rݒ��_����4-�ʠ�8���|k�|i�w�'
V�����g��
�[v�OJd�O��<������lD�����y��ޕ�`�	�E��E)% �������c:thpG���"�Z�u|��9�K�t� �,���t�� 0ç�q�L�h���P��"[ʙ��D�DGO���إY����9!o�%�!|�T[I�?9Iы��2�?��@���u�"��eڌ��x����>��7�R��<U$I��w��U��(����	���#O!����V*�t������N���X�<�q�E���G�����:<l°&OD��������W�.���[�V,�x���`g��W2��R��!\s�B�{"���+WT��^R�c���o�j|o����3s��9����޸I�II������N|���nfM.R]"e�Q�Xt_eJ��|i֦���S��B�e�C&ԫJ�3��O�j6�lS��/w}U��
�p**hxh��IC[O��G\+�DC9[�K��5��i�~Eֻ|4��b��m�*�@�.�9u�%e�v%����*?�IL�
����g>lik!�T!�e����.�[+���S�|q<�t��f�fpnR`S/WL���%���'���o&S\`�y_V���<Vg����`�'����W���g�N��}�Ь�#�gʣ�G�vIF_�>�2�ܔV�� <5�em�x,*�RS7:�ihO�ɫ�$�z"�Ga'Җ�1�����ɍ�h��v�,��Av�'rQ�tz� (���~����[�q�W��k>����<�[=Zks�|���e�O^%zr�cs��6ְ�5:��\�[꼽@���N�%�k�5��f��-��`��X����N�e�[�.��E�_�����QF�̥�V6�i)�:����Y���;K˺�ٚ4g"A�ѿBXLu}�)W׃ P��ID�X�_�]��T,�9�[%K[T�ʼ=������"C^�.�|�ξu�^�jc�O����b7;�U���G,v�ձ�&�]�����#.������!Z��1~d�I�{I���{�{�֠	lB��:$��̄F�B��~QH��r��Ȝo�D�ş�-etO��Z��fjտ)��!V����C���u�ӌҁ��,�Z�?��Ϫ2(�(�TH*�W�_3���^N"�XO����;�̵�j��a}�d~Z��4$`�����7�SG+���$;;���k�R�d����i��G~�Q�;��~��܈ó\o�g�u_w��^���t�i�3R �P~�ģ<�k�/]�+c^�}����.��	=L_�����@`�YAQ1i2�[� c���'O�wx�C���-[�͌s�Cer�u�:�� ���^����gIrY�phz�\�Y��KK��lxw\�0�,PMڹm��+�lY��W����uW_Sb[��y�ǲ$	�����׹RP�5����+�J/�(�M��~���H�uʕȶ�S1:��z3s�p���îb]z�2�Kl3�~�v���/i�M4���R�Ŝ���84�@z]�I�,�N~yJv�����'�v`�+G�4���VR�x�㥊G���G���q�G7,(h��@����v����5������y�@�.>i�(���E���)��D/���r��{���Kf�|��mۀi�ż�u��K�����v���gW�(x�����fJ59�ßE:LKs����Fw�D0�QX��Yb1�/��v=�2���Q��:0�E��Ky�$�ӷ�Zo�زdp] �|����ر �����^�=K�%!�����:�}*�� �Cu�Jm�����)>��\c� �頓Ț6�k����%���b�O"���z��Y��X��`N�F�âP	��CY�O�E�k뻀�h_��&�9$zh�� �h@���}7j,<##�_��D��c� ]�vi��s|g�b�����;׬���W���'Z���>M��ߒ��ē�yf�C�6d^������!?����N؄��7N�~E�=�<no�D��`'���Qk�am���(T-����c�_�����p�|B�;�gWf���x�G)N0!�yA��ƈ,u@�VD�jL$� �aY�4�����>���8�a��TWme�=�� %S���@X�E6#��A��˯@��U�A
�Њt���4�@�{�k-K�,l��1`K���&R�CH�SX�w��͠���H�3���r.b�UjL�7��=����*3��$��_FM�0��e7�F�^1|u^*��r ���r�ɵ���k�}�X��\�pn�Cu�4L�����$}'�R$��>}��9I�͛���p1�l�:���D�������2�M& 8,S֪�������N��31y��胰�����6�{�z��*�Mo��>5�Y��G�������1P������ T�k���,_+���4r"���3�K�Fʵyv	Ȕ��P0�
�W
|ӈ۪ۥXW�w���f6a��U�
��F�4	h��ZJ0�c�r���2�,�4��k@���g7�&�&(��˫�{q+��PN>�o.��o�)T�	�z��8*����w����V�N����A7��VC�Qa��I�4!�!OL7�N�G=�]���3@'m�����׺���Q�>�rI q�p�`�|���`,ܰ��������_ɷ�' b�?����l�����}"���H�S�|{i�}���8����|\2O�����T�weю�D�L�U~js���U���)%�E،"&�DI��_��HA�7q.�:F�wP���}��H�4u1��uD��H1/uL*<��.5�&����W�R�x��4'.^��w�R�	��,���e�4�	ӻ-ψ���2]��<�$|
��Z���確�WW�;���ʇk��Ak�r��4�N�͋TTXS�5g�y�Q���a-��@��|�u�!�����r�t"�f��$�i���4DE��L�6;}�{P��'Б���%�R/0K&���WQ�R�x��ȣ����7���j�!E�{D�(����_+��o�v��A ��-�3�e���TE�.>�#M�t�Z�RXI�Wx\ԾM�Gx{yZ���Dh��D��It��*�U�u�7�ZA�_��?����^�C�t����!*.c�]�n*�'@�$���g|���g�-T7��Hz����hOֻȨֶ�ix)�A��-ET
��K܀��gO�Aa�{��I^��R��=��G�������E��I�j�'�	Q�G�lt���A;��3X��|jΊ�'��$��[�q��܀��?Zӈ�K�4��ZҒ�jH0U��{|��z+J�����ƾ+���(*��ҏ?E6��5Jƞ�$J��G�"�e�=F/�V�k���]���ڕ�Ӳ��I �����H�a�~�/�1@�V{9vCDIġ�CX��6Z	�57�	+L\G`�'(�e��֭]��A0�����M���f�o|QJ#�'4T�=(�p���h��l�0e1Nh�ƫ�L�" Rڙ�FA7��ܯ�:�}������%�ν���|��J�eH�L���d��[��c9m�>�
�
�ԏJp��f�ٺ�K4`�������9�V�>���B�R���f��3�
�q*Y`>��:[�������1�g}yw�l��>�g&�P�\�!7Y�a=|˓[��>l���u0�m�ghs� a��ä��v��Tܕ��70;e��Ϸ���DN4��䘉�����v@/�y��K��p��(.�"��(>�_�G�wp����ƛ�ta�F��Q)y@
�zRմէ~���:ˎQ�"��摢D)D�b��;�G���-,K�aU�@��Z�'\���%ᛤ�g�F5�'\oO|��:Y~M�U8�=�$��!Oc��O��Jb�?T��Gg��	#���کp��(1 R�̀�aXFU��w(�w��6��He_*!��a$p{3�^~~�����B���ӝ�ڌ"�Om$��ه�d�:�nu��v^7�<�[h����"SU�Daڮ�о��� 'L�e�y���đױk��+�y����2C�BG�Ix�*�7�oޖ�]����!z
��Mn23\����i�[�B�E�ς>�?�ql�)z���=�pSꗏ�������T5�Dֽ�
%@;��4oX%S-eȳ�(@#�y�LH~�c���U2?�_���dAwfA� �C*��+:��m�2j��mx���)�[����� ε�_r�p�/�������r�~�;�sޏ��z�1L�{�Ob#�{l;{ˠꜭ�F`��1�ն�W�u�7K^�ڂ	��ú\Q�}iY��v�A/�`��$f�g�臽��{G���T�&�_����<QI�%GC�z|��㔮�}_~i�9_j*��A�>3E���J���ӣo1�{M#���QC78'���a��P�@!!�0��M\,75�J���X�/|��Ѷ���?�,]�٨�d uY�a7Y�gG�"�r�����h���=��>a�ݨƉN�7����mV]���Fy:X��y������e*HYO���v��68ԃz�KԖ�[�Hy���Dw��m�2���WVY�c�|�P���+7�; Y���B�1m��Zkm�;����Qt^���F�����?��1j�|����=(X�MG������]S��B�%gxȿ�0�f2c����>���������b��$j��Cn�Ǻ-��A�HPO�����������ę2P��.������CR�m�mম;���c��Xx��67+���;(��g=g��QR	��r��K>+ӗɳ6�O��;l��`y�|!���gf
A���-�Z�p7�o��S�`�&�G �&�8�V���6)����v��m�!(4D��r�sҵy����mT�֜ ��~�H�MU�	�0�g#�?�WˋoS4��1
/کJW���?:�ɱX�4��r��xG��W�
���0P9���Q��k�p�A��Q���63��\	�ݟ\zDj*�T�����ZL�u�M��?�U�)6�}�bj@�1f�q��E�Z�Zp)Ҡ#h�����Tp'���ܡҒ��#��lI]��o�o��V��XV���{���Sz��.�4)o2?Iˑz&OQ��%�x��-���F��C���i�T�ԷL^�X�%��"��J�X�#{D�r�{cs�Hp��
;���h�ϣ��}� 5�p��STZ�oL�!;���o{�������F�Usgu�DU�)��[�`�n�6�fɻ�(�z���j3߀����j�%<d�e,T��V��� 9���*�C�E���12{�����pF�l�VN��Lٞ!�;��C�Ȥ%��t�S�,�j$�oU&���6��w�ѩӔ�y���C��j�*1�����LhS�|�Z���>Kѩ��~�-#Er�=�����p��P>h��zY4�O��SMms*��f,����W��[Ϸb��{[�iV�A	4O����I8�M�3@�'��,�)z��=��%���ۅ�n&��
�`YlN�m�������~�?���XȂ����2}�"��gD��f4pv�ɒav`������ϕ�h�#P���1�L�����o�2������ &�൓��N� _�:�
ǈ��п����Gj�6�+VE��.� Z�f1�̉_��'u��>uY������ȍ��AN٩�/F�>*���Hw�4�`��/�Z�ܵf!_�t�ڋ6�D�V@�c����s�A���1�QX�mHb�����o(N��Aa�r֪��3����D}��m^�Ɂ�?�t����p.V�
ƫ}.�z���'&$��&4ݬ�䲰
<��t�	����Mv����րܕ�1�W�O��u��.~�n�p\QG����VZ���n�4�ɓ�h����K��|ݞ`灬XG�{Y 6������j0M~����A�l�󤽛����ɹB�99>�����W�0V��&���oxy�ްyU�j!�Z~�:��hC�^�:��N��_m�[�^q���A��M򻠎�;ai:��%̱�+���I8�	M�2&��z�6c>?}�ʩ�'�ѳ�(��U�Ʋ{"3N���,���AJ�����*xU�?4�B�H��E�$^�|�4����� ��k_}�2����0j;Q]M;�����G]r~%�T��%U�7Lid\��G�v��&	(�%#N��))cՋ"�w�hf̟��SMM�yd؆�x�/��T�b��yP����
�k�lM�J�Sd�z�!�ׯxH�ݤ :]�M�=X���H&̘�;[�^RQ��hLe��B��_�;.��p�=��'�ud�o!2��Dה͌`��P�X��\�7��X��~�g�\Ʒ�I�
%�!f������n
"Q&�D�C� CH�M����c���*��4��}'����oZ��Hg9�����q�}��6�����n�X�a���"������/�eT9eCsPƘ�z�p&��sfE��KRI�m�����ր����I[G63�V��>��n%�b�A��'����f�d���.�1�\x#������a-F�C������Dǝm�ZkJ����:���;){?x���&2hD��4E7�_�C;+���ෂ��J%��n��_��'	�=���A�K�h=!Eg���M�^*��_�F�B�Xv� ϙ�@K���PS��N��՟ՔF��E�q3B�Ӱ��ߎ���$e����=>����e�{�=���p�!�0@?��a&s8���N:�7����U�c�m�?�^<3|p~�Q/mFKI��2�y<���d:,3����
(癙��+p�}޿��ϙqZC5���.������W��?��Y���-���M^A}��$j���θ�5����ڄ'����7��\3z��4��̿���s�/��(w��C`݂-rxz�S���H�Ņ0<{�]f{Wm}����&�h8�]B"2<���<j=����Y,�>�b0T��+;��"���{�bx�5����L{�]C���u[B�%b$S0��x{��"Z�NT��A�L��b��G}ޣ���V&��"�6"�`��L.�S�j��D6��L���EWoOQG�SIP.�'|�}��w/U"����h�7����ײ=��y%�:��5MY�G�q�+%@S�&6rՈ�:^w89s^)���XF��d�Uëi5�2Z����^?���^q�"�5%(/c�� 
��lK��ڻu!���)w#����6_�	��^��}bY��aH+��MD�ҋ�=`����rI�u��!&��!d$Ė<����`��ka��0Ԅ��-��PM�b;@��E�V%���咧�|%�c_�o=��B�n kf����Xd����P���%[4c�sc��%�� d�W�f��7���0�B,��D��éS
�8�'%񾿟k�`�̳���wp�s���"�˺��� S�2�A˪,�e���#��&yx���c%kB`�F�y�ۮ���~�m7����2AkU�5_�x�i��G:�ں�յ\#[����k�w�R>�q��cr�(���������x��[����^�k���!��e=���=W��2�^ ��|�y�� �X ��qj�4)Ar��4K�&!�c��+�w�;��ԥq�E���;�m1�Y+�ep2�I�$Hi���~� ��>�P����|zUՔ��"'���l��;g�w>�\���f��^���[�['V����'�.L�5�g��4�T4=3y&ptY,�,����ǵU5��������SH����7��p\/fx�?�󻊺F�y0$��EG1�Cjr�Q ��)z�Q�z%��f2�`b�.��%2��F�|�$�h�dPE�O�ʽΨ�P�.(��2���-] x���d���驛�����)�0�|*aC����jX:L蓡*-��Qm�d��{uҬ��Z�siF���x�X����r��t�FѳI?���U��?�G�ۂ\M��p��[��.7r������R��tr/�����%�8�z���=[P���Z'	��u/s��/F z�LQ1#������o[b����?-b���|.Ca����̛u�*�:k�Щ&�س2��y�8�(�=U��Lxt(��PJ�^P�'�jt�&��okUE�kCV��RJp���Ɣd�4�P:��+�I�s�g+P*��f�A��B����������w�:�:]�c~�����w���W�T�.�ܕ�,	��`12�G�߭�m�8�ώ
G��@�:�6�_G��#�y�՗nB4����$?��T�f,i�oa�V�v|6��㈟k)�8���N��Ò��Zh�H޵!�*����� ���c�~���ix�eԪp'��[g��%�Ѓ�i�S&D�v���^\���9thF�G��Kแ�e_V^/�ͶN�G�ڶK��ZEٹ�:?��aя1�<J�㕗����>	ni�ܿ��ݖ3��Ӌ�J�\J��k|`_���f@�-簺�������p��3~�-�N>�hy)�K����z�g�� Q����5�.g5�5��X�G�`�jV/�� �78H��&��|ڹ��צ��$�f�q�4�D�݆ݒE�#B���I{��l:S��O*�ai
��N��z����f���>Gʩք�$�����)�PTUH1�w�(|q�=+K�����n�ۓ�y��D�sZ90��HJS6�be��H��᭾�Y��'VeAh��͎LFc6{*8�})�X�؜���P\wlC)[J>LF
��e�_����xRA�� O�����n-)��O�+�(���@1���/�s���N?�OM��"ھ�B�Gc�Ri2M � ����-�]1w~?˸�S����&O�X�m<您<�7M�����{�,ep�!�߅5�;3��e�8�C�LP��]/W��*�H�E�I�	ͷR�.��8�7���T��R]uޮ���j�Uˁ��'�z���lH��_FE�/�6�	wA8��UD%�4�[ N��X�BzQ�T��K��m���nyX�k_�Y���i��i^��M�-�	CH	_֪�A&������24�z7X���Ϳ�X�<;�h^��Aw����w�g0�^��=o�0ʪݕ,[���IJ �b����ր^cs�ZP�y�	��?Gk������&�H�r"[)λ*Cр��O�jw���|5JwuR9-`�j�
sQ��"3�tļ;f����AC5�9+��%=r�*\BLzy���n�M�{Y�X}�&���r�������=?v�E}�|�re"��ܤy�S��H#��
���x����F�iݘ��:��ٻ�9`��W�a�`�2#g��ty]������20��]O�k��ؤ:�?��1����ӛZ��9�p�>q�����^E؞�c5^%��;�g`L�:�Nws���%�t�й�v�sP��bY˻r��Z�zU�0�?�@'��4�T�F� �<͍�G�͊�7��9���RB�P/�%��*
Ln�)B1x��D���f��+���	�X�>;=��Z ʑ�pY�z�#���˚x�5)�E{�XLG�٫�Y�=|Q��h�8H Kv�JHMכ"J ��na�ƅ��ڕ^h��-JǄ�g������ɀL�6�K\F������J�/�o'![�Jh��DC�����q��J�m�w�u��W H@��F��V�<ְ���*N��>ya�C�uX#^dM���*������(���������`)|4܏��^��-ӷ��w���&}�������VHnSZ�V��ET6���8F��2{��>Jv�]�����.��{҆��h焰׃�mH�"�8�o�w�<�)���g߬�b�W�8���f����!��a�5oI���
��^����AFoS�Hm��
S٥��̗
��a�����.4~S	~��s��Xo���v./�x�P��w�<�1zЋQ�G���5�yL��*e�i�?ı 5m�N��a�UM�}vA`��^3U���:*����Mj��4NW��`-���2��/�Qeٱْ�>2Ё\N��ҵ����ŦDw��&@��k�_��+��_[����۰�l�Q4m���@��R�V�b�H%����2`zk5ܡ��?i�����Q�����p�(u��h��j����6�F^VIi��f�x
��ܨt�?�����M���`��H%�1��q$���#��B�t�k���B�U��̰g�68������u��ϗG��B���\�s�~�;b
1�d~�,�'6���朎��rj�w�i+\Q:�
֜�́E�� ��Tl:�}H�w&չ��q�������z�i���`�"I�!��������'�N_aNj���}�,�ЄoF�����^W#�����w��������*�!)�D�罰�1��bK�^X$� ���g5�#���mL����2�OƸ�/��mK�بקD�z3��{S �M���[��j��	LlD��j��
���pf�����-�޹;͎�O=��7�җ5V/�6J��kq��^4����i`/����ɶ�CxL��RW��#I��:�̉��6s�Yq����v�_[�,}���}��hݒtx�S���>�S�c�qF�޸G>���`z��V�*9���;����,����=�&���!�����jK��t+�B�4,O��`�|J�n*ݲ����Yg`\�+j�q�<WߠN�r
Kp_�No)uڱ�4�n�V�
��,���9C�q��qg���S�bM=&^���^I���Q�1�&F�\�e�R3�&y��s���BC�Q3�๣_� �s�L�'~��I�j��`��L�k���@�,	��"�^�*[��Fud].�p(0(�(���@f�t�XrL��y��a�\��<�G��9,�h�J�o��� �7v�P	��cs/�<W�>�c��0o��	2Q]��Tj���)r�M,X�b�~�S�0q�nD@[���B`υ���:��Z��uB�+$,�p	���1R�uC"�L���qn���(�����>��ߊ��=`���Fg���a p��ɀ���a�f�>|���"�A�ꃳt!c)29���������H���d�/R�;q�����
,��P5����3?�Z��.���85��*P?�A���X��EDm��+W4�U�Mu�*��Yg����-�ďo簋s�g,%]W�n�N�~4$��rH�7���Tq/�(htX����;]�i�w�+�(k�����I�z�
8V�q�q���m6���?��a�\����\9'��5o����]�w�1(��=q�����j����#��7~<w�K�q$g�29lG�ĝ��a� ��q�b�����PBƄ�,�}��NML�@�?��E���ə�bٿ�.���-�3 5S*����N�A��h!������~2%1�k�+#���OK�H�_�W�ƪ�24���i�8�Bg�`Bye���S�x�N���a&.�����7��/A#��.D�a
�~�m�
r���m�D���D����nV�27�<C���F�RS�*�C��\�^&�Y���C�ސ0gܣi����ԟw�	�v5��Z݋�K���Ks�S����������H�����6���z�V�"<D��y7�&D�R^v�ɀ(#Y;e�GH�y�˟(���/�3,T�2�f3Q��<����뷹;(���| ��L�˔�1�J�&P�tF�;z�AG�5�Q�_o��>@��^�w���0�(��c.�*|�>6F9A��������i��)ft@qڌO���eG�N�[�\��XN����\N)��E����Z/4~�nu��m����y��/[�AO���!���)j%%T�mI�z�X������O7�=.� 2�aqS�V�z:W��r����e����x�d�_��r���Q�B�l_"�Q��I8�GO"/\�c\��OW�eAب��J��{8,�	l�~lL�������Ч��/-�� K)���-n���޾�xlF��23$�V�2E���N�����_V�:f�rS��\�}�{��~�u��9�S�v�"T7(TK@{q�i.N�e=c��k�uC�S�%N(K�&��o$.@b7�%�f�Q��]���^�*N�_?��U�$頻O-����Ӏ�w!��Ei�Qy�=5{�߅�:��of��Fu &�B�( �,�z�.���þ�
`xǡ�o��IdY�@a<�y��*�U`2ޛ�I�RTHa�+�4�T>K��iHo`���$�!(��eEv�T��k��_����������m���c��!������}�\<׾�#��L(m��\�8.5��	_V�"&���ѫ�m�����0��?Ex�{�)h�v)(��c�w�!o��yR���z�.�T?Pb������j}o��m�߆@���g�!�hY��9�@����F�G)�ZJg*�u��@���ڶ���r��r������-lTZfp`L����E �WacOCUM��j+����$GN�y�#����XE;մ��ʿ��L�q�p2�˕g´�'�=�
�������	�UřB%9*�75��Ǌ82��I1O�v�哥��+ۯǮih_�8>�?��8t�B^<s�=4����I�uY������_�q��:����#.W	�h�~�Wη�� ��*��^����ᑼ�O2t��SY�H�S��`�H�@ف|������K`U A�{����YR6�`���JϿ�d�VQ��Y7�B�)��$�|�/U�� n]�u�k=��#}�p<=�k�J�1�������}R�e�d��ȕ��&���O�4�e���0`�}��Wf����|���K+T��{n��z�i�y�L�;Bz��π4�R��]���+�I�&�9����(��Ҳ#;^v�fy]v�D�-�rPg$��A��L��D�E�O-f@d�7��<�XI�.}Ԗ��ӑ�"z��{�wb!+N7~����d��U�I��5O��`�+�9�g����[Yk�<:� {Gp���0����:*Z>�����z<M���"c���"ⵟc�t�D�֩+i�Mp������~�D'AG��h��@��<+;��lw��3#��\�ޏ������ �
�V�2�j���6��󮳦hj��iΖ�j0+v�+��YD�-������	I�.0ˏ{T�2"��]ևV��;B�F��r2.�\��{vaJ��i"%�hu��X[�+��s����nw�Y�!�D1�lw��'I<￮(��.�~\���=�Y���ww�5�#W;�+�[O\�G�'���)��G�*��&@Vy(�+�,�Ԉ�ȧ0�b8�����I�]&�H�x�l� ��I�Vf���0�on�cG 횒x΄N�\���ĀcE�r
�L�o�03��P��X�Ԭ�k^̗�c3ոӼ]���S�H��튠���Kd=B�i�9�$�;n�j�)|M=Jz��=�;�G	XR�I���)ϐr���ɧ�Ѵn�٥�V��y�~��,}\C遇#��r�ߺa�= ��M3ƭYG#
˂6z��Cᑬ"Ҥv�g6��d���W��w:�C��k� t/���|��B�8�H��`ʉ�
l�dKK7����ѯk7��pb�\C�� pF&>�Z��돫K���5ί�I������Vt3e{u�(d��^J���L�&C�_͖zԲ�B'�(	���Kt�^�ف��#���zR4��[)BL�'�X�P͂D�]����4Cػ�8�o����8-Zt��벇��)�Z�F?^�[ b���Q�6F Yp�mD3�qGH����r8��{ϩ�X�#!��ҧ��9A����j�'�f�oW���'@~0+��9�����X
�.ӧ�K1Qd���`֩B�t�
b�E~�
6�d��$��8�D	v�t��v�����D(>b�x-������GQNX0�)��#���p:��j�j��ep2{�[�lO�Ϊn7�ϭ]�u���|�~���*�e�k`����p��J�� $vVt�+�uc��8_��G}B��.=U�{�J�ұ�Fo�@�N'���^�P���|�A۟Cɳ�3��ZVno�����;���@0ns�a:>��Z�xu��sK�k2��>����e=�h=�孉lT�� �
�J<��3�N�
�&���h��'�J��,�<�Ӏ�rV �Y[�]�r��z���]^D���O�y�����}�%ZV\l5��oS��Ns �:���#0ͼо�q��%�i�&^h`�Pmv�[�_eEpq���f�x ;f~���V�x���ج\���m�����G�X�S�$��Q<��
�s��&eh���-A6��@ԉ��D��yd��;<t��dӮY����wz|I(�KK�����Y���[\O�wc}�b��;�1�t�Z<R�c>�vL�r�цm3���O�<a�L�?�N�4��?���e_A�G{j;�:��"�9��Ӊ����SyZ��� ̖�b`/Ac����&W��Bm�~�]��	:�\ӱ���h���ҷey�t��r���OD���[g���GS=��m�)�%�󼽸�zg{�W�������"��ES�z��`.y��[��m��&ۗ��#��^��~�����S�
c��E*�D_m�'��c_|��ṿW���R#�<��X�~�S��D��b q�k��+Dr*D��S{��)��I>.bv�<Ӱ�Ѣ���K!6��Jn�	P<��zi�ݟ�Ѯ�h��T����1�&�b��}#sd:i���>9j�8Y��x����M
oYj��܌�Nׄ���EH�t�@|�`�4z�k˽�~LvU�V&�ܶ�
m��#c�	0,�e�%���!��c��'���l�;oF�!�Ɉ+ձ��q!�9TdP1-��h4m�Q�][֨���luY��G�ޙ0�_��L���x�������o�����
[2��<Lz�}n���~�s�0����P����Ҭ�Ң�eV���>��3}:��A��W5]	�K�e��wwV��@�t�pk0aa�t��)�Ь��k�)N
/�f��V��,��9�m�"=��n���[Y���G�`[?W: C���c�^�~���ڞ|��Y������:�<���S�z}���+���ۦ��^X �[�Wd�! �(�U�����91�I�X�tN�P�Q���n1�-�ML��b���:���S�L�O��߁�W��z�Pe�������l�b�׻��,�·��N����6Rh���C	����祑���g"���PMɚqzz�}�w�%ˢ�ޯ�d�bZ�>�\�]�@�����x�5f�b��i����z���h��vwMW7@�HV�Gr"�d`˼RVՍa���-�4|���9L&}����D��4�V��O2����.ݭ�)א�v+�_�#fn�����t�C�n�Mo)�v@���nF��.Mv��/g�^��ʨMLWeI�Y��(u�����q�Lʦ��f���#��smM�9J��$�������k��"��$�O?=u��������!9�&�V��L���Yj�_]�64��YAի&�?�?��d�hp�0GZƲj�`Ah��znF�d�s�����4��j���H ڕ�}^ҔNtE����8�C�o�`��RE�����h&g�?�OHW���B]~iH��4z����۶E�S >����T�	wû�O�uc$��m)U �XIW���Z��D�PK�s%Y� ��\G�I#�J*	�b�OO���q��/BA���� �"]}_�Wi�xd�znSM^�dw}�1�`��K�`�՞G��}�'p�4�����5d%}�ɍ�%�(1i�e���޴�(Yϳ�N���Ub	���$%@�1������bP b�ä�y�x��`��B%�E�p&��%���j��{xެVH��� DF�'�V��4ސ�+���XOj&/P�Ds
Ce��%R�����'�)�,�S%+Q��
ɍ!y��]+�|�]�}�A�i2�-h��Չ��^oe;��sc���A�{|�j�=�V�`�N���M��}�C��-�W �D�⇞�/�|Rt^��4T�ٛ���ڳ�}>����҄T@��F��|:Qe��Da-��=6<tͲ�ݴ�D�x��	����E��6��=�2c���,���Űp����s�w0/L���^�d}�Y�H\�!����Jʾ�E���T�R�+����+�;Pƞ>��#�^�XC���I��BGx�������7�a��g�`�4G��:�d�'���Gj��g9���E-͞�Wk���X؝���|_$�}J&9��ɭ�Y�9���%h�X3��t�J)�b]��Z@�_�$Be�)3�vo%���� e���N�z%h2x`�����HL��ΏDcM�A}P	Au~���ߓF�j�c��;z���c�d+JJ�Q����T���'�������������H\e�X�F���$ �!Є;_�_��3y��]w�����kq�ʭKh_�
k�(o������6r���	!G�F��?p��5�
R�e�qf.�S'&v�� ���.�Vt���Z-Ȧ�)|U���g݃�E��f_���v��;�X
9Qc$��1Ԟ� Q���/V:0}���s~�?3�*�Aj�Mn6{��~�2��p�|�G[fQ�Mq�ll�Je�����5U֡f�x����J
"3|ɸ>yA V�g���Z�,�:��c�B��̉�Ő4;�P��7�8��������C*���ђ��3u�����h0���y ˱}_#Lj�P�;���h��ӺAq����m��J���\K�ܾ��2�!�B>���d=8_�K.\+���Q�gz�<B���d��Sy�[d};��������@>�mỎ�9��f?F�A�)	*Љe� g��ٍO���Ӳ��W.���iL�[�&J춪��f�7��7�oFӠ��m'����������`d���~p`ݮ�8��������U����6S�������v����:Ga���C����vH���̑�*  �ۦ�sW�̵�ϢE�������Z�0���P����r_�9����u�%֮��Y�E��0�(b�̀i"!V���Q���RXư0|���٢�?Ld��Q]DV����eZ��W�E�����M�����'v'��Rf¡r	N��e#�s��%�N�7*��p��
�:�:~"��|��/z"��R�k[I�wC>� �,�b��-�Q��`p)�Ʊ����&^�z8�vVq�Qfb nDk�Q�q�<�u��7,��ԟ3)�b�N$���{����&���$��Ú��^�K�����	8{'9V.��"<�q�.G�ݟ�>����P*3x�f��B̎_�;�<Rn��<��;ɗ��V?��<]�v��8���?�� M�����&c#���s��lQ9����/�>C8�O���>%�OST���ɺ�d�&����O�v�z��7&/�_I�q����8�����|������d�У��+� Yx���! ��T���j.E�u!�ݜw4Y�Y��K*d��*Y�������߰�a�$��(��P*[�8?�`���u�<~�,E���!`��k�Ó�+�=�	�J�rP­�s�Y�Ji���?�T�?�Hn)�ʂ�璯�4��w��\J�8�	�y�W>���\fa�f�����22�C��� �?����H�;����C����Z��|�0��V���a�z��旹���]8pz�.>D�Ǖ�8�ѥVh�4p�����{��nu��?�3�C��b�'%���?�������?@Wٔ<���!��P ZW��8�'b�)**�Ĩ3,T�Nkd�R�'�ZZ'-P{T�i��9L��\�s3Wc9�!E"�/2�{m#ֺA4zh�EM�QN9�{��x֞pcy�74�3�m����ӭ��{)�5,��gY��
��{��"�7��kG��-Q��o�N�.������T�O'�G�����)���ER���'B#:��g��Z����m�9?�,+T#��o�S�-)j@�W��!�f�Ёb:,$ S��[�L�v��9�j�h��OɯM`���
���%u��� IFw$��RS��ݹM�@hS�j���8�%��yL��F	��_CԖ��߭n&�X�E�3&;����H��f�է8��\�6��=��:3q�@�9S�|v'hh|*�A�6;���IlE���!r�M�qR��D[-�Bc�-�:�L�Y'c`|`~�h��4,T��~�r��ms��%E�Q���� �C�@�ąV��y�w�i�8�w%�&5`�-�`P�����/��G�i��ݤ��&��+���;��&�nUZqZt�(c��M�zY;=O�>� �`K@�/uR)*�D�N�;|��,t.�b���j;V����-V"Vcο?!��I������d������]O��	���ո*���i�J����(�a���ne��.�9�;|c[�Zҗ�w�C�$!.�_�w/�|�s�p0L�E�-y�7A��&�8�����^܏���{� {?�c�N�&mER'�����H<�O�ŉu�=�ZY��Ț�ǆ]�WQ�C��;���=�Ǉa�AƔ����5R'�Q#��{����,���h:�?��V}�&�;c�;`,a��8�:a��0?��K8LO��C �U�c@*2�S@�![m�'(4��j!�)Px]����,f�ˀ>`w�T�}�m@�y�P�[U=m�|�Ҷ���?�@Ȁ1�΁�ǡ�ήŝ|�vC�XW���cC��:0F��%�X��\�$ʛ��\��}�@{��$x�gpf��&#m����k��AΈvt@�;酇7����#�i�E��܈h��LS��
�:�����%*h&���ۖ���wA��BT��u(#lk����y,	��X.�G67�<���I^�v��qI��_7Ѕ�Y�*��q�u���BK�12`�FV��:j3�7i����$���i�Ɓ�|"	H����	)�'�V'[s�އ���T�م	�-�CBN��>�H���#����:��0���/5W��<��Lj<�<��hB���,
��C�8x;�ۆ�����a�����_�y}9����@��l�S���R �UN���K�F7�|č[b1���#F��Uʷ�F��z�^���ѧ�H3n܀�w��Ha��b�s��YҼ����@�օGmp��#�ε��o8ӄ&gdi��@��(aߏ����7���&(�&@ ��G&�o�ɯS�"==����z�����7���V7�`�G#���{6���A+2�5�$u��잿��t%�	֒`;[hw�R�������������8jL\��X2�r�I�ɾ�QږyA�YQa&�p��.d�w�"a��Lt��MdC��Jƣ�\YM�O���+7@a�90���6�=}B��%���^S*��u�����O�qK�X{w� ���^g�ovd��+ڦ˼�b#���V�9�V�v�\�[�=��㍾p�JfE�X����z��u�Ԁ�OΧ�C��Ed΋�|�����F��=�j�V���X2�	�L�	=�r����$i���tj�7��E���0��Q���R�
U�05Xݍ��[�;ծ4~���l�r䧧&�53�$���v��S��'4>�o�+�+m�=0%2_�i�"H�����g:�t��|�sV�֩��
&ˤY�aF�̠?|n�������$�),E�wbʪ$�h���m�]�5p�8!��kv��Ď����׽��ߙ�t��f"W�g;��!��b#��H(cH��7��ߋ(����槃�Ƅ������+�H�A>��Wܥ��"�����z~K_9v6���,�9����lƄ���C]�SH�^�}_*��ɽ��$�i�)�����2XQ�a[����tq��W���`��cb,xU��@��p�0;,+�6إ�� �˛�|u���e��6#Uɹ91tMǀ�h_>O٘J*c����C4$����@��̗�-�ĉ�(�1��M.��y��;��ym�M�_P"w�c�b���+ԭe����Α�\���ky��N]��