��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�u����'�d�
�u1�4��s�>�s$,K���J�v�V���_���-b;���\9�Q�����NQ�t�Ft��p���i��4]i��H 6���WH�=�'t��Ė�����\#�	M��Rʋ��c��2f��1�k)�E�*�̱��g 8m���C��6�~c �M��HA���az�g_C�ԊX�}�����Cg\��?^�Մ�g&�]AU�<+z>�� �&80�(�~�>�'�	�zn����a9��q�pf�_7��e	�ܭ�$G,1#�8ܕ&Ii1'�gg*l���d��n2��5����j�7���_�ۑ%��2�a3H���q��"�AV����r��z���ݍۨ09���kd��S�����B�-m'Em-Kۘ0 �����AwĶ�`�r�^td�j\���(=b5?�eښѲ+��Oej3�o{şrV�M)�+����]��Q%#<�c���ut��O_j	[����({���N-�ڧ�� b�q��x,��=B��H.����v�+W�r~����n���i'�+�`P�F"��mI�'�C&!������� �k�����p�.="��K2#��9�\��嘔�l/�'G�b�3
#(Jk>_� hm���������*e+�Sn��BM��ex(-[�$Dck�r7���ʭde1H�;y����Aq�\I��i�h��j�p�� �],��$��E����c�ӹ�����:o�d٣�N���b���HS�4Z^T�F���_��!�e���U����Ψ�aFz��^#��r�@�+.�ɷ�$+7FO�z�3���2��U�}�<���s.�4�M��+`���'�'�=�qlNf�6eI�4��{�O=+~p���j���Hk�����r�oʓ�����We�:����J�<U��91�\�$�Z�8I���w�T��@Rd�}bRz&�hՂ?�4@bC!}}�l�1E���9צ^gS�!'�|�Q���Os2�[ve�Ƙ��Gue�+�fqnRn�*Q�p�܎����^K@��c�p���V�j1~���/!�[�ǥ��<����#hr�aSbk�=��̫|X|-i»��Q��_��XD�4�����*>�F�aNl|��.�x��om�'NH���Q۶f׮�d]�AXT=\�s�zG;]_���`�,������P���I$�y59��\9s�������9�;:��Hf�Rc��:٩d����B�(�.p�7_.�a�ܟ�=��*��.�0����4g^�1�*x�q���̎0z��X�ΞXf���䖮� 
����V�a����lCG�75�������ާ��a��ٟ$j�_������I;�W�ب��к8�[�~]���.p�J�S*q$$�kI�EY�k��P�$n��!�	��A�t��c
V�;�l��v�^��Am�[o��߅��B�y	���'/�V4��̦|����S���MG��R�y��iv�D�U�Hr�=�����Y��cd>�ҹ.�����.��O"�m�Q�6�7����+�f.�C���W���Xς;�|�a͙��O.&N��tl�� ܕ��G$�6��j��^!
Tm�*������~��ذ�R�ln8e�~�"~�	U�&����bJ��>{�P�oq�9v�k�`I�L��oF��5����\e��Qs�/�X��OD�HT���%:�`�-'�Ǭ/V>���o���0F��<L�Qz�;%����;G�o눾Og�}8�ʃ�^��ٴ�@DԵ�F�c�	]c�}`�y��l��V�̽ �?�|�GV!���6o��?�2��Wk)���;*��G�iւ����H�I;�
�b�yl})�A?O�8G��b}��ʑ�m𮆆�[E�[ic<w�K��-�5�)F-�˱1�":JfK�r�dzL���7`,k����O���X,�P�1�?�����G,�@W71Mǀ�1�G����<��̊#�H��>N��Ә�B����'ZKbIx?���.������l�+K̄�[��F�`�m��Q����U�p��Ks��N���Ò%�A�b�>�B�/p�A
�]J<�ȅ�L`��(#��N���Lp��>��\.E°b��"�C���r�m�����gmv�ܟ���7��;:�<8Ƶ��)� D��G�C�3�`�P�C�hX��4>���֩��I=���r�t�3��� 8�` � z/kZ����)l�%`{H��>RR�؛�3�n7���5^�=W�@y�s)�N���;����*5�]\?Sh�Bm�2�X��fg+D�j]�K
�nGVW����c�����P�㚌�����[����n���O%��Rc�f)@�:���wa?�I�p����u~?C�����i�%!�OG��3	!)|Z�������m�X!Be�!���E�]�bѓHH}���J+�(���K�����CY����o��M�N��0_a�v�?��8�.̲�>x��Z'�q4�*m��yt��e�a�
о����lq�WI�����u��w4Y+Nk�`��_������Y���_���Ǵ�r�j5�qn�K�AD�wW0��ZU$�X�,�T��K,�JQ��PmA�$-4(�V��a����jC�7��А"�񭢪A�ߠ�5A5�]�(������Ek1�ڋ���C�n�iȻy����N��a�z�ZO.I�����x�2��La6�@�WpKہT��9ܔ'6~�ǣI�TA�>���QTx6df8���z.��&��$�_�zP�g@U�y�q�uZ"��M:iw���!
6�5ǵ~�YD(X�E;�@��s���ln{@��m��q�!�s���ͬͨ���"���ҿ��Ko����b?� PÇ�U4����q^Z�&긟
GȂ�-q!x�
��*����P�H���~A׽\�V/Rxg�����p���q �Gvʺ;�^�tJ}�!�;�i�Q��簵�O�s86=�.����v��K�G�]ZJq���ɓB�y��`�k��A06zNY�|Q�0y͊�g�Zٶ��ǃ�X�pcrik�D5�_E ����;Z��ߤ�;���"7t��t���5�U�ӯ@��9����7�}Kp� ߿�����(42�}3�FMGX�G�a��1dQ��=�iR�������=��j�k�Gj��'�9�Z����l�d:/mV�0tEWM�� vC#��7�$�uf��U�1����"
��� �=7Wj��ݯM�6��U�w�b\�b�S�A-���t�Ux7�����o���Ŗu3��=i�z�r�����`�	��3L?l_о5�b��n`�+�V���$^!������h�����L�+�����j�rn���[B*ISYLEwt�^���f���Ӏ�t����	��Y�P�?�MJ�Xul �n�b���C�͵Cb�f��cA>$\;g��9�%J"�.�I�ݍ��}h������R�{�R��{�YR�ucŖ�aT��s#�s�-�����ٛͶ���j�D@{��)��!�OȖ���b�w���V�p>�JO<�Ft2Ի�K�i��GֶC],�h'�)Ԕx��1g�Y���������ER���c2t;�#-���!瓞�!�o�D��C�1��1FUE�~����-�t��b7��1VA$H n���A�:�qu5m���u��\(=K:���5̽��F�<��e��SB7��a���>�ڔ7�'��jPl��#g)I�ػ�g�7L�������5e��D�����QP�n�l 3�^Q�7��)<%߯ ����2��"�l�|
�.�.NUI�T]q����������ņ���t�rƲ顮�Cz.
.3^2q�Ĳ��R|\x��3<7���F�,�1SI F�Ha��?�oe�q$�@0j�Se�c�x^�z�w�`N�q������uia��m�����'�>�@@m%x�W8�-0o6L���$�J�ez�[�J�.k��jc Y���^���d''�3p�n��=�!k�r+�_��~
<���c�{���{�a)Pv5�)J�2^�yV?Sw���ũ���n���:t;j������sJؼ�5��g��G��p�J�iŲ�۪�SE��z�ky�T����2��#�ZH1t�M#�a�}Vl2Ǜ�ϤT��\�����+k.�볋�V��-z��C���P��wh-󴿶��������}D�<��h~�h_�HO�1%�A�8C�.�@���V�:R��zC�҉�6W�Z�M�Y�C��G;�y�}1pj���\�,��_��,l2���L�@)�#
FC�o������o�'n�U� �!���T���,2P����Uqu�ykǹغZ���[��Ø�+��|�]X�0!���o�#Z�4/PN�iG���19�8�7br���j���<�֪D�A���$W���E@B���SxT�ͷ+��d�B��5
!���b�4�!�� [�a�Q �k�/3�/Ux��p��8�T���'RK��^���^�2oG�O�>O7���Fꪹ0p���� $��Z��5�' S(C��W������T`sJ	<�r �zwS��=�q�A<���=�C���Ϫ������Z�h3