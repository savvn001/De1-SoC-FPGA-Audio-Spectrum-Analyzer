-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
INP4Zw8FqLGp6K4QU2AHil84Hsc01tnDUTOqw5CF9qYxYWZEhTu+uzX0TjDQjpGafdpX19gQR4sx
a9B7PD1AVpijbUPdRZAi4BF+KbP5GeS97yYkacd/y8tS1E+xvtex52HMN9X1aH/iACDAAqxG1qLV
CX+8jg1YpriJc/yd0pnVoCDAcKHlY7SxqlskV7B4dYFErmtMHdECOr6GJZZXx2YhvsEh85bLNt2F
yESnuNRnANWnzIi7AfpOt7qjjKgLzd/dxs9RETcDdsz1uPLXx0D9XnfAMbowlOKORA+HNr5nA56J
kuBoYwBY+VrmR5z6vwYC8drZu1pS47rLXuwKvg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
2op2r94vuEVreouboyr19w6BTAMDXZuLewFECG73Cn4ODeOpdiHEcLFAgRsRxamY/7VeJMMjhx4G
pgS2KTytEOtVz6hJNdttCTpY2rDMwGABmqgiB0acGMMd+zfetsBLKa8Nmj68jOJsViGPSWs4z+S8
E18+7bTUKsecJOTb5jlBsA/YSwI03Ft/dpO3Pbb9OK/2Yaai0IGOTEmD2kL+jUqCscklCPCcCHfi
pXxKzhWCH1eUqbj/QnKD+5wUQkmmpriV6wdbZm/5jql1kjDMsPcYufI10B26fdbcm+gYNvTWnAky
y5dCsCVuDqkFAwBjgyQNte41Rboa9u/kFX1du6Lv9qol1ehHLkQ6p5KOm8dsQ6jBsN8SWca4cZKi
WWFHX5Ng/yjQ1N5uOP4mX38R1bt1CQwwKaKLSjwmRBUAcEbTYI5GVm9omRPmiNBcBvMOuUbS5fdS
nCPKy1rbd7eCtArNIGBkFXRhiKmnWq7RJatJux658Y+geZUXnIfjzSJqm1XJN6T12x4wd2A1Epc7
hywT+PylV+pRiGXBaYxSzNj78g25eGVyZks+27hiHJJuUSRAtP8vqSEvSaK8rF1Zvohz9ZJfn7wr
DFZPIrpeY89AUuflAmAMUVV9fFY3Eu9omHVCh/5IWGmQ/DrhyJxcqDVOtC2VHoFHxKDj7dm+6qnV
C88J9mJaWYbon6/G8frLKxPuTU3Uu68+Uip35Px55q8zJknN3ZUI05qWzSZXVUPIRkQv78jGiXG7
yA9Ki0YFNNDDyvM7mhqEJE+dFUS13qYDkxTg67w1KvcjDQQIxF3+HolWqAiddMUFTvGQMx8fRqgn
DcPPki6t24uiKKVoLtWblDnb93qMf8/SfbN+JySaDWwdkxydB0AwuNMQgFb0YPTTAzdeU02vQtgf
kg2kFJs52c/Q8/Pw+Yx/UYzT/9odCRa0K1kYGqOf/O9tyv/UQYl4YIKKAsIHLW5D+Vk40oAnGM/l
E36zv+fIM48P0R6SixDR05E1Iwd60RxsWc9xjiRh5w4rF/QMM5xXDuXhwPNpwYOdbFFRTNdpmXID
RVLQJfYEjfb1lHidoNsNNTv3DeyqngceMsIOODpAGLWC6Hnr/Te3oXFNLBcTL9/OZZUkqD47gkHg
xwrebUt55Dtd/Qy4kyYFw+B3FeSgDCmO8z4OeXstEfJE7dupd0f+UfvuO1VpwmoBaYqI9q7XiuJQ
OZ7JwvDfGA3JIXH0eLxcXchgKdqHLtmuoiKbN/EOAf8gvZ4SHaNfXV4nKNuMQXALgDNoavDVn4jV
dgxSAOY1JeRm0EmB3GzmA0Qc2uXSyXmt8ve+xNUNrmWj474CJLqrgigfUHBc8dhg/UB1uH4C44Ba
zimKEAxciXv8mGLHyfTECLiHcrukITylRmTqz0afjKrxyd7XyOKvrQN1Pyyqs58pbizafsEdoLSp
T/Cfv1SJaPk6nUdnnhXsNNe03peirvT2/maj5iVkfxA+NG9ILSs1wI1x+DNbFTi5vPCe+SZzQXjE
RwCdFTj+8laGjE8wctZtdNoxe1z/AgUshMFNWLQAl5c8h2g32FRCID2c3ne3IL6y1KgOzG0dlDJi
HKIbL3u++p56W3jYGjCZfYFML21xYEnxUd0BFqvMLcGbmWWTSU8YoMwKj2IPHDpMS3y4Mfta0CCd
yhYXResGg/kB7/xHEO9KOVrjSpMtqjgXmfy7cF3mdl2f/wTAha6rWWwPekkMXAE4l37rabo1P2bH
dcSjJYSwaU8uQKXUrcot0sh0+DXifrv/XUxZRuZg2eqAcj1UvI6TGHL1H8ceGR3Fu/0x7fPNlNtf
ZHr5se4miLDE3canGRpQSXhM/qEnVdIezC78kK5hCvZ4iEul39/vpCdlLZMvMADyjjmkBqGIpkGL
tuMuibLqWM70txFoBbe3yQbxa0gAuDftOX3uUhTYfP+aj/5s6cMZKJdkYJKr2T/dMSBmUVfMr4oh
+bGVkCPsKeW9Rbbugrx5tjbbx4oH4JGa5NL5NRDP4Jh18zHm+1B7cgQhXuZBK7yo6ieh9qup3kZO
8aWCwKt/39FHntyMxd6lqYRNp2ay9v58uCztleWg0jMtjiJm6mUwyrXs/jWeqjUs9i5RrxlFuOx/
73DTPc7T+fTWo6MMYh+E0x57VHpEExEM00ncWpMhUTnSmyqdZrBEKpYErmRCtbfnzpa+Y49Ks+RE
5p+dp7yLcUQ3eDDuMhf90NrLWDbCpdOn0aFS4FHCyz1X/VhhdHysmd7p81zUkPShdMirHNFpGTdC
K+NmVRb7xMEcCcNPmuXKkeFuabPVI23gCezkTCN6eaurB1ePtZtro0OKfEhsFUaIgWkN4BfznjXg
L1slGCgieZmL1pXVaOJ3kpkckRDyC6JdzJZiKYwNC+21phT8J1WyQNK/1NH+3dJ/5l8SiOOyklqm
Si+YLYQVtm8IRd7J0EgS7E5NucYRS4Jj4A8ttHIeVmQcUebSSySvvfS1lNPTI3M+JrQBmmXaulub
xeEsFwIwfs1rr6cbGOBKiQSYwJju2E1Z9HUjEdSA1rgzPb3nGexLQapEc2JQKymZ254JeX6Lro6+
GvgGPkN5zZarXOnGUw1fQBEHr781j8Ro6iTmPhIUwpSbDXefR5a3Jmt0teVajbPdsXD6CdE+e8AY
zlqcnsdGDn8ostqLMP3N/L3wQgeZ/Zmzr2WT9skaSxCISGOqwOO7ein4x2UcXYm6mvKV4YzlqfNr
PktCPY4ynO4qZocVsk4VCickx+C1C52Ei4sVjgQR5vU9fi9XPXnn8jf1WICtxP70M2rKuuLT6lhG
31/QlFx4N/aqeu1Y0UW8D8eIUxAJXdMJxF4xfmTFjyhr8QcWbbSmOSkwEafl5DGh2RsJlzMWXkH8
y/96D/AdduT++OgOb09yY3H54AUZu/sSmFXI/Rjq6l0j3/4acdw1Z176q7/vQ37Zp/k3lgrfXIOM
tE8SoBDbVsqSBjfsEkiMChn4dRuP598t+Vacyuui1SGIWOILbUSdRggrCBCPCDwVzUqo+jN38Xgh
j3nprjgztXfnHL136nZrl47U8WiKvlzeyH1jLZph709Lk3b8dPZVGytmn+EwS4BmGRyNA2UfUlwT
rwgrKrruTGmKwMij2vtg5aoffB6eOhlQDKgqPDyprhsPbUt9KdSc1a8Ehh+WlhRTO14j2DnfTMpO
CXX9Q/0lK3kpqDpUph2nlmrr+4uevHrW0ypS+7kN9/eRxlyTmjsbk2hHhs1zp8Zr8JdUsi8ejWTY
cP4wJ7LbvOQBw0HT09QyRS8AZGjbZXYRMZUWfthzlKKXsHh2qn/TMw7Ig97ejFdAkqbqf0oCIXKP
XWvhT87CNUEcgJxNIeYKU4a2IV3E/o7npieX7ipwYU9p3ZcorIjku5o6gLlnfsEAtR/+LR46bXQG
mso+PMuODPsgQRiTFLaV8rM1PrjTr6v02dUTHttNgbHH/vvM0qAvGvYCkZDqALJrdCYzfMJt5pPn
Wk9Xe1Wru2LKkAQST4GW8QZJpKCYLT/xvBJfGruzWWIq4O5UQBVzxJKbGfs33aavvQ1isrEsxS+N
//qKp+LF+Lbe3nTB1EereFBtAnbjuoYghC7UzcGHQaobleBBKulo9MZreYAv2DOKw39mEg7F0uBx
pO4SH2NhPkZLbsYhOtqJ4Mo9R7ART41NJbp5SFreEY0Vxjg1HWAszewj/r0YeK69Ag2UI3ErsVwz
9b6lay5yn6LDanIpj9EF4R+c5fPCEZS5Qdnk/FKXVBPxoZH4RlD+wGnLuu4wItkt3XCaNL5d9KmD
g7OvpWFaYx4iiaVF2Q1sBmEmNK66jOAPfLkUMWuNOujJE1ksdHaMU6INCdw57u2abxikaCgmG37W
5VsgKCD2fORrrIS+k1kf1i67r59SJhiB+z6pUoa6WgO/iVSr32zx3dUDM+mX9akwpZjSjFh9WvDi
pv7EUXrd9q2kmw4DUyp2mbXH8/7AbN43fuq1bkHqc6MsQKwHl8qN2GkonIQpknomEBc254WIQFxb
CuFpsMCQNyPxuwnhp0ar7TtK3fLusDzkZkf1eU5KAvLoLWOyXInZ4ajY0G1Z9DUNu2iWKXHPZLel
rSBlz4eWuiA6M0LdjAT+vbuAmJKTSGJ/rBo9fkWYmu+74ceQ+56wS4UPgOJX+V2QNXJ6N0fgyLsG
pnfPSRLN8+098StL7H9GrWROTa/ZffaMzFBEyCNqhJczYSwkvpe2e4WE9qPn4H3FqsZ+NQWqfObe
xbx0nQYXCYAV8vMT/eXM6C33d4lRf+WpS+o38sNKjGCZwYg/V9SIeRv0sThwb/ZwPAStqDfNQ9Tk
f71HZg0qXGPcor4qm0kEP/kXgCkEQVcwmtHBh7kVA3jbGrGUOrlMhhUtyrYgonx891NMMQp6jFN0
s+rvT2i0auLndjjTkCpU1LY52Hsoj1ierktljH1s9ExpenUyswiQlLKK0O1V4nKWcwbIS5ZSSi9a
qDfeDOr+cvThj43KmvgXKLm5ZlUEGOX7YZmHId/R5H0uheg8vAV33rkwvj8jdVwmTc3B7JLmBmH4
bTosSVNR5saUdTrBD1B7qy5XnaoYs85XmcCWRbMGnfA7FkwMotFZDE7r8eDOHUG/j6BirR5mbq+/
JL5czt+8EjS7Y25H6RPDB9GH1qPHo47tnCvgpUAkj1o+q867q3A9RsTvTBEb56OjboUBWoUdaeBH
1IBJvlHRROd8LGOrKJLQF+3MPFD8N/qKTHEFxHIGPm8ZBH4AzIiIMKHi06XSpofwOKYrB8phu6el
hlXA8fvz/7ythTNvu/x7dxJvuObO+ts82nC7ra2PZo/qdi0LGFMsny6IjusGD7XfpEyVoq+qv/8q
Z1Gr8MfZ2+YyjBdaNKF8OGAkpRSVvnv1UIvHf6ePNBQ8cNLNm/6ViULXM2l176VnI4r7LFfm0DCA
O/MBPvmx7++OZhArLigzT1mpnS+GO/Uk5C8SyUmLPcOfrpZ7wdEOOp3CznKyVi9+CRl/UuD5jImq
/iVjFgvgZ/iPXLXEI1JiH4SHzY+CXFRDWToiBk2/tkgFqL2tWzU9L3Fp7BxMMFUVEFHBHhHORcyk
PWJXATQ2xqWjr00e5hFla04DtORXmZ7m9MzVgtz7rUaukhDagWsTUvY6M6KHqnnzbf4p3nkFdvRx
tZYCE1B57kZg/p/TRVGDrjhNxcigC/j3TqjE16+4Ap/smEb/qx9W+UPL2NAO7R2MtbZTCWGG0CfD
0EqO/t7n3ZzLj4Y80p1BMRftLwwNVr7hvwSCIWZx6/2JLKu/E1GB6xTQIXh/J1OA+QzzMz6JmZYS
r4s7FREyhUPobFBFjZmq2g3JyqjxxAqRZzLYxkfif8Q8lF9Ho3tTFx46TPBI1UK2bve8diMUn70y
jPhbfbbgVWrE/ZQ8dQP4uoPXuxfuMsUJOUIB/x5+UqClB5I1jkfUHIFxsebMPxVW83FvRKFz2ECj
T0GY0Vs8tzHdCqvVMAQRKbAV1ISHQCWiTEBdPWkP9rCG4h/SvSycyu6hFT+/VvqUG6xDSq5tg44J
AOlKpxDSzTUqIZqhvQgpvyLsoHph8p6XdObddRl8/tf7ODZHgVE877l72Bh3Er0Wx5DE+zol0tOj
kXF2ZgfIL9Er6kBNUdJ6dQGwHb0W5GGNRiVJh5QbGyjnwd4zssc+bnbvNPXyC0VH5mFpr9DkSZNO
TV/y8Wq1nMAfy3LbTuo/Q8cVFcP7Qaz3aM3MHc0Cf0AzRB+5X1VYDXyuhDechrkjdQkseifndmdY
Lxai3t+KbvrqI4oXSz0phDRSQSARDCJ/mS3UMTerFXg+TCXSZdXA1GjI33gv1Br3KE0gwwhLz41l
+FM8IdbV754Gn+eG6tUYOJu4OAI+JO0QkpCqQIBNtyUTj+7TZ6o6DTUY3eIqcrlShIsCb5YpHrQn
KS3PaPD4+FuxPveZrypADgmn0D36SvBM7jZcTBfc66ir6Je+rJBfkpIikimQo2AnMqwT0RUUsPZo
+QL7o9kfEkMbFUWSsSM5A/eqezmplYSfKz+R3JE89tSB8+dKyla9A5dtgN/Rr6cqtWeSzFvRCwVt
2b1Tn5uAIu/6TRXDk0JVq0OB08Lma0hlQJfrrxqcpb8doysvXtrjkQJe9EF8MSyy9WygessOtWeq
uCha60EFEGWXd6tL5k16SHHOgiNEUJOIYni2Q3X5LglD7sVW580bmtQVpeIztUwaLE9Z/hKstg9i
cVPARZhCQhy4gEm6EnTt5C8XwJm1q5/s3xy5r3dbGT/3uMuucxMHtoP/TIYLUCM1wAoTw+/cydzy
ALhA427NnlaX4XXARuew8MbPbyFPM9nu5WT87jHCAOO0lFkzGmCdne5sZN2EC3DUOZuj5NRXu0mR
xKu0KVPay7+NNH8iczv2P15CJYIokfQAleLi+GK9hWY0UEZFBqRh4H/vEOHiAPU4BTkTIK0X/uIB
b0m5/UV4K0B8f33x+PesDNpn7jScPIAPLyUrTHQwofAinsiboRInj9OS30MS9z8xoZAtl8HLpUfl
1w4S+cVBpxR+ra0IG9+0V1PWpB4d/pUYpDx761nvFKqDTvnPga/vr422e+om9z9i4T2TaIxwvejo
QXpxeZ3h+/+79q50Ve48eU9qzEqiq9NVF3AO9RY2B2WU7YziGP9U8P41h1Dt6TuVvRV9OOKE4ICE
l+U3at/3F/1OlXdE/zNr3HiG9rojBCWDGktCC6pPFymQ5yg6Q/gg9N9wDDPZSPpD/dXOGOcb21oI
MejN3kpEXFCMROYNCIoNN1XlaUqeVX2wweMSNwNdMJKLekKcCch3NEAPmGKO1J/G9M8yYBdmGmE1
+p8ujg6cww4rOkOCUJS3hcYSHLBZArYv7hcL2/VecjsiU29g1UjR3xCWLdz+VPsdKaRhil7o79+L
6nyB12i8pvqUuq1HSQq0HpADhrXueHOy5a+IMmcHMkX5PXvtjBCSOp1aSCUgdhuRMNdXA0T9vXRI
2PV64Yz6RpWe9lasA98FDqcGBDjp0kY5l7QmUqb0kpyCp3+otb8K+SFdmLxihxVQv+sR1uzv/Mkv
K4d4s8V8SDfN4NHxhLv1MouO7ou6FIZpast065G8BeZWqvFgyyKPhiiR/1UBrQvnHgluDVzQltka
UU1MMUwi+m+UaX9FrdXwcF+Eo9RhxXuJpmeQRplTkVJUifYzj9qSjaMc/lIKn6J0ZN4x8iAz54M9
QT7AqD18u+7hOjsyLOvkHX5OWH/LPAKYbBcLSck0DMYZj9VvhpCEq9bey75qhbJbawEaNTWlAwLH
hETi0ZsTOOmDUF8Rs9I3+pDUGlawPhRxQZuTSXK1IwDrJMkpzUuNgitGABC/TgvyUAWRzpwwskZ0
DlRIOL+wy6PPAoFJaP5qNKbJ0fZA5uCkeJXyU7g/irQyBsAIej0tj/rcy4dGyWuld/vMA5SNlRsQ
fUvkdXssGgtlK1XadP0Zncw8S3olQ37mlBZC2ZSkUH72NQgOBkvgKFDZwfrzA7NRXXYS5770dMox
S2v1XtW9eU+YFd1DPfcACuT3FxTX6wdHHCnD/G2IkmKkKj1upxhQvNVOyjaFAAoj1nZCWz7SRdFQ
tzeu+uvelQ1BvE+pE4k7NQ4YhnNitc7trldf4Oni0D3eevbNRRIL4bYVpHzDNhZfL1iraRKtfhQp
wyAR7fYoU+T0t6TQeThn89nbqCBAAMqaYVtGZgbE/NHNKDoQiPde3H7Zx5VWL3JuSuG6rTbEXKwp
mkdREmivLWHQJqUwu80dOrtn2idgT48z16WBrpepPoxx5xkli+pW+LIAzg/RuWZz9O9bAdAzvpel
ovBFga33JeB2utosErxIbP/piqElAvDh9cAo4hA1nXfWyWBAVKJj/WTcqQUFM2BRPFTtjzFosVgM
H+cLqJ0V0/I3FRDsEfiYDqbCohb8F7SdDzSCDzVA7/3qKn9VNcV39GFMRn/CE/uGg+5RSeEIKhE4
JIytxeRob/cQYUzjEB6PqConW7lhTQ/jQydr8sL184WbscOReFcJS2EbpgVup81B0Uuu6JIcsJ14
Xi0NFki60GuHBGTss7cWC+LdZ4bEG1Cp5V1FsI9m2WPGGETEKhAD4vgxmRgBF2j50YGSBRIjUnDV
OweSmD8q0FPdQjelTyhGW8Ci9YMzX7BMAwxPsfqePeJFolq+w+WMguVmNjcxySifTDCczDE3YnGj
XqIGjGrJAgcturuOd2iwTtlPnBnXuRN6vyggmlsanAZpNAd4aHMu11wjCs2sSyBS+wJJ2ZrQAQ12
Tr+/4L2MAKOz/g4wYCsqMaxTWYXRR7pZ64d/L9epPDjv3yULBUCFQa0IAwHEb74NHGSx9++wsloM
QLGQbAKc0rlXEWebwdgzRLlhf+3b91lcVACItn96/tgxUGd1O5bzmYcq3Dn+jgV8bcXXji+KDQSn
E4qIpAZDlCOSi3Inw8dgT6iGSTmgggsuCeh5hO7dvgjp3KRQuDLqnwF68dKL0NN9Ml9TvJj74T9x
hxnRW57cPFut92qv8LIMM5kMF9V+heeRreJDXTufSNli8Pp1CCPLaF4QZZAhrmlg4gG+xLy4o5Uk
+VKF9K+YfMuhEWzM8jVzfivcYOfEkUUxEtQoHn6y5YQU8fFdtybBEXEpOAzYVtDfKzH+33w5jEVr
wUtCuj1m3/2gmLeaXiPS+vPK6f2WKZ1ABLalwk9n17hh/27BB0xPy0ANoN4I5oKIJrAjnizshoML
TYKBqBPfqpNFxAPCjnO8KqsTRk/wrETbyfMNqxGUaoTA85LuwK5J62dMxxUOF0cLPg3o0QKDqnVs
wJ3ICv2Do29ncIJe/8zIOEDKsDkwRKvEdl37EsJwk73Y+2H3nFmKzJhUEP+qdXt3jAse37hGxZ6A
mkrV0E0B0Cmt8ZsoIrjBiUWjmsmzwLE2PcNm/+4DJ7XSFuh17nQ8fzZ0u9AWDywXVaDb/S9l0BLT
5tyh8o6AEQySFOLh765pkEpjTrRk1524tbgm5XIpLPhwJ2+VSNViMOO3u3P7n4HuK2mF1R2dbBz6
rJ1z/8zY6MwIW2GciCM5YwWN9MTPyOsGCmZDrO1AuJrMSrWB+5isigmvmrtwHhvdKIw0klzmLYs6
NY2ll7gufJi30jWXloWTxQSLhfgQpGjO0g5AkPAJDtOykl/PhubqAJOAYecXK76ai5nDXi+sU4Vs
NOwA+Rvtc3LNRGY67sQnKdiTGYC/oFBErIYivf9KFR18gBmCdcHQGyVZOLDn8V8VU26kuPBqArGP
nXh0FvndHgg4+9nQBVM2kveNNAyuEdCrpApYYQ8WFZGzU9eINYJAfj8R7mHbDiIOvOrpjg238wG1
UiZit64VSbFQeD6YHOQG70E5shzJQO9G5nkJX5DVyr5sHgL7m/dn5M4WrDhOJnDPRvzdEVoRFXlR
+5qKhFCK9EfA0OtufnYLzCmkRzXcQug0l7qeAiyQwhfZmN3wOOlX2RYcCfYqdZLg3TU/+UBdAR0e
3NcDbrga67SGUzXtt4hN0SKqCTK8X37hX/oo9QJbTU7Y2g6rNi4I/Mb1AKH0HcO5n1QfrDEv0kAi
xChdWbt9n87i3+FUKimlKrFsSz3XIV1eL0QA5E0sOSGdHd1huMkI2tdkCKwU7giICtl2JmF46R1R
RXN30ZmPPSh6otnl/D+1WkJMo0QrHTz7Yuw3noaY6/x9QpE0T5YAWMY/1ADkZZp+zmAjSry4P18o
fsmPVSgn14Kbj4++VUSz7D+ZB/riHcEAm1c1Ng5/3aSeVC1g6IA0QEOoaHaOGsUJ8HQcfTGLHu/u
ffeKAP+hg46ehLLgsXmtzBlXxSMKwyE7TFxYrYb4iSWW2qiU0a3rqY+X5kb9ZZHAt2cJzElIlwjj
8o0hEeCzYyVj3UTPGe7tKMrZ+xrUlBxfn8NBtqmQneO0ElJ/KO6lya8qgzccYvqdKqsLf3txze+1
97+epyXvQWPineOSY/UDTFONFlawmNrSKXAqiN0APQ+zOGaokUDnxGt9WYd6yhBbGzJ1Hzhc9P90
mPOrFEdNCUgqr1QcNKgWE4/gCWOOFj1RT+lKmWybtuk/xaOI3HT9fcwqLos+4GMeyiw9hxk4DGSJ
Pg+o1WMlfFSwxcOzS2Qx04/o+Mtb0wx+eK2MVY//bnr0YJXlIhUAzuDxIXB8qg2mTWUYk0S85pio
IrlfNey6dPtc9bl+kP5qw+vH0dwdCsVWRMVFvBId36P3bekV9/Eie+tozDrP4g7ex6/5p/Q8Jqyz
2C7gI7m9WzV4vRTiYNvY6CqauI4Mmgz1r2tm5NyPOuD5ePMAraTrSw/GdO7Eic/iNjAUVUEN9Sh9
zOJHLVAyxi9zDIa+gQXz99NixNi4lhcF7tkjBR2/uhHWEYLoIY+9ctzGfq6DaPlQ0JfWbJl0h2PN
jU7xQYB5X8q4lDX4dfTNgjxU/2r3HPa0ktzt6cJzxf8UPfDmfGetVr3Vny7z7soD30JZv9k6w2hb
KImFLI+7wTSc8dqMxnmMkpJ4XOmyr448AQq3Shl0MIJndhXwk69Sn9ngikVhgZ3nYFt/0DPd4Ylg
97r2JFxMO0aI8oA89l2f6OOjkEOVNByZLnS8dMjIUi5rXWgUniTX196rSIPH1iQ8VhGTLAGkvduR
fMF1IzqIHY7MXeIhTRl8Ks6cJHg9ojH1Ug/jGJBpdFKUKhBW1KI5GiiLFDHU7avSU2xz5HTkZ08P
h9YsggUTuTp3A+eXdYC2DRLor3u4d2gTCHhzALIUw6pleliBh8PzSdxhc/hKU8mcAKnM5LEKhTyU
pl3YTymDmu8y5SKpo+6JVmsvMN4v/BJSr4tfmfr65RIKE2vSIqqALHtDOVZlSxwsa+2gmElXyoH9
NY4XEFrFpmPqXyxRDwMd52+693QPoUOmO/Kv/E6yQfwShHHm7NsIAUCkNsfzYCfDdDHVnp66EMhk
WXB0KjgoA5jQgqiXYXrQ5SX9Dn2X9jqAi4Z7gCI1zHwrfBNwuZyjULKkDUMFZNchAPWtNRcw1wix
OnB7KSydyQNpuKxqUuALd56LEkabVymKaGpxRg+x8z4NTi4wufj4/LbG4AnxFkOqFe9uMrk7a3QE
xzwDIwSzV8zJ+jKWLgtsNQzPUB0JKEW8TpkYUiQ4UOm5fxvo1QBddWSrQRP+yNTRs9U+3rIXAIsO
H5QKsuU1NY6BmXm3L775luUx2Yzq4cLb2k+QKnKoSvy9+/z3lllZAQWl/q3nMSLhBtKsBk2mFnf4
ajFw2Gnl0pjp2s5vAmwn6zX/xlwUJONq7eHqETX5kMa7QDxUiiTr2lSF86sdQsLWKH1mukqUEF2C
Vrle36Q8uQ36uiJhc9dJNRSSMYmvfF21cFylcx4OC2fbmSbHzScigOf1B+Ibx7OG78MvhYMy4VUC
0E20+5Klgj+u9Irtsdqww6yJiTG+XcW90Ss4f3rVWJhde7h9QXarKaQb99LAnTOTnTfpBrPyQxfB
KglRbGpuA1yEDPK/1FJq9KjD4/AMu8iVtrob215t+0c+YT3RziZAPDS1JDR7eoY1dNK+S2EPUxlT
BdE7uXIlZR/ShxvtqPx47m18+r0XljLv8HtpE+jWuGbH3C86wAuLYFktxzH3zHfs3j3yiUrLvGeU
mrpT7VcGg5kFbswmrYOPjKE1xarpP014b9pHptIfRUKXOYcIQwf+1c9X1Z5gt3zg6aE2IqaMhutf
M/haT30IKpzN7OXNg5zgnP1fVLKOzCRLyBm9NBFOvLTI4jEhuiVaswxAbwzPFg/i3ijXup1OMb0t
FMk5cdbhemeuG6kE49SUtT49T+4YIbdeXMREsEN6HZhyUrjnyMjvXmYfpdKTnudtVouOU4tVZ7BU
Ci5Jn5o+reg7EoLQPD/dleU4SjYaLatUkNZB4mUsvHv91RGYLjRl/X+LSUJqhE7ZqGCkXwTYleqZ
n6St7cfVwKmt+FxysHK+RMVn9sqEmhopI3UETjXcO2sKAq/hFo4i1YY2RfXiGP9gf7HLU2D2FjjB
oFidTLGe0MA4ZVWNsecCdBFKutaZokqg3tTZCnKWIa2O7v8/Jpa+pGzwezxEMvVs/x4QQ2sAklHy
PiTdHkrSqkTx7uXn3Y1LDF70SuOFFkDJJyYE1YWdLX8pJcVrbnG3jCMdLcHH6WqBOI3V7w9M48gB
TPAiB2mXsQOpZyr09eYDIwHOuxz2LlVXwwkNw5Fao+QbotmJsXtg4tEDlZmb772n3x3uonPZY+Oz
0cd6nWAfm8TLe3fDYx51EFvbGTXb+l+0OsheHo+Xgx3jS2KUeWCVVpTuTS6uK6ZoDzY73R0HdDlE
RGRxhJ7p6Nt0YqM8qDE2j2pjM9cxBA5VNNIAP7WR0jJQSUEce65rojyG5EmmeKglL4JKN0oKAmQV
bt3XoSLMDuDZvlpHTW36BuFVGdVI0I4HpFwzSx4E8SsKbQd2SWSbd4vnRzpC9EyfymfGVBmlPuL3
joB/za/50M8dalF09aB6RNpiKBDoChBV2cuNiAFdgq3ddPvcm0OJYm5d1bsDYCI7nbqP7jtFA2ZN
ZzILNYaPeXP2MsUcCweeYH/ZPGlNOG/BbHpwlAQ8/LoyccLkoOsE9iTtC+Ry1WSQLERROPZ/Ehkv
bR/sREAtTXoBDaB97DOd8vvdHRDSjtjwj6E5aB61eHO0MDSHHdmaHyYDKkjMkFqezYtEhcK/bhqR
bBD1lGRhMBK026AMwssFeUxC7bwiZSqa6EpMC7VDoSMKCzEekjJ24DvVbabmsPKg2p/elRJ6HZ4r
8k9B0iVodjMY+G0q06+hn4O9nuRjpYqdezr6Sdd2ZGZEQ8UWNjFOLdYkeMwvAiWNobpy+h5J/UxS
YAjfT5bakWVLUmqH4xx95gNOhHXvbuKcLJm9GpGOLvm8e26RBOGnKmzx3ag3CbSf6SsTC9FqpnQK
c9HdfQdpvzX2Oikgsdn4XV5LmfT/NQtG02UdI1QH21vgrOfx2AYFdc5BTnl2of32voGFF6CmMR9h
HHJ5ZBNu+4iIVZw3dcTLW6VBnoqvTwd2GGsdewrXX2nbrCaTNCQHPGGpMESNsIu3bczcmIbpxixA
Tn4ncZ7FybRjJdi6PEUyqOW/xEkg1Rai8BKOcXlCEX96NpOxd0csdGw9zYv1WHAkopxi2XY06R2E
gua8FkSEpnEjPzEfuewDYC+P8jszmG8WG2DCJB47rQVytpmV02MzHmH8AAG98nGJ+LF/6cAN76ON
VsDwb9xf6oB/nbKnyvcDGQZS7mk90nujwMpInxt9xgURgHsj2gdi4liGb398uLXOM4gsPLQpUFZN
PfrPGkdmZk9R8BDzUb5NOAI4fWgpxMWWL60MPzqGiZBNKv3URK2EhBX/6ohSpMJbfzdWb4xo91OH
URTb0H6lDNglxCnJLYsPS9jat4nd8LtYCc8/vy0jOHJti+FQEswt7/ZnzLDnw34yKKcVHt9nEL//
UhTitoP7cueIFcbfyUvNfFjmm9aAgPt9cm6DNCIa+bFMgO1ekaIsSJ7JqPrtfifhdia3ZF6Gm4Q3
ncgyFvGYzwe0bYqgnb7EOrDudoLI95asvxf3/dHCibHqwDtfHL0Tsauf2Js989Plu3Q4T8etRxPa
S4+qlyJJCJCt4bfym2cEUGLEKTufnFJgvSChK4ATNL+9GAn1YMxKRLM2GLdV3p00tqfAL+1IOQbk
mwzDjPmBBsQii4SbWzPKhY+nRoYayZZwzCmuh8h3AX+Qw4aeF9cyMFFIqsEiwhxJTDz1OstmlkCa
29qUwll1Bnx4PiPjUB4y8tZRcb262NDBnuIyoVOoysvPZh5Ioqk2N4Z1jZom09vbuN/eQd4cMkXF
PXGPeh/M8RJd2OwWNbw0Pq/0WHcYpbbLKnCOCoO8gEj1bG3OZUebQUkaVZBSTRw+evvtGPY9sFQ5
k1AmVoklDS6D+QypG/A8+XXTWO0XbpKI5Wy0NHXLo9R0BM74Kw0oqG8GLdPPa2ytVkvglCaSt3mw
RUcaKUV5hK31eQYaunXSB0V2vkUIqyVk42c4M0+KcDXTSc5IBlrOSoK1VA5OZgcYe9C+xRHTlYOZ
mBem4BAs5jmeh9SNh99mjDJd0/P+e2p2XkiJdrM2ZmpKGIRvRKhVFyX+sp5SRgTGit7XMOOixoiX
U/TRwPqjSUhsBotVstezBhLBJKDkzO38yv4oMW9uNJa46YOYnrzLLNvbYInmi/OixsiFOyfjoKYM
PosDeN84sGo5LoLhN4aS7gfaFSK4sVuftVQhJCddxN3gU0+n+kOhtFUWSb/o5ih30yL7XLudyGlL
omTuQtR+uSWOPQDtzraKyBmeY/DpyWqeiw0tHycGhk7v2NT6/VHl82wHKIxlxHOu1HpZ/n7++vO8
ylsSRfNyNJLjv+IA4aETlHDoxMwkj70v06/DX0URSZUbn++dfp2mvdLns+g9YBFvWHNGFn46zVnW
klInGqts1WDeEAHH2sA1p6VJPqQbB9vllr98t9S4m0sfiPfQhm5Q5DDonStLHmSch43zQn1Or365
CsUcpsJAToufcpzK28YdGYlucUCGkG5ZIwDGR8ewCogEb5135Psv2HmpB3yvI8KtQ5MrYYQ2yOtl
kXJrWKQ/8bmaLmNI6QKszxOdzyH7nAt12KiMoeX2MUggf7GE9xfTj4brGjevuJW/44B8cSMiS3KD
XAbJY2RPYhjGrJMmnuP8uayIVB3Gxj1eNP3ykfXqltBqhj1F2VfHyxmxow3uNjRxsACot6xPbLlT
IsxVerHmRLz2Ca8miHoBASJlEb0IcI0mIocwIbmvyo8Y2wQlyRMo81FA5l+lD1SNaUAoIzWmEIpw
O5uqOQp3OHXqryV2flUagRScSZuG0adwTaH2mDVQbFJf4WmBbD6Q1+PX3Bvq3rgK1/08S7K95xeS
VuhIF9IoypM8rF/GtWZblOF+NFzCmcvd3pAKOinh9RMb5o3S7vh2Sls66SUjY2dC26MB5FNnP0c7
p1l1+HU/enXP2vYsq9aonV3zIYQyJDO4fKnVBqkRA15EmKk1lfdsDHyPCrGCjnf+kT1Sj3lTt7CA
SsHQ/QU8d4gtzUNCi37AsXIsDCV64AbpkImsYiawUFlyPeuA5IuVXgXHZswOeOwzA6Weh2lBc6iw
PLOm92reSWMQpG7l5lr0DztxK9/SDo0ca6B1c7v1LeQ/0jctDQtQ+P/xo2LcGbJhMUYI9X8PNT2k
oPM5iJQINckImrq//SSBsZS+tAX4881DeM2p+3lBGrPdz3WEAdZPE25DGBdvND/ukd09paXoHytP
Ip+qPeJ2/AYzxI4FfIQCsZp2sBoK/4abiKtX86Fg91kcnYCxrMmOpm1tkF5mY1yXBTiN419Otdtr
yXZFzWjc3Py+PmR+37Ycj0MexaY9NMBwVHPHUrx7FTFtXqIg/ppwoDtGDkR1o2CZpOu/Tq6HPPSf
rPmvIuIfoL4Di/W8DAJV8hIDwau31q2qFtJ2N2YX5em5dSHNWrb0YdchACDI9L5kG51Q86xAXu2g
ehR9UjujkTmZ8TzlEctxGxLNrYIRGjErSDPY6Z2Sr6MkO966URdZThotqSz7+c+xMv3hEzf/nH5p
H5k/7V7DhsH0bTfqYq9kYObduRIddiCQZjiwgw4vpf0M18a82i5hhJfw9pVwq2PeotI5ALfSFvE4
3O63LLHXb+aPO/Q40XwheVFWoHCJ/5Mewc3Zgg3IQjVi7gluZUOiNdfsW9NpcwFJ585c3dQgdynI
FJ4UM6p8I3ISln74nXKI2qeuuScR6xBcQmYLMFncv/fIgsMkEBBNRwkUt3/EAnu78zgv2GWKvfK+
paZh9u7qT/bZYLSzCKpkdrDfT+bKMtoXM7wpax5Bc3bP1dA2XVcrAR8CmD08tASrOygO19Z+ixHR
ZL5IynKeQQ+xgLkfJAEARQZBr/N8iZkiDbyaQYKefUekJLktakjpPtnIZkPhj1ZyxmCTHhG8d9fV
VG5NaUBJITRv3pHSPIR2yPgCZACWj+SNLuo5tWxfpc4Qje6lzcmnxTCKAqILxsHWD0HUTrR+gEEE
RAwCAAiV0n8j1e6r754xcLlftvxmVx6jmjRaUGMhCu8UEFrUORFQxZSxM6zAmp9KDAv8+ZpKEQ3f
cRo2vp6hQ9VRxorFY/hcdh7lSq7FnSotTPejW36EFR/waNFWUtL2z9JGR/UjSHKEgrqdqo14d4eD
TfittKgKX5nCbFNvFBE+I0WC+CQg+ms8c9TyjJ17Ga0QFBgAz4MqMYK6B8aKIpvEWRnHmP470m/K
ZmXN8fbT9bEiN4YE1+D5eqe0T9/T+5Q9g452jkbquuMHHR+FfKuLp5NZWkQXOBAFbqDC1YdDV/Sd
XBmqwXKGhiSoQ7FlfTQnFrK/mJJz8Y7R3qUZzIPrl4WaSgtTSD4z3jkdtLhkziqHWdZ6q+TaJDLa
RIHdX6PoCfHd8RoAAKku4JEEIpTboFpUGehEFmkMqRPJwFaQz2lKkCrbAtWsNYQUSfSHpvT2Zxea
lTlJ9RADH9K4IDIqg+kySa2UgdYKyc8mk9i0NkXULVuXj34tv2+lTgxcAIcPjeDCNz7i6rLRPUSr
NBNDrsdYDsPZNv6+uEK7Xjzu7DOOUPdPUHklNfymh65BExdIohyy59ZLGJymo2Vw73xyiO8bdfe2
/6ZoIezYJNbDIcE8VkIINohOGWgk0I/7FqIvmJEQZzQhGcxNnFAagwTjsC3/aHWTnCA05TWLqJkM
MUw7tADkgHdd0g/yXklvt2SYETAPmVyHyVEdavwzIvqYjJs9A8Z+c9kcj5F70A/mmb5rbeNksbKH
g1Hu27I6Yyrr7yXHuzDstsjkkz+CUDjsJoiOYNIULdqp2Lw0Q3UQyo4GD/lxtz39gzAALkZe1qHM
pCECKCkSf1Xsr8F7+0VJUTGERUeSZkQwAVQdPG5XAvLbm62WV/5YZGZXBbnhMyRKq70UOyLlyG03
mW4G8KeZN+oupF8fs/kSbiGH6bbgTHTq3C9EW25Dm98K5IIAJZkGLQpiDgOpy+K/fdDtXErs/Cms
HfR55CSq9XlgrEijymhSyjJ2SSPxok8Dniulv9zfeSFFo9D6/9/S1dUCiJhg7AD2NFNh75o87ABY
0mq4y+nTvyLnLrI84j/HfWgdeaIxIcwKMC7Qzknajc5lnMbL+6LkreaiMTKk1TfHPDxf6nXmo4fI
lRjaHnaPXS0imcyymUMYyQ9fKonkhXoIkbinl6eVFW9B68zYjWlPeheNdC8+qYUe5GwiIL//OdDG
zjuPrUoilF91rEmC7+Ts46Uc6jlwGZeWYNjCPhcF6jZJneZCcghrQ+G/tjHbDwhiJ7ZkFI2omkdu
x5ul6Sji2xX/5JKZcDlD+2cGeSuNl2YCG3erSjtvbmC2ROKi89zOQEk9eoMZs48S3uUSUnKw8PZg
F9VBAJljbJfWo0SLlLouzBmg4YfHF9kmkjNVHjKDecKnaiRhz3MMhdHJpYMVyqSRRN8MaKvpRjY7
gDl9DRm4M1ExVYn2mePlzIWSsey/n5JWq7x+kuBAgIBdFdujcW5FXlJB/84NjJmhK+WXQrL29cPf
gx8+dfkyGZfijYAUXEURfa9sy0m0d9ckv3AW6S3tYUjKB6TZmyai9G5I91033x6OWfZFpPQN5ITC
0JdP8m1mxzB8W1/aw7VVLY87rRQEUidYtXGy1qe1DFteA7nD4N5/goYEUCC5Ap+mevqV/PZRFFO6
ZQZXM6Dw4lmmKCRON3hOebIK0s6IGv5ijvU6UqOKiDHhSg7C3iONmf37JGReBjZ+f4grTMGK+ATO
nXpetULt3q4nN4sAWEwJMalF1zelj7DTt8wn0o5RIl7RGK1RSqdGVUKlPTcCoejLQ05xeaGebvdY
3W2GBRPbt2S57Kq88WLRy/zz3xN2/1JxqAeP6YsekGVQSn7Hu6N9tmtldAfbgvJtiB1MEq/DxFFg
0dHt9uWEQ5lTL2u94AW/58aV8JYkwjvwSSbtMVCOlfOxwFXuBx+Ju7OyC0H9WqwATZKgjPAuWqrL
hXgINiC0Elh1VaBNX92lI2pwdzde6YNVfSy+mZRFTHcBtxRZ6PCOvTu5Iayh/vswLSYybpZeIEmY
wvgofj51m8RAoLNWI/AcfhYyvnEaR75a8QisRJyQEhTYPJsgeSk+KF3H0M2Bx/3q3AZ5khq2Tayq
UA3m8XA5eBwzpBqAjVWYX7KcOLPAYIU+E/XWK5IlMankUYoV42GbIhMMMiYv9GtTD54YTBvdWE4g
iKIpoPOt9++Eim72U6GxacUviTTyecBMc9pwIdiF5Hu8eXM9m6Li0qsOVQoyD9rpxOYDTnwGQ/mM
CZBQC34rcg0NJKlUbiU+FKvdL6Z6FHczMyZsnzVmbawoL5XgPCI+YM477f2L+jdF2jyryQQIUgrA
DgaVaBm8qWNWzx54YnRSwZbRK6LOUZv2UP8xbsCOP0n4Dg08dqAchu2NzoCO5yVoB3ObvOsqt2L+
ovWNz3Hc7wr/y9/hs9mfRw+0QVqj4on2E0oaSSSfNTZJP7toZem5C9szLCRJTPIbAgq/4mbZx279
se+GWslFJ0hcZ6qSWNBN6r7L+yIyvxZPshAXmdcz8RALUPOxkc77NwEERq6IYu/ZnR0OpOsQ9g9C
EvPMxLOJguFgcyDYX9npXWr6D5sCMtnBs7ZEr6lty8tIku6NX3nKK8VAZIrUk9WZ05MGMwNiF8eq
wJWzcK+jypCVtie1ULH3R88/Y5s5+pFBbQKsw7/h6lHbY+MY97OxmSYlGm5kDhUgFcJWTqsLKANo
CNyGnC2uNZULi8M6WefL6+KGoomR2Ric8QH+b2rQhhnXIVBFsXX2bjB6Pk/hNNiuU6Y/8aD0ds/n
9dVO7wTl7efS/fpoRhI+PKIXcYe5zP5lypzfLG7hefrgGnDTszvCHehx7RYgRuDkoWx1kcQi/iu4
o1NuyjCXS/Hl48b8cdu3+2cpwmWTRUeRYZ022D3wYpnuVHFO8gr1Ds3NTLo6OBrdoC2mbeQ6I0qR
tApHHG7bSDVPdbghQSZBDQvyHfYcIjeUNjaTEjnoEryF4XKFrOcpwxh4GIUTF/fzsBpQAJK+OvHN
jAN3VwSMZq84sn8R8o4R6uJXggSdwmDzthwEO/OBJXDzqKxzHmdoLtZ6JBKpUD1Cb4JSgez97+6H
XMP872uP5pMdPFCId+kRdzWQO1KSRgHAODYOylURwDQiULU9RJ83/hnLL7T3mfR8XAdl1dhQzni3
q3SiNciICDqtxL1ylGQ2J9uvb46cm7nIyHghMogUWz/WkFCcd+f7929sSWdVxs9iA07OXIOrpEPX
dD0LpCTct0c/zBafeWq+BfYXYmQwUmNdWxd9a6uqtHtwp/WavHLwIda/wncfsN1+JIzF5F8q3Msf
B1UBI3GnsFYejFFhO4f0SkgIwkN/NPXl2uVTQ88RyLzi05t3h3lxqoXhFfhBue2JBY2UbpC8AQvd
bTCNsweMK3a2CMZdAsct6T1kekeS55P3gjKQ6Drc+wJI3KH2HrkDW6dTfvbFmsxa5PvpNl9xW2/X
g7dsivzGpdyQZHFSdbV1sTJgn2oJEmorc7H1oaE7XvoYA251qRIfxXkG7ElYuIrXX4A5CB6fsQ7N
DucBwLaDX1xT3QvtZRnqC/To2oJpOVufuo/Io+nEW6Bzb2JryrSgNfenfzQyeP7NMtflXMBJSECL
aRym2/AwTwE7/ZlBmtANsTYlkoOGOXThSrNbV+5NxSa+Ad8VyQ/8gBSy/Bt9pS8RxmppJA+5qMDJ
pgc09j6hwmGqXzXThfUB2em2FRq/JeGItiuW6qO/9wZGwxh5jwqqVRXitwJr3KGaSak69nFX7oQ2
I8Jz/V1mmbREA84Uk/hhKU1My0ERT3zIOTn16C30e5tZxUaYulhkEuRqgceTqD2nzDddWNXaCNL2
LPAvhPPdJVfpyun8Zf3rcJKs0JaTWkRNRFp0gjP0VgjqxSzipodEi9zymxbpGnPW6128cvh/mO5t
1mBe6oetEj4MD60l3qsLV0ObiT5Tbe2KIRsWg3DuyZ0svRMVdaJvT88kTPHBWSYtkS0H/KrZCVUs
YlSzKpKGrEs8+hKHW9eJ3TS2vUht4dXGn2LPILyIATdBCH5ihDlxWc6TKegB3pCajOiYmLp9l/Sy
PGTeUdLYWNLQKja6BHd3YV1/cSOqCmlfcdj639MP3yJPVQtOezPxHyIr13LWtret3uFCyS8VqAVC
NIVEceLEvfGtzVGQVPiU/xLv1O2laDjBTUqQ35ouDKJouPS2QNdZwHaWSsU093sJLkT/anojOs0d
UfD2ltGoIgP+1UEphl8To+IOOGDElW2Jg8+f6D0q1PbLFGESwLH4rcIXmU34T/PzIl3RSVXWCiG5
OJjHt72eJZ46x1VP/fc1lOJxeS059UrBuKUS6ZzcNHPokdhkg3XQjt5N7UlC4m1gir8/F+k3UaCt
rZ7fXvr9frmthEd75TUtfLtK9ASoL+/9k/IliAMjowPhfa71Yuhnp16kLFXbIqHUD5FezkppUmts
z7AS8HKqsfxHU2urbuEyc7YLqoGD7OvWjghGUnCqe5EdYWfWvt1Ud9Kj4w0mwgd09Lce+Lh9EE4g
/wRlIpApfJDLleGXCKHT4gX2L0Fna0EvM6KQV4y7YHowV+oJ7EwpfPvJ7jweflowym6Ie7myBgHN
g7ERrSjq31K5GZ4dxXZe4/vUvC370ktIK+9AlsESsXjT99NyvoUDJsMbb6QjsgxQmtLS2j8XrYTd
4kZ9+BO6bRhHDTzTue/+lZGxcKzdMh00Zk2dpfqYi1s6zwDEUSt33b2NUyWVBJLldvZYULj7d1uC
C6dJ8OJK2u+7vmmx3Z7jBqDE/8CEyncKSB7eXat1VmZkW8UK7u5wFrCbwkUbtIj2OuqBbOIqguO+
h54BODMpFNfEyY4DONRtaDy0jq/E+AbfwKPqXTw7Z87xG10zHGXnPYVDGQtSsYfNmHUEfGqBoEuW
5st/FmrAIC47tSL3HRfnSJi+BDfZmonn9ejoSyAgMdk9bfki5QHzBk9fuJyvpjED9v23nvKi/8Vg
RpWaM1mkHeTrZ56eykMFXHU8nVHdCGyQTXBewnBmRZ/BtngraA4+yPmE+yllVyKeAh/O4bH9aKPl
WFmYHjV9P3XCfRt9wfupBm+ooWfTG+i/rykIfyX6YAZWxjWGwbhPGl7zRK0yGBdfzKatQ/39wmTT
czyUsICxddzaeb6QownieyS8upfcLphARh2ddICFAJ0PMWgtLizDMW72jAY1wxJYD8+aXfX3GqqO
jIGgu6rggzTyQ+RlDJ/3O4LqV6+YbBrEYwufR+cYoUrN0YHr0Q10yBDyeWtQ8B7MdZSolKAEY0tp
iNfLmJ+oU90s5K9ukhU/i4Vj23a0aAfFYAbS15vHelChPwVmlucku8D+j4r29542Cw2059GcfhkN
Qh0EG2wLxQtUhEIySnDqD/3sbqaeYFzGyS/ELPSz9JwVah+q/YZ6Z38zo/7Y2U0k7cKJYghEYijJ
f/I5REwTc/H7eNmDdkHPyxn8PdRD3GjBsBMwjZGpxhU56yGJ4NRlbXq0iYqtyoBl0Bu9jrGDmjjD
IRtPD9Ox7FE3aDp7K9PzoBUa+ZzDrRhzQCvowmXrFuhaDRBMDhkziGqkWvHnxx8fIe1fJu2bkDLZ
7l0+A9olJD91x5uZ4LK3ptq744mkhngwj5erZQyGNLJnXIZ5zu0BV3xhSz1mw+QHAhpYLy5ruwH2
nw0Z9GdF5dCAQPrlFdvLRaE//tQjP2KXRdg+iQRPVljlds1r13M429msoxdrSNlbcCwbEf7ZFXcb
ayyfJL2I3gs8ZRc0Q0ImyjP+2UpSJvbGTKoA8yViPRyzkJRGSTe7kS5sNLbs9B18+mUFUrPoMZA4
fIcLKmEL/u/NQaFf8KFI6iGZ8NNnis0RS30mQs2/NJI8O9R73FvfykRE8sumb5S5piCykgQFzIk9
g8XEt4WRBuzLZY0fYzBo2nei9T6P1+u2CWw6Hp3sfLrQ/xAKxke+iDrdIrCmVP05biniI5Q+1p6O
XXq6mrvGnK+azhpm6YCYh3ytxcT+zAJY6yNlpJoOAPuEeRh8nzoSD9o9GkTLqIonqlSYc+YoMhAx
Y53nwd/iYEqTl2bzO0qD3F3MWk3TYvDPLJ6cew1I7T4j7M7Wk0CM3uFGKFtBRst0PdpUxuBmwnVa
8yq4/xbSWO40/wls0Ocr/cf1TQTVY64E462BhrPbUnL2RCGfgdfMLskOQhU6mkVFtTZjpCBm0T5n
1jmDXjjaWbwIVW82kGZMuYfsax1NN9GkdV1vnbzEy+OLWjCFHtT2IZS6isDpuU2nVzVfi1g0X3Xn
aNGzZZsFyKPyprziv/HOY+gR1u6UV88PC04lD8TPuBxW4PVEh/7bELSCwRQ9NfgiAnMbATsE3+GB
aCZOnMJCcS2bRbcRKM84mS2E7A5terBBFgm/d9QMS1zWQ9S2gzfkPTE8wizjf34CElAIhImZrSl8
YDt25wOMn0iPpA9MkWPuCxfMQ1vVM35001vx2M4cnQDOJsb7GGVTiGA9MDMHDHIACdJydxG7c9Dw
4mqCnRI63q2ePwdwRVdxdMv+eUVlIt6KaHuWpkoqqawbrA8a8/fwHylHKfQZhO4F14yIKVY5/LNM
gyZp1Sx5rsmNpHgqleY+bXPRgZS+l+Jfd57mejH5NIx0AMafZLA7gwATfdg/P+frPA0st6ARWOek
7sfogm6/d9GkCTdZsEnJW5txnEZrlcUJ9LIT68q2XM7xE1r3MIzEoTUyqatzucts/T38Vub+U87p
BVfes0hsm3R9MaUlg/sA59C+HD3ErIOgWqhRY6k2EKAMenuPgihyMtfa94/nwU94jnBx4rWXLftA
OQJq7AlqotpB06w7UFaTs59RunC8a2ccKUozI9i34TzF5WFqT9yJzWXlSrUNI8bWvapFgSR6PgHK
Xqm8/l/YE61cJsb6zmh2RAGHTwhLf8QgbgLJqz+7ByEVKE1xz8TCQSqsaKojjWXBIXJtqLcXyV+h
x5zzmeaPnxeBtuQAjCMjfmD8P8kHqEP93joOtXWl0DCi6yIbftI1ev9q9KSgMfoMyjH7ilQ1w8r+
P/uFv1as6rCozNzS2IuKjimziRCNoJ7w3oo4YwP06ysA+jbhtxv/P9l7ge1NkgjgpNMz2I6OVsiw
8EhDXW4FOLbnvwGNVFeP3wHEEUpykj88yjOJO70vnmmGP1yjfgIM24EhUcjauUUs04Ej0Y7M2WHO
UHUL5tvX3hnFisJoQyxh4zfzdlRW9bYNQVvNAOQiK0ANt795MGtD6rlm10kE6+cztbp4KHUUgNYn
n753HrFbFkg4NAf5ImfR3I2LGudy0C7/+Z7BlxKyLj1SpHxwTRpC43KJ4cgcoalrY1n//4zquCSm
85KtR8CSSrBvbVUvP6S+MZVz1675UrGzC36YQTECwIHPUGns0CjfLxdTk+p8konROsUATlJPw6vd
V5OciLERHlWNYJnyje/KHhORoXzyGF3TPNmdR1xOKnvHcnfraRM2MuyA1oATrs80B2ODllhX3Ecf
8rABKJDuiSm9CbxZZGPBPesCfKQYwXm2K3RWDqYnnLrEgv/xjh+dgBNcJvtEoiDq4Czm9HEbhb/C
bans4E9/IPDlBfjYcAPmSpSKkaoRqoS658KztKNOAbCLDksAPitg2+c/e4FYIIAEwzR5VRNvL1mb
Ss4bzRqAbrf5KlvieUFtHwpY97NDfkv+Blr1pGoKwChefHyTDJPWWtK3CTgS5/JURASCRrMS4zI5
MiJbEv9ErCfwfxIOEMxIPuX/3QooCFnYiH3EKWiI4AAGWbpNIUYfeX6D0WST5d79YnDH+JIcIZEW
pMjpO+wKuqxI0dbdVP388bS1RRZJX4x+PkTjDMQNZvh9K2H5LsXlxTUgh+i+jrVyeCt6sk8hEnjQ
iEdgk3DItAh0w3CgPD236GtghSubdCCVB+18LDSE79NJRByjHbrDKQ1n5pOpG758S1ExYuPJLG6D
/Xf62UDcyklHT1L2617Pe7/iZNh5LIKHOlOA5HD7fBGzO+80Uvnrmk5O6yMYxYrmURE3Md/TmZPR
UuHQqUSzOAipU95h+yThDitnpof47SxQuVPRCbHHmKgzYRdGw6FRi84pI8SblndXVZhVjW6Zyozw
CZO/C/psIKiwKwz8WTdc6J5WJMUVZ5KysHZkEzeydy0nrkLt1ujL3MDw2Hc6SefILvcmrdvHlDj5
hND9dOWPDCRNxBcu3Zp5IQJJq03ps1qhvvE2Hieh2HO6VkyW01rw0EJOdbxyRKS4v+xTliqaUnfN
lbYHg7J+yUjKvFDGRaGe2KIpEgZLmcpq82uAtEMw9Z0XmLPpt3e91643nHdJHMS+typJns36HkyZ
7SbW8xzkzZyrAa7cfV8bkMcLAWr2JlAo4PgADLTY/cxnXpW0Zl1Qz2y54kZq2wHgRYWtS0bfv+oQ
WW9tbcxRp/BILIPX0J8dGaIEo/BHhlQPUP4gSvhadFQl1O1PYfl/fG/iMFe9z4Lq9ejQCs8QiBHn
hXR3HDWx6bFG3yINrsFd3rwVX4paL5LeyLlZUPbGJgchDngCwKnETM4ygCpn3O656z7ToKbSuwlM
owmFM6cbQk3nnIBzCy6hO43Qe4fIZfqwcI40E0HjG2QP1t6zX1f0jV89iKLYUnZqI4TjKsaXX6Cm
5yhcERuu30UXj48OTkMJvVINVvmZFwjlC9H+/wrJAUi22zSGchE0ENv4ioI2llvv4+X3b4Cs/kgS
dbPq51bZo+thjOVZq1PE8R+9kUayhtNOe/BnXufZ/utUMMoiPtUUL4JgnCilJrl9G7O8v9PfAidg
/Ql1nq99cZoAXxdO7mRb0eLdNcRxZ3OhS71YBJSofF+vfP3p0HwGR6rCSwlH8cJaoQp6jplG7SZ6
rW/4RtEbwTRNXrSvxpqWSoqQwnhZ7Ofm6SfZ/nbbL2bkCthvU9v9sf/D1KvLq093WKPRfgbaQLOn
IHl10+KI7dc0N6PXlmYeN5MDD7DxiyWx9tDgWy0fwjxU8mAQuU3f45Y+RanaBDcEkKIcJ/xx/LOZ
3Zlnp0OaGDDH52bSEKq6PelJrQTgqSZU73wJ7szBFIjH6pyU3MBDHdsyVboEsJG/ILe/G16+imj/
dI0Z8VyNYgc+XMzz6ZRQQGIl4kuGz0OBC6uQdij8J7agznGGPTT+MDhO3MkPa+bdHuvxI//8/npq
ddm/lP8BAIi18clWgWEv2cnEIMR10ZLVnGWWZe/286BSJN9hXyjc8xTRcmOX7GuCvWjqggI42iMl
eGBHdWNj9jTYe7mlTc8kVmE9iEOEGTuPXrRwjYOGr4r8uvcQ0jZBj2LRZl5zu50VMU66jMkB1yWe
uStboqFY2un9aC5L+UC5KLqbBP7AqRzSTUNULFGbcBcABZnXpMHLynBzXg52vu+NaExwKArTCqTj
GhjGQrhXoWZBMXrudVqqJjEtTAJI/Ew4F4S8AE8fLWDOrBDUiCOXMZqWGGrKbvqCovPMPun94Ljn
lRKlXsPCjCr8vb2OmUuYGoioq78xPMwbvWhWsuFGizkbnGw+HJqJ2WxVxMOB1Ir9G4Iz74dqJ2+1
ijnRAjZtgtDZzzUExRXfIA0tQP6/DTNNifHkmx/vcqICeJOZvMf9akpN/KisVfKKs+2j2jTsnH7u
4mRk0p4zi82qAbPotIfqz/auqBwozfrUzwVZhss9204WW2khd66ZPSGPZDL0wIx+AuEG7OPhZUUK
8M2ACJk3GQDeg7OdX94JnbiRGSrTZiTNTEXV6hXj0BOvGeFQ4XkHL2WFLjGuTSsITWf3umUbrpIf
DbHw1nnsI+Ezy8EyYojBt+K4QqNOzddsQWvdijKGA161l2hL6jAhuxsNNNL4LfbcwoKnVuWNgSjJ
8EA+KhlkT9VkI6BlI4uIjdw/Olg3+5OaLAkFWSdq/GMecJkMHYmFltg0/k97uFni7bbSAC8usCEc
IfsIUtp07HrRo7go1T+toHYzwpicVHyOF8is6revjTDo6GGbzFDKcBMpzJLThQejgA9aj/3gKxdr
/aGA813ewxBfJoqEqf0vMacX1w+EnnEeVKknXdxQM44Z9fBr70E7AjhI1IVRmqq/XmkqRbdwaYLB
MLdWoZ85j7v48LNgsdbzGu64v2DTQZLDG0QCcqrysavoN/rr1fsj0oGajRnOdG28XzLKK5J7TmXf
841AfL/T3/vT8mrEJYzAA/8m8zmviMZ9qq7vq63RpERhtZ8YyrQyhEeiDVO3hmkeTsBhO2FO8UdF
jGSJ0N/V/TvUDclUTUbrD1Fwq1xLElyy9BPjAa6Rr9y2+UNAPUQhLz65V41C5oFjsz/sU2MHchh9
marQDpHg68okCwMxqziqWpR9fincmIzM+yDqMgn6yliRoCPtsFUbKaZ757qXKeC6ibTj0M6VSLje
sdEaXcB1AkwsC2ZQlD3CzM8JZUXUJNzzT9A0im5Cns/lwyaRLZtx1OLGd46pfCia6dpMv1/CuuhF
AHc+hLzITF1qzghoBW5vFdduI5kwcMeHwTnjoubZagT7SZ5M6fZVoNOpy8cdR3Ad71mqEouMa2ZW
SRwDxmcxGNnn7m6XZScbRKgmA1yEigM7UQTrtGszYl9iUJs7TEzWW80EQ9rP+JHIASDhWf2g+l+G
MA0DWIimXkFmQm/BM/4J6XwCwTMpkqNKMh7vQAbUwHPFSSkwuGVTlyg2JtZsXFFqSVQaxrqZMXIb
WbFC25mokrSXp8HkCktPQRhtnSStlFG2a+sFwvmbRdzqCCwZcIaMP78Ly43aGR5DDSIJL13QJCAa
1MREEWHYbO9+ja2Viy3+LyCDmyIedaiJQa5Cam4ZjX85MphvQtFpcd1pD2Ku7GVaSf/OeAj4Pkdn
lS86HOQ8zYb7x1G5QNDjt8mgopZB1cZDBo5DzqUL4LsH4mh0ob03WSGy8YNqMyRpY10ggj87ysWB
4W/t6HYtqEBVbpb2KtZgoBuuTPX2xlea6vqGZimiolgVh6bDH8EpG70vFDgKjMVmrnKho5L06oWZ
sDN8SoAK/QmvipJiBNyAWTTIdLmsvyxAE4xGEZld0T7fEwOkZ+Y69OdLT3/atp8zcVw6a9AzGyao
RqXTj/GJyoSERrOVyE97cqjomew+qb7drEWpm/9MucA67tjptSCK59SKrR0Hb9IVRLE/pB0XW3lp
4KvpK6ccYTaEAczURu5W/iPLdiz7F9mniQzehrA1tBCj9NjdhFR65+pW3BkdIe71sWJho1uWRwB2
LyShLm6e3IYMC7Bnrt6s6COhkzEj1iGbNeVmEBiqtUjzUKkm3sHn3eFFC+2lS2ioICD2SrUaM1On
5pJOfNTHPgPD0XhkjEyXIUtjVeYINCkrM4lZlFHXp1ecnEvomi/WnEPVKTBiVU+5B9ifY/aj63dY
qNS2vHqUgAoEJgTdNvKjAaVsyfPIGYgPI0j3cZOjNI0mVT+1GR6zEEvU5GcJg7OUZ1rJYbj+nDGj
+zdANn4EnYYeKsBuIR9CNFQ5DcaCWDb0ecLDa7pNC02ZOYP7zkayVV6s6qBIQzlJzmXTfGLJLPsU
r8Fj/HSzSfU5a3HHYIHskCLSSbvAN+b+siup4ZOo8rhtx25fXGfZUcRZsRqMt0sbMx86gvOnUVWc
/AIb/RgaPBR88EjTccRtvEPVxwBZkdz97+cbqL7dD2hk5zy++6V9q5KA8Tm8Yccxq/SktcaItc3i
xwHKuSE8tVUz5FGPOsC5gK4DWGsVJ32F0339931InSlk4K7mh0VwkoeG3m+gjop+YJFl6Q8ktZe7
dg5jfGZ6jl5CS7boafcMnZP3+KKIK3SU+bnOtYSUQtV3Qw6hgXCmozym7MiepT8TzV/KJFchottf
u6vbRGtukiGUafiOh9qvoaM+hJY3OcnOnjhpVXCKyqdwvm8rdz1Oo1F3mEWZGDvT1u0CzyEBYZKl
sT1DBH7EWp+FWHE+eSrgLqhtloCu/O7rL9r2tgdK0czq0tm6/7EPLcgaMRh2jUGuiW0S9I45tgF/
cLouyzvLbzKhzymC5BE4MdZE56yiCpUU27O44Fq9R5GrjWJCxQREEAtf9J2yiImymw81tK5kfJ69
z7XigdKEVcb5Myizqo0ul6meUrZk9Brcxvv1Qm3jjs1GVdwcDlegaWsMObm9QaBX2jUJD3lOQK5p
ks4IavF3szRr3VwqFcCSFdOGmdvhF+RDj+TpOr6vcfhbqqozWEDy6Z2hzxLcQL8T1IuKrapn+RNn
BpPZXftlhoTr2wFSz/SJiALpw+LMBkE8GQrmxk1bycMovLbakiBVdp2HpR5woX1nzgamGrrHh54I
YFa+zTg4zBt9m5IL0qDM2sHyZqh7z1jiHWSrM+RVS8Q6fct3ciSsZBm5tKcj+BqcHYMTz2fna1d2
6wA2VwqV9btCM9ZzQg2jJbb4S4NW/HgEEPEwHXkaa4t4cnep9k11jgX5FigEs7Obc1HVoIl+ZcUB
K/YnVLIGnjBqOauqeyDwodGNC0OZevjgTIRw8L3lRKn1Pc29dlrzK7KrtGIjwthaCJLTg2KAUp/y
ivT2gmRU4T9PnhyJKxPzG0i82bTxURAkOyo1B8ubqCjjMSgz28iuat24i0BVifK3uAxlpd5exgLW
tUnMd9bMhZOmK+LQ5WQjpx37xSB6E+Y24IRgcajK9VfupTQZiy8mrAxmyHsRHW/htcS/wyY1zwO+
fPHZ8OpLI9X6WrpzAsKLkWLHHE5y71csxNaH0UoVLYpbJcWfwWNfnyFgEL8LN/IjLgbGg8QWiqu2
+xTep4g/KWo2NA9Ff5DPKApC+mggturjOJsn1avZff/KLoaombJiW4qO0Ab4FcvBlYEh56ZDMV16
GpYFauyO6wfKmXhGf9rumnYfrJyhtAhRniCpRDeSndKovVOctQyyOLPk423HoyVxl9PACDeLHevO
K997EONRpTrRtHSSvzIU3AMglFCbG+YaUgpxVfcBnnzQxBg5rfWpIcQmVGyi5uiA1VmmH5zohDKk
1aaHoIoB+QC933b6JD3MCXVIXTESxghQbBi6G9jX842wHRlCpz1vr7Hwjfs38RX5rbAJKDXTvG5O
98mahyvNB/H1Y3BJfOJf97YoEZfd1I1opSufnQ3isV0o3NhoBAhWw2bVtvzVW9jSEPyaqiz/EmFh
ZDB8pw0R6nuCII+Foy1sbpp81g/h4Xir1NFNSUNlCV5evRD0jKBcmWBuv7LNO16f+5ivd9hyOkcb
0pupu/5q5hhN6EDuCmsghb7IKycUC4o44MezmBh3/j5elrlke12cYVmTv/datoPejN+ICvjCLMR4
9y86tM9YsADuA2tYf5B6yz6Y3PDGR0aqW299sHV92S+93ZeETF6ZqAqKqvx1b5rfoD8RDL6UDHQ9
d+XP0MROE5dcRSOPVuXz3kYQg4cs43AZ8YDGnGlG2M4je0+/UEh16Js5ZrR1IVSu4n/xfSR3t4c3
Rc7O8AtbYaIWAE/CXTNoHcaV8+shzJrtnvM4hpcKLa4fbibdZIT4QdwvD045iJrS4Bb7+09Ulo5O
4FIz0aeuLy4v6RxaLBf4HLhcvGQDtuBI6I8ND/1Kyoye6YUK0iCaiyskVEVin3Zj78lVg8SyzwnV
0VUHeK9oiJJWhBbdCSswHPoqM4E6TZ9sIqT+QLx5x/4jSjOBK0e72MYGqRCZAXUaI9QaJYOSBrJ1
ukqIp3T9J0iz77Q4IFf4sOG10M2p1bErj4E1dRxfUtYBZ1HdAoONLmPgVBh5suWMhkOTaFZh6JN1
2DdcDqR79c4U1xl6Fmlh8PLxbFT08v/QlsFg0+i+1RggfVQswzUnKBGpoeA/x4TdNQa/fct8DNVN
6RiDDC8t59qDwnfD+mmyAA0zl1tZr2mpBsUhFDTaz6WiJSzwCVWY6T+SzJ16qN/8fxsCfAodTGrG
V0NWmwvoWKc+c7uCJ2OWDe+MXXwKn7Scrk3oblsoyDmm/OwkglHcxY1gDeepzcGIITCXjhJAKVyg
WOyqkJfhXzry9Xy62ZJ/ctE591tRY9lMMBGm+nnbAVIjZZ1Ov63UH2C4htiPctE61LyHmIepj47l
mCjyv6ZaOpEOQEqhuW2Bi/i53K3h/4m9JvV7uMorvlgb1fNzwfTF1EdT3yUcRIQn4K1Jmw9t/+SR
IgbyzWGkf6kwAOtbxBiNlcOW42+wpy9u8Y657MH8uDdFvdcaJnVKt0MuQX9TDnM0JAYFrjuZTryN
RKNg6vvdE7dG1QQjJdivRGI7TVqRTC4zygexVU0ul907rBZqkJ//Djej73wyxSx9xz4BrCOgnXoW
uyDJWyy0PPNzLZlm+DKwii5vZH1ND8IlFdnAfCQoU2vdRKNkOTK/k2TgglHyo8S2uncq3NKh36b2
Wu/6BsEum1x5RDd8AeigpEtasxUIEXcwunf26bIlfxlFMSxFDhap2vul6Nb6U6vN3OppeKpkxD4s
F9VJznahNqyz7PTVcqmjKM0LfUEEmBgI/ZixEdl/sSx6SjQV47ary3UaycD3GYJE0zGVdwVH8ntv
6rQ4oXMs08s4/QXst9GgGpZsvQrbeH4yR1ZkTgYUXpXHlqWy6G8k+JNP/1HwSQZNN0NQt6hOM80p
YYc8oXkiAQKnKD32T8TjbpZgTdTKwLXDkyodZRgsmHaTXIx6Y9zF0sJD9l+u7vICq7VL5aVCLi84
h0Zbb9u9jEbbypP3aTs/5DqNY8NoFjuP1uZO60kPx5jPU7UB9OySaXRWyMbe0J02fGpH6cGd/flQ
xHJOz93TJFInxnQuecR8VqJpNgZlZKsHxClrvnH0FBLox66qkw46mS6WwmIM+cM4cqkeacVNVyKO
aRrRe4IjpwAbQECIm41EX3OUxT47AATA1wiFY0OHazCVVcx3Ys7dTxHGDDJStnhSWPU0+ib5zqFF
5UccWIZOZSATuyzlIdxEvjNlkdeIp5vJaU4sZzhEo+fMsNzTOOCLzHC2rX0qrVQQ8R46NroZLRDN
tJ1+5mniL6FWFM22N/GiskCXdRhXjIM2+jqpLPpty6inSaiWARMJZWd/ZouhgClq4G3AHWdxoTkk
BHRZWkrHTExpiywJIRL7Sk9mcFb/mttppbaafB4ZgdUrvMTQAtlCx9Zfrret3gevavTBzH/HVZpH
vhvD7ZsMQbKkS+DFckezN981VIMrt3gbGIYVHrfm817Wk/9W3dC4kzXGsK8X54W9QYJeawFBzrZ7
6xnZV7AZ0LUNLlrFYjrimIHuiRd09qXKgAeQuQRSa0aQzO7NFvwW6CpLV7AltAMimN6oG/z6aZ+D
wfT0/3iT3bEOy8z/G+K6eO64Cn6p413FKZ4D8icQyO2UY9ufo09LuDGSyVhXUjaWyemcBrQO6HxM
Nk3IuIdsyHAgIDCkj3PO/dN1WrgEjJ5cNtM5+Ei/ulhVfzBnen64uK2qYMTBYE7ZuIu5KP2+kQ8r
61D92yt09NGagwUG70C1qwzlJe+UIHSYv3/7GeLG+KdsBkOKAW9+XgyWP7hAZhSJKoDCY6vl7wHW
0cu6t/+xY+RIXr9EsMbWc5dlPtS3YOX5Jfxsb8fgIGmA5QHMJ++Dl85iqUnj/+YPIdNG9U6xYdZL
euasx9kOFQ+E4vIYphAqZNrez5ZVWVE7ev77Xh+ttDzTNyjckVUF4nOv2IiJN0vrIj8/oaQS5m/w
0Uz/idn1dDn8v1i3wz4noVxmWNbCBR9BIIuEYPxuGCZvx/a44R8eWtajJ3IteTTzzZRSig6hSMJo
ZfDruF+1IDKREhjn22N7skBpALSAeB5o+oaqsU3+Njwr4erc3QzF8PrRly4X4L/LMr031Gu+Gh4f
AGj8+5nMNv6m30adL9BsRNuuGjYVkAVqpqzyum1lAiOBgMqUej2uMcI3fw9Vt4qOXdGcxKnzauuK
qB+KSULmz9qcLE3acI9WRSJqxH4o7rQ85JTGMLVapdGzKZa3xdHxFFIQV5OMCo7gJwuFBssnfF0L
BTrWtem4wuC7VDcXEciXfo7tYrx5LAGlgMK7CMl5J52j5k7QWhlbKJqowCNX0e+NxAQO4NmLYOIk
506NnLi/60t/Mf3u2sjujjO+CTslzuGaRGZPiRLjGfuTo23+IG3JeXgPk7nVJmw/uu9ZDHQrWjdw
3yzQizHrt1G0uBuqVxYLRh+OMXid+gXh5oL/5B7phxK790jFWRKzMeVXT021N/ZMOHdyNe8IH20p
fMP3Xdkgqd2EoJZ16g9rmD4Yvq8pCmM/8egXT3zLoc+oq3OKLrYvzVYcqDnP8kyPrYBCXDb7+Lti
dbMCZJwmJd1XKU3VQXB1Zl632MnrA812qecJt5gyMjmQSIlFfTYHFVEIGooxD3MLkWebRA1/nHIs
HXojMMWrnfZooL16I8p+xPOfsa/aoY296Or4DalFxPA7wYmBdpWYkCbzgZVIEwndr1hR/iRS0jD6
KCIcxDgRkomKSCICaLA4OBL8umPckpKfDta4sSfsDD+DROn5Hl4Z5+eY8qBy13bC5FcJSR49yQ1Q
xsFItUX9Tw+b4/EQ0xM5RK69m2MI7YOlSx8UNYFMPeS/nBj+h6vJjvI18jq7S0fYs4RnJUdXhg/3
lsWBghVipzhNQvPVCXdcbJBZsIlD5WQjvun+MJdoS2rZSpXhzYXdEAqwfJ4pkOb6vhSRXsgN2hIs
YdElvB31UJHnJSyvwvWWVboGmChstwSe4P9CPomNCRSsMGNxQHbqhMRDQ0/EtylYRnzNM0yIqgRq
VxSD5iMWA/tUNe924a6CGHIj+YVa0wBLJ8h5TBPxPsv9rkS80T0Q/3IeTBmOyYPFgd3KpGWxqROM
xtLkYqo2Ou+nSvmL6j4HCQUqRM8x4lJcc/TTKJ0+405ez0Pul0vBn2ajsjQFc2AI5/rUqewY+k6r
tMa5eJxMpMrFlZjLhLOTThJV7GiDTMeMrR6G7fh72c/RSSxDHfx9g9Qo1Vs8onU5gxJ1vikaryEs
/TQYRzAdruU0Kw12Mxt6WdUR+9NBUuSCOIaU4V5zU+806iPo6zQ6MBeEf227t/k+GpVTwBTTjMwW
F1xSvvcC6qevIszOlegDEgbYAGsDv35+6NH/t0iMacxr3++wSciUHX4fCC1sjFNT6MKXh52dkc9D
BMhl6o9v4RERl9BFPD1O9PaYBQfFmiImBdEf76shsKFSwjKISGboXPHJyLIHYt3sCXmgeKkUB28s
GYUz8ZE9jkQv1TgLdKCxqNVgV88nlrzJQUBJphP/gxw7Lc3Wwy37FnS4FZjvy3gykdF4+fznC86j
WP5q3v+vAzZjUMq8/825l0XBTUVPFD3nChvhKrm5/JcHVRyD3CsTDh814K35uwO40lowwKnuBXVF
4fuYD1Iqhs0TsW12/dM8+M0tUI+mQFBX+9ipQMSYkFlHEc4Ee79cnbcY7wjc6IMObGtZXslvGIsH
zuocgK/2n92e0Hzw/zBZ1YpGVURJOY+9ZqTdT+HD6jbKUIIb/t6UGhRYQk1AsRqzRY5b/H+piBgu
WuuNQ2g70V60OAn4JkxvX+Bo7tq3Vl2Jp/tFJB/lKgsme8RbgP6NNWYGNN5OpoyhPE7jmDjdKzMN
wgJ77km8JerWuv4IsCfsRzhB8i90c8EhLq8yDqqbyXoCZiW7kbx+ReM1HCVbYMgdDM9CcauWEorG
BExOAZWE1iRCdK7wAngoUTzxrdEOlvJLlE4GqJfiqfCGGSciQayZyKlQ3czBvtti+GEqfS+Xnt2E
0/xQRhBo4TWrDarqmE/e/Io+MVVEONmY0/tmeTf/CcwMuFtEyFgsMY0C6lQBEKN2/wEGwB6vh3Ip
Cs7DIKzCljpq6GDlzazmWHn8TzyJP4aoJ8gE4Sv2FTW2kHlbq7BwRJ+6j3txw38hhdUiNEg8AHL3
ggJp97YdVs0uCcp5xM7X3oAS1XsUzaXJsH+FLnJtUretZhspCrYAhGTuHGu3xFfTdlEVC5GTUpLC
m4Whqr9+cM4WMs+qC1NZ4JfUTAF8gBTHavsJj8wIUwEMQUlQMeWIKNg4+LBpCkqHidLCwOXhFSI3
JdwKlsMIwaha2UVfK9f7n27ORIMlkyK85yov1X5KjaT867ych6hLj8m3BweoNC6oTL22DqjsDzCq
suCf9rsO8p2UB9z5qpXtmYtX86CiYW3iQRGPvTlH237eByHgd07SgOIrNxI65UhWZ0IM8f6GOP84
nZZAO6b5LCIDgHw9MO3xSVZkCvLhnOt3uNMSB7g0rkiJn1zONfB5JXyDRIAfEu7UgQKoziT6wCCv
XGQTRq6NjCF0d1twfdvZVH+uXEkJfNbrMDIGeNHO7E8ycRR/PmFWRPFT83kpcXfdSA91x6c1iyLd
5KuaAevc7CF9VkyTttFlvK0uXCnORyK84pJEzu+Eq6wh8GJly8iSrfEbqaT6Nr1nX74dL0noeIsT
k+Mrq0PluM2cZ+V9bp5t7AdQNsxrUsqOZk4HVKDaocLYPju8NGktNzTWFVN3iw0y9gayIE8lpZNO
k57zshtOBExvZ1l3Bg8PZoVm+eKj8dZ6QzYhaVMrbqpSkr27f5jeS+p8mkeCEVnMxnMtVBfDx84Y
fIwfpI89wJ4likVCOngCI7dyPnF3clLVSYJJlGsfkzE5tly/zUAy/E6mWBCn04G+rSY6nrsu0axz
gFePyKPnoHhaWYlPHHZKj8UobDKGZyN+C5ke6TP68Vp3oI4+AHKCGVR02Eo0id+LlTOyd83XDUgo
dJxeKb9rF3cy+CqSj1uvrwSr86fGhrdlblTT73whzF5NtMtfwPy9CvGbnQX9lsIYpuA8+kJESTB6
Suh2cCI8eyxwwT0MCUbj8bGs7r7nUFHEvg0jUHF6C7C9+OJYfEw6Bu7Y6cuNB/qiTzaW1HmJvvVL
jqpFO/ltwJ7QAPnUrHNayQq1PVL+mXngK1BXOwjna0rSX2sDIOBzGhCvAV/C686TSCQMaSLeaJOQ
2GK2acw2aev6j1ovr99jmBVab8+I0P+O7j/mmFMy8PsvIQfC652ba8SWMGSoWJ1O0LtzcRjii24z
ayktcA2xxW2Gngo4DFWF1u+JUAYwPD6z5ssF4av08xo7NSQvFrUTXSpvSW4Nq2oaoPno4tbmoY9+
9UQ8EDZJKYzVU45vNzyMJ4X2jcTn0HAYSFtFp0HUtOn7CmU7aHfGdU4vtw12DRCoMUU75PUx5pGF
5eXl+cWy4yU3fVwR4HaiNeio/Uh+8Qhbk8AuUsP8Vu/1UzrumOLKOBEnB4rgmjsoEGr3ohHNoXID
Rs/rjDHUzPto5MexI0Gstc7xNlDT19idExMDCC3sS942bu0spDMpVT+gMP2PLEAstWjHTnXhtFQV
I/xHkQjNfTCCoT6FL1T9gPPfxrfX97uNFNbTXcoutLYzipjeqig6p4BDIWagQsOqubeoU+pn70Ob
fF6Uyo5puIIocdUPfdbJN0z2LBOSBp+1/G55G7dwr+m7dXko0yBtxTf59jZjXEgDqKDVrkBRva2E
9bjcoAAOgRBgVDhqRQQV0WPuiCdy+GR+aMbGJT49JxpTrMkV9zkEeSBgvHSdcthf921VKBqrCz2C
h2GpVLtnun5PxezB5RoVRWGLkaijTkI0sjrzQGQeVibrDnia743GiptpBvzUVYWDfgyl0ghxRYcT
XKNju1PIJvnWlPj1QTQkt924AqgD1VsnEfyOzTts4u6/WE3Rfg1Kg55wkSzblMZ0E6auGvuHCZvd
MRbmeSEcvpvGLMRVN2QmkRDffgrzF/9tSrB6ZhJBdpEyVHoU/uTF/0pp/y4yWAMBGF2sefmrptee
Unqh1KAwEpZ8Y5ahPmisw9uaXF//WU9qNgn1UDNF4dVyuaWC0Ypix8/VCf+IvzOmKdBw8SPLE3Ym
TZ5y5Dl1z0SFc3X58zFKQ16HnE7Y9QX0Q97D/j5ihtq/s7sPWygrF9zatV1Dv3fncXOVXhxxvbDm
FbceGeBfw7V4HOjeP6PzJ3SxRv3wVehalX8FMCk+f1e+kiOQMF3gmPqB7GjfuftSR5+y1je+wPK2
41kkG4EZzeVGtauk6x07rhlAZdFYpRn+ACQdyOM/oUkwBFMN2jflXWVO3sxtcWER0Erc3K3A5lkq
EBSrZhFpJcN50YS5IwG3ggUrUJzTFWYiXEbvtH2bksQRtHOKQtKP2CxaIlVaBzhEumZbgqQA0kAe
iM5q2WkrqplPSrezf/91JdvMfs4etd1pDz4fkbOvfOuqfur4iCWH9FCyPPi5qWwMIOWf65WpYej5
YUrLJJPPpedUEKFDt22zQ50k6QPOWibzB5zajK2cSvzEAx5VJNfnqyxcVDNbx3g3K0FBDTKsflu+
Nkyn6OKnmdfTcIwxOne7ZxhkcTT42hbsDj9cSYKEd+ekZdZ36CbrjlHyQ80yPL0M51ndS8gMD2ne
cOmKMlDUq6/7vOpTuTCTrufDd8A4ij0FTMH4sRlMHw8nmC0bua17A7GJ3kdQCIZVKmSfcOY0s0xv
LNBDgnFCcim/utnwsTRxH0A5tClzPDzUswZFWun43ElFaBPOiAgLHWn49T5CaajjbJDwXXifgQVz
9LyE/yTiMvdokCKIO8lEjljaUgoAC9AJ5IPiKMBEZ+Ibm+9merCjy8BvDmHVyi0/zsGb7+YU4C4P
xFPKE4ITm8ytpitAGb7bpeC57ord/5zYI6GV77+YsQ6miRu9jbxejzp3RYL1I+xtWqTigQN0KKez
kCwosYoL/sGVhmP/Km//viGg3b2u8WQemkr6r3LYJwazEIU56CyeDURl3lDEzbT7qe6zICnC/8GI
npvSX15WlZllaHt6YHdGT4VJmGPWCkXekfRIE3WRU/q0QwbCZ0FDG3MZyIMn6tb+VM5L4cYkk+Bi
YcHPYRXEgNcos7UfplP1BBGeMf0BjXE9jIyr2WpGQ1imlIAWLUn8zENao5vOZ0qw06ezlZzWP9YJ
lZTyPT4OjEiZrAUGABY4ZZbhA+r5SFHFwpRBhD7MDb7RTTosHBPqGRv5SL2lTKWCWtBmImzRV58G
svbIw6OjqL3aUf0bhCJQFoV9UnlRDkjosqq4GoDLSNV+o2PAW5gQvZugeUdddaMOAmgPsTPFt/Kr
Q5fF/3EziNFm2R4szOBkCy8Hm2o+eQpeVzQT0HNQYIed0YKgi/oa2Zx4r4ZXOfG7tyMnq0jSb1pd
56pTIMpOfBBkm/6/EoD39S8SYwOuf/eSZBjzzUW8C9Duf5GWacjHOrwz4vErbudzW6EXpkCOIWZ5
cPTIPuQ9b/C1PB/7DcmBfK/BpGIe1KhvO0wIFvTq9+mNkbuFVjinbuMdfUkPziOf6SjdKsiUO2D7
l9A0w0auiYhIo4SnfMOYEGsXcrjERys5XtpB+F1IkIkwCcAAHhjVWj68hH/J9JggW3bJ6WejnBuE
GL3avg5xCPofN512TkZ5OYcssEQ9lE+M/s2rOpQMrvadXk5njDCM8GDuQs7ioEAgqiKv+kT3L0mK
jKFa8Zw3qvocVqkipRFkR7suyZmPpjUDddb4Eilm8oo9tMw5x5ZNqmdT6u5uNxVxll2OacZ3iXCd
8DoBBFOZ8d/3S8L655SbVDCKo0lcshuXCu31z4TbPxPz6FoPQd1XVDuNMi2p3HiqBfJ8sMZ5/dG+
4uCNB5d9ReHv5ZhF/eqWevVJMfsmZwk+IZK3NHMZlnBXMtWhr3v4xvctLTqnfveQ8zwkRXI+W2z0
dUf5n1ncEBnUN/QICTVUj/0cBQl4M1hqTerWBUSm6fxB39GlKHgFPvk8vTpfTPrW0msU+k6KaL5X
/K32R3UngTKyJhdMz0qvFhvRGvWsm7NMWuIrvPyCvrji6V6IRTkqYCcA+EasqMcf1DX5kDNddlrY
oDfvW818ePS3V0eQRHqkh+bazecuDPfADhuwQGPkna9KPdLQpxcNENS3CZA0K3iFxjD7TIMb+J7e
70fwBf/WInXNvYRgBXP6Ib2JOcmmTb86i00fToK95YzoUuBwwgCsforsxEVU4zosFuRbGe44m3/L
woKZEAX+VS8rrwSCG5d1HnJBHJ7tSnigm4jJwLqx2LQHLCRxJQtlQaS9WGFuiV6OuTYUhXXEd5yH
NjnoYtBNjivXIM+l2DXCZ22S8rD23+B0XhbqAr/YyMNb6+qsFMn5MBHYNTBP2tfnmFSUq6Ncm6wM
a2nq4fBg/1+9vTvpkfWVu7OCqOUjaePYLu564sktTk7+9vMjVLJarQwZvhj8Dobb/l0AOHBc3U1s
2tg6Ns3K/iBKIS0Vm/nP6OcFanILVAQi9R3m5FPK1f0e3/59FOlT/2OSW0eFEwNj252jpLSGp+8n
CmOsKgtDwXQx5lmv/k6VpA+ydjYn7MoPuFlWHExFsvXAiesoYYq6ZEPsFdgnjp0aI2SKHn5Eu3UP
XsKpwIeDmCgt+QL0kZu4U9uha4r9EmpIMC+iBfy/KGffZo2vVCrRZwxav1qw+7xMl1xmFggKJA5G
b+eBS8l4RVPdiLUlZ5xVzWvO/OPO0S0iknDZG2bw1TdxrjZ/4wLXE5uCOAkGzNaN3F4vOeEZXfD8
dLchAdMhJaYMQNrI72mNd4ORY9AqznDHRvnDJDSKxqHt68qbrJGfNweUjMPEPwynYIDXc+lboz7u
ksq694qOMAHHTWecCNpJfi966LbTvNns4KITLEeDZz9g70VEnCm1P50xblKLCL+1HHWMLIdqyQhE
vDNYQtVp2xwVtje+/i5yfbAjbEbQa1Ucy2LdBOtdareva7pvgeX4WvCFfZrrufRixONzMUvGd9Vc
hiSaa/jJv4eqBVoSG2ZMvur6VvqcWvKls0Odd6jXfT7qoPoENn4rkC91hYWz89/wMF69Ghu3GOyz
9neKkyutUv9+Lj7JjtFYd8q8zfSY3b0Sg8+j/5mSpx/XGmnJiJw+QgOv/5I3OIM6E+aMm+H6U/W9
NH0VsjCqVhXk+mMxzvGnfs4Rn+PiiI5e6K8BIXWZoGI85rk5IejUojg3JejXpWjStrBQB8UPMoPY
8pW1nIXy4qhp+7ZQGOFzH247CofXqJYDQykOCWVXLnqilByyon0sujbhgmFywwgUOD0Qy46q3TOk
aFJWW26CVRfRo/OZxnwD54Y//CP8BsAEaGb88+NRRWO2r5HErTLS6kfDUl1ML06DYPCq9iQvir+p
iQ2qIe+4nzGodUkSJEfAWmJo1WxoilZR7cCjXB+yN8582SV0ED0qsB86YIpem8k5BkRV10hOJUBL
enLI7qGR3ggvHGMwrnlP7e+JVfVuCtRpaQbLOIQZCiB07dcvN4LzRnky8UUGceY4DcfY8ugQPT5r
Gh6Oj3h/nWurvg7B8Gqmj/hbuSfv1tp7JMiraYcG9GhjGCR4Hmbh1dUQBRxBeKF/dUA1A/6QM9T7
8wfRzSHuRAXUCpflyvz1ovzKFeS+L4XeFpYuhBuwvk5l0dZkRfmVLnP6UkaROU0czGraWzklKKwS
vQPRHBdub5ksoFto3uOGGSKgkiQL1mcEPxORFMi3vlcEllHQxM+oUCZahov/8BSLZ5fzAZJ1q7qA
yLBGCgLDSDaSzTOxs0ZIe4Vdj7aF1BNkE4kt7PNX50nEeTiSQGBp7qqN1a8EOOyXNNQgvwYSt0DD
b1pBgcXLjG+u0hvB/5T1mRiMU5gkmBMMNBKCB53CBb0s5BYC5zzJ3o5g36h/rsjZr4YZdesMrpG1
T9c66qzGE6GqFt9g6BrGKB5Wg/T2anYnXt5WS6ewfmse1sh3rtJhDS2BYb16O2uFmJHb5mHbkjW/
zofHWpykdnRu/kiIh+xZWttlNh4eYeQzv6otzVDLgr8o4LR/88/CC+GTI6AJW06cT1jeX36mEJwR
hkMYeC31r5fvhX1Bt6SaoAVfUcqHeJDwkNh/PLLQG15PE5P2X0de0lHvVot53zhsg9nnFtvWn3J3
7ZjsKFuxKajykFFclXESCpyJwcYxRRQQMBCdknThlp2I/Uurx3tF+CV0NdAQrOybOg2eTxAbOTKK
QURlE6dHTxuKu08cGfki1hdrSNobBH6wpPxeFbUudoXJgptqGvlOosLrXVxHAQnl7RuoXAnVdAzj
YJMAdpSQeOfm6eTG1Jjj4gj8CBdr66XsvtdlYvOzKviDNfLoeVdq02/ZUgOcRC5OKL2EhmKfOfz/
EZpGO58u0rLoK/nNIleipg9AtN5TYnmuQ9UpxGfoCWcFDYXRAddlUOt91KqPSGXdXG+mFv1DRe9K
Umavf/KCtQCoIUL9vW+zWFLlIu3RJ6oImbDJjNbKp525AO6bIGtap887bxQFFPhtCy+xbUZ3RYbR
k1IOoAAMZJXpeRMI6gRWrVBEGdXX8PB/XE3Lw+q8wcIGdWIp3+W47y91ApR8/+jM2XDYic5zAeGj
R3sqUmLxhwQf35T5eTCwRAeI80Ic
`protect end_protected
