-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AG8fTuUiKS6iXOlSRysRveH67W40mx0m/Cjx9ITFU5uCFGOzwuFno933Kxiwor5kRXeHPls/lY/L
iYJEVJFT28f236yvOYrn3XlQq/q5e7iWfGagFW16tDnSJpL/wzmF89PTxZx6Sxbnk6OkNDk0dhBL
6HWuhdd2BvOfs97FnHeQTXSTkgR1iiZoZPl+ONsyHuQnw+4QNpqbIOgNYqZoF/ItwB0P5fqeXzKR
L9Rn0O3Uwds8umgd/kRon+A643nxcj0SpFoB9iKvjLFaV55ydcLwbQcxZPY1hSht8kyrunIALIQ9
1i/0rvqSbZBGQ9J/qnnRJHlN4ki76sh2wZFtjA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
F1j/ENNoIluamb+vHHMgRJ/d6rGENkYyh2QuFyvgwZlu/ZmuUE+ZpFf+X+arQRRgMVpWiI7IuBrz
gSuruaLfDwSjXM9a01C0mGZCLZqeaZqYAqDwrFlyhfu/d92B+YYXGK0mLexgUHoeBioZIeY7lFyY
wxLWvyAKluy0xnzTdQyCJxDKCSYyoBCTfRxlbW5YMSZwGazY3uCLcpMNzeHB3GCJuqWGvV+uyrCH
0a/3iBRCzVtX9UmfzbqBdU+ARh6VGYjhH3tx9Il/jYwfT49Yh1jWc6+YZF54MqV93aIJkBWEoilq
nYMQpmUJjjvhU1fT1ACS3JmWP7B6mthsY3g3klCYO8vhin58CSacM4Sp95NT1NJvVQn32PJFWbgE
G7dn7srPdHWP0j5iUrNEUX/FhWLSBHzmz2uTBTPljTt6TgKSlRJHQsUxbPIEzWiJSGWhOHbdO9V6
7uOi2KVWBHFSNVsO2f/VMKKQrGIBECO/3fHEevXLrh858ckJFS3Cq3KnhcA60OM2ohZ0sVWo2zbT
rS7BERcz+c68g+OkEC6SVFEPuiHZJ+AJmds4enbP1FPWpugHTNfL9f7oOEl2DwNINWdTEn+0xawR
Xk9ssEn1Eu/QvGIZHD1fhXC2usKkOGo+AjN67lrnDi7BknJ8/YwrEuCoZh+xjhDD7H7zscxAO6uT
S7Hkz3/8ySixPsqzZtNd6mLbRMHoqS030gDygOp8kIzRR0p/QAfbukaqUtIK3BPmb+rRn3tKyFIA
eZArFIrkRldVrK6s7v/cLgpw9FGaDuXsv1UQSjK2FQhRlubSm7aDHL/i7sTTVG1kXJ4cbE1TKCM9
bA+veYOQ6wkxRQt5X8jq+igfVkFcdgJcCuqJ/HAT+j9Tcf9VT+6HscGtUYHC6w/nYJQY0caXouZg
Pilp+yYSGeC5oNJmgSHN/d3cEORyuvsKlu87upVwXXhdifasfDkEpjt/JpRsMRXV+bGcvzZq0ukJ
9kHRwC4/r7NjFCefPREfuLxWDtDmCWOVPOznQ8LnXXGPmLlRSH9uy5cl+JM3TnV2O+59WOx25/KY
rDDFfQ7x1C/Quo4GINYimPWYeQiownfpx1If5CvdoPO7Fq+B6cJi40ZVLjGYv56ypRk4Sy88SKtw
MFF2eHMHsLv0mXsZN3UsWahvR8fOA4IdOrDtfWWQytlKhDGbyONzSESP60loh2ojDbzbH9s+hvJ1
j5nB5RRykwd3auxNe3lSAfDfE65P9BK8TmbNCuYR/hUzh+J7RH8vFeoRO6N8OyMpUxSu5X0l2toD
J0/LrnxnmCfxknD6TO9+o6V3EOZk9PL7vGq3F+H+4XMhM8Zr0JccreVUJB4GF5Ysn2KhdkEKyXrH
zr22wsb8T+MM0jVT2R+4/SUchMP9MFmP/c50Dn9ZoeJLa4PBNbifGLQdE76l9MjMcCXBM20+uy2O
MMLLL2Zqs4AMVasBnq+iqdEA+D/ewef9RyjpT6F1/OJ9aJqP5mzMS/oPw6LANNkZWZhsMy9uKh8R
2axEk1oSO3OmvCeh+hLNWAyjlrrLLk3OcDChDnBfqzatyEHodsokWlK13gTxo+qjsA630sRR/e2F
4NLQxNAtACplPOeRTEnoIl8ZhdHw983DyN//5YuMQVZMK8yS78YPdrFY/yLPEGbOK9f7S0R80ggp
XWp8XEuphquLT0X0b9Syw2naAqWFgc6Inu0Lh/urZoznfWks6Oz64hmm61LlND109bvG/zLytIAF
5xneCKjKP5BXoBrJhmvcwHx9yqz1lobHSsxGa5DNgnCtZHsOCJUfpA8i59/ynnRg0QEz0Ka8RKo3
/12glhZa2XPGIK6ZM2QaqZL87TUgMmK9vBLZ7e0bG73JNe39gbuEuirUT5GoXCp23CUwclGGjwhH
O5dpCm049Hs5vDNpmAg05blGRpa3ZGOhFhbDkGjy+mwGX3DBPO9v6n9a08H0B1zI6L/rydqYqD8k
ealvGXe65KkvnS+pRuXTN/TxpPia7twpokCWqZDDPT04zWeI8H14aSTi1Skq78XyKHCcsUQh8O7r
AYYrmhhkaMfJT44U33WYFWQXIv8Ih70FBel/hy1+6The43wCQlKy7RP6HtS22xdfePz6tt87U9Pg
ZHopWsnaa/g6OAYxQ0XmYgsq+vGshyXIXZrvVHmzqfbNOqOz1YwwwpMLoNIHbBm8NG4RP4Qh28GB
YHZU46W/naf3w9TYAOo9h98mevw/m01b6EL7kFifkw+rcavR+0ARunnBpuqFnuIjotUdJMDSD55x
buV9jUq5m8CZTWuiERduCYd7eebqkq8ve3W2tlMycTF3sgD2KmLy7ssr3Fq2Ttt91HIswtMwQB7N
ownMLfuXWbsCaYI1YTF0OvjkC/kVmUDXk6bmDWraD1DGpw8GpDvQXXpZZWiVmXe6B8LohmGRTV3r
1W3cC4R7R9gTT1580sn24/LrbPWvOmk0O7au+4vbOPvwtMge0/Y19oFqPYScfsCr7l9WVPC8hZ5y
IxQB6lJXR+UXw6FGsXnAWLY+WCIbhHwwkpAsNtzj1Vz4F5Ml34+sO/9L/zpYpXCQRXuS74z9xOvg
e1/GJ+JCO/VbNAOS+db6ocD0PlDFQ/mc8QW4BLblob9/vSeBh/LEHqj14maF5ltmod2Dd8J1PCre
F5BeS+ByXnFbdxcxy/icc7UMTAYkfi65epBmsKX2F4jb21MGgr7tFguKOGQzZeTb07O2Ih6u5dbn
df+hpZMW+Kvls+uKtsez0Ny3IRsZjMLopTC88YICEYNO9+U/36wVl4zR4h/RTUYrTdhVhwE4oLGC
LW9LdgXxayCmo4/rfcnVFs1GO7JNPVCB08ti4Y5BbGB/XHD9V3ye7MTGZuvzTmCjmfbaHtTah4uc
IEfE66fcahE3GddbH5K4OakflzAPJL8gZ3aUd6ufqKj/9euhSUvQkQ45b5PpikCAGw+Ay4VaV+Zb
P1xqlBZ8b45avDw/7lZysuscmzWyzEKc4EH7A3l8fsri8taJRvydQVCRciky1LEn8btYlkL1v6eg
Cn2DzdQFoa1+7rqCZjNK51CvluZqB7+eMx+lIRm9U4FeehmnAl0on4dJKa986xmk0nzcliJaxG26
UCUqclkrW289VbvYAFwK4DPQpKFOk8RC85NCOo5dpv7Rlzr8Gu8e7+Fsv1MwG4NDtJXoh38Xiib8
8k1KP8iMAg9wFa97tTbYb+XaDTitz0pHicv8XcZ2MCoqzV7/K3s8DmYY5siQ8UCeyQCRW0S+zgxN
3RUUjQ1iTN4Z0WTVC17WDp/mxU6jzMi+IxZWPhUW8T/bHLSR/PKnyNunNWGvqR3AJGI9kOZAKqeP
UW+HfNEcXELUTJ1tyCfKYeHZxS7TXKX1dQpE+lsx/OXhABTQgg0dqILysq2C0FGzZHCnBwLWdn5R
0JQw89Rq0UX74DBW+EmBz6y5NB+3JzXSk5cigDdBNvIV0/cAkPSXunURmpHgfY1LvT7GcUDsmSPz
iS/dhpraLYe8Nez5fFEJ2/OMeudS4+XiGHTnaK/BPslpZC6QhBfTFSnjU9Fh6zlPEBUc2gq6fH1V
Kb6sj6WEYoadqcaOHITOwmblfyXVdN5t9NKnXiOBzkzmLfG0qhjHkaI3JXeXfwyDLGgA+4eeIV8x
FVx7KHAi9H7OcFEaDEn//hZqNA0athmxMIi0nvrLl2dbKKTpXzWQi9BaBIWn2wzzZpkuOPlZmmB7
nVfJuJeoYEK9TA0iFfLYwyiZD3rs2AtEjwecFvsvY3GI1aXeFqPBFMDIklLhMJCRo14ZhXA38Tyy
cw/09Oh9JfigIG/fpTick9PnLDWXmPSLZNr/L5BsanxaQGWfgYfVu+B0EqH1CHcQRkbkhvhl/1+q
j9Y6vBwQ2H8LZAsBnJfz00JMSkHi0J1J0XK/ADLaisk6kF430TTKHq0ltd/oi5ID/DuMMBWIC9WS
TgpPsT5P7qe4gbAvBT2WT5EM5IFJ3NtgXJ8itBRzPEYDj3Vqv9DSUO1XccAd/pDaYOKEvzapXifR
OVsPc6UvET2sTRAptJO0Q1ZaNnqOCR0Pgf2F2Oag5i0z+RSNgJq+C+IEjibZDoFiUQq8PxQb6yxR
u2hnvv4FJWuoO0QbiMbeOQ0exIr27PcTuqnPqdl2zGseAAizIbzDZVcfiXZnbalfCYITuogtFxvn
ZMEOygepxae930DzjCS/oqJougNGZ0v36b0zA3r+Y8eCnvOPAVwzZAHQDcItv+OYNMVnYW5J7GqT
tekV4Frp0JnQi3J/Z+WE6PhAhF5F8L6iDg+rNHWAP+OKIPcZ4FKLXT49HTmb166+uewzykw26e3L
f8mkJZdcN313X08D1te67j1sXNkuObzMVd+cd4/4fyGm8vZNJSeI/AHZzM0v5rXAkxs64F6FhV1p
O9Penj/HnwbB+rT9ROvDQzGNz1FpO5hAjVYbVZufeDjb7ASo2r+FwpiUXQK6Av89ooYy/3U5yKsi
+T/UlI0H77EyZ0GJ5QgOwAyPGjXt311VCWBR2gJwcdVpSNryGV4OqJsdxrvHGKaLlJ94iMchhUU6
DhfZmNTeL5Xix1bA+9owD42oBmrYHiju7uzYdIMnEhqmmvaiufwLUV82CcQibnpxNUouHhpnNiPY
9lbJfZhxi7cQCA67rBAJcJSLRSxxpeZmcndNCJH7Kk0uTDG+DTUxR7fZAzUHS46RoFy+2IToGchl
x9Mna277xBErp1Th+idHRlF2SWO3TqEyGUiWrjTRdB9kidr3lYa4JPoVf+WLK34lKHouXUfny2De
f4fMF5y9s+9GlVkP9o8f/WgZl2+Zb2BzT5yjWl+N9/w8tWgKa/JHVk6EZjv7rBholyKf4S+JpuG2
7/nu4ZoCdVtyYi/RidbbscL3bPmW8r1HHCCLzarwN+q5KgjD+uy9V6trhd6olfyK38e3kLRKrAAp
Ylnc8T2AloSeRzUBe9XRRDbWHPwQmga4pDR4macRZ4ZX8LUA6bbhxDWp6UCNDOZxXyP5JMcfu0mr
i/zrVbpm5rctAde71W2kJU7A+FbiaRU3quJLtBSmQnBBScV9gylwePGwh2IP+sup5WqJW17eO1Em
BeVY5WXLxFgXRpR6W3Tv8Sv8vdSzzhUvmr908tAo69xTeP5+4pfPw5IFH1pfhUcvfiBcmeKsiGVf
+P1Wruk44lyQlKrhF39nTaip4sDEj0p0DckI6GT0ejkdU6cM4XXWU6kIUMDfWNt/kHL003qKzAa6
Eixgep/t8qvQEtQN1oTNtR/1jz7gzYsK1mkDcNzToTkqQCXPwPHtctOfPylbjK1SVhbe2DW9FFal
Mqo4uVFO83INRZ3/4ccIdI5XsIiw6FxzZKz5O/d3Vp4FEW2+IqODo3dPdnnQsbh2GSuTrWRv9kKO
4L6iUO4crGdjBmhYfxvkg6Qe79mTAwCqsmI4Jw2h5LV4mnbDCVAWQekhT89JoDOyFtwRKVvXx0FS
AjrY6F5oT2ZjC8FdAQtwor4mbEkfUDSz4WnNGkJYi5qXJhQmcDGyrZvjWo7aOGYCOjsaOKXTrdgv
mCtrS4ymLnNAg1D4JaRpSfNikkzrOrICvjVvX+QHnXpND7yuK08OoZAs5vMNwrcb56rM3jxa5yGM
BlO5w0ZeJEkwx5jthVgY5eWIPVg1g/wlOcu9gi6DIZlaAnqDq+gZNQgtKDa2QodI3cuqafkxidQ0
5frQ2QQzguvi6gtFiqeLxHm6eSxLQEjl43hGn+aIXguMpK9lhOrkhiwYeCVY5RtoPGiHNw71k2KE
dUGJfRCtQhFhuTFoDWlxJGuo/UIGrW2VC3rG2184Be+lhbqHu6Tb4g5Shb2pBWL0c6xuUoy5xc1c
fK37HjKHWCBu0hA+0rZq/ZIX1YIB/ofrLlORqCazfbBCxmr5JQM5aiybyzUYEKakngPUm0iWn4Pc
2fw3CVt/n3ljhxZYkV6R65uVHb6Ryu/jXlAGuJzAoNxKpPugeOfZgLsYnf1pS4vcoBvHECzn8XKo
hR+N8Gt8vQciG7/BFxZcD/0yU7JBttWe+m7YzpZ7rwrcy3oqI77c3MAbYUxuCxjY7YCfg5V6i4Xx
RszrUx/IAkVH/SbiU881vasynXeRj3MMvyQbuiAkynMOnwL+0i/yYi6Et6s0K2bHqRikkbY+SjMO
VzIu3rdddkah4hLAPSrzAZwxDLsSoqn7jIPY7Jd3lvdPiyfY49C2GQ8zYtAQWhB7+bKYVAHugZkO
E6HaSEryRSsCHhu6N5XB4l8WABHQ73rDhJpBWRHb4e74mSA97JfokvEJe2pGSPxjFKS+nAQZyMUt
RuVArcyu/Kles3gvHO7FjuzALXGpso7w2oJfGBtEUrIIsg/SG+tym+6YiJYyRpcE3Q5Dlx5dfX0N
bAs87LVCj318AQN2uhNskR4DbNW6Ht65QE7IXrG7/Ldvb2yePjlCFomX9CC9QwdjqlRCJiPKSpuw
1uU7gacQgqxs/mYyy1LnkvfBIAFoRiewdxBynAnEeitIsnU+4ZlsWEEbFQeKDrxDp1iJBMrQRxBF
Kj8AAdIi5TRv1avDgKKKXr0NXP3rU5R/IRi3KbQLoRk7rAujVwtENbEHDIsQGz9N1rk5H/Wc1te/
VBvaFJLjn180vf0avDb9y7Em+90avd0t0TLM8UWLvIHI4S88MDxS1hp7xzbocUCUx/5Gtgn5jrco
Mg8j4ZsTqORwkMzOuRZX0dROKE6wjNXRaPNXCpdoT35Vbi8vx0DUzSmov5EGwtpNbyld3d76lCBX
WwzeDXdamzUw/PC32o+BQQrE9TR2fz6VGPyiadgHGRxGRbJiooejbjfs+9XZ+lK3fWImlAAII3fX
ioXw8mWdemAWhrBxSzWHSxl1VSwmcxLmr4W4g5f/A8hV/cJkL5V3CEhwcKWDM4pyynXaY5ff6V5Q
R04rI2t/xXlU7ypsugRkIERPLCEvDkraI29we/3qMGC0+01PdtKjXXAuyukOMWsRO5KX1Ilvf1O8
474j8kdkL6SVc+2C3vhruCCPBr9KxpkRk62kBAiCVINLyjUmz/ew4Gf0zO4XeTi1bbqxvHoVvYbV
uJWyNybSsfV8bdAgnCLjI2ulWbxUGkwBoUuVk1UOpM3Xo7BvPWeRBfyR4n1C3TnmMMYpenNG8t3j
gYcjvi+dHJROBiX6rvcVK4ta8WvXOpAMubBzWA+NaXKNDydQU5ZHFCg6+cjr7BnV2fKrlVU7DtHU
M7C37RY4YSeHDcIhzDQfmWhPyd/tHiAwQz7pN5lE+xd+wFkfgieW3ZaTGpxWKvsa0NwUrXP43fIH
/bQSdyqrOyXHyhxI4s4iZdFUcoq+FFHnGTm+74Nuc1aMN3vJhGN3lNq3XNRf/VFmyfSWzIMX2IUR
TnQAG8m6ietfA0sY/wmVq4qFVu81lKYB/EEQGICLYJDoGt5uPk/YYrTu/kgRZw3jEsjmh6GpIH4Y
LH6r3tiE1G9x2fffuOrRn2GJYbQZHiejWFswvnib6rw6HjWLqS/aYGjSrK0U2AT025+50AdzQrlp
QUb0mt251uS52+p9wJOhPa4b/APdXBgFsIporBRvnJZQkiI3jWRj9kSpLmlj/CzjQ7ssKufhDntI
XYWe8S1c/zrk+acdFhlTnmFP5SUvuSizNS3wYZtWgMMpHF/bqOmAGwW/7iajZjb4M9lKJ88PAv7c
gfByjcwwrsDCG5rHx1Uuu1dWySZKfThA7lYhEy//Qhb9MDstVQzqKY/3cytUdpeIlwoRqGSNiB/l
v10NWmAgIvWuNhZJc9wjga4wHFSTTkftg04fNdzJPuDpn0Sccc+M0s7bIZJivQh4GJKvl7JKGwM1
j8PP/37S9h0J9qbtia5Bnvg/1Zq/xEK2NMd8KTtP8AUdiLXzo7nRL8RI1jOhRjbeiNkWY34FHHjh
MB5Xww2FcycsnBmeFC4ISPF/V3Autv+Fs05CzMOZid9EWk4ZCt0wF9W18yvfbz1hE/V0s+NvX33c
drSfSN49ryzfGfAy1Nj+SSWsh1WfLA1/zV4EOn6wDeRWB3a6vNiM2esx1LXFBEVBckoOvj8aYt5l
nrifDtz2Rdh8TkIskWzhDbmtj6Q7WT3xoqYR4Rw+8OQvc3rllyLxLaw0TUBVizsgKASZjDJc9odA
GoPSpLHgbgqaJkpm39plojSgHBJeXmj3YJMfMRR8Km5YIVSRT4X+cI2VTl56iHFMjbUJEu3LtpyJ
bLIIMvUt5E36XT1z4hxGy1CzPorszHXY8JRjoNnrlpS/SVTtgOLJPCAGKrCG8kvJkJ8/UrwB+pJ2
7T6FxvN8m25YA0QtQwW4dR8gGL+9POtNMsenM4i5Mp3M2bTBhf1fqndSYrZo2+TVItJN0Jdkcp4S
FYcJ045GyP3rmaTzJrNrDwVEfU11oxKFiTy+sc2vLPL7BFhZLg7e5IcVO7ZZ23RzeAEjvUYIkkRn
X5y1LynhWy5znuj0mTGIl2dSrLgPLDfipbrowL8Hy5v9IDglU95Q1MV2uSmq8RtrZBXtrn5JcfTH
xqxz/IY+ersStdAuuSAZWG1+y6J7tDqENpTieVMLBUmCibxx/pe+KZEGyiOkSpiTKF1IP9PhvqiM
b2CbsFUS2eB1T4xDO/kNzX83DzBB/wRciXTqKljpUbdHd1Gq0kJGIYtFWxivgjKpGACb+kzO7o/T
7Kucpa8+hO/rDveXQD1oZXiAuXr09dHMGXV4EdRtrhUjMI3go2qoH2ksBXBqXuWuRhq+Ff0Ix1ES
r+reuW8mNk74w0BSoF0B9b9CiqR4pZyFQs4jMbDiKNjbfbDpTa/zedbyOLxNvPip34Rvq868ESo9
dmSWBW9briCMIInDpm0wciPkhLlZRZA6o0D4+tn9AYPTlnkwPbmr7RRVyJqSB9Gr7R6lBVOrwL5y
R1Er6zCPzjASw5dxUqKuVqyUrdcoyTtw0+NEPLJoLxe5741mEDrgT3jRE/jHaGmw/VPEXgJvqtZu
K/3gqnOSArdNxK/A2NY0fnzBLahOKQ99m0xZs4BIlmtrcC9G/QExMqnslNpKZYQRMWGvO5OciDZ7
hob36pdSY0gUxaLMJDwa9Ltn4kM44aeKZ6RbyyU33Ed1dXvbRMUTIDNQHpDbFEb4EqIh3+C6W1dq
3HJJLP8mR6EsKaoXTrhQayDNCRaYja9Y2ngLKKhglsEX1yYPTN3OOrAheXiH1K7SFFQClTNL6pfi
Nt3LGaoghjZCwdxk1NFHlRdSxbVtLfn330lFHFPah8WmjRSh0NKHsvugXEfPE5/hfASSPWULlpUj
cHiZaa/olNFwBKsSudO2py3gjunKyTDLdQg9KjnNeZJtXu+ZmY+Dao02Vz23OoS4oqYWsfVrJ/jP
zTxhgRWtuF0j+IIsJBDf+RKxrHik8ei83+pFAd0w4WM63Avia87tZVbIE9v6t6eO/dLVi41sVGXn
FiGiK9/YK0jXkgExIv8jPS++u6AyfNu7ZKJOXAth4dgXK+q/Mweu2myjw09UVBm8P4Euh43GEVp7
pM/+soQBtm3EBhd8dABmH0QziE1y2D9z8Eu5HI/kWCAdMoutDK3sLHwwH52KizuLrnq/MoJIsiu+
WP0Ma0qXhVupgc4j8VuMrUUCiUa5ZwSALw5ThlgKPJQmUTFMfNcM2NDVLDgKlYwCU02o0jXY4Qux
MKW8duNECKPM0zoeuhTqgEY6PKFNcBMoDPbZfKZaZy9Onm9/ZVc0Id2VgmX+jAuNDYx+wD6NJ3v/
v35xr7Jy/Pb5gpt9badH5mzSKP0A5q/s2xciPHqF3bcS3S7TyPGDLMYtFdqx9V5x9Di/Bx1Gfle7
EPDQNqBVimwCIvFPybr2nq7SKPSqI0vHkyQaFiNvqGqThj0xXHVvVT1cM9DE19IbI0/W6aW+gRNy
cVOyrPhp2H1VYFAWEltR4t6u8KhK9CdDNPvelQFdWTWtcRfgDrAr5QHM8uuTicoHzb2/giDMD3TR
OmLUywJQ28oHEg8F19nR/ttyG3B8FBmVgra2DAV8qX+64Os79tRo7VFMxJMLZr1oKQQPqveXR14M
bqF/Kr/FMMSFrIY5DbUUhYjko7Ptt+EJsh3almkE+fbiDMIRZHjH/fMRq6DpkL4CJyMOin0UDZC+
RSTr0befs82xNFbaZAVaj45d6Ieykib/Cil6GPWCe/5aONPyHilIGkr1BrWfr0sKy7XaOsDecNCX
t5gnzETsW+yfDAZ89karrmlKXvyJk9NGDsc5DKbWGnI3s1trXCJUflRCtHFS83kSx8I0c2JZgA/G
QyC+xV0YUO/an3FT1+ccxcIss20sCcu3cMQMEuesuiq9+hT5dy1xk81UbRoNPBUkQs97TRbtrmOs
zajCBO3p17EQ0DDP9EWQaFBymhVX72JQUI0enazWJYixT8hKKFQs+FUELNFDITtzerUZXh0JZ3oV
fHn17+A38KWH/pXAtSnB28+Y+0Tgi/7tpxgo7pdFm1ZlisM2ePvH4YZJpD/15HiS/Wp2kBmBZqmo
K230C7McNsm8oCyJMxmh3ZnuKkyUi28JaOl8iJjxGkC1NwLVAdit5HcEdxmYqfMZmcczN3oHAaLh
pnaIRVDNvkc2xgsEZTqzfXfzJEigyv5Kd2jFQLZlUBZcATdXlujzCW/ZX4kNJ37mW6E+WSNy/727
mQV/05wCIHZNNYZ+0FXrbPcxKS2BJAnjLJ8bfUqce3JlMnV6ryZH3q6uPhhy3EtbyWzEM4r5PjEQ
r3jnHLhyJE4Oj/MDksIYbgVkrxPqHSuthi/eBG7S43xiaDpRmeT1fzfLsmkRTrURL+PF2w26sZkw
hIyPsk33RGrhv/2tY9qI7QUgzKrSsJHmJSX1sNyOi3IWpagm/b0uXVQCEcC7APZvWTfy7PX3IHDX
9ckqR956WHilQDyImw3p32E9Yw98SKy2ZnyLTL5/2n483kkkqoHRNd48xC/316OV44bJ6u7Dmv8u
2mFO5qig/zuPtG6rjp5ggA432XrkT1M9I4s1HhCG+XrFg4KPNNLt8W/05Y2zomW4DNLnjiO6zw98
HMaPzQCGCnzfE4xqXaFVMJjj9/LjKsaICwJ6Uuz9lr4m2bzjCI1o7CLYrSR76CMi7HT29YSXvwlN
hcasKWRPQLYIfRHRQHm2dllZdz0p8BajkIXHCdTqdH92mGrOONbq7B4lE8FU5znL8ftPsPdv45lC
FuOduMaahNRQPekYYQ1aqrKSfT9X2Oy65mzTCvrz36pjUMHXBzKOlshYBo2LgORtX36tOcy4nRHj
w9Ucjx+3rQ+rWD3sMh1mqLpyqOj8e87KDW7SGDkzKydrgUSE4v3mR6pSymbsWSSzLLP89VNYTgQ6
xUHHjNgUhaNAx60FjCRQrN+rDJVkM+JDAAKOHKZ5SnP0Lfs+H7xK50JMV7pgeNRyW6cP8NfZoFAZ
EkFvnjBwSJiFCA5iyyKeiXWQJNYzIEYHpcRmQrK5cfgvFoRLTa791jwFdMbTsgv1/I+ybrhlY1sH
ycoSYIo8lZVkd4mbFZcTMXmLwTIDGp3EyOIGLKzopZT+s9VuKsludMp5MUAkxtZBR2+2gKKzvKMm
70HcXWf4bytdohFdBlqd04do/+6sntYvj5gj54f1PMu0CiXYmREBcTZAb4fAERwtqTTxzGH1iHBu
vfo1FHGIEkG8WPwPQuSjDapc9xuZKcC5j2A4TR1eF2vtTVkcYvwwFJIjib248Vz4IF1IhyWxJV6f
RUyO7ObGe5SSe9HyvrMGk12PIwCDGXfX1IF/imy39ZMUZkzKzxM2PpA4mRyNUwbXmJyp5tT93R/2
O4XpZBFRqAWo0z6hABvxPpSF6qDzmRn72JPDa0vCzhvgHWSWmp1D4kIrEdNIoRw2HWVoOgdtuwxf
O8RXAqbKMnCbjtUoUfdNOO6B9ypkZIHDICmpOFafgymzFwh6XQTWEfyMRcoYJ2Mt5mBJnnKP51v8
VwsM6jivTPtnOgqQ0e5Iw6AR9JlON8/RzW0w/IC8GhxTJHpIAQXoG1Up/3vl/q6NUNrGrZMXCCMT
ufTJmWE+YjJW39aYS5BIdIqygWB2c4kvw7seIfuhXjDAVuS0a7b9Ish4xb9umrgIypXKAalQY912
sj7gq2/X7/BkJI2LZ61lAxogGXKUStlJYCgnTnAAEuRUHVGH/J467uMoQDRIyHUJgRVHO2qFDnHe
Nijp6LoGU+iFzcqzxQb0N+V1kAtFXDr0rt2V9HMeagpYzkkdwtZqkz8MUgM0BkFSdNBJEqlxYg4y
8hFZY7Mx7CcM2+b+TXOoEnfrfs+Tk31h7MSnOoqQ4Ip3XPbb45dSmeCN9V1JahhEqjE22j4MGWfX
xpnlVctcOnn8d8jm/3re462gRTCcD/pp0OfNmHiXGF3qpeDZDpEBQA7R2DFtR9kRcrEsEwMJUeDE
Fv0MhXrbWmmfXqspsYLiI/Z7r3ZCmuWkxC/7Za8s7tC24LHiqCX5l7rozt5y4T4IO1U77rscj6zZ
Q9XLMx7Ntt/OF1BUb23ldYIwFEEa6tupb5W0p4SFm9IftKHWZgn3oVkfF+Jo3i5biyvCgwtBDoyK
4InPCpsqwGmx/QBvdYXSqB/nV6mNWarf4/W9aoF6Yxq/Unx5/y5fdj0QVmt2ehrQsq6Br7jQVRFW
oRdjNWYb8y6/tvuTWy5UOfCP95dZ0k5Zl9xf8rgjsQt2+PEo5vold9u1Vef6YIJOFFxjxJ8j5yxu
4dTB39sSGjgUK4nibQV+ok7q1aJfGp61OcSdajki88Il4xUiA0UMFwA5Vg5JWYU3k2ml/G/dXy2e
m68H8zbKfaP+k1KJLZjlSCS4TznmfhR6LbZuZuNk6eLem5BiLv4EIY5lRNXtlevzbmx0HQaiaqCn
wxFqcbi03qpYVPeTD1ldOT7vhuFvuF3AHF/eFp26kIUp/2r0QXHuRBOM2P8OtKLLMRbFoQvZUe7W
2L+Rm5U1hBb0RRXnipctYxQaiFthXYoU6GgwOvdUDEedi9CWVq69i5HIFnv6RZd3Srxi6o7tSWlg
/TsxIAvtp66tLDEinSsYLUrT63gx0RciiPS+Mnd6rEYVavoJn8MdbK6KtkwOpeXZ8jC/DhRZcODq
EnEEI8vDsl30adpHGRPWyBdOyIfYUF2B80q/vs97F1tIpVjBi3dbXRmjr9iRIpID7NF/NgE1BKmt
QJarI0zTWZ01gGIQPdBAoWllyr0oQnAOmbWBgULId66De18tqXp6FTwEZZtN0i6zjOwhS0Hvlds8
fnNmEl1Pz1w3RXwNJs5n4VWdjj6w52Tv7nhgBsXJKjSpO8b8wS2QguWr/YXWEhIWsFXhvt9M2fcs
r1PFSmDmgbjZbNAqS5Fi77Z+QbdRFgMFwY4r6CfWV/lcl0VrNwBJfsya74qUlm/tYlamrVbK1lir
xlTa6buJvTMyDN6gQMXGuGCjTkCE0RQC8OOPOejTLDR7bLVX/tt4UwGkfUY4yyyGkeIaT+BTH1f/
KeX4dqrp4UQEP9x4l3B9j4XBFpgxJuLnC7vHQOVx/GuwEhdvvKCt0Kk6f5g8lO3vIA3y/1Z4ZkHD
gN5ahffjC7AgfG414J87FpjUXf3140JJacjFDwirNZxBH7IGh3D1F/ip3Zm1z2puTh8q8KFaFD6e
ly5djtLbhQVzvihA6J6afPzpTrO/yXh90wT05dg+R7a4Fgf988iPSCIRd8NpAU4gd3sZtGTyL3jy
lMikSv6XpxvH73hCA2fgUwzQs+S5kBrN6VxodlA4LdXzzUF0I7SjGQixjqB28NvQl5YtUfkD5urJ
70QJJpHw3wDppZKnz8R83y4Tq2cHM1PU98RDSUaFdZYkKwEcLfnlxdsOK6xl9uXXPznxPEG3BzYI
WALTznyHX40xtHqBK2NSreJRFFxYEerMInoY4INvZeLZ97j2xL1iY7HiWvU1KCWVOJZ9s9kBJmTd
gcJpyqZG0HQWzrfTgrGe+2JJBjV8VcBb7sgr61seCr6FjwpcMHxzDoowllesUe+gbqQmNYlmppzw
CbbcEROkGcScHakCB0sW+xzeaETzmGgh5QQ+OGKXM4pcBkQkq+ZeCqr+5i+uqQuVrAwAZOoq+GPa
f7CrvNTmvt9rLngg5p1mcceWTOSZ2QBkX18s8sUKBcP7lkytDHG1I21RWz9l5WcV2y89dFQ678bc
mtw/UUOYdHnCWvJ4ui5t0+GN2TF0Yfitr5us6zS5Af6sSV4DxyudbUZa8xy+EC+x1Qf5BX6nTycw
zbSYzsLu31pud0iJY0M2x9b90anKvHxzHgoX40e/nUGk4W3sSmXWzcJ2d49Qf77l2uf8rUAEK2qt
I7ihjEKVu81dtcSMa7BEITJLD1QgBf1pp5FDPLfLhkIxN1XgdWzVfIwDoT1gVIjo81BrEOO7OIgA
BiOcj9l7Oa+YKq6d788FuUZdabLznlAW1oj9H7pRLHBy8MtLzUTvUgLSXCJL6pmWGlFPkarpAkaw
qRUDx5ROobm5i0cdOA9WkHSookrCH+LkYeMbj9u16IPUH3bXWSP4LROOLtg+wPJW7c+d8gfKJjSV
aZMD03fZZd/9cpz88nuqJcK4smACpgv5zXGba16eCcvgIUQsyvGqivJLHctc3Euu6pI04F4qKHGP
Ub7DTd4MmuDRDPFii2phvmNEpkxWyiB0/AEM3WijDcbhWMunGQNdqpMpR34J4vyxiL7GfrMIh2/8
L3/+9+1/aBib55rIv+qrHg77hZQDZlCCHCBvLpodZSMfWM4valezsAWY6nWQXyGs9xv+X+OaM4xw
b7Z+hho41nuAH++EqW8TsqC9zs7ar9el6VTEQLA0VskDGDrtG+ubD5Y/y4n5k8A3+A4hmKbTHiCh
ofo16BFsRqOqcQbKfLx1oCNuL1/OxtaTsebFcX69SFSOrxeuxzvQ6+u8ggrtRH3CZxxnLtxvAR7K
cxiwJiyGrppM/nH2twRi+ISNpH/DsVhpBZH1v3eI2ilIxxwq9oFf6XV7yxq/TiGQU/DTJ8RsSz+z
EgUSFzHKRULCNDi7QBOMgfwZYQNoNGCuW6qYFPR4DwHvcZ0IKURO7rq5MAMOo6LUQdaDwNKl5/Dr
viPq4tXugmx6nMF0Yn7qn/q4dNiuq6yQkwXv5FrcRLBgJ12w8Chd1hOEQouFbC5ykD2DgU4V30IM
Xlkr8dOcH5u/Lif7PfLs8Zv/Q5OLWgWQReovKMeALq7C4Qu3r8OFZ/Jzv+w2ttyGncTs4nupPoYD
KUVQYS9zE/ryHcPThSUZ70O0ZqcY66OMeb3e7gLUzsSrIpNoSuxyIL66gw2K+gpL2rR+XuTMsQeW
xJlXE/Lxs1vhTpCMFxj7BkrrnYj7f0pDYYnD5bvnsfWK1urEC2cXAPgmp+V4aeV9vpI6A+NKH37w
Hqf4hw+Gz5Nud3T4vGxWU7/sIxYNXwojbgvW2GC4ZjRd6whgOnggZFZm7PdJjDcmvIJ11VYgDi+S
ExNd6OnQCK3JMH44IebUupxiKGi1sf9F2XGC52DXy69kiImUbdhDjMoRxEk4uP5Jyn3BfO3lEdoY
+sG0JWNiCC4uI2W3aTlGeNtGib6z41ThMN31PJOW/Ps9gDKr5UpIztq3qzKXBLubrpR+5Vm9nui3
ZiA7yZDktDW6AlgTUBzLibmowm3TWXiXsNVf3Rdorght93k6D2Dq+63tTrQYzODChpsWLhBwolN6
szz0qvFcU8KyX/9FNYYiK99T9o1FoRnatZyEWxuyDa/8iwvbSkQ0ze9xJK5Iq2l0W6ykpO56kSNf
32oNCb+8NLGW30l+lvoBVCY6cdeAiJEYU9Lg7n5xk+Ip4mg8/6+WvJBMXkG1/S1H3tNJ7nvWFOIP
iLvmQIcGUaI0xiYVCz2/NlMHFrVqFvgXAVIdS4gr1/yDgeWtEWRum+S5/64QjSupMvTfA4d0AwIG
57oOB7vB7uCwXUNFbzCowVbXHcW6gsbOrAruzUbYicwd6dSayBt1zV8QHWA2ZGpse0oXJQRbZ/cD
MQ0s4RQahlzrXNYME116hMDkGTWlkHOvzyZTHkG0KIMtCNGHqWzRDAiVWFMzz0kLwfBh8k3x8U/3
IEyKcg/GL7L7uhLuf5rbyBZ2TgjcVr1VF2HmtLIhq7Varv+CuD3f/Y6XilReeUYJOc8R+f4mA1cK
IfwAdVMEUd8ikcEXB8cw3Wek1CegMyLF4WhQugUvNG6/2q7mpwYxtoRzKx8IFDLpvGRXK8JAbrvu
1kCGScfzKHZw/RsZX+znpPvUCBPxElbdxoP2em/jNNt48XTMDgbHIBva/mQEl+IAuxprOjPsFNBM
jslfZBML1y6Tr04LJ9kQ3qj7l8U2UmHDMYfdttg7+qrcgtnuGqS70IPL6O5bcaPwlNwU6CD3U8U8
5yV+oXus/4sy3Lgl6TQa4ZNq/uMflxSIMkyFO+8qlnsgMMrKme9hLP64GjctP5vUBqKc7F+FtXXe
5bi2FMz8qvDan/5S0m6TV247aLtbjvAhx7vsEMK3qLK+ZrljrXl+XEpRfVplMLw9Zm7lUOFe+Qsl
wGjEMHi3AzkV2N87yLmsx6G5W40b8wNQ+88d8mF6lhwJBWi9T0YfRXAN4cAPAdD2fuin0iAD9exx
jX7PqgCPpCUU+ceG5F6L95EKrLOBvIC2FTygmw+DMiQAQeK+JhI1oentoUabUR4ODheERqBx+q3U
qaFWgdixOjtx4roOtgebp0l8zYh2e45sqngY4G4vylJt+twproEF567mcmKdpojUFT3aDtxYFjlY
7HsZZ74dpLQjQx8BFwsM8YOwC1dEkHeOPp8v6OJK2VVcPHIrG/Qm7nPF8+qfug1m54Coy57p2ECT
eylBWSNj+2h90R25t78muO1CSYHKxx7JlW36wsKI6mfckRAikdE5TGn8PYzPfvJ3IKKh+1qk9V3T
jWcfieNnwka5cyogVn7baL6v1VFYm5X1E+TTvaKk1vxO0r9AmTI5QmX9K1mCcuFIRhEESybnoAr6
QCOJvBc4cX1DR4oINWx2UdW6XeqvGXo8TFmbj4feW2uhc181UdViIuuKjv/MORN4mHSB5N35A8Yf
QaaDvgbf1U0YKVZeGrWOW6OYSfVuJaUdrq5HCnGCMdaNgsiEDFZfoTndhGay3r40c+8H1UkJbv8W
ynWNEH4DAKrK4Gd5loGeiWeMSC8A1l7mwmsA/kdabCPUKilrrANAAEyZnhLkFfxUH0b39t1WpoVK
YfLyNf2XzTWLQKW0LwefEZRekAgMNwdKMeSaHmtcn52/Ltw56tIs3oOckuZdr0hk2znxW03FTgCp
nN+9B9ik1Ytb561NN3UMIAYpgGL5Rn95YJCm+zMPYJFFkiu7m/9CKmoU7PU5Be0eVSb6t3SAFNLp
rDIhDYAK+8KjMF7PV7qUNX3wPgaXGe2AjgA3cgI+B7xo97VRd56Ylv1Bg67fhTcnkEqnM4wbHeC6
CqCkTDw85OB1e/6HyeoqFzijWl7ZzmFcC02a5A+TDWMRRqAiWdDlu9LJ4baF8rmaf3G9oDSmFqcZ
tPFqt+VGleguAFb5sqVy9wj9f5jtaF0bUGJxpwUZtikjOtNt4uQcBaZCINR3U4CATpRSSY9FDlu8
4ERz3HMh//o1Ym9Y9b+P5TqoauuGerAsOl3oDPgYkuLscpfwdZic/hGVv2fnGZc2rKDWOeTgDlyX
SSiEnysDLb2lXOYHB5b6o3XT9FGOCsLFTNlbQUw/u1FAZnKIee6JKeIZRm3HWJi16Eo2oMS8xD2P
tXiCls3ApnNxyCb0S+zBKWd0r+QNakeKIhRMxK/gxyQjekQxI2uY/MrR5Xir1hcOx4s6D/TXB4qs
Xwkw0eNYFWqZ2MkSyKVG9ltyborgvG8WCzTcbZ5P8pRxjOiZOvmx3odm4cv3tQRU3OalL6+m9n1y
tmyBRSBWtmTWhAT/ZXcT4Os9q/lo/Nsj4xZc1SswLEfnRnxrcUsz3nceh2ke3ox35wCYi/wL7b/9
nKeujnfxGiiZ/7Ys4TNB7K+h2kygak3C3IlE7fNpZRiSqVXBh3t1tuGSPF6N8xVLLQ6LiYOJlMEL
kIizMx4SNGWOrKI0cppWpCStL7T5UOb1fkh4k0Z5F37EG894j5u/PNWSHCerYO69lFvcfPR9mVtQ
hta/nDtJMsOTfXUQjTOHkaS3HxMAfOYa1ZR9wC8lrrWU8H2dDaTSRnvrr9F4SM0vr3p7+P2xMB7M
7TudIFpYuQGhaGG9I+hPQszT4Y5Q2loOG8mP0kRwN9jRw8Y7+44Zq+zIiXUGw1dXWYDGGvRM84g1
RuSE1QfuXPK/WTmz2HiFe2hLNxqkazsF50phFOFeM5IjIqU+TNgMscwU0QSV4AsrdLg3pGxLskK1
egnPTRQKTu6+kM0C+i9zvMGrxkq8cZFSm4syy0UTHFKnBN9dKZsepNgKiDsI5M0XoQfZU/uppdHc
ughd3u+JgrN/ODUQ2tHpsyBRZmURIZloIpFQR7VBUWGgYDPtJRJFOooOVecE5lT1e9Olb089K3AB
JTevVLrMfaHjiHky5/CnaiQMNthOZyTlCD7OaIIPSk69R1neOOufIP3xnDDpNhHxW1HdHOo2F+Ny
iLlPMBEjQ+lkQAyYckSMO0/xpg8E+pYisJ0RgNYyxMNpgplbMGRXxOYONKV0GTNQbkqDaOnrMfZS
fGGX1/wdVj1Q2/5SThXmiEUY4W9UGjop93UUZa4P7VgRlXNKZ5rOCEXYColjo1dBJqAeAEE8eLey
XEb8xB8IEoFZwyWnHpbsgSF35gojUfkwk/vFernxWGbErEKRSZQDxjjjfClc9Cn8HfR/k4/7tWWU
ccAemKsEOn65AceYjS1YuE4EtUeBC3ZPgGilNinRj8fMTiK6OAEzDS/5/YfS783bb8cWb7C+QqhW
0AZHCSAoDt1bE8FlziqYWIvgjguKyvvM/0hlOZHkYdWGh6Nh9AbaKDjhDfS53mFq1mwYw1rXqUrJ
TCTMEk7B5DPDgm8qSqC2tj33qPHY+2Vss4a3k7oo+9KT+jPYJkeFk/tpoc6HEB+cn0SuJvtGh2UU
DX9eFPUt5Yn6LlGeZxJN5qUyxK+4ep9/ThSa9ZkzxiPpc9O1JVEp6j29u3CtgBICciSDbQ8g/zah
SNmCtdcrUF7mK8AAEDauzWOiVGmDeqNIfsi7Up2BMT1eQ/0tYvFNg4xTnDjM0g5K9dWwxDFb52US
+q98Q14vLHIpw3p8WOKejFe1nkBe5uvncAg5uHO0/lHfchTZGjPHSDyN86VxQny2GcOwxZBJqy2h
cHGNJBYzI4atAW2dSUBkmqfhm9WXfTBh9QaSKbrvkcoKYnQDtS90oGw66jipWD26dI9hKLR9OUW+
Uw1tsGOC62mgXbZkekn6fmTO1UyQdbP6Zv6fIixiWuqdkRwRxzAb1Idgm3TNAXGDsbG2B8FDSQvo
bBWY0FIYuAmEBHEcZX0I4eLLHmRK+J82DPdCFEWm9b9v0TsZphTDXV8SU5SetYtrOsm18JV8Qo8j
at3mGmeo/GZ3/pqI/dTVTGHr5ylQYZzManQU2OpbBKb8+XO6UDUwgIbFGNXZZTHO1D+By7q9oKic
ZGPLQYiymPtZVnqAFtbeWkLJqtXXSMQNfy0N8CXXa1oYGN9hfEpn7JaK6kjxhN/csylZkofkr6IZ
d7hs91nXjw34JyWinl5qDNpv1022hfs5+EK3QAgOnKMfy0J5d1fYqBkhhPeeNE5cLICx4O+SncYY
ykFMh0AYtgCJ4PwpwME9hrxEr5F4umQy6egPWJS4XF9zK3V2nqZwAoUvpwaigvJ2eErPWDf33TNn
W9DWSiB8gqDHzMhde4jNaOcrct4CClybOK9guZCutKaZvrK+j5qK1hX3sQazE8E71ET37+7kFvw9
WxPF7p+whZFJm4I3eIpClYTOMak/ClamAzixBZ3ByFOiuuq8Jj4otm6u9BVSE2+6tl+cbEmm1RJa
a++KoWGh4kn/YK3USzoOBZAMqrChrNCATSPxbasx75BekUzLavtjvF3FZsODmXJZFGb7vQDfIAnB
A2CHdo9b0q0p5WB1JYYKgkdoRH4I1d/5GhJA/sxPQTRWZHoA6+qmRt+jGOX7p6zc6PDXbG8ADjhm
rb62k5z1Fzk4jaXVV7BKHX42XEZejAJBVzsD8wkv9gcPMu/bkxwD0dBMEnkz+2YbgQmB70Tn9P0c
bLXCjvW8uxWvO70vCfkwr8cv5Nx8AtiE1USi3e+L3awiWFMJkqMwmP20S06gdaPrgsMTxw0BJq0R
zBKhA9agW79CPFDbn1tfxn0fZ/yjY/+M22aYWaxwG14JAlcc4ggSxdHOXUJHpBPkmdBLfMDJCTfV
4ltJOSZzJcR/MfcQFfOQ/kpAPzPKrN2Ok4n397NiSTz4Zv18y47aGvEMYhb5vYLRipOjiNUlTyI+
q3CAxT5wFYnwsB5vsuQ/fHn3+oBOWPiZlGhCfG92f5xgIH5axD+el134iIMkBWZHAhsp65gFLptS
bGerZrxjv/TQcJl4rtrYL4/amcmUm2fceIwDbNa6zWwV8UzwTi5Ce+Gt7k0o3hBEpyG9vQsE8blO
wmqnISMD3M8c9yuug2RATUL4/Jgk451esyE5NPXeJ84mvm8gzwJWgSoYHF3y8k2EuvJwLTkktC6Z
D+WyRbNVvXVSl8CDCXr9nAmBrxUQjaIPefR0o8xKBxJehLFvEddIJiy96DEWU3j/B7P/+UuJBU+D
1zKy/8/Ef2moyyEiHe/s1pgBKkaTxEijNcttK9ZxsIvJHAMZEhjK/RljZH1TiIn2Tc0TsaOkYkBZ
05m16t/2bhaLqUytWT7pntOGX9jZHr+xarwfnrvqqzfDuYMNjWiwcO0YsOnzjTNTVdCPCAqXYNQs
Pch25WwUnBg70LLWDTQsME3IAqn3iWqKDXXTEKvcl0BoC37fS/bM/99d7dUAm58gz/Z7jO6GMmb9
65Q6EtcEakqP6vlfCk/qmKgmSkFboNYtpVz+ZG17/q4hVNZYWuhYCMwYHPlkFJlX3pUJs5TIw4bA
7CRr5yJj6JDjJq9UpaYTSz1JK8kWwBFctysgqbjxXxJKKy5OHGc9xkiVRkVwY6KO2ftdHgbc4b7w
9VFeOrJLqvyRqymvT0xOqTI0WHHGnMDMUoii0rCzf5BWcFoUjyU5xjmoQwfNNt7Jwe9Ycpf/PUvJ
09B9MVtC/H041DOOxyDI9HWg/t+b8/YhRCQ/FDKGHwRTPLFOnv16eF4ZW36UjNfTQ7vEBaCYfZ5H
u1hXVIS5JjgQWnx/bw4Kq2fpjCL9g3FE6ZF9TiHMkoj7LTwozeIUln3Gznx3MT7zwRGduHqaKGhY
06iEsZ4HFM9Xs0/6/Otdj1JnF9GNHtHwXOrco8JEakscQddDmaKJbT56saFWUf/LRH19HrYB2Vv0
whbWjrTnHIdoufTD+a2zguYP1dFKg0JWzaVywsE585uyy/nGTwcGh19Ax0KOLpzBv6aUhbJ4kSEx
eiT1b1ZpPfNBvh0FQkOh6RAgdaKGCOaeqmxmtcM+y451qHVaZsTwwQlNxWeoaGlib2GcvUUIHqLl
BbNvwHNS/jpsNa8/wfNuFAgha3JaxLluddINjyv+p85Px9g1F/9Lpqv9ICQOD8MLFrvd8oxFTTyl
QYu+UUdOumwOelo1xldSXdWSBHU+Td4oHERYoyIkqyqKcsDE55dLdOzjfNddTrqBeqquEr51kSf4
GlMMLXgAHxOU4kiFWkDzfGqv9X3WQpBebqcYAVhI+Aop8oCo6ph3wOo+uMTzfPRaMFgbEpFH7NWK
JNOBpiQsVZ9+OL7FAk7e1shUZ8ct34L9wcBveDPfWjhQ6CtfZ8LfezdAmFnOPaXNVsADJH9XiYi4
2ivIEt4Jv48VHe6V45T1oquDZhpiRlFkdA5IR/cLIw/RMDPYal5ORUgCHFlgkNe2Le1vhI7Hi9G9
0xuWUAM1RBkYaIMr22QkoCPQh9VRivoaugEfYcsLpB0MrQDuerkKY98qX/ERrwuKojI+0MnQLO5n
Dit/0tpETn94waNLsPDpCF0iAMql0B8TI1daryhqrGmS0WpG3crOMlvjnnkJRuqrs43diOcJIuzh
kq/oZUT5rnCmMZrDmOQForg2Jk1uwj+gN/jkoraVQhIrxcpfgfh25YgOnFo4skM4MrKuJiE0yhqu
bPQiLs8UQ+xNvo7VTO3wA/3hbYdkcayhzcMajonXh/QJlZDLjPzJnJaC/teOoAPzVrlfeiV1REmD
ajHC79Df1aJUfHnrjnoAS4cXTJC27l7LFvMu4ntvWLgOJqU+tOjjIKFUyw/5cNMWpQ0fGcbDopJz
+W3wFWdcipZQtZU6IZRAfvxoxn3pk0W6x6iEV9gRanQuxGQ15b5i5OG4NJF7ex1v9f97pN1GRBzn
S7ttfJpa2xFFkE9UxeMMl06uBSJkxbdahOqjwJfP4NLdMXn0CMekaIgsyd16c/mZcktI5loYdc4W
cOmNVtGxII867lGZuiuP9xftkmcQmtXKvynikn+ce2aKb+bXpeaN5P8xpxE34Ib5ewTM1ismXm7b
129FBjQQDQX0q3PseeEMJl9tOQDzKhKTkvxJPnXWkNK+w50yQkmOKzfp+Dc1clDR6NECCCZ4EVMM
BOzH/Zvh5NihiP3/XVXEn2b1D0bkMvr2KFjJHR69hUmGNWup6amQa/VVZAKCruDjGl6ivkAEZCgA
9AyZ/15yYae0m0prO5JQKwL7ubMb6QpmCtOq4D/vzWw5uTkjwkw07m58+HAAa8+hzwtyKBfcNxp8
2rYTi9per/tGYCD8d0gfy8V7jZ4SkML2C8ncYBMJKkEEDY6CQL3GXRdLlG3EW0kXIXAsf/mcvtNg
ZfnfBQSczQtvlc9wJtnJ+P1LJxlxhT6UigPVYj9dwVY7WZ4EcMbT2OBWWYQuJ7aKc7axzpcvmPiK
H3g8A+QJN8yS/1+P26D3RseFIH5uYi7GDK8GiV/yUWQzND1kYl85fZQSlVVioeM6JxRLm5QXXlTT
akVvQL+wXQXac5z+1tx3/gl7vaPJ7fCgQqCj7DOThvTnfjMrqClXNES5Wxi5F8BPAtk43qqed6ZE
5ZEyKEI/fqHDXHrxkLfGfDa7+2GnjlzKuV+YqiG2mWvEntB4j3vk9Sgm6ogTqql4ha1vCWBaahMh
Zm1IuzqOdU6Ogk4jvquEPFSP3KS26StHVcZ6A5YxiCGsPV4u41plV3KlP2tRU/B4FpE3nmbQLH0s
W/1hmQNstVxkVopPGsQK6LS5x1cE0p1Zz5ihJGoh7bEldZFxVC0pRxMm1DXhSYPEgUzceTAbkqVh
NzLTYSy5gmPMktyiSdTGXBnZn+MQDmcuLYcqDtI6TmYqSvtdV2/rGPDcSzjWBwfU9OAtcpeoRmp2
fdwGbwNIh9k6lKDkTl0VWCvVoiBNqRzwZtjPB0P0Io4eSnhLTr59QDfksZtNDudIefbkqV3GhDlG
wKmtlIJpwEd20kNIjhAeeJLo1TJiv0pebkUn7Z4vo3JDOp8Ht86M9nTPdjsoPmB9UPicTQfTFCvO
BH0EVEpHxW6Xsr4p4x1lMzWrNJ2plahXAR9r0oOvx9OwdV5B8c1vOBgx1l2oDfDKgYRqZXbsxp6p
WrcbUXPAvLKQCDXHhAGHPjMGFXgRZT9jRoQkCwg9AGXEWRLoY9qOA1WgLhD7I3hj0ymuOE+cTrjQ
4w7P0XX8narHFIQv3XhPTD98uiJuR4R9aubi8yQvkBcPWba+j6jNO7SSgZKt6nL73x+r3Et8dz/C
DeQL/MgquUArK/Uvy1gOun9TXkUeYhdiyQLVDde+Lu8e5tlXXsI0zlBn9UvOZqw+uDi7x5cf1Wta
ZkyClUoYw0BkpjF6gOTNSKzG/HvLLoOo43RqwAP3k88WxsFAmlDJDemAxcvxGpHuyIKT9IvUFJG9
waHD0587pAh29AkL/dJY+7T9zh4qEvgkcYlLjGOYJ4ebSwY9zGCBgE6narBlVqzhwwCfuOPLuTMc
zF6cviBBnPScnGwb3Ffr0gpywV2nAcMAFvufBWjL4TBtwdefU3HSbv7dGzeBiofDeCqeiwtJUxuQ
wxVo2BUYHLWHyd9ZwePVttoEKZfmGTK3kYO8gMAFxKXgpaZQqQwTMTSSaQLlInHCGJ4PAuL/+hP7
sjHEoUMXg3AdBkkC24tRSbG+UQNk6rXxFIwUEB9Oi42Ckb2FQQNH55KqKxUHPV2NiCJ+8pP/UKcb
Py2c8kNP8gmylSWplxJz9sUJRPV/d0OxowRSyKkfGvNbW9dEKQE0vcZ0QL5227+U1Pc5T1PofYid
aB1uAsyqaburemtbX0cayjVK4tCn5FNpKPVYv4t6UoEgpbz4s6WMHTczkl96Zbl7spZkvmTjiiKF
Nu5kCPcR2YPIocdx0Er5CYKqb5Hs8X06ojli+SHS3TuEDP/3l/H42kksbR/6y3gvORSemxWwwrwh
MdbqcE5ja0fmYma29YUvIRY7LHV0rhMvY6apsKIQ3VEASYgnWU8+9Qn30+tzGAvAtpusGQDvk0KT
TRB42NDog0R4PgzR4SQNuXbN5RMAnesAxMXPIA5D1eQE1VitmVaQni7gGJ1fJlXThadYL84nsnZw
+iFS6AkzyM6lZsR7t3i6xfUlxbaO7QIn5rX4wTlVRtQNGUmcJmGwOXsuTQ6wx/WBRUi9IHpCAUT9
I7MTwfvTmL2cnRZcGEm52c7998c53SogpeRm8lP//LiNs3CVEtMvrS0fZ54jJQEWmb4zWjBu7Y2p
Bxs9XwTt9/CPzjMgPD8quqoXquyhTC720Df+TjBIMPrHYYnumCApfnEhAPSfr7CQ/Pc/pCIAXloO
+jsLzxxZNSVu0Lo20HX0ZyQGWCO4R9bWjEHeijRee/KtDoDinrHQrlqDWtwvjyVoJiBtlsiH7l3q
u8tGSZnVFuGJq4zDnzKaeYrsRkGk/J9t4o8sYq489ac6BkQ5GPexQ1OObiP/5A+qPI2DzUuY0J8F
fAXMrjQNgL6+A8nLga4ghuQAZId0U8L5CUqo0eo23LaqkM9gk8uTxo7Z/QRt+w+5vV4onofLbVoa
hoIQXoJJXV6alp9P0Uu/uHC7jMZnTd8QAonY+EeQniyvvUUlxdQfkGtsOc8CIiu00WzLowutbn82
QxbW6wF9ih5kOw/8ELNMwpK65vDeOsC450A3SJBPLRKuCDj/l08sDx0GWlHRjKcOwpXCwdtcFEEi
Qh6W68u8tAmpOsfl57a6Ax2mZ5e8lZ6GRueATljdVixXmPmWOjo4t5DCE75Q/oWmtd3dFMmnpiGH
wIbdPSBUsg5tsz2hdB6FT1ZG1KLGl8jyFnwbGpkwirm5xlhEh4fyA5leSzVO2sKipG38B7RXSag4
s84w6dEgoXC5GuXFxHrBitKFh6UoxYXVw9l0EABaGSaw1fLoa7kJ4afilUTqq0MYeswyD9nne5Gm
s15Tvi+0HM+WUCxtTYedpUB7C85P5qIK0r+wLiERSSUMhpyropwV2QWsgD1Ln8kAlNx98A582VJb
DCreGmSPYb6FfOsmt4KFjTkOb6jkJJw0GZYEXrMjI76t+HW1Qz6j72qQgY/n3d+MApMlLOejSou6
vu1AgKZKnbU9CnEg8dvoNQgNL5PGbYqqqplbjrQ6eiv9aEk0mYYupkvip4UdKL5fPlnudCGUq70N
dr81Ewh8sdSw4v89NgKc/9e43ruQ9u6T+fzpa6x4vMxdkTU0cJHTckSi+zHRABru6yT5zGXIBqmU
2fGIFuJFGMGdwiwekz5SMPBi2g7IApzUAlONla9okb5r5/nEYOxu/O6KpDrgtwT3v/hy67jqtyIg
+XWfQZ9Q++PCps+dgzcNTPGL7qotf6WGWtvH8DAsvMrsB2gKBl3O9uOeC20gAlS5CuB2sPpLV07A
uaRPLcbA/sRnLvFmlDZ6UgW0oYxbOofQFc9E4Y3Wr/xyPnLMxGisikYGvi4VaVB93ALI95sTT/Ik
T32+DpHcu0f1+Yfe3wqfLAD2n11fxGNOC45/sMfc/tQt2DSd3/SIDIhUPdZYHP6p4b53apS1Cv7X
6ffw4Qr9Ona1nRqBckO0rcSHl0AuWU6gOtSgjgeyxwDw99bQi2wM2SCxwG7F+DFCSwOBHlkBT2CY
+0GwHWF01NFbhtUQ6ZXVGMYHNlGLyTz0TF6mHKU+0DdeXUxCCnFGLQzvRVidot+j6rthrP/eVq8O
txN8vZ7bhXMtbz134ZhL5AIG2e945JGbiVuBaMbbhwZ2/3F5SED8lq0b9B9qVzdvQVJ33yxxoc2O
Bcw0On8l0VZbZaZdxwdrMN04GkRsgiVa0ua0ygcS3TP/yJ/hTM8yupQSkEqYNlhfjscgxVY9ZfJh
L3uMYl2/u0bETRkcSKniU+cxWObuj5ljvTMR1PyXBGNHKKL74jcYZU8otp8/uICwjeA8XqHnuyCe
m4PMiRI6cN3QvO2vtv7Ah1lpNxNIeyfxhDTspmkrjqs15B+RQS28TjirKSCG0hKwypPbMQUsmfUn
htFWb8fX+f0ktPUDVX3UMGA5wptfNjqtl7unmZ/zni/+3Br4cliRiZ0Q9rPgjhpYiv9sgn2KXhlk
yDSqCyJII0LzXrdPpECRgHz9AEUn+Z1aaVylM03O8MULnrVDb4iIJtjtY1Vizw/GH+4wtU6sF75c
4KRdq5KSM6uDBTOtYu4pI9NdSNrwwfbMTYpjP+pCmB4RQ00SeYJi6XbzYBDyT6E85tmysocKbNHF
q2I9stnm8jMr6ZFliRRXi4HPVhPbHh1oPO3XXM/lsf3A7l6osvph6kuQlObNyHAQUu7RI0v2BlbJ
YwPb2n8j/YEMagYZ3l5+iJP/g8X3/5nkuFxslBnIgFwrqz1yADJ5Hp9owWu6mLZWlorMoRxrfPW7
QkP2Vy0FqhMEdY8+lIe/l2us+pP0IkjDkNbKf2hc/YjMN0hrtJBAAR71wyWCzSK0/m6QY5pmdQEJ
5pug6EE+lcmBq5TIwGFnbjbEFlnHMsRZBZrbxj3wQJEfVrKmVCpRgXMI1AzNwtCtKWEZAx0oBqF+
xWjT3MDjdAE+7zlH/5FLWKmOQsIjcv8v0QM5bZSY9PIfw4bCkSnp9B4clFyKI0EmnzIgkwyY+Ovh
KE3/npnB6XALniM4ncVv7liTLMb+l9w/VinM9hsuMuVES+Yb2ri5UwJW8/dnJhIKWCV+b5BDyojp
2xOko/SI5R4QZE1efRT62kpA0TaL+aIBaqSwN4a8P1Cr+9DSpTpDh13pw66vlSSKEQ4PhnLd1eR5
T/uFu0BuRfQHJq/Alj6enpxUCkhHtR6VLXfa5aAKYAxdXrENug8DVatEaQMlEbG+P2WOoVLManoU
eQM5A89GHJTWPP0BbCFF/XEIcbX4gnqyEyDLpLzH5PUq5TJ79/TPtNPFxzOWyfaDDRTiWWx8Gj1i
oeBXbrPeRwuz/Ti+2WKsMRtImRJOtjh8WrJEJ3eHO9TUL2Kjzqk5hbjQYQZwiEuH4EYhsTwq7igC
hpl/uMAQVlESkwey2kEm47VCiM//cjI4dyMxFWshr642w11+ITlX7AJ6fQHzDLv6KEJtIsUB3U58
xcAKvOpbb/rdRhunlP8zAM7doUqiFUO0cCVTr8qt+E4rRv5JlYFkvVcM+ChwDx+6R7aHYg5aux2M
qN4+ZcCoNXEqvsd1yAxGWH/Bfdp17JKwQOBZqsOkQ1e8AofqBke4HjzQ8df36AvbpuvlptWCXLhk
JgitdBd96metcgFUsvCQRhlQYWcbXBbfcmL9gPdyVTLZXbR4WPlQB22U9GvEYO7grIQxM59lyLlM
GMkOIX6xFHfzvBqwCOVlrDkuMRH9SuMkL4K7813hV61Y4T8oPvt7ZtAPOy9b09dBkhlkYWHLs7yF
Hn8=
`protect end_protected
