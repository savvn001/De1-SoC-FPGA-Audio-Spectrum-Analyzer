-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i4K5oQJ5WabRT8MzXDFrT9TbDAc6KH2jSKCAIsuzNDGc2Op3a1ujI14Djn+AlZqKKfM4Z5tI1mVy
hzD1f2bTLjVwuVhecB9E7swCUK3yfIK8o1NU+xKN98nPNkHnhBr0DqvpPfco9W76EFICQ90l++D4
J+BDumG3DpZ6rEG+XbdBaAO+LT/uXyxcW+wFV9MjWOXuPatLsb1Jhhai0l4L9d3HZpmJk1/hBAG2
u1ZH5gXrDiBtslPP8C+Lea0rioY2zbMoaVE0kGNm+tTo6qt4dhWsDmVen6E9Bbkc+TbmRmaIealH
oL2d1Yigo+HRbzkdXGnjIdxSDlrrHUuI/oIrjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
vv3YBbAQwxSB6KDL0e2KyEmsYZYhsrbPqhKfQuyHqk7q25tEhIVL4TtmpglZd+xLgFP4frAW10ns
+MtB3UXYPc8T+RrxYLsB9ZkjV4wtXISBJXy1foT71xfXkdPM818DK/V/LH9/IfMgebGf1niTgDoQ
y/2LNsn1AMSHCj9AZYvaKXcaqqHcrm5s52gt6qEPStPb/zZAEhHHOoK+8p28HpdLgJhpBuN8QorW
DzYJHUDkFypqgSxsDU3DzPobajzfVBMPpTCHdS3Ik6aB5QwTS/W/QxswZKWl6YbegsgjpYmyCetV
BzSeAFQAs4OYlFcttRPsaicldZZX4BN6I0PKoFy61MuJ2PrNdcY8mupkkSe6muWo+LqGscGHAb1n
NgTT+1B0kbpB79LbxzhMV5p7P/Zie/yljo2Dr5R2RPrYOOwCJtqaIDsdRdVLo3C37WrWQ9M+gI4q
UjI1lMG6zXuTL6Hqj3H49kbZ+1QB9hzaD3lT7Cs8MgaycIahNp409Yd0qpD7Xa+ILnNOZ0tzrgE9
kgzVxpN1kGL4FsHss6lgCLoN8DCp5aiap2h+5WUFBkOo5NXPRIvKgPJaVAgBdLUACDr7itfULj+J
UQIbrRAoSWIpkhsqteW5+8NDjHzvb5UCK2FU9IgJFJUNoPg9Y4A7zavxbG+EI8PIJWEBPJu1xhzq
ZNUkKupnIvAeg6hpA5+4gFwd0IyroFvYJH0aGYHwLnS6GFBPwNPasbHCj2O9e5I38hheKlHmXQ6P
xzI5PtyOtDmmOgknUndv6VA86CSG59N5MUe6uGPs4xIxgxoHGSTlSacun8ogmelXY+lv4wsvrFdF
4UDKjlNjxqW3MMfrxe86kceRUaN60633JkD3+i5GwGDHeW2OA8H+P8opbvzYsIwMgjdRSpQ3pOEo
jyga3L8mazwKPsAQW+s93ewVS0lgaxoB2fX/krHYiGUJKOZj4kYNHCx1OL4liOMrCQrKNd2AaEBo
Cb4g7wCWQoNAPiIpNXJwLALys5mXtdgR6nF+Z8m7pgY6FdVxb+czJCKuGD9FpidMfKtVP65fNJ47
Pv++bWA1jiHm9Jl1tS06CNyM2SpTLYUfGXawtlZyBKciMiHj+Hn+tmKcjO3iFGGb3SyczMm5adt7
Ru82Vn/ckntBAjqefBMpvHedO9nPS6OixElWEPIniU+XUV6lWcrAXQ3f1TXiPK+VkT45tEuXlhIC
RgXhUFYWA3YgML8iIn+Wnpo4gOLvteKLZR/6w/fczlrrcthj7Wx2D6TLfMXp5gdTMKfS5tdWkXSj
k9ZF+gRDm/ahKAdLFcNVIbs1Xtt31v9s5qA0vTqbma94W+WGtWkYnFjJADfrXarADSAS2SqqufqW
fS+1XVbgSuxdsweeM/J2/JFbtjDY1pWKxFwBZTs63JYZFdOd/OBgWYSwiqRl3ie5zfvc3NNQbwNf
05Pz9zjhgWWk0hK+iddcY0HQ2FskiF+gKfUt44Ws0ni2S0whikbGhLy3VWXIzPS9hOWi9TJaKzqK
NosfoEKjBWo2u0a9LLQ8v81FCfps9HDdZR5wBWIgHlx1IcwTW2QIIjzv2N6gH2PDRlNdfTaT8LYM
9w4u2tE8dX8W9nxRxSYjxLGpiQiTM1lmGusIJnjSZCKs3jg1ByH5Hbo2+0txm4/6tKn96kP6BPOK
/L+kuWiIv3ykSO7K38nZUQF3PLc0r1hoUe/JZlpVnys1m6RwAszIS4o4cBmqTGCWzoeLUOTZ7fZO
mknVwlPfbJwYFgwj9nl8irk2ZycE9v2uQOWvbLWD4n4kc0+kPn1n6GzHNzD4Nar34Jg8GHF8JtFv
tKJGvrqnD5BKZPRU32N21iDccK2b+h+7nxVxfV5BY/egiiYTBlS7sC5jZdtbpCoIdSinJBGSdE1n
8xFEKmClVl/bGZTiXM6iTSbPCqXIeXAS/SMpfcYZke4Lmt0YdCf3tFkTpf/LY65yov8iXNDlefOS
We0m1pTbGXfcQlTFHYcKLqlkuRPugOaSvnN27FnAam8Fd5DyCgGUrN0GEAtuU0YzUO15cUlNsRRn
rs786HZ+HZ3La6T7TXdGA3jigVnoIeTfH3yI6xaEugCEx+p0VDc/3EdvsyclSQu1bSmMrEx3cPuj
Eve8zVA8ryE+frnGF9Tcq9JqsVh8JNgDonipFUkX64FK3NnTrJIzQqx01eqYjUd3VgTKvyuojQS3
qcmvLQKTzpmq3GtlsuBZklyPS/wyYxnU8uDUE4XCJA+3icSdX36mPluFSMl6anOjDlQ8xxAOAKeP
eKpIhmZpb00a9JcVkL2OoTB7DoZOhPFpMby3GpSSZD+IxOORFOIAy68bhZGaOUC3yl/LGu+rH4Se
zgFa6Uu++W0tnVC2FEsUHMJgLFOO2o5jtOggbt7w4YKtdROHqDknO2DqljXc1pEQMhIHHr0RS2g9
z6OrXhjC3mPM6SdG//dD87I9/Ee3Fk2UI4o+HVx+FRjKkI3J/2hNmshNwoRHs2B+4DUbgmp3/iMN
JhASXh2LcBI086JA5u4kLABOSoa5gQ5hLnlczFsra4YQJuOr9x1M327dziCQQ02wZai4Pcg8L4Zk
tmsPPS/dcWprJ9qEXqV5Y9S6ZfuqkjGmiV+PivfG2Bnzsn13k5mdU3ArkgLtv+7IdazBnt85onpR
UcJ1RvJne0jhtNHu3rRa7eoJwZQtahBm4jBbRoQGuquvxHZ+EZEkLRhaPye6brztLn4+lDGWu70J
jmRl59i1Z9B9WxwjOGQx2xjq/2bIVigrAoQHpNN6COUtNCNENArcRInNM1LmFWOt/+g+bP+WgVEa
Bvy/Yu9yvj/MLZgnnB/ErrNM/v35hCQ9XgF0fz7AHIIPaGUSEKgcIVbxJxYOH0t07y5rDOynrMpu
0xR2aVP4tv5KnJtu2r8H6oAihM/tHqDeE5rCI0geuul+LxEkWOJo68PZHFxqHmaGnWAV2zBaX/Hg
WXAUvrmByY5tHdQrRgjcGfWIe1GDRnaJT0SHJWZjxDGGHT74KQkoyuEGypinCU6SC4ElIaIPr6PB
vDg3hcVB+dxjFqr7H2YNB0LB4ypr1qv/lhtWqIj0p8nsNYVMrWAdSEO9JqCFdF5rD+HoOJao3Ze2
5DWnRxfDZGEOcQdD9XBt3ENmDH/N6vmJ6Jd1b+eDyb5igaqQ5izJTmZxvw9bomoOP29+X7F91glA
CHbfGeL6gN6+qBpl9aD3nQFnfU/PqBucGEoomWXEDo7jFAhskH0dxHLbOeeyYrbvPPsXZp82AQbF
0SoqbHSSErZ18aqMm5cmKr5qLWkmh6BnTjHLcfiN9zva3P6Koe1/EqM4ymkTJU/+go2tCNaJwUsO
fmkdV23xFAmeGtwN8iY6vwvpVU3U/zNcZhGC+wswJemvl3PXPvE36wx6QMipuQIuCxBW+a1ZHvid
iJ5zqaXKZZ2KirI20pzU+CbX/8jj89sV3boKWq9WwUqfnUDHnK/2bCMaEYWmokLvcubA6ipbXyoy
k/MKsUu4uPIRzhljKvtjq/MrzM/3ax5qWy6yIWJZOgUtXfrmOtZ7fQBail6svoIkr0KDO/frzgL+
zgWnRUWMTApk5D/fBDTpdyMR1SeR/sLgueJcVt4fk5ZUwNpZvUeLZZREsC4zbWsmbnIcspRbFT11
T1SCOOAphopt9OJZ59xkxkqIRBMtmJ8ygg9fE4iIEKmI93ZjAucIMi7bABey6YMdoaBWeZrltAIs
bzLggpCnXMzSAhh0yegRxrwGZTEnSkoMZWzFuvEDU+MaeWl5sU6/FMxBMkrXwhu5IZ4PTvCu+GWk
WretShDBIsHHiEwx2mH39CqAYeA1iZjvOxLfTL4tjKVb5pj9wTkk2xgQEoChruAaL8/ZD+G/w8s6
ieZCync0ETri/kgSO17deFjlj37AJEbvfRl0An6kVg0WuZSCXyqLoam7obISGRpCLTTciG3HB3be
0KwwIdZ0wGzH9MS+IUNFmhcI5PbemuQxFwUZMltD+L5fsVsOMs6eK3UoWR0c28B/4gRiGl3QjFJI
La8Gurt7UDg1y1SHCMfSff4fDY6SyCtthLw+iJumtM/3GBG8ERIifOT3/tBMA168Xir1pwzNp9NZ
7I6e5cMUeQqc5jAxfVCr6FETjIXVEZbZR8bwvndhcIul8TSwBdLX/km8QGT594SLKAtLqrC3iZ+h
mbqbInAzQ1OtOAuk9qD3Jd0tVGv4XrHPXRMMzbTK9ikGwG6wb5K3O4pD8IFhnv+qhmeOA00XodCo
mD0c+7S+babxEcUx0zlZo2HdTdTt0t7l19HBrJEKigrYJSmKxmx9qiefcFZMnIcwwwo5D94WhuVd
KGfbTlxs9Pec4OAX2Bv5Dx3CndN3OQYu73QlthWQYv/9YrdzDSIqHB2P/qWk2cOczkOzGfBnobut
YPck0YTqOGdhbaPB/SaislUGBnzw+rTWxc26SRoFG54q2C6q38PC7ipRA7t+28f299jMkZsoTGKc
mnII55UOOWgBkO/sLH1XQFT/NqJINWOQcW2+4t/0YvGn1+3GO3hjN+iwjwuzWK/nwFR44sGP8v84
yaj9SnKXa/Y+6KkijSpzTMTchtiDUA2fpMs38S7OnvE6zwnEUT8bDMhuJW/EKuHei8U3sG+A++vZ
jjJuu+8bm/fZjTUuJg4p5SXCYJKIRRvSijW5Y94QH4udC0/MGqs2LknQ373ziFrHOPe/3O1acaOj
oLQS2oS7PXPpS+Jkjp4cMLAwR3soIA3mUDCqZHX57RNAace8/ra9+C9/uoS2FqGxknkg3NtSeAKr
+07MNAHym7cfLlkOHZ+YDKgCTZCnFhaft1Y4IRJwkvQHx8Jy6i7QYUynMcrYkBYVypizcKH+Crwc
KrEHXEZwF/y273z+whglb8yCuW5a8/DRzVfWs1TB6jnR4rNg1XYYgToQXwYrL92Wgn8z07J2inmt
38yfOB/cXzmdzEp8AoV6hKk3IlAHdHswMrMGU/j0LIPIubMVMIpvkTW1Nhe32sgqTJEGF++AZBAA
paWMvrNH2ELj5iV4NJUwD3CSEj7clUgR1kUb5hIZhNssGl0ufjndiqN9wEA7mf8M90a+fzbXsqyv
Lj2uCXArlPdS7+zTC7gNvYRQctPbSWDUrjG5SvTExfMURDW9XC0BMGrKLjIuPbwDkmntidF2fnJm
TX5Y1bBZLRsmZt67bXncfS+jQxYoGTBrWAaj/ZB1I5aveKzC/KgQDSO4zYM2GDVdx3Qm0AoAk34Y
WGiqlU6Y7PKgUCwHLbo0QQpb+wTfdQaOGreGMux+tnNgdNAnyD0KtkShC6cDCnBPmM5iBIYdm8vL
OIDUFjFRNwuytDP7+JzgOdC8jQaRyvv9V/QK42+93b4NSCwk3xtTgq0z3qV7xhYR1JGvfMPmDIW9
3KfRmW6DEzviGAn5Anu4vO2tcrNnCf5RDYHZE6L9/DyQDYVMPX2HcFd+Hu1OF49BE0t+CcV5LgE+
0KZhtm8iZayR9mHhIh4u8FhzuXLIVHSKQwOQmSL6uU6Px2uvZl1aMULqPxRDEDjzL8l+hA95R6Jn
9/NTVvEV3KPqCP4PM/PgCXrK2Al3KXwvX68KW2ZlZnVn1CWEgxFLk53VkbA+1xRgqN47T8G6s8v5
vy7esUn/lktCGXVuWBRQ4dI5nAXKdyg9XvVAb1tmSDt79q0zSMEz/QMfQHBJ9/sQ6K0XrHLGGYu4
HJ/9UkrMxbauOxdr5znHjS035OqUpHxE5ApEf1fs2jsO2mqqDnxV6t2kj9nbIRFgozNSsyrbi0Hj
IXPTcSs8EDqQ7x/5lToOgAEyDNN9QG0zj9wfS+XVRH5gGJfyJxlw0TsOrLLVHWjA2z++3qDMIxXs
iQrsjDAuk4bnDYyeptO7c2IJO50kRmrJy074isGAkwXL6uaSxj/80S5w2GZ2ZkpPyF+pLjxEJi9L
iBv/pvhzqc5PeDQoCE9Iv2PaY+8lO19Mzvj2DYgf+TLjv/iRrt0uRMIt3UwoK7hwit/JqesVwt5x
wO6B1JmvhlwHNDaP9ZSsgIeGFtZTNWHjziVn5U+Q4b2QQT/2aYXwwaooHWblp2tGqp/uutN+8QWF
X25DWPFlpIwDY2QS99Pp0paYHiLF98pPGEhHZSiB6nVLAuwlt3+ABKrLJFQU4cY3Q0NbDsZZ7EvN
/FEIftw+KA0QlmRDZ1UjvVgWWtzYi2NiWfXeDMJnFk56M1Dqy5EwwdQ43kSDyuLFZWs7Bnpvoy4H
f0jQCzsrJDFB7ejoCayjwejq4n2ElFJGL7NifFHV3lafH4uce4hQF/4Zux0D0utV0e2PqDAEtstO
91egQHTK7w3o5NvwdkT+56rM523z3pw1CU99TZ7w8Z/Ti7BgnxlhWmKYZJRBcNtf9GtUr1ID5tlV
EmdTFdVzvYT44caisf6G8uacUQG70CAkLOedC3GkUUpjsQNiMb8NcUwoH+5dE3i7Xbunr/Gg3yM9
2hEffDROHD7MomSvoEdDqF+Dxu99JkOkwcekNdNjeHZb/etM3SEJoWtdINjlO4c5xXsQ18WDDctU
yz2ytAksMu2Nhnq8J4pSA5nJNjSuAtFvJXNmFxa9FoRJhVsvz9dQSOwLRY+Q02FKQ1kQkN6VhFqj
JVjQw10N5xvGOtYwpvhYVv4T70OdtniCczQWJzR1OkTfYJlKwgNNkGMILY9aPdn6kJIxRkUUh40c
M0dJgaP+rlPNmEuDOZsc934bXe6ATdCAM5i4gXKqRGylheS0h3QcRqoKeKVxyLvhaAc8OFAr3cXE
nK2O2iNw7VTAifGQeL/d1/gXrBxdqBtuOBg5Db+WF/UDEEWvtjceqawZs3awvtxUM/KhuZxUZ1vF
g9DYrDJzZ/dptz+WHZjmFbdu7RhWMSj1iGE1E8PtUfZJrkoibwbeX5orYDI6pXqTai0pPFobqNAh
RpMi60B/NfPmwRYymzUTNe9Q6CwIjnoWocoE5IG57DLjRewlNxmvicYBs8SpyXHWixVjiWx+CgRZ
hDHFUWABgN84Y2HeAFitiqoqKBRtU075iOA+T1leBqYWz5LHLI8oMnZ/FdW813RM3HRXgztzb0oG
vIQuxPuO4zT9A0JpgizTzhdN2INGLDdwWCr5pRqy0cQ6s46NFlC24nwpbD0WQcVLMHJGNFpMFaOH
mxcoI6up7GJK7GyHi3WHkpPj6C5NASB8Qu/rr9W1aNcVva8EYcuY0SJYvAh8T974Uq5FoxVs3MTw
4NS+zBaT093iyaqN4xuVxEJh4x6qm0weFGFeb1yjh4L/HFCFP5W6KNknIbQ8WY73Ss3zDjBoTt3Y
3SPuwkVU4trIDSoEirpwvNfmb13z3cl/4zYLKYXI1uwObVTuXtn7f3a0hYijvEwhS2k7fvWmHxtx
3XHWBweEXX9uZ7Su0BevnrqtnHjXS2lb+ZlLlfiKLBsDB+yrSTllC0Oal63jfDqPS50lEfLslo3U
bz1t38yvy+foiPh/cLD5ok9pYeRv6qijS9GMYvVfbL9OAgohFoncUWRCoVrXmAWu+4/VL+glQdzW
3DShUlbxzdw4LFbYeTKYx4tEtz01MSXC8+2+UzGVQAM6k+HpM4ThGqVshfjaMDDuMfNpDxv9TXel
IiDzPdu8n/uAlABx+YB2lTIKswqaA9FWkaN2ktqItV/YXChzOyWgcxQriuEkjXrJIIFBNcugk2Wa
AP241FnNXVPb7d9yLFD+tO1wYjOFCj7dDHulq3EspKK5ByL/IfwkNzspYGIqdDraZSNZInHlt/Ru
Vi6KaLFPSSi/HGbO3+OLJHy/Y9/GFAftaHORS5tYJwwLsKfPMgEXMdjtLrUapAMDkL3GIJ+7WSqk
x9PhVJ2muwmmOG8WWS/CdgBaT8V1KahmHc1IfHewm95jxlK3YeqeKewWOM8+IiBVj15GtBhWcKtc
d+/dyv1cHyms1hA9E4m85AhvWKznPCW3epGzXtkH3SX2rdo7cyrd/x98zTb/dT2IsE25iSK54Rup
7Z1+6iBOltehuJTMHsseY2L9MQFYNhxa57o8w+5wYpOE1OkpsopHNN0P5xfUgqZ0HOmaejBb4fWU
QDK/SKrRsBR32hLXxA8kkRhTViFyJhbH0Mn6LZWFIlafOSXTioTcpYq2QijZXJ25HRvS36CkgiUJ
XkFWPCkAK9BSw7T36IaLr3Zs6XshC162tK9yTDX6bdRg2qkWx61APOTq3Ev5kkG6mfVlQlLwzsrf
4/F+bsQT+BJPtmFLW7ETB7wqcTfRqAb+QHXzMU+V1ji0jNqHz0eGPC+5uLS20EZqeD7B4tkvzWg3
B//Poh488aRJVLIBBDSRv+FUlsHZJ90y7Mh96dTsH0XoBWVyVDq057vYS8HVrrJi5lL2KMvhGlJH
r9wkQKeQ3+/y1YYD2Ht3N5/vqOVkkxbBdCsCj+64GN9ufZ4CBLMsxHKWIwHDBOtZA5h04xk1NrTh
uYqWTfO6jpEpx/GFC7Y7JAVXr+IbYPyl4iIJ4tMAuLX2mnW+FOH8BReWjiol3GenCo7YPX52G6i8
Cp2g7IsPZjvX0CH5BUTBheSA5L4SEQaPvLYDJ88n9PH/S5b3LOE6qC4EfrAKNWHUWot9EzDlt5bw
m+aDDPq5VZ3QnAcrEhdBA9ZnyUpYHlkOB/4eTd4ydKoVYaSq0Ax/GGGJAUpXeq6oQXUluTbDtY7H
OEUM9x9xQwvUv9szJsGd0+ytTrlBXjaOA9baemdTQJHqZuhvvnTcIxLSZ9KaRvRL42MqA8akoy79
eGUaupP2qhKUbzyMmX0D/roF5xqsaVPTll7PkKquTyb3wzpbnwmFm5pYGoe7E6BvPQ+JAYC+Hatf
8MDuokr/TzrPO7+0mTDk0mxE+CcODus9UuMT0l+f37nzwSKy8tTv8Zs7hdAVJJ0bXfVaXBp9rvBx
CY93slsA2uh2Av/E59LFnB3zdinfB94KDPBfr1MDeJLWxOMXVSdxlRKM/NusT0cETf+1ShPWroxt
wqDQgR7b1xAkRLWpnUTFugJ1Z/J+OV8LveEu8ZBxIV6qngiLdmQniyxv80awX2AXY3bfSJ8hyK4F
LFvgyMG4J+5eP/FMO4xVgTBxorEuV1CJuYKlVwernzWZRyhpcnAr8w9XPyIUowP1LP3MHZsFxlPb
d9bV99ZnHw2WLPVvgcS6tlfBaXfNXVo2PhKXAwriF4ThXRbqVCMW5HybCnvuvCT2yyhbBvnpSkYN
yfOROKzLHgn7DY1jzTK9gSjseZqwD9UwDbVn8skvrY1eQRAAZxFBS5Gkpfqm5TqVkCEWs9bDRIgw
zL4vrRQlNSxhOo5+sax2pFyC9jxPmiyU1asfIxksoQcyS1XGF3o/M7sbOZ5zzePpFPQf/FBDAhLJ
3gNCEYcEhHzrN3Uel92naSODxubQ19rzOLhtfqdlACJtA/B5zUoqF9kgXOSCvFsJpYjUWH/gNRiE
Y/cQBonlAbDi0hhjZ0DkaHMDE9/nJiz3DPQUnZ2JQ1nMRadlrCytrgpioQnA7jSPJdzXWzUfuZ6/
ogUhvl4TvIOydMoQ2U4T/yLcdkogVc2eojxkPkqvLt3QAL4pb97NKeUv/kdO/O2xj54WxHRTFf52
7yC52cPy8mIfZp+vhVy2YcmiYeRW8xK/q7e34bFmkQ3n22Az55zY2yC5QdxhbeVIxl3lJ5ygc7+0
nI6zVlFitPG3uNbolF3TMRpqI/MjtcJsGpabtdY9C2mxLJPfWu3e1IR9YVOrsoXxGHLZQZ359nrv
9vbFaqmXKKvneiEp703QiN3rTyYpCpo/Jv0p3qmB4GFgS8ikF6lu66hFP4HrPIw6gjM2gdK2Cj3q
sDpGdtzskLtSMgU48wy6IOkPJFT7o2vwqznMZ073GZn8onmeTyhVYr8OkxLgu8XJXPzDnoxfs5Lc
I+1MjYIrt3spIercqR5UU3qjmxBXVkXapsWKV64zlAwuA16Nc4erVpLHskEuh7FRZYryQy3HQMja
yHa2PxrmO6JNZ8FvWHpp6QyRwOw6pT6bhOoqRixb5ayyCx2iAIC+i/EKFmlRFW8oofupvlxQwBlS
D5Vw9X0el9nI396BXWS02jZC1dbxlDiAGDB+NsptQBq3NBja2NAd2RfcwsNqo4VDtoDnt7PHhWO3
WJKhwSr3byPva6V7GwsUbYcC/pb9TFJpdpL7kVvFVz5EBZvItpHI2c1EHmZKUykkmkyD1Gi/gy3X
+zZDD6EO50YaulKTyX66PVm62sPWhoOUR63V7gY6WJWRGRWdKFMEGmaNN82Ny8Keu37ezPOInkAU
K+p7wG3USUcpRDP29oaZa/wBnyTMsujmJK9CBLj4b01DMLEtwxOamtoVydgcfXSDnAoWAEfmbV7X
InR3csCsXOQP2W20sNkl2sL6sacZB6txnc2nJKWJvopxJzIXCqlBRtY1MYS3t352FBlqnajyVlon
JLZw49Cjq8+tu1JREM+/RHMFqjc9xl1mMuugxM5ziusoZvkOhVHrQGrpEe9iiwqSuV1WJUv3dh3b
wBR1RqhmIycGG7G3/xapOjWdXe72VZmFwjZ6nW4Z6KDCuWMSDglyR+aT546xKa6aIwrL347fDjtx
zvQvJUBmHi7NjU2BiYUViUudmeHIwCay8AJVyqfdXM0AG6AW4H5WbDcEi5DkkkIWzvqFcgv7Smme
ykqmPEfHJtal1zREtz82TeDa7m1WyxQidffyNVx4+x4/zB5646eWk6C3gLZclqZkTvKNC8KWjKZ2
z46CD5bkgiRMeiZObXy9hTgZcn5gRaJ2JFQ9nzK4l2bqjbeRYu6yIbAUqS5M8OSLwqjNy6XD6ac7
+/tqpUwFvNSQmAZKShx89lX8DHy+0vlIOcqBHUeRHAJReftszKwch5D+2Kk+oFQ0WAT8/rXTYJnf
5v8/SXA4jW9B1Fdxtjmmw/ZljV7xNeRoMWXUSRkB8/e55bocfsOtzHPI8AvC6/xgn9nCZKKlfU2C
i4NDbGfpNm7YDjOfCgEO0TnSIBeYEyC1cyIrf2bXvcoTxI05/yrKh2lz/dUa+cPrtrbkOwgDva1o
gcgV4wKavxRg9nchpC/jkb1Adc7noYQNGXhFoJBTnUR/v+z9UCYrfMbRw0Movp8gzKBtoy7Cbzzo
XowDn+jrxPtf6PGCbpMfwki0olB1sAa9BSyVoAx0uUSIz0mL/2bK6cGJIqup3p0ye9wkOfVzpxTU
9Dy7Mq3QiJ+tgQOy6vKRE6jau/qGTwDuf3wfDI/+3EESnY6t98E/2K2ZCYUuFj8RppgwWx/JDV2V
mhub+wTh3YD/qbJV/7UsyNIS2XWN0HWI4fo9IX2EoIm3Uh9NlnurRGvBI4NVR4MkhfU2m060bty7
b7JbyJBnKD9TkDmH1dYZiOf0rusDhgX+xJuRJbxTzhATwtB9NQwaPlnnWc2tYqcTPM3x1bc6ioF/
Hzx4KMPllR5Beie8Zp3bpCoN+fsIkEeTiFnOl8mYzJkVUV1nXgSpqsjfRuGhxdXhhNIsVM4LODsM
NiG3ITtWbpbJQiPUgl5CmB/H6gjKbvUCVKKH8Er0aP3/nZzNevtfrSjQJP39sKq8tWQg7/dc6+tJ
3hY/YL7nEKnBAsW8fVbgkG685ioyfIYrChtqusDOmfjhkTjHluzeSxTZquZ+hQgDbWKPYaVmw41m
4vNXBZTOnKyDjToVrC6kfG1M6baLEugP2wWdT+E9ef1ii9WbhQ3m9i74Ta6/s/01pQkTlgRFqV1y
h61aylann4SoaXr7+Mbu20Q3iPDeEwJ+bt+u/zj0kI98JN18vZWaoeguRaj78ZWfCAQiBkmVqFGL
gm4fPWRIjuXGrsiOuXBAfNzhFvSrq/vo8OvK03a0F1759jNXA5sdWuFppFJlOI8fnsUl64ZHsBEv
4umhR7JL9rwJLhHfYoJ4iA65SPkBckgD7IlRKLAGDKUSSFQQQD19SSj+MV4NvyaEfRSjV4FihX4U
YIC2ra2JDGF6rDIPCvoPO0p7S2xNEj0ptCG066+wE/LvF0WokmxWm9EGFXvraZ10ohBoik+sTbnF
qiCWlLFXd5GwvG9xr2th9LHuF49Gj1hpPrN3f5drkouJ82wEbG4HFsNRaL5H6jiVuiU4pI0nE3yL
xkCNa5hH/QF6E7HUDv9xdzHBNMiuKBOLZNVDP+grgqr7V/zk21hmrPx8IVYyJ5uRq4T9bSANMA9q
Uz5/sP42KF7XDL8D/YEeIsc7v9KX5McBjh2oWBZfvem4W7b+hyU+JFdD8bUk/SIVzHbEA3J7pEPh
TeJNhBtmIaggzmwqsnoUZglWPICBT3L/U5XOJv4X6KfqJv9InmMSZEtS4sJzPexGeStgjS7ga1uS
xCeaApyRHT0MYA4ukPTLD9BhJkWlq21xXIMkFBQJApGgLH0cgq08NszBhyvtrEHsNr/V9xHRcvpR
Bk4Bk0XCJMDmLv3WlSLRoc7IQElafSpV9Y2/4MaofJiuUPeZYqGlXhNXphzEUbwNKl7F6KPrDekX
Z+io0xZO34QWCRh0ax9FqdXK7kwYVS4LRPteUsodRx3bwt4qgsKTV4Poc8PTxQx4dbj/efLIOxm7
77yEH4VSiGup1lIwQH7g3L6VhP9wdjWmJwoiffn2p5RTE1GQ4rHvFvWUOGF4h5VD7I80cMb1BfEN
b7jMNZty6LmMLr3PjF1LZi5A8LVaDRoLkvedpVrxpm4G3lWJhhMCJQipQaGA+UsceQw1XQ2gJ4Wh
DmRpAxdKPofMlMqljMp8+82jBu+TAtTqO9N1/k5I74frENe2V/uPnrUsXlyZlBv8ZwK3p5OIyFdO
sMSJJjOKMBYAJEdBAoq6d0uPyviq05QcxwROF1VwAEpfxqiyCUEa1FTT/mX8Gekfs/JkwRkeHAne
T0c5fdT9w2yFavnvgb8ZPecU+0oABsIqycfu62YMTlB0ZU5t0/uQOsEF9kh1yPItIABQY8Jp6w0z
1VJRL3qwWJaf9cLlpewmICv664klD5yIcftSbO3zdD/LG86qyRloTng74B1WKBjvB8cJw6H6gJPw
UqZ5KCiFBogqlq1s1K9jBAR2E5UzUuhekTivGZ5qgul/TMAg7T/DmN/kZjksQdmZb0WYpy7u0yUs
7bbgv5/6ug1ox1eoJJLFOP8FvuLvGfNePS7Ajuk0P3WjAv1Ys3M7D37TmuDn0AXV4Ve0xjB7qXdd
G+YyzbFjADgD/biEdUO3AvG3VSLJOmkbqJXG3dkTdJjHbGk/sWFMP0lzbaYEtZqBvBz86gtxhvbY
KxjaStIE3ZZ1WpZgZQYrsaKSKKvkORqnPmsIfG3Q6a6I9NgE8lZnzQ8nx1JNJgJ8BGN5AFpRSTQf
Rz3eGWVQ6UKDSmZDxv5C0C9wd1qQCW1EUFHCIwy+0AL3iB+hqzbH5tBRdxaMchIT3WZvJ/ol8wTT
IfWHsxJF4y0/LD9PA+9h+XiLRemNe6dyjex6MmipRPyUTB1OFryYlOz4CS0k8Nt8vp2AcQX35lg8
xDTkvPXwL9cRgKh4qaJ0JYP+Aa2YOEvBXu1RDNPg0FTE4aPazntQdDTE2ZQtWuARkn3J5aHzIF+f
mWibYUJ07QZYbWbGKYeoZj6zWUUPcTlPsUIcW75K4qREKlLUnQ0BRx5S8svq5NYYOBVKzq2WKHZO
Pj811E1k+I3s+QoJps/No6tr9CwWhUgrZrgtFUunJ3CWEX+jzY3NjqAbCAkhXFwlpgIeV1Ne86P8
19nx755KGx9cMdoENuNPmlYvOzxoJQGfwapB1l8TCsRW9FzbwAXK/WO0YSP5JfJuE1hqex7PtXEC
QXQV59naYfxPoaNbsKzu9zWq8FDiIdsuyeFMFDR2OKzKuzRbZPe8xe+qIEABTmZb9YRhw1IWKaqH
hYF+ILGOI/cMgrjAPEFd5jWHVPm9mMY9GcFHP+QsiEp9aEDHxEoEAqbU60eXFKZnxJeVvs5B19T4
L58+DpJ5Swd2+RoDchim9JBYISs/wc+vCDRKUhEDBkPkiNdR4TR4dkYIj0pXr6PSBSY93HfyhnTx
B4kO2hoWOCssVQ5CY4nKxFLSt6Xn45wHnrKenQ5HGNZeJ6OKwpBsyQuNaw2yj4Vy+umRClj1I6ij
5+gCYg88LEdhgkz4/0jBCYFzp1dDeanQDG07Q5e7P+V4JQmjU1odXM9xETbHhuNAO2NetQSSrTY2
ArKikYWPtbg4ecWbEC7Ww0VhUGtMqTxhmSdwRs2fXHT6NnvmXjCYTxz5qrlrckwtBluA1Uru5oiO
u1wNq1Z5WFcSgI1RDlFxYz5YZohwo9H8WMK7rKSxSnaqV7iPEV+dCEKSngBvn4rDTHsoGMmnhI67
yTFr86K/m/7F447uMy2+QVlhjSzypoVxPri5u3e2DWqd+XJLllkbRjZvichbCtBEXOKZ7Mtn0BWF
wwoApYqF0VauaPAswdQdfQsEepOPKgWnW7vTBAAapK5PAcwafO0HNoe2iwy9daph0SAXfAnW9izH
PRGUsqiSFzRayGVTaZbuP+KKyMIqThEa560qFxZmWiRwjqaLYwzaGdbrn5A3AxErUlwDPhoMwL4K
dVBpavdMeQTVyzP1CcKztJjPTC4mWoQphPKzk74FAAFB9PQLMHYwGYDgWndFhr8Qirsn4f9gYD7e
u6HU76IruEhZAGkjbjyru6l+uCabhFAokKJCVpRwOszjAwbk90VHJsdvsSgWAhCfZsXTskQ9zms/
VCrbOYOWy/DF2H5+ak4DgwJd1zPEONn0li8LRkQrV/gVAEYHtK4JiDIwkUe/mwFP+FGlCFxR07rw
tHlHeqNJg5zd5z9TYLGE0xnXmEUh7WBa0Hgr67jIdiUI1gqrA+Kpu9jKSQgv2rVdqS3hX1w489vQ
AG9IrgrjdskitZzDG6JRaCq98xglP9857jhBkwAYOKNSxj6muQHyDxY6/ioqFP5PEaUa4Ko8CQlg
IvQmr964VCVCHgzpA4TVjZPEzZpGNpMxCjnL7q6DlLMDjMYjpkNsT4GVGg4w7cDCldr8DUZAqqc2
+FiPzAw/+v5Q1ppJY5ATw914c68R8lmqYtPmjTmky3oBU5XHZKG+7EvHaGokvtusXaoBQ1hRneC2
Ixkr01pOS5T9THpmDbh9r/NWxKKizkt5C30nVBzvP9Jv3vz0x4NLw24WHKv6JYAoyrsQpJnLpg1R
aymT6bH9paGScSS1+wX4qogGkwObHx5R9s9EBM6r15yRVbZuFqqSk0DkE8WCMXZEuULVEog+XBXl
AN9VQ34pYrH1QBrYGwEs1kXnfdrGkXcUUrEi335q2zlm7RnimZwueYHwHnGUcl7GF50P56+AyvO4
gJ+lgoqQ+UwMgrsDuBNAIr+PDFqUSMegOxd08bO0fuCgiXGPfwQ07w93TH/KOOePUf58nDDHXef/
Ym+gEBOJx+JfCQV/X2AvegsRxEtXKQtmts0wfyiu9yXgjCpMWLP/nSFcg2+NRJBAxbtwHz9woTKf
LUJnOjLmTzuP/f0AHliBe3g/zxzjzEbSWPMxa3DHClcAqKHusuSfmCA2qRA9JD48Hr5wpg+YCaqf
GAafEsVicf4862BZ+0OoCrtK9ozoZB0R8E3BcmKP5jdB+YpM3U1+PFt70aXsaZ+c5UYvAVV7xanA
KbvvxLxvtRIieuaWEcmTScyElfgx0wk4rIBiK/9prN3orVtJ3JgEOo1i2HQbN0WjREyb40oOlsOh
0ImtrYDY2uwIX3nu7XckT0PHLf9ytA2spKohS8lkPjgy6u8uIbuOYJp1SdXtMnQCkmRLmDegvXjV
G+KG34B+h+qMBkl05tU3f2VBxySlhMLZrLmyo7w2Wbu5V8hQWKKViVHlVwOhbdqxbCCmK10PxhND
w214vPX0DC4snmlcS3eszmnvKGDPVGu9N4OYh+iOjtwiZwnJ0Xtt14u/jo2cqK5IL1l3NHjsUR0b
+pgj88bNunJjSPDERZnP4LnW7ictPXlbHVTwuW3DF+A0nZTdRBQuew+kSYPt73/P2DSzegW6+w0a
T5ML7zNGjEXSRGDs10zFOaAl2XB2EHSkrvX69sSkO+Py0KH0H8SWJrYVXDuM6Kv4lmB6uhXGSwH+
gaqirUkB6XGEX5E3GecYXRs5BmNqqVl4dBrDylcuevBKuIx/GknWBwrvPP2cdy+F7cITPr54twnn
1unLTFYmr/6XAf0gu9xuKBDAyX9c70yxPEi0fxahMbGsD7QnE3ox2mTccsLMKOMZ13BaMHnd6h9H
W4JiqQLqKaLUPb31YlYVq1kgAvNGTYxdxnZ9GAkRYsNJQCR78jDnXLEO2jCLJKnyN5HUBk6oNGHM
txIl3cLDphTeKNG+3dj1SJlw8lWn9ZVPIpE4ssPJZpvipyUW/FKdPBS10Pz+VfGt6ZQ5clTTKGuk
54KOC5R1rDCHKeMcjv2sylR4lIweJvqIM7GgS1OxEtBsnTQlQlN28zbL3Zd716ZPDAU1WLZ4jN6t
lljAKCRX0sT65eyHN6ek05wxFK9zrpI1taVqC9yXw+Hj5pUJCXnF+H7QWYmwXEwTD2ZOCd7nD8X1
2uf3FA+X36NccbreF2HaJP0eCPh5cxTpkwEfw9W2E3VhkAKywpy4Aya6qr1CbLKbaqHL4PQA/RMP
Ktl9YFz+14xnnr2BIEvioOWhj4Z9eSCpPVgJFlzkY6eZxXxjebP+nnVEw01+Sbes2ubDjNgNuNpI
wdWoh2WMxaUYukjxnYp+Ec8rFhsXlkY/o/W6UV/5Quk1X91LJSIoXAkfILteGetpeCSyfHicF8M6
WQa/wiKVgk+DYPXxe+nPFD3vxFQZ4qgLYK45euJO1Ijold3aWoRK8VZPI492QlJiDJm/n1PrrMo9
WqB6EhdKTF9gn+xdUdIGoSC1VaO0TsAAfx30gYNrYsZ7h+Gh7CoaiW94JYFMMko7DnuV04lVHPwf
40ZYDM2J9Au+yNNl8fjdcX7nS1DRcVKc6wliblOgVNZnpv4f7lyDzglYrkZY4VNmdFc++7iQG8di
jjqMVOQNmlWII8r+EEZbqZ73t1ZZtjpATbgOWmaaUCaJ/7jUsXBXiaTTbNGQqe/NRXYfTS8KXKWq
5PX3fIwA3oEtY2S9f1cP9djmVTt1dQqbDyoD9YcRRVPMiUQXoBovskMA/lFPca4j2hFY5u6T5sPk
rbnr+O8Sjj85VcAM2GKRvH+kQ7/1iXaiDGZOyNBgcoVAUbiA6eUvLQeH3/n1xcx7RPSxHIPr9mLe
YxA8vpWZePdxrns5AEGtSqH821XHbcqjfeIxzd5KLg+hyLFihCYNk06QhCqVMWglhMv2wz7rmyzl
Aj6x6eYqd5UM5OMxOxWrOrJH/mKu7Y/X62F9XhJEkFdYTAnQ/Brkl50U/A5Jqj/tZcMRU1aO9x4/
L2yZaQ/fdb5Nz4cLiESS6NxacAA0CloNo/FfSoVipc0vrj/Rp65c8/vuSztM5Mu78iV2tozfT0Qc
vjB9Nm5RZdM7+eF3C2NLRpK1XZ5e2u5OazdoYv6Sbc5fBCx3pexWVnkQaRj94E0pjGPwnGHNHMjx
1KIhVDywVmDryy3V4OYjVFgoaNFYZXErozPnOpM7k7/3bAAXRKc/Tv41VFoL59Jl5G+U/27slfYI
RFUCfT/2/KuTLJXGwDfqxTFFyu0upQi3NOD2bB02LqWcUYe0fs3dOJzrYggKeAFMW3bnIFD60UZ0
XaaOEG88mgx2jrp0DBWe8EZl5kumyLiFPgJqbf/xoFyYSKVi3Maz+JWxzCmFjm3Vx3sgb6mkNGHY
0QEqq1qR34us/WyL9ZQNuYrPhLIgtx0mifubtneIrXk2Mp23xdp/QiH05yYDTZn9Tfj2Iw75IJtE
oCVmqDi0Xsre3pWiJDvSNJMdX5iOgFMVd223HnzSIZn+qRiZmEZVgb/BSA1zEHjDNvXyUqM94AwE
8XZVHTTPStUnjkMc8tYdoTDIe7iyQvKmlUrgc4Il6ZFhWz1Av0C1nNpk0ldb6KvtsSWIhUFIC07c
QBLU6U0h0sxRoOdP1o0ShdJ8NGq3F2nm8yc9oQ2wFJpDUek5zONRwp5+na88rdT8Z31Q8vVVX3Lp
03f31ytFrda1iSThlARFQ2ob8M8iyQLl22FsrC3p7K4T4MJWfLI1NoQZbTVcVEqlwNwzqG4AkdRf
Ag+05bUXcwneCH1H9/NH5FP6RMVBtcUia3F+XD15mfzrMgxIFiXiL/2fFayBmYuw9bIy4LiOHoOM
0ynAGBC8g/EG+hIVlOxsAvIVYImLiXAqCX6E+ka57zdXwPl6duDimQC9bfrrf+mHCsXW/cW1B5pU
ZVZI5Zps9kHPBcd81WIZ82VwQmvyYJEEhNkUitnfcqNv/8dX+UWEX5q3FcpAsueh9gy2DOjdz/I3
X2J0tQKrLfFZS68a2QfTQV4WQcJpXlyySFm8vRBUsYGwX/VDjizybgVudhYk+i28MqPLsG9mCjCq
ssg5u1OrhhsiOQr/P/c9O3wSjYdDB4qX78aBAsF1Itbye/dmno4gfrLKXZtMLgGBuLqZ+Xy0nck6
B2FMQDdf7jy11FYxotUKcKcTcrGI6U8MRUPUu2GoeUxuIQF2AcLKBsTXEAxaBy3EHKZZqzS7QQMQ
lJp1CgJwr7PEDX42PFZxzR8Icq1ofV0WWkLZ6ZD8pRSqazTzuesSnNaqg0c+80UnQSD2ie7UZZbX
9Nt1tR6Usq/aqqvSy4SiNX0rSsMGcsuQXRSuf60OlRVR59udDQm+qnYE5a1Qxqm+kZGBQaKzgYTV
4xjDczeImGI6QPDhsMBnVQjjnJuTQmeyHe5jCpFdCaycPYyADM/aKrwfSTMbXMRWJtXC27cYSaVG
IsfAAosKaAR+T4cmKZlO4dPtRqA7JchGGw1Eq0HaIDzfeS3T6YF3paxaypw/TZOzkmQksjaVp41f
VttOFd7qrjdW89Xba5qSVnaYSAbK3PocTfYR8Aq6tB1hZDLmfd9QpIS7L4CRMqW/PDblk6dkr41X
kc9JqeZsvPttHSYKpRR93ONHMpmLZWd8ddJCafNh0Qg11NUosiXu2n+yfUi3L9w/ywoeGnRVm8Xh
OcGsBLYNC/Eu4pPMVjExf52uAdKFW++nJRlMXUUsvN1nkOm/m2O5gNp7rVYO+HawmC+4uq/rElHu
u4i0jFQHiXxdVeeKvgxTMFrFLoy1rDNFdD3+ESycJM3tdiA4h+lzMfJA03lvYjOLpr0ugZ2PzyZP
eBShqn00aUGyWK5luFXH9SvLau2oExbn3yRN8tOzye8u5l8JB4sXs0SURUg378xxVXOcP1hqkSne
19F/0f4k5Z5c42BlmnaxjRSGzr1u0NkmJNCATspvVx7BmFMDQKJaUrjsKLo0XU/CWoXWQbJaVGan
b3Jdj1zDqX9jEk1guiFCJsUjT1Xx9HJaalyuR7jMIgpp77sqbu2vnnmM7u3yNR5vVqUGu+1sJR1w
JufVtQ7hFqbNAQoGX9Ws3ePaGE09V28hAgyIL2SXaxjpPcsSwuk99TcqTd/+bbfKMPa2Ae1Y6Dli
1mXFAlcjAsjgh4xkIIVGdS30gIFHuhLmT7uvjVtaEyjE5J/Cc5tqplj5WJ+VSBOnXua4wX48pP2G
hsHcy1ZPGpniNCymh9+0A3vCEmeLgoLHo2leC5J10dQDRzTbjGsEHmsROBj8rGEoBOXFZDQkEXB0
q3iwx3yeGffYQ1AQI710Z7Khs59GIIeARBb1QxA/Ri+SGyUiOoqdHA3FHrTfH7qxbFZF228aoATO
i/BuZPi/gvr4tdxF4lyz0KZbXQYFY6CZgtnBEJ/1LAAPosmtr92bsNlHCJ7WmXbvXR61NjUwiiMO
Vn7lX/9v864TI4NyoaCDZHKRDu2bXFTvpvp7CtLcB0SDegz2bit03UDX2iZ+aT4Zmu5H1TTh+yp0
x7a9W57UlohBYClJyv+xH/WQTlFJdq/fKFLEl9aE8e/Ci8kqRfggRiIMxhkxfCz7a383aI2eg1GX
AfIqs+SDjzbt6REh4Hfiqp5s3g0NhwxD8OneYgrXYult7/xAmAVcQ/cw0DWTR4q8S1mVpFy6oZJ0
KE3UQi1E6GYWPxa6v1zGIKEUMa1/wGZLDldQib62C7+u+gRb8oF5mDGpI4vWN2kWrxL8GH3SgIpy
W5rAq8moriVK9P1Qs9qtot/CAa/iXo1O2ABLKbD7L66TGxMxmPJj7masZurQvI0zww1P/mv6ZGv4
Tzi/imzHLpV0BLf0KZkwkjW0smf7nPy02JS0g5Vk0IKonSNcF0yC5dGdj5Bro1Tl8jyvpV+ITXba
ZxmobOLeJmFnp3iz3ns9jz0AAqafLy5sJevikgIeMlBguVrcOY48DU3k4o0ad6hhMQ6ccXjnM+Vn
lxZ2fdXcXrnhxzqEjCg8oRhvhXsXyoLjotEVEKJftfHPgju83z7GpMKuIt2e8j6dLR1tXW704FS8
8Ah84rEinD3IvbJPFbtiRlwFI6XbqSLj+0RBELcdyXsfr6fJapsSoK0Az+bC8ZjcrIYOS6ybBDhO
5ia30ENTMeWPAy2h8anEbY9SjFdYXcvWyfNXDprQqBNU0m7EQ+SwUe9WqaIWIP9dDInFfp15QGjM
HWL/fJq4TH5TIUXx9bNQV2TcOEqycxMSS1zmsVBGALpIOXFcbJKyHWS6RsGlguuz5ptNuw5QaQiA
ccQd6gALArJIiuvilztpauAxJw5tyS3Sve6f++sYKWCTJXK3w1JQNgA6/RjazHlq6PX0o3o4G5DH
tj6tHeyib+yl6bBTc9qBWzCJNB+/KlsMQGejmYIYEb69RNRP2Ylat+QYr4NjeWJLZB1NuByrwvFd
UQdbosUKIbMDS2mX5yctea9fclWTLIIBgBO7JGuQb8PDYAUuliVzU3dqKICN6F0Zmi7pUGHsLBJb
r9D08WXBWkuY9KsqY8kkarfhxZcw4QSUtc/tFdfXD/N5GoaAAWA8fYVHuiOq19ttLoB/hSuudDTa
JakdaRnQxDLzlU/JSFolC+W90TzNjU6lIc96fLbSmGEFEHJa+iIZBfXOwIo+BhvlITs0STy46ia0
ixBpKvycqU4B1s3yfD6snInd6f7ynk1W1uoasoPOMHdrxw2PQnGdKOFPRLc81biSTMgdZxjdd6NF
3qd3XEi786zQOjTVMk39QkulnR9RCPsSs+sngb1ma8IJfqPsO3baM2mVCG+cXaHBV7gONxvDgRmt
OaUSVmZUXW9/m+1Ga0qtCMO7r/HYQgJ8xVtKHySNGn7bg8fJWpDZisuGiH0xfEyjecgJE1qxkVpW
0N4RMkjJdFb9ghAxTNCWkiOjIapoHBumI0TQYBg47eGrMs3yiw3oUG8CAongwTS4zccIza2mYm3D
dePblB8l+iSo5yvw72NTXtUo1MZ8QkzmwJ9EinJMgtoNB8WduWZyl3drTZGknxSm57MB6J+Zu/HZ
vnI/2J5brZfSiqdhUsjRd5aEmp9QrsPcNGxIEUPQPd+kc376+rCtUMcm8gQHFia5ntYn1CXwPpus
6z2HanmoBZ6YUHLz+nD6r8+EITb70xZ4r9Gu8RL/KH5TMcwknb7XYoKN3obapywKd4ViThzp4JSD
03tF9+fKUFIxxAACcx8tc1m3ZqMU1mUdC2lYjOZMAx6uFK0Mh+k+zyVMuiPKDvz+BvZJdj5e1nDU
VsFGu9HEErQXbi72LfT29GB+OT8e6HRMLTUjgc+69XjLgn4zpD0YPpGSE5DxskRSs8e0kRCSMCLq
anuvzQLB5aPy7iLT+CughOaLkw1pWL3R09RrPj6v4ujN38chkbA0MuFHMDY9Baj41aQNiZX5TVO7
ZfdbOqlbwMKrWGJoX3kT3kR67mm3R16FeIBHXNcriDmQl6eWGZSipKKZ2SRNwlZAbg/samMF75Q+
Y0mHWOO/14+05sVCddUzGoiJ+tKJcNNLKbq1EDhMh5N7K3llxW2Gk6jyL7dytG2RO9R5DRXObLpe
ElBSPU0GxGmdvZBf6c/n+YY86LLekvBLA2Xha4iG1IjZ2s0qKZ1j2kedcV1LjN0jFljwbm7MSayn
wROzdbLMEU6Pd9XOtgD+fmHyJStCq9RKLWpgPU1nrl0HDnaK6NOzOODvSNHcOk7D9uiRqJjKDlCE
oybxHVCa4ZM+4w7evWjstrf741viKLoG1e+03Ucg6ZYXfMToTekBfS8RNynpQFrd3x53icIOF3W8
kZ7zhVY05O+PdeBSwfpR/ct7u+vDWgLZWDErdtFK8L5VewMru4LgtdNlEt/3gBbOtwfuQJz7HzUn
5aVyTsnvdjecuhyvX9W4QyssXzydq0eHAs3YZLSPYL/NImTFSIjFUJVcK2h9UpDpftIRhiqk/hW/
i9LRSlz73vyM6clTdFdW9tVkROMW0f1XfyUFql1ZXiTBBKkR7cDSmP+AjZ+5Ecz6w3uNzKSaGIel
pWVYPJ+2U+vAxQUy10bySjmh0xmKuKMd0PLj56Wh34TJzcB8wnqvzxxJ1/QUwvh9e5YSj6yfz/Qb
008e2EFtonWSk3Vrm72h02mB0ALcK5tqFrkPzNOpgB/P+v/CD1NzsVXmuAWUVkcvK88e1vyujNY4
FExPpAZ5ZATmHwNI3IelS30v2WhzU9H8VZRXTcUHU1SMjE+wPVC35q8CxLR9NuG7kr8kuUVFZ2xV
D/kEWLFoiWetkk/tdKIXCBJyverm9pe7W9qi8xR3G6SKYVPd/xkwddu9r6JDp2vfEBhfNTXFRSkC
pgZcIHT+2p0oIZqPZ5LadINQ+x236zmSuguyAL3pppaUhYjXtp+D5QUu2w1VlMzN+F/Qf8eAbbzF
g3k8SjgInOWW4AV0y4Xee/xq94OA1aDHDQYSxqfwhHgo/0O4S/5CYuaufvfGNNsrz+TqopIU0ccH
2sQI8jzfpCafxptVeWGRLjYyFgcccG3/izy8q/f9nzBY3fLkZr3ixGFJdvwsmIvQM8BS4DcJB+K2
6MUgN3iFLMiLFDBlAqDCq5tlytxH0660JK56S2UVFTE/G8EtsmkdV/EIcvxshhAUUEIG4/KMcLvV
Yh6w6XVzTUOhfA78rwZdDvPQ9GhYDJSrC1ZBe4W0E3cyXfC2ujBBwRf+3VtYr448MonMxFaFMtwd
7PEGFkdYRffI8qEk4gwIvmaRWLp5b0mz3agXEY9ijmZdyBG1gFJufmAFyFaiI9vM6EIa8pnIrAR3
BAn5u4M1zh/y4IGxpWeQZ6icyF4Zdtnryj5m6l6+SFcfv9UxeQa0IfCtJfumAXD/iTMIWqB91y+z
iTeIsTyMX8J6QFoldxKOO4GWSle0WKBvI0cBrKdW93fUqK2WbOj/77kWR7Nss4FdPsAC4l6wTJ4r
/8yz/iXzKNlID0JD9ZrJGdVxWKEXTyJie6E/YGIwYSZKYnBytKDIqABDpQGquaVMFOJSNuJNRBgZ
mqym6stHMqyT+oiHN2j013a67che/wxCLkuBTUVz6L217b31/CTU9pjS55qzfhJ1vO/ltpmbbNEi
SMlukO2XCpoK5EIuxHBnqowpsw341zsfagsbWmf3SeK3LY/j9SzMcaxeileEohJjcYZ2hDPm8tas
4hdFtfCjQuh6D8IJAeaxt9zvQOH0SZ8NAvks9sSOxRUKdV3IcGglPRGVmay34nmoZ9EE7IvMXmDt
IC5S8hXOEvvwxDtSaNEdSC7ajStaykoQ5Uhfy7xjdEjqMPAayRnsBVgEgxdJXzSDJ2FOXEcbR3Ar
87ZggO8XI9RJA+tJQyL+71Ef/uaPNzeJ3nnoBW9gEyqYVQ/FnLMc18JJHJ0BUHdJnoVMDhvCvjss
J+iSgLgLH8dreJQKDs4ccdjEI7a16RHSBcZ306y61RNWxKlDZ9e/azXR0ZzwlZHyAgQPWHuU8G/A
wdMscNl8lDkrnw98uoCNdRw8pt6jX+q8pV36BfjwnQ75HTV66BoiSvvyjPV4WZ/DfdPIBUKIC0zY
FExZUyreXCzU0ErSEPfqYdGcSWZjtQivWX58c9FfGJUa4ajoTy5TYNsZ+8xh6V8BuUQab0mkJepZ
i57LinHAoE5BUWoJdTFrr2H8hpmeOC7V+cOd9bWozjIR3QUptj1NDKNwKrDzZ/FWyq1I4DOfw4VE
bbsLbyhBuGFFa2Ltv00zZnyYOXYEpi3jQ6Qv0fLavh0IzxaPWu7QvwNCRggh7yiAhr1iLO7g6yTt
n7tfVwvwWxO73VzPDhyzqYOw9PEHmIkKjh33IEf1WroIn93JzItMhS7dpIQzbFL57K1Hi/l6eu0w
RkGPZmMvKOaxBihGAj6kIfUaD3IxU6IrMddA2SVJdgOjxWSSi+ThRfJ7DJRDqISVaxoQHj9R29bE
FZ2GgkBeslxjbeCbnGJt58bJSNYc/DVwuk4v7PzNZT2dIyI78YtGC8HQEX1C4VKV3qA9HOAZYTh1
kKaZ3B1zeOGzpAAgdRwgHzJB2y15v2DvUYsy0/4hUPZhLF2qVjbvWYPfWvh3c95KHZlsvXVPf52m
vD9CwKpXHoaVY0NWZ8QxA7JZZ/Y3XhG6Xl68docReJiOZRJ3PcrNCmFs2pBVR0YP8vDkbfeHZtoz
FFTG1gO+uRl86m6CvWnrEBuZU28/QRGyvNoe4/a7S3hWpoc4jmAHGX2NtvbFiKQsmOj1omVecsro
w7nwAvvNwJ2AUWdEtwk75p1JpR0UW33XO8nI6SW+WMOu+0eWp3VWrIXA2rcX06iyJWYuUNsLOd58
Qh8wCll4nrEUwwZRmLQxqXXQxl8Rf80UCJUmbPW8mLUeVBuEKgzW7oHM8+XxA5M/XJJHt1Gfx6Qt
sy3hzwT+19Bn/s5yn8ouDHRW7+DaKP4LpACJOK7xk3CTp8qfST52DLA3CP1gjISo/TSthaTaU+VW
z8G1aWEpXspQIOs8akAIVeGGmI/3zSW3oqnXUkMLqEJh6tkte7iEUumU7IKkNal11/WcicwTFz6q
vhoyP7k4RMws3hpGtnCR98NkZxYRt9++68Es2aAU1exK04qtmUOnoDPxVztb32+FN5aiR096K+Ug
NUq47U9pKy83QgSUQRF7jt4cLJVbavQNaJHRqj+CEqFTiwctALMEcLDppBl5+CqCsEDFSIl1od/B
UVsf8YYr4gr+BdIAW6kbZ5Fe3fmSs/XDr4XDSUUJ8YVL6q22GpFrpZeYsUHkC4WnuIcBLOiDaJCQ
9NMg5IP+bDp0NzdOaS8q8aNAuhD8z77gGNA9Vi8n8OqF8oRUVwNztHhqdQQo7JL5OXWeAzoKf1zI
tl55EmcPM0f953fHoC7W+cHsBerKMYny7XuizZJ3mtInqtPHWW4KtqlufSLcZpFYtSOYNzjR+v2y
n0/38WhKeDJHpGek623qlPMeJnkTdbpNcl6ojZ5hdhTomv9/DwwVwfEdQTT2BVOCvvcSpuTuLoRo
Pq1nuOsOYVWVNjWW2JY/50Y54BOKc6vFtGXMd2i1KYHHcMaTw1iklg6B9Q2I2PbYXblJCNQjEZdP
5yTtmOhYIf7e8ZUbCEkzYCY/EwkA9zU28QWldWc479hUt/i9P/tXQBrL0BT8GRx5Fz3sq2OHmKPH
NkOFkk0BmRrWtEJ6F9x44B1ZN5wBX2R5PsqFRWsXV/joOm0eotG41vFesleNcWqf9uZpW6cDH1aU
s7cwWTs9mmlcCkfEVd2q1zxFeVyK2odF8ohKDW+LNyxUWvsvaWs+wy1kvg71wJqAFRjmIV67szKa
Cc8CiSPN/0HfD/xG3xcRTDAz+dhznHH3sXQPFolCHGIvztVIiA8ZdhfE7GAWRAg773T2BVJsfX+Z
MBIuMQjIiep5VY8fJ3dLWgRkzgtaGWpg/8MwS9BvaddozRmS1dqszFk9qPKSxeHMklMJIRjjvrbv
USpWn2I51dieSd9oNPZQrpUpLqXS+fPPIAPMsdxUFiAIODLEaLvoxIPm9b91UMDF+FhECydn0xG5
xWKBlTR0y4Iva+6ofFHAytQ2hR+P4ZkQDbNHyDvp9UHNyYnIA0Rs0tKdyriYRzJnB/Tt2NMg18ej
ZoklB/tQHm0ITyRJ/Uy0hvAOgiiFuHEWhYWFpQf4ZhNu09Lsnu3pJtn8mtV816OFKCksPwCQwmbU
Cc08vvE3GgWLSCBCRSc4DHsIngSg38x/RJzBj76BeqqCQDq4blll7lJdzLLa7m1MgI6GsGQsqMAw
dK5s+WC/brEIqg00jCospr4QP4qdeaG2sIvbmoBn18FHSNiosG1IMWvEsLE79i8lGdFnmDx/yPXN
Js2ylnqVXfNElFAV1yRWUqauCXDYtO7k/HjIS0q31FCCTF7AOWxHPZXw1IM3CiPpx0L7idiyMdsm
i9GZk8P+Onk/WsB1WQOik6cSwN/90eXpzytxiwpKtIga+AXv5EDMBvDVlxZbaFozrMgjOwXLN8yk
wxJE1Zhvc9yCkkWuYzRkjEB5xaJ80q8ehZUoPTvwQet303Huk1MKigDaYU57J42WX1tjwJytDCt9
I+wNd93OZlozBe1R8Dth4Hxo0Z2ERik3/Fi7zsidXDWZDKiIAj7F7K5RouVg4FZ9oAArdx7fQ/ri
98MMlrZkA9DU9/AW43Xnsua8fGc41pDELcNr4HOi2mn2t3q5JoE0l3XSm45FKc9toh2lJDCR2gei
Z3vFBuxfDJLLJTpyt8La8Yk8AUyCcHbGeejrfjMP/SQMB+8rPcJtnvmPLs3A4yHsb7y7Dx/LUZB9
3pHFVxrXBRUIkk5eneoND4E41Vr1nyIMARfK1earo+CVH8JdL4Z1M6uBIkHFkFfovtF5fPEeoWAG
pwzYArKi3T4Wo1ZGe/HdbbKkdHkjtrblXaYxuVLfTonFRgQZOxLYyiWuCgT7ODqa/APe+3AMHEAJ
Q2SNnC5sIE2/7byr/3Btm97gIF8s/TLS3u1GHf7nigr2tyVrWnSzDavJ0kuL1VHAEZfeGMshB75u
HYI59OBCH88nTlJN4khcy9pAYxgG1RnzF/2M8EVZSxHSZTHsnTF6Jlsfu2RB+ALaQLI5Mievc80b
VCVSDSa2IzOkt7015yAS7QLJHWizitBigTAIf2JqEQWFifJthPBxEVYlhG1mFo5iNq3UHM6EbgYR
QDATweoi69aq69MFREE47eLRCAfzujkBjrP1TQ/Hkg+k2uOWKi/QvojJCvfT1nJ7h5dWqIYbm+48
uzmfB+/gycsZGmrMfXNKLWarEx1ottcmrl/t59cQsrieKC7Cxj/GOQ9DyxJB8rfn3n/4uP65sInf
5puwT5g9o37y+k+MRYLJ+ampSXBWqSuY80DFRZqNKtsRu9Hs3GdnC8oIhbDzP3trtV2ZxLfHRfTD
tgGuz+7ee+0xlsIw1DpSiQZLJOR06HQoHXIpluVsj5Y+x4/m8gKhahgie7WD5tej3lL/q9/1HwKf
Z6dx7DrEPqG67HtcFuXTPZtJ+Mw3vxbXJy4fDVOhDO+Sd2Kip6ujW6DBiHHM9zttfNavrwbGdj/O
qH5swnZrgnt+CqixzLdY4Ne1kOYLUHsYRlEit21PtBnwX+5O/tPiD4FWWcM1cwVYBpO5Hi+Bfjb1
2o2WzMzbRFBA462V5vVSkpLU1wSlznwXeQyeQbDFAUBMib0pohvZKaLVmnJfmzqJzIfBBlQoEpsJ
2m83SWjzbSUvktb0hBSi2PhsO1e8HQaU7y/EiEmDGfbWP5a7s2dXzxZSUh8FvKcsdROnGrK7TC7k
rtKChtFYNfvnAtm1XdHFAR1Q2re7NUn/JYPmkHGbudINizCzAOBZgUWd42X1h88BfyrovXjrjy5r
R9D1BrNvmwnoCafhg7NJdxe77BFuVAopC6H9b8/axk+m0Qws3+FHKSI+sq2adlAvi8WETEm8kQKr
0CJyNc328qyMvsQ93iOGpJqtQNws1Gp6r1oF2Zls6nIaVQgQSNZI26GPyYzAV51UC1BaKR1qcCSW
timzaSFyY0xRxrgrzsca8IkD6Dj1Vc7Dr2DJFRUC+Klz3K1vP4bgjaBXbGndM+wE49EGxo8nOQD2
LgITxvBKvPoT7xkTkSQCg0XJqdz+/8LiZPBLLSycaXqfv2FpfOvRBJzAGXwieNc7TzWSq0FsQAyZ
wbLqipnUAzdR+uV6AsKlZxDQqVju7CutH7XP3jkihJGTUcq2dkrEOf3Z9Nw3WSy5M5tv5BXopJcu
L0jo0tobaPpoacZquuETbwngtgvbcPw/5XzbsnYTNvURF0YiW24i8F7JS3hYFpEdbMI6VSRV8ie1
rK1J0rn/yrVZceL3x2U253XJshhRNdRB0wbpL2Pr/3yKUTymUeo9SloiHK1ZdnG4gI2v3II6llWu
Wu8FXXHDyoOT1t0zAX0mDYXcXHNmeGaNLqlTMuQcogGnJSlDjhnmkAZ7kWx5xQgqt1TQ1jSQu1Mi
beNLeGTbEDoZKhMd6GGioEv1c9QIELiGXcGJgLRD22FZxR8sjicLrq1KYIxjERjiVXyAmu1jQW1Z
cbevKNlZ/oMHHs/td32vOiIxInpiwhMTcVbnLr7/C111Bydyk8VQXYCBNwihpcOWWJ1SxT6YK8UK
4HUAxPGC858XGkSfOdQDpO0dv2uWtps15/FnPl0K5T1rYZkDg4HEs5lRaNYbcIhlwdHvLAGy3cdI
rH2ZUnZUJSC1kIXcAIOJQcwW3jNi2xlACQMzUGfiUINc1QcGlb36ALc8BApeJHXXHbTU/prWCcWu
AN+/c3kWvUwIWwW2dRhFuY7f1KoRz7Ji9BD5+gQTO1PLAQOsOkn5pdQdaB/JDdLZd+ARx/7mfPI6
O7Ur49BAiwiT8lmsyJAz2KhmoL/egVL9EXEzlJkK1QllXf/f9+gELB6BbYQ+VyqssYpcc4hTplUz
3rf+S1Pb9LgpWTeskz4eJdIjqIIjsijlQUxen2qEfmT1pRyaMb5CUayWYIcO3ryVT4KBr2KRHdTU
atqNewTP1Qx2gGgupkbooz59dl/bOyz4qQ6JDoIefEk+lMCmilXb33Hy3tqYM696Ur6LkToRgFIA
4cNUpWhsxG52eGV4awZDNMa9jEOET0kcTEaBID/C1Sp5a1vNS6dNmKAVCrH2Ro/gPvHiP3puHwLj
a2kgMGYHXZ3qlxnU2o8nB97iHYHpArpMnxZZuPma/lNJ1zktAzN8CPtTkZIZMR8bcAsyxFvnekF/
VJtK1ZYsF+pFRp4JR0VwULaCTxj7nzqzUw8g+RmTWZBodanyvttsyuhuHwTQ1r5C91h3bm15NbeL
zRi0xog4dxUPKch2vSYewpLkHgPvuhqmls3rVvnIQeV0JIg+PLoIdjZNzpuaxhiYCeXT500VNQvp
f+zAttcJkdZjv+vySIH7m1e1ZfcTdgclMvUtCOg1UaWc7OYuj6d/kBfk3pUN8qTgsXr2kxnzofjg
F5fgz7V1B5jOjzg1mF3coOKMXomeX5RI+64EhxcVoc4PIK/TRuL38k6eKjVr4QHuN3xsF0wT3Yz5
J9zI3unqloao43kbd7gbnhmyrtnLsPyEc2/4EvjMskSAffqGexuaSmzYpWb2hVX7dRgZRqxByypW
hlRwuXWc6WdME7zwGXU3Kbao1EEV6LLwhmHeFozmsOtUy5disxPUmsDrCEmCLNsrjEGX0g04gjga
KNTOa0x4neyj8xmj5M9pwTI3xy2iTCCZNGIZubrwOzIChlGiSGigriF8/rg1HqiTwRv0q7koaKAT
kHQr0312g+cqv9Yrs9fd2cC06tncybnTjMd6VK6DpkBnAocnmGiy1fLofCiyi5FO7CKiUC1tDFOu
dMIxIjOxKFIAV1lu4tWs1OrP9hEUxqpkxPOLE91Qf7kkgc3vXAEV0UmEJeWhwxsMhjIPs4nvYqTJ
e8De4wSkiylHd5YCIasUID1jxfmUljuumiR8LxV4ebJoOq2wR1fz50hyOZgS2JQekl23JNHiWSEm
Zl9DdIEip1GBUq9XYYKDh6M6MuwaBwMTsX9aBmuJaS+K29WY8vEldmRQ09MuaswX/nlRhZrAKUAp
a1knWefggtFsXrS7abfXWiA2HIAyiQrWdo9b9jchRIZ7IkWVaGxrkf2gMvN3DgHR83bOEpdXjiTD
XRGmBlG6XO85HnlHz7hnTibuMHbVgf68XAxVimUTaUWUSMw2X6bnxdtu1ZYbxPrZriPKO7czHywW
4DGR6ugR4k31ZzyTPVDGkZTOnul/fhfZwsO1ur7+S7Z4HbNHP7pEBRim6zdVLAE7S/6Z3ZAQ2F2V
A8VuvjTTPjxmrcNM196eY6I/wnHODobSUoZteNrMIJXPExNiAGfXJn1fxnIvUbxm9+kgwZ6cQUej
Ogbp/Ufalf4nN1QRsK0EuO/yNbDdLoHhJu7oxSPuJvam3F3Dz+Mw3wK2PxRMGw7YA3n4x1Z4Bvsu
Lu9XzuOGJV/eglC0YlAGZtDpgjcxuwmBwD3zrzN0Q+pYXXnMT2Fuw81oIQc1J4AWNN/s2ERIgonh
+sLaPAM8f7MXJsvQtnrCseaIxCZMjPKBvqDA+FswZAm0KpzXStmUKfOhE3UQ0HxTgo1nFDOPgqO8
vQZf9YSyk8FqnJO6zQp7jHNIJNWfReuaNQWqV76zc6WcImJ8y5xa+fMcyA5+LADzsFkZeyMYLWfX
9pYIFWAjWXURrG0KESJe/d4BM/+FmsLYy0O88eRIRig+Ilz3/DjDUyWfDWngLpK2eBwz/2m/scoY
h3TXOVb2J7t0cdfNKDyxLJdHRvobnXg4qtgJjlofBtpahQWp/jf+EuKUHF/F+GsaW9RDzl+8deRg
H6o2y7piWhPNse+DIPNEKAp2aH8/ZEZAtWVlllCIMCz9hTZjAu0OVW5wewF0Rk89KePDtNWS6f35
ui6NW0/uEVuZjJZ+OJ8YI72e78fw6Ufo7hwrq4OstjMbnuofkEGyhniuOXl5CVtf6r890wSbCde+
9ZAiKa/QXnNCOix7jy7Gyf2EIpvRbg8dq3JuOZKHgQfRELE02szJdfF99HMnRzSNgpqzE8dgSGyA
W560FFlcnr0oVbB88VbowtZ8j72Nr/tfOrCSppITvUdzFq0DLEsmMiEXLAdDhGQJ6T8NUlf/Khge
iq4YNqDekKfYH2iZWVJu9YUc86FcC2VA7oCT0RwTpi+Y5yNyFCWp9xOw0F8zWYz3ddj136Dp2PJE
N3gHokmBlLD7ZTHzK4Vpwlr5hgK0qj2dnzsjZmOpwEqwmZbuaBq8JGmbY+KKD7V27GXEam1+OD1G
YdBwUXPamtC71WdNZAUt5eiUbmGnD6ob1jbtAWlvGVLJiyvp/NLIZyW7AYXKRhAg73rJcuOg6vSb
bhRwRF1D/CTr1uiuMhljJNpQoeTKAUM5SxsDGr/R0nPp5KJ6kxR70mcvCaE20tYJAkN++FSFpphl
peU9T+X0DjwaxaiF2Febl5EZZk2r2t9OE4Ev+679shBAMYcIeM9fZoKIPvRvSACBofsV5yBX08Y8
GqXY6wLF0Jw4Lq57dfHsIRZqr5gMWtiTVXMpyEuh5U/C3pCQdLu11XutMdpFSrCc0LcWObnJ30Gb
7NVu3cM6PE/nVHJoe7VzufeO7JzkSvBqzzFAeV3q8jXtzaz6E/9JPPAltwqc/45nI2a9QGcwvTv7
zELLUCUEtX5C67SvoGY6HTgmUhqj7l2Z7m9x/UAf6rIt66HBQ865S4mDShKqvi4sqvJX6xUbv4uO
N/QXnCTxOjzjbRnQxw5G6dTW7CgUAwPCtuSuDy47ZzdnygPHyPLX7pHQ1uefYUeFvM7HoKWresal
2OBYF7079rUvE7nfHzg1EvFcnoy7PNrYQkiS+2UmdfsDAbRX4h+Op7fHNCgdVKvCqVZXSL9U2N6s
18VAazH3YwBqQFexDQcs3kaHta1TY7gAKQ7Z6sLOcCSIZoNZh7aLEVvuW9BNy6jr6YRgKfd8YcuX
P2/smklCB6EDQagJviktazfPh4seUFWyoPYpJ8Aign2ZwbLfceQoE78XXZuA5e3EJXFQsNayL6TC
rYFSkvqkU/1QOp6waQGMCrqnR9+5M4QDIvf1l8VBq4JgFsn2nXvucMVITsExqQ9KOyExASE5dmMR
7OCo2VVGFF34i2VeSCFwgrmY/Rw6/DOTzP8LRloGjAVbW1N0D5RN4/07olKVio7xHqR2f9aKYJiC
C1T1duHST3wBdJixNFoOJzpw+b3wjpEWlYeqWrldRBpKD4aOdW7z4mJ+sTpPfdfAVb3NA9J9ivOi
BpbvRCDAI6yaqx0VRF5BWSahL64sMbOpqfOCcoFYO/gOTBNti2VBjAy/qspYh72aD79hjvKLFU47
o0b4IlbPPtvSroDKbEAdqExmJN8DD3VAiE3RttxX8JmOQ5CyeMWogOhkmHpQw/7Racb9f8Yfnh3v
xHQ8NmO5uLEQxxGyU4o8xYdCGgbr6oATwbGtH43f0n343VZD+y2WpRXUfmND8bP7Um5LnDZA4Df5
EXJI/51V6FZ0l38C+mh8qcAdCJK3eKUVJ4HqMveel1PCnfI8IxsCrxZY6IXsuFVJXF7ELp1IxyrA
QuKONXs9j6RPCraSSLl07G7UX7zKmoZJIZZvz3KhZtwsMFGEorstLhqxJ/xfoLhJi9yM84K9ZPZ8
+6G67CFtfxDjtfIX53+bCNPNePE3eIyyv96oPGC/vQ2cHH5tt6ikkjer5IcaREtn4MF3nAvYMuzV
/Yt5yXucSpMS4si9Xl6VRsPxZHZ8RGFrg+62cN7fsMqZe2pus0ZUMCUD2GdvhG/FY8NcN7c4ax2Y
1FlEc9LtRKF4EBYejHfdVyi+Do6MFqEMXqUj4K95NvqLeexAbcgpzwz1RUm+NRuP3ah72WXgD98u
ojR9sCcW2iWkGsB3km1lFqRW6qZF2O2M4ZtLmLDlUjPMTVX6V2fsyBDhqk0ozy6c/MOwkruBD4Mb
h1EjHXzhtVAyiYkuLFWBNs2C8CZx8dV0/YGdDAdDOHOuWXKe9cRfJ2pRTe+oNjZgSsofhtibnb9a
pYP22A/GAqOi3AsWi64tc4H9BaTRS2YOHH0wazW+3+80WhpGNXDWb6fXZOU4yeJg3ClzBX7ihFs+
n+BWlKQB1x4LgS8D5Fp3LGmpppiQ/AFQf6PIRTx6s8fdhxA+E/EfhamO2VFF5d5uzsA256wq/DPG
Flne2HW/tJ3YaQT+OCHyYekSXXJnclEuJcC69UVrnCy4t0Cb1ARVKi6o1bCCr5FB2mYrBxtp5jT+
wEN1ElPCeo2YbBptSAJQegdgIe+/EO11u0JRZF9iedyez/eUtl2B0jZ4V4sACT8U/GO+x65N8xMP
ngNcenQy65nOYRg+iI9kcw/Y2gXgTbrFIOgI0YPqiApYZN7ojuGYMxR/rLCIa7Qz+DNJJOJDdn1Y
13/0kNjSVbZuGoV6KSaHejhsZnZKmFX3T2LofUHoOYvz30gCu8D6FBA+VNLmki18lxWDSYMTOO4u
Y+m2OjQ6qBpnJnhNXLDSOiKZQvJ9JXFdRwD67LChHkBjD0LdgB8nqECBFJTbH/BTjpCXhtL5xmZS
RWYENpNvoPrLYaOe2B2Ajq5IGRuDPFKU8Qml91yM9U8JEId4UrNbIqLrCXIBLJLDB1O0x2/h89rj
w/GYd0pc9t8jd2Zs8iNKLW+gBisiUhj/YQOcAWHfcV+G2MZPZ6t7Dtyxgc067Xxlx725kqU3TrPI
3sh6EcNG1TgSeFj1tpftVAlJ8xNbTP4OiUY4zzS8XZGNU0koebWJJ3cR9kp3Bc9GubF1sHZU7Blf
zX9UiKWe/OysUF1VzcCAmQb6N+Rhw/51ElBxtTLNs2mnddZ/K/Z84FHT56F30VjrBeVEsevaIt1v
oXcpU3whfutirKXYTkNNw4gzIDpD/Tz8GckZe2W3bHicP+qrJZ/TJ6Q6lB8RP28Qq2vr0H78g+vc
6zyZc2B1+QeHxuBAgxFFL6jraV+XaH4vF5QBmiUnbAh4WNWlH7NDOBByfTs/FIkssGXqLq6LalsH
ELvg/y4jPgKTWDDCv/zbDpgJdV7Fj+qPRuYF3LXFhCK5wjXlHy9lioBx0NtIuEk8RfKgVkj5STdy
M9amtQ5aC7ld+7EXzYPs+YjYtgt/IVwGwrl4fYEAfqmfZJ945Dnu3eEmx9ozDn0eiXJy6X1sshJk
jby6Tc0ZqPpDlqAO82kiJnZwoShl+/XAqkscdf1+WRDhUjM6uwJW7Av+uC+9sEhHUylfaiiAm6ni
tVvolePVs/3t95R5scgtTC1mV08uatDqUqafwy4R1km0mWpFEgPTpelzsie9S4lesra7FJYrLNEu
JdjNo2tKcov9cJEKU1j0Ow7v3FQpeyYxLu20MujbQzbhJpMxmEq+3MGFyxTYH7DuTQJRG27XqXtj
d3w0isl1+eYFZ5qynu8hMQBi8yaxD3BOq0GJ6CeI++9WSC9rPR9Roq9JAD2cwxXjfbpnrXJOdlXy
hVWre7k8zUUJKrcgurB5i3eHuU84M3OKkclEt7xlDnIhtetyGXWEphfdY2hY4pCfz1JtnqNMbwj4
F6GZH0Y0ybXKwV53KS/p3/ylcEZiWg+Iq2X7Ohd0IHUtWfNIf+aKswU+WSq1lrz7vzHugRY7cvul
l1Fd8l0MRwocrvI8+gDOtLrWyNzED/kSgxonQne24q9X23um+tyK78UupOr4xALqrJddpUmFTLvj
1C+Tt6ummvLAyYwppFYPgnxN0oK+25AMPoHOPqfI4i075M34Qpo4PFwlvacecfZ8ycQ44IYioy1X
cAQ52hv8TLNCat7gXULQoRwTvdtTlu7fnw4ivByvTpnV6dl/8b+3PBi+m4nTdl8nfEX+ZBl+QULz
9o3yG/4GxnnIzV4YHESmOtH9cpaNSe3cZmRda/nczTkjt3pxYA5wt+QScgzzBDJTBlytslsrGdqM
/EyaBIW3XzR/237PpirJIc8rLBQgYT0WtHJLk5vcIQ7vUjmS3EpncZ8R7DSFXeVxhcCm9aKLMI9l
6K5PYSiJXc0eEzMIq4iVptpjWfzJIj3PijIv1aBXtVYiZzmP8TDxz6xng1FCFAWPDzMPHgWGqro6
pljrtk7/sWufSndH/w1tLWBvs8/klb2tHyGwUnkc6mL82MvSEeTmFoJlIhcSIzyKg6PKhJeBHyx1
KnqiCvefOSZF+/j4UpEr7/Ba29Y1N4ytRKlxAQ9djmoo0WuUL+M7xRWl8Ulq2OrjecCbgTqFk7wG
QEhCAhsSoO2r4VQ1q+HsWF3dK+W0BXNHWK0rqo76AoXY9yPRmRlkod8L9yLWKbGcsJAC2zbEs7NQ
VUTt1J9W1ln5O2hQzmyR/zLfIoFiz1ldQa4u3Z4uj2cesMAsuEwoH0Fp4/9IitT8Kybj7kFncyRJ
JQ2i1u66UduIXXan1mN+8Hg3VkjgL+eCYNf9Ifsal9YntQatFuqmL4Crb2IMSpD0+jr4vUUrwQtK
DGWf8gbogpN4GrhFrvGFQX6gizL7AluONpCjewc9NH87WE6MKeYgN7uDDNpONqxoZ9mfXJ9XBPEH
sKJ4gpDLGJjIF2/GUfhzx//K+174CsM5LB/eJ+szu717jUjKicCYrR7+mMAQtGl93clx8dWdy8Ba
gfWmIK3T1gjmAghnx12U8gG/twqGikEjZglLYJzxPi8V7p7p3hJKuptstAR9zCaA+IsWHnEolo8r
TD99s5SAKMWTa56lxY2Hz2/EZgIz7Y5FvWkNYhO9cuib+oBn9ss/VH07kU45BO8fWoTNxM7bCKdY
D7xf8crnWAQNpNh1lJuPRdZFcp93C64E09rNQyD4LwN9G4QvNimqGxxo3OC2P3UgzI0DUC+Ybr69
UAX54jLaZiWXEpARY157lmhWsPd5CAJhwJtBR0jMymdYnnPxzy4xEVMWcN1EPydc3QVJPVSYtMjZ
5zRB9Smt4h14n2GJmShggnO1QQnUMITZ4D3EbZh3w05ifiZWhpp4s9iY1bkLbUmo+AfhKFbcsWVk
g1k16bneYebi/4ej/rUCDyrLhSOblV6Vwvy6SMLkldK+tRjrBTBHVlxApx7fQrnzek76JNF4HNpP
+0Jh7QBAKJRvxvsqWPbZnwjorR3Mk3ETuGTRJwKHEicc5JNdVdHZeT8JJhsl0pR+1C2czRSHiLh/
qsQNU4DS3yZdjR/tIFQk3p+appZd5nwrPv5yV2eXQWafvIcscaNISQ9N5RcC9X3ywGkw4dxiURPf
38m8fj4+OhOnouRFB95KM1SyrG4NEX/eVl2DfArm7ytHvS2a+j5f2dAHpzCtlElRaBSbSww8oAq2
5QMBWmPJcQ2xR2cxgQJg2jNADX0KRsrdbJ9PTJkbyo3qVKgp/YFJO2I7l9u+2pOskxMkj0X2kkB7
/VXC8p2FoJRFnvALKzzV6ZzhwL8qs22H0jlEivzOnaC/+ktTWTXy9eS7eSIDVp+K72C8UXYnor5t
uFnb1BMt+gL9QPml9sIF3WiMHYyV5IEW6wZ/3ZYf4xwLvWdBYIDjvBtmivNc2Kg2DyxhGBnjImWK
OodYAZix21rygy7Z6QjFvejxzA4N4o0TKRhw+0w0OzInCqsKibCm/3glVTZi5tecZY47hLgSHpDc
xQA/FjTVZt4O4FZxL2ib9MtL8DNPU7qCGTnoFBBtzqCqg8oAe9r/zpQPcKC9Ut4zuQCHZlYgNbWt
XsIyvRtKWMUoIWf20lVdyZaLgTdlrF18b1piavBkHkXnfmOUz9uV8PlzcUm5Y3H9EJL8JNwWRzYP
zKitF2jgnx0WH9RRFhiYR9gyYXsk46B4QVjK+w5mSIQsynRfheowmg8tS2M9msZ5aNHdvsP2jQQY
1zXArV9lNYjAX/AgZfRCSmwcQmmpHd2PawQKGqotCm9ZHEzElP4lDTzwYyg/uW2XEqim9Di2Rq62
fO2iy/tOx6EaSNKKxCOFi4C4PpMnnycDwBQYDMnrq8T5SY6B11FZzEwytR2qLepuecKjP0JVHY2K
LumJ+hUJ/tA+Rs5vnSF4gmK34LBDb5k7O0w4d1t6FlENDZ6TnPmyd3N/ylcqMFLlj2oQYbdVquig
YtCUPWdLYBqs6VoBgDfBpxNqdp5AA8BEasyHpLzYnWPcRYkrYmqUp66plfBAIpVydCYt2srDkfx5
vpcfubfiPNjnjxh7+gG7WdGpfGJs0kspi/o/JFFgTHa8/U4y4XUqkkuUvfu3XfIt30C4RGr05k/X
1UX6xItkJeRH/0xWPlN0Xh51k141496mQ7WBLTiYK9oMKysK8X2YbUsLo78gyqrkcy+RbsIkvech
0I/GD2ZhWBs+rGpYAEWx/VA5M3OIBeF3nLc2sQLNUMB/B3yV3M+/fHis02P2kJGmR+SRkrF7Fwie
i8JRwMxmKNaWl1MKTCMtITGe404oKu6qHvzq4/o9YwupjAmB24VTQnkB1pxetONzou5bqqN0hLHh
BsyXkIihyJe0YkjdaP/FJ6Gt3FLunAIl8NmgRkgpxHkIDGzvk5ikpSFH48Q5Z+Z5blm2h0MT5kKk
XkNEQT4YtuvodT+XgMYcjD/ccOT5ZffTTgtxCPIDudytXY9ZwAVQcaO5j0H2X2CXGqxkFkKvqmXU
qHJhaOKOF9m+8FpjTEzT7X4zR5OsLjEnKzM4Y1alNFFL4UwWC9YCkFrYK6Kac68pivOfhh4IwnNw
1jojlQia58RRL90+SG2B8++gnRsDilU+I7xQbVQ/5Vkcla4eQa4N6yE3syctk6GIAUDf4fYQRA0u
ss7GY8jTGXrVlZII8SSukUtglgaVRsjJ4CQuX7YjzMUtIE5X8LcB7/OEM3doHttq0YzW2z5ld2DZ
2bS39CrHhGuXXf9GIZup8zYX2LC6bpBFMG30niD14ThZuKdeWnudJueMoMh/6K8KrXwzJFB1lCHO
cl/jS7TdUXeBLwSl0T3oOJzEQo7B3yZSS1Ty2QQ39LndrGnb/WmeKd6BUyJwUkor0jepwTgwNEzn
hYVeLJEoq5dSDJPy6iG8nnIHcpc379a4SptUus96qh37klmL4fodvAHaD2Kmfiv/2wdtHDaY5Cq2
vI/HrhMdr2wTLeqK2Mc48DhEyZJho2DW5b9FXDGE/vTVDIecSM9kheac/+M4BOY/3/fmnZvpFX13
DiqLOGaUHWRO/o6cU5/1iUpulThedXermiW++IC8CaGD43645dEDGiKyb/2+NIHdnzM2CCTjUQmd
X1fptVPjmqOShnZOAHmApQ4osRP55RB4xNB6FEMGWeWJ0MCo7+vApD+zEz+qQxLSiSVKs5whfns/
L8GDkhYymuRz81LPLTP9di5PZgpAvZEozQt1go0CulCW1rJAnkcq55Welf4rTO09MWEeaNQJwdel
1PGR3YVvMYCJhNDVvxwkDB6F1fZfOkRXgn9FPl61EjRZmiG6O18gHfg/m5Vh/x6AOpMjiYyIUe6v
V6H/Xq9QEfcr1U3av4tvUE9V/+VTt+/UZXhrWzJX2UysUn0P2QzuYioyE55OyE8QD5kN5lskvBRE
GjnyJP2NOIaAbHjO1o7h3c6+0NU5XY4Zxm8fPgqKlVWlbMN6LAsTB8k4Q9jxp+1Qy4zkkj+hGWCN
XS57rujx2BlQaHxh518x7JVTS+nHzj6U2IW1Ycn69NX4OXiVKonFh9ULkUVWTQEliVnmBtlCC8zc
HZ0akABNZ1MuC3O/QWL/SzTedD2Wk1O9TjtiZ8LmWfnGUIx5iNLovJKPq9zjU/P1ScqzC4tz/EEO
uocVyW+eXS0Qreh+zI6RJJ6S2+wREPuAKGYetlxxwKq7YpnYpmvS+thSqRoj5W4UmXTmiv5NUbSN
sxBjE3B7uFLQQT1F0kIHtSgUsXGLVhd1OXOdnPCbzfR5s9HMjRE+L/bx9hu97W/ftRKv3J5rMHOE
o4fThNnQ2E4HRy73tAwVk7CBzWDBIpy79ZUA4hJe/+zdWBfh0WiCQXWgYBvAHfGG2n6yjxGkxqG+
jEibR1PkbbGbrtsi+K+YfZU589mTTm4UqYZljouCkUmGeeyu/3jDL23hJPljQudann1T1eSS7HW7
wkYGS7s7LvGIZfToYzxwN5DHjUGZPUywRX5Y2VLlCGU0B9aC5gTGuE+tZhZAZJjK/XO/vYh9n75c
ybCa7GnDpvwGQk1MOaV7hxkbgA1QEUSEIWF6SvD3keMmEvE2P77se7qBppv5lM1dLqTlxHW8UOoS
ZAnfcC3XbCmuXJte7xxtCD9BF5Y2j0i02ATOJTq/SJMBwEmhuxCj8+e2jqXmH/8w+2529nF2ehp2
UhyFGmMWwe4XyNg52XMxJMx5tYwQ1T/yqM3sV8JuBe+7dsxZEzqJEck9W01hkbYeyJmftSzdX864
v+IPkvHL+Ke3kiKsen5+xHvhegFKGnzeSjOOWl2nVUI6EvQ66mZyAglL45BZhjFeyHFzbmie2Bls
9B5pRuJvdr2/TENR4n1Wj5neIHF0URDZgXsXOYMr+X0dOBhan7Bwvmbr1XQg+btihore/5hUgUqJ
BsPqLGu/jYASvPtWIcrDiaNrPD/E0GbPTSHaIwa7RMT0/S3p5ULakWJM+R3wAuvQgaB3Q04kU4U2
z2e6u+sI/6JbebTq/qYK9C0WdPQoF1NOw0pqCk2ex2Vb8OMo/PsJ6W4ZWswOa2fyBmVdEDOuIhTq
oTTmA8AwZPGArhoxeLQFGdMxytPvHq0AdPEDWOtBpB48SAYxYjj9Ifc0m4ejd1g5Wbl1eHkqXA7N
E7JpsngHGiHCakrGL73yhtKXAeihcBQfhf8JGetY1l/FZ3ujEp1eB4ZlY9AIMj4AqiPnv7IiqzVg
1WK+hyRIRTem/FdPeWXmSLHJbhq5qRTwiyoax4xRYtvTwKyhaVHmK2QPqtgbHp7S1ShgjpWeQLee
inEAH/X4jQU3OlnODWhfeWSZQ38lRZjHtBNUHjEyktyicboCx3FfLiLqcdCBQstCfD6+g24PMQ12
WDcgpSftayl9XmvzfUcKNB+DsUS72huA4/Y/+EU5/dEpGLZQnspW2URIrhyt6+Gr00LZ51QLdhaI
wKWWoR37iNqJ/FCR13GCPSeNXPjm/ScSrsKp9wB4v8559R/D/OrGr4TOIFiVu08WYOkt3uD6XMgE
uENgJF7xICqIia9n+hdxkiGyrpqXY3Q9kPwbn+4q+e/1E/eCjVrlPSsIb3iC55xlNT9+PtBw5nW+
WniM2UaKuvLNyLD2wZFiSUogjRcpKUF3Z5S9LYxC9UjymJRdaUaPuaTqr6qL/4s8yRq3LlLY8P4I
WwDSb/SqKxGbaF4KQLQzhC0Urin8TpgVAD70BTgPsYcxp6N3leacGjPYEg7hgpKA1bSdpC4MEg68
tac7OzgeFxUIp4ISohaLEYEa9AdKrxnrxbz0vq9cU/ul2oOBQ0gMzN00MsHvBKinepZSGbh8v97Q
bRt5vpiFEaLvo51OQWgAtUvi1Ab9QJtMlgvRnVWXvgWIRYpCHRmGkfOvr86SN59rHX+UUCdPLs/R
oaznRI/5UCukgwwUN64kGYo89rH4dH/p1BM+mlZV0z1QQ1TSa4ui1H9yNTH4KW4b8G22SmWxidyb
8MxpnB75z6NbfDL1sh4kIq1Y0LKHxjdtG/VdTgV7GNmd0kfLp3c0tKIZesITVCuB8qOQGz6NPe0t
Glr0TStdxVKi24i9Me6s6vcvlN/hj7sEiDBy4PijR+CfKqcY6wFlUDqKTEb4QVk2uZ4s+jregwma
NMAIiVm1HaD20PYXUww0ZQeLeVGbkhKXpn9t2N1a51G1HarcjFSj0/NLgVowZzpHzZg98fOpZG+4
dxvULvrHX0TNW4+uPhe8WQnPtPBY6CZQhbj6oJT8CBnRxdYJtYG5VprJcQVD2omnQmOlZ6P1bX89
rzB67Xxv5T1S3VP/NUHS/DqStCLRScltmYPHHwX/6Fl01hW55+jkhXB3W+IRwDDh8PxYi7naP+jW
jYe37NyAgaFk4Xk1jfmPCiJoAOvsxdaID8lH5ZzonP4DA3u5ovnojuxgkSVAzKeZViYYjx3hOIA5
oxouqrq7/0X8TIQ7brABeSDdiP6wNwAHeaVTxPm+VfaxbrbLluRR+ZQ9lrLD8SypcU9ly2FXLrL2
Swr7sBBSd7026k+l4kcibGS8413x+sffczOjld1qWN+rypuL+qfZ8AVedZZGpo0EtyAxkld9TT8C
0ZiYF35kjKjNF3IgRPCIAW3CTWAm3PMugMk3boFYJN4SH8eTPrOviuCKGEHbl/qobcPQ/Vetnocy
XyEhScx7uzhpmkNmKU3K/TJiEjfPEbivcLzXdB2vlOfqgjChXBMoiFYG/i/YYL2IOVY/w1DRcqBH
B5XHCDRTv4Jvd22gShpbNFKaopUYL1Ia/x/mIDhf85Z7vNn4Vxfri2iVkzeUTA8Tegjy2ckjsqD4
KUqW6RZ0rcnQl3kDYGfSB9FYib3Iosouu5yM+QXX8uq3C5TBuv21HRBwV7+WMa9lToLju8aHdsIh
KrW4SwKJyrD37uVW/hPP82238iOUqO+vz2J7hgr1njPwnnNoMp2aljpOUCgTUGBa/pWT6qlJP+It
u0+vbsja9oMSslKTk4Exgn9KM+9cEZE79ZnAorXe5APDIO3suxvKP5OeXnJGo2pCPdzdTowbXJmT
ZZLtH6Z+tZHHizKf/rHPruVPyDe/bgPxx/2QIak56w4ClCuxrAmIjAA6lrlCwfX6+7/Oy8lM7tkQ
kwS3AFHPCBIHsDlUFGNsP/Hifg0jRk1fOBzhNDtvT/0vA5TTNVRnAIUzcHWPWRNtZHUNhb42Kd0/
UpJ5ZBfh1GTYRzPDl5wC+ZG5afkos+WAn+/VfIoUvHgG8BtscSI5HO1b6JC0ZgHcyiqe4mJiWEEG
882bdFYpXn3h645ZMFuE5U+oYx6kA/d4FBQF68RiyR9P0QrlVAYJjEPdbRn1cNJSLLECWFq6LMk5
7s7vZZ4foGOQEdkuvY4Vk3N5CLTNQP3Pjr4LJu/vCTE/hJ1hsb+tLfdajrNdmRg7tNKymrjUURRz
k/F2VID9gohTgGBYRgrHTRAVQMKp/UWIgKD+V0o7NdXUpUGFzaK3vo831YHcBsNfAdF2Yipkd79K
99P3Rw0r6Q+zRTHOvDrMif+ahlEYa/GUfGjqi1+WFdhZJKESpQAAbXP8sKfqKyi3/54jDD2xfEKW
yy9kH+ymtTl4flP6pNnrpFwE58tTOPLo5/4lKtEVqsaWoJwJFOJh/7T5khQ3LTCH3M543SYxYL4b
XYFQbe8NtzJEShVyqN3Xhy+pdsWcqoqDYlma2JI9BTukxg+NJs57R9e5NaXlLPlyTuhPwSwfclDK
Fi0DPMWCsRnOhJu6kRoNZTlJesauX//1OG9FHVk13rY3Y+VjFVEJwAaFfdh5bjUHUgxDfauhZxZl
CD23/1++WnraU/n7Y3kB1EiJdUm3SiGRwYYbdKM/gJ4WWNW/ildOYwnMQB4KWHD6V54jzqiyGD3p
M8nOqIHUWHAktDwvyNYak9Kt+qDpY0qCleij7GGw6NfvATrHcULL4jXFXqa6gOCOII/QeBcrSG+q
EnpCAUV3LtY2A97iyAAiGHkfvbQS69TEkkmeQQhuHUcxRawbUBnWaTw0IBZPm71Z97b1uwqRR5zU
3GDwI+ThMZNDgpiQRKZKg9+bSIAgoXzueWjEqR1HYCNFSySs3/43o23uSYshVb5lZunNxGnt9Knf
daQP47Vdkb0A0LS1mBAEwsmCLjbRFK2LXE0gzO2lejrcBBodXL72lc66vJn24m/j/cH76PuyCZWv
1WbxRSlkTd7AQxOHRKI5yrUnDdundl0gmRW2s0OGrcsw+dO4+wT2rewm/LJURpPBCWpa/hbmodx4
6dA/A/ETd3GxI0NZvYSObAPhmHbn2AMlMyn+jOMJwaf+TrjOBGrwIvve0Aqdr1ZwhnohQDGTZy3X
aHYij+/0Hmky8scT3ow3U1Em/zzmduB9nHeKhY3PLA+Tu9XtEb5j4RpbCQEzkAsZ0jLDWy63JvF6
4C1dFVOfxLOkAHPfVooPkFq8THzexOfukinqjDnVd/XWT15DHTLh0+uigbFF2AHd4Z6PsjFpTwdN
ZKelEYQuOgNTCXjRXfjnjvwiAVLYONLLtcsLbhWjSBjn88Wjw2fRVPJgGsnQW9oN0HmR2Vl6ZFDt
KK21xMIUsW55zn4po7JZkYM4K14v8IYPx+Y7dFvNH09NfXsiI4mz/twryS3TU+Gdol3bn2m0fRM6
W7PZAdRz0Kd2oreuk1VxoDhKCjeUiBeqkINIJpc5w5W6kpMXtVnaDPidyp5NX5wzHYZNy4x5GZ+A
aivCgsKS7+m7f2lQYuxiZdrpq+ZDQaXcELSg2dNhn/EzeAvTrfYvDys7K4xiZtKiAzxOFWsjFvbL
ALdDAGcjIohYRgl0lSChWW4nRsWIGAYtmQ+JB8RRpDnVenl3WztMpIZ1d55yq9RSjTog9LI1uMsw
AMiescV6g8TCi5pcK8w6vVa/eO2Ze7MvVD9Mw81N9sK2FHfvPN9YesG//eiCMn989MFi/wiwXOnI
nY7P1SYtIof72y1AdilJjsEf2Diu7hZmaIhv3smI84UHzxyQFGEIlgHjSQXMSIu0qQ7qhYmrPMxg
xBfr7XL2OAwYtC/Y+Uy/VTjDVOgxLbe629pP0OtsexD/AHPSbvJ9gd8htVedB6K7OQDNjUFOpDVH
rodWCnS32EsWMN/cmBkRTwcBqZ7H2t8E+djDOY2OINRV7GQLeyMGIXPBUmFIubrK4MDOB7Xz/4AY
GmISjMToWGgjVSkdq8iV51+ObG6MEPiiS1nY20UKGuwrtyGghTOY7xt1QBPSzRmch52aZFo5czEi
7RSBdi9vk2Mka7w0b4f1+6zLG95rRHZPKC12rtkKkTI2b1RjA7tcSbB2Vic57EC6dTzLhKu876Ps
cmXIU3g+MDQO0qmpDRjBwzP7y2XHEvtIS4ep74UiDWvHRErzB5tKZsnhjxtnbixZ//jeogImgZ3I
4ZsDZKs+tqw9XGEaoJLj2f1JjB3yhsGHInECehMpssD0ELdnqpLGSLWYBtW23IA+2glEwvAgTPAD
mhkSHvGrerESdyf8PWB8VR+yD/YhzV1cFCScisBV1Q5vgXZZUXbvF29Hnxr5t4gwINi76UAZaaMg
mGALVahVHHA3kii0GvVep/IBlwmzHim/EI/Hgtn0Pwj9xFQTNUvsfP3x1fyMde2fkQZwmKQ+S/IE
pEzl37x4iXpbOvW472BT5aZ6wvOMYhoKTS00/BIMam5mJm8kwY7lInnd5kYE6qltZDPIvenry6v8
YMziSRZANASd6w/GNEeWDr6dHssttTz3YiB/oix/o+fD9n6XrN+ebZlZ+JZDZym8x+rL7GaevWAW
tLeLg3aEHShBStQ8ithGiLVfVM9V5q8ZoyPbHFrp/YdDanKGNm1YXVuxH10q4NF/gq6xiTnthNzT
BVTnB68fjVOUW3nazz/pFgtJA1u6P5426W7RPo6H7qW+r3fqDK19ZKZHACEWA8ksMw9m5Z7Gfjq5
fkD4v6rKMYdJvH5kfSC798yszH5YwYbJUMPdWHpGxiJhbSTBQZkHuaY2EkvmyDerX/SuJe+pTdOC
wXT/RejKCokoPnA9M3szHBq0o31j9uXDnXY3M8AplrESTFyZ992yDyX2dy73tS6LEU8kt7OyZQkT
pw7K3Nk9TB1Wae10473gSRqSF3ZJ9GUeTJsLVkUpVQBPsjD6jx4X/oDDMkUMJbhMyxNpPm+4ye3z
SSfpwLJCSZaEtb8RVH0sq3RY9RCi/3L/hdyUOh2slt5co/oi+BzmnLASo9uN8Fqmemwe201h/VMa
cqjEq5RIdwDY46vVWWjXP5hpWUVaqulJZMplScX51tPt2eFumDKLORBH4g+0Q3EfF1hjX96ZjRUz
f2BHimsK2HISNxwW+Kp3+9DVH2gNhDVHuRPXPXtW9MWGJD6ridMRJ9PgiZBOms6aIsTfbo3wW/SQ
eSn9kJVU4WvQc3ctoIYxsp1kF+fwiCCWs0iWSvVWDJq4bdC+pdFVntV2sbE3AxlqLAWVFhKnyw2l
dHCIxkO8jtMXOimT4g4+f4NPxcpmnAnY/vs5Lnrmm00sLuJ6JAf0kyBxmpZV4S7Unyn3REFdf4mW
hesw1fJQjTUxxBeuPbLCCmhCRvzMpZrQ04ejypqD9Y/tTHLhowI3l+CeO+mT9ii0Agq53ojtgT87
CAgksRBYK8NjrhctlEaiD03csaIFORpPIa2LmhXpbNxY1yv+3f+y8aWoxLRWWy1SgDK6r/II/Wnu
LD7PAuvOw9Kq2yZpiTHRXrGopJMlYqHGIb5/RrPZ/OEqOlcY4EcjLGiuVOpwo9YC3zqVnTC3kfao
J4j7ifwyBruhBdkK3tani62P77rVKjUKKb+37jVM6GG2RyeZ/v0HrW/aWzRg6aEH3/vDoxZY1C21
RxTFYTO2RC4ckwS6T66laNn45e9eG1EcEegEzZmbV1g7WrIdIS4jEtmEn97Bt3Wo0a4BmmnuoIcK
wvYB48ewySbNSCkSFc7d1UZbpjYxMc9mTWdO5HsDjsrnaxJAyNUQvdJhtcs7m0ZuL94u9m0kh0MF
Ax/zagoiiGa5iiW8CEprdEbhw8hPQr/0P95h3oZ5Pj+87ft/dR+xpeEPn6G9XpB9nd3JUlVOoFxS
Yl91aaS+52kb3x2OoZEcLm2Q7C1WjvrT6CnelG92ukgd4SV2bb1BK3ofGdgSbQloeLfjDp9clTIM
/VejndGxh+fOCB0yEqmhkZR+n0lE1nL7Pi4scV+660ErRMPYT4v89b1vk+q6e5RfyMfNy2FZ7dlt
k1KlYYSJLSmmh8VtT151kao4XCpy6Ty9geLnB8uBuV+YhezcHYKNZTYf+Qv86H2smlCksnbGgCyv
LrgVCwcjJkev1A2M5G+ybofAIOVMh1oY5H3MXjNuFQN+GdEbGWfYEBRgOQ3Hl49806kFRdj5wtu5
xs+dTK9fM/EkiKh3I3Noy1LNJG5JRhcnxrv51tmshz1/C3snhV8B30ce5ISkwdPqLVxZnoLWPvnt
VdpQfD6cln/pVGeQe4d34JewpYzSlTX4tnu9fZRlk4k6whVY70T81r69dDcUPZan5GkALNtqOQI7
7RUCHFUJbNc6E/0Fyep5X5A/6nJkjimO73N6kgHauchKizS2oZiSNAm8F7rmkzX29OqeldqKsyrA
q4ypfy6asdwjt7flJedaeRjf6mgQ6qsDkKLzNMazG+VK/Pt9xw3rpOTpZN90+obO4V5O1WGueP5G
jxeN4gmWZeIfOlVwr6BLOeLMComb8HjGrjjbrZgeoeRCKYy8bDINCB7GQikl7zkfWPN/Tvtb2qqo
+95NknrMT6Tkgf+BEX62gp8iNBqmYZQiYTNu6Kw+3/54ZB+HwvhqQ8DaQ+MIHIgIKjxJpRj42EYL
B5cp+qvqn48jxyfJs1Hi3uF+PZPJ137TaU2/eAtB10RTT+bIq5oAycAxzsVF9wT29u7kEMas400f
B6q7XxQ4XXmKINnGiXsN+q3r8Wh/6xw6zHiAp6KbhEpvIykKJiyqFCXZwJm0ZYJVksrJ0i1kwm+8
TQZAMl2Y1CPy+W3FdkBOdXRLaWT6wDiMRGAWtSaATTpK4a8V1RjuReXs8kDbykB41N7WN43sfG7t
bLowM42rARul4Rtmq/qykgJsq8qTRW0+ux822JYm/Pu1u+gp1fqi6zQXCxbssmAiGIMDp+1KqsCm
kvBaUD0RDl+6Bxjs3wAxyeDf1T+MouVoHmkwTo5VPENQYzLZbdma1GnixzkdZhAgU4/Qb5O4btEB
nzWvdDCARmxtRWUx0+c3+aDAHe5Dj/6rcocjVZC1vbMpvzcD1+DwQe4hPFc7NCj0vbOLFV7JnFXX
RdAK493Kregp+ZDKIrlUW9H7j8JgHnKKyq24GTU47GwoTZp79Gogtv6oXJCaYCEJ1I8Y9QOM9x5X
jG1mD4z595mgrewUH2KdsTXKtxgko20dvYL5f2mr9+u/JMfVhWAu8X2XbrPX00iOMazou7dQ+AxP
SiMT0Nk2HvCh9/ERO+QxiN1LK8ba6ed116QN+Ri/d/KAVzDZ/zSV1PM4feu7opSc414wp9B+4HmY
rRFhf4SXmiQ0aOYt1c/3UlI5Tk/tiV6F9m2QZzE0nzTkaXb2fH00sczXs7BMlVHP0FQ58sksOguw
IjItVW/pNJWteaF8s+MaXyGwSoeOmg/xXY37btN9Sn1kETfWyB6ULiSbNwxQOZVCKf66fbo4JuUY
mJ7iOPDAEv7E9m2SAjAjg/halBbekjBPnmrrWyAbH61Da4OeO8kxgPpb8ozFzJjq1sbRke2pOdSV
kXiC2pPUKSiXxENnQzOPVjXdVzrcfuKG56L5EmIHtzEqqfbxCwMdubViAhcOFoP+xzITT0lRUCEE
0lDlGRDQcdd3lYIJ3wlGjsP5Uo7sLMUuw+6Icw0fwjeKtSgMpp08SncaBlVf81xs/3VPT/JklFHm
j3q/UjyqqCPGZu4qVrITtiyq3IONM70H/DQdRHwbnfPHPiMQq1idXbJ1XK2Aa34JYrlbiuA1cMsO
oCIu6/tYgqRAxr53g96jd/2Xis9Z6GSrwCmZvPIo0dwFueTGHLR+J0i2ai7d+taZoZa1tj3/q1iR
/75kftbaBsdHrKXhhSs/k8617d6c/lfC6LCLN5QY7xao28wB5JQbxIQC70AnLCJ5nmBVgZRoq10Z
OD+qApVxNJjKhx5dgIECAyoIilywZlaoGymOzrO2qK/RmB+MR0vMfH1oUh0I+4L7kgvOdELMuXvp
UXEV7gv7Z/Po6EpvwwH/785u/3z3mkRjaj1DPUTSde+WQjjAH9QZ78T/GuyR71VvUVk02ux52hmD
TfitKc9WLlEJJhP4L1dc3J6OJ66MIoZzb8JnKrjMhUbL3dUyMrqUX5+M7BC6G/6yhuPJ7j+TrCeq
3pJ0T1q9axdBYplqihhVYTeQNXdXpJDSn4zmaHyMURepozRgohyDES7IDkO+QBeWXE2/YdqUVGzW
Ued0hif+FqhFN1bOhfi0KBTeQqJJnGW3v2CkVHqrNkeiMDqSVgy714Biux1UXn9V3AyA+/MyB2tE
sSVNZ8rp4YJTcyH3ETKSNChhsrJIRGM4avKJJK31PKaVU6IAlvYylwC7LbDEBi80Wh6YN9ycgQXP
VBHIxwJDu8p/xrjn1OWKmwNAOc7Fzc5j2yDx0V2uc3iKs904cdyJJ+MThobI/XbBSak5QGcXCVIA
dFtwns00tlI0dIUTrkuAR/964tuvgYyJzP24BVPsz7IeZXAkboCceflIIs4t7f1AdsuvGV6TkuaE
DNPzMyIXF21svCj76VPC/buInI9WerNwCeLCoKBgKe3JOGCVjWe9UAO0Pxh5G0ExjoDY1lm6tpv/
Y8sbouGAqDeaL0SafERAXlNSPbvmZKVv6Xyiox5FSFgdFwFyXcAbxK1+jRFJRPbkQOtxz3m/JDtd
8N83qD2cnHlSigQI7y3ODFbDdqq0a/AkBBFn1FAfXLAsGe4Miwghplt7DVtkOTWT7cGH0uPBjnY5
1AObdSAgmedOAzSAJz6YRtvEHr8MKxIQ5k2oWjMEEeNwhh+CmyjSAyOsYzA7UOPf3L6ilIZTtmcS
eEvKpykvjgjAbMbdyTGiRT+6px91vU2Atj0ACVYJhuxVdVDvSUgGESQ3klVJWoV4yhBQUqK08JbP
8dSwMaVwBD+hCEonS+wDQJT6rJnfYUHRqwm8zCp4fJlu90H3R3Z6Jx9402zlMCTReo0vTdprFD0i
voj5ohmHQHJrkK16vuBlNQTownM4SaIyEFZ6JxaCo8UFoD+nzLwAuoBRA1grgGCkBF45yNfzshGi
TRcOheY0D7PnBdTf+7CVkBRfGp5giUzqLK6bxe3ykAA0WX+UtuZSfBhK+olc63s+pHfdSnM43sjm
mvQbne9zXTkSUoYzZ1VCXBZqFwTYIzMHiEHn5SH/fEYjFzTv8g3ZiNSIiQlyqguqGjO9LTYAmIm1
kUELUITCNNdV9ba77Ap7jBb0A4U2BfT/f59sTokowBrusSYFrW0+ChVQyMFG9XFmSWH4lDMR+aBc
tA2uae/H2/zDbeofCUnRnaVGHQrtfB5lp9w3VJPXaeNmNaoi6PaneXSdgVkj+IflKx7K0sdO8N7L
AYtcYRZblN8AfWYhmYSMwFub98my/Yv2vYEAK3Gj24mpcxgysjJNfdvp96iQllmhLnEcWad8XVYA
j5BpzNT4FoNJDy3CYrN5GywPQTnqs0DvnqJRc0iP44oi055tCaS63ot6KO/1FRy0uNs8B4KOE1p/
LhWoCGWdC5+9KcUtpf3PZiAVIWrG7cvsPJHRQEz5L5AzmTAeds86DWXNdyWlXuRZSWWa43rz0b2U
926JDT2MmITVfhcs1450oBbCYxznEsCBTVlKKWhJeqdH9LmIi4FmD3aGRlskYB8QIjfVCQIer5HS
iacYPTO0vVUffPryZbjZQA26VtkaM4AKkCkBKwuk5eUMtj2XCXLDqZm+2hP271ScaUoPgrF4ktmE
4T6lfLBwn7SDE/Y/AQCMZ+70eJaCtDZr833OmQykST4B83mzxgvXPTjfXSvo88+O97MHM7RMtIh6
nqO6x1tjhB1yaRq6Yrwr4voxOIvQ/C79WS5VbXatuBgylFRk4op2mkYDvw2X4TzvBecOypn+DHu+
/yOYZ7Tw7qMzcJuOlq3z7apKiTD3Cte0tSa2XuVh6vkmqkJmG876tByjeTiUhOBPQgMMss3weMeg
RTdLkO4NzSFmjLOkCisjj6FgymWkP89+7ygzn7XEpt42gwjwxFQwfONAqfuHssPVXj2Pmr+1aLs8
vCbr8ux//FGoiHEiXY6emJ2PcSnUqx5pKl0fkUPon65N6Nex9Kuhrzg8KzHa6DZk+z4pHaEHkMB5
EtUqfmDYYc9iaOz9jryMRUaU/AMKCx/8MRfe4UWxK9P6JTIHNj4P3hNgmmUTN8nHnxloYphb0KS/
Jmda2BOV+Hk56uC/qF+AwTqfxIIEMaIZaF2DlhKbmV4sr2p9VHIPr2fgH8+SPiSH5AAnjLfs1VBx
+z1dslWZ9lBIXqn6n/ZkalJ6QDh88pEOUh7I22icclH7PdyMUarYHhLKOsTSfvQ7hIGI/cUz1mEW
wpiLdzEIcUUw5ASbzDBd5H7SPLG5N8Nj7c50yBYBTJg9MxbCHhGlG4dQIAxOcfRh1K1j9xUjffb5
mdapAcb/LTSHIXGZm+d7Dv57JNDh3CPL/tJ2oPE7GyiyIIw4PInkShMR2bq/IfJTcgoJ/sqYOAbM
JzMoV+vZMLKq8ZQ1aua1nZxjugaHkuwFZGdxBIcWB4Dn1pjwGEmDJcPQdUWcJx5kYugciyGGRJKn
tiCqXcwSA+RxSpxWDQkaclzghjetG/Q2s4wDgc9cJUfGlUNRNh1NSxZyscb1HJAsFSioDCSgiQkW
AaMJe3QieeVjwnxNG+6AQJWhdg7DUtgXgEO6GmKdb1rtA6C599gm2ARSiAi7TxTIrjV59UWDr6+k
+ZkzXjwkkb9aRLIuXyQ45nINJ6Hi/kVKnfhHwBJ/Wdh0RBJPfRJoYOxIRssGYiGtBElgXH5q5izR
jI3ijPX4Hc9lSNyvFr6YroOuatc5sp4/WmyrEK93b2735iIRD086SMXa9ltsBd2l7koISfE/f1pb
3T6Ap7G8BaWoSsjrLtdSiuzc89uYR644oBL1Wsv/+bccGAgAs61CGxsSYWePZIhJC0baq8VWprGM
mHAhtxJBl2EenmRF6yk0B1oCKS8FEtiKLxQMmHGFOzOD0LN6mcJUwHKsCO0FtI6DrkWGWHXel0BF
RAOuyvKIBX0a9/jGqY7VHSVEzPik+utnwPbEpYQXy42PLaeOpHdAlyLHCY+MLblK57oBpiZEkRRN
jj7z/TaKVfNLdTHPaGHg/6iyseRoSwbYZzgdtvQ4rDZeM41qXhlIsCvCUKA62Bz4PYs8Abs/MSoq
vWiZ+JWN+6YvyQD4SJWoOMKOe4uTbcjZr0/znxWWohl2kXQNfqbHR+aZPBjIXp34uXL0ytqMa5FD
CQX37f0Qh1iOvjN4Ia9OhnUIrNBLg/mP/KCWuoreRfZO12g28qUIUPPZipWvLkGBmm52MCzL+hqY
Qd8DH8DivcIJiqSoFghPNWfgm2BZPIlBUmxKzCtDOqdhdE8JrPqnXKo24w5ZWVuUEM4ZUvmLLlqX
HxZCyIKaZ5I17GgxSPNxLMWoIKoKEPWbtA0bP8ZMtUphkVOCu25ZEbzkaOitlvuLVJbu9Yh0qcSe
IvV19A6D5zlPtDJ0VCkQ4nIR73Lkg+V3ZiiZt79Nc34QcrwICyaFtd1K2jub5Ots6WQOHLOGtWPs
3CYrf50aXRql1ChG/C31d3RlEgxxRniswyLjovsly1McoricSM9LdnJBcpADn3iCLNK7dyN4E9oe
fKOxOThzUHDDSb5roRZGPO1a1l6ixEowSQWKs3Tay1OAMwNaTuqsragMNyOlTopxVg/kdR+6pJix
xFKiWjkce/wWrIdJ8kzykRZbwIY3cPvahDpevcjiRLNW+J2X4Ycn6D5y8pfeVVvm+MP2aZa4GMZM
Tz3fsjR0u9l8YO98sI+rRBkNe6Wz9pLitmxk1cPe1hCiM/AZiAsYwpAPCCuBuqGA/KvR2iiWLtAJ
B4SHmUHUynLSHztGB/V2dZtsFeGCb4AybPHZvHTDDkKFnp9usZzrr2vW6j5dVShjQGDudxaexavO
KwrD4Z8/0n7l7D7OA9iUEYwe1JfmPwfr8+jdU0A36NnY8HvaukeF/yKbJKZvo2KO+gd2BEwdDP0v
0siCAXcnwmBgLSccw38WT84NKNQ6wylPcAIWNAmbIr1f0sq4dLY+Uv2rmhVPdqSaT5m7i5Fm9Cqz
534CQAyaeKfLSZaFcC8Rwwdomvyq4YBJSVD0hpG/A1AMk4lmPHm7J9B/xUzlWD8x1xJMYcd/bCVV
eb3f3nYADx4r4l/3XSvf0PLAUCyA/QqhHVOuR4l1HtBeVcutMlJiFT5a6DMDbp1UCEDNBrc+hFi3
bPAJzuwONwUpW/HprsZbEv12BZCf5pbN1aPnJieKyIpKJ2wBMM20nLPFTh5T6K3ON5C/qBqVF2zV
vohHV7S+0ZPoMNSCO2X9mrAgd3KA42CM1ZCMunojqK+hm8xYkVjByitejBY2W0Bh9P+JwRG+vwAb
CmEz/66+kWyaQkA6pt/Jzsi8c2xFwnqlu0UPJEHMli3bHqxLuQvuzmgWR4o8Ok4EsYOQ825LEXO/
X7rvEMlLubEqPKtowGuiOLMNqlEp/A0A2A/pyXFGjaIyRnZAO/8w2SKmuK8Tj4Y2M2vyaiVAcvV9
9VPtftXH5qFqTIkuT8RFbG9xFochPH5BkA47JWfBCTAMsFIAPpfjZzN7qD0Z47PnuirbKda+iLHZ
94wIcI+IyM/JAW31EXXTqktrtl0lb1sbdNbL4qiHCcoYdGzLt2R8bzvGnBHLdto8sVAYl2Ao7Hye
j7aWZVxqAHfL4Wf9xnI1yv4gh9EwTOlvCWoYTy1uD+okfXFhJ4SupJZY6dbRkKWHv49627bConoe
ve6D01MmmWbDZU8TBToQaaqGiacuJQLGcPhidtqHGQqdXCffzcdlnzpMHciAYyxr1RNlrARZK+Bb
rYdrWrUBMyhVjF20JMzFwozLtGkcqF3HQEtWFGKZIuJ6DKdzReiV8eOIRpOzkEtyFDynTEGxbsDT
q9LnUZlKklt/3smPCdXWXTRxrKsDhr3/UZBrnvC5JcdU4nKxNh52tRSMtQ/jZOxi5TbZycRLxLre
g6ew5X6TkOsRGH2OZlWrBsA3lhnsWbEZxR9MzTkZweXlG18v0w+s3gENL53cIQjpb+1Es3o3kxhj
8E4Nyfxss0ZLOLPGJ3/HxZkA30oS9eTMDaEbln59Zly8WLedgE7vKGKSjRvuD9xThOpn5pX63vrr
IQdaTOkcwc5u4+wlZ4qe52WXQUEMbBBlDM/g2wCmMgZD5bPXtmcDulopTmjkkDEL946kwqenletT
5C4wuD2wiXTThbMhF/vtWzZn7QndVhEIrOKwbo+XUVlz2zDnfyfEkPOwjmyRb5qGzJOWX3Luybar
Lircl1ISAwf56oDtvn80zIXL39P7QKyB0Hfcl105E0LMB98swh5YxxG8Tjc0ehWss5zt/9F6u7d9
PBe+C1S7wYvC4aPUl7MrUdtVCVgB942eKTTBjlQ/qZuwNDdVVKIOSnPc9BoWTy5GbnL4wdeg7cjm
qDKWsa85FsMF1kjV95jkyVqRM+LglrGLOTwJW6zyMMY5uKQrRKWG2PAXAy1okW6Wnvpqk+4Lx7Ge
6HydMfApPod05Qf605oVwuYQUV6nuT1oQ0An4rmCm2/XR+hLfborgrdzUJxi/FXOX/3dkS3rVgcp
yO52PigRvuvYWKtglNX6wkIZXQSz4qTwaEeHsQ+m69XPSlzj0ZvBUGuvXVhwSCuRMcJz4dG2rHFA
6G4xGYeJW6NzfypHzmk/FO8TbCCLKeg0NSj11wwqUKD6Zuu7UtoZ9sk5zQChiVv0r9SvDyQG18K1
upMRi8IhMWVmAFiLVDp4hpNa4oi8anoNXhFWL4+3u5zqmB7ExF2FZdHkkEUvBgkIa/TSV9EsXXIs
z7a2z8MtVwkLOqkfr6wznGmVy4k5a8V5k2D3SkyJulJSoN21pfhSrXDroX+Tc6NLlBkvhxliMLpL
ILYiYGb62VW/8Tk5tgbW93EMyGHeGIB79Waawj8kkJ0BTn6HUEyj5HUXWpzkbnXlDaELRy+ZG6YA
+BkU9eZYxdi9XLKmUT+/8PwsAc8PyUEYyyQid5TvqUEMuRDuPlP9Jz6UMINPKwt6Ru95rPES+UZe
AornJa8T/OAg3yRvjp6vZt7Ys4it7K5P6AHbW1PL8mqO+OlXK36L5Zl6vEtwU08Ssryp+a5LpGVB
NVvv+HgzcFM7YjozzO27H206p9SNxkOCzLB36EsjiAdXWhPibszWakHDFOhf+mX8AU0PEfQMqnfx
KuzARmAbMvyVHWqBPztFB2hqFylmYDWUvUGuL613cKRixgajaGMEOUzH4fr2uBRhcFClHLEdI6mA
xq+dRr0SDdXaljnTe5PPL4uwt9JtkW9Eb/sfwuiAcWcUKv2BcFBC5ht6nrnkJKhfftj2NAKIcmZO
orkYy90veSlbrS+XgpPMcrs/xEJAQEmAV/iL+aJmoLDHbtN92cMhbGxnjzz/pbmSlxr8T27swt65
QOwM3RFJJUq/adbmD4sx2JhtLZ1NlcLr00+lCTTO4boQNaBEiq74Tqb5ZOL/Jlv29z6/iQMKHLli
PR9nW5CRC2AqNyecxs7Ldfe1/0VhpNoBPPP3hiHUs4nJSimo4cP9npk5T+86/hFWDZ5XkmWVGOuY
NMXyZj5TvjjnCchWK1x8ZesZlNWs6WQEsMuI2gjenfnYpZo9CimaOmZnb19gF5vwN4uKn8kTy9aM
A5GgcX8l5Cbe4TNoMZPecYat4TfBsw8QyumYvNoHxgqEdmDzv4jwSFd+4VcLg6ie+PAChd4OJsq5
b+8Ug4X0Q+q5Qnpo9AFnQ1lYqoCVDqp3AMJn4bGmEbEw6S/Pg2wsrozDUPg2jO20TdPjLbdMwD6q
efpsahu8I9yraSDdtttv1zIGwjMAOVHmo4zGVX4eC7prmccDfDBmb5bfzG1fo8H197NksOMAFJo3
PoyA9n/dlGwAWmypxX+abXDBB1djNHgYbtHE4ydr1qGjUFtRup9JjJF0//a62pJ9b0W98QNkx629
dhF4u5ZAG6+T/0rinLG44EeD6DpnjLOXrd2bDMp/v2A6+xE6cqhJVjX8vFkRNfOGAH8kllRW5LZD
199mVzvSoWg3tPjHZUlvwZhlvObRM9S+7w62XOulqlnODPehya8uF26UZXp/kzl/9rhT1UlxgZU9
JD0shVN3R6dWdZmL/FNu0ZvuRyxqkezsa7MXsvci/ObeSYwIuzcF4l13keSBzbZ0eEFCrDJ+gtKI
8nUYGdoochv6v3hZ+BD0taE1ZcnC8nNMDzi4W8+MgptnjlOoP7JBPf4jJIXZ4CPXsZN7jV1cwmok
zgIJzvvJLLQoRgSdR0bnv1dldcX9ILFm9drscr9xq7v4Y4rik5vG0gor/rlqiTBKkvJwYIWKVt2D
BXBg5q+oBwsgQ1g/s7ml0pmwypSQcmGU8Rye/dEFzfQ8mcBvjwE6uH+DS6uAKJcevtc6c4FfJTgY
3oJ1MHlCWupUM7cEbfmEjrjXkJ2EqJGZ8MJqm1W5kvbUIz+2eBLWJ8QvTum6mERVsRYRF5WQFsEL
3sKEPxy4ZSr7Wwd94l+vWNKq5oTOmgz1i5qQSoFbX352ZkIOWt+MDHqBOr5i+3XfKOQIBuYOJmjs
x8Lxse6+ySof625+XUXTc2GsPePdfdbOA30mtIZHKUQKROKuKG1QqRQ/BMGoZNHTNX19l4VoS18V
KGGfY03Jr1lZ/iKD7O71zu/RGOmt9iD+hKbDHIQUsd6mssnpfLSM/5hmZpF4hrR4hYM6zchjVUmK
8L/0iUQ3yCTcLylXXwF6YUyf0XJqLsOLkHKcZPWwVF+GWsavwN8TBQDAgyExt8UaUZCEZsZV1HzM
oYhwpKnGiPFgzJTZAMwu4RvBj9Bb6P9TUBqPdqtIj+H0uJto8xZOL8GapL2bYr+SM46M8eFYlZKf
QGzJ2MD/foIiYuWT8nZrLoKg27z+b+NvDFKP+fJrxwInnxmJrulLq8rHV2V9vEKKd2h73XH4xuAE
uRlRT+StSqZDMH7kB6wiaHRctbgghN4msqGrHj8viiuseJPtJ6ps0qVHrnmZLeM0gwjhF1gTJUi8
XOMI8+CMaKEpo9TnYHdbFHHmOTb/KEQYgPAdDYSReuA3rHvdmSMF898jmYIEH+13nKMxn/WymM1/
t3/cEhr7g6/9zfGmxMwOcZPcEtqpY+ja6YWPVY5xnT6C1yLBebEXHYDm1koaL7fQIjGzQaoXVulr
d9plZUMvxk1OhorU4unk7o6d1RZil8msW+TKmlMKHQRGlR1uzyArkk6uWRcG9aBCXHAWYMG+4LAP
Uaf3QIym1E+NLbxCKhmvFAzdkrqMVwsycwUn6jup+DG8UNoKm50L9XBcutv4VMLSmI0WHSA5O9nM
C+/2/1fjpZt38epxRML0g+vIhwvb7qSi1GdT8wm1iq6mFWrbDbm/k+EzR3BjluxmnCPs+55T03qG
lRWq+SIJRhY5K/YWIX6M2o6CcZ4VyeNgXsAP/7yGlFTEpdgAs6/UVlrm5qYFHDVZKSkCBd0wpm5Z
TYX1Lu7D4Flo5jRwJP6jXJNHmH+VCVkPq2iRVcxSnXS1iT4/HXMMybyNUg33p1FrdLSUcMciHuG0
reGpYDaXSkU/KxIPs+9e2BBaq2/4aSDBwqgsD95FufqzPhGoPhXy6bnFtOsFiqWfWjNBVwk8ZpAd
nicC+zc9JcOTNWf03J+rqXTXPciGsSZJD3K2FYhz/+tA8HMNqjN1b1IzwLkVELuTMo7qzmqj7iN2
WM6YWUbJ/5yxQ2xbawyTo9HAsW3U3lIWwYwdKzpBWn30z7d70rx7W5te9oJj2SV3c25KVTw4HbUb
bnmLtHnqY+46Sjin+wjlM7sTG38UEDsavn+Cnh0x15HcVlnWgtJ4tugGf534trHAv+ykoEx6pOnO
QHWr4wcNd1c7vKwKSzR42rlxFnceLMFXxSvYcIli/ZXQkwVt0i3OBmVgP137CDc/N4HpApiOc65p
AadbpnhUDZzfKGEkFKQlheoDZssap00plh6utPiZOhTj+nqhR2SlOCpdR9FEtEvOXIbCJm/lrYFj
/YQYtsjHPtvWvJbikT8EH2TOzbJva0wf/9MrKxtLw15wABKTS6O6xfMjHg3NvT+yLv5XrxHpO/8n
ZqOGisVevHKwFcTt8aTI59DucGqv7LQfZMDL4Ce1rLf65/trCTSKZMse4qh732hH33yyNo2ogadI
hXHF+/35VI+J+qF8a6JMeR9UyciqKLteZN//oPjYgnvW42Z+fgSvIo+EVsYuWXUrBVGljC1l8jRF
CBKgTtjfbxR/P10ILgwUtyZQ6fjyFW4wcmd31oyaVKJibxuzW2j06YRu8t4zg/AwQQfCh8kKlXDD
z62LWwQK+CnCPKfGrC8Y+O5CgRGnCEdAVgn6Xt2ckO2UxXs1dWi7i5Oz/6+PVqSa1eT9LifKXWqv
IiTiS85v3ltE9jJUJY7ARQqXk9BAJeUmOwATIbslH8DGDxKzH/Zd1eYU2soFrmSdFPiTBWxifgwn
taHuiSXr9wovNE14VSxUocmfl8mkyZZiEK2iGoQjQ6/O0l/zj7OiGJAIRX0NOq7qQSEDQkfo4Shx
zV6XXPOIf0at5XXbyon3yMYCCTCuJfxyuSI/xLKX6QoEnnSXuVHUs1joUNzVBhYZcQfko4fn0zTv
sgZp4CKNG3CZ9bTXXNb5ktqQ0QhwQrSCMGkn5OGeV/ClVHbmprQQmCiIwQPy/Ub5+EtILzqC9TUt
wnMfMPTDOFpPPBB/fWndqVYXkS20uOTwkDk6l2GGEbZVMh5pHvzxKeZ57lYXKBCkoQQTPR8oEStw
e8aOFAh31imWbz1bx/fU9dsJJdjkgpoKAN2WJm2kQAy5+mISh/MgXT0RIgz05C+u0BA2JKbDrNCs
baxomJsZ5lm/wQ22fMrAtWyuvDfNrvaLMqd01BEpFv0K/bFPPiDGfrZOpamCldhx+9hy/13oVwfp
eD+83uScLfVRm/1Flof9HlSRgdjrUyKAmzqfs5Rd7RtTDN8Orx8qhNyQqTw7apaToL1+F4/NTQMq
JMRQGRc+jYDhATelIb0Hu8Kq5pKGT2YIpU59zbP69gChgyVI8e19MIED+BoITU8VimsviEoFgT2R
QcDhuk0DqsE/l2xZzjnSQOi7G/KzhtfNl8d+xnReeOzeLvHa1P2Rrds8ocJU52pdgS5g0Zhz+rDf
OPBRB5XSRZBa5Y/qEhWAfQb2XJ8S2pKHkkNVngXXB5QCi9fMBtNsiPjLOdkT1sL09o/JtMj2RHJZ
8P1DCLohsh3tE1VZTWjrhpPPndn2yCCejkYpJox5PHQcYdWipoZQMFGS9Z0Ft3XmGNzeBxL4kwjI
yq+t+MQBUfUYFbmTfbD+kdTow6vT07dequfyaBqcVb325pYU/1u2t/Jr1IROTl6frIbjVBUdQJT0
7muklk0hMGbUc6rMNpAk7m5ZiUDHmDPC2pZfqlsL5RPyQJRdXLmfg125nluISaGUvfkcVgmbXPFu
i4cc57EoJY4V+oJCt5BYUWeNsOJsoxTIW4DE3TmrkW2a5ShUHBCroZJ8o96eeNV8Q0zUGHQDiHdL
UfA/GVeSNTV3LQENYibU3LxEi/bSmVR/gRjqV/0w8XmuRehpofssue7iEoRs/1tkTGQcdQMuEaW9
gMGi5Usn6VZjHZgWWP9DX04kosZF/JIhEKohmRSNBDM/FrQMp9W6y2Y8TgSq1TwlI6HZoj302p+K
21UDpwYL4HwHwiMS67felosEWwXkgmOluGhAQj22iL0Niow5l3WHFPwO83JOaGmfjuWlbbdDEeo7
mJkhdip3RhbWuHUtjihIid3yEcO1SUhE+byo33urnPa6xfoRI0OppOnjoyTrEFAfHunUMWyqx7RN
bngUPFClNriXtNFWdJRJEznZvIjKvnUWhoMl6OysIJpA6si+arRpoN2XEz/ImBRWlrYejVlxgZQG
g0v6M6KZSt2VAs/tpVBTrzSAYqggBseQ4czoypnJ8UvkkO8Ornuqu1zljozqd1Qb41DfNVdeNNPb
cLEd8P6ZyfTQo0SK5wzcxxUm3rtQqJqLxt3in3irHe2x+MnUS1folh79TD80Lw5RT5p+IYU4uZpm
lVUxDWbwo2sP8LH3OCSVBuG4sRuiNg9rrYAqy2WCWLVJDa3hiyvRSHuIFrpbFuIDy7upvxse4F3i
pjRVdJnE0rKyvW4hTPyJX3ULqRqncBREBHRbUk411PnqRk2AXC/yQ01Z5J4fHiuZLYGQY1GYZmmr
t/axkUP/LHS6GeizU2vf/JgCvxSFCC57uBxXoqlFRtlWYVsZdjieM2e+5Pnv9uWJG+nuDMXZyDSb
fvIgjyJuQEohRIqJud275WhuTIIrV1QVNuBTRX4sDwYYVoAVf2G9iW6h/K03qTNPkLhF9pNQlNj/
yyZvCSZwUOCgb2dcK8YtuDZ/tzO2BrKS/9xeiIARNna8etunKyBFJOElQL8xqA67CiQpz6BY6xZV
9S79ekpaY6Nwoq1vOPc/A0GFIHj4N75dp3810Q0zkaJSNikNU1heaoLyf33LZHreHHpBkVQ0JaOl
d2BECzhNWNbYj5YOM6TekQqqmwbY8ylgR6Q8MFmURu0XniNwMmKSeXAmKZRR2cl4tUaeXYso/arQ
nYkzCkh99XxKeEJCfc7NW2j3vd4GEXRnLymOt4IhsXn/N6a/v8hPEfXd6fyxH+CvgiF6tJaW4REQ
psSXJ3xh0wnC0jdKSghepUlNQPE0Q3vgptffhgPxd3e2KtTZfnil9j9Gy2/CE7tmDyHiUULp2EF/
/6NlDvpyROTk/BadTK2PC5G+Rd7sEDvZK9uuxLpaIxwr50kerJfRSwmb0x5lRC90AZwjlHHnpwj4
mvi5YGhOOIkeczuIjI4MlzvwFBTC2N9nLPAI1QbGtTJxlG3iQSg9LRaQRaqwnbj3L98r7Oxpp0qD
/U3TrrmYUYmH8+op4+L7Eybz8TUEcVFqPjsnmqlKnDODoxQ3ckyAE38HN26bxKwhaToEC+Nr9E4/
wXCW+Jqur5C0lrXuuMSLQmFthDj5JkJNcmm582Z77x+DPOdAepMwKfS94EES52wgoqNkTl3lo8hH
H5a7Z7+zFNDCrQVW0kpvyAp+GZakc5bNjqDGTHQRHJoKq5RBP/x3PsixPm5/YSuB6QqyKwiwr4Rr
BzOeBfluVE/qSKKvxpB7QCoUNF+k5lYN4NseNPw+TvLhDwZYNiWqPe0f74bG1MY3GiVZXnTiqNzR
5G6J3foxd8mJWPgqB17c6XMBb/aE6FkgQuYI36WvE8+XWXLDX0eV0wQaxhdgb4ga8PibIOc0sgN/
DfjrLMXyGSrl0Rx54VbzYUiAdeFmD2Mou9V7NjzvqLhyA9kZ9g5TtUcn1nkIj0/EaiJtV8yxmvGP
J/9l/WmzApCES5txbHmu+WCjaF9v5ZbpmXcsAi9FmcQWqIGBzi7Rz5BS1YC3soAE0zALa9erlnLq
+ltgJf0pQQpQsTlrhtCW+e/1uDPzAT60WiN202Lwm9upugzZciVUByKj0ouJ/gIg/e4zDhQsQ3ql
yh9jK0uzAkr2XR7DT2Sy/Ry3dlLihWwzuHLtJhZFMSw52Fh5q2o/dMYK9ZNv29VU1KgYewxzKNEM
dmPTGoDkupxL7Y09l9IYyq5QgqkR0A8DoZAE/6IQDEAM9R0bhRWlCD085DmUGWazamEWaOmn16W4
OqTn3DQxDcaRz0U4aOl0gSnogZ31dHfVyeSfEMViIydTOi/bcJt+4xhYYMGwAeI8JP3I3nbgWL8R
BU4/xvIG4C0GlpVTBF+n7qsQrztPE0yKmq0HDoQTr97zZ2io8nZowC6/tkJ3psq1RofhTf3p0m+l
EoBLenBU099/Bdm9vADpN8iJOo05JVeYMIzW5gaj9uMUPl7hu/SoGyBVaUpP4J2wBxwEfjcYFBB1
hVTRmhSKFeCyz0FUTL3t9cCn/NS3GLs4184zQY0SdCqo/y6JbsrmahSIl0rgw4bRUNS/uF9uayhr
OgWzg3cGy6JKLExaf0VZflPSVjS5VkaHWzOFe3dzeEKwpH4iVbLkh8vQedtkyovO37zq/sghfmxH
xneTslBItVxUEBfZgo2bTj/+qGizIMMKd3+VR2/iAQDPiXRIRibQ4dvguuxK16lLShh60pcd07Fr
iCoZDIIigsutGdo7Hu2EGfxYqpiTaFafqIUs9YqvFbA06/9UVs6BjYLNeS1s8bcLJed6e+ZHo6ke
Fw+M22I+ZF7N/1G8Fp1eocSCSERl3yImPMTkvaA+s72J1RlGMnYOCrkqBY1whOqQlqAju8LPRzHn
ql5RJJQ+HnWbU40reeye5KFwIN55vNXMVd3wmtKow1pompZDB62Uxx6iaB5p86nQDGidwPNKIWx5
KvE0l3dt9LM53CjvEqAumTs84q/c83rl/2SVMsq0gHfOUxnJJBhXcOZxYAvwGe4h74AvGlobyaVj
UHWNUbnOAmid7kehbUIltnYWoJoqEcJ6IQK9FC8Qk7OeTU07kTw3krEtAw/qGyWXYPzYWNMB8QcF
0K1tdGQjB3djw7uu5iszwW/jft3FJ3xCzRPSuETgNmsAl6jB3kWgjg1gI/GfW8PnVP43qjDkMg5D
wUNCRrF9NkQiRftkeNZr5mxQVLf5TzaS3RCxo+1iON5kqYrc9Giso1hOKEOmgk/sXctYqNvQKhil
umH3ikktX/8Psb7lh/XqododjisiK8XqOFGn0f239yLjcr/dHtYSgDNwaz6I38PDIPpEunBSdSnB
+WZ9MlucWmEL2lKGDpJvz2r4+coJliBNIyUtcD0rD43GFI204BpEsH4M6h6i9nPif4drYxhu/M18
XeHYn8Nl3lWl8JdWA0qBGdY1LM9W4WQPdfc7iP+FixU3wbNI3AuBxspfj7rw9OpvbX+MKIrcTWNr
oQp8Yt93RgOjNN0iWkn8uPkV7OHtBndixotZ/vaLkD2FAdSdNXGm6I51wQPPxha2mcQ9pGZHsUKG
prcSO5KuE9ZRvebicgpznh6o8rvabLGCCQN//CIEwKkumNSSAmP8P5Yxfr+SdKWk+C+H9XzE9JGp
OcSU3W2uLqN8UB1CXM+CIbJ7kNx89XNpCDRagzO+47C+OVxAIwFTr9yQUAt+fNFYv997+IgGVAco
pWr2ZVTHVoshfQzUiKAi3krE0WL91ZkLzv+poLevi3yAFDE5A/C1CNW2KK8h5kL3eXIIHGC5jcCi
4TV8ekqvwewYOCPGMPg3P35d8GWERlL3MSvH0vPbNCUWwyNk3Qg+iGzqLBvi9D+7uNCCVtDmLSuy
PslYOsh/hVVtpiNz6r33IASR9xh9lIVzU+h6s+nb4UKu+qWwkWj7nt+cFv57pgvP7CgAPp6bCAVP
/XJcPi//POpoHC4WjMptKGWzxVv9saD25MeZfl98KrV3M4/K/raORBkIArk0HSjJe+4z0D3ObBRD
5ymgLcNGE0xb0sBNPin890J2W8cNxG817+nhB/51CJAWwnih8Kc0pfQKoppFNH3OBzY7CUqvLLbw
vORLJEu9kssficezjc+4mLi9bGvdAnuuHImiZN57BwkJnjE9ZSWoFPpnGza0TapMGlZG7qpH3RoR
ym+Hj+xpWmxMQ7pHCqSyLyiz1KrLAFacrJxExJ4/k/BZowhb0f9Ot6TJWjp3g9k5viYoydejtyTy
xWNNRUjNsPZpTxYOW+ge6uplnrRBcJz1dIWd16PPh0lV05hjgY6bonc+Y6yOjgssrHEYogNv4nI1
uDXDBm5SWVoxaGnQ4IpkqSAv0nQW59hk8bFqc5oU6IOImvhHj5AT9pkCkBZkhFqVlnGoxS06PZxm
jZlMpNiD9F9QsJaV5WmEzexIpQjr6ON04Fus3E6hQx9u6GNTS0WpIR02rUp1KH1PJ0kvqgutI2vc
btTI8u37EBcpZ0TzZDKEA4DPplktmjYZX3i9q6n7/c6pAqUvZvJratQ5v32tfv6EeBwABN6xU2pv
G9JVx+IZSQav+EAg83pGlTgD3m0RZ987A7I88NTfJqJWdr0xk7hPePp81VQtif1lDohw7Htq2d9W
rMddHJZ0O92XmvN8+PXvN4YRK+J2lcoY41SPtR7uPsHzEv+QfH8So/eZa5qCtX3J8fCO4J776yRg
e2k0saoNuoO2usVQ8qD+loRjAnh7osmUfmW2/e6pDVi8K18WLl+L88MUkEzWwYWCe8QXkEXTfcAo
i5wBgp4Y2hzp4lFFPX8QCWr8bbRgZI6Q1nNWB4g/GSSfsYDbJPxhNzkvPN47YWPSDTBMRsyFhNom
1ajag7XtXzmbc/ogVBumSBfOWCqX+iOZnorwQ/Vho5Phw4C58xY3PF+C+XaZX7AdwzQg0hHPxNWW
qRXW/pxytvOah6CCeFtfJ7aZu+jvs8tf3huijGurHR364M3ovpilVcrzTAgFsIl7fs+F1Bzyhm3k
TF2Xr4RpSpxrzuSViZKWQuY/1uAJkZqtKgvr2YNEGoz5KmIO/Gv3GbRIRNNM2LzsQFYW9AD279u8
YwBgowx0069K3rYg68rMwq8eQ34KbcQO9FzzG4q6lpHXrJwg0q+SzkGdBLGAUnEdPiz2Zry6P/Ki
B0y+QX1ZyWXNnpHNCF77NoPeN+qSG6sOv82XaCXisePETKVixO6sCX/G7GQdDdqhgRLZ2S10/Lv6
6fmyGXPi9iETD12AtI0xKDWCFPkLjg41dIdZM2JBX/w4j2g3cpMmyYkWBuzdA6jRpBevJ7yStIn8
/N8zluNd6kny1KOWA/UogAGwEiLdIqZRMlCdjBCMqwhtX4Sq5vUiQvMPEL8K1t6Llpbyk+nonFbA
3m+GwjGqNlMb58ErJjN0Nov2S43hpBD34iDtWgeweBHIys7Iz9Bes5oNQtshAB0Xy4FQ6454QxW/
9zi4wwsHuSh7yKxam5/7WkYBjXtC+VGwJBA2KGOtkGwtpG6gD1koq01l7LAiwBHf3kLwZz908uBE
QMzDHvp2uUKT7vHWRNHxK6t8MUabsqd1deOGOZwqOREKJ05SScA7EyGFASa4dogxd94HZGbuPsQy
QV/qgeqj3s09XQY8VPQ0RZ3csQQUaJ0kOTo3Lh2BjTKnfKBzmR/wvXRsHdx6LDPLYXAofQdZJ9+b
V8jmNH5/G4iBFkAyVhhO1lVelVZxFb16G2IGI9T3OYqYJdV5pG/hya6QXh5Apfzy0BMGT420f6x7
x3pEePXSk7Tq53uVy2Inq1pQ6DcWFxUktvFXPmtK567mf0OznBodl6ra/nbVLb3H/f+5gPVy1oE+
08nekHmmQNzWc+T5y4C3QkSzOazNuR9MVKcFmUyzgdI9Es9Rqk4sCtN7I2G5oQHwqCctTyJ1/Olg
MyvO8f/jbvmbBJtt5hWjsjCPrRqJ2FgGYE21YrE90/IZn6gEErrNspuqN4bElWEDL1GL0LMXwVsz
1LlE+Axx2BDrV6Jqscv6vIwaIIJv2FeuBuml2ID1UZ7wYodTGwhtd0h4L/ECAs4Lvqjo75iewQoG
AlQQfwuNWzPqvPydwZnZ0Gcwtsq9HzfdBpOBQ5US/ws24pxiLObRrtBsdCUVMxGT/VLdkvR9EoAX
/HCS7t3rumLIEuzct4LsX7vq8zJpEHhz1jd7Dz6HvqmcMkK5MPt3IxSTZHRFg/BOGrtdPYZSIoOk
J8YtI7KLxBpDv9EtsgOeAKU92hCJDWILWs6mJ5dn/1QyMGJ3YTdwMKxm5CTNrtjBKDjfIqn7MaDM
yUxZcgkPy9UJ0WKl7EJsVSzjF7uiuBz/rQyJH/OgIFpEfHqXEdzxr+KjivlOqrQ1qDqkpc1V6hgW
2NAOZfg+a/k+DpozMzD9XiqUR6aRJ/5jVqAWmh0kcYzpv9R7aLonO6tJ29GpjrJEBjzD3jWZTPAs
AT6x3STeA7l1ACZ9+vOORSdn+Y7mC7BEDuBh51+fhneY8zjq1NkeOvWVxZYe8lmZp9mwCAoJdVlN
qGnFmFiOZ99QtcUNoePX7qEj5VV7jWS/DmVkTPJUKXhWL+JmjtEJvpRb0aHbX5Bnjo+try6aisfU
ZvBNnozrMLGZOWCu3i5fyWANekv5u6utj7rkQ5oaLW8JCvvpp82rc7+MD8DFW0DgPPPj95jcz/SQ
O44kEi1HqaShP4h9X7trEKsFm2TYzcQosaod8z7Khlp6wGc5U/GbicpAOxakOWA9xJ35Rs8sM+hU
/MCBAEU6ziEt+fj5OW3RpHJOHGkqYwRAl6qbfRpGl1wieaxSy8BZq279kGrSGlABQ3nVeBNn+wv/
KzJex8Ayzuuf3nCmayuhBsml+XaIsA2GiIf3zb8O8rinRD6PpL7jNGgOBdywTHPNTKdekzjaQ4de
5cJsxFapiyglFaxp1FizhldtvqXLM4HjGHv75Cq87WnJ7gRbxRQ/tiMPkU9SllwkZ6WE1kiZRtPg
9+Ir7TavIHoArMKWQOkKZxzFvso2VPtWDDasMliTqy75ZScQV1Bao9VzPvuzkPcnfn06tUejyN4P
6RVTJgrzfFRvImwv/nr8RbiMnmctjWohVv43yMKoQOaCiVdbDUhtZghdO0cJc9FY3FU2uXti3UJc
7DLT/uvIcJi2itI6OT7X6kjECGoxQuqQhiMdCtPTtdn0XFuUSMgfWGqOf4DRHSP2VcMekw7/48oc
Trq15A7pqnI+HAQPko1EZzaYAQ6o9XDMDWcv8wvAUFp/YIO5Eqj4bcA8S82CUgOF4LKuTqG85ZQr
BHuF4ext9mdf2LlVDqAFIV1PqwtXWNrPfBYcv2HGokNm6E3DG8ezOshALRF2bN3jRnA390H/M6bJ
+YdAi316TVrV3fePuMFgGyPffG5jRl7k4i9UyHM1S1sMKHZR0QSr0qPVx432Ij5ew18qJ3RzH+Z9
iTxtO5LgfG3D8WtYAtV6oKtPMDjAD1ipa6EFaaExGFJLVEOZXd9Op9HkRu8tGNWE3KpNYaCzAuXi
sGjJrfoy3utQWf5yDUFPyQdG/wNJhw2P5QqnDIUikzCBcK6wVqntSiT4O+fGHuWr6+RT0gY9sfGE
9GCEiyZj0RibHlmj5qAmc06LzJXvUYYtEFiEjl1pOJ7dvmm/9Mz1/tqf7dzMGCFShFr5L8/cfC9R
QSRDjHj0Dm9U/RE1zYOSrEJIt8aUrJJWvzHkCUu6Nk/jg7IrQCQS1VgBUj4hODlB6q5tb61Dt25Z
fkSlBuvkqCtTL1XmhUAEIRajfhuFKjULuJNm91EqFjH8vlkp2xLzXMJOPM0OHjUF+0eJPT6kcMrd
VufBuFNCDDW/COgOfVFkbHilNkYxXKcphwVvQYj3PcLfysqF0JrMK+xlX+ObI3DfFDY1QFc1vLxc
29kL3nZe4Zj+VGEYoAp2tNN3xpfp12l/2me1tUBfkoxHriMnVNjtcc8Q0UTI6gOsxl7GE8iCsYzQ
1YHeS4FfTA6+AVQJ+G+j47376/LuziC3OW4VncSg5kb4V0oo0dtWVu1peGcFjkC8J8zhAJJxmgMJ
jqpU/HXY1zmdthkR+LGDkYgcwNg/2r1DYqYRga7BEZ5YJTH/7AuFGJuNf+EybbQovK+rj23KDbWi
99lR/ccArgvpiGttLsgkSJMnXPl2cDQxUYKKZNWr0S3OCOa0rueVNwRuAjDdSjEqkyHjtOzkRb/2
jznvKA2u/tfT+oEOeqXxJHtDYy/K4FaGIlS/ipf6NeQERi9RX2gB7PDMMOahk77LamdmYkCRdoj3
VpOyAXnVs3TdYzRmsE1YvujZi6UJNsWiRSUAUUn2ttCpwQW2sQODudHRA/LfYrSiBf4sZ+o4NlRM
DVzihijdDPRd16vBSaw2dqEUuh+5Fxe39OLF5yeUHxavRJVSBteDf5WP8QcZQm385d8XjZ2Jp/CB
6lkCM1da+NGNhOYvWX73fGh91MQKTwn+gWbm8Yh904qiXeHSjqchXpnsSduXpSdFBi9tRUKO1MML
Qv07tmgiYvMWfAJGhA6o6Z7owHqPUp+n3bGSt6AF8Lq7AT+ddBfUCUR78zeOwD3nvNfpZ21H+rzl
MBGFtntq1KJ4y2k5PQme/7ZFLy1xhHAVCZQycqSIpbh9v8gjJKsVCz0RygI4pBJ6x/KRfa6t6vJk
ZH8dfFPr8Ewnl/hTmByimqIcMmkB0lU1Ph8dGirJcPs6ESG7emoI9mq/JbBg4A4GQpUkwj56u2Jp
rcpB0LOAUCRv+ML3O2tpjAGx/vMZnvGH7pP9H4m61mQttOjIAq0SNfm5zIXN2m2dvuWRGfLH0DDW
/f16juBvZxkVP1a8oCLtZCv9uLP0VkKNTZJ1hVZLF7/ighEnTWZ/N8CDiwf9KMmdKEU9Bwvfy4mi
hQyNwkj4FUKDbQpl1bz9JppOVwyUq9gOLc+fvJ+gfh849GvZAl1o79OOYlUECqrJ9f5LWcgjO7q8
8wi5s9tJe9YN/2y2giWG/pYi4+8QEN9d7gvyvLJZ9sWs19EbN4yGwGZPbSx2bwNedqu5ANk/xvu4
oem9vqXALidGghHXXlCDF+PsXZMqkWYEg8KRGjvVXwLg7uVL4ceo5SOnhvpRnPyMSbDwhkVnSmKb
slaBcp2kcKlfyu118BbHGvk878xFFok3qGGUjxz8Jsr/6LvJcYcKBNupW8/C/vzZugaMjlK5D7y9
4vnZsrtEBEu/aQIeZDdu8P8rFOUE0ymegJO89QqMULEg0bbkbkppFL79M1Icxj+s9Lin/9dHwXSq
BDqBwIGlXV+WCL9VRm26FBEVR0RWtTKFIsNz0+u2L4ySGYFEbMXh7O0HYG8suOINs+yWEe7WJtZn
/9L66d4VISr73AjOfL/5KyEDhLliwg8mXAS/+z0Hzmr6SCwW65Bas/5IPcpal9+6ImlOEbvlApP/
tulMkkX0OFKrSiENGpdr7z/YCZhqrjXN0emvqmXsyc9zQ9bJCvgg2R6SNcbKy4B8CRoUINxLU9uI
l97bKa8Dcm39esIH6+gwhLmjcgrpgQ4ZVSBEl/3wjUYJcfW034w7bKBijcUe0woAvXLxKfvvn8kd
A+s4xph7BQTY7KyERn3uNxRcAjZOGf+vnmLXc2nG77j6wVPiiM7FAKC9TU5oTB5Sfw+l+WlNCRmy
j6YQlx9CpjVBbN4AWegm1yh+P+HOG3I6nqPE7vTk26+yMYZmKyOh+mnCr2YcaN3L8pi/3NsrISl2
GGXM19/B9EetNCrhZkj0I4qlnv7pgwXHMLVUzfGU2SB+FACz0PsBPVDe0u54rE9M8KLcSyJmaC3T
SIjxJOnKhHG80twlD8FCi9X5fpF3QsjHpULznJjgkaXjVdMkNrVLHwwn0+xVpD3x+baaSDdLqOR1
ttQLxCMaetz9sGJ7oz75epzANAyx9M9hpC59dfbhVPdGUO1fuNo/Ff3I8RreUQnIgVGj928On/1G
HAaC7Uq8J+CjUAARQ2RpJLGL2aEjszXjD19U2PQkUqYvnkhu/EHxWcqCP4O7zkwAo+AxLYV1QS2o
KkgqRNrh6RVkG9pavTxJ/8/As+gjVrMCfUAgtJ9jnqSuVe3dZ49fqp/aG/ZCS7Z6VB27El9q7Sy4
xd1rDGiJGwmMzkZM/hugyytltOPiUe6A+fe6GEjF7zHig6+OJxHCyQBGvyu+ecyu6/dYOxYtuuU/
mPUrg2+43wdVznJZa/dSXSs9PyShyTF/3QZiWVPPTBI1qp6vDzSzrraPthoDj5fDcJkyq9iEYDGu
l4LpzYDC0yCjX4ha+iB/ObnySbgiti3eevKnBHZo2UWWPdabH9L3I6rB6/Mf99hP3SGt2S+c4it8
sBx+5MJclRx2fg9MfMbU56RKPDOkiXC3uyMisJLZE8O3EM7EolXGmlNkr7ONYwtxu8rqIBPvNMOi
JEuUZOtregLhTL+l/cJkacpCLND2vfaIMnEZQ8Jul2hp18xuynAdN6gBBDHKufmvZ6KhB+Tv2QOt
fpNKoqUfHVe/mOF7ukzQwT81mGBNhxdh3NR+QfU54iprBsz/ClZP01wUiu4Oqd+JS6pyYHDGeIsC
BterUV2jpPNW6k7n+Rhr2A64hgf/EGKmhJkPHXhx7ehdJwr9G6g05xhiHihEnYzpiGIY1MwQKM/h
FnLdmYEovtQ45FmtPhj+0uoaIKoAmNLCKmKRRHsVk///e9gHmqXZ/nj6QTJ9n8zOh+C13Xk7eGOe
ToTfrEQJMktB/8b04XOasZK7i95oYBBLzh7WK8v2wZd9lvMFY51//2v6Qt99WgTjfLHQ4ik4ck8a
BiLV0CUhPwvHcCxdLB09Q858JcLFtM+6iKu0777kTHt5NiQvNoJOIdQGcTbnHhsZ1MwtmHkyxdwS
ZQlHpN1Adl+UgKesw+IQ0CeOnitL5MsMZrTusRKIkBahWxPOLuU6FXdLsSG4OtvNNjM4DuJ26taB
7lYixE7gpPXK+LTsB/4H4oRHAvry0GPXZ4RsEl7z/0quEUudG+1PQG31jTv/W43Egpvw36Is3/Jn
yKCd9aeq7JdQJFdztOR1J8R3LAo2qWzxLO9l+O4VWhu5Qx/WpGkzlivYDq7i8Mn3JDnD4qeWjV1v
a14OEAcclNxSqy/vX4vMb9LPDmKGNdsHYlQe+qixU6nxqov7ld9xwol25HfFT9W/Jc6Rue7YV09g
hUBZHgtBCZApK/QA32mPuvieMn1/BL/phxw2sQt9YCmJW1ZMd7Cb53UPeBtcDh9FVfBuy/Egy0RK
x6oefTYVITvjDz85Ia+yrX+T2AKnAwWKVwTTFnFWY31LIG4s5CAeIz8o3MMfmrQPNv9kheJqnmhU
AhoSmqonfmY/goRLoywe3QmtOH7SNYiMr4qFnX5iOJROY1yDGt3Bxv+dnfYs3jqY+de7LQxCy4ci
Z5OAsWcdHI2d+qj3CR+zPn8ZsMy0qL2B9KXXXLpkodYuBx08YMoDhkSWtFq0YBfmM8VEHRq8F5QM
J3/3lS/D74Js3HCMmJMXTNkR3lY+SjHtqUYnZXd9iPZDM+RJLjJT1BgjKDMABJU27+EkKbfhompE
aRTgvqRWRho3iIO8MgoQ0qx7XQbxVh50/6oA2wtVpEgv7ixrQvP1f7NUIWd8D+rGU1ggf+ITm0ti
TZerXL4imhLRXid9EzmdoOdTp3YAaJBU/I14BFNA4vqWB79bItQjrb3OuYE9o5C94g3UsmOTygVL
XIvhY4Lcvnu4mOJUd8PfvwPEgNpVda6SxrL/D8p084K9hfc+/G4bXdcfG9jHnMBEoCpW/JXSCabu
HGCa1Rhc4YSZi1wylufq0LFH2W01ynIUIesxKDQ6/KwVy9ih45BN86Z9YbaFssrafqOln4yiWUrS
OSP6zgQdQwvLrbQqMUDwBLbmyj7A5kMsDnvFJu0Mj6Ae61W8DSYJhEw7hvHxo6zOyX7/mE7g3zwO
MeN2/XjY4CaMhsgC2qJ+/ET15to/xU5dcAo7n+mrh/dM2GTAFJT2a4ZpMfXZTDZJ1+5PuKfXfgk2
aXYN2Ggj9xKcwwA98Lg4Pz1funJL3qUzp0K8rWFQyvWVntofXJZm19g6R/qHOgxw5bzYkLh4YHXm
x5jAE7e0VCVRj/IYxAJkv4vVqJffCNCJt1BAjoq3OkOM3OE/ph6s/ShHjJerK2tMDq94wKCS/E1h
5bRPvpL9XA8tAlX864e0IbBsk/TE/yEHBoewnEeNIBKqKykXQNJw+AaNw+xQAjpoH2LbcY4G4NGq
zg5OP1gVB+zhfVi2Ozm/khVHCu6PnzfRzNzmxeuYQ0jHW3tI/5+MhALJIqv/e1avwAtOHb4LcPhj
11oNHdETePsVaEzlcJEUDukrhTC6qybdP36gPPlAmDmbexIPUmCg8QjOZ5pix9r+zrAvVAFTX8l2
DW124L5xAsoV3lWp1MrXzmkQ+5LVoe14LUybx0IOWcL38Zl+BSCVtNnzgkfEDKcUk7SRNvlx9L5B
mRLRpqfs+hkZRjx1W+keOTxrQD7ERDsWQwNbZTCnhdgnBLrTDIvpgfudad2PxX5mDmQv6MYiZG19
GAD0HX0Gv9rNbSFrdGNzNsLzVgh/ZF9zQIW0HR+FhtN9Pc3uS0YoscL8Lz4/++XZlDpAn0y7qUTj
elPB4dUeiCJepqCGlKu2b4KGozx4g9MLCt4d2p1qb8MnMUCb2XmLFgsuG4L848trvnKUxYJOWki3
YGEA+lstSxluqT3/daZgmr0z8B91Sz2fnk/Wk1BApBVTmkkpYheaVJhf3WeHy5I4rQPaK3S8KqTz
5s7ly8KrQlNJ/2aPq6v3l003zOl2hj2GSxeVQz1oHJiTUqN6FUR0hQRjURp/5XbBkcYCV1JTG3IV
15FN4+OZYUw4144QTKI1na+ampJKvp2LIfAErX6uiKcDtXBmpD528GKRc1NroyUfQvFI6Ot3oOat
q47E0hT4IpGUoZ6cvudeQoQG5GHEyoPDMoL8315ChJto/xCo+l5pPwSxvG/lRO43iRPPBlPGyCDP
TLvk9DaefYffieDxYGuh6EcZqJyxt3KRv/ZlyAfW25jhhxqZScnqPKApnf5i+815F5xsCqnwj/mi
7BAI85B0QLAHN6P4GmUHL94CWu6nv3Ky7xzOoT9tt5puBfZtEa3jqhrWcusQArPEbunpFP8yJ9pl
b9Ws6Fu/doEOX7bR63Yh5fgncCL6pEw3LtG8UK+tvReF3VylNUWlrGjqJB/UrRt6OOdtUctevu9c
WrxcELMXKFOhX3XyVYzBGkT1xqAGseuW/68+FW/kwSHol1o8z0isI1nVsY0Z4wrYugnVdn4f8Ssi
jy180tcTn1sptr8WaBmKvm9CzgPlBtaX1as6dC2jdd0dyq6xxHKXAfQhjeFtoBNaMWp7vdUIR2km
yxzL21b5rapZUcQuXY4Spvg210oVUp1J41yZAv632LYzYlgPjBVaapDm2yUK0CgniwVZoT0TOkVp
6xxDNcWuPTesTXimgBljxt+sQn/yKCZq8cU3O5MilyrNhqf+fZVmZiVweVvQk+WKnul1wUNnHKmE
Me3GQ0rybRpIOUeNM8rkQCzhzIKt7yL8mnNlITmPc8oe3zJDDlMEeuCkNmhb7xxfEnhvUnba1T4i
XBAA6tVeGH/Usb1WavW8o+hfRqoUwwX1qiVynfc0dKYCP2ED4urX98iE4UQ3cgW0IbPyzvLyWqhE
1P8gmitfhxqlb5zUdDE5j5mIM1OdZeMRiQvTt/u8Epp2XKqxQWrtuyJBR3AaliBylwfGgnv8fdHf
7pOix58mmEkvV56KHeHsLE3osUeSsJSYAev/pr+RG3swJhufxMg610YmSTYGBX0NQ3Qp0CIU6YM1
fKq26QOFT7VgXghYDpiRQDl33ZWr5MWWaH61K/whCQiQfTKvuulFR2V7ID0ZrGvD/Nrf842qxU8d
hL/1U5/gQ156MLYeCtO/EzQx1WnENiJkLvbd+w0Feg5x213uQO7V5vvy3FH8xpHQCtg1MYMcv8Bb
+eMdp0sP3A1RDUJa4EqotzH+5P+Jsddl0ZaXI7Q4W2Ya62WQzGI9zNVABVsCxSH70vh6YQ6ffWwJ
+nJ513wafcNfND7Ihd2cTqFkJC44adizlb08JjoVcLV60sFkiTJpg9qxI9OEUGijlraL0m+PibbZ
A0Wdf/81cUGXvDNYB53JxM+p85hJ9c0KQCXj7vfiLPCp7np8Ksnd27YJlB4+sW0QSb2LTXHree7C
93G/vnHcyAX3ag8VmH9eTbcBmpE0OIy2J4oV7kPq7yomllJ7qzLe3LD5zCSPeT125eCrdrhjOnz3
cHhw0RSfa+axdFXf5aIJqYjmzyNILYYN+VFfSJz/kFmfFXY3BY4CmPl/YuUAKQm6fMERw6uR4sxK
tnRp235vVQrDVUIJjWYH4mcgSz9XAf8nqR2RyV2CXP8uJ3VXMicu7GU5RFVaNWoGpQzOSnPw3vV8
4DmW/Sg7s29M7qo36U+nOK0QG61Pa6xpGoBYCybEW8CAcfjlMO61gOSmOyfZC/wtSirLvogcvD2D
3N0+2O6x8BLB9oXaSrB26KpDyFyW9lMKtGfjqyCgoIGePV+bvgfqSQEI6ONp76o1ZRYHKr/nZxOs
rh3QSTdIbgJg3uYG3VdIJTaFYmitfq6K71+5OxN8TY/l7JPcKDr/qazVr5Gpvs6gpotaoowAiZSA
n7tQYnBgy67beNwFDRK47p0MffBknuISFqj+R0hf7poDg/L2+v/MpCEZvLKXMCooUgseM5ns7+sQ
wB+H+VtVnNcy9r77rTl2E2KOt8IeYIM+izSTlB0tVdgqP8MUhX20RPjslnJCKrdqu9UiZtVjya7m
eyS5a49xfol+plE3k7oHbAw+jz1A/ROC+O/qzTTyFR0mhNEYz+M9QExu6H5X0+GT5VWEDlwGuvJA
pZB8mlbpHLPGl2MmFXpE14Sh8G4AaT4WY0snwQrlWpEppgsMicZP9u17MQDHTKyeH2IPiQgctpDp
vybrXulsYOGA//1dxR/auVLdLuPI/yXhq6W04J3caUSt3MEEI0MS0iKWC08QOHDp8VN7JJiaP0tL
1M134tx7D8P4WFWpbzwj0mBG7ppDOLKv3uF7hwmwrj6vggX3UOg/00cgC8XJv1Vb1abGaHTxn2em
6YaLRYRzWsB5kKZT3QTJ4rXEn8F8qGvI0g0x1Op1vye8MnXFMJ2L5yVh3ZZXNXH9Xph7GRG76KSg
ZAWO6RIgyWYWc0aUEaUiHgFTdCdmry99o9rbycjvj5ARNKjwXKvYQraZGSeIhxd5T60Iyvb6QK+o
u3iNoWbRNQWAsQkI97BB2rlu6NJBiGFJ4iwbIOOTR0Y4FFSqvus4DAQQ6pBzh1FFf1VVkeV31x9g
CpP9qQvF68oFegyYpxMy8Hw+9VPplv0PiDYQTAya6onsGpZ9CRe+OyjO9VsyYXXC+VOb23SJ/JXP
g85iu2hMDXqF9ELRfWDvLU6El8Bvvy71wLnLTcnLwRLAo1R2vZQfp53NsfPzkYK/r1bvDX9A9itI
X0SqgwN5+fEMmekVv2FElx4v9RMM9f12dmpp8lndOxh/+MziXHUAZIwnEdyrkL6v2QrGxeZZ9Ej7
JBNbXLN1wiktE/COyyi0jlXVRWFmNvqo21IAaAra1//j7AK5DA3RCDPb36QXyTEg+JQ0jYY2LlPa
6Nhx61JouGLaML03rHh+jHO8uUK+Rv5UtZbfMHD5lBBsgNBNPKbxZZry9zsfziOSd44Kg1bNUsnX
WEm3eh5B1EGnvUN6K50R44CZzONp91udWHWktBbCF+U9QomC4xWoG30yfWBNqBQD2P+QHFwdVcr5
CN0XqEwUyHzFjy8UeGABxlI5SlSnlY8O+S1c/hfs3An6JCv9SinFzaee8r7h2usAtfNKBMFPWVqL
EDNPMvxORwHWWXTa6ceXgPv7JrNyIJ8tA+LgB9LY6xEhvPKXzqq1O3dqm8UIFuV8utdGkq7TLVLf
fEUbahINo8uwxlaZx87K92XG2iWNi6LD/n7TgHzjrlMRJM6jV7fmyGL8JsxLyVEbE+MlnJnxOwTf
NkG8b+sGH3/rqewCZ4PF3PAAYycGiDFtslh3einb9lPrFXHJ33AStHBe5JIMbs3gCtNF9QbjkuFa
URUl2Bsg2HGXQtjBoVLyaXTDz8RfWuJtBgl5U7L5toR39Ds6Q4GGymsgvHyggEZYMumeLFsxR9VX
CH34AiRj0cBGJgPne+yuiflGEYoAJ5tFbAFOgwmIDUrEfGgk2JZq7G7tNIFMUJMJdHMfDThnjpfo
ixubhNmphxuntZeuuU3r9yE+oBMh4lNZte0bkZ98qyLPawEzQTztML37GIbhIG0ef5LQeDHBjb8i
N+G0rKiKlzItH5KKerSctVFiocbBprVngOzfKK1vdBtxiYnB4tH2F4K/Vtd7CAn9CrqbvI3Vt5MM
SBsLjIUOqQVAdzRt6AdZBb8kzIr6eeqFwagK8J5SuNJtaWtqt9cKltqm08UnFeOGE13+qFlJ8J/2
l2HVEC2lIo/vhkI7LqiZ2xyka5kfZJB+9lcW3rRsEqWUYZQG4Gk62NNLNEm7FExrWcAWeGXJ1eiW
SQ+zS8T63DLPRHUxsaT2SggSdWApVUHnCDVR75juWPFBzbDKY0Yuo91L8T4UgsEOTKiOZ7mqc9v8
kyelx9TXK8oaZq67L9tjBrk6BXjXDAc+Bmtz34pQ+Zj8QpPNHMxv05RFGagfm4bArmarxawfJvJ9
xjscS8X3Ii2buOTBYdr/ex3lOsFD+e70jBCq5ICndj56n2skdEOEumswLpXiDomKKOrD8d7uotCE
BNOGM9aZjiQ6VVOt26OLNHN3uniGbdW7XW55CAjGaii66ly9zROi0LYAtNA7xjPlL/JQIdlUkJEB
q+fevW1MfbpDlMuYA98+7m9fnHYkTM/ddwrc4tWJSQisIqFioUjkeW1cUK645IYlLaprRzMomDV9
5y+1s6ouAAkScqeJ+p+MIZXNSrv1TVv1tRQMyZuUWXULOG/2Yp5kRhu2Lta0kaNemmUwKvydh2Ls
LVGv0KfiQEfe70NgesJvE3ElAtzB8gVe33ajbbW15zMOCdYpHf2N//RHpGeSBAgO39jlc4ok60BD
aICZ6marIJuPN6QeyLGPxWFLWq38P5HKij12JjBDMLYjpKLwDyhqn9v/EW2shwT9eAo4o5yO+d5e
unG3HObSu+LdBI80xGUvd2S8XjSyt/3dduDyEQyBcXZ6cnc6UoeV2D9zXxmRwaoxTwACmzjtI1xY
96skD4B+RJlJXnDV4gaNd/19+C4qTFtYFvvJdSIOu5B3adgs/mpHqJg9PWy5px49O4NNdEmpTHw+
fCdFNDYf/BWYAp4XuFryFCMAKXZU9UIpr/lrcEqBNkDBfpctgwHprJbKNdYQAfHCmdgbLpKxIqB3
58lPt1ezGr8uM8XrYdkPGZnU/gwZrTu/A0UzQornsT2N+FBDvsOMy6qX3qQfa9Pr3fPyaRl2IHqu
l03t1NUdT0fyWxFCOxsXlK/iD8R2kocNc70emzTqVsrztbxdTl8vyVZtQJbUWZHEjvAimbSvzbUs
fqlj3qvSJKrzlNdL9bE6mRDUIiV4ajfAhgFf/pEJOsJLYLdSLRofb4XhUvmLKiH+IOu9Ngwjpi4B
o5RFcdxE0qv7QqnQSlGD6aYOmUjFWL1j/I4Rv8iH5ExIgtkYrbl17U5Y1G8UD+mLzcs+6QbEvMWJ
ES2PJzzVFolhDlDOa/U9LelJMPlvOdBIZitS9V8XKtJvUPbRgdsDe/2ZlcZTXhq1na103ZJN0+Zq
AzrTgRLfGUJeYTQcW0W98GCtXWCdAITxc3NdM+79sQDUwJG6hzKu+6Vo6fYauJp54wmn+rBmGwwg
AZglhba/DWcTiiytUcyj0mqy27erDjUDDwQySCT/OOg5ZQhdt5mmSQX8FyHnf+8HfTaADxnJw9UK
s0QnvdoEY47pyPjTISADnCC02VNQHRiN08BPZ6ehAE4JYCe24gnWCrV7XPO4F1dOHZrHojt/Ni3x
001XXzpIwVgyVrJm6YjzkSyjKic8MspcBENyiald5W5FlxGCRVSFxPyx/QA3413Nvuz+Xy4Nc6TJ
ASq0FshLhV0XtZjzZk832wjXcStXQ5jliGBLake6tBVscPmlVJx/Uwhw3k8uNzs67MHsAB7goh6k
v83v0eayBgPXsMQQ9DvXItAelZ73tfH+xXbEGCJO/9OaUXx5/VyM3F8alpp7jIrnaZSTb6tq9T0O
4bU+BE+xAgXyGjijdM0wG3wgdyhou8UCcQue1q7dI7GUmjkr+vD/Daz1M0h4NUtgWGyLRh1IAUEk
RyMuuXMM3bkGIbLuBoyc4FSBZJZ4UqDiwG8q8NSGQXbc0//PklGVdf7j2EWFrabtzAO8F93j1A1c
aFeXYxYbPqV2AF8EiWZ4TN3jDajnJT4RjyOKuRLfPiEVAPQQ+r7MrMWIK0FmPgruU+wzwwfzxSTq
SID8vL0WLrq1Gx5ZdMOIfnDksmnOIczLKkFi6Ih44sZHsdZa7rTZWkqSI+OwztlY0bmtcwPZSv9f
gtXYMgzgLuVuBRTgtzflY1zzK7ibAObVpgHLXed1hkJS82xMt3V54Dg6hfb3n+2lmTOYaec2rKQE
hMjQzQmCL0Cb5gvowTEdMvsPOnz6nIqWMnBRKRvwO4aO5qV8tR1tUXWiVHBkslqrUDari3X+oH3G
GV2XtznutPE8gFfN3VQGbiwEIOW+Jt9NXcpZ85kJ+5cIFCGnxRPGa8kZhvALyL3iFeJxIC70ZKS+
/gGya8oGtfgtuObbJaQS0LX9/UGUnhC2mNJimKKcivs8xEsiFxpzWsc9e9oedRxkOpSPtdpeR0Qa
jkhSjCjLf3sMJ5ARXxNvnzbbzZu7u5zHmFRv79jP59/Hi/LRI65373PpiXkQIfP6ea7GuSxWgj2m
dCLWDRfOck3ha/PxaVpLe6WzcD6lHxRglVQWAyZgp2kIcsoxMzQruLO+jKNdY05Ec9yne6UkSsYy
d+ET6RJYd0eSPBEL3Dnj6zGqhY+N+0QfJabjQM2AyEEFd4JWlh/RDphP15SrHDyXPE04K7AYBtNW
adr61Daf9b92C0wUA88htxpZPWEC2/MiOBo04gMAIjiRiU1qa9bKFnOFm9zG0RJLSvl61Pw2/Klj
/IQjMj5iMj5BSbw09wumLCCWG3yp82LvFmpcg+ZZBy3F/RnX4W1t7w6BXxz0I8vUZ5i5NHw0rsGl
sWMSewGiyjy4+SwMbaoNgyP8Chz0EZWfuDK5RmDKzPs4gddmaVSwGRTmwC3YvUxoFcTkjzSgl8e8
sJ7AXL9dN7uuD118xjvoF9HI9mEFUNSzZItbcm6a31d85cOZHlS4r627p1njrgysJf6tarCQdbvf
jSX6HOz3y//l3A/snAsJO1Fcw4bi29RjDsKOQH2xpVBZ/9Mt4VDJo0M60UGdg39B9moHyWFHTfcd
lvW4WfsXgQnY/Ix4vWY+dx2RzcFuJA/fUtmdQOgNIcYZnjxTcZf3OtUQf+mdsg8dPM7EdVZn4wGq
fdLwH33sWdpqWK3jFbfRkNG0BOjZZqVczjMUc1LEtH5XJPAy2qiehO+sqXp1HM1R68at5idfNd91
T/Jk1Xw88w9vNbTOTbDGmzCfemCwMYHKevwvouHhp8qShIUyLbNJl4W11kjI9pfSw/T+hJ6BNjBv
I4XJNQHGPtGoB0cMdXYIGtcl6A1oUa8RDgaiJPgMs+EQ8o0R2csSBd17Tx/PAs3Nzmgd7xQDjCR0
ENvGca54b0rHFwFNyEbqmC3rIqf3MdvHS3vvT2qaJhxDJHL9dJtUg9NAhFI9toDVEdvT0H+GY1U9
LpUskwZuqO+dDfKn14lCIEGtPrCPcoKrWPBe2eAci49XToQw0ZwkROIHMX4iQLAmBuNbag5uWOCn
4IIdS1Tkvzki1Ykj0ontGG1x0st00vUtbeDcgDKULBWgFGkajIA2klBokZCwa9H0wUTnnDEXZUKu
PyI6ArEeyd1ykom4JOEzT0QECDbTVjT+TVcu4QbgzncLHx8HvG4UmZNU38avUqo3SJ1RA/XOxhFI
+tdvn5LmD3jb5wf085bfFIE55V12kSJbhy3jTaE/MWVG/H2Z99TM5mCE+Pgrj0hnQnbIObHE1inJ
H47FSsbHyeGnGJTDRqFC5bG/L4GfXvMwLa12mMm+Bpx6DKHjwDGXxGXGWxVArnhjVX6AiI8cWuis
OBROjCIeaUqdGW9bOkhwftdaybgampaRcSsDnNBoe7cWKy+Bx9uac4s0wHFL7WR6K73FQXXvwXxK
Iv9VC5BdVp9CSM5kENuJm8PHRNjQvCqx4QmVS9ICweFouLJikWJsURvcJex5rwq2V0NpRQJJBJdl
BSc665u3rRYbbRTy+0DWCcR10zASQxc2whj0P3Ertr4zJr+PVO5pNfvQejDcV63MOpL6UJqkSQuk
EqYSEVPibXcBpbiWPyIy+QU0wdqwRfeWuPZX3C+C8LUhJhYIhyhckzA4fuI5hqIKLhbOEmkzGEcQ
QPa4eFBNLDFRf08FpvGhP5SJ3x0ANHx5RlGiI1SAsOtaqFTTzu4rgw6ohev23s6uAShOlcyYeXmn
N1S090WAhDYV/zJ2Jt3sTsKWYWLkuNWVlPV+ZOBivNiqozh5ZD3bGT3Hld6qCJ8P1VgoNmrWkeVg
b/Wy6ou4ySVrLbQHwPWc2/YcEAcYXaPV+E8XV2A8ZATYrv6shRGNWGrNhJhDIf5YcRzBAMxMM+Sr
wxypgECOmWO8S1CSNDIX6+B/FzCOeaWyBF5je+8/OByBig/cGCP7uMjCnPQOd8Anx38x70grZGju
/alltLfxmg+/AL/CFaHPHEwWtlhmaMcZ40zr55eSoabDIwUJF0SMml3qVTQ2BCvg7lJsgPetiJEE
32sEgIWCcYLMwTMK3YzsS55QJxxaQUzfrm4qFkTriCqQoWuRcIwRRCXnU/nVQB2hJ4oPpqdoke8K
+jL4bHVwKeFeT8kpFQnrRCI5e8+GTtSEHH2lvonSa1XjFrRbMmQzy5HTH64B8hYwKiDajw8C4K7k
jq1VzXlzX7QRNxea+GEY+hA7iDb7nfYnIbh1QJ/nwVTQ0JZ3lCdAVj0/s1mc2twO4n9bxI3HaWt7
dqyFY6S3aoTvIQSxxXRvuECH48XEmBNn4GIxiogUvyS22vhst3xnrAvM2PFQ33qq4KU7IgZUW7bH
wdRC++JHMW0rnVtT0b8mKJL6pjWR3Dk9r7cO1VGhRyPBTYuqF1SK02QhKUMaxSLOjX6OxlvpH34J
XrShFBqNnFHJYJUU4VY1ZcveWwog82nGUM4CMK/p3FiTOlPtcVQvqXNWHaLB8NIonqA2SY7a6TfD
C1AxRf8xr2aTlZAL3T+15DAkh+7f455nLuySjFgGCmHgJfbTWyoKhwoenWquoGa+VFIZvCJOJ1BL
u5eCqYuhg61AvcBWsv2jJ2b7t797/GZrBcTeXFKu0raL4uPnJ437d8PWLBbIgHfdAzFN7ktvEIKh
CA/LNy7TlVzNzSSqpaLZkjOXGWZvT+zaqosFBKu4dgQWH3yfI/EjckF+JqjAFMyhfLj5gTJRd5CL
4TWf78iYBvMoCX3M3FqebYFtQqx7JUPuXqc/LU83z2J4grjXznCgbi/BubMwB6wmfOCHi10kr5I0
ccthV0Q41dGBEZas9JTF9yiDjdSmpXDarGRT1A1Yjxz5I3JEDDYPAhz9HwnnvAuMhrNMQ9gwdLjB
K53SPv2oa4Se5X67T7TWJBG+f2uWALUChwC3tX8b5QjJ1QVY8cpOQ1+B+GhD7uzDvjzWieAQIHA4
FgETZLw8FnsQhIHue8H4MPRa4pKJLBHHwE2LEgt7/BdQTLMvUSNrRQP+HEF0m+WUtKMf2OCXy5x+
LZgs75n1hgV7GL517rjA7mfaBkiFtgc56lNhCsxmb6lPU2bHHyX7dC3szSaogkRiXAhoE5wz3HBz
4FN67/EFRTqPdyTGoU0Z3nvePywUTEEX4Sz6CnXLAWyKRXYPg3fBOMGEQm1HVX66wx7gAxJzpGiD
xZgsTdcc6wOrOOdPsN60D2nMN37rHdDfHPHonZPzYQf5BdgNfpgZo3lZZ7fgsxmCHmNfwWBtulkY
2BkVGKqgYSeEFZTTIYmpFypTmQN8ijdO7HghSHSIU4aRMlr9TcqyRxZo/vAR89jC8S7wU+8W/1l0
6NRq15Yw2YjTEb/iTicuY6lA5a1Yni/Q0DkSVT7hdm9szREW8bFjmFuiYgWMceQwaB9PIJWSDP2S
Ne0wW65ZkwjqFfMR4h3Mb/UsGEzCZxrUvY9s4jL4ZheoFxQMo2InSmkTUvjkIoqaGy9RKMVbaIJY
zxJ/iXjHluqJlQPh6IfQySEKd1xFJubawjBM6KBwGdWTjpqJk9UunRfJeWXkv+BEUVV0Vrr7qeEP
AkTJszuwIENMtrdCIBt91D88jSA5d447XVGLllUK10hwtwmeNKbreg5JOGo5fxU2jKQsKhrnSPgA
iRgJy6DrAgAdIXMadmvXvXh56fQC3iDKrTnK38OxQau6R1RwA4oF+iuN0olt3gmpX+d4brEKGUQi
0I0BS9k/6qn9LFhJ75uCt+kosEu5HbXyRZhfWhxyN7l7TeRP76zv5Wc251G3dgtPoz5bb9AnoHCw
qc0TUihrJD5kEdqd238F2vKcFyrz4XzXjOda+ZvPwASbI7m1spdSLipXDGzHNXgTy0L6P808ZPVu
RhjrY1oYuXjX+yWWbDM/cbKj6wXbO+cfM/69HiMZPYXXYbjYqJou7w0vYyCaXdESoP+9RBPBznyI
dCAUeIn3ngsslMbTIwwid1zPwAyO1piA9+WsIPlpgFNy0/qgUkl4p83EVsUM90lIfJxhxTun68QD
jxJWFuy7imVgfwP8UEcmYfdVOXVKpCHq1MWSTGpZFECji2HbYpSGI27ZpdCXsffpgGyBhU2UwLrW
4WNH0I6LfC7X/HHAvX3xm0ZAnaPILZG0fLRdJaUw89SpWOpElYd4tMzwDjKbiuTzN2T2QrJT77Fj
UpiSa5RcCc7R7XbwLA2BVoMFvFoHKkNO4Dq6l/hoIZXy8tQmlwPzbc/daK6IKGPAW4Q6/3etLtWj
jYoK0FhSDBfMf1IpTStXZ6d/pw1UFS7Teqn59M4tWyitKGerZ8VQMKYEjgHoXjXeFccRZD+rrLBq
RCg71uSW6UGi09Ul/srFqqHls7Lp/jG4Q7yFvg/SoM6BW6nOJxwhnK7EESUa+cZTpcDVs2yTHsk7
l9piSXmtI4GLgGCNbhK+Mi3OrXbSIIPvB3hR83tt9+YpxY3S8ztQq64E4/YDCTCuvhMROF/4E11p
Q7LlrvoIbbfGC3Nx0u6KSXCwz0Q5d7xDBNWYOxp1jwWaixkQu22W0mcd9iawdO+MWeMnM2AQYwP5
pl3gxO/k6AHcFxHi65c+7bYVO2IYSpxJXq0PWuRyRaApPyg+lTqCFHwQxIZVX5Ovl8d0DCbBQCO6
Cmy3xRM+8n8YWB1KaHVdDxXyt9AhJ0xfjXCeK7+WjiynLfbC3izYrLxny0KofVQVejYwfyxRkHKr
je062A8x2+Ir068mGQZexQhpAnK9W/D8XNknT4O0q3hLjbRRDSW7gopFaSBvvQ3e1jXv389qKNBn
jlJphU5Fsinlfs5BpUss8gQmkmOq03P/u9IMKCqhrTnpovQCAJ+E5m5Ph4YSFmfspO/CvCu+P5Ty
rsl/wH7l/1qkxkQe7TMn97zBIfJ52PImsH8ElFJy7BgttjjE1vUa7Y55BYLaFAVgMBpbDMTgwN1O
7LhdMJdxk0WXZZ+ak7tCQnTHYspavXGEJQ9al4d9Q8ggO6UoQCwU8SSIEp+6P9/sZA2Ieg9Qh2Jz
d2PFwwEtZ0WpzsA4wFmnMlpxujvlzId6zn02DNjeqyZerJUUThtD31nr+zT987q97cPddcnMzDss
bzMhNxLMiQmKWBFQPKgAj8JLYRhHq/poICtpSQTV++Oc8eRBIXrgWP3t64cUiSmdOdHnJs2TMQP8
8vUdE3pc4aL4n1dSYBvCj/Qb842IO0cFM7j4JmGVR5Pft8QGeqNaU4iEt+a8MorhWYUvFxNJcPDk
KTTZ9dJO958k5JFdkj49hiAXwdxMIYerJix9575ylz29unlfPFtnD9orZuvif/q/+NNthDABoIgX
RXObgKePdpatsWbunHRSVhPcFd24s+Rd7GMkV0sROniXwdH/sCuWVQDMOMfeJwSZOcXkeLvEfdzT
neR1cKE9mAeaKQAzAJDVu2wkxhE/MchnCd2PCALgwwjrU7u2UVgTiLIgYjEmODzVykqQTwsGYx6t
nIwoiXxNLjGWUEVgk/KYHEsqxFiy34sz6BycwCBegr7lMJa5kF1xRXCt/+4qWnNkP6GS8582MNhV
rjYul5dKKCLhvA5cfH0Eve093Zy9SP3yVgHe8gkwxBzywwnBCpCxG5nYXf0mp74bbTVXo4YTq0Ct
6SBo9xLUJpmjw2Ct6r9m+ZqIxB3W9kl5App2fWZWny7MZVSxS2EN3oPS6WQiqSPZm6wuhCAY9E9S
rx0uj/uXLEV3XkZZWAD1qtKyMnYOBfmaJ2ImZYkn7qP3QXreuF5vTws1rcpSw4cI4SjtULCiWKHI
xW947byH8syWRCFxpyMZhswLI2lnuI0LC9bQSYmWqPsbautaYZSPT6iTWmhgN+tFasnGngDikRZg
s/oWcj84ZUj1yrHMliPCePkh9Io7oMHYHgnX0vkFTiTOIdrVTDlACgcEYZGE9ospA5dCpJHdqMgU
lIlMQjGfym3qTGfVxGX4gDcYkDoucqGUdETIx+LKPzOZPk0lgCNDBcDxLqg/D2ZU4UnoWOVTdIV+
Gcved/KJY9/INgNKz7LT3m0QMkgIv6CoCg0yMY5IC6tJqMydkL6BuJ8r7dRk+HQsBDokRc5+kwme
utSuMrKvncJzCde8+2A+PSOEqQrsoa4kIT+YDjG2R5Blu1FUEcA1VWrtkK10o2AV5GYJjX80Vk4C
WF6/7LHFMU3cN/0fkNfqEizq/iLdxaIv8YKy0UfWnCrgg9KfVcfTTyH7qVgsyHqFk5rpmy0CSAhX
Dj73eP2uKv/M1FK1U1R8jsD7Kgbvz9VlU6ZUrYIkvi4i8tQxyFD0fyLp1fb5Yrp/+GmNAno0aOtH
Zo5V45631qCCp76alynM9PVLqCOih+UlfRt/wGJdd7gWI8PVi8rlB8z/CD1i2fkJm3w6gDaQuQoK
ZPivF+dPsHDwbau5OX/TIwxwFZfOi24YhSS4w9kM7b/pUUEld+Jgjm+pcqYy+Vvwl+Pd/zLOrjm0
oE8rbVw6/M5R1kij+zxDyP8Z10n9u8Ds8ChcEsoyLwPOm/k3u6U+9krzHgyNvb647jrm7bFJmkMn
/pTVtwQcDEa5n6wRVqb1mT91FLQcYD4a2PFSs/mNqd7nVHyZoN0j9//wYQsSaFOFGyx+qXPMzI7x
0SfBa4OcWJGWSKKH5ffnkluG8+4ZKNujIGacdrn+gQHlCNyoaKiOPN2Z+y2C7uRTRAWByqCaVAsf
9TfBx5c6HccAj3tldZHX2PVmixiRA+6TR2OuViMvnClM105icp0OP4yZpw4GwFft4vchKkQCGq9M
4LkEdoyhb0uRF/VQ1B3yxBcKWzHjDGMr5XMbVmVjd4DivhtncpYA7vQPGPnEeIAdLXAEZBbqVNWB
O8XEbTJc0JWEFfJgrW/8UbKGeb8NQdYNCTK86FTghePxrAHHLJJXIA5ts37nINmn7CPfJioYfVZ4
utCiZXJyG9BPSsNkD+UZpYIn2gd0/q8hG1RmC9kCfq6tn7DffVfwW7tq2Wzldn6ezRsSBAH5j7zg
ZuHrHsyvrP4R0kNiQl0lmHdgj7COgp7bTMCj6pLvljx3n+oot7s3Pv5bWiOzpZmK1OO7TDVvp586
V+FBwFeHQ+VV4CKlGp/zP+NhtdTqOtRYqy7HmO/9gIvZB4IupRo0Z2B5JXAz6Nm5jxodYNHOsgXs
g/0hPaRreKbaYZNwrZ7Sr0XMYgCgpQIuBFlF90YcxqtrvUrDj4zMcTVj3OZ89kQQ3M8MoX71Cfwo
ythbLI23rYj/bQ6jbONWOkJULWr4hY5ZuOr/Y0Vu21LpqnWQIjfeXbrMK/978C1vxM1wWZx9tF8I
FmAeDrIbsv8bU2UzclPBlo6gALADbufPz5jCqpZoruSswlm3qth8hqHVCqm+9pociVRrnThGJuhN
C5Sgh9K3dvVx6Irc/lyCNRUlg/+fhxVq71RG9tQ7eoTc6PVWo1uSe/rkzsDggV7mNE5/IcvYnvpc
M5b4HR6WRtn+us9cr1iE1LQJzezFS+rmbriFt2ke5NWp8ZUENpix9/GgVg+kvsSGYp4hJe44D6ws
cZX3IACiFvpjNIOiBlfrI/6slPSMsy1rBadY5vdsGpjAkFtJ1u4hiE0RUPcU9L+6LHVqIsJHzxPv
AhWPYxSeyGLWR5wKNpcWSlwJxxoslXOg40Xz40zjzXcn7cwEeJxR/VAHdq7qFwkjWZXs9Oc6365u
OGFS+xJ9+akGFtI+tc/OhxGqmWfMZguMPuk0sdan0S1u+uRxN7TlfnL5PXwVv1e6a1v7mHVmfJrM
HNwCg1ztCs+4vFmToj5J4iijhpdCEd/p7/BPQjchTN0Mt3VjfHa+UkwCNf8BEyQ+CtB7oHEVyVOy
9rjK6txmryfVlEw/7BLGj9wdTrcy59K1I3nsELAlNyjlh8k68Yk4xXc3R1ObKc3JWRyqnteOrBlZ
weuuB7ByxedyFiUZuS3Kk3CtlTXWZtrMDSiJLw8JtXAUsfDsRUus0P7jbc8y1co/+FHoJei/Q+bH
5EG1uvgmSKk2l2cqdofmDF/Jxx/BGGjcYIuKVjUGo6Y31vH6tvTGL+Fh7iQClxmGzbZetSW0oRUR
3+vuVGQPiUSFQGF+dvKTehmaVVL6kFksILqJFOI/UvNPTc9nEVzR41cRe/KYs/sfnIKHr7xbVrsQ
soJQS50dlJfQLSSJ+X0fjqBrYKCUSeNiJkBs+4f15lmSjZShirOQhOlqoxBLGGqY9WGbT2Ts/RD7
xTlzq3zZOlUPTzyslXu+svQjUV00bKWYwwRvtOChqiWg0zXOkoCbT+DBFPKoKG5WqVm+IP9ncEOD
fMxUoYZ7qrurPruQdsddMRZAetgkoT+DYFbw8q8o53nAD3xDm1GLgDtXsMeZsX6iFI7G0BU6AuFv
wRtYlxKNQHumBLCM7/4SlVdSy/tUSiDN5XTa8uDW0pF7AATaJN0fxkTo/krcpFtSfMWx8g79/v61
zHAGSX+iLyb8ek1N/whNzZ22b2BPklduylbJEO731AXPNVlnZDrdMb864vIzEfdLKlb7UxbIUcUz
642uVN9rxTS5PaYzJAfUR6boxsBB4g1YYHKGEPaUioTW4dScEV0aDk6y2Bzy1mr4qUzwkRzYeifL
cYbOYYvYcNmJfyx4X3/A2K9jfAhtf5tqZnPIOYsJFots1TIMtedCEkTjwfMFxuTDkGdZg59AONVA
OfhW/FSuS12UZERH4FFbexaxqPx0hREG+NwDilJS+oTseVSCYe/WQq2WmUwqfa3FUv0YUUauVFJx
tXBETklh5u1B7z69RvR9ifL0m019mi+t8WtYaY1qsv6+gZ2pf5f4vTH3+tqPUJ9z0sSFA5YTtBCg
PV82BfzxvHemCjnguQT3X41X9j1ZqhB3qlbF1ICSAKOIlSLmwuznbR/DFHM1TBwbxWlbN6nriSu5
Um55O9zXf4Nc/+uw5PrPZzeexpRJ8xsvB8L52tTrxQeQ/wxRoTngRjuq1La2PRNfXxYGD1qawQ14
8pqzHgpkT622Vxf/E2qEOeblTTbwf010uGjd1zPqpmgGG6cvJtM7WXnUc8LJhZ3LHiG1WAz/Zats
FdkG3u3wekFZWB+FhzC0Z5btcyxWmuAb+uMT4wWXyujVPEl7LxVsSGvK7L8xvF6JQVuXCRI3XzQf
/uO1bvepA+n13aCZed+sWVedtlevGXBIckqfAFgbe+qEbguwO3JMytv9UwLySXV7+dMAuwsI3waW
fQcOK6BR+PCFAxfvf7D9kennFvuJPpBeUupM1UVgNL7hkBB2p3zlErrD5GII0BvLS2aqbrS/cJFi
w++ZDUOy/azD6NHLGJYLKf9iDBJvS3h7PWmQn4sywuKnVKXjI6Kjf+jpHGhVmh+udBm+zBGWz4CQ
uvCVxh4qR1r+5v3y7ggS1igGFnh2bNTV3t8QX26WURefT/GLgedSExlZ/kECjT0Yt1OVaexLhrAV
8MhjBFypa7IFv5yKBG9tfxk2SPqagCuMHuVcZ0ZhyifRsqIvuPPOEPmbaPKZAqr89gr3SuBfOn4j
sg4LQf9VS8qoUZEYL8A7jggj2TJg2esE8xWqqZ0Msb0FLwgsZ+AVEnIOYDWalZShQXRE4L5+NgR+
Gz/G+PMkTmV08Bl4d6BbXQhZOsxU+4Ens1Yj7/D1uxPybnE7aOTa/tSAn23xnzeS4B563x/FgbAb
4DBCodu9aAXq1D7VpKLJwZQ1QmyEocTBQITcXE7lhWuLZWGEWhU4JOkbhAas2H/lEQVkhwli3RcV
TEHPEVMvtUCZQyQlvQwN+BlPZa/EKxUeYsruri6Frmz+9FeTL0KYSQTRs5VlQi9DMgGECvU/dDNX
yp8QIGiM74vKn4jb3mVzbzo1KXUwXLs6tuGgEtTzuf8HcP7Ckcg2WCNkfW/MxaVas+7drYMQUzHl
jSI2In850uWzi8AJiapuPhtmOW8AXGaTwh+H/tGoF8KA/z6dzOM2ejD0oBTE498ZWiPIwOZIUgwh
VTY/A6asmmYE8hpw0p65A6603nn1mu9cHPXJPHADYv3yZ5eTA8l43tOsCGCCjaPN9psxuV1B2HiZ
oZkzSuLLfU+s7FtkCakthSxqQo7TifDOD8vkGDGkMa70TfryUZzE2x7rLy6foAblFXPIULsgHEk0
SRcZkNzgn4hGO8WpnBFoSDvd1YVUtqvifzQ41m+H25324Ewq+C3e+TlV6GWxytthyiUPFMPz8etK
vhch28WLjIRHjkmyuqZ0288auo7z9SwC89GvKfBdE/axA7ZlheR2x3W7m31MMXSola3aSkE1p1RH
Ci39Zm5zVNRNUckVk21fnosXXftu4fLa6XAF6ytEeCU9xFcchY3EwP7ne87PBvuF1i9ufGXV9oN4
/ff/7F930zoWG58a2ibW8qg2y5PVB6x02lSQlxTTYehbfEIuSosc+62nvWHL/9J7Ze2VCjmqzioa
tPx51H6rHw0HUtosZ4ZDu2mMFsBaM1vQgf7rl2rwdBFQG76MM1LoONXWFRENJlf3MO8T7c670JRU
WQwNTdC7UF8KgOv7SyyGMVI7Y/lmjxw90CcPX4hrjLTMUP+WhORfAxMtOrDGaWyK3F6MhAIIjWat
8L8APDWZAUD5Sp/DCleaov5VUZ5LsU3ssB6fkPwPXlds+CYlgCTFgyo9w/Wcb/TeMkedEmorPJLO
oqpBKya4IxtAXEWBS+Rc5NwA9MPYIyN0c6NHTziNo5Weje7Xj1PQKLlr++Km7foESSvf8ij2myjV
lCzKIP1DOcri2/By3Jzz/vslkFCMKH2G2p0Y3VHIwlzGjmwVYCqPwx6FS8GfuLjyouPyEjXtDqMc
JHKdr8ngGManqXMzvxT7DND/chVuVuwXTTzBE4yNGLurKIgMzaCFyZ4ZilNLceKlDStWPg2NJ3lo
j548AwFwqTdnExc1PfL5ePNA+UgX+3bcrT6Mk1kxAdldG73fJiHjOzFCRURzNdic1aZCm6JpWlJQ
BDtB9cWEXYdz9ctJtfLez8DAHjScuxfZgyjl+e3BMNq4sPZfVccO1wEa4Sxj4Jyj7ma+uodhvuEe
dxMHyZDI/sOV9MWC/uTVB9szf09QERhFzkzn7MizoadCQM239qWtRMkYxpV1HayPJO/CgNlVcLG4
R44TkfmbuqHc9ArQVge8nqCBIaNpSXFZTK3Dh/EHYQP/UK3JwHA7+tmH8+R0bIbgow9yBM7yYkl/
2Ds2D70rD5ph02QVwlBdrS+fKXAi1CbOBA97HsdTFkOhYUp+0NeHlmbhfzjRUGOIWl8NOnM4PpqC
0aVWUJ5/Ku7qHydphSmz0lsMTI/pZy401JpPuSlgAwshByP6im69fknkzPly9H9B9bPN570AeSd/
kR51A4Twby9j13SZKvQK7t69K3iVZQJ995PUaJ2vSJzGwIEQnYXWVMC3BDzB0x0W6r9ERHO7QA/C
HAob0dzMZTnRY0W32NtB4L3cJaZtN8jlGUcrv8G5ah9kWSuRXOuQ+Nzs2SZD+QxcYpSRywcrmxIn
kp+4GhlqO8SvOjmRSnBdDYBbRcaxV9mFIRd8qagnuCNY90cTmylpDSNAQcrwWM3SZKfzx8hZr2QM
oPtfY5yOuRldauVlI/p5nbPsBADit9QdE2qm7hDqzQC3gPhnn6kqrBmo12q3XqF6hMDX9JCbsim9
FAIhEKV20My8OI1tmDV080fIwO5SoPdsoSARNV9fib5sICYnz3F13nSVU+Jw9FnenMFgpWke/q2V
uBduY6WA0b83y4FjET/XL4Wmlb2au5IQJruqj9VMBrFvfnfTk7bBu7a8hponbjFYhGyGRS9VpaOI
NmWIMUm9n/PeJJlflFVAlzdaJ48l84R65POcN75crT3O0WlhXpmSrqw6DvxI4DIerwlA8WCRB0gn
2RUPo3mla57SwzFKi3gh3orZfv3W/2OvgjuizGcRCw20P8t9hjuJUfp9jJXc3otJYOS/YraRgWb2
iT5GXo1LFT7Al/9k2Uan/xOCeJS9p0tb7Hpk8WGl8hEnzeFSpmE8rgNDaDpkHuvHltKL4aeuNBqE
3wAu3OvTgG1sSII/7Uv3qys504b11k0LnRPkrvwomKrD1cYaKpgH89rVSOn4ypApmoCqUhSgBMIN
dPJxzKJ86G+2xA2upp0oIolQs4l2DjpS29rlINBG0EcaLUTo7BgZ2cSedA+Wx2eJUv5wch/j7tfy
G8abAj5y0cPZsz35F7g3mcNES9gHSXRX+SnouBSvAQ16z2+adxc08VI+PM4aVzOE8IWVF/f1LkL9
sPfCCoe5OKTn0nR4858ozwH+GWav7HU2AXkMZk9UnaOSEl/1VIcbOWns2di1DOLnPMvYODytxfhb
64wUjXAubTYxXX2ceE9G2WxRmQYKWxHiziEbFdMyB6A4ZJPnABp2yFaUOgeAQKFFRTZAMbzHOtKp
wDr8R46Ay5XVnUY/uqAuWfDqe3znlY2J0XR6HvHCyUwpRLB3Y+H+jnEG4HOuI+xI3zUAXSJiDHKv
WEl4LQm8r6DoASbqSadQGZmOurT5+QFicKw1fgetMn+sD9ql5PrCd4KObseQXrtqR19r+14roQFN
lUVp0dBoUTjC11h5MXYhBx3y4niPMJyypM6AOz7LVYEKuOKuJ3lq5cwCT9u2U/kjo9cyuyi1N1bO
NfU2XMabSgueTXNXb/yvK2icQCeWJtsnqpnbbRASr6uXYPPQpMgFIfsAvDZa0oY2+cz8YHA014gi
dpPDgbHOsQlKCbgOsPgUOOSW96K4v6f1EFUTcoSNxEgfSIoteykH3QQcAd4LmGk7yWcVDrYIm/5E
8edEXfyATJ3fGdS3nJQviza5/Blv85L6o5RVic59bGCT0LdApz5RjKDVJTJu97cXRFf8S+VahsYZ
xKstrmLjXE7FdqNlN8t9NsTwJ+bMTSxlw+VDyulSs+eWE/uNu6vIjLq/IqPIX/P8zKR45C86Vq7t
8g7vRQ1NN6a+V9hMtImJVSxWe4yWFErrnyhnrAqKDewLvNXhS3mnZqxrlfzIzIH77vt8ODIth+87
S4CXx4FZyja8ijBx2EH0Efm9RjxvVpXkTLJU44lSxKrB2WquRWcMClVHJALWM+zS2gMAZHjj7nVK
sutzuCt66xI88ZJW/6UF577cNo7kfUoksHSbW+cGR46U+fTNTb1fReKIYe0qgsR5M8hOPQS5JXh9
BYpA+Y4woqsK097lMIrtqH6VHJnDUS7mti5QZPxgvUQEjmSFqwYku4zTPqJwUdr1HIuepDzPzyU4
g5b5CK9zx7tKtvwUCIkLYBBilZeElHuSlCTq11j84eY7YbTKmcObFEV8JfNwsAtp89B9E8fkuUcd
E5pd5OCoYbf0jzlCmyGiay5jt4o0+66OWXaGy3Yn4E7Xt9BzTn0XHcyRjKUCv492/2dqQ39HUUQ8
KYdwerH0rqgIJlOQZVO+/dx5XI2Vip/Dj3ejt48vvRti7vqoaoEoyjhJK3o5pe1SETlkBJJ6DJdU
lOz+aRlA/57RiM3AzFMs67m2hZ47uuWvnwHeLOPntIXTaOxTU5vQyICYxPxPqv0Omrf3bJu8gNB6
czZdHQ4epoLSyvp56/DXDsdOsONCuNwWhalAwtU+/AmyzQsToXkQFCMwaVIsM9YshI0wgEWJZwXF
ZBgGuXoKtH2j6Nk2tb5Srr6CvgKcuL27eP4jkOieyEwR8XRR3VbjUc0fNhXJk74VxjTYMFrvsxyx
Q96MjbtMsZyCp73ON9E2mUjCtdBWgbMB1sVtc2vBhDb9kVobF7Wr4UBb7GtTjPP1Jg4rRD0eJAU0
nIA/3AcL68Ml52O8hltl/gLo88Z7e9PU744UIFjpOGQLi9bwV5F2ndH0yuipH3EmZoYEEL9SSFvl
1UlE0aB8U8C2/e6TUZ0EECvJBghkR3R6wvzZ3m7qfgr3U0WCF91uSSuk6P9KUMRax7bzc9yQE0L0
NhC+aK4LczaU1s/KSu2/NIKZZ8iult1kGqDCFw9de4x6VZByKNtUExqRPIfAi7rOqotPIhg6Jy5X
P2I2xI5Wwl/gI1wOMNmvAK9P8M3csdigDma4Ys9lIOe6bZb2y64oS/DOYuY3ZGPc9jfbWkNArr25
A0hLxyjaEoopucpvnWOxVp0l7QK59OaHS1EsN7ljF1y2aVs5KERPMp4nDsqoJ1/wSgUIVAnqJ1uU
4MU7fqQ6r3toagZ51qBDA6C8B3oFCNjKwc2ZqVRPITMUttUagIanowlvd45u6ud9Fhv5pceg3xDs
VQn0lwPIMrBobujKe/EQ2kUAWeuKjtpjh+sEQRWORJ5pMdFRbH674SzQBxy7o1qJDwE715j3WpPR
9bm1kTmEDl0rIz3RJQryPCgEn7GCxfKUAdN68Ch2B9FmHUpDR/Wxzi+QS67LNqzEWSvnezLx7TTw
8vS8QZSJV+qpO8cPVb8DXs8EvdUS+w6Rm3RVAxe36MesL9mWJjMAH2t3FqhY1WuMFpeXy3Ad3egq
gEbSFxHJlpnDicGcsj58ziXrPkiiw50u/jgEr4ge3cGZQ8//awC780OtkqPivOoWswM0c3rZXme4
n/RRTWB0b2r8bp4b7VlwUzBuM2wuZKFPKYsFH3fjU3vzfqt9v4THZ5xyN/NMeXOmVnCNN8HWoH19
pgjHlC2uei/ZUG9i3Fw8DYtzQ7axBWeOgkNnJEHmSVQESLL6XirkVjmK7MSkA/nhYTE7ypTt6LTn
z5e8laFuwJnDcO1usTgLWfRRpNqXwUoBI6bpflJL/RZN7XOgRiTdPmIaV2glE7Jw/815olxxh1Eu
oHZQu+dPKKKBiBW2BV2+etdIIqRqeBXG/dkVKWymmfquT0y3i3LPAY0Iq4SoWSRu1FoOjnqmOSRG
qSW6xtAGO0m9ioZa9TYdys6ChX+xMpMwVr2sHaOygAnOzd7DuAORhY31gyioPxVLzTgnm71nIfmX
HWHGRSN83SyvlRlrNY2jfMzgcPPeW5X7GG9HdbeJzZtywvtVl+hHaZzD0ASpTnq9CpNxak3Vykb4
ZFuB+FeDSKSa0oBti3qaR65sZDbzEpzwIpvyJ6aBCOfQTE8bWfVKWocXC0u8wPjBUsSryze+PWTz
i9GSMhpuqdXDkGWlNQ6HxrWsCl/nWpftmFCts2pFpE7ZGRd0JdVAPyYibQAl26O7ANLxYgTgEXX4
9otlMwB6POyKxW46LJR3ianUvImuyZ/X1ND/11gyEMxUqduQEpLxBh8sWqA4XZrHnRCzEJEdBzaU
7IYJzATcrjVfP9fnH4SbgW613hfXqLQeSclhlGh9XRzS1XPUUptifwdgQULHe2xyUkEijVC+o/uk
YG0hejehaEDpkOVfpwRfXwcBMDrRfwGyFMNyJPFUJv6u6lAZhMc0ninRjx8ktbnXqy7G7P7Fgy6U
Fg/W4ZZDkqYz6oZuodNKcBVGKO3JpzlF2aoIhox4llRt1PKtjqHZ6xx+QBtYyAzHn4Tr8fzvE+7t
UssSTvJHZklo73FTri1SwiLF6Z+ME2zL8qdraHBAHObFHMhJ7t3w+PquSfu67I9QIKsHcxhcbhqg
jHvgJIvNNUTLvSKWFqCcQuE5gaY1N/ZXxmXp3zq6R2BSodDUHJ6bpGWLizVYwCvBVF08svjwJkDw
Bt16WSUFvuMBiP1Dqi53WVPNkASWqerE7kS0Q2zL/L8jG9QYcX1lI63VWruyQWusa+2BmAERCdKF
/gXBEw+7cjKeQQQLNgzdTPSMEz0GIvkhYlg1IdSfs06tIjQ2y4YoKoVc60/g7uk39rCDYBcJ4OPx
JKkfOXauElsUNy8Sdcby+lurF+mPF6AN8nQbuIRTOHHreb7EnFoeTu41+vTexq8QShfNCinYanTY
hTsMjDtnIa3aWS4RtW5Q2xldzETorfrvNK5992eDbtiNZBPci4G6O8pC6vfh4cI5/tudwOFfkBtb
S5A2xpLe/ZcEcdVglu/gpY1Fi+vS1cDhrnRazSpp1wMp4d33CBbnTCagMBXob55U0rYrsTZdSquj
jIIJ9K4oqnzbQWrWBjUAp06tPI9glyLfmhWOZGGqWYaZOHVmwsZ/ehxW+Xmec5Pr9GbeImI/alRQ
r97xLv5GGcmC+pztzswvH1LglN95GkSxHU5N7IDrfoiGSuFkg4jrrnKY1Qt3E2VJObRuA/sDNJ32
MG2ZJkgfREDWbPhTODLk/pdVREr4Lpt19s5s4rdghLr7v5lGFFCLQyxQ/y3qSINCSTJxod5chv1a
cbGoaxTWPLDk2EgA41e62+Gjao264hNwemIBi5X1Vx4SCzqu+xDZxcMfjRSUr/XNpjvNDahcUmKy
k7Kp/uPnAuACS0wBKYVJZSc5/Me/368JbpPKqG3ZTmPIz1JPQ4K6BKWxiENRC8xp7sLe58E20RSS
mOJd2FPz9TESkLx6m97lqNr7zuqt178JvRqbQf5eORXHbdqD0iHrePv+CBMZfs87yhX1Vj70M7ll
W5iQphJdUdn5SZkg8hBIPDcjeTWp7z2D13BoyR92ZQqH5RH8FFmvAE/JxqLr5pfJ1j9yFCaJrgKh
KS4jye4HybWlsSJEYMhIDp2hupP0izV4tonn1x90M3Hfp3P6TBec64zgtEkVWioGP5b0HhCrxSfq
RsaM27ch8PvaISF/xJfRTTwLFfIhFWead8D6tiE9R9YSZWKASFAFEPz3+46zeu9jl5S8WV/mPLoe
d6GSlvaKrpU4my+Eu3Z+5vFDvdX6lfczuSTrMJQqzSd2KmJA24tUDBzg7641JRk9c/GV/ytaEd5t
FO41+vi6Nh6Za9/Hi/lVU6HUx7yuCBwB68LFkU85ApETbQkejfccLDlcZ9nWWlUfy9Bz9E5tWuK8
uj7f6/9zkNKhiazHAB+CsD2ggmJHZOGrQAxrYKlzJP1mkq2D7EiqQ0NsWhqD3kQYyIcMI0mEGw5P
4Y1C3hl+1R5OsyLr0Yi45NAp102BagSj9BuM6k3fGcRK1nAenYB/l26yQDNBi7a+LkI/ZaBlcKni
IlrdVxCj8R/CuzOD3aQE7VvyfAXh8iq4ApiNnO/FC7RC5Ys18IQJ5nmgqaLQGI0jV7F1s8XeyQZ2
ET012JYThVBoxsXP/AqpcyIGI4KKXk1HsQIP6bfJM7Nj10y9KUmkIpPgg4taNVnXNyrkuZDqUnzG
WPkiNareZYHd8GwWmUBftaQayil6vL5M8DliX6Tcq9B4zUx5/j681YTiL42RQJEGv3rYkl7Fn9qm
61so51XIQnqYC2dVJWiLAIdzyXu9x8HIjqmKz0yah7FGxIxrH5IJ2PgfB7fBrgsFhi3l2LiL9ilZ
D4bj7K9/5aXitU67GguV7SG9sTYjeWl68EitK6DeaVrx1Zux8WhgjKzhyYTZoqYkjG8qSdMEUYsM
cu1FbLP4HaIjL9vDURes83fLqBomLtjertZxO8eKv52Qn610aQmkk9g4t64jvcpehvtHoTlsdS4s
SSqz77CIoZisfmjIhMHOZIkyqNTD/kp+g3b49TO9fWFENrjGJJAawp5QSOJR7B1oE+lJegqPZWtp
wZgLLyDxdJ6C5sXKm+UkcZZi4lc5UKXps2WVBH9nExEbISCqhBP8HvUtTrgmID3f1qBrP5akm5Jf
nSH7h9sM16IiUs5x0bdS1XBa/SRmqn3bcVszt34PdVOB3scCGm+bjGSLzlR3yVeLFNuzwa67l0uc
43GuNVKzQbSGFLj5c+kC5ZPbqoWo2CFuWt+Tu4cmwxr6ZZbl7r8Fb4rVG5v7U0YA4jpPQ7QlGEWU
RzNioE+hCLxyaA+FEYSbeQYKfQhN+FNmVzTi+BeD3Q+3d4RMDLn9qEZdHvB6qaa0bXETw+ffcM2R
G8sgBb037Js87WYSfXa1YDboScySFGHaFVTz+bNUv4rbOo+wKLS2WBbeIWibx3cAbkRJldKqyj9W
ji1ZXYlMYiMlwwyg0v8/EDgi4T7RVth2LAcqwDpCavEgD4ton5II25ojsj3e34ASgdTyxQ7+EVCW
lCPTfEHxXoncD2Fx3f9bEoJK74kXT6sm5ZltxEJ2Bn+yyUA+sJ/6bA8WqwRoZJYVFOKAt4WmgIEI
2NF1enEFB0CQ3rWalKqXmbcbXzwbEIvDz02Hu2TA4ry6j+zlgZxrXM61xsajzlTGjgsZiSATRo6I
CMDWku+OjI5VCwnNJ9WDnqjN1dloQ+YmYOwkGcqjBW5zNN7eGif3n2rhkcu/0LNSkEELDC2WEAuP
s3yQ/JQrJKjKsHfNFCKPk2t8TIyVOdKlQD+thCkSrM8XXD2gkw7AqJJT7JNfVDbud/RL5jd+pUj6
mBI4/kfm6vRcYM4Icw6ANoXQ7dHvHC655EAcyDYcKTQ6hJsazcsuMQoEg90wR9rDZna/jyk1hp5B
Pf06uvKXTjAdjxbMv51lVkMgaaM+296JXF4pPkmRfD+U7VIWB/pGNfnwwkkLhCAkTR68PytQRB4b
+UDEHEupca2HqIkVjki5hb/f/pbscR4syXFgYaGHL0BqNUnz9wI7E86TXOHhiXXNmQeNjBjorWoy
L4/3WSdH5Zqd3aX1SJbPHWwJ3EKxdDxkK77IMbvM+svM3pijP1wY55IkgMlp+4pRiYXUBq9Pa1Db
c4foQ4APp3I7mvacKIWA7GZfU4msjBebn2Ns1jbMhaJsBFDxpzJGCWOubahSjJAAnCEXt5IbCbEd
Ypb6fyTbYk4c9ODWILBLZtgmM/mFoIXA3jNL/faU+DCMYmMR+215J7JWQ4McMAgBF3gPTYBhDMNh
aL/FC4MfNI32+a3BPi8YzjWjk0Z9XUQqYO0ZsYPlkb6+uJ4dKt04atW3vXqFXNg9c0ZK9FgLnqvv
f6XHQjK5r9l5T92L8M5IihzHCrTy40qLAPsO5vOgB1n73tMZ5sJoWcPbYqdt+0mX2+vCsTxZNGpe
2h6SMmSv2Z+sC4ID+4kTgdsrNwqBH60H7b1oG1yOORguyU7nNmOik20nIcKozND1vswnLMelLAtL
XZs280Hr8xB7oGH3VGrdxWLGPkB2FLY2zqDV7VPmNsWuWXVOVqC7veN4FfYslOQDZ9k5/XI3vk6g
d7LrgKxnar68/JDeJecli5WErbub40gUR7we4u3TbEu0Tx48WKhNjK/zR9wow55/jhjYYiT5KKj5
DmZknGl/qQrlM60ym4+KferXxVeDmZZ2mcYX7XZNqTVrHBUBEWp47up92ZzqpJWaSMz2MNyPnXEi
bOelgM2qFKdyJ+EQzVE4EcRri0p3+JwksmuISbkJKjuXY1Gon/ukJ+AAG3p145Bvc0dpwvzE0X+J
gFouovYgHgL3qKOGDJcdLI3pK3CYg/qYQmMxMj1H92qT3vqpaKD7E9gtz+ZPsOKQbLvlha1LrNN0
8CoWZWtpOoHTAqAUUe9Wp7vDp6+Eix45BG0NP1jbYJwZ3An+ClgYfNFjs+cnug7nutueEk1RIaMt
/d/ZEGcQM+RsJMmhV7Y8gxfy+Rjbx9IO9KyFS7r5s22sjW375kUmP8wGssoKgBJFVSaWY6qTbaWP
eRfln2BZj3pQ64nbVY7h3HFnCALk4SjvfVpB8nte+OYcGyTpusIJuKRHot1aTnLRHe5Yb9dErt59
uEwhGR2H7f3ydNrE9w89+AWPZKT37VOFvp7CUrYMFmH9Fm5G7hRY50oFy1lhVujOZqvzcicMs2t4
H5JPYXnJQnVHdc7LKSssfdC3f9lHYUyocFqUNiMGJ/clJWnd/HfqQEHAV/4d6AE0oZXtr13xStJx
aawqMdf21tViu4phWGaqIt3Pbbp+UIjulgHypQ6SlvAndzPE/MObHFlYcKTIfEABF2lkTNDv6pAj
q8eVkxGOF6oRpdN+Tu9tkMJpPSdMDhcFI6xJu4mmN/aAjkigzuYcV19qDnRt1xVnC2lxIyci0lSg
gSZ/Y/2PSO81ZXtHqCRhX622Y36oeNseXo/DEirxVFW+7kaHqrRlf+5uF3r/t7CpXdIUAJTX1hUI
eQdsQoNUnSbd4DuTDT1sSn1Lx5zapYkngx08d59aJvLwyQc5mXkqwNEgbk7CRmAdm+UlYSldyNWe
DWjesGvh4QVI+tetDlhOSSrs1K6gu7myowtp6HjMKPSjKwCW4xh83v7lqK/R2d3kAXvehw8XjU4B
g7SHEx2R5odE8/LDPM+qixP8CBSUzMoiZi9zMmun8KlX9J1t8Jv8ZsLChKlO6JoK/9HvMS0V/sAf
bIsOLQzd/SnQw6j49VLwcFE7zo5LwIJADs1lK9VK15TczafNLkgpK5g4zCtds1H5XEdGu+CjqYkF
iOaxITBd9sNExFo1GK01hGlrMrfR4YD7vWEPbbsiK7D8ZcbIq5fPq6TP7IfjrWwPrnQfiE3H0Ws3
kw6NSRu5eG5Sx8St8usTYn4RJZGiyzN/mj1UBQfr9yv64bRE4O8eUWTy1ZnQ/6nsbo5ICRqnn0rp
Rks774I6WY5BbvC8rs4naDVrU/V46vvZJ80QhkSz716xdkwsW7ND8xPagMNyi+c9vMNCPFUBgHmX
FUHmfvqVvxMTzBfDH+4KdChfs6jJVu8c5FM3BD1nJv/Zj97c4TarpqimD5f8e2xIvxMxxpTIoz80
uOEgAhOwO7jEEwl9Cr/83o5fgEy+xI7EUcagdpKQTnI1F5VZt+i4bAP8X/O9+EOAWAOVCHf68mPB
oNp/iPHGK2pSxTWKBXveCgLnb5QkAaVGtB7/nGMarpL47RPclAsuSH8YG5mK4l+Im4hnS7/ZVkwY
OxoYIu0gsl6mkTLlRzfVP71Omu8+eLo2OMASLBYSF0p2mApo9UbzlgLmVV0fTQQl8mliMHbuG63y
JlPIhA0rGeSAkzzPBsKGqwBO2rmQd4HYqnP8+W3Lt30D6iwB+8JvgEBHxe7xsSwrbjUtvJwpwgm8
C9q30QpjQywxkQtAOo07T31Vwh+ANacpre8bQG86fyWlwrqO6bKMqHPcE2a8RQRSs6eVBLNRnF2n
zxgfeWvYAC6LcJBTWWjoUOGgd45EOBozXeDESoG8Gz/zTvnRzIq6Z+ITD5FXFnmehPLwU4CyeL6M
KBKIvS1fRv7eNfBmdsA7dfxkGiia+VZV4jRVZL8jIpnt5AZRzpAWWvsosTpvUNi4agyuCqQgUkBt
9nf+hMCn2plO3+ZfA6otmm907uvnRpkD4zWg/c+PdaoWfMnlf+sjppAROZP5/041uNAYBp9YwBK7
M7h9bz2xEcEZoTbOqRZwnnaXUGpyjoxh5zvTH2OTNfDidNcKd63Q1elmb7rQ39OgdnGCtr0xXD+W
8Rv17Z+q6npUComfkmbUmQZbCMkRVvnKG3KDL+/w/54J9CDtJoHMDTKv/1CkYsQ7qOSh5tmGJ4D7
N7G5FIPe03HX9UCre7zjqySW6ooxkz45aGWc75nHeE5phK5x2T0t1z+1dgC8z5tr8hDOIcxsjq6P
dIy1p22exRsskt2TKmc7VuVm93zeZ5dO54TCM87qMXDBWjBwQtKrALzRZJZJZGlkX5DpE9aMOTMD
yuuS46o3MApOABk6Qwi+hfqKiaBCyGwYJbfdzSk5o6RAHMnjoOp0KadLI/F9GBFxUD4Sn8Wi57Gq
o0X0or+d/sUz1ZiB1fpjP4mS9TeOy76fvu3gso6DYuWQcbWAqne6uK/xVuzTfkL2LaSy5GKyLPII
kNZqyiFZhKly/4hgsmD5zLzWgrc4xqonGq7gJArOnsNUTL+GxWyjtiQYK3LhwyR9vqDIjTkr9eLs
3iddjBn+c2coNZ3zj3pU6r7I0RS4iyn3X4ByufLLsW42Ct4Rs3+ZPmSfG5gQT7+g2UTtrNr3yMy7
JcRo6UJBFPGiqACX/nLFvpOcbNLn+pvbQD7zTlWNvdBmPmbjbTs9Y+QcGhDpIosmynM+wURpFFCJ
1pmY/dFCBIckkEpv0ucSSNQlkVV8Tvx4UtWrcBpC/GDzb9W/HaiKtM5kiYy95uSBwj+WTP9/EDrp
UEv8n/4Ygmc1vsNBY4bBPA5etexF8LLYA7+mLxpy0nY2tNaCDJHXJbVmYBHQ3dlk6N+cZtp9QkEf
scI3nLK8WKHB7BXpygMIa0OMA5jX1dPNOclNbaYv6Vf5gvyegy3gzmzMtiIeeXskcphud9EJKhae
QNWKScmYJ7io8XFe/OUQDzhukbTFY1GY1JNPI5VhCLFp2uFtPyY6hjt9ctHVvlGFdhbEg4VxpmGV
RFtQpg6O2ibTxbB12UuFPpvECtV8Ntf6B0/gbv2fTPWjdn6oQnkZAfas2T0nx5aqHAbAK0MBx7c+
PL76iSC5WTyxRa/k+U9iJIUmdx/5vGlSmYmSFV6NV/LQhWEd1VLN+vXLmm7GnsHgqxwHDNRxGrsJ
fDs3a8gX/5X1N8yfkx/6PikTfXFVKb55Mqjcb8I6x3yVh/+lVBGueMxuKSAzBrv/Ja72iy2KCKIY
qQiiVGjlF48CrOFWQ6fPPnLyfokEf/oGwEp3bBe2OgTvuIyd+I+JLvKdlOjctiMBrjh+bEDY4VBa
taBFODyGc3WqIF3mWTY/BSHRVSZ7xT9FAygFLwQidK/8l9vcBm2GviCDY8X1Ub1qDpQApoCVa1S3
I1oltVIiiX2OFo19ECk1PGG0gSdhWvvJHjfRYpItlOoMM8e3YUsYxHsiCMOOlU9ZkCZ3bHsJ4s4+
g+romJLu2o3ABph2rjPDSfwl6CcWuZE4fsyBuW4G1SMSi1MQYyPbh/IhcAAM5NNPRkU792UzW3go
uSAz2F4sfkvEHVxIkv1o3wCjDhrysmkSO80DTCTpDj+ofmzT5Phb8iItKJ3HPesxolxbLLACMEIB
Q3iuYLSlGGxqXp8YTnEtAo8EdvmH2/LMCHQi1ecsSEdEyNkx5Ijs+Xuf7c4Mft5yKWunLM13qZA5
X9UvuI3Oxwtqv6pMKXmLljrLgkyJqoNAL9siEH+Keyh+TRCGSHl68tze2oNWx2pMRh57EDb7lwXe
SXOT2Ju2OstGRcRJm5ISNZGTkWnK1TIjB0txcoqGql2n8NCNSzMFC48caqb0opVEk9PP6/Ryndd8
cEGPoTpr7EWmUUB41+fajfDix7g/08Cs2UzdebP/wXKkZNmOmwDEbIN3OrZl57OLU7ZaOj37yIXs
Fqm7MS1bw0mcahRIUwMVj0vXeeDx+bA0SkiPASgZm3L3+tXfM3xIcNV6D1AokoPoUApuCmGUgnSw
EgRQT7D3lhJcrnKQIcVP4f/Y1HlVSB+q+xJmxirgo8pQNDklGBsz2Svu4XIW02XLCIs0Y8IZQaKx
tTkHr4sWbnU+MiGnRj+pmP9UI0PzmYbcg3qRtrCt+NaVMzxKiUAiB1JrVRkxrhN6HuQqjAh5dkIw
rFr61+a0qeZ/ShJDNXpeygervRC7g6DOIvoGAHnqDt9o42MOw6alS9XW5a+Ev61PQ9AGqfNs9of4
24tv72QfZHUz1SytaYPNkStrLuF8mOgiCh3qoWrLd/dj2LMIr/fMXZNgU9k+90mKPeuGkHhv34+8
D3/qqbtG7YY+9UDJrKaTb214dHBItVepSIPjtHW1ko5AqV3TrcRYfHHKh/MXaNx2Xw4tW0ZuB3yI
WHEG4BtsDfLqmnfs9F0AjbpbY01b+GBX9IUlZISISm+ehuS52yjbxNEUftWo+SwxN6CBr3LDe1zK
NqilhUs8MT8AVqU2SthOGVkYu8ncx1AkJBhh5zrBdDk8F0uUmLQHiNnwSnqxx3VnGAWMEvBoof95
1sY5Xw+GKd6gh24TdF1BBKg0+UNegCCQwmr4BO1GN2k75Da2MNMI0GcFDCiRmzE906KFIOzAETnS
Zca6RH94XBlb4f60hejwv5gIX0+N2FDtyMp3T12z6Bh/jJx6VYiGoktaSUcQziecv8oQ8pk4CN2s
o9mJduqJfnSuumgyWqcn1scKx6RnVvisCt/v9Z4d5mLqi3v+VgsdYBdE3TKkO18vY0oDoYS5Mv+S
Kf2O2JTgmxmAA/lxup7yXdpUAyWld7HXFcA2/XHFOzN0J8LC1ccCy6evlUGiaP10Y5n2vyuzZcLH
qV2N4+9/F6olWTru+a4hHB5xbSmED0V3u78Z6aM+Zk1cjNpbKu0rX8oe+sbkTD01rGlBHd535Tw3
OzXfmNKnNkCMNWKWdWG6ow55qPWxAdDOhw2z6hkYGdNPoTxTPFhsFjmDfYYNMjaGw5UgK2rhNL8R
eedmi/5qB/sLBYPlcYq4H3X5WrgIej9QgSYb1wRj3I1sh55qAC8mJwhZHd110tpEreQXyttkrck0
CpqvxEHfvp/55/zs3LZPq2MQGKYE0geckIk8KbjnrEk1eBysPBRvPPCgjTRKeUFN2bIWhM7aeXXv
76kuMb/l+hl5uraryQZIoG6SoiYzmQyx+mRQVdx9ffdys4tmiUgl9th0WeCk5qY70OwP1gmPLoE7
lGaQtAlQCtMOI+DqPfZ9uXD6HIB+4PjQMiz0h3OljQNG/CC6E0Sb9uv1WeFCY92aef1QWYrQXlA/
Z9P+2VOwgu73emjbilAFyGqZEV5ckKfYXvNDG3LqVtc//fm009oiAmZNKJEvBSNUovrTCv78xsAp
hKmPGDD+gFkDIjMTt7neDwicoiWhSwh78ikxCCYw9IHGxLqrcnJ+jrmSucXGqisq9t3A6ZJB2TI8
RCgcmeGaMkfBk/x+8PBVgxpJ5+TgOolj5XpHYRjVPykZxwIO6Ru2dHIw1LFgKgtn2o2sGkIerZV8
s2WAlir1VpvhXKFxAIX7Eg9fcA1we0watQDWS/85n7Zk5apDBV52TMG9EUJEEVeALB9kPWbKs9wS
mXhlVp2pmQAx0CBpwbTsW3V9mO+4rq/RuFdIH5yFjn41EERRbCDUZlnnAdSIkoHqbgm3ztgaskEE
eRLkioIXevDtrZKAtxM3eQ6ehHYqrcXUqyrA8AoYvJg33NYtdtNguttLed/Mo8RmZuCjsqqSu+dU
kw/zG+NcWUjLXfN8NjckMhx0f3TbJhm5kkpYBGafO3KpKAz8Szx6QKQ9eaPoaIw6ldvLdab2HKNh
NwTl33/Di9K1xeu/4tt9tFJWACkl8fwGLPzNydgG03BU7b4cd3cmjmSCWxsW13bNMnPD1t704Kxs
rXUmjaE4IYExYWQNqFAwcpkJNt9cL0lEbFbTTAQTaD6wBeCRkXxi4hR4o4l28DCk6R95O3mPACfa
gnuBquDoxTqsllrbOkWH3o0i/okSC+6FrSRdVh/nkiuFzMIYwvB/En7/Y0h3yHUczJ9DYGioWbYa
Z3vz6BKM0zn+XwV48eFgbh+m7CfvUQu0keujRfp1zhJCdAHe0qPynaZFe/Xo6wLWWUU7r2cjn/ec
aR+HwM9c0x40wbbqfzGud1HBs/d+9V9Rn/bjDQAnKBTgBN/Wd3cpDjDJ52YY/DJH2grt8GiyK8hl
HW1V7rRYAea2G9F+TLMCqpEOiP03CJWlv4qmzWCmwuzpva0BCTHx469g2qb4eNVQ8VB1ghodSd6j
TW7Q+V839qObWErGDUCAjdcMPVhh921sPEkfO5xYPwNaY/hKFIQCYmb5FDux0Scy8KVS5zXQcHEz
2V0dCLUwrgQM5lkYYSLtorY/x+Qwn2vT5o8VPzkR4N1XfLO8klRtU+ecOfO86L4NGddLXNKbBbUC
cHebUIf/9D8Xt6/n83ru1aPBaPLiLCI8f2eIkzr+/wNfOU2HWq7NI/vOKUg5cXfIJFY2VKCLRKHb
ENwiypYoWvFYy5ads6u1M+Fovlmueg+kEKTgzw1559E3uPcuBU573UYab8NDocr3I5tkdX3v5203
0PUN27UJwQkUQ/K3Z/sItVxNTGBUEsl1wAGbFkaI9FkWkJn+fT9VO6490Vg+wP2aO92bhH2g3ixQ
j8sQWnoL1a42aEhLmVNTTkCiu/pcKGtM9zDMHOdDX+ubnLOu/zUi3uG4nTcc/OBtA9jWTXYQDN1y
Z1XZdVpcT9DHM7LdyV2uItWuk7yJ5ng2uHdlnTP/Gaa+z7hlTNwDlWbPYJSDZkF3eGWfvYV9vktc
NKNishGJ4LAhIpy4E+7yf0VgzhrvyW/pU0yCt7YymTqmSV58Qb/mW2asz9Y3OgvvopCSv96clUWR
GxoMs2t+aYtOlkMmwnhQniDxaOQWyRo4v7AYR+WbrToT8cwXCpOKyTw3JV7PdB8Pa2OU0S+kBsmH
E5EW6/RBS0UGrZADnU/xuQ2s3Bq8ILzPibfNP8yaF4Q0h81tCzNMj3rlgotTMqLsJ6sHSs0ZygRG
Y+4nLQMvFEhgJG5quP2DNL/DCD5LfYdmDW1TwDTjH8r+5mFd8Vzn9s5eDsko5jBaTcsIWDMu7vMP
uGdc6bvMVpGvBl2sNZQ1N30ZuycWq9DFfurl61/olne7xIHk7t2FJn3JrRSY0F2qFQBoL2MXP6gF
Vqxjcp4ehHRF08EcwEpmrntitfPWmi45uLtPtj6fqnIzvX9+oA4bPVhlmePYBfZ8i4Omt/80+2zH
eJgEmeWhEZ0VU1gvk1EcjOTy1m08JPsI5EMqWpBABUzVyueCWeDcGKI8c1YqI54aEO9Ba/OZEcog
Pxs5cej84V0TPuaZloJXN/4B0BOmt3VHyoW7FZaMd13KZq0ROHklCP3uUmgL+kP0kYdBnqKQRuRy
yKkcOtPgh5J81TBG4p2+Q9czt3MrHBW69/K+FsPJ96AF3dxUR/5plLNdSatIvJC2Ggc/ju/KLTMD
t4Wt1znrmS6/TUTFldZCtn1fFYAA4paCJpp2a0jVteFrle/IhT0isZZaHo37uKVgLuTeXx0wNekn
H/tqatghgluQDARyUJl5rN4aCd3J5s2ynRx0wWgXkx9UmY/7tOMzzpoKq+W7YgsnDWXv0AeGAXqV
Q4CbzvU/3e30TPdSgZqLUT2O5/gL9nmTbdQY7rmmkng7t0wz7CzAcIaoDzCKjm497UPQluc+555i
ddEps97cBAtjHlCaBoOo8uu37p+m5eCWOVGwp9U670pZdRIVHamP22xmrWetSBNAB0xaE/FLPGqZ
cnwKVCAGopaZEuwbbfpWnr2X59rkeCFwO3E4xdiz/JJ5D/H411av5oHPch9itJtmQDN1FD/UhiNi
INFU3VCgfsRhRm3hZZ99XHg7SoqRVIIVBd7zU85cT9Y2d3X8GVsx1ADHCgoMT/gqB9PsBoAiAYmB
8/Rf2QtHEG/PkybR8YDii9h5g8eKiScEu2T2zP5mQc92BCwe63zaf3LzcZqIwAjcyll5uTSgcTnA
ehupZNJRTMXJs/qGdyZHFdWfiPU2+phWrRPnVUQp30HTBeeaCFnLezb6Gr9VohJU4berAn1TPBOr
8AMs04hLoMpTkJV9razR+oV4MiV721fD8GPyOxn/XU0GZXNbLrKyCnDFx2DteVk49A360Yh6FvlK
WxHdblcyPvpHEbZyv3ctOe7iri3MasD/thzSo7shmj/te/53dh6m5RcLvnZRNyHPzmIAT0fr69xZ
V1xJ2oAAxXIilwnnhrJqY7OgIDJMVNp+/Jbf8Yf/WKHJqcEvtQYx+O5O8f/PSjHdW/uoxh3ChDBn
4afrgeF9ysIjvI+2Hu9CLBeMueIB5aLWz/8eCdBdlGqwasqHHrF8S9blHAM6Ji9k8iCy6qNQNj3W
WpZ/fRVmnYjF/2hqSnxbt2/jkADE66Zs92yGJGir4vd+XYqJOrZTB1qYes+63xO2hwDNhOYzNmi/
+W2wqRE6XasddGuCjkb//2CzEBN1YNmwPTSi+kU8hyVMncYp4VvGcE0uuS3rVHGSjWMHk0LxqAwT
4pBWIDZ8U8lKk4z1unuU+BsSuM6U9TjUpOFGVz3bDPMPZcHstLr+cIb8kwE136PKMCu644lru91h
7CyBms803J6fKMZeBYv1faKbkR78c/UWPdaAsHZUJPFdeV4ZeGujrE53gkShfqYjPDnZvesnfbMB
TKX0fVBN6HxKdnXTEym7Y4ULjhTby++wmi9CE055mjICq8oi69l0sAldlquSCm+HMHGsBIelB5xf
2jyoqd4yc/p4a8oyvrxojLRF/7Jw42/tHQz4MTDavslJ59gya3+d5vgs/89KK72f+6vS0UB4n4ZE
/nVlLs95ZH4xHbo0K4FuBbGC2944cH9+Qe3G3e0sT9xQJKIQOFzdjPVTbb+hy/mu9lmA8TuvJ8ql
aE6bzfajRM5j/ImoyLvUqKKzxUhUZRGiUjt6r+AjK91bwjQapjLIVcKxRJJpPZkkMBeyhI3T1jtV
sZ4enyA9WHiSqoRbX0Bw1QKOx7Nb5BvblhjjtDjIAmPd84kMP+k/Pb5JUc8WaDArA4mZ58fGHKjr
tj1p7TlOrz+I/bnZTbJ+VfLhRPtJR2BGgoCgeVQ7LDyhNyXnlt86mHkvmyiV9MdLnqGqDNAM0U1I
HWUSGdjYT0tTN0wU1I1oKVrSCIfeZCdKar4ONRoJ3wWBBBZdC8cz4WRPLoKd09BXwMzpyzraCimw
7F7MO2zYaHfc061V9VKSVN1N3bGy4v3q2TGntgoQ29sWWqCKXY1r1lf/r8azX8aJly4eeOBNgMUI
4aXu3a1fGVumn2M87Ky5dP83DKhe1zUhcb/DuSVHP4aFw0E8KIll6jQSxNRe0m3UFjdwqvvM/eID
AqhUNQCCCBfg5fCZVdGzl4k7ofRu7SL9JGr3ZohOYSiL9Ym7yc9D2xnDY6h2DYNdi6k/FBqEI+qY
xTvZoSurf53OY24UnDHv5DvvKfqCyr8SsZJJZgifgMTEQcugLhhMsSafqxcaamRLc1eYTDxzpyZO
oCTkUbtNSrolWOrt64AYTsk5zRtwHBV1yiqzLHF/GoZopN+XtdMFD9SQ5Em0iGL25j8Ao2TjZmz+
dR/xZ/hkwrY7y6xaxdlIGWutRsdp+28teTV8JCb+aMYKoCjOTgvG09CmVR+Uy3/K5ICkhoD0xL4d
ZsvBlxhqV0M2AUFN8VPy0LqEizh+tgpaJDaHuoUgPhLcjrmnYJZe685jgC/Tge/g4UM4P9fmMGUI
MRaU4QXmzqWlooGcmcHDoMipml7JW7El5uHN+mloCLeXu0cEnfwU0i35G3PZ79pqc0SMfcbChcHA
52R37nza7NIc+1SFnHmNEa6d12O7Nr/IPYjuxOxnhLgi2GabkyF1tZMjOO3cHH0pRiv4+8a4tzUs
XQs9c08Gj1p2QlJSbw+zRLX391DJUTKSUF+iv+Hnqc14MHr7HlHQ8B2uLMjlPq9hMCnPxUSn4yEz
NlqRvR/lHUvdP5u4Y3djWuQG40z2ULBLMcZZQVpWg07CRr8gPeDBuZTxbQHcGrMn4Tyy9k+LyP7i
+j2Pf+pxVmcUoGBhLzEBd6EnLp2BnUA+msVwIKty/Hc/nSbdgTztnsRmJpnESA4qC3KKtvpBV/cs
6y6+H+nNORd0y1u7qqEVEuVALEkMZimP8h99mQRFkFj4NpDyBysGnmqiER2hlgtx16drW1M67d2J
uCerYEVg/+6VXjde4tqEfISDP6yQ2tQeyXllW38eoxueLnLu9znpu6fYlgHTo5wiaziNwfn/kDi1
LneNPSYM17CkThZ/GHMgMCOXrSj29LL9TtYOwo1kKoD5iR+0SS4h7hIxKrT7x+oWa6uXFJ61g2zV
UYPdLvg//JfFyIo+EMsKolJ0WYPaV6lM6+LpfIBlQE/bLjmpESQR5HtVr4oJxJeTtkit7rwwO2ZT
AoFYtfyDLrMYkFvLBQONMA0dRTl00CyTyS6ZSN8ZRuNJphVt7uQJnz19MB84EWz/mRyrgJ2ygNoQ
Aan4WHSBxIfIeB9T5o1CJq9F9mBhuqmslDEPul4iH02gEzqkKfO+rf/Gs6HCyZFYH6ukoSEeADl3
25VDWGYLzMZtzjV++S+pUSBx2r311gmXkTPGQBKiwABU8S3w7RetMBkiR3CQyfS+0pLFzPj1ruoB
qR7dT67tPp71EPgiASB6xG1PGl/TopTDbDhqiFb10X1IZ7rDYe9iIGu7MIYt0BWpJplZgyHe8jtU
U2gjrJ4LuJUwqnI7E1LJc/t2lZNjR6Q2o8V/jWz2N35LivHAZccrnnLwzbnj7ApMmbo0uF+h1SMv
DpG53V6G+OWGkeBOpQDU2eTuUhQ+mxotGp3ACgWqYBahWzGfuXh02gfC9LLsd6UxOEpZVHi1ccic
EEPzNti6DwnkVdyDCThGZvehxvVl89D7/w/E+Prb6Td3mJ8Zi6tsG8PX83ei3jZFc/0vfQIXVQJV
sJowhLh3zw+2M3Ez/KSrBUb+lruc/td0LG4Vt9f1usz8bVi1ou+oEHI7g/yP3wuVTaUHhI9/dh8Z
sApXK/6K2KvRlQUPZi4TKLb/+CFXcZMZDGNbUAH0pnwENJbdjNmh4z0EpidYPqa6ZZBmjDMixIpH
g6FCfgxPTVLCXx0xJ0WqAy1MB9/ja5ZOwNodkUoRX23DLVzULmIVWwyE6en4cJrvm/7sirNJsuQs
Vu69PnSwudy4rcgrLR5oBulwDnWvC1oi+fVJMWcKkEC+t7xnNN0YE8kELTaiglqACm4CuQFhlFRQ
DvMYur7UtagZS4B/L6q0jgBSmFdx6gqDUIbXbWYw6/Tqh2Oj06Mpfvk/1eolyypVTLOxnl5vRSYd
GxqVpRrWt/yXAvNthY9KeYID9rw0cHbipkzK/tXJshDSqrsNmJirDmhjDRiWeG3sEuQPmdSMLo6q
baGTnpoaxAl29HYi2O+CODvzv9U+zOJnlD9OyPgoR5v5NSwAZ8QIVM4sxrMmxwVkY3fbUJ6SuPOE
R2s7G0g1A7NsIQgjfs4uiUrQj+SWbliLGrAHsuGdUZ/xBwd9utJOlP6LoMujif61EGPHAPFcnND0
8wVqOUiW17tB5V+99ICse15Fn9xR0DC8eXWWR1sEtcP5VypjSBtSZKgywuVyuYYVwN+5HWaC+xeQ
Z52+UhZS9a+xAoHBzgD35Z4XJ+7YOck4l7epGjYQH6Jmtq963ehDMq2RK35jONOYijQpZ7MruCKX
LXel15sjc5eYPxlnFGPx/IYbGRSSxet4qgHUSeOyu4inEKbrKvGwLAurHykK7nOvXsGzSZzBhG4c
K/SjyePxM303rikiuZJQuT9buBoMcX0rEaaAHaVYTI7f0nHsJPVrClnX4fckbUE4RGfnUrLVmc4G
RryB1gOV+kuwLLhYM9xpjgx7R4KxdMRFadfM4akId1jCLBr06hSOQQvR90d6FqfBtbpAzFUkoZNg
bBL/sZ0Qm48E4Qrp+s5kvpeblp13ZRgzNAIgqjFUfk12e0cGhhHP7cOoOJxeT5RHIu/wM7Ac5LT4
bNmzvus4EWp/em6+gCM0CkbUlgKLb80pIvaZllSYCdRa/H2e639rvV80530hprvyVOxX16lvAa9W
UlUYtT3DVF9SBG7eEWp6EcrIASLts4khgZYV9PLcK3CKvFZH/C3F2n/8g92m67SwJGzCQKI7WYv8
7kBZkyhMwjrj/ZmqAth62ICNYo8owMQOw4/G6ihcR+8Y61pQu3lH7yROYjMMh7vYtXbM7WEN1tWN
HMP1uzqnEsUzbxMFXec9wBTxHz9mY3d/LfrvtTKdS6I8XoN2koHwQ/QOrWuj+jsGIpphcdxzgM3u
36XsZqUJ80sZHXoIcXyEu5RhhaL7sNPFCKk5/HKcIYgjKSjUAktx1KClaUDSm1fEIY7SpMi6OjiG
mONTCVQ50PZgaM9jDaAxR1uI3Y8v+dgq8DyRLTpVPDqfcKQkIsGCys+Lh58UxM2fPjvUerWtMITc
D2ZBzPp43gSv5eF5QMRHG1fG7eL8fDRC+pleOWHiETbFmX0hKgoDTw95cYJ0TknIevF5uYKkOMj/
48xe5GAQuQDNIuJ5C1edgE6Dk1gufFD8Rn2GnScvqyPwtno3xHwuVjbcfhxDAdS27FNK2QgWJIUP
ORbL+UXWJnxIaNRYCqhpegcTLRbxtpCWPegBkXJv4Y9d0KQvU4tn1V9OjKWsYJd6/48Jc+Lu4LtM
B335fLrW43iWwvhRWF2+r+0I0hQl0NmTDCTmkNjXgnbSCnlCo5y4P/muyl6rLeoNvFur9cP3OJED
2syG8hI9xbjDxE1ddE4dpgm1h/MvwnNKYGtXAXZrzlJmv9dIYH8M81HA3e9cnNWQkvao0N0+pu4k
PCbdnvfDbshqUDlZn6RbkBzT3/IB+dL4n1p6rU/VYfZtrnGBBs32Hoon0aVC5F7EXJdStJTkdWkJ
ktEZ+UVMmM2q4MOPw/grlF/uhnRYGVFo+HLJQVVel59rPfDsrbtoBj9mbfJRb0UOYdk9O22sCGvd
Lec2UcEgurxpP5DFlcuTIVl38zh69daNOsQuRsWI0f/EUZOfEIgA6HDu4bq8rx+zm5yJTmciNDM0
THGG59NHNA82xW9+ghAGGcqbEXWHnVAaZnvwRRYDHhLDjuzWvkeSCTaOd9rhSJW/Uut0lhtkz11v
EOFmBHOhQo4g/nxaOvYx1RCBLlTZqvhpFzq9jr29/MW4OwrHkSD29PA0ca99yTQRUBxhKBczrR+j
HUBxy261zK7KnT//XK6KcgyG6FGU8StyQ0tmCCwYtofpQx16NAvuxKPS9w5z5mlf005NtMoT8AfZ
pyLwZ4ls+A1/VjXuEEV0gDIb0ny5Hox1+NJuvHOi9bIk4yvetb/7wBxfJLi2wrnIM2hZNBX6m8qU
pGWiIDqG0JUbkNpwzRTwYiZqy66Nf0G5m17ZpST0y+CeXQERBi19V3D/29o/fKuUgwShL71G4khW
h/roCAMNiaulPURjcxmlborSwY4PxoJaZUoq/D3YWv6Zt7LgbnFUbq9N5qIX6WfEycPY+seprAnL
7q0J0rBdezLs3ZuavJPSYjYhBHVoQSQLNFH+Nw9NC4BPiqFELkfS/So1Ytuqmxi0yega5eq0WxNW
zWu7mddxx2BtekheeHsd7WMPVw+F84jK2T/9XzBBtpYqMnK02NR/ZMhqdoeAH8219/iEwK28mnqF
5GpmR1kRVd36BMabbytlOsBHMTd5TFNmD9tosKwba7DfFa5IXEcDNKUsJ9+vRPIAOw1UKyC6Kqiu
5VMCKqmrFAgUzwU7l0ARvmzyUHVP1xTYnNuz1QHPpIezhc8lxd74enpyXtmq0VOSr6ignsAAuDCi
oNQ2wO48lYxGaeOu4xRgcsfEwBlMp8Aa7G3IDWDQUBnopcTS+0IsjyZF9alSAQ6KebfRMzPluw4e
NlGr6+9XUEWsRBz95EwJevXGo9UqoPmN1y5iPGFFEeQ8JcF4eSEb14ejklBXvzgFnYf7N16/cZEA
opNldXryWUNyeetYinDpNYytTfNXyFb8bB0wN3Ohkx28zslEzGurEUkC6ULqPWwL2C5E+MVEeWBj
xOPCi9Aes2NSLcrlTfaQVID0TyucFjdQW+/EoyCahAgzhWN+wWmgXAL+jgKyVgM+dkcsVpCFC5DH
Z+NlcCg37c/I1PeVRgdTYXIhTZHP81A/dFhXEaKuX/h6JFhGWK3qDOc9DuJnThEnZRzkXpj1CdgZ
qb/GrXBSKdtyGaW7+7DdW4x7IP+YWa16mdfDLW/ClIPvoktra64BmoWw9l+ANiz5goPJpVdZHT0t
OA1r1dYt16FgO0L5mHct0BA54s43xtsswwEsEY06ggQ03NonWI0x82eywkx4HfkOJANYd7+oVLMJ
HTnueTIEMV3d5tGjOciPlv9y1M3thP9u9UYrtluOoNw5Vybwe0sU0CqVNieFRIe5lZGeOTTEPZ3N
MQV98d1M2gyjT8HuwZBkhT8TfH37rAzseAswm9tK6LsFptdLklorUpbOtRXzRW9J5dI6FCmUSQwX
kVcivUr8IHAIe+EH6z0CylQw3DGB+rUiBFO2bHaEt2JYcbRQ/+VTG52xGqpYpBxDlCW7dI9Urp0R
Lwyzi88VHS1n//qPuCyAaVi/lLXnzsHyAw2NGmBukovqq985qX6sD/BihO0haQKvYnl2tU4shEzv
Czd2LaGtOO8/kcF56pJWWYTp9Prh6fQOSW5njv2TBzZy8r6G4D73SlbeAdbpUW4/Vr9cHJRNHp+r
eDKOZho0bJo/vhi9Ymsnjq4+D5yjyH1XZy4kBBe6q4I9Dit3atZtxhzICIZ2kq+iR34deGg9mI2P
la5ZU8v6P78Q7UMEih1n0P9Pw8wYznE+vRajvKntMCFTzFTn0bVr/MLSELbhO6kTGiow3WoReOnY
9HgW5ppg4q6FM/t3uAI1zl6bYeAvHKLRofGHrpJnLnypBKbjJJs2BYvWNtvRkuIpiNAfMERXGx0u
YbfmleW2gkPVkJELxqzmFG2ThLYLEPPBdsjvj+Q8CYLzpzhNNXaC6g3vF6uHCsY4i+PUz64Hb5du
gCq/VYKrVkCcGosapz7W5GPK50GH+xWxow3iAuQdsqMUH9Sh0le5VIH50HDqQZ2ALcyUmH9fQgW/
f37ZPif3MZ+TjYMSLLQU99igWeWYLvImhzaNaHBIOi3QwwasDNWPpUDRWqgCwGWeusy7I+N3hQka
pm//yQV+vwKPHYB183qHkcEvaj2vo6ER+2+S35rdc2XDHLYzc+Cl9mKTygOPvgasHDHmYuHuwmIT
dThX5mB8/VEM7nAN1yPCC2ZxVrdHo2N5eiCem2qEgHAigTKyQhVt10rzIRq+KNQPNSYdBJ6yrxSd
iDMRsvpuIKdt0KzTHVj5Qa8sWQhUmVSUAD+KGWWkvqoX9CsQsyjz2xwo4EIgTEJLEiDRSRk2wOMQ
yaTroFTyhinSnvClg8PW7+RVuZY+BQltkruTdR31T2KvdjLm+I+iyBN4+afiiBXIRlyHHhQ/FxIr
RwSrzfsKCnV5tts1SoK/jFFdBMeCzSikxURS5f8ix+uKxab8N4ky/2kt1VuAUF3B0bB4NaHkxR4I
Yss4naDu0BfhmmCU7KRmrBT2Zu8p7rzgWqa8UGUnUrELcoQBRGzlQjCjS1xXqqapCy//TIyhjUzL
gSYa8i2dmQIIQ82ZpiFJzD2NYaR2ZwM19csv1itmXTojXoNjd5p3rcP/qWt1jdqBQPqdl4r2MKPj
lfRkR8YATYVoMF/uQuwUKFA89u5JZTupzPL1Fy38MGEAqH+KzOfZUXCUmZ70wGLli6UOXdufJgqm
aMIA72L7DcsnkediO+VyOojwulMiZLn3xfTwlixySPyNdcjeiIWQee6pNZLgWGT+KlPZ3xVskZjK
dT8Rb+I9KbjlAEVxoKJ5Dq21ET4g/khdAg1KX/EAHtOFdxdndjVjwhPZGuCTLFElwfCP/XCXJFUH
9mdFSC59Taaw/pQinPlFqIfsGVw7+gDDbiKZTpmmpWR4FLitUquGB9soGw+VeHJOgmC9oRomLbke
lxBoktH8fEOwWsk8UMwDEYBbWsKuColZrjXYD+PPRC9W2mLNevZObrGjoaO95u+DUWB1xhiXNXAr
91aPJAxiKUL2y25Rux8QwBrhJuI4Z9Ijh/lBDiO5xJcDQHyG4xsTU7f0BdMorM1wUaIUgdlXed19
WA57Wy1LdX/WQI4fp84NjGMqeOhM12SZgzfKa/NcNfVaWSCHRoIZ1LmbxAgRxtfvhaG7jEkQ5gP0
P0cSIqQdPScnVD5662DlYeMGhz/7l28MsJByXOgeXCO0KPFHJdY2PqGKbbAyYucGhB5Z2A9ptZ0c
mB6CLvqpdj2wI4/QxCwFta9K448I1adow9y5YTjTyqyb6ztpL5XSsSS0PzOYB+qz5SGeYfm3+K12
vxBFg6cOlI9765WLZ2T4mxXu16qt1STUS7udx0BW3RZo7SxlxLVwRby+jR0FCONT22hNrouC9yB4
H4LokB8pMUnW3xqRC3fWUPLXX0AVNxlVLy+mbAK/wtT9t47kFje5IhQsQXj5VejSoZGGYHHJTxlD
Of22+oafT4+x05oFGED2QtLZvUBhFI36kpPbi6ROvR0gXlqGFtFXCq19HZIz0RYeQgwS9emCWPLD
szyI6Gbz/2xOh1ddHMo95/WxM/UkPHyWN1R7A2CJvvRg/b09U9nhrP4NBuMU0BpnQKpZb5LIhNEW
pPSws3KTwvDsHd16La+5LlxdR/6zDGDttbOrNwmAqTOQ8O/AdXvotZUSDiAI9qyU+6T5bS612cWP
l8Bwhx7d3T2EsyJwAIg21OyKXddLmzAWBdfnRqwJ67C4a8If8Wmm6W113nDUauysCNJKH7YdMPqu
O3ZEvh95Hbz+z99+C3ExVrSIGRorqLf8b7SylZeW8+ficvhkwJvlsgTYLouph0ABwuKejLHUVhHI
EaYBj6DXYOd10gc1tBuz5iTHMDjYiwsbicMwnrfvukS7OPRJLhEZG3RDCOIknKcTPqYea/RbMMf2
Wkc768dnWZeUeF33LdqENcvDdlwO9WgcBrV1IgnZGgkQSzYo9kcWU0Y0oNoJNp+mV/Orq62vFzum
9IPVyXEzbkebUuQB+Dg+H9Wmbci5oeXw5gtkU2GRr1VYKmCnHg7Lsez68lOxQsGUHgXEu95PrigJ
0gF/EtwgfAb2d5slVGHYmG694kbixTEEie1yoAg7Rw67xl9lZH/IIgw31NAdm7rM1/r7RJ1yudIX
ef7l4ErmHuZI9tCvk/BLgcxa/j9N0s45E6sox72PHjjo8LHM0+Kb2zjpW4Ml74MDxAKdM8zpgoao
CposAa852et5C9WCRhxRRwOzrjCTjuhtsCLLKx2lwiIzQA4LW1odHM393zSJzIlrOQEa58Mmho8r
BNwrBHInNKxcu3FAyU6orX0XFlez+RbiDbNP2l4hIi7PS8mALCAW0/1X+8NVMcrEztLTB4sNzsLo
iH/xpY5R8WgbPyY0ftmE4wvh4fOuUxdpyr4P5jfxQkbM49rLnrd8TbrVqX1NisDrR8paTVkrbaDR
iRj8LdllzaIPEVBAJnFaBzX4s954WTqRMIp+j8VLxY+sQD6zZUpHV0aEDxIgoBNxaXyC5v7DcvMc
cn+yO3jVfLW6k6ZgBlYWEfdrZaMUHyksqxLVzi+hBjBsDjAc1CnJD/Yj6ALZJip9hQabtc1KRMPb
hEXIXDwQ+taLmbSuk9UvtgRugIkY+lLyDUxfUcDCRZKghQvESu3+ka2u7h51V3f2QQwzjjF5IK0C
ZasYBuz7m6hZHvL42Ea+aND8O5p/wuHUyNfh0AwDW0chzcvJQ7a+oNg/sphU1bRa/AZjZGQ5Mqme
TLyOayf8FpUC5L3EbSQQE0twuKEBrZ5bztUQYtXw2vb4ZgWBhgtvejQEPwTqCAd7GYmJiKBJZGr8
VSUg0XkNhEnn188aF6p3WHpAj8EykTHLxwxuYE0sSI6kUKGd6XHfXNtD8sn9Wm5jScnU51wkeWIf
fd2PZrXvpxIdLvUeNLxLFgn/cIAC9bZ1ZxSezDqM6tGNOTR6C7iaFL5mVY4l7FX98z4TsB+Sbk/n
ZPCKAcFZNJ/j/vWbeG8PXc+fWZXHYa/x1BTrRmDQt091nKoqxvqck2PlcRYR05iKtvjOSgjc69Vv
L+Uw0TJPQUQMx4vy5BoPTfXuJ+TDBGmkMWI/J+6rdAjKP1VWrWXxPgfeq3DYVL0BnMYNbZE8filb
Oenubkg0qRBEl+270Ywd5+j14FPxzsaka9D0g0vzBso9e5B96fhUd3IRMNlrQRxYSS1xUb4emfm+
qs2HpHZRAOuT0jY/teYij1BhDRo7ocUpmTnfpCmCAfwTmPh1o6hgrsoTs4SLdWc1eonVA+PobgqT
4YY1WZHEbwwTa60KnQXrcpS9dlA41VDes1odZhYhS6Db+CeO9kr7R7pp9EmmkfFLmIv15Bv6TO36
a1aOqTGD4DvQmGgkOApl9T7WaXc2cc+spLQ9bd7crLv93on0aatFGS2ZQ4w3NoIeXnYyIQSeJI3r
/K5Ek5FQUkeIypP7jaz3G98j4M2GnRx3nAB+7DlCfHLc3P2LFTF97D9+N83xuVVYCzg0JSnAfa5c
+7CrHD9DlQcxdXI+jLyGZb8bJuVn98mYjAqNDnIGPktIg1Yi6iAkLbgVGp9iXBtikFmV8giuHouo
bCBAMRcCDXRhJeUlsq6QWWUyo0QZKw46veDSaEORAyC6a1+B6vU1ON7atWskLOFGig0ipVxEf/GU
d2B9pgZBJ6van0JMjRGqUYLdxVj/xhRiRDZJNYJzVe9zw4cxxuTquQ0QD5ggUEd5PckH5ednYX3J
dZzm0EPumrSPYZqHBmKI6G4AhO/s8NofyaekRTughtU1F1U6ekNfBzWd78aTmjOOcJWO60zVc8Pi
73tbofrSHJXlrcMj1QOGZ7eTn4XRzp7yQW4XEhNLYscHP6J/0Ny4aOGMisHlS5JqJFQfBWVKEiCC
5am/6W/hM5YT6fGVTs5Ijx3tTZDBymFtgFal5v/5MYccHtnqWbLNpQfbpMfa+xjwqNJf+L8ZzidY
vF2R5MoLMwoXgZiH4ezkyaZGP7F97zbKV/fyyjn3SS009TCXC1Q/SlDMxL3WWkfKaOAE/E9bZ0a1
aFD7k/R39KkVDJSGyQKNOlPuuDM0bJ4zKZZ+4B5vG/kuYkW7wLJb7I+4LMqIItfWcz8tUbPkTYXv
j3FsXEB/X3QaejZqLeZDILQgs7cJ6OmjC9H73kQxTM6IecQSl95Xa2zi+grPe36/4GrJ8bADQsZF
Fa5O1+lSxkjhIMjGZnLMW5CRq5W/xJ5rtQvsAZu7YVkokp7E9J4JjgO1UgRpSMG4h7bEXOKUOg/6
1ayB+8fylvnpg4Sy79tNU4LWE7oEkp653S5qWDOemLVl6MR4TN+wtCx5RWTOHAil/vj/rhOf2CXx
uEVx7EItgmRpoYHjhGB0yW2R5saT+eSpp2KHONgFCKDJlDm1tP5iFS4wBwoPifKzm14aMw4sjs51
2A6H7LMlSpLOAdO6iS7BcqVUQw0CKvbDdzY0jxc9x4CAPpsDsRh48ne8Yf35cW8dJQYcNcTTJYgs
je23jJ8GCh62ZcAo6vAp6JtKtlWIe7hVBqxthofcXriC07ITH59ga7n6U43WkrU5Q0vzbw021pkB
HtFgWHGhah3noHZ4vT0=
`protect end_protected
