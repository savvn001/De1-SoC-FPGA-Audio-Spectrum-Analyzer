��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	dm,g�@h%I���UF���!�/G:�~dZ��^�M���,D��O*vo��W\6E*��SQI6��$�B��9HW"�q��p�xt�sӯ��`����Ȇ�B�6Y*����b@-\��IB������e~JK؟�m����e~O8���fmCϟ����H�cH��Ԇc�EAV$��wX|�����i5�X#������ݑ���f�8�Um�K}�2l�~<y���2����������ccHܟ��H$ ���0����èH����~��!�a�b�@S����<����(�ϩ���P3��~�<�O;�㷷JH|,�lG��IY�%G\��Үᖥ��ƉN�(Lu��W�1n�ӵF���,���݅�W�3������e��H]��8@WEST�[����!����f��[��P�?̵r6�+��#����j��
Љ�L]�����U��c(�}�	g�E%x,~ر��� ��@�/��-+>6��C��N��w�1q�1e�v9~8lǾ���ѧ��jm>���簌�^��O�N܀���Âi���������L�{^��?�\��E1���)
l�#��x����_>3�U9eSѲ� �&�ۭ�RC�u�pM���;ѻF-K(8�ч��1d��˧l�X�*#���K����U��Q���F`��@G�u���:/��c�)i�lg�{�W�	p��]z؂h�a��W&t���(���3�S'�[��(Ӧ'3������i������#ʅ�����/���q���Ε����U3�I�q�ds��w:�j}??H�>�E���e����%_s��2Z�ak��m�\�쥸���Ⱥ�S�I�Q�4y` ��M�,�`]��5�G1Ħ(�L�Ϳvg�}�m�0C��b+H�#��oE�ux��e����SH"���j�����v���e:�Z���c��3�SM�Z�IK���kث_:�?s�5���O� 2iѕ��N{���@K�}���>a�3FG.���%#1����᮸�CD
���"u�_�y�������ܩ��q �
�:��K0Λ[���=�:1�2�����{�T�;�: "c��X8� ���
0�(F���-��\@�ʓ�oA	"Hm0Ƚ�ʘ]q�}�i��Eӝ����7i��D�p��|���ǌ �=�ToE�#�	��VwFо���D��
���<i��Z��)��6匾�>���� c&{�G�ϟBG�K�K�Xκ�F��2�Q4��l"�q���[F�8�ϩ�I�8O�hd��hd�J`8�Z&��O��W�����W������_�\�S�6���S��E �;�K툷3Z=`���?7�-���'"��}�� ,Ɗ��椶4�@{\$3��m4�h�'�E�	l�a(=3�O�*c�.�����k��,Z=����W3kdg	��vx���臶+Q��L�EbM�r�J� �!S�$�n$e�h�����㙦������F��N3)t�@�U>����2L\y�ڮ�Y��BW�b/%���f�i���D`� U~�u��dB�Z�2s0�ŝ�zx�X�%r&�dCH[(<��ԛ`/ߊ8� +{�?�d����R�{�����K��gY^!�p�i�E׎��Q��|�hI���P3��v+)DW�9�fk*�k����<w�� ��]��d+qy�d��������P��o7��ǡ��2��\�Q֐���Ȓ�a�(�	;%�0�MNr=��RdGNGd�Qӎ
(�=���j�O�T&��͞���
{���G_/|ݥ�
ˆ�X�`�r�Y�����6B�5����=R���C���@�a�`C"݆kz
2����q��l�Ng�$Qcj�[EUb?3x7ϒ��7��F�	�}rZi!7 2*�x�X�յL���Ҁ[���z�!�Zoε:j�^�����	߸e��I�:�ҹ`P�(�m�k#���@x�ɥ��Bj��i�\bɍb8�0D=f��>-����_�,��On��dhk���X�2��t�`#�P�5��֦�Q���u_7`۠B�-��1���zRv��!��2�{٪�kdG8�~�QNG���cyV�Q�Uwe��0���/+3]�4a���7<F���TK�ؐ�X$>#V
IGA@����[~�H����!xY)��@����-D?-���6�mǔ�c�i>z&;��cE��"���@+$Q�ݟ)P�I�!-pf��&;}�1��=����j�qJb�V��J�Kɩ߸��G#�yS�����b�lG�͹�cX�YkO&A[6o*����
Ԅӑ���ܔ"���^��;���ҷ�ea���J%u�q��'�e�9p��\�*O�r;R;RF|�\�����B�W�}�y�.ʆ$C܅�rN�k�X6��:g��hE�J���?�����1�r�u^�������1�ۑ�'La�X���3 ���@�����1��1������[Rś50�~p_J	o�i�3L4C+��oR���-0�ǜp�P��B��E�9����ق���<�:�3�ZcV��.Ұ6��R�\�n�'E��[�0��-�S`vy5�T�ZTK�n�*��e\���/�ҋVs�J٩8�L$���L�{T�=%�oR��63�ԃ��z���@bE�wG�Mg��/�M�ZZ3t�����%  v�-&$���y��U�^�Q2Vs����ZJ� �x+�ǈ�`���KZRT"��!0���=ܶ������j}Ǹ�r�{B�}P���K��u)ϗ������i�n&�L�6��,�����3xW�}�9Ǩ�/�72�̇��=G?�v�|t�E�;Nia��$����{��q"��eFt����7SK_�# �v����/�xo\l�w-.SA��w3I�����)��"M�%xk÷%�s�g�ʊ�m��\��Z� ��-s�x�!u �gYG��T����o�SE��%�0��4��(��m��epW������#�����5#��i`�
�%�s|,�<ŪF��f������#¼�P1�O>a�(�) <,޲
T�	ht�����֢g���	�����C�$>ߵ�+6�8O��R�1�����4G���
?h����H�醺9U�9+n><n�Y}��xF��s���ޘ"�k/�����e:r������إ�a��	���۹���7.n5���PܰGdW� Ӡ)g&������&��r�E�H��fż�k��Ǟ�V�iH�0�P�al���C��5a m;��c�4.��g s{ݵ�ɣXR�sr_���3s>��4� �l	6�^x�I)���KP [4�_���,-�T�k�t��5����4�~I����CY�H�RAW���?�q{sq���#��B I�I�6�;]����C!�p^�����=:~?Ѫ�k���_6^��)3�E�͹$�!e�A$.㸃u	.yw���������D��8�
d�kԴ���v�
�':���X�O1���wq|�D�C���{I��vJ��A��%Rȑ~�ܼ!�4|����ר����P.�E��GjB���'���S_����+���U�H��f>��n�l,�Wp.���0������p���ȜM���:�̔7�`�*Ŵ&��z�A]�4D��0I^�.�y��<��x|��G�*�e��2���OK-�4r��=[�/�zhp��d�h�-\l�l^M��8�T�"���,~�i�z�lw���I���kZ�g���5����|�y۪���2B�B��@� �c+˚p{Jo��T7?��ی�꺱�e��w0��6\(�E�n�F��{�d���S��L��鑠ر���� �}��kP󗳏y��������z��'	G�VUs��tH_���f;F��2��E���n��ݎ��Y�o�*���nͧ�	��D��p���d�)pDd�-�S��M��(��1��� �̠�=cR�Yw���o"m��9X���:'����A		���C���#A"�8\B2b3�!`��M��j�c��(*>�S� l��k��5Y�%�k���aR�{��h	σ�?%��r��XG[�0jz�#��cme�>c��m��:Te"��Ǚ �ɚ����e"�6�.�� ��N{�)�,��I=���w�c���3l܉�:-I���F���ԅ��Z��4��R9��q�>:���4�"Yv`�Z'�$���*tƖVt�G^��{��N�r2xc��өu~� �!J�E��%��G�gXw�#��򎏛c3��,(�L�*Í��;>� p�'
�u`��zY�Qd��"v�㣄e��K�k� �.G���4A��+TO��-]�!���2�)��D��۶,q�VN:e� Ӑ���WRJW=���|~���O�vƶ��T�!��U�>����[���4^	n�-'.`�
c��s��;�q�.�5VVɦd���2_����ԡ6��ûu|I6(��� _�\(���G���9�b���2)"7��h	ǬQ��>s���3s���w�喰2e��&�����-w(����iW�h�no$���Hg��o��5<O���	^0�������訄���O����"�:��2wK�jY[��}ݭLB� [�@���.�#�G��>��o2k�{�W��d��KBq�<#6�f�F�\�����>�&�5�盌�L${<&��Y@
Dm��|{��98���5�y��a��
AG�&���XܸE-�S���:&�j��j�$��W`M�ȼ@�
��M���:��`��v��:�h���<l
`�}���I��D9�1���0Ǉ*N3#�Q�|���/Ŭ��҇>��h��+�Q�,t�SV�����%s����Jq��b��XT~E*ϼ�+���v��@[��;�A��t����䰨��U��ͬ�[�;tfm��jgm^4�Ud� ���"&���D�&��z�t�$Sק�N�G�v������+�h/:��J'��0�BKHh��q�ҌR�7k�.qΞF�j"�P��Cs
��~��T���l�y�j.lxڂl���c&s(@�߻������J��M�<���FΪ��2��"�H�U���J��R�F�V8hͯ�
(	��k���T�̽�ݴ�L��?�va���zn~���bn�uz{b0cV󌎐��L��nDC���~��Ě]��l-�~�����!I`�}8����=+���S�{)�?�yW#8�Ӎ �� ��i�����I��m����ϸ��"�C-����V��|�^?�u�@!��h�JG(2Αם�i<�~�P3핀{v�_�³P�$p��L�a�����}"٣�+���
��^m�t��60���G��j �OX�3>�?T��qv"���Tk9�9�iɷ�ǌmY��[��1;0�R�YGA;V\i)�C��+M�wr��"\���w
�sT��mP��._v�h��&�K���d#��Ӥ^�B���4�[%͊R�.���`�N�U�Ov	����.\�d])-	��e!m�g�&u׍	��i��a��`��b?=`�FJ�����b� @�B�^�:�`cg�
�f#�SS[�a&���
R�Ĩ��4��~�@t���6h��0�K�Cdh9�t�~z�S-�	%��%��E@�Ì/�����C{`E��4��r�u�oP�8$��j)(��n{%�M���(��{�b�$�oaw��-��,�=f�g����v�Ջ���D�~�W���r�?f�ٝ-��ה��!�'����ɨ'��tmG�	ச�x���Q�/���:�0{�HR�Ty��SuK�K��k�8
{+����L��)m�, ZGH��s�е� �S���x�C���*��иn�a�M�g���ƣ(���"����{�ڙ*]�+q��r�=/E`���r{�~9��uΜ��*7"E�LW)��%���Dў7"1�'9y)��jP��[���e�w�ڌQ]��|"W�1l[�ɾ��L]��e{���l�P�#a�v/\���,e�I���$��я ��?q
Y��uZ���d��R�B���Z���o�)W?���~2Z ��!&G�J�|+����%#z6TD�EI�F�x-�Z+Ǳ�H~	QMz�u.�<��[���fý�ف�C��d�Ԍx��)㓬J��:�U ��i`J���Xx��	XL��\���vE3>	�N��Q-P��9�e�wglD��z��B�N=Pi��ײ��y��RU]%X7痫�73R]zN2�-���"\�p2@?��/� ��-�B�k��Pʕǲ�-\s)��;"X�l�E�sF�[>�l�\�5)��z��?l<���+[x)�i����|4������gXNU@��]>j�y�����c6��D�X[�#�-:-�#2��T��V���;��J���%E[J\گ�49d���^�ک���4\����f1wCyz�^Y��k5@"s1��5�/����@`̴4$|N���$Á��<c��ﮃ:p���"�d�	n�B���a�'B�i1�=Wv��t�2dQ9�s�y��2�Xl^a�:�J_�!Tk^��^9��t�X�o���(�]���-7�۽g���Ţ�#�%7f�-�G-�!������+Qp�&L0���؍�?�D���֧�kg!x+���vp���~X<��I����gu)0匏�4W�����$Ԥ4M��r�۠���Y��/��c�v�2Y��ՓB-�~`6)�X���@�6T�!�mȲ���(z-�^>�3�'���"�@��m�-9\V�%c�<k���z�K�U���ܐ)���q9Λ��[֗��vQ4zE�X��@���Rq�ɍ�.ܬ	��?��+`�W�wB6�"�y��������� ��rM��Y ��T�$�v�O�/[S�.�ǆ�����yX�ܪ.�L1�`p�$'�;	��3J<�@�����\�$�leԓJ�����@��	߲��Pv2�1�AY���a3~2}��uL���֑O��ޖ��?{��*#m [��.��̅r��Q�bqWQZ����,$�R�!-��b�P���a� �#��X�٥�4��z=�z?
�h&�}st\+�B�ZȢU�o��6r�"�'&8��ơ�sK��h��	 ���/����ݨ�q�¼/ŽT5_p�|?�P�"\/!`b/�����0;S�=�c�����{�
��r�"�B�?A�]*��s׼�W�%�i���;��(�&�?� ��C 2:sbヌ��2L�m7�z�QC�A�au"�+S@w�;�2�w/,}�P��h���ȩ����k�-N���j�@���">!P�Ry�*�Ґ�������9n;��-�b���U�Gxm�X���3li��I���4 ;���I�b�u��|�L"���^n�N���v.�"e�b���_�E��ϑ��@��Ũ��pPUFC?�@�^�XK;h3�6��MS�b[��fdi��>ڥ7�o)ٻ)66����q��<u���{F�Կ�p`o'�B/���؟\h�%�"R��VD��8L�#nc�Ӗ?��2���a)tV�M	�<F�L���9Х�z/J�`e�>���5�o����r��+����ŽX�=O���"5�F�)�e�!����n=����@4��e0	���-���!Fd,[xٍ>�mLq@<�O�m�֏���Z���&-I8J� K�
���;70�gh�&��lj���S��Q�敵�zاK�*Y(,z�Tu->��=$z��^c��Z�8Jgu)�p��X �ջ�$�ۅY�AX�A�,5�<�E�Y��?�>��JM��ku?��5��� �gmPO�
�#]��:[���=<���
IL��>	��|�[�T��뇀ːwv�:>ͽӦ�ě�@����w�l��3L��SM�l����o׀U;���U�n.��P��%��wɑ�����Ai�_(�߅�G��_�u�J���x�9M��}R�[k�i�(
M.T�ٝ��q �~�^����;��飩P�ViY#U�l�C�޳�Ց2�
�r��������22�v�JQ�pKj�Q.��BJ��C��}f�����(9�%~��?��q�h�"K�	�����YY(�O8}��^���`4.�q�qh��%��l�(f8R��\�f��mש����Ւ����^�\��·Y�0p��E�� ?�;���=�'_���?*$Vǥ??2��zVLG�V�ݱ\K���y�a�?���&cF��$xr�	�����	��	�k(�L2J5BBgh��[X�.|���G���>�8nYe���ح���3�Ee�bO�0��� {>��U�l��L����[Ű6�T�<Ġ�W��  ���=��aP'����Z�u�a��UI�~0i��2EQ�M����`���.J�0�#]N�չ�J�e�I�+᭽�-�HpFQ]���'OM���T��2I��e5��B(�'"��@x�B$1L5L��ÒUfƛ]���ǷA���9�%��<x����	�� 0���b?Z'�M~|�x�Ikz�Yh6>'��4+ߜ�,��zu-ȰQ�.�OX��'��+��,��d=Ԓ;��cr?-v�Ͼ���I�]��B���Ok^_|�z)������C{,~u����s�
��3<����:U���'$�g��D�*�]-��7�	\�`�����Q�@Y�(��.Ax)r9� $��؂b���2�!���*�D��,�E��o�/����� .����m���n�^��W!$S���ψ)3��ɪg5�&sFb+x.�b���~�Q�pU�B̼R万�Ka��V� �P!�$���>k�E ����r&���T��_�G;r��u:.�M��l�kp9�"�H��Q�N\u������_�#�MȐb���?|���ZVO湍3�ޅ��G��b�����8"�c���#���FTԅ�Wӌ(�{�4A�V���Hb�rr��+\T�Õ�xE��% <��
�rxMC!�r��:ֺ��wtK�DVFk�sp��j��]8Gta�;�-���"ş�Fv�O�������`F
����#V	�Z�R{��Jt�yL����v�Y��HO�Hב�~���bv���BN�وm;$,\�!��h:=`Z����g'���������6���τ�.�P68���|mѤrfEz�-!��M�5�מ{�t��{����
������mݳ�{�N�A�UH`����z���0N9�*��"��'��<Qڔ h�Mg<u�Sj�����7�.��<�Ҧ�w5)��5�;�(fZ˿8�S(�PN9�`UH����։��ˤNp��8x0�	�ZObj�?�g�S��.�Il/*9�u����)�+�@��-`{(�W�t��ȹ�e\�Kgb�Za�����fv%<_��KLj�]/E]���W�J�:���~1����)��2��V0{��}N�^�?�]d�IK����7H��?B�H19�WC}ߑ��MN%D����)צD�w}��=��1�Zl�<FN����4_|]�M띘�p�����_tfӫ�Ab��B��]%X��-�oij�#Nu!-�#ў�O�� -�Dhȫտ�V ��?��==�u?m�Q��;�m�B���P��g6�[�Li�4[��u0�rop�G�����w��,9�'���Xn�z���j���L�����w=��=�A�y����Ə�@=Н�tH��;�)e�B10��\��Y���\;�r������3�N�ɄO��\r?�$6�l��h�tX��K�tu�����b��J,f�Xs�R�\�h" �"���L��񐖷@� '��jDxg#���S��#�a�4p
f�V����X��ǠG�5of-�?E���M�����[L��JqiPY T�֑�#�^)���apg
=J��Z�|�����&���3T�EE�"�s���4�H:����;ra�t��%�2�@�4� �R9Z�"�3��e���������,�YZ��I�
|�Y���5�4f�b%��s������`�e�႒{ǚ[Ym;CbW��"Y({���К�M����#b5����0	fff'�fxwE�B��l.�#��b�tά��EGRB�O���D,Ml&ࡇ���_�'��S�^*�JPg��%BN�NZ���k�/)9b����cY�؊_m�۵}�/�6�㇫��?m3in��K`�u�<\ɒ��VNDK�# }~�rL8����5iZ��2����1vt(M6�ajn��\�PpY@>-��nZ����)	U�ӻ���$�Kv{�r����mt�7i}��#��]7�Ϸ��@B�Rف�[&E���lλ3�w ��څl�d���]62Qx�g8(O]�
�u��8��~K4Ogk>Q��&
�=�`��8E�bG+ٝ������&��.Rf`|f�F�.��V`�J�G
6 W1�wu)�~Ij
�U��r5�S�X�6l���і���챏��п�K�Xɑ�=����j��	�Է�o4��5�d#�`$��ϸr&����;mNwņ���۫3��4�a�� �i{X�֟����)����$I�e�퇨��e�Jh�h�.gEG������j:٩�����i_Vp����_�S$�o��kW�PcB��k�˰+��3�0��j?�����_"y����_��tX3�5���_�%��L/�M}o� ^\�|�xP�VDo����W���J�D4K&v�r��׋�K�樍<��i	CG�2��R���jX�"K�E)G��O�C���q�ԭ!�À�q�F�Qm�`/U Q�:fu�&١��%�|
�AyL�ż|`���cm�����#K���}�����R�u��FH2)��S����U\����Pwl��\���z������H ���P����:D�j���� �|~!��a���]-A��3�LFG`��,yQ���,g����6h�	�W_�<y�G2��MQ>L~=šp��KT��.�uo��25����K�4��#�f����V3�^]��N*%À�ގ���粢=穘�u�}4�?�L?4�o����M��_���%|˩��Z\s�Q�]����(eȬ�1��*�S �9s,V_i������U} >Gf�x�����#1���f
8%*�ӗ�B�,Z�L5p�7�Rrn�&����tk�N���Eks[�A��q�j���߫z0t&��$V$���G#��yݚW�Nܓ��^��OڻE�L$�����������(�O��I$aD2J��\s��p4=�I�[���4�3�U�����/�һ;>+��.Z���3pm4"�|�,@-[����~ ��EM֦�%2��Ա����av���Y�p�̥�~:<�u�6M���z���d��� r����e��3]I�)�U�j30�H^�] ,Ȥ�C��M��uϡ\ �!���5h<�hwJ�߁M	�W�Q[�;��l�Ѱ0gYx�W$7�Wy�p紾���8�B	��Q�X�� }�Pqr��b"��N�Ӥ�O�N3^��1��,_�<s��c��d���v��s �D6I����o�y#�+���	�T(�����P}$r��P�zm�ˁ1�0Y�%H��������	#�Q=%��̥rs�2��\���K��W���h�T�
�8�!�5��
�m��7�F�m�5�3���	�<�b�D�cN����:���������S'��Xh��9Qnի t|�m���^r^2 ���-�/'�rk������/�0��������㵟��=�P�98�S')��|3$\ "-F"���Q�$�S~���uzaT2<�l�V|V��f0<�?�>tv!&��W�/_���(e�]�C��0��=P"��+�G� O7D��w��Fߑ[�5�o��5F�)����E���*��6{�nS���L� �����]�&��>�{qr� Ne�n۞� M�c�}s;ڢ�=�sN)qR�� ����@bh���[�;8h`�:L>xd�P�w/6ZF���)?�C�+1���4mΖ����;���C�CRZ�C7`Г��1�!NQ�fu~�P�}�����l����%�16����x�)�7���,��P�KF9R�u���3�k?�����7�Ź8������B�5dx��|N�I�kt��uO/���V� ��}݃��g�>07�(0k��RNgG�+�����_y���J=pi\�]S�T�
�"��܍���X'�S��3t�E�o��_�;χN�Dl��H��xL!��(���IO���"���o�7Pp�B :Ƈs#x�xB ܕ�2u�$���mb?�}}�"#Nq�:�K�>��B�d�ׁ�d0�I��;.o�0G��w���>�Ō᳟x:���n�*�����Γr� 5�|���6�{dx�8��
0�{*���������H�:�,� @c<<<��ɰ��)J�hM>Դ������9��`���5`*��j���r�PǼ=�,g�G~�ݶs�L(��SoP��"���dlHyq#��:�� �Jy|�k��t�U7�Y�\{�Ҳ����C�t��6#�7tf�ꐥ�ͼ;�Va*��E ����F��g��H�I/;=2cC���J-K�/��e�*tS���U��0Kl�2�h�[,��B���w�,I�ܥŻ;ͷbƵ�F=�Z���o���ƪ^y{�c{.%j�]@!�P�3�����}��(3Dv���B�5�(�=�T�d��g��@�[�޿R��,A��d��h1�B5M�V�R�jj��i����}g$۳>l�-%�"�h�����?\���jS^pz.[a��O�%t[�{{mMP�-�{��,(s��� :�l�	y�����Je���Y�d�2�u�ՠ�o F�~]�l3Cc��r
]ô��K���9���&3[�!�C�-��G�Ҙ�
i6���'�N�X���F��	���GPG�ǴCo6�"y.s�TV�YP�8_K��c���n�>�#���=7�J��Y�����c�H�5%ͱ4�n�hQ1��LV�g�e
��Ry �yӁ����KeC[$ƚ�o�zľ�5/ �|��w9|<V��?z�#Б�L����'!��!g�5w�u����?�g��M�����2-����gǕE(f����f�>�e����CpM1?��<�n+Q�>^
��@<��BS,�{H�M�S��	J��*-�����:��꘾����d��h�'�J�礽۩�����T��Ŵ?$RN ٢��Z��e���{�*��1<H�\��+.D�"v�^�����{B�r~�f<)�!�Х��}�*��[}e�8�����q���y6����~�)/������U����!���;��nM��V�@�W�y�=�F�NJ�(w�Jۉ+�-��n4��kJB+��FW������&���i�B1'Qe���K�s���)Lgg�I|��o�Ѓ�4]%D_��6,�o�ggP��]s���S�"�f><����٪���Qh(��]��@�I!�Р���<UZ�vc�wR�oЏJ�o����r�B|h�i�DW܂���V͔W��ɝ��v�=8�`��S�J���<��j�LHϕ?n���u?��	��K������b6�V���t1Ei������BA�ܓ��y',R�	LvG�}t����$�.o�����`/�.ߍwIzgT���Q6	4��x&�	n���{ E�����@jrT��4ك�����j+6_:kۘ� ��(�t5��P4'�����+��z^�kt�T�3�o��f>Jή8K��a�.Z3>ĽA��zy%rh�M��䃒��Y#�Z:�1g}65�´��e$ǉ�||��P���dG��7D����N0`@C�5�obe?���P���c[�[y�M�����B���"&R�ƌ5���M��t��=�jRW?D�h����&ǒ�� �HhqL����RL�B���"�{:����@�-�N7C��+�}�����md�i�oD���$�.}G~���HIhHRݤ�}_`�:R�D�(OY4�u�������5��]�o�����O f�ti������)���0ޗ���k`��+=A��^p��(B�?pTA��RaB�4��#ˣZ-,�mpr�A�� ��Kf�4��f��/�}��D@WB5B�?��.�3�ϖ��oW���I �V�7�Ĳ��:��D��?��x����T���˘��Jܟ{����ʂ� �O�(t7�0ߣ���-�j�-0�R~�B6p����\���
��o��{��%9,y���)4SJ#��Ї�w$8�	
��ʊv���"I���e�BR0i���j����c�T.�L��lYВnn]�^2kt��S�h���3�ڐ���V_[��
�b���������ua>�u����C!���J���EP�$7�8�����;VV7l/���t��T��1��<_�F�x�����1{c[o6��X�(�� ��z�rԑ��8���Ő`m`żm}�T�}��Y�qz�9�P{�V�զ�NO[��M}5�]̌L�Em�^�0���@�3,C��ê����N,���=Ku���V�8�l�F�Nlq`H>�:v��#<�
��t��Xi��2��<�>C�IN��$Zj2db<����%��;7���;��Gv^ Bj+6ζ�x�u^�,���BMP�� e��o�v���#
�����.�S�P#O\��� �o��>�j}{kC��qU�!i�p��ND�v��#>���h��|��o.x�P\��\�V
MY��X/~�Vz�R��^�ы��HH����/b���΋�����ȈpA�p�hr����扙��I��,�+����u�&h��jg1��vV�3�������q�o�3�������# �`�ԭ(����*����ˁ{C��W��	�C�|]��x[L��Ba��ӛ��ɊBw�,�V�1u�wH���a���M����ԟތ&�'���"�(JNѧʅ�)zt~���MXI.��ɔgDF����n+��?���a�~:��8���#�_8Իl���V��6-�%Q��w�m�#�f�Uv\[�MX>��>��%9�þ��1FB�����{+� �A�NBC'���*|��"p�P`Yr�*hUd%��V��K���� $n՞�TgUu���H�&@V���Y��<I�oI�kH���4(*��rS�qN�v��vM�]��:yk�Y�ϩ� �����B5�8�2ĵNh�M~��"��Ͷ&�h���r?H��+�P�G]�%�N�#]��W�@�^y-��e�k�CS�����^2��d��@��\¥\���jgE�.i��;�f5a�K�*Ǉ/�~�Ʉ<y�O0,x�ןRaR��:�m�ѝ��?�d��T}"�(�@�u*��H�E|(�NVt�-��x�U���%���|ïd���X�-6�tۄ���Q�!YRb�,��JSm�#욖3�
I	�X�&�z/fD��޷�%�o��Ї�ۜ:��ث�C·�@{�?�!�ez�S>ˊhH�<��I3,zj�c��3���<^`٨|Y4���p�D9Pv�޷�ԉ��h0?���v�7��rl;̜]��!����i�>�8U��iQ�.b�H�?���b�1Y�	Q��e��9W6�#����󉲛�Mx� ���0�;�wF$��������0��g?u�H�֚�Tz��.[�]Ky(Vѣ�p�w���H�"V�g~��Xʋ�R��Ey��~]@ß���WӰ3p�潶0��X!z�����G���歀U��|����l%��Z qk ��ͦ���`���[fM֙�,jG2F�y���!��q�Bz�g2���I��X,=�?O~�$f��\2���b���;�=Y���L$�U3�
�욺;�J�q���	��a6ح�`���-�;�X��U���Ayט�l�G�?d7��%�FV�����U��균"��"����޹����[CL\�����p>|Fe�P�]����[�4^�O늧�3k��'�d�sD���*�巍�ћ�v���PՇec�&�lk�޽D��b�4��;-]4��t�1���5�زx�k��Vwu�X�m>�'�E`9��G�6� ��&�dE9��̈��o�D����0�b��O��4�"��a+'y�9�,|)"������FA*�F}�t��E	�v.����#�Y�0Sd�l� �����ft��=�Z�:�F�� $d�`��?� 	�H���8�8~���/U����t�B��jaP:���fE$�����DU�Ew�:�������z��B��4��O�j����{��wx����}}*1a���q;m~�Jg��`�r���ǹl(�řW~!_��
������ ��V���Ê=�*h>�_پ�\�S�k�0�M�{儖tJ�f�(-��,r����)��N(���K慘����-P�s����~��K�#��*��gq��~,P�6]AQV5Leˇ8\����9���%k 2��'v4?~���g����TY/I�{��f�ʣJI��)"�X�=z��/�6�bM���f��V�7�jD�,Q�D��
�wN2d7��|RTF�|��<4�S���G#�:�5�q� �O�H qu��5 ��d�x�Q�z��	����nuu8�N0w5�����n��<�oϯ��THr-���@�����Č�^���Jp`2Wg�w�&��H(�}��o>(r-Tj��xh)�#y)��
��Rڵ=KQ���!S��b�H;����|��� �"N�swW�)��z|��1y���+	)�䀗]��wZ?:�b�R~FD�5ٚJݦ��֦�þ����Dy���9�iHx~���:�3m�5��Y>eZh�nĀP��������Ř��~�3/�`�{;�w�$������L��9�Y]�l�0P�Qj��ޡ���q���\����g�%�&�����tH�LN1-���%W��4���vF5��^w�+4��	ڞ%B�X�~�����~5�D�6� �6��Z=�93�X{`m�쬄Q$�\#L%%��[
H�ǗM�ڜ���v |�/�A��g�`�j��r��H�y���d���v���a���`ŀ����7�%lM��)v�c?����<�=;���Ύ�+MuR��>������~*s����3�ju���L�<Ɯ�,g��q8$���cd�ս0���g�sI�����
JNWD����檒
Z��as�@?�;���_�)�S�FT���z��ħл�9x�i�Te�Bst�������t��b�JR|d�6?���sGs�'�<	sZ�C�/�} 㪽1~�|����	i�V
�ėxt5Ƶf��+���X�q  و��+~��?�>3��qi���KV
������K�}�?���ӭ1�7��iu���
L���R��[�g��w��M�tYt>�B��S���%�{:�y���e�_�VPS
mty��*�MM�� Jro�\�+T�">4�)I�p%CQ�(���1��
����	��}�[G!ՑUگ{%}��X�N&^��,ݘT*���qOao9*],w-������\����X�v��c`��*�uD���BGcKU��=(n+R(����������0�r�Q*��#O4��u��4n��q��t2��͘c�u�KNĥ��Ϫ,(�#�Q�LU�[u�v��`/3�$8�=P2��(�ԮM������sб���PV14��W�F����#}�Y�A�WK/h	��M�G��$wo�lJ'FU]����t6ѿ�ݓ�c%m&/4K����j\����v+xM�x������hњ���@�㯬6�
����KJٚv�����}ñ�S������*�v��13ǖm���QB��.�=W	;����/ ����������pC<�ћJ�7�d4d��z�P9$��(WbE�H��
������0���c�c���}�:=�N;����l\��b�~�3Kg��ߪ8�����~�a0+�!i	9rӚ��M�`�2�xB_�1�_):<��Ȗ��idg��>�Ǖ��j�I>R����Ɏ��9��)ru:6�R��jLu���Q	p���,L��ڪh���S?� ����!|4�E>���M�D �-0�
�1��c�Z�����p�M����E��]���˺\��-���֙YW(���(��ݜ)�W�OŪYq��G�ͭ9|9�f^�=4��X�͛�k�b���%m3^,�$=.��6�H.�Km���u貪�fu��C��P-Q�h���5M�H�jO� ����d9�z���Zp�ry��%�>�E�;�|V W��
��-e��+����6�FǄ< �����d@Z�t��7�y"[���oB�Y�J��̳E:H$�u��~���Kl��u�S��ӐZ��,�sr� ��]��$�C�n�2 ���ad�?H�ѥ�h!s,9.���YE��s��mv�ΐ
��T�\&8�)�(�m͎���R�W���D}r��2�N���1qk�P����bG!�1��&������ȤN~]��a6�]P�d&��4����2���60[A)/Ob%rV$�!�ag�y��u��''�#8��X�ꋀ�?��i�/w�A|ǵ����,�x�f�s�?蠢�O�jd����M�<�&;��o��׏�_��TIB�qi,E�^x�<�a:Μ�@�0`5�l0����C��
2.� ����Mk���*>1����ce"�ߺ����+e��VhϮ&���Ro�����~���R$(��`�������W��I&Q�t@����W?�0�Z��a��C7�b���+�.\;��4x��d�I҆̿ۺ�T����t[�d�q��gX����P��������0�v��ݍ��4�U�3��˳��9i3k�gJ?���Ѵ���PV�ŚUAʀ�V����9/7�qX.���S��'3�k]����(�/{��8�zs����1���67c��u�L���CGFu:��n�Q�������2�3�n6��z���1"77��G�S����o!%X���'K��)�{E���A|���r����K��1�� QV�����Y������;�|�׮�����9��Ou�Tз>�y���3{:��`�W$z�S7�š`�
{?��w�Ō0��&�����A]��8"W]-*�|���HK�I�[w����[���*�ե�7v�*�=���B)qt��s�l�8Y��WU_60��&_�,��n=$�oWg��goO����횾��	C6�эr��'��^��߱������`�����y1b㢤Z���=�T�f��)���8	�����׋@����&�VwoИ"-�.��{5h�/;�f��8wc���2]-����O�}��j��F�Ru6l�@I�'���~�X�K� ��[�q��mkI�ѷ;�Qk��f�Dy՞�[���}���=���>�qZ�I×0Vߎ����Aa۾�X[.��Ե�{��Z9k꽼"��-��U�<��7J���7=�Ebr�*�z�����Wn���~` �|Y��ԇ�="�!���6��r���a<蘹#�3|��t6)6�U0���H���S]��FCs6_��3�Y�D��(�ݖe���o�3+�P�;ʨ�]�\��L��3̧:�7٠[�׽�K��(cJ����e�=�B�Kɨ���lb��ff���n�0��J5_����9�
6F�~���i!��s�˄]�7�k�/3a���)��#���=�L�;<����u%d�6­����xx�P���&S�
��ޥgf�m�������ڝ+v���R�6���~sι���a�^��;�%m7a�uS�$\����������79��DY�$�h��}�˰p��4��f�m}�EE�ƺ�;4W����lkƯ�mG9��b7Cu/m�t����u�/N�c���=�Rv�����&�"u����o��|��ߝ�x6B[@����y���u��7FuJ��1 ���.2��гc�o/H��w�!��l��R>o��A�{��<�ω@���X�f���������8�iK���X��\*p]L4d~#+`r`:�	����LI��p��H
�i�>�c��u8m(P&��C����+|�v�I�F�B}���<@G�\����
܈���׍0�Uh��H�(��Yr�܂^T�gqW/7����Igd�mV�Q�P{ùɝ�r�	-'��\�f�&�5k,�^q/)i�){=i��S�K�ڠ�$i�W%�-VX��t$Y1��X������$���3�!�h�'�J%?��]X��V��r0U������p9T�~�G��0?�� �:z�M���uA8��c�^�����1C1x]���ϨQ��Z��~�����}�n�:����	)�V{X����K$*����ؽ��p
�U��{�	y_x�H��qU�.��*g�����qe�?���@�D�	�|N�ճ�=��>A6�KU��l�wusP���nP:�巕� ��J&פz:�U�Se=6D��.�����Hߺ�zɄ�u�Ug���Ґ<8���w��T�/dNC��W��͔E��/�{�5�ek��0(؜�'٤���$߀s��x�Bu-�� ���F�x�S��g?|�ȁ-�a*畽g�����mP�\�N�$n/�,�#3�3�7E�%L�p�����m�7�����jL��Ĵ�Z�%'��N���>c��҆����I�k+# H@_"��t��jo��Vѡ ��W��ߖu�N"�&��&�k��$�}�Ւ��v���F�(b���,��t��|8�D�6�nn V;�NQ��n�z���\���L����9!�Gw��<���r�b0��]!�G�4HU6.j��~F��C;ڊE`\���w[�MU��zЊ�slD Q��.���,��^�SmЫuM�4�f�p�?�	o��cs[��[ã�V���u]+uQ���c� H���׬�2n*�qSD/",~���ǘM����o�{��� a"Z �걨�'�M0��{̴��[4	V
R�����$gy���L��_�ӧ%�$��]��P~�u���'�mn��R��-���[�aݖ#��K��U�7Ij��+~�oq���uo:��J,�����E������x� [gz�ǭFa��I����d�:�(��9�A�\�~&/�c��:�5@I}#I/G[Z��޳��^SY+��`WqW��Hځq:�%��qx�� ���T�����2L��%a
�R�&0��Z�}��Oon���3�&��� ��d��齿�5�' T:�)N�E'b�=���u�[Qʾc�1RPG�E�zE��>��c���!
�2����Z��ϝ��CQS�r�+�w��Гv	�+������&Yڝ;b��r`���f�ZUw?�2������]��\ӳV��������ɪ�!��O�Vϳ�0�,�Q�{:t�ũ|��'˿�]�l���Ɠ&̷>.�s�(�����t"��7��ե���(��c��F�1�G�?m��Jlv���d�{�hG'�X3Rtk��]�S>�N}W���D���;_}K�>f�\��
���cZ�0:���S��@ߒ�Zg���g�lm�U�o�d� �� R�C4��c2�%���ov'�uC~��e^�L��ҁ��s���H�+�-G�r]#� ce�C��+ӈ���N �y,�_��S	�� o]�׏��P�f���c���Wd4_n�����ʦ6"��ϐeyb��MVw� ���AN��幢�Q��<�*[+�]��R#�Y��'[0�����eڜ��Guͱ���F,Q�em�cwե^��"�L�GCO�-Ӊ-�[D�Y�K.��V�x�dc=�������+��ҵ׀�l�`���}^" �?
�`������1Շd:s!�:(�뎼J�L�[^�{0-�Q q�k\���~E�fU��%��e�a}���9HB	ר|�T��X�������H��@$�V����d^�R����	�4��D6�:��n��CfZCsW�d[|o�.P��K�Bx�[l2�s�&���`�m��)����S�{���4/(�}*�`�b��<���Rm��Z�~ �]���o��ţ��S���G��V�*z{��Y�w%�a�<��0�b����&����$?>� �ޢ�~�J�2��<���b���)D�g|�4-K�C	���O)r}��t.P��Ѯee�c�h�t�;�E�ߋ�C��pz��6� "v:�����L5y9z�ޑ�9�I�J7[�i��%$7�j�g�M���y��{���Q4��Zhh=���L�]�r |�X�0�&<�JMP-s%�/\��Qh~{�P/�x��b;� z��J�{.��%������������H{N����D��p[�5`��xRQ)�����-��}��'!l�@����7r��.#���<�N�r5NT�MU��G��i,(���yv��߰�K{o���t�}r�(��H���B�i�J��$&�i�� B=ih�v�7t("�EsK}�C�g�OD_{)$QJВ��)qV���+�X�5T�;���#=_�U�4�%|���?��P����n}m
8퉟b~����4t��m[[�r9�$_��2�2�+�D҃|�b�F:�� I_=�G��7�ohL�&�L��:��	�d��h��zMӺ�}��I6�1K�\�1�Ւ��-Z|f�`w�M��8d
�p��eydd�BtY7QPD�*ݨA��Ӂ�
g*{��G�D%;�[A�E���3,6��$ �Z�&�B�	-7�����MяS��R��ә�}��Y��P�z7�47���h�Ѐ,i��T��U�o�#��R��Q	f�nH~7�L�e8^J��b�(�P��,��wRr��v���Y|FܫYȨրU�G����˒!�f�Z'���U K��W�Q�P�k���c��	I\�J�������ż��eh��%�$�<R�T�~�+vUT��_��3$�1�wE��Ӎ������&U�qa��N�5�ٹ��-�׆oB9�T ��-��Hʩ�z��۹"Ѡ�]���)����`>q�&>R%<A�����IWZA���ឆe~>��_݇3<�����m����혉���CK晊�z�/<3�1��#ڛS�:�O����I��L�Ï�BOj�'+��n�Q�h��|��#�n�uL�G"���&�����Mƅ��k;�n�-���z}fu����N�aL���U��`t�#))��O���jr��0�3 >��ƀ�a�b��@�,���zʚ�S��pT��rݡ�2�~r9�Ύ���"��Jz$�`��nDB�� GB��I���B7K�%P,o�&�i�����z2�=	Pa�ٖ�9_��\�ct����/����fL-U I��G����*�\��v��R  ��D�"9���$��4CI�D,_��0�#��#�s�v���e*˰�\�]��3AW���E�e�jb�!�.QRq�������XS����N�āo��rl�� %3��c"�{t�˵��홖lD9M��g��I�K�F#&�CĶ�x�����ؖ�{�`Q��d�� (e�g[Ѷ8���GT�`��"��I���;V
�Q��������lf�1�>�FdJBqz�*�J�&2K"8�F�ny�م�kvt�"����b�7�<�Ē��g�%~�q�ܲ�K�����l�c�1!���l�� �Y凝H��(!�?Qq�6�ؑe����Vl�9Ɔ�J�Yi%^�L)��gA`n-Q �Y&��1w[;����D�Ǔܖ�����n��PՊm��S�|��\ꐟ��yQ�{C������qԎ�BKA��¬'n����.�&!��x�o=��~ 6�}T�&~��~�W揦P*ј��|�-=�<D����j�i�-�� /����:�b�^e1�l#�����f�N(��`�hQt�T�������U��0�QşᣨO�9e��ނwRy`�:�+ �3��`����u�j�����~z0�g	,�H�Xy�<R�5��#�g�p�(-�]P��~O�v6�{=9֖p���cM���_b�q:
�/��"� MS�qs���i�� ��>ogb*E���}w�c��+�T���~-�/�-�2�/D���R�<���x������<RF����X�_�P��%��g�~���j_�K���U	ߗu�T<e;�c�\�OA�dr�%��h2�bkhÒ?�r����yϷ�ph����� 6���DY�|� ��u�<���ڥ�<]
������_|-E#�����%[�_,�$��Tc��L��h7�ˏ:*0Ã}m�ц
������6v-����H���ůM������R���jK@mj;�.[�ݻF��m �w8�fV0w�e�tFt�o� :�w�5����k�a��޹q|J�@�Tc��ֽ�v|=�mh-P�9�-%2���E�����L$L�x���#_y�['K��t��|��	d��	f1�I㢨|����z�[9\�݈)�)G��0 l=uA��aOl��M�aV�-��U���QV��<C �d�R�s�l�@DU�؛�g��Oii�_ggv���6T\t|���X�8� ��=�fM��:������`î,�ψ~D\����{�?Rʆ]~����{���/U�&m�w�7�*�̀�{���M�����N��_�����.K��y����е"����lFfj׮�a���ʁ4	f#���)?�F#4���Ve�����?߸q信SBK;V�McD�J�S���Lr!5�V�Cҧ�rx'�w@v�wPj����cN�6�k�4����WyM��Jd�BǅW1�C^�0���opú�x�DW���~�f�{3u���6�� Yh<��Q�+�wy���P�S�s�/!�/�!K�?�8�8�����F�V匬M���edy)��#]�NT�̗H�L��f ���W}ѻD�%e�]U�C����ceT�|0�׷)�㨲�j��;u[���8M�<-��dFG�6�Y�3CŸJ1a���=!��O2jjD7�B���2��T�s�������Mz��T38.����?$��A�e�sj��k	�BFj���k?)F�-ܴ�ܾؼ�<�4��tB�+�z:�����5w؄��i��a�-�]�����1�93;
�K�W&��ާi��
��0�4��o�v�<N��h4����?��p�N��qyO�?��>�
�+Tfմ^�{���ķ��Bl��y�k�O�OO�<$�� f�j��b��WV{;�F�X�+�mQ�i.���*c$3I�-�a[�F���	���Y��y	+���p�}�!�x[z�D]��Y����c�[w,�t�JD������I��ھ@cX��K$I��@�q4���h�Z��C���*l�c�TB����~p�ބZ *sI��7[j���� �L5͖/��8�q�*�_�㆟}�-n��)%��)�&�@��]]��E�U�G�!�ERA�L��ow�M�(D� �"r���g��y"��I��猋���ك-q��b�I�n�Hi���f0*�d,�a^������>i��Р�Ðt����۞�ʳK�5
>����;��ʊx���n�S�	����'��)��� �|9YdJ��<���Qx(�pd�Dǉ�jꔠ��,��>K����p���2=�C���|����X����*�@�5�B�-�~>�-d(E^P��~~�Xÿf�m��L�BX�֞�O�u�p�=ñ��9����}���@�qD�|�<�F{�@�����h mzh�:�.�L�z?�G��/f3�:-�x:��H��9\)�6��@��N�J��?�����V�@`_�C��O�W�Ю�e��C][��Stm���� ��Q6ɡE1�I�x�Ky�^�2Yp"Wg�*,f��	t�'S�2ٹUq	����$"=�?B8�o�+G��
�.!�zZ���Q�?�y��H�Q:��lӹ_�No8C�F�t�$ 	���\L�qJC7��KN����G���J�BGR����m�Թ�%3���+����!���J�����o~1���Ш��?��&�/]4����8#��n;�0|Xؾp�����G��$�d{����w���ܛ���5�ҥ�+��m�º���v��KŃ��W��C7�r̅��c��EX������*e/�f��UFX��p"Y���3'��T����ä�-σ��#�{��*>l�y��s|��P��&��x5x������(+�Z��>�p�T7���Ә��&ƛ�ynӸ��%B0�O�!K~���q��0mI��o�>46�҂Q*<��@�Ų��}�? ��\y���b�c��G����i����q�}v�WҺs��YŔ2��-�4��G(f���c(,.���H�D�\�z��C�ũqg�"�zWw�N��t��R���-^ �A����ZG��F�'�>=���AiW��e:ս'w�%d:��ED�f����f_�}T���� ���e��?~7��֡�kcwD+I�h �+�a�j�5Y�t���9Û^v,E��C�|t�G���� �T�i5�X3�e&es5�1����CRʌ�`�q��7B��f�9��Y4�Z����.�G ��	�x��%X!��� �'����l|d����vQ�ꦦ@J�?��[}��T����'r��s����~�?c���`�Ȥ˒�S�Ei~��1P+��0�iL��dA9H����鄐k�|*w����ߴ�i]e�	L�5�Gm���o�ں$JY����D��T.���'@hf�kY�vۄ�1�m{��4��L/;wQ�#+Ѕ��zTw�I+�5����փݚ	H�yP��g�#\-c�H���|⦰|��d��I_<�<Ж�k��Wf��@1���!h��;��3�r���:@��\����p?4:*}�Z*�%���O"�%���p���'�y/���2=r!���緵��D�x �K`G�ҙO�[v���{��J}��\[�k#�=��B���ٿ�켣�}c����ړ
��qʩ�(����M`�������3+�p���'����F1"0���l݊�L&��o���˷<��߹:B�˹�8�j����R�4,��xr>P/�ͪ���(k��l%;�9M���=$�i���"�V(w�K�@�2��s������[�ۦ�ϛS�+R|0��S�?bR痕n��\��0�m�wQm�z�h�jU~��Jf���te�[�D���kԅj�y�b4 ��?FcI �zu�UcMC�H��ӭ#Cl?���,�Z7��R0N�dX���[����ʘ_5KY���d4y���VC��0Ѱپz�ǞdN�|h�y�f���l�K���vQ���A�X��$�r.�\�g�#99D�o^-�<C�޵��'p��	��vD-�8MZ迷S �q<�Y���ᴅ:#ut*�GrNll��)� ���IR���
~$o���E�	����~����rK ~y��{�7q�LSr�Q?�.J��j|)ps3M�WZ��f͑��,�8]��L��缓<BP~��#v�Ky$Uv��5���n���Js�qI^�O��1��K���U�+6{'���]ߢ����� m�n��wWnw���v4�My��92ˇ.۹�II̴V����!�"��Z7�[���1�Ж닂҃��[��\�o֙t.�L�\�`��C�g�����J ���ke���9ڌ���WC�g�簊�g�UG 55�GxB�#_0G��$�n4�,Uc��4����X�F�ӑ���$��<��EȤZ�=S����H�*X��KMܧy�9	�\��[��E�����v�T?0�rc�&<%�q8]�M��5���o;�*�H�C��8�̾aJ�T�H��
n�����@�ԣB�@at��w\Q��tՆ���,7���4v�v3��0�x��G:�,��S�|��	O07�{�J���\W���;���M|-Y���ºV�g	�ٙ�Id|U���e]�7u��1w�>|Ӛ1A`w~��I�����F`	V����6�5+�Y�a��k^�^�0']���@i^������W> ���c}S37ūn��!`�������̽7��&��\5���l�w,�V�w���,e�w�ݼ��Ú�.`fw�G ���&����g��NآV��2��*��Jg�9٤C��'���P�%I���k��	��nmߨ�0�tjgd�����k-h��䮚v?Ǔl*+�E�S0SL�J�^�_�� �D3;(S/��K4�m�%�	���B#�D�\C-� �a�=[��U�������\��Ь�H��6{e�_��h��`�L�z��&w:=���4U�L��&d���dI]ڨ���$�,����3�>X7z1YY��oͶݩP₎���o�L����A����ZLX~�C��B(�j�%��(eVWk�0Km�~t�r�$5C*��+��տ��\� U��_�lۄr������T�b�p���C�h� }��b�B`6׮��p9@�!�k{5�RT�l儍�N�G��W��Ԇ(o"� !���3����l�~a;&a]�w8��b��a"m���nR͔,e�7�ظ���3Ơ�]��=�����ĬsD����S�&Ir�U�Jټ̽�F��!��`�ڌ�Oy���NϿC���0���D�����?���G!���y��4�����L��8�e��؉ya�Q�@�\�
0�@�6$[�=�b���4�j�;���l9~<R�CK���]z�����CO-���T��*��C��Zch��cii���e��nǚnaP��C��(�Q����~�)%���Ox�ܔ����w ;�9c�ʯ��i�nQ�.��C�������=�^�$a̰*�f�1IX���%m�����	+��p	@vVV_.��)H���S�2���XGטT��(�a���E���]�����
�w摪3^�I��>���H���Ӊ����>��v�b �����sY*#Xh��R.�9�@�ܰ���G�/9WUAj�V�)P3;�$��Q�^���ߍ���N�ު���S�?�!�s����=�����y�}�Id(�
;��X�����ͪ<���݊�3�k(Ȉ�7����ʪ�c���>�FG�� �2���cpꢸ,m{�[�����@Ȳ��P��`hw�����t�#�"�H���{H�����R�ݴ��:�s��� ��N������B[�f��E7��:��S;�6�J���2�7����'�f�퇌� ʙ@PD�+�q�N �P ��ͺ.�q��Y�"��*ߩN��.��x�@�n��,�C���vsg��&��3��ƅV��XHVj?�<���m}�4��sʍ����k�w����r�A*�e���!Q�t!��_�\��mmL����'G|�}��)�8!h.�����%����%j���)��sݐ��ʽ�_q�G��`y��'��`��f6�j��AC��Viɖ�Lmd�8k y�;��+��)~��0���(�y ���z��T�h���8�W��yo�r�������b��g�C��vb��ZE��Aw]s��F)���{��
�w��^�Ǌ|y"((�����Es
Zӱ4WbI᳦��/*�.wD�DB����f��T�o#�[�# uv#���F�7InlxI^ k����G;�=@�c�oT�?�H�˞�)��u^�7b���W��K�|���4�{y���0�`�IK�=�Z�8����19T�+�.O���3�Di�����U�]{�n�v�]������$i�F��و�˻K�H��]�����m�8�$<K�C+j��`�#F���]߮�iGh�ऍQ�����9��:=������YP`����8���jl^��O�ߧP�X��u/�3ᄹ~2�V�=�&�v6� �w�ᛄ#�W�<rEB��XT�4P�X�������A����?%���!����=��vR߻i���L�+iExtK���`�A��U`�o���`N�'�,Ø��@ql�.��f��Z��Rf�퍬hCh/���0Y���қeCp^���|���l��qFpUW���{��=���;j{w��FT�l'���=]�ޠW	�y��ƚ��鉋v�;߀iz^�x�l�
N'�r��ʹǘ�h
u�JA�I�cˣ�H2ǑLgd���]s+}gk$Ă��ދ,H��cvM Pf���L�޵��YR}LPH����\:Q�Cz�:����q>
�/B��p��׍X`����%��ƋJ� tѴv`�L��v|�*L�=h��~����#%��R|Ψ��G�^��N����bQ%�9��l�w��嫔�b��`	�ф�n%�-����n��\�F(��OF��#fƵ�Ƶ�b����i�q� �z����#�_+p��	=�=��ܣ�I�Ջ?N��DJg�JM���Nq�W&zA�z쓌\�ǌ4��e��N��@_K�F��^��'��f^�p�c�:V�c0���ä��23���<�7��#wG-(�=�����T5�Ua}��Psk�|���_IK�B����o����[HWxK�)�{�S��(z#�ʼT��ƅX��3��N�*���"�%��d(�
������,���q�h���Sյ�`��ŷ1)4L�j��'R�B6��:d�w
��j�lmN_�n�_�&HI�T��T�'��K�S�	�/�^��!�yٌ�)}V��o;&)�X9�X�-e�Q;�Cr>��������p�z%�H�+��rj�����Y6]�~˕�aϐ�/E=�Y(z���W,Q�ܫ�WcH��e�]H
Y��)L7R�6y-��,�Lc��?��۾F;�=8�iS�S�p5��cO�_Ě�T��0�t���yYTq�a9�5�)C8A�[� �/%�w�ܯ���	i�Gx&�$ �^9��%;�Y����\����hY�x�P���A���A�u؜!*�OЁ��#�U��Ld�����L��&"�Vj��;hC,�m��o^(f#i"Q�c%�'��s�!E��1�%�(�ܐ�A_�pEy��{�9F1�>��A� <*���K�>����ƒ�	57 t��@�O��+N�*l�gTD¼���F�9k�2q�e�����i���Z`�cH�yŕ��c��!6*��{�ZG�o�"��7z��V�Vi#���fb�z�R�{<�w��_10!�0e�]3V9vQ��`�@���Y~18�/s�R�)d+����.���M��F?�0�27*�i(}�dv.�Nt8�	��;���FR�)5��SוU�9������{�[�f�9���xm�^{՞���]t7����p�Յ�1==9מ�[DP�*�j��K��v��j�@��n�f�θu������Ƀ<w��a�KA���y�hE�o�D�5��"����"�]P� �Pʫh��a��/}�4�1�(�ͮ�Ej�ʅ�6�TF��>:�k����R��lc��FE�i��O�o�7������Z��yy���D+I�}��cj�^Иػ�R%�mR�T��cI�Y��@Q��b�@6:�D4a���^�>��S3	+�w{(�b>E+��*��h�@^	���%��=�|W�b�ad�$AU��
[�ة	,��؞��~Z=B����,��U���%�����#��PBmUw$�)F3:J�����"7D@C�ΨI9��8�1�V�潛�6�&���2t�����*)G�c�w� ���ĭ���o:��;�cW"X���
3����H���4Uva	��=衵u �aV�@��~��:`��py�.���i$���J�o:3������ ��\��I�m�|�������jeuB��D{P�d���؈E�R�q��ő�D�S1i�	n��ݭ9_�'���0�w����H_��{sFϬ���.�;�-j�7��_�_D�t=F��$�X F��_E\��>
n h��c�/�anLA�Y��*������B����,ӱ��4��hi$,x��hi�?Ϋ�v����%w)���@C��P�&b�og�g�q�լ�#�P�����$�勯��M���ܴ��y�Twz�7��Vf��Z��'��p��Y+�/��'��5��uD
�]�HT�]nWnw��v�Œ/c�KzP�ݏ�6��dW���n�	�ϩ�������|O�4��0{������y×�N���$��>��;��{����eVG�A�D�����x��"�d�����6�)>��9�T��\��b�ϧ�B[x,��� ��;ͧ�nCyf���5�4n�׮H���%���0k͇����~�?+�&X�ɣ�7ݩ�h��:dZFn*>�U~�����/5hI7ERc����_n]��?!ݳVGG��l�WM8�!���/�xu�ss��6�T�������h�l�������a��(�J��g�ےZ8�n(LN��ޭ��dV��>�f(d~� Q�o������6����۠�\�Ծ�G����T6u��ڬ���g�	��+pd�w ��{
Qڸ"�LN&�"M6'?��i��-I����`��p��4�|&.м�;���5KmM5��rD�/���X#kN�$\˯�R�\�x�s���*�����܅W�P�(5����m80sFs��\/��x,s�ϋ�h��/�h�)��F�E����0����M6,O��
����+�Ʉ���>w�^����8���m咑d�7A��3ʈo�9<9�5�j��Q�YQ�U��As���Y� ����-7zV�����<�jZ�#��	�G�G����y��!�|�����H�;�����X��2�Ju�c$}XQ��xCu�T�W��D����Ȕ\_6��:�V$���c��/��=��{�0�_�A��qp�&mV84#�j]�&kv9���Z��:�s�������H�s"��1�:��F8�Ɔ7y��8���g��>�Ǹ��[��^᫧a��ƅ�Dx�gBwpP*�;�F�*7P0�}J����@���ufiJ��u��u�?1Y�X ���o��o���{�6֥]�ڗ}�chL�4��(?�оR]��ƶ������Ԣ�E�.i!�Pߓ������\�u�Qch�F�DӦ{@'wx�q��˳n-�|E��70[�-�X�9'eQ�<uD�{�a�gY��\�`?�r�J�W���&��& ��4v�8v �/���i��`�-�g(l΃"�HGj��ȵݫZ��Pv�蝩-I�Q:����{eY��u�u��{�/���z����V$�h E�?��ΐhy�}k�s9����c�C�o��7(#�aƠ��wGh�;W<��hZJ�Q�7�ح���c���yF7��<5}M
�L�%x�Q�]|I��*��C���H�������a<j���\�R�ש�i]՛cE�B�W`����p���'s��04x�P��_f��\����)1i�T���ԏ�S�o�U��#^ɦ8��b�A�\�x�C*c�s�:vG$CH���n3R�ٿ'x��C�'��Xpj@Z��Q��T.��N99�u�5�A����"�5{/�e�ġw崿�;d�ǃA���%Gm}f�=��F�����X���G�����1���gwK���q���^+%3
|���#���_�I;��I�0�+���QHqu��o®o����=�`�R�SF98'�B,[ӕ��x�E���Y���g�CR���}k8��HQ�9)���3J{9���[zo��~"'z�8�4㸭�I����-���<�,�lsd�bR�L����rf�)��~Y�X�b�L��^Ø->N,�i�@ՠ�[��&��:!r�7��tI|�R}5=��m��B� UC���\��=fT�Փ�i�W2X��1x��k�.Y�L�k2��{����hH��5h�F1>@���/�ˎ��V�s��$�C{�9I:�TQ�jh/7���?8	�/��T���lG��x��䴈���=��-[��\H���P��O��#��a`[�3:)���{�����:k}�[��=>(�I�/��ұ�>��3���X�h�Ŷ1���S��v\�qB��]�eg}�ݳ���t"��;�ςD�YXA�(����!�I�3C�Ue��9$�6u=��g|H	�ĉg	��S��PUu0��:��7X�a+�˾�;¼�W���K��/Ȃ���t�¶}g��O�������!�Dv�ƕ�0j`�#o!�Yb\+����G Hw7W�}�5�7�d���58�S���@>m�%0\��v�{Ei+��I�ٖ�w�29�#��I�= �4���v�Q@��B&,k�h���������X��˚�AԿ�%�v���3���=���^�a�x�qׯ���58u��TM<����z�42�^��e����w�T��i��=��P���KT�֘���`�L-)��?���[2�<!��� D藒h��$�6�N'�nR[*�`m5�55��y���Ͻ����_ŉ��{1��P}�,T�<~<d[�1.�s�k}����E;��k�$���7f�ǴƏ��-O�&���1?�p3���nhh�dUo>�q�X\>�}m�U�n�V^x�7�i�w�F����ڗYs���Yk%Wя}���� 87m���,L���Rcn ���͡�29��W�=
���F����1!�ǁ�7�����Q=��j��Yd.ѫ9xn�ܣ;���.9���[�@���3�c�=U�ӓ��|L⓹�L���M�/�� �nWe�I�I������I`%�ƃj�)�r��k��J�F��%~��Z��Y�#�|މ)Sȁ0�V�w�ч�.�u����bg�s�v���%����ʎ�`���� �u�{����ܹ
��z&B��(�,��D�A��cA�Ë���{�y��SG隂���u���'O���:e&.��tC��*#N�K}o8+��Gn��R��V�7��m�O���o~�V��}ZN�oѾ��s���Yo�������4PP�Ԋ&���+B,�˹�|o$s�"�ѿ�A��8�lݻq	!�8�zy3w�E�����1��q�C�G�U�f��w�^�����$���6x�Ts��n����1����c.���S����t��K�(eN�n��������Gn��_Ǘ��}�ۀ���J�;S�Z3��'����
������.ʚe4�;�KlH��mel��`�_���Ԣ���SW�����d�������ڇ���0�1�:�c�أ0��S�LL�Ա�i��DO���{65hr����p��
����}u~���okZ�U����b�+����{�}ةUY�]h�E�N+�D`*�mZǿ��{6�QE�f� �>�O�HAU�� �DV�u2��P���u�'Zj}ؾ��!N���(�7Z�8�����P� ��
�ccoo���L�+�Nf��RW���6t�8^(���$YH���f�YZ�������[oj�!�'L a�`G�Z�[�7Њ�./$���>�y�ݵL�+>H�l�"?uxA祿��]h˨?6���v����b��NQK�B�rW;"���#Ɔ�<�������r���0D��J6��{p����4�����W���1;!���n"��[�W^��k=�z�8����t��`U=�b����q4bB��Q�h�p�L�up�j���_5yݐ/}^�>a�x��g��Mw\]�0�5$�/�B"��]w���V��)���ԁ[[ qν�z�H�Pu��c%$ȕ���R;�6J7U����a�]۶1y�mK'�P��J��]�q$��Y���$�Sݦឺ��.1&��� � $� �,V���穥܈&7�� ���Q�"UWK8�)�x��fHۀ5���!��8�I��=��x&�a�L�Q5���Y�w	��H��C���H ��<�/�F��=Wv4�}-�rsS�c�K�Ԛ���|tv�����B��z���Τ��������)c�nmx�y<�%�����]��K�< �(���DD��P�	=��ꎎ�%w�
V�A[�Z03X����ei`9K�=^گ7g��=�`,X�0u����<�	�2F����6m��Bg����`�-Ґ�cD'�_}����܋3\S�+�& �f)��� �4�x� p[��}�P��^_a���pV/�\Էq�ľ'/�^��Y��>db��'�ﶧg27�ˌ٩D!UD�Я�v��t0G�Ne� JȂq	��j]��ۿ�n ��SDc+F���fh9a&dG"�^���P;�n�Q�>2���N(P��DKZ�
�T��ɳ�%�����f��T�� L�=�?̷����X���3R��7��r���O�y�d�s�,��W���0X�t�u��ζ��#{V�8PoС���j/��u��W	���!"�V��l*�M�[\Pny�k?rŏ���9��^$dn�����'��;� � ���6rW^]��R����1��������3B�pg� n�W�#.�ݪ����PK�ȔC=�l�Z��$*uO��_�B�؟66��6���7��{�J�y�{d��ʳo��`XfRGvH�� �t��-[�<�����Uc���q��G�^���؇�ù|�&�{|�0����f�&_�����J؂�ɫ�pR�ЋX@�t����vm�\�!��5��i����?;�R	 �����!F���3��Ӑ�*��i�u��{L��w�Ӂex?H��r��	4^�t�鰜M�w��[�<K���)I��]kDp����8Ń&  �0G1e����]����6������3wKO�'�+Tk�VkN�0)��_�, � �5�jXf�eb��;~�$��#���}8<��g3��,|ɕ��e?�`C��t��{�� ��!�57U86{Q�Ȱ.��zo]�����*pU��v#�ģj6mUY�֮sA+�Ӹ����ț���+�g�D��X�弐�n���ȇ@ê}�JF�TcfB�h	B��Q,�k��[�}�g_�Nl�x&ks9B��QT ��X��z�ߛ���}`AS����uU��-���%���U�oJN�@P}Ï�T��=(n�B�rш�y�4f��קe�:�A�z��ܳU7u�XҜ!�������2q94l_��n�n:�P�7�0 l.�=O���d�� ��X2��Al=8m�]J�<�cr-��ŏg�}˔G..��m76w�{�?gs���T��&�)��|���|+b�����?d�Nn޽m��7�j�"��Qx�6���saG�B6TU$m���S݋Sk&�T�*��#�(kb��)I�����I��EC�FB�&�5��mA%� ���{=aB:߳��z���57��u��T��uLu�:eB� ���e,�,Ţ����I_��� ��*�B�~��ύ!ǐ�|~������>�P�$G��6���~h)K���1�O�!T�
��?��-��JԶ���<l�v���t��8�Lm�$�/i������P�w詚m=�ԃ*E��+\���AŬZ/��3ֵ�^OR��لD��\�:����z��_�. ���
ɫ���Mz���e��[��Z\R����نmR	��y3S��$��F��������O��^4�:1�pz_N�ߩZ��btO�?�=3Y������u�"�@o>%&U��7��e��Q
���>s%�� %�FU��b�jg�IŎ%�>��Yg����^B�.O������P��}�F?���Vk�YAS!`�������r�z�B���#�V�_�7K?���5�g@�F��)-2*�\���W�$���R��<ee��pO>*�$N?{#�ozd/�)p��>
䤁��(ʞ�����FL��4i�8���B��܆�	[��_�L��8��:�r���F���4�a�hESl��Al���/�n�K��'�W���Uʄ�K���\�ӑ�>Qfx��,&h��`B�M�H���g�F_T��|eU���z@��fv?QCȎ�
�� }���
�HR���z��{�*oR�M��9ޱ��bD�<��d�I�[s��Z�A�=��qU���ל��IY'd5�ϙe�:��*�45��l��ҸGn?f��óc��`?b	��c��������K�(ݳi�7�;v��F^�|�L��Z�8"DՃQ�p��,^���`ʡ��6��i)�U��#���(@¿��i;�A|c�@�f.�۰rNڟ&�aw+/�#~��]�.L+ |�;T��>o�k�D��2��SUj1 �/�X�>7�;#ڥ"�Me]�9	���Z!���m�QA�h�����N�Z)�)�z>��p��vv�NM��E�g�dI�� ���2�M��,8.��m�i�D���	zsʋԐ��Fe�ͅ��x<��x��f���k0ٽ�v#��-�2V¹='��-�"M� !)��Pjv��ls�.�]�RhY>���Do^�a,0nPa���6y�����?�&���\��%b��)Ѐ}�:m����
��C��V�ն�����r���,Xb��`��u4��R��?��9���O��jX:��q��i�Ն�oU��N���2x��}\�J��խ �:}}�S�kuy�~�ǂ>q.S
:$��"�C�ڞ�g	��L�g
]��Eģ���N��XpJ!�4��&�Q�s��1'X��]�	ਸ�z͠)�U=�2cAa��5�����2)��*����0�L%t������.�S�X�J3vt��>@ޞ�N��ʭ`H� $ך�"a'c�srC\��$�i:������*̑�]Q��xK#m$�w��_��:�.q*qE�P��������|Æ�0�=|W�Ra�_@���e��w���熟�Mu1�w��dg3i�//o��QN�W����>o�֮��h��oڀPt�F�䝰(��o+z�<�>TL�O��s
==vz�՝c��83����.���VJ}<>m�'�(�<��=d���u9���4�x�޼p��˧m�����}����w�FOB�%� P �Ť��k�b-/yR�[�<#e����D�����c�5GgL��� B/��r^5Ļ���"����:��N�3�C�h�D���4�^SPܕX5dr�%�䇰���y3p!�p�@����P�iP+ҮG2�H�T��y�k���%� ϪGA�Qh:�q���,g��:�ŷd�1|T*���_�_\��7�.��Z��5�����yzỈ(Z���Y۬W��|�#C'���_����K	�>2�=���A@�e�!#t�����8TY������k��^Gl�"o�"�N衃#��2yf��3I�j��w�Fk��y���'�av1\����͡Xl��72z�����Kur�����_���ĳ�)XC��n{�X�7�o�8�(ӣ�,�W�׋��76�io��kH�H���-��s�����7lWx��P�EU��'�kxFO�a|�Rc�PE�FO���!�<#���[����Ou
�%��h��3�05' ��� 4�D *���%�w�$G��e�1�.�s��'WUu�ww�Z�͖��ɲf�Gڴ?��~�������g$+�&���Cq?�wo;�s�\W�*�	��.una[��@�+�@=O������K�ktt"����92��dǩo��d:q�ki,��UxLBV��l��x�W�A�\���+�$��l.�����|
g�;U�kb�4�V�\ۘ��'�AhP�I P�n3���XU���m�5���Г6��ݷ5������*��]�_���8��'Hm�����e.���+��G񼴨E���V�4a(�)���o�-�n�������Ϩ�'[*�)%���Q'$L ĎTe�ҥ�qU�n2*��3?�� �ݪe���da���J_ >�.�\�b1J+��1n����tk�����I�lsy�~�����5��lH���7��A��\�J!Kۮ��=�Dc�8e�H�m{��j�|y>�'�:�W]�c��֒$���U�7}�Gb�3I�A�r������E�2�ҩL(I�N��(�H�X�ѯ�I��F���],ԉ/��˨h�Ŵ�/2
;�Hq�Sߣ���K�a.�u���S�0�Y{�Pw*zwT��I�ѐ�#�3�T�q󫖗6s�F�_���>lV����<1������`$,�OTu�S	K��ݲI0@���!KX����E���Ў�~��E h֋s�	K~���/$�!9
��R����k%�o�va�~*Ej�U�;�����s�4ȹ�X��'.Fx��	�1��
�$��Y��C�%�0{BӅ�En�۴�0uu��㚘_��T��ś���rQ��)�#�ֺU��B�V�v�n��:3a0���'Q����ZV�9o%1:R���ř�S��J_����R>b�	�j���"�@1iB�$b�=�seX<����}h:�7jF�i���-�4xF������i1{Qr�ğ�>��rԗ��}�XQ�R�47��h`�;���J���(��%H�9�0�@�~�����1�q/y�Xg�hra|���Eڪ��H5��C�4�beSm��#�5wu��v\Qr��0^��P�9�LQ�gk����|�]� �>����������i�On�4U�å`޸�5�C�G��ɨ����L��)��}�^Rtx5�D~�k�Q�8����x�H`�k
�˽�>e�a?��X#��MHK�l�,�=�^_��<��@�K��;���Ӌ�%^ל�7d�]����FTP�K])���8�.(Xg`�U��>J�Yk��� ���,�{���۸4lǜ� �C�I��:�s�y�\��ڱ�eZ�b���/��?��RB�Ŭ��o�lLӪ#zp�G�ZxzHc�Ɣ�S�c������l�ѲE!Ż�I�ǯ����U���<�I��ͣ(� ���"N�{lX!_cR�I�+z�����/Z���,nN��%���g�]��5�舍ht�t��P�ٜ�2X�f�%c<���P��چ���XĜ̌�+Ы��ǒj��5�0���+��"��ܦ����0����%�G,w�&���y��:6��������nkO�p� �0�^�F�S�S���x���>�$���؁�'���CQ���k�5)p�K��3Y̥-�`Y���9��kV��g�;��1����;���
�T��٬&/�N��hW�z�$�#��zǦ7�jJ0��e�g��'��'Bg�u��I�F|�@�VX6�8r�	<���Պk�Ӈ�J%�C����j�6���[�G�����Z���d�J:�"��|y�86K�εd�%(�n�Y�잉L�@!�Pu����=&���^
Lu^2�����P�9��C	'�)�5yp��S{N(C��sP�V�ЫH���(��!s"rf�PL1X0��R���G(  Z��M�g�SN�4�;�^�4~]�dF�_4l���C0��XMa��'k���Dҷ��y`p!F:�=M�R:����6�Pd�#M�5���f��˰��h�TQ)�8�̀�F*aF�m{ �YB�p{$�Ԇ5(�>ӏ;?UI�$;ټ�����@��Db�����M�!��=��$�xt�w��nG�]A��G(TN��󃶿 �m�Ҥyd��6�پe��I��e|��h�*�|�pn��'-�] �]�(���ԯͩY~S1���V����+�Z�EnG����Kđ�m~�����_В�HJ�*���f��.U�y��J���I�h��;�̶%*o��P�t$d�!�@У��;
!�wJ�:�s����D�έ&���ʡ2�sG̝A>Q_Eu����� 5�	���ʷ���&�#�#@��yֻ�i��殍]���yj�S�;�� 7���/���=����j)U�RPX�I�M��ґ�6p<[pL�G��)1y��>�|��1��m�6B��N�:��$�AE�Y¨�Zv�R���!����e4�b̜F��[s��ޖ�1�r�{�|�K#��+�U���,ri䚹hP��ƣ�}���'ŀx���W�|xʁKf�D����f���]`�����2!����C�o��Z��P�	�/�hZ�(�r�s�K�g�����ڼiKR����s�
e�:;Q��!#�U!���jQ�_�!G�����72�ɋ��<�8}���k��v%?�@��T`����\�w�k��O$	$b9{���0ITI�.6k�{y���m��q$�Vc�������������v�9\�4wU;�6��`B����]�cF�3�N�!��c+6�{��nc��P�)���vgE���)d�����zs����ҮH�p�\��E�AE"+�P�X�(uH�.�z�@�8��d��h��(�U���]��� Y�28�z:�
~��=�L��o�$�������^ q��Vg�;��ը�1�O�/`�"�b*�jv���dk_��-�ίhD�w�XSU�p���&�U���zkxb�u�� �ߟ����j�K~�z��E�Ŗ5����x��ve�����|R���h������8,�cY�0��Z�ƕp�!.V���&$��k/�2��*�\��� Z4��з�
�ϪŀO����P=�(�y�j 0�#�B��H�U��2a�u�8��f����j���D� 0d�����A��`@���Q�-���C���	����V���!��(n�ze9tZ���ȍ���w��V��(t�<��X�{
{�jԜ�W�L��}�ΛK��i7��2'HAE�v��Ԕ�8��tɍ��z��.��o\N2P��.�X� Y�]aUތ��Kg�����_���u��R)��a$y[�t��F_6O"x��2V�a36���×�R��6q��E]��\��#c�P��#q�c����Zi����܂��@*-I|\�،=l�6"�Y�����$�A���%����+�cۗY�aX��vvtp�/3������26�l��N��$��(L!@Ŭ�Y �گ��w~i	���_��|x#�z����`�5i�A�8��ڴ�tn@�y�����|OxS����&b�뼸�|4�#g!N4����V��5Zv�v�i���|8
T���X��I�1�hr�D�tJ�#��3؛V�c �;���/��hx���=�v@�����󇀣'�V)m>��<sf����'H���|e��e,ɝi����<0�����ͽ����]E$�PDh�x�<�7B�](�zF�)�jOZ��1��M��6�6^ ��ki@@%N�E�g\�(�N|��R@>N$�b�i1��"���p!"sh���ܬ� )U�aP���D�.:)a9;[a�����0%���E����1Zp����՚K�y�ᕐ�����±ya ��c	=9e��㧈�-w�]nΝ��(r��d@&��.)qWʜF���cڷw,9�ǿ�=�̑xw^�iK�b3k¹qX��E!�҄	�C��I�n ���S�Q����b(��&[ޖ;���+&�O�],Ea��I�I5R��Y~��4c�|�I���N?�"j�åe����;���O|�� ��V��8�'� ��xR`c�_k
�wF�Q�F��t��0��X���t8��Ya4�	{��P\��T���+U��5TA���D>W����I)�*g|)dW�<u<*5R�P)��g%�yK�������c�eu����cvÆ�~�����$'�S)�y
�Q������a��	��*��V�|�b��̆	cp8�0�$e*�|,�m��,�������:�ѝ@��Ƕ���iv�st$
'�:2���KLa�����]�4G
��&x���3�8V��,���i~��\�nOڠ3f�J�q��4�(����~�O&No�8���+R��������wJCqy�x�,f��6{(ae�IdK����E3�#	�;�z&_����]��g5�]˶�#�*�&5��ph��	�m�N��z���ѧ��Po��O�_�N�]E.o1*��M���x����Uz�ww�}ȷ5��a>y���2ٰ�*��󕞷�3q��m�e|I1�Z�������0�s~ק%�\�o����&?�㯳�®{S-i#��Z:��3���V*����;ǵ�E,yB���	����ȇ� �G�������Q�j���tO�0�~�q����3�9 gYl�+�Ao\�^�"��?9}������ �%��r._��O����k�����ŭQ���$F�K4N��V�4�J���Y! ���S���7�}�ۡ�j���@��v:V߳�2���R�>��ϡ����߬�E�׾'�Lhb��V����y4a:�!�AA�aԲ�U7�Ph����\)����9N�P��t���.c��Th���E��S�@�=ݒ���5��lZ��mo)�l�~H�E܋8�U M9`�r��	[tb� ۽�j��^m�7Qk�G��`��d�<�W�ށL"���K�s�Y����3F=�B���`.Ӳ�V3*g\z!<�Yk/q�ul���45#���E�����sH8g%��m�s�zꎮHkL���ID��*'�(@�b���S�w�E3��f���fXV@�1WV�D��)��A6˹�ȗ�޽vMS��5��X��C����{?��ߩu3�l�C�OR5KUR��qʪF|����X1.l��)���]xL�� f�x>*��(��M�Q@V-z� �,�"��u�srG��x���}�vY��ۆǁ�W/��pQ��p�'"��ˆ�A%9$���+���:�	��jQ�EB����X��~�Z�瑤�g�F��?Q�[��c�ϡ����>J�hV��/���
r��}�`{�kj��.30E�5���@��������G�,v���8�b�B�*ƹD�0���b��R:����*�ÞɖY�w�*	����㒦ţd��VT�/#����+�.�+�X�dx�M]��2M;���	��8��̫�ɂǐ���P�м2�{�6/~'����X�h(L#^���2�%ّ�"��:-�*Y����O��7�|*����	�ρ����ā���Ϲ�ǵSKY���6HȣLxO/�ˀâ� �Kk��C�'�}q��i� 3��l���������pRC7�����!����",`֓�2���IVD}�1�;*��*1�L/ѕ���Q~e#��b�{hx�;��YJQX-�+�N�| A_<_�?f7�9*	����u��J9a�hX?��MmkPžvŝ�H_m�
��Z�yl��w��2>�#Qv�'޵C��Ƿ�9��o���~b%[�C-(<����)G[��~�"���l��	P�w���|Q�X�0:��3���S��鍫G�|�J��F��d�#㣈96PCTC);�8���w�A	�oI�*�N�x[\��3Xy�����d�����xY_��PU?4�+2N7�jH��8�K������\�8�[�c)��8ƨbl�Jg�(6���'�`�X֖�=����)�`(�G`���ǣYq�2��,�v���@�9X�B~7 �ZF���j��2�xlӳ̬-�܎�*�T�v�r�e4U`��9�̂u[�'$J+���n�S�&ڹ�U�Q�W�?ý��F>��M*�l'��Pm*�#(�k���S�T"s#<ݨB���t8�4F�x�����:�TqlA޳���Y����*Z�$Eـb��l)y]�?�I�`%�;/�zl��+���WE�rz�����'S�i4�'�!ǋ:k�h�ٮ)�V�ۨ��6ܐ<U䩆�5���v���j�d=�ݣ�ed���<����G�I6e��r;=�����@�_��fD�^����C�y���UȂ��{��E��ŝE�S:L+���+�!#E��~��%»����P�H��W;hU�[�����֊��G%�	���5�:��c�٨���]ة�8&)�}��\��A}��X�Jv	8�G�K��X�Mp���;KU�$�����vW���Rն�]�����n�[>2mxe��`n����}
��@�vTZ ��~yZv��G�AXF���h;�n諰u����O�1/Pp��s1j�<q�U���g��n"��}{k��c4���ee�)ۣz����t|Av����,E�����
��Da4�j�Ž!pΧ�S"����x��PӘ�y:јq��'�v�^`������0�ɏ���ROs��Q�:z;�AK�[����)R����MZƧȔ����Ab��a���<�&"ț��E�z�1����{M����Ls��J�\��;�?W&�(���� �-J�}D��y�qv��̥��X�]�_������bJ��!m��iT����a��h���g�ƮR��[9�f�q�"�Ş�Xs��@S9�Y�fV�S�aمQ��SW���+p��0C��{��)ۑ���WowƊ���ڒ�I�n���Ͷd
|wL�A
K�����M�٢<AV��a�v�$�Ô9�'y�����Կ��0������p�����,B^ɻo�g�S:G~�*�Wցl���A�qX�����j ���t�F�S��')`��nX(>)yX:XC�;�`�aR���L.ME�eʕt9���7pK�݀�ӧt~9F�G&`�f�0���C�]�mxM�8��!G!g��N!�$����!�77�^С?y<~?)C<��{!��!�BJ��nI���8�\�D��BK���bҚ6*�e�g-�^�	�P��ˡ�c�C2}at���ܗ�&bI��#�5lM�J�+�-�2/S��������Ff
	����O��VQw;�~O(�i��+εX۱��)�T�T|�r$y�	Vˮ���ӛon�Kwl���!G;L�w�R!�}���]�,.F,=K��d�����,�/�k�-���d^�i�-��I@�O�2	y����t�ȚbM���;�=�(��7$X&c��C�c�;�y�#��7b�
d�	)yw��	7��ح:f���#ْq��Cfd��{��6x4:�g9��<�#��˝.�Ǌ��e����k�/�þh5d+&�eu$Tb�=ɐRCi������.d(��.��G��D�_��ϲp�0��9s.���PĂr��Z��2r?*?�Q^��p��tkѶ��|��,����_�[
�4�8��X) B� ��H��=~zd��-�h�i�=,��*���t^�k?�5��!�kx쿊E\�:���(<S"?8C�M��07Y����lh(`"�\�Z4͜��F�mT����h���1�{�u,#�/+W|���竜��<
㑅ʭ����9Cz0Rcd�픪���mH�����DR��f��â��Av�\�����/�tW��MQ��-@i(.	m��8���i|^��P�/�?	�	o���NEd7��A��*K`e^����RS�7�hC�!V|G;ܪ.��`�����2�U���~��0�k��C�.	I�_��豮C9~�I��՛�m2����ԫ���0�ܟ�Ø�t�Γ(�p��@[Y��K�����
���N��/7������SD�����v����'I
̜{("�-ـi�W����
�,wӅ]E@f���>���/��?�������T�&��Dv�@��\��3���J;����e��`�8�5����ꎗ�(���]_����Z_��SP���+��;�IőBW~&�}0��i��WXZ����$^b"���o6-��x��%�)��A��wv�
v<�"I֏f�jطF�� ���i��SAL�cw��\�����O6'C5������7�Az��Z� u���&��XEڰ�16��i�0�S��g��5�gt��Kx?�=ۅ�$ʖ�}���n���|d'Qb4��-�|�y8�9����������ǚ���z���)�B@|��ah�L�������8���6�������+>G�n��4�]�^��K�X��u���8&�³����S')7�F�F��P���PṢ�Ej�U�B��M�	�u$�]��	D���1�C���O��yz��k���}���um��_�2s�$����x�����؛b?�N�R;�L��|9VL��'N̊B�u�Sνr�X���A�W_\�)�C��,�yNC�S��l���rv/�$(z��Ɲ[�����^���{T?Tr�b�ࢪ̝]c	W��y��vt��o��̉ �K50V���J��k'��:�㺚m����a�b�8�_pp<?S-�B{γ�y��l��tr/V�M����GX 8��Q�O!���<�����
`�?�&�~��S�w�^/0�Mvs��;Hߣ|�V~�7��������&�@�%:E֢ܴP`�c��=�D�tC�o�zY����+ ΃��R����'DfSɳ��"K�c��#���
��1�ڇ��/i}T��e�� �w �<=�'=B<�(���{ Yt W��
���#�
��;9cӹ$�Zo��S��C=�mUb1�k�X�r�{(�@�d�q��`�NP�A�=�m��9X���2O�e�(���T3�AE#Ԏ�����Զ;¨���seŋ���5�:+���i�z�,��Z��_&��4X�o��4xt��#l�K�0~!���5ɾ��<)(1u;82}#��)moX<��⒏��2L쭳�]�b9�r�3��̆��5��fϞ��vH��X�n#c����[Iv�˨��2��Rt��E�bu+��:j.w��>�pHyh]S�����&Cu� ��T#�i��ؼ��!Uc.�a��g< c�}�-�8>{���z٘kw1�+.�QG+T?��ﻺq �?jR��o��W=%Z�w��/���%Q����^ڧ�|a;XX<��P
�0��������K��F���Q�^>���c�D�P�&Yp��DB��w/��A�~z*2,Խ	�l�0��n�Ly�2�:(�1߸B!^,z��~�Nߛ��"U��BL�m���˽|�s:�]���W����J��c�5���Ǔ���2R��i8�N�^��&�u�$G�d��=�M)��"��!oE��%Z9	N~9�$�'m�����l�%NhV��[*�Y~z��t��K`�)u?/g�~��C�iL�}cN䷞� w�q�M)
��ſ�;P�=��T!R��tK�T��ڝ9����mI�U������i�r�*H�&Ho�ք�_?2�
yXg�U�Ɓ98+��cŵ|���1��ǲ/�O}r�n��� .H���$���\���Vl����X��3ǁ����a�C���G+f�Yc!�IS�LD���2��o��YG=��ep�WqW�q��>���a$�V�M���8��'߻h�)!�Ѳv�ޕ$���*A-�pZ��)�}�,jw	{rȹJMNBS�=�@�19��`��|"����9���+��WV�"Pd���7[�v]���I)� ���xY��縄�L*@4N� č�����mft��$Rr���s㘾� ���X;�/�_�f7~��x��]b�$���m���c"Ȇv9}� ��8sϱ�̘������c�,ƶ-����|���z�	aS/�d*�����;���?(�z��?̕���A�J�� ��Y��O�!a����<y�+�����AuS��P�s},Xh�TsϲN����#�?#6C �s�ʨ�1c0Fτ.��;��������G!�\^l3$�K�2�SѾ�kfu��.ف�4J�7���ud�j���{:��_8C��K��XD�T��e���V�R�h�skm�V�mF�5�uz-���W
��V���5�+�����}<�P���Yل՗J y_&f����6Y]�I�N��,g��R��邼��*�H1M����zh���S�l34�X��Y�?=\`���M�4E��/??�m2�J�U>&-lo����)����	�s_����������q��[����y��@F2���0�1���aE,�0̺�9|}N���X�ҧ	\��C�C-���* �ԠǇ��p�TZ>B�_u ��l~?qp�5�5X��+W@?���'u_��3~_[G���!�8�̎Iu��;�!aV������λ���X�������Ml1~�m~�,�R�_�f=;�E8��Sᩮ�`�q�0q`Bҩr(�����~�5wFB6ukUw��S�qVK;�^{: �s>	H�؜��ƷO�o$	W��ݘu��ʮ��+�ˏ�BC�'�����$�3Ė�b�`��'�r<�V;;^�;(���(����W1Oc��6��q�r�4!mh�G�(Қc�5x3Q����R��.ǚB��O�8��n$F�۳���`�	���3,\��E�&��6�{wVo������׳11F}>���]z�.��>ad��	zU*]����قKi�$��暚�`hA�ng�b�TT.�nα/��:���Abk������y�o��oA��o�84�6�	�K��.)��\I%j^	�{���`�l�7D���u�������u腡�!�W%})IL5(���U�Q�\�SiJ�P��&�!tj+ćW�'�[�}���6��F�Ӫ�:L�q�+v��T� �M���J<���#T�:[�r��(��3*<��cJK��h�g�qS1@�,g�&��]���8���q�/R@�%�j^ͺ������G�|��8��HT��k:м�*I�Ѱh�N��`D3�B�(�vt�0���G&Qs	IPN%�Sr��w0kPd���)M��x~��~�<��]3'a�c��pV�ۂ���J�3�cq�d L;˚�Sml���u 3t��ՆjU'��I#����5�1�^iϩ�O���;���_y� �Z(0\�.Ǆy��#�[�S�Ġ����X2��=r�$�׻.�U��`v�8�3�������z	�YO>�>���Y�#T�b7�@/��/D�i|^�S@]� ��肉G�`)�����N
�����O+a���^a�9�] �G(g�nx �TGY�7��oE���ߕ�kH�dck�b� ��U�����fq_E�*w^� ��n�D��?x@��V*_g�(����~�p_	p���o�H���'L�2$W��f��͵8�����9�i���W�kj���ʛ]'�?��E�E&�o5$9��`D�-ԙg�)���|�7tØ���E��,���C��G�y���c���w)����B�/���3�.R���}�`!IP'��e�{&HQg5Ł��x����9=_bp-KP���k��Ҁ��׾�@��5�}-��
F3�::������c��KY&��:�e�������HJ�[oY�5y0��0p�|�k��rJN�����A�F����h	��z��n�g�g2?W���k8L�
�VHm�ݫ1K�G��:�KV�C}�9�<��1%�� *U�8���\�s~����PiAÄ&�<M��.U�^�vM��8F'@�涡�׸�,��ѯc��=�}�Q9��ɩ%t��]Ap�{=g!Yg������8� ��2����x.X�>H�~ ��-��0�ue,��f�T��b��ý��2���ҿ���{��ܔ��VW2��ւ5%�,#�n\0�H� C�z��l�NR�QM��h��M-8C�j7�|��wDs��g�ʮ�p�x�@��]�*�a�劶z���	8���g�}���0e����V�$T�QKRy%"�6�|�r��|e=�7��p�/��u�>wy�ɧ	F8'Hj����J9N
���X����>��u�A/b߇Gf�e���(����Si�����t�����7�.��q׿70L�`K��=\U��[��%�$ʤH�a�p�k��SHع�p,iB�k5�������Aj��W����9�����[��|M�9$(�pq���x�K�K����@'�a�����S��:�j�0���������}�~w�͝Yk��Q>5�&�h��G�j�<����O�V�����d4cXF����5�;��W�3�iإ�_���e��GNh�H���oS�]:���=Q\fԩ$��Ľ��w�ו�Z�K9���0g�����c�y�QO[�~�%m�KyHU�ҭ8!�eY1�@Y!�9Ub���sD�<���D��]#7��W��X귿H|�U,,���Mh�h�nx¢�7��"�t����5D�#9�����7o�O�>�#P�$���P4 ����O59J��緑��-S�wM�>;��0�8e�oŶ�yR�.4��d�'��#��>�n_D�Ţ\�6l#̸x�v�``(T��1�X/�{x�F�LΑ�I�	������o-�P�%�Z����F�%HM�,��e/I=�����ܤ���c��%��h�4���cN5��\k2�ߦD��p�X�bY��i�'����@�ײ��ɐ�a�6��ܐ��� 2e9erFUj�M&���B��:!D�x���1�ЉVU���1�P�ٔqž2��D!5F���yE!J}�u$����/�:���_)f�n@W����8h:2�8����? 8PU�?�)�����e�s'*���m�j��_x.�8�0��ԖC��yx��7���E�$�����(�m�J��כw������tY��d�l��\���K�ܝ�����'�hwh#����������H�����?!n�i����^���YL��o"�� �$S�>o�|Zif�O�`�۷Vm�G[x��k�5���i@�S+��%�%ΰ�ƍ&&�5B'������_`���,�C 8j��{v0��|��@1��*�ŪG��̥��o��y��Z;�@؄t�%�_N�8�"1�s���{�Q���q�2�BY����+����ᕥ�6���qX6��^ื��%� Jm~9Plԁ/��8�Zw��s��1����~����z�RGC�|�n���|����D)H{GkI�[R�E#&�=UN��X�$-��w�E��� �\BZl`�yS�F�B 5��*�~H�F����j@[�w��T�#ǸIi�����y\x�Qg���JO�x�(�q�B][5� z��#«8��fN�t���{_=�ɆUJ�GdW�W��ٳ��c�k�z�IT/¦B�qX�"�!8Ⅺ��7 >L{j)
�&���3���yh�]kO����{�������G�Z��q�N�6��9�G%%|G�4��I��`\�,��i�	"gPz��� >J�.=��z;��H_����aBV�ɓ��8�����hQ�Tx�%����p��dj~��@���������8��Q���bPeXÞ��3�v�2C��<�)��RЖ�E8�[��T���j�R�`(� n�'�E���a;��w��_�����Ӏ6�> <��QR�i����E�G1��!���,f�t24	I�00�U4څv���x[V���c���O3�W��/C>��}�X
-�c����RAo�����2�88 %:���m��m�޽���Wɻ��_��+.�9�t�a��6d�[?�|�f,O왞�� �P?q�)5���lRj*�*��(/¡�o!k��[o]��W�Xgj%�X�B�! |H&̚�5t�&،�0�u��x����0�jԹ�TչRZ��ȠO�d~X�#|�-�Z
�U����,*&��.�&��tu��.V�ێ��l|��5�jP�`�(Ƭ�$����8�t}��l0w��i�	��_�����Bg���"d,�3�
��\�JJ�|A�x!BXC��5�5�@4@��k�u	Bΐ��2\��h*W�޳*����^�}W-�ȝ���X�ж��o���('S�G�]��Qv_6
*�6bT���b	��(������Eg��-%ܢ⵺������O!��ct(Jn��|�}�;��C��=�o���>�m,��	��R�ݨ�����e)�ĜeǽJ*���nGuK�SAB��ጁ⎏�>�m�_�Cl=M��u�kw&NY�p���h) �Uz�G1[��:�N��I�3���,/̋�q��Eh��u࿱n�x�F;��n_s9�F���Ղ[���n�,�� ��`�nDl���.a��b2�3< a�����+��������>a�?j�&��Pf!���"^W�PE4�TQ�W��m:I��>��!93���!�P�[��r=Q0��@���p1	_��>����d�r��G?t3�餿	�����@K���!��LNf�o/��`uqi���7/J��	����O[��F�^��g<�\D���0����W�A r�Q�)���	A2����������a��
��e�!��DU��m�{>O���y�S$t�1���If�Oz�5](]~�y禩�>�q��X���=�µ�a|�!e�KT�h(q��"����F�0c��mo]�(�Ώv�����Ԕy %�J�k�]��-5y~.��w<�X�t�2W�~����I�B0�zE��(Ν�K�ԭa�uZ�g�}#~Ye�@=a��e��x���d��?�`؉�/�po�?y��i�r��3�+�ݓ��:Y0�
h�k'@�+j��=c���X��I�c $�R�'-���a��EwX�N��b8 1]G��zT��ٓp�*e��e��
��&,��z�ɋNTfcz<6��-n#�i�*q�e��v2^���h��]�:S>��pB��
�Qe��蝄��[*F��<����D���i���v��2��(�B�~3�2��^�F��^�W�7!�޸�����l�Pc��C�3t��W{�w�����l��{y��:�|�,�)�ld��JDAL}��0%���;��=Y��v�՟��)nٌ?���r�!�N�o���%S�!���>�^��&Zi]�����!�C�"�����]Ht�	��cA�.����f%��c$���e*�-�o��7n�xJ-�u��&^��pbV�rL��̓�%6	?@��	�d�)߭+n�r�п�V�F�:��hs�8P��Y �c,���|z�$��c�q	�G4Jd[�dn���E�E{����c@aB�,�Ό
@�i��;z�x�l���-��;�L��������xƉ��4���]�UF�3[	�qKz�3�I��t�6$r����Q��ŘP��>��W$R���R�^e_)1�Ә��|i%
\��� ,��D����*X�!��b"��9Z���V���h�c��tF�H}pI�����=Q����?��*z�<���xi�ҟ'���Di�����V����+߲��<m�dJ���G%?���h���� x��}.��n�p�AG4�;�.ʳ��mR|�fJN���&δ���&߀q`R�2�{��u�zP&�|��1�՜��5{#�wtek��ꖞ1��^e����ܺ�B(+ȾV����.��x�ZM�Q�;��!��'6m
�q�w�l��A8�G�6��`�i���{qE�/��|A`����_B<G�5@POߴ\}^��j@?��xQ�?�r2��
ʥ~�9<�	@5��)e-�ɳ��?�inV�31��B5?�#�t�|<Kv���N?�y����ZƩn��DҢ��2�	��w��Ҏ��CI?����JMin��AEh����%釈Gf�tD���πŇ�*Q|J�|S�X�S�y	����J�����mn�e���Qq�I:r�ޞ��LnR?*�}�ǡ;S�qQ����
�L@���[�'��z�rcNTz��sԑv��9񜮰!Ws��Je�Ԕ�[p����A@�2B��*� m�ic����?nq��}Y�Q	Z|ΰ���t��@�)��~ɍ��(�4�~�>���������b
X���mQ����$�%�M�G����cv�!��g�(������C�(ȿD�&�G�Ϛ�eM�����%E��X�����T��'|�XzI�C���X�r�X�*�;bU>�*�,ot���ӻG��J�Tө�u�q�[����d�7=�1�۸�v������.iJ�Ǖ<�r���T�G��k,wl�Kf�R+V &t��wI�[�Eq��f�~��8+%I`�J~�d&C���qi��jC/&!�\w��g�@k���!�[�_<�xſ��7Sr�.3����-*N�j�~&�޿j�%�?���?�G�R:3c���=8����х@�h�D/����{�M w�3,) ( g�zHaw�Hrb�e�X��6h�2����<��a<��?d����S�8Q�R�d�p�5�Ǒ��/�}�c���D	�0���5cdt6�,6P~� i~7��S"(w�|V`����!V.Ԙ����i��s���W?�ĸ������w(�����7�)���,㕣����+�Z0-0��:��~�N^F���;�v�Ԕ䰾�	�J�d=��6
@��W�u7��g��<�DDc�1��Q]
G�K�?+O'R#w���1�I�p6 *�?��I�W4�j�Y�w���l��V@�?���.(�h�1�b�#56��=����a�)f�k��f(�xo(	���o�l3�
��aVw��*?��%`�rZ�m�,`3qW)�� 14A<��P� �Z��{_����}�W��H��W{n�(Ζ���_�
ف�G�����WIj� �mo�T�V�#�	�r�T����@X1l-���퍷�����T'��̼�lj'����vz�nԿq�d�+��I���%��;�z����N|�I�.���,��.S��\��z��Ӏ����7R_�:�����$[�#�/' �����9�ķu�%Edb��4��Oy�W����4y�����Ѷ�Z*8=�_!s���mO���*q�C�K¥-u)��J�LH�H�<�e;��iAi���NT�1.Ed�.5{^��B�:i
C��J�)��6�a��,���������������ɣe��Y��!qD��X��ahhAkC��ý���6h��@�?��i���X`psd���x�?�E���v�	��E�wSj����R::�Q�׷~iZ���O�L.�JK,d8�0�4�؎���i�"���(�� ˁ=�	��C�,}I��׭:uM
|��l���@b�A��z���
9���x����s����0�����*����%x�N)�NV��&:T(\_{EĶ���T
�*L��5���x/mt���h�R�����%u�cKf�\�h%}��:2���f�@����UO��k	n~|�t��L�i-[22r��U��䃪k���%��R��$��)��VN�N�a�5� 2+���a�����$m��@��iC���_�`��+t���$�E��x�;EhM\c�S��-�KV�E\�p�8���:��V�(��%x.����K�Z�o�
#�"]y����dHN��_�M}�HC�����L����I�������ᬍ�(%��5Iz� ��5�,U�#�ٍň�
W^����1�D���3�PQŸɥ/S����E65�RK�دE��Y�>.��eg��ioDQ��<��?{`��qόL�D�<q��Ao��V<�a��tK �h�S�L|:4�;��J�w>張���<�J,c�6���U�`��7����4G��=	Z�T�����$,Lt5�T��-[�|�ۂ�Vfi��y��b����Mz��fud4_����c*����CjFF������@)�O�=��l�%�h)	�j�̶x %�i����z��#�K�(dې�|֎G�h�:T��'��슼t�T�fĮ%�>��ww�<Uʬ��5��NE��*�#���������j`�}b�z,My��7��,�f)��ahg���/#��
����#�֐��@����g�]hŞ��8c1� W�8�ٚ��e#${���b��Z�_��q ǰ��H���%ser�z����s��l���k�*��#9�V�B��'m�'��
I�N����E�Y�?k��{b���d��`�%�/�������<.��~�oA�娠��"Se��-���N@ �J�=�����#&w��k��H���	��-#���ܩR�p-k۹�*��\N���m��`A4��9�����S�e��>��,2�����ψy�P]gf��ǅ�7��}=��G	G"�U�ajU�m�����|�FD��u�#z���S����R�1ѯ�p镕O���#�P4�<�N@j�bF�-���9*�|��Q�|�{_�������.����.��
���J�J�P�f��PcTɪ4Y2I#��b��|��ͪ4l���8�}�K�%D�������	I8Il���^���иP<��� 3��3��޺�'S�-��M�05U=��q����3��iZ��%
��R��$�6��8���g�� �h V�Io�]]ϑP�t�]�g���|�,u	�:�Mf�`iS��2��]T ��ՊC�'�j%��g��6�O�>�c�{���槂H�jE�xV���$vJO���8�갏C��c��N�0y�ǉ�W�?J�䴐?\JA�d衈x��\7�i�J�~�c���v�ƺ�/� ���x_��� �y�hX��jF�yzszx�b�eg��<�W������Pd�}([���$�Bg�]���O&�<9I-Ф���kYZ���2�'�����?N��z��Ans?(��N��jX��^gp{#4�4��:,=�D{�Lcy��N��t���΄ŋ0� ���:��1L �q�3�����%���%/�ʮ�q�X;p�1�u��( h6ؘI-��
�&N���0xuNkKS�{)��j��a&[���?��	�˽[�a%Vȭt��I����Ǭ�o}Co�v��J�)�h!e ���HdcE}J%	�%�t�����uM�����-���G\:�"o�A"u>!��0�JE�Ƃ����L��]�D��C(̿Q�A�����Ƌ�,�W�	�È������@�Oi�j���w�nB�vC2޶��j��
s�-=9���9l7�`'��w���c��!㖻�	�Y���*�g뗉��`!�kuIJH�ye1��ﻧ[OÖ���}6���!��ǟ��FE1�	>��-���O@x"]�n�����I�v��ڏ��g>�ϙ��t ���mB����ۿ�cI(]@(�^˃��p����À�= �U�������F|dko�F�[�������Y̫�Z�aɹ�'"`8���.G�6��^��)n5�E:����1���	�����yS6��J2B�+u�U ���4��dg%9۰ex|�a���[��k������,\�.�}E\���V�����Xmy���I,�7%�"��ݻ7����>�����b��)�b������	������s���*U��Sv���iڹ��/?�`:.Lԫ�p��I�Me��դ��7R�y�v�����HW�r���Q�#���hh����d���t�S����迉VY�9�ڛ�VF���̳�����T�S'ZCq!��03f��O,���]�k�|��
�/2��-a�o@M{�.wM�G��#�(�_�c�9�ǫ�����z���sr��������7�Ӥ*���`3/���_������
m.�ɵ�*86��(��0Nm�X/2����~��R,�f�/��!/��ˣ%S�5���1�}�jx�P@�݉��w���3Fӓ��-���f0�*�R�����	��OG}�i����Y�KQmd��Qr�7$�����瀟�y��� �hR�����m��Ew%�C�+�
Er%�����Ͼ�U�.�!+Q�P���!�;�6
\v��Vr_�����S�%�b
	�I0�)l3�>��l�a;G��3�'n�β��q;YC/�L��v�/UG�.X�^�9�oNˤȳ�W)%��A�ݜ���R)�ޔwnx�ƭv%��݄�P`<��l���Q�ˈ3�Bm��&HB�u&�%��d*����> �RQ@�"?�ڟ|�+ܟ;?�̵g1J�e�p�.�]� ~��MoM�b@���D���N���|_i>:X��t��=���@L�jl��$@�SA��=nQ�*GJ��s=|�|j���r#��S�~� **h8�	���d�SUN���}ir��z�|qI�q��2I$�y�jM"Mĭ~AB<W�1�C�tX`~N?z��@V�7���a֢�_�t� .�3�Q� ]���_T�;��xǜ�*s�Pm�� IoQ�jgN���Ad�a��5��sv��8/�6�	k�"s+v���D�2b2��Mz�3W&4�ky��<��6�T��3
�'�W3)G�(�֕���D�e&;R��,��S��0ݾ�4~����h�	�
!�G~����K�Ի>X��G'�a�^�be�	�d��l�嫳8Gw��r��h�b����Cb)	x���g��'b_���wl���X�e^�L])�L��G������ˬ�Y���$�I����D��D;������der]�۴��C�j��ܚ�^��3��z]'�բ�ǍP�=z�j(�����Q)ߜ����ֶ�U����XR)92��꡼�=������@�! ����j�R���΃7��^r+F����7ވ���������!��]����߀nE�fS)c�^�1b�꾷3I�ni&�-��9��s��
�p�)�Բ;h3�8gz�T>;A���[8x���?�B65�l�Y�p1��K���J��R1��Ǳ�Ǳ?���*ĝD�5�%H33��vN"�q�O9Y18���4�dÖ��b�<�N�A�E�8E�3�DëZ� QS�e�s~���ŏ�!\��4	�iV�2�D&v�TN7�� �~+�Ӵ����������tTƗ��6P�ǹ�DY���G��<+�eB�8��gd��T%�A�Rq��� NU����m�R����%>9��s�n_hc5[7Ԫ��9S�uQ��r�5��3¢�����͔n�"@�������;"y�7�P-oe��)����^��6������>�Ror��#X�!�
�a#盰�ϣdҤ���Sj��4fQ\oE��1�b⇈��%�K��;K���*���{����D�9lg�X�6��W�u\'������ ��j�Y#_r�X�>!�U�{P�Π��ύ���qj	M�!�e���4[�?�$�A�K�O$]%Ɋ��u�x�@[��D��(F��c)⎠"�R�᧲GB>��p Εй���oU<9N��v����ɫ���4�8\)RH�>�!^���ua<q���jLf9bډs�G}���+�󅬁�i�/�x��G��Iq<��&M��p������`���5,2ﰼK��>���r��b#�����C���9��a��H��+�����SZR8����F�I3�h��%Z�Jk��]Rn�%j/�z�U�l԰�������˿��6�J� ��+��y��������Y�}l]3Px߅44��%Sᡭ����'qһ@�e�J��}��;����d�P�~��D��0�G�s+��_w��#J��۫!�Ly\��Ϗ�_n$���O�U���`%�L����b3�b�EF���Ʌ�h��$5����k�G���"��������Z14c�8V�@+�
�3D���1�P�`�-`��Қ�s:�m�?+pxZ�]Zi����c�Pȇ��M��
�)�Ƹ�cI�1���ߝU?�]�� �~4���|�~�������v�ůD~5��V6j˷گQy��pD��:	"�l���
<��3u(#!�'��R��}jt:V(&Ə�y/�Y)�|�au�R�j$5(�D��~|��0ܻsXS
���E>�K�@���Y&��r��F���7m% �"l��:&�$��(��H���f�\S��q@z����E�B������k�k�f���1��^�癬2�-lt[�)��oBٜ��/T_�]Q�0�@3/ӬNs�:�5��a���(�����=�"����d2v�Y�Y�[��@c7&��S*�񖮱���m.t3#��:�\�� j[:W�uGe�I�b*ZZ�Gul�����,�W�ʤHp��ho�a��/�˙Y���[�0�^��b������u)��vD����Rn����%�ԥo������K�o�9�/��
fI^OF�TE��e�
���"<�^�$��[j)�T\����0��|� {+~N�lS����,+P��[�+R*�c+?��LٝE�<��l�/�>�pZ�������g�oa��P�C@{N��t�I���.�̯�#�8���`0���u�fSm��]��"�,x�_"swç�������C��e�Bd.�'�z��7Z�j>7�� ^�2�H�X�2t�׸�������U��ط����H%+Y��������w�^�'�8������˙���R������c�e�BI��l��l��o�h��7Z�q����j��a�ܥ#��U�-�z�0�\���Á�c��Yx\�=����U'ˉ̚�ub��p����t����-
"�-_��Ԓ�j�A9����2NLRS
p��/�0iE��z�	���@�H�dڤ�#W�
�>��>�`aF����,<]>��pi����V�iz��rq�#@`�&���/�|�գ�4a�3r�f	E���ŗb�&뛗�T��Ԓ�Rx���1)�
`�^�L*H�w$F<�J�4Yi-�jzw����i��S6p��N��d�aJ�D���G/�/��=�����L�\2����R�냢���|�^.p�3פ|�6��;23�,�&]����2x�=ه�+Z�4L��+�c:בѽ�3W�rn���71��{+N�!r�@��E+��x�2O=n�H�ɏ���K]>���(z�w��]�4�ԢD��" �.t�>0��AV���f��YV��>&1�v�P���O��5�9j�'�R:ē���=r3��|%d��|ր�hY��A�Gc貔�,� ��g8��FМ��b��>/�S��v��s[,;����.D�����M{��<	�y�i/p�4��x�~7��d9�{Ϩz�	_����������|���h|#y��\���7�#�����Ӡ	�阅�A�~�X��A�X0��1�?�%pM���]I "�R;�S�إޅ�0�����F0�rqe���)RP�-ʉ%����R=�@����q
8V)5P�]�)H`7�(R���%��N��Sl����fh
)DDm��x��qs��z���*��\�)����a�4�y�2�`��%�j�4a׹��r�ue��eJߩx�:2�G������@L��b�R+e@��4k1}t'9͈%u�($��<�F�/�:�QM�M�NV�t7&���E]���	���"�&�o�S\N0���!7)��҆�V��lhD(�(M�GD6���3�N�Y�Nƀ, �V)�&�d���[z�'.xQ���z�)-��������Hنb����H��"�g4�� �F+��n�?�^��&3����wHJ�I��b���-��!��Fv�����#��Zֳzu�=��\�cW�M=O2%�*���[࿔���4T���.��>��P���*�V%8��j�t��U�R��?9\���5�z�^�����f��"�{Q�F��6���&��ZZ���D�B�;bcE6����u*O03WY2�M�!#��6w�����'�(h��A�� �)��{t��Z�[rx�֟�Z!p(��XD0���D����d�6$糖�K�A��Eݘp�qK륕�#^��o.K��c�?�������p��&E�lz��j*�j�;�(O,#� �^k�x3p����E�HL�='8���V�!l���d��AS���[!�h�2���J��XOIgt���v�����モ�N��+(�5n�vo�$2a������SRR�/���ș����zA��^����H���Pٷ0�!� L�(=S	X3)�����mދ�!��-��kDb��3��Wæ���/�B^�"k�\;�ހa���o�����)n{k5����%	�a'޹B�4a�K�;<�� [��ż��JȬ��&2���®!Ř�6���I�ST����d��������r	r'%\���%�]��v��>�k�X@��[�������?��G_S�<̨���uYw�)�r?�v���?Y�_
N�u�#�e�vPh�Nd�4;`�٪�6�-i{L��X;�,D �jV���{��
�)\�?� M�tX�ep�N��u���g���\:4���.��߶1&�W�B��o,&�^33MŸ@D/�KP�/!�l��n�T%[֣�cg?0�)�u�k�͠Bfk��A��篋Жm_�*���E]�j�_�R��b�uI��m�����m�^���#��2h��t�SoYk�AtOA���&'���p�\�R/��������'W*���܅�������mˈjz}�ج퉼}�ދP�@܍��&�L��)/~B�Z��g�*b�bdZ��&������B�0c1����rb}��a�� ���ƅ�*zx�"�hziJa{P",�V�L���# ��������`U-�Ǉx�~�N���JLN]��h�|���~-� `����)+�ZO,�W��S�k�D�?4׆������jF.�:�Ǧ�����?���x`�� �]5ŋ��F�
�/�`�L�bmAx��W�HhAF��T]6t`�:����q���p�\�r1:u�I�:`���ͺ� (���J8�2&1�X4%��t�!m���3�A�֏bkl�΃�G���Y 96�B����?�O�l������x����G̲r�
/_x1q8`���=Mז�o��3)���e���>��!�i�k�N��Aa��o�o�����Sǁ�jj+�(V�nbؼ$O�F����C4�עe�FGV�7���q�X��ݷE��E�R�аL]���G���`D���.��������[��ܬ�c�u��H�RrVU�8���{T+���5��]b�n���� l��a�`�y+9}d01��\������Q�?�?v��	���ʄ4ت���r�� ��>䯈���e�H�׸PI��%�2��]�CՒu>Jܤ��љ^ƖR����v>U`�|)�S�͐tD<"�vF4w��8m �"��@f�t83FKfq�����}�A��ɜWx1B\\�`��qE^Z���;㨐B��o��Mrcv�`���wb�?Xb�Od�=/���٩�x
�Q��RC�"k�o9�z@��v�����Ϛ�ۡc�Mȵ򥤮A������^&FIʰ��	����	��3��_̥O�Ǐ�2 �:���}�c���#`��"^��(������g��$�\2�R�32�B��r��\O$��}��5�zL�jUP�<a�f͆������4u<7���41�B�׺�Ѳ��J�����E$`�p�C�̺�R1����:X��
 �Ks��w]�'j�Q�=Vz&�GA9z8A^�Q�;IP����e`K;��B
R���2�8q��쌻k��vg���l�;k��x>�uO��6��6�eH��Йy�W<4�u�K����N癏X�BԛLWœiS$��!Z� ��M��k�o�U$��-o�����Q1'����"0U^5�}�.{�X�8���܀o��g�@ �ֲ�)R���	�ES�L���F�Z'�c��ԥq�0��.���޾�y8�s�P�&/�|�b�w"�;���B���cB�!�M��?�(�ۢk�34�	����x|?�xHpH��ћ�<h�C�\�O�`�Y������	?|ӡw}+�}��]c�d��L4�d�+2�
+�"�>O.��r�t�Sꂽ%��	���ˋVkѼ��H8EKggm}ȃ�nu�A�؝��l��`7����������C��`U����QS��S��,Is�'���@��-7 W0K�&<�F�'����@�c@u��o<�9L��Ǽ�i�[E�~H];�P�������J��F$�F>�/I,��(h��_��	 �\N����Es����m+46F6Sz�{��|�ho}�l�e�s�vK�lo���/��r�,�����Qi0�:��X��A�vu�fA�`>�p���Gd}����V~8m8)��鮜Ѽ�)>���8�Ub��OxV�=����xz�j�sCWD���)�$����yGe��w�V�N�� bOױ��0S��,�[i�-���~<�s�;��e�����\����w��Q2�r����
i�/ ����H�T��-i�w0��v�?p��E�B5��P3�3�Q���qw�P0�ð�������Aa�?pNB����IU+d}���At̴��m��A�*K��)�(f?�߂��سD����d,��/���>\զ0%͕1b�c��K~Y��ְ0���(�R��i�峂F��0�L�G�P6Å�d�~6�Dʁz�r0]�f��O1��_���1�Ԑ;'�kM�U<@s𤠬��l7uO\B���c}�+f���'�ȩ�o->됐�j	��f���~�wa3ۍ�1�$��F��e�����)���u��h�*:k�uC���>���\��(ֵnBT)RksMIUl���U��-k���~��Tg @����x��	�'�靖�5�QGע1�Ty��tso��p�t�67�����*��J?a�I��`,6���Y%Z�?��D���̓�����уg�|�35�U'~st����>���q�,�Hn�c�4E�Dx(�4�q���F����Q�?)����5���	�vhd�8�xӘ���-P=������]?{<mx<�&b�1�UͿ�F�M�.Q�o���ѤjN�څ�1��P�.�R>��W)�!�5C�pw�w������04P���f��A�����-Ơ�48�X\蜋�;dH��#i�э[8^{D$�	n�Y��l}nJ��{$1�a%Aس�y�
M�xޔ�#� ݿ����V�:��D�<F�ײ�����~#�~z��wX>*I<������U^����(��:���v�>�/��%�c~��ٓB�޽���mǙu{-�	7�|��9��i�%�]��c
��c"	j62`�q>v�:!g�B,WO�}���0H7!u]�@2�Q¢N��k�P�ߥ��#�-b�e�w^q����� ��^�'���6ڹ����zu�������REh�.xrI�f<= }��ޮ�3�-�~O��v6J�J	a�G��m0!RtN�5��<��ё�����O�0�%8m�ɒu��l�ݱI��ބɏ��o�UϨU�>@���j�\X�&L%%`��⌇�g.�yZ}��K����Yn�e��:���X�� #�Y�/x�B*:�uw��\�S����+��{1CY�3��r����O���.Ä�>إ9(�"�)bd�:{rfd��%	����ާ�Z��@��좝���Y9>�m&�	�6 ��lbT:T� ���?�5I8FȿX"IS�7D�{��?QV�vz�2����f�d��0��4�9�O�όeN��M7[���&�7�r���_ƶFm�Է�\�*���@�rQ��Ҙ`�D�5�햚��93%\x�S�Ǐ�Ծ�p����$��g�ݠW��v��iFO�At)>��7|��O
����2���{c�+g�p�J�3L��n�]�z@�>����-+Vr"�i�:���޹�n?'��җ�N�?��N7`)��LFd13,*�M3d5�^�aMtL>��.���XN��s�l0�`G`Ol�A[��{�-�F�9�=xJY���C� GV�p��8h/����^/�m�zB١-�j���O����J�E�A5�7`V6ycZ����%�ɔ>1,<ˠ���H�`*����}��CV)�A�d�e����pf�h"Ea�^1r�+�ʙ�ؑ
ʓԨ�^O:�����	 ��M>xrb��"��ƞ�v��<ܒ`y�4~]�aē�Mg_󴬀�iH��pq��;��ߐJҊ6��I2�䑩Q��c殜��o�"�	.%�ǧ��w�v���6�Mj4��d: �XQ�T
�Qͮ��Z'�j0!ɰ/m=���M��>B�M#�*$����=l۪��o�}��KnG msDIF0aAw�pI��l�]��6ˤڴB�j9�O�6�|�C��Wtt�}����E�a�=2@��9��A�"MԾ�� F�B!��$UV�IFt��l���i���L��.W�O�Wћ�^�?�R��sÃ��	���xg�\`�A}%r���H���0_!�ZEQ�H{���|�|��ޥ-E]�J&�LIƙL��x���:�[�P}� ]�<)W,턜!���ەW8���ĸ.�����>x�&�T3��^'�G!��t�S�I5�j�>��iÁ~��I�-��x�mP�cj-=7�C�&�pI���3�n@E�YT٥�-�ԕ�=%��x"ź+�ޚߏ�?�1Hf��>¿+g&��e	9ۅ��q�MA ��|����r1[�=&V�d�h����1�ɜ��BY��6���@�Zʿd�Uφ�2'&�ZF`ퟙW:�������R�a�^v*���ΔU��v<�O�9�Ш�ad����~��꾯�=N}��§'̋i,{h�>��P@iΉ-Ʈ�����{�	&���F��_�߂�G[�"��b�?ZFߪUe-�e�_�"���}1=R6{������V�����2�8�%fXe��f�q����`&&�/�4`e���%�}