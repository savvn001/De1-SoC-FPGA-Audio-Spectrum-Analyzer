-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ijs5TfsZyEdpun13qqfcxyPyaKUGaStZK0VCczrkvMjcbhp5Ioqmm2wt+deMM8xg3p1CMbZjrnCB
VWFOZDsr+6fyWivzGWFRZoCUgbqChktrtsmiZh+qNbZK2RJNQrDop7RH4idPF4BbpFm762CN57wF
B44VXxq2jUvG9lQKf93pF/1J0iGnkq8gouDO/LADlUjkoyFP0SEfrcEKxuOY1Ywq0wTrhkisnW7u
2weAup1WtGlKgrc94V4W+qNnZe1ZmkJCrdB5xIiYbAyOkeemOWgnvbxz3sTLUZsHAv23BSC8lucE
4eY9Pwhn3EAg0YV4eF6g6GNWqmIlWNGeYexdyQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3008)
`protect data_block
j5k3mKqnGKaInflA7siZv9J1ImgmwdrzidKmF+4zh7S4IamxTbZVdvKLhWaRMVBQhBkvEzqwx1D3
gsOLQ0g0EaqaoIRGe/UJWcEx6JKiSf0+h3WTc5Ywwci/W1KXTpOWS34+3RkBaLi8OmFpYPygNV3D
K8Ypj28s5iTZ+TlyXh4JYnvGtjZ1hM8TVcMbjOGCgv3bB8QW7gYFmSHVVpEstHm3Bqwj8zuytuz7
26Jpx9+Lo20hNVhd9ABU0KEAaaCnC9ftQ/VObbys9tYJBTeOLjdNbABJMrjq/VZvpowk/sD3oBtP
7+/qxslGK1IByFN6tVohNx6O/nnCr4pGtXwzR7cSTcNyM7nW2H0D1dJbq1OmEP4v9tutCtFeRsrL
y+UqioMrS06wAuv5iCR8fQ1vKYZiK2cCgAG7SsTOaOJx5UrWY6d3aEMw8y7j+wuZxBHFoaGc3X8K
FlBxdwyL+0h9kdRegEZbQgHINaDKzy6ToH1+eMTVKWa3g92tTe73BVjNGNFpLyH+BYb/Oln5zAZW
Vu+eR5I7myRPD8SD75gmsqntZP54OQar19wY8f25U8uxZvbM0157uMvWmVnjZDT5wY/navi9uYH7
X9mzDdMz/K738P9D5IW6diA1s1V9/mTgMT4mw5mU0GMDyfnV3f6G6939KDvGr9DB7J0ENwr1x+lM
IPua0gPNUhmbM2N//+Cbc87aq2RwMoyiX/Lf3vJFfPgFdGA/Uz0yLHHzWfpSnmT/d4ZbQsJCmWmB
mDsjswT6lxqqBWoDhUJeb1vsOuOVIn9lHz20gnLZU8+KyimcKNULg1992aR29+W2Oh7T013ysYxg
hPe+ThNcZFqXXmnRMnZC3FKwoPu8Dvc9geke78ZSz6ZffYkfwxse3JbRBczSU352g01vZg1WBSgG
9SO7BnKrdzOeMiwQTdyhr/t8Sm8JD0yjkyBUG0zbaV9EXewJW2IB4BT9+lXJiPnY29hb0wRbap1s
mfvtAh+LXIeMcRuW+3P+jprOPtRbBiZ+N+znrMSJ/3gvG7hzhE0ZvE8mZF2Q9CB7Axd5qNN9clQA
l8nWVaQYAsovzl1vb8kp+jGx1HEZaZFndRIYoA8PgEf6BGIAHukfql+TF6Tk5qdsxIfdaWumCEaG
BNJvLtY0UL1hZvaXUz2iLh1mOfz6X9/rC2wxfyo8XEc997m/SkC9DEgLOTogPkp5e0IvUH/CAhiA
Ex0VG6YJiXHc8ARxExvToc0O3c61mORDRYJxhjJqP4zqICspAf3IVyYVFavceEgMo9nk3CGw/KPq
DcXVJx2lxGLtoqXGFkZTUcMtZi8HBDxPeibelqgjyQiP5Jbqgtuy/O7jhPWs6RYrPNTGYXq5HCd7
5u+9HWU1aIbhfREOGOyesR5eUyjM5p7faUD3aAVWT31fzHpgIhqMMOLtKF++4Eny/zX5Cec4iOwj
65ZWPSp8/A4E/KZDV8WU0Zc/PsjkAEiPEpadrjdDK3bYSlagn2Tt6faQUtBRNbAQAJXcEJ//ju4D
c5IJ+NuHaz9O8AKTJZmAakrRmt45FmwRq5gD/mwyGan53pDDOqV/pTGQnRvYbVAdYWWdSQkD3kF2
3jtxhJYLX8Vb1qif+9EkhltkLQviUYu7zmGymhlBVHPYP5quVfHPOMF/jzUJ4jyVNKxDTlBp6oCh
rTE4h3FNFpWe36ZwJRx6yj3lRPQAitLmiaYAEftZ8HMb1gXRxqGM3kzo1Wmz+j6hxbIyJLOMMwwd
CoJaNgpHGMnAMjvpgw+CXikXeds+t0aDl9VWvjFhBx1Yms48yGOy3VE1kRTmcOPjd0nDFYU8f6MT
9NzI20DlXDMol0xva5SOU7RHOKUln2Ff1tqYml/dI5Ea/+MWnWuhNQABbqdaw8xXdEjk8qDQJiJy
lL16utBJ2iI5qQhQRYNMC7Yo1tqj6GZ1Xl1Tgvqiinv75FdKKn76t9+EPwA9ecxUtnNCf8vvuR30
o/YX0gRUwAKpMn1Bodo6bwUKXzaGgAIhtW0NQI3Ts/vlafk60SpdxM8v/thGKPTW4DUQ+x3cO+g3
RBuxJERsG5K6PobGbKmjZDUDc05EfKKPdLkt9kyD00ru1+LjPoMU30hmU79ZkUzOCtBIVHaS9FUW
H9q2UC0lVF7AX3s35XvRG08Mt9QymrJ/S7inyDITtMDt8if3igoBiMKf2z6uKMNyiXMwPPiUFP5A
BPj58dTbjYh0dO/XpLCzsNSC5QjGQ96Cjw8RNtRwjLnetyE01c5RyoT1HnlOmK0bAyaNuYYMMPD2
GGnWYa4lgPS8xIZ9uCH14MPIexgs0WF1l3vJ+H1lH2B9tigD21/KLZrFPm76LwLoCh+LzNNyNGI4
HONLh1IaClBQzLrhD6sYsQw2eu2WL5UrGa9UIgkgaMGRgWOdfjnOOlp0yrWuqjQJmLF3YhCjNTcY
RWuN9TI6tgYsv7BpN/SLL6jHKhnEy+BmSjuzKHBXGDpxnw1yw3ekuWllI7sRvU+UM5Tiiyiw5twN
bF1YiLSpgeU8CSs1IsrdyHtyhLQ+n+1ha4Rs8FSsHGMu5T5/0eFTY+7WmlwzlRPkbfViyzvHidVQ
6o2vaqeEBpSFlXJD4og+H3Bvuzo/oMR5/AFyUCZvuLVIFvTtcnykSsrqKa9Nz0xTM/7S4ZmVqUSr
TYklvcB5ag1wtlCMg/Ek57nO6PLDtv3bjN+u0fI0fJBRcxFcqeC7XodSltJFOjFBnc69cvQLcn2N
Ghwygm7DVPBihUgQQ2hOLYlMXC/A9tE8sWtvL/pkHBEwANQ7P3sad40ugt2YvJGbVeCFpPoTd9MS
Ocm/xsE7+5PEKLvmGvnkarn+U4BIL3ZOagOvV0Z7QsMrJlCOioWWX2Thj3bP5DNLkkbLVaKiryEs
t76Ic2Z32+r25PPXuuZNaFc5h5JGQB7EwOI6DIYO+Q6vIAvDa+4+ziMIYDCNBViLUzjwO8tEbr7Y
ysaw4ChY61bQhaqBX2e0DOrFYtsd3xn/YANC+dAOhGIMGAA09ff257zNDDRLDqPLx6T3RUKxrYPE
2c2CneoJZK7ZVBJZ8sN7CvG1bObybuTTC+fu37MxMrAZcXJXEjLymtC9HNYENmRdgL6PVvU7i45H
r/AMLHCOhYUGWlG6cnW9ydUFRHCluuqT0i3rLLLr2IwLUf+4xQH59cyRvEK7eAcbvQ9jhLK+VbQf
XtUPzPecX8xvhsE63OH9U1rGpQVbi21EjA5POa097YqupHsSKqGz3mUUiU4v635NsXTwiGX02mdp
EMOg9253qt3DN0K3HZW24X9K2pFFQmlDWdFG5H4txHlq9tlOjs9ujR/30qaccnzsTQBY1VHZLwC5
oqhq9AkAbZssaSa9hVDqWXJeRUjjiroStgUtxNCiGIuAtI4WclP4njLqe05tDKa9Ms189dMQGVKa
fT7+cvA3JYRnfNPZwhZG9cTd1PzHjcHkb1ZkFiZIx+CrroR4oDRVd3SzkjKn3JQ4cyhGbtGdSiqh
winjBT2+zNxK4n2B6g5oZFuhhlcfPq7apDD+lPi2h3Z9fdRPUeKrpyoBw3fcx8p0nsnv/tWfobq2
SO/pdSw2QHBrgzWOse4WsD8RuSk6JK1gRaUuB7YosdJUZaBbRhsiHZ+w5odlcU8Udrnil5Zwrl13
G2vYSZP4hCjTMMTJ8sFYpaNfRpcfAlslz0eSQ9J+43AEKUK8oz5XW7h5chnXED1rewbfQoN11rbF
qVn5javzoLDpO+u4BEtzQ73QXS55YVtUPIutUiBpNT8cfPNxqYlogyKwor3fXmtlK5v60n6SaPvP
WxBeiyyZ1THnccRHrRLqiudf2JutZ7+rUiyA6OhLsj9hYTpfiHu81ZXro3XmC1rOJMUYxhNM2zgr
kKLAVKHupU0za2PCfOmHF0AUeU3aUJWL6gEmupc00NF0j6i9KcoHLac2slclPWPR4hrbTkQpy4/B
RWBjL5Ut0cz/179khgyzxCGbY2YyLZ386sm5JasPwP+5wscd/n5pjiOac/4=
`protect end_protected
