��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�:6�E^'�2J�d���S�[`���G�T�H�<[��!�4k��ﶜ�rʞ �n��e��Bt�0
(�i�M�M�l���u�DT���'����TK�CC���Z
d�CW�.N����c�+T�w�m�m��J�7�	����	7
�P�n�yɠ�~�'cM(���d��b�;kj��	���TޤԱ(�
��ѓS9k� ���ۓ��f�����W`?S���F���=��N@����$���֯*@�Q�]���F�J�_��`���g<����$�S�qk��'
*f �x8zz&T��n1Y���_���aF>fY7��� ���P֎e���*O6���ʎ~,�@�!�q�Ix�n�w��l�rX�{��9E0�;(u�}��YC���|<��]U{�L|���Z���բ�|��Ũ��V3KW�%�TI.��w=�X��aѣ���m�%X�I�N�|�����K� �!�$�I$zʣ�k.'�g�m�7�׎9%�#��/JN-$R��-����^ݩ��� lt�
���P�/X��m�FE�� �Ʃ_�]�_�K��gh��|����?�mM�
�C�	_y������M�OT�)��o-P����^_N����,x(�-�V"0��J-/�̴���w �����q�ߔQ4꥽]����fݭ鰺0�F�~|�q2��l��%W�⟻�#�*���g*��e�n�SLE*�/���H:�}�7[_�5WƲ��+ư�	2{�=�_�?��~�b^����7��|zjN���5{�f+K�n��RRՑ7`�230;0H�s��e�Xя 3����5,(�q2*�gD���Rl��
���e���y��@�KR�����K�����-��M���#)��,�B?���Y��T�AH�&iF������z&�g�l?���/�.P��3��n���w�#3���X`� ��͈5Ҥ�2������Ҏ��ܹp�8��Vo�k�Ϲ�Z��M����F��>@Ü��(��E�V�f�l�(��hkXaC����az���j�����"Q�ӖKa��W�G�a��b�L�����^h�Vrv���܋X��E<�[����q �����F۽�.��4�˒�K��x��8�W�9c�k��by&x[��CjߣU���P87&�rȺ��tW%�3])�+����e�yn�tNQ��Nx0�˜=6 ���1WI���*�,�4�v��G\)�kz�N���G�}ʘ6*ױ}+!Ty���/�-Ɠ1��Ui��-1�ݳ���:B��@*0?�TRv��Wp��<s+�d�Na)A���3�DATpZ�X��l����� q�����b��A�����_��^~���q_���M�ö�4�t j=*Se��y�EC�f�P�=* �u�[������,�}r��U����0�Bm����4�M!�S� '��?4t���y�~6n�
r͠��`'�N��l����z�W �v�m�@�"�Fp����s����,�Y�; ���叿x|���`��Q2A*����v�&�3���8NCoǃ^g�PY/Z���$X�o�p�E"7ͧ򻓁Gȏm+>�1R3���'}����"����j�'�	K����`��,I��n�u-O�#h�;�O�S���/��6f�}�e0&�|R�p%����%)TB�3h�%d3�c��RZ{����f	���((<���L�U��hKrGO��q8�0�o:�1_@rE[�V����B�ͪPҦMlh�^�j'�_���9{��q֭�[|X"d��5����/V�I���y��^��ӢƠ�TU��!�	�uRx�S����Enm�Bښ����W)gߔ3X#�����T���N8��?��;X#�l�!���(D�]�s�)�a��]�iʢp /(������4�� V)���;C=$��t�or߰S�hBlǴ�õ~rD�1��\iiesyu�t���=�9rP�6D[�c�������E�����G�8g�����l�^HZ�2����j��Z���%��6]���W�[Q��0��������[�h����DΛz\jg���t�!����E�e,?�;Y��ih\ ��dv^����$K	4-@m�l+Ior���Jg�@T�c�`�i�`!$я�n�Ln�j��L��7��b���}�k�rw'� �ѥT�g-ߍ��� yJ(�fe-BY}��";Q��#t^_|k�g=��]+��~@����r�S^���{ʚ�S>��z�
y���dZE��[_�:�a�i�連�k)&~�"�M�{O���ei�p� ����j^�62�*�	�B�[a�Ez��ο������8'|\+�ǘ��������z���~�蝈L���{�.4����>j��P�2�P��S�2���F׎�a��R�
���FI�i<���2���&�2�5D��4ϡ[%��]zP�%Wu���k6
���X�|@�
�L*�I��u�{a�(�u
M%��������[��-��f�N�*�ǻX(�s��� ��]Ϲ��k�S��	�1�?3�z+��1x�d�;G�ĤQN�߯+z���RL���I:� y���n�ծ\�N�Wa�7��.��@�;k�Df`R#k?�/=�y�}&���r%��|8E�"�23��T�@Ю@R��?.��ƕ9���m#��Z����x`�t�&���>��D�=�Uݝ���f4F��b
:�n�O�w�:�,.ϣ쬥�0L��U`��y���ɟ ��-[WKkF�[a��F�E��j!9�p�C)�)R0U��7��t��9�h��=׊P�P�1T�����1z#���tm��6�\�U;��?�aX��O����$��Z�0��L5럾(�����!�oH,�:����_#�<��&�n���W�@%A^���gp�*�d�H�hj�ֲKu�#z�j# ��9���f�-��6삫��wT�F�������O����~�hN�	�i��}/Q�I�t�|�C�;�����O�1c�|	��!+�����t �Zsa�/�
r=�� )��z���H.:'o����`�}ή��K0�G�?�|�9�J�앥������Q���*[>�W0�̛��q��Y񠽏�G%E�c 6�D�lr��݆�?���aЛ��4gЖ8��ɬhn���,/W6+��pfk��-(���	��	J��j�"�d��hV���C�3J�nN�H��ܚW"�#}��f�C6zs>݁�_1�L �q�j8�k�u��=Q�c�)e�6� �?�HP��zã8���َz=K�;m��B��e��c�=�	��4u�.�am����(s���M�s��ӆ(>H�췱n��<�'��8ƨf!�=(Z�U�1��Ȗj���	8�@��Qh��M*��>�:�O��K^���4���A�y���:Ћڶ��u�
�{7�s$Ѫ�L���C�I@,	mct�dϘ��&φIΐ�	Ψ��Vq���M�1�Iۘ��8��kf��je0�$����V1��nFd
tg����FN9~4��d�0� j#oƢ�"ϭORI��Z����ϊ�ka�~��JNv�L����̛^a���&`�ǵ���H�RӚj4.	���H�����hΉ�+������i�7���[W+���M��GX�P�R�T�hK�K]���/�Tt,b?;Ρ%��nUu����$p�	xu�&K�Hz?�Q!I�DH��&F*XӠ����{qN���˻��?j_(��Z�j�6�v�/��B"�Ns��]Uð{`�����bq���Z��W(��a�.̻4{7�b���K�̘$��x4���!1�*��E�3R蘄�	R��tS(��T�A9㜴��e�_�c(*?6? �����K���AO�A��1�R�������~��)��6���#C'�R��v���쭻x�Q�����Q��z�l{e�2G��Lε�85"ݪX��x�.�WR�z�г'��������e]��@�z�Gנ(.~�V�*ᓊ�H�t��غ�XΣ�o!��b�U���xH8[m��y%oއ
?��r�v� /�� �6 ��%�r r�By4K3��+���Q��C����cJ[��B���"f;	��Xkcb���7��N��0��4��x�0��7�єO<}5$��zJ0;wBE(q1uOƍV�,Ǝ��_�>��� |�C�J'�t�	@���?� ����[>$��,�&\:�^]{�EF�D����N�x!,�5c���_Jkt��U�@ĺ��x����w�_XU?Z�l/�iÈW�MP��KŐ�԰���y�\s�)h��{�=�m��ɂҰ�������	�پ��}��iY�ӫն˟KtME �>�o��=�9u�E��.n{
�y��ym��W!Ԣ�:4grЉ�Is��4��Ŕ!�(73m�X9���~`Y�tV~��dn�U���C��#�����g�����"�tm[�]��m����J�!Oy,��Y(�0J�-LJr��D���(Y�CV�b�81�M]x�{]�2п��6��j��l�=��lp�E������ZU��l����\b|I����%�s���3N��m��!�q}����>����n$0H�jq�-=U;�����2�M�(�4��?�ph�9��%~NX2aw#'*Q�6�[Z��>K-\�#�[��$H�.|�b�\�JY�����)�G���^kO��,����KW�2�n+0����q^��M��]LV?���?�����h��Bõ��2�+)�Ɏ>$�f����Ⱦ8���:2���*S���+�� ;�}��X��܋x�D��Tz=�z�L� (�|����P(�����k�g���ܗ���}H|�����  Sɉ�/^0cm�o�Z_\K�D(}�:<��o<[͒�Z�����U�	d��~�R���nF~;�s�1��.}��}|%R�]�&F����α!I�A2X��!v�:�Ye�N#
��f�N������=������0�]-�Ϋ�J���.���3����Jx:�i6F4rt�K���w=�f���CdAխ�"̀;�O���z�O�QD�;#a���x��l��pw�0xZ���U���!���~�vQ� ��Q+�h�b {�F��V��3��ɇ��o ޑMb��:(`���?uD��K�#t��*//���R��@���N;Q�҅���ws����t��@
�wCvH�~?U'Utj����g}7�p�V�@�@�r���*���#H�����n�'+7��8�Ţ��%yiׯ%3h��X-l�,�n����cw�2+�K��7ʓ�p���\�xkۯ눣/�ֱ\}�.�{���S����5���D��8pe���F���tm���k&�V�z`c��WxtX�Us�C!Ϝi��?W��8�4.���!����k��i��\��²nh�6.�[�v�)O~(���%�i�����;�g?M�S���xd�DÏ���4%O=J����)�־T,ܿ
{��8�?�/9iY��<��a����l���Wy8|<p0~�`N��#	i�IDg[�r�Y��LL?e����3���AS�a����.\�A'�h����9�:!��ݬ��� CNm�I�{����sY,^�����w����B��M#i�A�?�=�J�$�8�J&[������K`�0jf���s |q3O������E\�f[��$�֪�B�ݱ�0�b��.�gHC��΀x}��"�L��6�en�۲Ii��4"���6D��d�X�+��aE�&�Əo��Z*�� �p ~]��Ѡp����W0"G��&������9C��40��%_��3xj���nު���y�\bwN2��2,�x���5�V�%�_QѹO�2%d(9�$���X���؜b���鄩��V*"?���������۰��ZC����j�i8q����-g��@��@3����[Ep�_h���Eh�Sg�h�tA�A�S9>�.~Q��`p>E�Ka f�GLdm835��;¶�\��:�Xd<�4UڃX:|-�L�=(r�N�4��[E���W����(� -r{�����Ӆ:^�����ė;��m�%-`g�'P��\ʖX�3���e����L��2q|*��.'{���CN����j���M��l�R��s�0D����N�X�vi�k��_��-dw24��mv�̞��Y��X�Z@�w)� A��Ҩ��;���hd5�GX��up8�%u�,�&g{��D;R�N�r��f�W6\��#�E�rm�r9���~}����F_h��)���W�ft�`+��&�/]�h��hj��G.,�) &I	�*�ÃZ �_XG��[���m�����%ծ8հ�L�9��ET��8>ā��~cSg�W/���锦�ځ؏X�kA�K�����by6�-0�r�Uh�	�0���5��j���2T��z���&���B�<�r�om��1���Y�w�N�:|�j�uaJi�FS���R:S=��C�e"���zS�1���#0�Ԡ56k^O�Qv�4�C����^����C+�v�9���޳9M�8j��UTj��7> &�}~a��
i��{;�v�������R#Y�DQ����~���s�!�?�M|��V�m�]����r/{�b�}�C.H�$�W�'H��(�N�N�h9+{`��uH���N��	��@�|�H�?Qt}�"�ޱ�
 :�xW}���95���gms[�c�i1��oN����M.R�X�q6�φ�"�Y$��v�dbT��H�a,d{�].s�Lp�ggt̎uY���]���&�����MY)�C����g�Xie,���P4t⎉c����? @*c��x�r��T����}��5
�C[/���l�A[=v��n����d�C�Awzb�|WZ�B��#��Ԣ����� uh�:�����x�)N��˩�>���؃�����Nj����bѽ[�RA{W��P̶(���? ����l�6��!S{�@I��L�F��?S3Q�� [-~H+�~��������� =>�&I( 3���6�}�>2����3�Qn�q���4ԫr��_>��	� �u�1|�H��q�ׄE4wv6�r*<䠰=��
|���\0�+	��8q�#V@WڥD���GdpN� 
�|aەK����@�K�+W$}ʗEd>��NL�4Uu�]L����o_���
��*~�>;j��]j9�6�8Y�i�4�WL��I/�]�
_ՑR���q>/�9������_e'��IhKb�
�V4��*Wg�,���n~v4n�p �x�0$<ǣ�ͼ<�K����Ai��D��h��C-a C{����kM�N�qZrKi{90�S&B�j�Y]��L=�v��G���?�3L������u�G M���&~�:����mZ���J�(��n����l��L��iJ��o���e"=�
:�ˍ�.T'8���0��x��`3�hhL�x%��frPOFF`\B�r�č��0$�Rf�E�ɏ�AE_��\������r��j��Rӝޅ
݃h���	����ɽ�6�W���KDU�û�t�H�<�&>�1<\&���Z�$0�0
�S1����\A��M���H���&|��-qT�����JLW%b��v�p��Q���,2��;����������G ��lӋC-�[F�}��yP���m�p*�Ԗ[Ribh�.�'�&wC{����M��d2� 6/Fh��י�"�Y�sF�pU0֚���%V#Od� DL�Q8�ka�蝘�2@I9��>�����	[.Ы��Q^x:��up��j�mP����ǋ�Ҭb��K�~����6C�q��I���^�t)��lE����v��mm��k�.!�i�����p(�|����ql���ځ X �n|8n4�@���&Y ڤ�C��w�<B��#b�>�+��:_z'�R??�jUu_j�Y�t�9���[����[�B�ؗ�<a��7�s�6["h��ʲ=�tpM�^�O'J3%��r�ҟ���1ⳗ"�N����$�ʆ�r��@T�hA���W�� �ʹ�4a�>S����\�sE蘙!��¢#���R�"F�*�_B���jh����?!m�ۚ��`��[��y�R��yIJ��/|W�5�Y�܌���Jp� d���:�is��M�1-�Y�6����U�bŚ[: q�ꍆ~��8�t��6���`ճ����f�l�⬔�uUO�_F$��[��&��=���+���fK�(��Z��?Ǫ��d�R��?����Li���A�4d&��a���0)��<n3�wn�
z�S�����/U(��k�@~�[����X��m�k$�{P,���:�zC�8�Q5�Kx�Z����Y��'�TZ,����?Q�i��y�E閟��pհ��)'���4�E�79+�)ls�Ѹ���3��iTӔQ�� wB�J�?�k�O�q �y�)��XS�Zܯ͊]x�5=��r�}� x*�/
+���j���S�N�+)W�p��ګ9s�ԡ7/
ڵ����l;�$���<&�Sb4SI.D�~:��H�n�,O�j/�`�~�~�׮W7 Tg�BX�|% �ŉB�t:�y��!�1s`�7��������&p��3�9 Ѥ~�n��90t����l��c�;��1w������4���M	 m��#|���_(J�i.l�z_�����|X�=xm�=IQ�cX
,D<i�?O������<��E�R��&�-�;��x�h�ޤ�	�l�L��1FJ�1��,v#��`L����oS�d�N�.,�X�8H��:>ܘM�}�a�Ru�H�*��v�X��] �rk�QNm(-�7Y�d���fGM2Z�LOlS;_����5�Y5A�@T�� (JS�{PS�f̵���輛C{L&,�H���K~P)&�H��V�h���"v��\"F��oe+��6� s� d���#T_�%��'�$�ؐg�V�xޅ�iխs{ŷr�5��m�u�fú�'R�:^	1�վ���F�.޹M��s��T���X�D%�J�LO�4����pOP,S�i���a����![��?O����R���t�#Q(<(���-Di��'����SKxeW/
��"'�cNeIb�eh�{�g��B�p�h�"����)�tO\�d��	T�L�g�����y8 )��h�ٸ���%4}��9��r�	�	�Ԩd��q���E���D�Qf���>���AMY܀��n�ԃ])ʂ���$jXw�J�6��~2�Y��)z*Y�������h�ח�ӗ>E0�w���^�4'6�a�JIL~���x;d}"|'r�@_�S��P�����U��)���j=�.H%��p�)���|�Ĺ^��D�A6Y齆�	�n��Ђ���NT��B�S�5�<+��L Eb}|� J �_ӭgϏ�T�>Mk�}��G*B;{�}����.���/PK�HD?���h�{�s���.��گ�.�a?bט����#��x}�x��s��ț�sKl�$��Y�" ��_'h�Y��ܲ ��o���4��)}f����/�1���ޯ׼�Z\z�m�&�5kj�]�	�f�`��XZ���нB�?�l�),)�5]��UJ�U|}��&����A{�Є�r d�P:6����R9��-P>�_��a3��`<����K���e�'�#����� Z�+*r?�l�fz5џ ��*�F���`y~'i�v��7̐FE���%N��Y?�_� ��(��,�D������`�80Ł&��X�J�c@h}ä�>��yӕ�O�"���J�߃$�1�G�س�r���F���V?4E�g�$�Wd�� ��1�Q�$�@���#޻��߹}7���(y�Ms;�Y����Dӷ�Э�O��)������;�J�\���HG�:1�G+yC��-�=�GJ^���,G��¢�`�@y��h�9��l���J�\��8�������/����9�à]�,� 딫�e7�٤�X�t���蓛Xdq1V{��K��k��慩�yN*����y�Hl��7EmFZ��I/)B&Z� ]
�A��Q�2�eV4��_�&��q�xab��}
LԜ�K�!ťO�nfD?,�Q'�iO�%�N"X�!S�R���.j-�Y�(^��<��(ȶ�yʸh������T�K��E�!�S]�W	O���s���y�3�E��)�0T*��抔8�o߻���/��[�HG���8Dt_��.������D)*\P`��x$YP[�1Ww��+�?��~�!2���\�ǁ#���}�Ap���~�	� 5>��m�g�������*Ubׅ&�A� f^���	\��x�u��D�[�n�7齈f
�j�ҷu��ec3��Qm�)�X�f�󘖄� �0�w���6"/��GaR�Kp"�z6�/�lƉr{(�!C�݉O	뻔�>wq_��SZu{T�2`�D��&�%���v&b�RI	SΔ!��^��4A�۲��������!G����i��*79�P���rb,sY�2Ļ@��$��M��>�bRbٽ�HY��{���ͫ���Ǿ�wX����+���	��힢�����\ $i�X�D?8�*P�nK�`
����b� ,q	�%GQD;�h�)��^���/��ea��BV?�I.�@�9�APs��c�\�wApθ��`�:T��Mڏ z��s2�h���bä����m�g�X�n��7��/�e��_�p�5t��Q�4k��!�E��<k����H��l<��K{D��+�=�#�,���{�o݁F�򋒝lܵD�X]�B0�]r<s�hz)u�����'�z,!]=:�����t��O��-X�54!������RebE�6�z]D(x!d�Q=��D�(�ot�9E�G��dotI^Z� ��-sh�:��ݷIK썔�/�����!��>��,�e<H�O�[�66�qyޅ��NL7t����TR��M5�����sލ�n�L�͹d�1�p���~��R̓�?/��j����ǚiy���6��h���x�E��Ժ�W���[�R\q��9IMZ�9�����-�G�^��
��+�Jb� ���N�Z�N��٥�;���.���)~��/��5<m���O�ntN�B�[J���`�O<H�]�%E~�������JJH`1���-l+�P�8��d�H�M-�=�9��(��GT���bGWwBe�:���!m���zc8�$+�ZM7w���IA?1��nõU}�ɧ��h��W��N�1�(`$�inNe�~�;�-{؝X�}:�@�<��c���56Q?y�@}�|f/B:�3t�c����u�`q5�(��S�6z$S�>��<�3؝�;�ښ���M�t$���z�/�$�c�?[E	���7#(�3m�ǭ��|;����}�x�`����v%h�]��NVYS3�j�]���kzN4򐵀%;{?�S��'y�5�?%��rU+�5h\�*9�. ��mBV����~JoE�4�� %��c��GQP��)[�7%�����]��5�����TM�l�Tq@��R487�
�F�#J,�u�����[̙$��m"Xf]S����.���$N�=�Fpz�u]���x���)�`!ok��5��p��ٳ�M����U���?�'ˀF/)ye��Q�ئun�Tr&�1`gFaW�r��(����̜�~i��1W�������2<az_�X�6D��lF�*�.ff�'�+�+��h�u���w�	!�.I�Z%�|�
�2�ޢ�	�O�4	#w�̷�IR����9�UE\�N����,h�p�l�(�'t�����w�l�+�������p`'+�F�,
b��X�+�)�� ����§>UaRT�PY��ẏ�30�!'���K�g��f�H\�/�e]�Y+#B�b�?�:���<�U�L[7�X/+�CG�ŏ_A$�����T�y�����f�O�`���.,�� ۭ����TV���±�μa�����.>H��6Va�c;U���Aӕga��y�:�f3����B;G�ț~�W��wM���oK7{��tR�0�^�E����;���v- �i]ڲ��D�CHD�r}K}7�գ��\�g
�{�34}�ӽ�ny�E%!TE��N�Y�����(tvA�r�����8'%��x�B��ο�03��oL��n�����,d��=��/ʙ�H�vS=W4:�/��h𮆪'�����Ѝ�i%Z����]�JY��-�0�#��W[#�;4)�gB��|����h�hp-GJد:E`�3fEm46)iq#����VgkfÅ$��/3�ۓ(^rE��{�J���Q�����S�h�c�W}�h�Y�a��/�?��H�~�d�=�1c[��`�0�YdF�22�Q�Q+d��c˻�HE�`�"*6�Rw5KYB��S���>�S��/�,Y{�����0yyk�J����Z>���V椿�a��`�^Ӌ�\y�L1>iQ:�R���Z��ٓFͫx�`�HG��M
� U��)��7��!�]�mT���&1�1��b���V���U��IPt��\�Z�O�� ��+gP'�q10�ʿ�b*w�2^>=��*��pBP5���m��,�]�bۣO��=���bo6㧂�TG�v%5@�w�$�~8F��/�Y,��t�eh�ʼ2 ��u��y(��h�ል����v ��g8m$�}�8{^�sG�����W��;�2cf%>6I6�d�Dz��2 s���&T�-��/�B\`qk�Ҕk˜�i��"��%��OlKz\hE��\%S�a�v���x�(x �@/�C�;*�v�L̀`�ex[�����G.�������ٞV�H¢Cp Ő ܰ�N��5v_+Ƣ#�13�����<��y�i�$ks��X� wv�\�f�n$y�,E%�EjߖO��!4���������ݨ��k�R5�4�Źc}!9��pDE�BV�2�-!��ik��8a�*l���UUW������Q*I�A=��n�N�L���T��ȿ�F�N���*��M_�ן�"[�dz�B��2~Z���U��k
��X ��_���B������o�έ^xGk�"�b�~�\i�@C!��4]��;����>�u{2�;`UP�s��v��*t�s�����ڱ�o�<�Z�S��ӹ+�4��ܥ�E[��]�#`�MP,��I��벡\R�nl�*��$'�H��+��[+��)�/��X�d��%�������_�A���ϸ�s4��FZ �z�Z�D�R��>۳��S���q�H�)$�C����@6���)�[�sL�ѽ�]l�L�AcSA�(�d;Xܧj��Vr4�&�\d�L?\�[��F1�&3bڽ�ݲ�Y�|g�;��燝)J�1���� �^F�m�h뼸�c���l��ª�9�	"#������?�􂬥P�W�kPe��,�����8L��u��r7:4��O��ؒ���YKjr��1�#�#jZ~$�-c�[�[]ޘv5Thg�+R�&�II=\n��"u ӯc��|�-�4��L����UtTRF��I{g��a���ny�D�hW!�/z ��dn�k*a1�s��ؤk�.�����^�H����8�2����[��(��D��KF�=/�:��i�s�ЀwLF�vv��M���N��94�!,RO3W����%��+%��q&w鳍gbû�7����ec�%Db�6
�I�z���/� Ac�ρ���Yɛ��Ž�(�WNሄ��^TSm�%0����q��q����)��#�SVؑ�����_J�=�1�$�y�nm����#��miF_��>�-_�V��8���h���PXZ!�>�B�<��!j)��v���A��IurN�{6C}Ew+��4���l�G���6�B��2���	�N>(\���_�Chh�^L��i�	��?'%l��y	��.�ф��Z�g�|*l��(��t�����v�,)8 �
�s�y�c�R��j |@3� ܌>\�ȣܦ��V���+Mzq�+.��7�e�5c�Q����n��B8��ǴX�&,G/����=��#H�l�*�Ζ�Z�qf;�!ط-f4[q���v=M5��]&���`�B��mQ<���¿Ǒ���?�ʳ���o�s_+/,%�6�dnY����u�S)Ƹ��,�m=�ͱ�b��'��s��pԱ�����J��EN�L�� xo��5��0~���� �>EЃ�E z��F�#�wc�V�#�Ty1&,�(W��{�6Jɯ>Vc�$0�� ί�<@�N�Ñ��5Z���loAT�潯,~X�X����n�X�-b�dn���\����M_����Z
� �Xi�l'�?�b��A�����T?�)،�Xd��� c��� ��t6�2�p��pNKS谀!=��w)<`i<a��I�gC�/ƿ5���X�M�w�MC	CF�c�*�[M~M�_��`�NB��y�i�	di�18�~Q��
��˾�tcR�\Y4n����d��<�p�����K�P�)�і���O���Wd�0U3fR3��A��h�x��~�}|RM��v��8�ߟ��y���7!��o�Aù0Fߋ �tS9�j�)tr~t��U"�zs]�69@�{�=w���|��������M+׻އE�5I9Ƃ�ǳ�!Ɋ�4�)��>-�5H8��}�~W�9�߿��݈�$�X�S�?E��.�vM����Q'
Áp��+jex��~?�v���EIVz	�t>2VL�a�� �.�]��.����\C	wv;��ý5��1G�	��r?�-���:'�*:���S��0���n�x�M��p��P4Ⳁ����=�S!>%��R���� ꁶc`8�n%�3�0��u��%�h�59�6��<.K�U.��,����y�uh�[�������YR7����޿Q
��4ry��<h��K�]0��T��a��t"�G�8����e�dCtp����T��MB�S0�jPz�?�YeT.��"D(���3���*��sY�HP�CZmn	��Ͳњ� R��&P��k<��GZ��Z��6>�ڛ�t���=���嚽�s��+L�����4x/u0��ld���LA{Iu���C%���d�.��;b�ݠ��L���V�F�Iʞ�C}�i��Icg|텙5���i��L��������6z��@���0܎Dz��<�x�sWlڬ�DH������H�Ѕ>�?��F�g�\#>Uk�Aa�rfB�����������<�Z��.\Ǟ{�>�6��q#;��+v�I�-���)��H�nCYY�Z�uFC��ΪiҌ¼p"�����pa̬����O�0o���>Qͫ����^uk���R�x�L��-�Ozfr�~��W��OA/�꼨�k��a���Ȗ�/����Ę���j�i��D��+7]�5:���"�P:�����9f`j?Qv�W �L�:��@S��2�*g��k.�!n#-!x�&�]A,ñ<�H�$t�����,z���D�_-�@|Y�NR��S�v�]8އz6���dz��L�p�{Bz�}���Vّ���r4�D�|&��8�E}�.�uF��cV�?m��:NuS���>�$0���g�wH�Zf�I��ߑ�`��+�2�c8!j;]��{3���t�ɹI��G���a��B��|� ��w�WL;$�pX-Y�$W ˕R����\�7
��[l�	Hn�i>�G�uG������ǫ�dI��Q"z^�t�J��<����������/4|�aFD����|��T=�}5�ku(�<���I)<.Pqj����Nn�"l����8�f�^S�ov*KCd�?N	���Q�_��Э?/�,���U�`��I��ᱲ���d_hxR>~�9[���)�-Ǟ������Z�����j��c�Z4�)7��!�_+�+�D�����|���舮�[3_��Q'-�ڸW�tWr1n�âE��0��[k`����-x�d����;�9���-�����|�ʇꪦa�Vײ�(cKd�cho��bM1}<v�!~`Ra �#&`�'�~��QÙM��D�9zT�w��������ɜ�uC��-�s�1������,ڑ�/��T�'�b�~��R	�	J������qi��춟�{��"�K�8���SɈt!>����-2�����-����_�E���d�����A�&l���g����a~��2�:R�|#"Sց�@4���A�ϡc u��y*s�W�E�^�� �m���8�wn�z�g�0f=����3	�D�ܗ�^�%�ϸ!�̅K�$�k�P2���%�;��l��͇L�NM�$7��T�����X��`�LO\�Z�5̳���L:�9j�P뭒f�a�%�
���
�(8�S����ujyR�g/����H���_�3�lR��R&V%���W�{l"�'��7�i\(���YZȡ���_����Ҷ9�곖���W��Q�m���Ȅ�K�=7�-{aLՀD3i�$Nܠ����|���0}W)S\ߎ4�8�Jӆh�UH�&i�,s�3,A4ZÎ�T��2^ǩ��z׆����X�!�o���9��T�����eF�?��r-�^�d:!vܻ\˓=ǭn*����O���/0��q)/#�K����-S�czk"����'g@�N�5�b���1%0V`=���O����R"Fn�t��>z�C3��vx�#Vuu�k^��Uk�I\-䱅�!�t�$�B)xŐv�h}h��;t� ��/fP�eVC�	��\�:=ÉE�Se�5g͝��ƀ��%r���H�'T���Ǹ���\�w6��_�<�$%�J=YK;
�����ƺ���4-�J�j�w��S��7���M�>���ys�.�^���p�7���N�N�)�/b��_w�=���X��3��H�VVJǅ?�4Z�\�tR�Pq�d���';b�`��S���h�ʂ�O2fuh���I�SS�g��y5/=��`����S:�p
�>�:?XN/���uԙ6���3_�%伫2ݏ[=e���6t�[
�ŰJqp�z�T�x� R�_i����5,�"g����!|{�zZx�$�:��ց@��T`�(�Dp��90/��N�^n����J��w���-�	�~L�z8� ?��@�7ی�$�3�cT'����zj�8��DJ:%j9��!�V�i:/��i��<d���r�:�4<��R���,tͷ=�w��>���a-eGMȼ#�D����g�r\v����Χ�Xn#](�Z;}�D�:c�<�)�f��P��ŜR��Kj�>Y%W����m_R#�/�^�/J� �jJ������]���֬��_g��HX�m�\��[��u���S�Й�r�7��G��xWm!9��7�	WeQS �;�SN���S�OO�_|7E��?��1���XS�8v����_�S��²��v5~
@��6����<�X�$D6���GS�=���ϩ�F���v*$D@�\�_Eꇢ��4�"�խdR�K�o	�76�q��Q�\M���TQl^j�v3E���P�nUAI'[aU�C?���&j��r�hX��ƾ3!l$3�@؄����Rd��H����|���j���U" �Tp���x�ah>���B��3b�\����%�}7b�ŝ܋�f0��bY�����_(�)u:pi�(�8��, ��N�XA�PL���M^8= �*Y�q��M�+u4�k�����Zs�[Ě�y��0/�Z��L#U�$�P�M9�T]���{ ��c/��q/�!03Ou-�E�_6��ۊ|����!gP͖7���+cx�]f%5q�	b��.H��R��2�n�Q�]˥@��sB�EKf�NZ?�H���� ;X�nȯ+1Qd�Ֆ$
�;�;H��x�`�VU�=��3�V��?4�a�-%�]���M�n��j,�ؙ2�d��Dl.����Q"c�&�@-"����0d�?eF&��\bW��V�%o+ⴥ�Ŧݢ:{5��*8;���aT^�)�㳗��"u5��� ��[�ɎN\���
=���U��H�?��1�,䒰���p�V���}^q8�T`�l��m#[����6`?4�=.#3�����2���7���a92�xǌ�50}����7��?l������s츼A��z��d���]��jb�����q���=�i���z�+%�Z�CPE��0��?.1�ry܃����x�֏w+��9j��?����?�G�oI�H? %�%b�7h�y#��:�@�g�ȫ�CX��� _��|����Ɛ��E�pP{��8f����7�:��T�~<��T�W�����"|g'L���DQ���ͻ@	S�cR/$����F�%	�C&2�87�}�&�Q����6����q{n&L�'Cr{Z20��3���������+43���Yi����u=|�hp�5v�����a3�ݥ0���E�S�B$'ݜD�ԘW �����O׭�0�HF�}>%�m��O��~��w�y�[ze�d�E��-��E��lE �[A;��Z��H>�5�:FP�T>Nq7���7~��VRJ��Qt>����	�ͧ��7��V�]��M*��v�G�/8�]�!W����)��T�������+�F�JF�m}+�m�֒���	�����py@�5����g��?l츝R���$�dH1
��rG����G�Ѫj���m�&e�9l�_E���e���
�`��H5DFG�C*��[6�z�.%��l}<����Dn]��o�BIn�e4�U9w4}#?E�׫�m��P.��bdH2��}��:��9\3�5y�xvܱ;�����z�Ef� l�Ů8,d��V���Ә��^�K_�e/�����^��>p�@��~��1y�zG�]�
eA�\��!�}❻�ޓ^��ala�W��c;i��'s�[�8�s2	Ym���o��0�8�M^�h�����]VC�c��4B/.|���t�G�xg���/�zd.�0d��{Jo=��^09hEv�$f����z�Bz ���U�C�	Q]����W�t�Q�?zG������j@9N/H�ǃA²�9z��~Y�c&��V�!��#���
�	�N�{�]�_}�o5�ݎc��3%���f�����^vfr�쾯����DC���N�H�~�j�,�p����4`������-z:����M�O�����s��-�sF����dVG�"�a��E�=V_��������eCԨ�G����/�r17��fv��4�F�ZֶS��ʨ�E�P$؆��
�,���zh���'C�i�]Iz��v����p�Y6I&.j���N�<ht��HvQfl=���s�,G�K���y����B��S�87a)����z�wT!���r+ԫ3a�s�Ib`<W����q�����v8B�Ii5k��Q�=Lv);qcdM�.T̡��!5�>3@i���fCL��&�T����b?�ҟ������b��ä�B�\ �E��e�A5��2��N^/9}��v�̢t39�l�`3�e��O�1�sN��v��I=��]����d�B
��-3x�'q���ݯ۔)i�x �s8���?�0->��V��A�i�I��N6��&	�t���(y3����]�۳���K��d
�_է�,X�Ց�6s�p9�4��u��쉊��j�ҍ×�{dE�y���1��}\՛�c�殐\����*��RQ��:Fu���n��C�XA�.�A�޾�=�L{(�NF,QG� pc�/F��i�j��M������ꁡ+����TH�HP��e��G0��k�Y�S�ƅT�Hz$�5�Z�,�0�Fh��DK٭ԲO��K�_�J2��- P�iI�~I�a���\���ܜ��l��25H2g�"T��0z��Z� �=�qeV�y��q�,��`B���HN��E��6o�T�M'��:!�36N8A�f&&�u;��v Y��g�idS��2ck}t��9���
�4�DbZ�uP�@)�Mw@���m1'����y�"�2<�`��;��\�ѐ|,
��E����n�kq��#&�g���M�Ɲ���I;䈍��l1���TV����Ҹ��Z��%�6���c$���ϩ������z��c6~+b*xLؠ|�B�������S2�\�QC2���v"���[�4������$b�����U�����;|z��.R2=nS\Z�NE��MpA��?!x�2���O��I0���N��-�ʴ�l���Jj	7D|7}M������'����Λ6�-Jԁ/�*�]�5��d�["����T{6�A<��^�O\B�Y؂E��,�o?��6��{t=��/����id�T�?�E�� "��#���0�a|5�cF&t_�͑�($�C�#��P3���D���1So0ڇ�[-��	!9�*"���� �y�qC�5�憴H�7���շ�[C�s��vƤ��j�6���v,���ӈ�}D7�	,�w}���?�P$�%����.�NĄey����"똇8R���(X3@��Ň|G�����f������1�=06��d+�4���}����Йs��m;�<�� ����q�,�J����Y��A���������}�8/Ȍ'�b�g�]A~�@K��q3tae�`��"��AXu*˪!]�Ġ�u ��t�1@	�]�φ���w�˦A��r���BJ�ĔyUSyV�đ.,tt������S&qG��[S�@�ıC�������ˏ��i�/��&��T�«��#�?���祉��m$h��A3�����9h�v�i�|#B��Y�s��e�{ ~��Q���۴���ΝbC�ui�r)���r�a�EuSɳ_�
&f�߯���A��
]{���|��]h�!c*l&�idҤ�"���\��֥����w׈V�Է5�N�?�Kv�KQ/�6�B��Xj�G���� R�|@��T��
0s�(Zyy�%74	k.pqnٍA�2c����-@(����a;�l__��*E���a����e-����>� �{5eE6�1%L��6xB`2�n�~�i��x��8���Dn��7KK�a�(h�5�v��fs�!+�^T��7k���+c(>���84V��;%��6l��<�ߓt�M��m伂�VT䦎��F8�WG$t��7��w�4
��TSs��3E���T&�����:b\�s��ݳ+<�\�>ׄ�Bd��>�5�Y������	�#��! H�!QjGR�}�_�2��2���ߝ�|����m0c��voJS�[�ĻH
�dS���/2tc	Q�c辕�1u��9���i�x�����L�j���g�#�Q�R�#�YNW���A�O�����8�cR8cJq�{j�s=���t�l��D��
�x��h��XS�aj�y�k�/��Q�� <����]�?��098�ÇO6k�v��$�I�ɔ�>��:U �^���1�$���;n����I�V{_\7�m�%������P`��HZ؟wGzPկ�G��A�Ѫ�B��k�yP��>W7�t6ed1�'���ʘ|�H��EC�����v�������jJ�}2� �c(;O��{{���mg�T#mqO�{H�E�==���ru������{~�An��#�r�(R��)j Ӆ,���"~�d�F>��*"������ڹ~��8�
ƪF˝9TQ ��޽1F��$4ғ����P�I*D�A+#PBh�j+ :����)� ��ʨ�^���Q��5|mJ��(��U��
���h4�]��b�����"��Y���	�./A5h�&냚�NF�D�Q����h՛Rl�����W>�K�e$4c�����ٛ+��hu�NI�Cb�RA}�����E�nQ��{�Ц|`�ސ��t�T"v׸/Y��f�����KN��7�@��0���CM�,e,m�e��c����{�+D��#�w�ر0-�"p>�g�Y���Oh-�uhf�xeʝ�)@.�ب7:���	����O��x����O�~���T�:°M��&��cƜi邏�oO��vB1�� �!*;̡�SR:�#1��fjʳ��k��ŝ�O|%��jl������)%����▇J�W�wg�6�?�-�ۘQ�\��P��?\��m�׉з�EE}4��A-&��Ҍ��f�+�����;�rhV*�����f/��wd �*�����`���ɍ%3��slI�4^qX��6�l:��$Q�oI��p9���Q��S��;��'T!�9T���@db�ϻEm@�j2�5H*&��]4JA=8��J��I�V#O�ln~�>;֑�f|t����1�o-v��
�צ������:��U'�~G������В�bT��b����>͸���D����1,��v5W5vy��T�Ȟrz[��X`����6L_	�o����KL��f"p!�]�жX7~�Ú�h밟O��$�}��N��GA�ؽm�L��}%=
��u�Z�w[�}x3�ߐ��ԿQ'�ڣ�θ���^u�MLmbq�[ï���5=@^z�5OFO�L{ R�_sj&�X�eo�00D����:�[�ɐ���������[���op2�4�w�p��_^��]�g@�i4��/�V�	�{����πmD˧�����X^G���n&�fЯ=�#X����b�9��M�D���y�>�/o�"؇��G�6Z����Mtl�ӓُ�Ŏ"�z#Vmȵyo8e��9���K*��$�@�DA�!GXL"^�>���I�&�D�xF��/�����ލ>�gGj�"�xi�A���Cfs�D���-�w_�|%�3\�|����V��?d���򧑪�Bŝ|�e�b�k���7k	�9�8�u�.�ES�2�n�3���\�4���D`��E6N�|M�a\÷�p��(�`i�;te�~�=��>����iU�v��]��]������r~�ǲ�Ir/���~ɾs�GiU*�O�3'5�QA|��K쵁J�k5Zn��q{�YmA�ʱZ:�.h
��N�5�C5���We��"���{r��+ȅ��`�^�+�ם.�b8�">C:Ӡ��;M���N����1�	�jy=��׵'k����tTp�J]���y�1Er�H����R�Eqd_��]�4��a�=�g/�3`ܵ�52��?p��,�T��j���Fi�/X���̄�B�]o��3'Yqӷ �.��lk�0t�[�.j.�GZ5��\�=�����]�k0#��^��[�/��CCm��k]������������I�Ӽ���]�z�X�[D��r��ڌ[�	!���-����tSbD�������%ӷ�q�+H��y�Z��OqP�����
�2��D��A �B�'}0��` �B�x��ؒS�V}���đR��Gp>�+i����qc�R*Q/�*dH�%�O�/��[�%�lL��K+����Q�*��O:�,�{�QE.��a(��&�+�2��������x�����Q��|���pI���˘��VB�ڒ���� `(`A[���6~KW��Xd���e7�cb�����/U��s�Lzh{�ܟn���$�[��^�ԍ�wF�k	@\-�0�A�^Z��D�Oy�`N��¦�x��KE���J5ʱ<�t%�!$���X!�T�0��-K���jdێ��*���њ����& ��wh���բ��ǚj��zV�!�w�~p ��Xcw\m!��NG�Į&��3S~è��9���m�H����F�u��[+���3����W.m���<8O`ǃ�ʏ�t�e}`X��!J{1`�\�})�\~Uļ��2�_����{VL�	DYz"�M��3�2�-��o�� ��U���@���/����Q�~���Tٱ�=��M�v2<φ�@�x��)r2�x]���W�[{�n� ��=���`-�߇�Z�2kqX���gz���Bō��*x��5L������9�;����"[�`���n
= yɂ�Zm��S}�*�%\B9<٥��u��kCT�9U�i�v�N挪���tՓA �=�9s���Stm�zVPa���Pw�`��K��d�j��f=��
�!�5�����9fkv{�'&�A�1h�R(V>���=zRs�Nl��g���,�^2�uʡt�Haᐎ�>gN�����tT���[B���ƈN���?�����t@��	�x���"��B��5ăs��A=��h,u��b8�.�J�s�"}*�W�G �R����#W���8M{�%���Kk�À�������79@�/"��]p�'��;ۚ���&Q���7Ö����5�-G��#|���u����ɧ�[`��U��l���AVWWe��[a��B�l��� fL��m �s�
>7���-�o}Ӱe�z�O��m~h��~���� `ƢWq��&4i����������@ta;Ԑ#+L-N`��+�OU�C8�;T*3+������Ǧ����4�VJ�¦�WCn9	�w]և��;I|�s���ȱ
/�x�L[uX2l0T,ú���.�~U[b��ypL_�f�{.�.���<�A����h�2e��3���zq4#=�Q���"��&B�A�����X=��&���þb.�pU:0��N���4]�?����v�R���Z��Cߚ��j~�Vy�Vj�f
o���T�'"i7����:"����]��G�,�gj��LcuNќu�`V|�m@��d�/��Ou���@���[ q�w�Utp��/nԺ-���D�ݽ'Hc�����P:1u���8{Zq
}�e �_y.�5i_%�0�y�f/�
��E��2�F��iCN�y�����i6*��;f��B���U;�<��#�ݨ$�3hV��L�_yY�G9����6O��|{�-�9c�AFt�����}<y'�N����e���������4_��,2����6""�>2;�2��9Q���k�k����WD�u}�u׋�l�Tʧ��%-TY,~&���>����k�ˍ�NO.�B��p���d噱&IP�}M��*hA��yN$F[�>�x��<�\���,�`�;A/�v+��]�����W�2l�ʦ�t�G�L�#D���E������V
�)�z��a�s��RE�E"��]v~�&�,�ok�K���Z����e\�Ys�F{�t
r�Qy9TJ��c+r�w�3y�s���7����[���m\�#�٦1kkb��9<��צ�S����o\�7M��F�l0��uZ��	T����
���z����h�X���Go*�x��_��}���ڤݪ��c��IZo��˴��k;o��ל,Bd���� ��.���E��|�1��Ȓd�ɟ�,_j='����?^^������;�
�<����I���}��d�H�-ȑH��Ӧ�U�S�V��&�"s7�-8��ed	�Ѳ�^��n�cGa$�q��z\G�� Y��%U�Y߾=�{,�#�$��-��jgb��=��
 �h�R�c�'ł�����g8 �!G�U���K�yG���M���픤����q���H1{�����X�N��O�����Å�;n|�}�]S���k���!��\g�A����2�ϲGf�����
������Y#�l#ci2�e^RT�?7�Rh�ࡅ;���z�?J�v\?�~�r��5��t�qB�.W`�Ñ�A@�K{����Đ?\0洐 I�?�	PK�����Y�K���8!��<_(�K}3�9�.*2������y~'�ڴ���I���}�ڲ
t��M�z��6_	�!BJ4xC��K.u�m�6��4cs���%���������D�Si��qI=����/rśl��7�g���z%�)$9橷����Ҙ�����L��uv�����t_��v
2?~2Q�Tj�d_^R�� G@�ej3��'H��v�a���Ɋ���I�S]��4���:�`��v�j��6k�/�vy^$��U�8-��E���ֹ1ϛ��|Ɠ|��z��6~�oHoX��m=��Ew*�n�����+y~��ĈR�m�hw��t�+
;H�������C��\��:��%�ڀ�1���1T����
I��O[� �* �Y��o�#����2*j^����w/vi�~p��"xں�G0{���ue��<��Q���l��,��us�^�`?�y}U���Vq)t���ӗ�k����KYm]e�U�����j�e��<w�F�AMg��?�1�v���5��,����T����d�(��!��ԆQ��G+������A=߻ ������
��棅H�v��ܔɶ!�@d�	|���k)�iM7�$� �4�Wy�:_I��>fh{Ƃ�6*īh0�+�c���T��|Ǩ.��:7��_�[��>=���Z瑜�&��`\�n��}f�<���!��h�@G~��0��Ha���:r ͎YA3�ʀ��i��Xp��EXSz�$��>�CwB��ʊ����-��α������m���S�MG�+��Id���wܵ��57���}|&(�$me.��~#F}�rTX���Li����@�6�kA-_������<�|U�k� ��a�E2�h�,�C'G8 `�2�����/z0�#n����e�#/\��d�C�� �4����������~��Y\T"&���?Ѭ6YG(}�����B������?��ܐ\�!I֠U�h_�B��'2Y#m7��?5����b�=��8Ns���V��X��ӏ�:��"�BR_9h�Dq�g���h����VL�p�_h�2d�
}3�8v}���eVyqM��Ec����5��Lqa��s�4�6�_m/��<����p��v{e�a䣤:�d. @m����	��h�{�ɘ��?fg���Yz�E�h�t���YW�1�9t�6��?��:�	��/&;�<�@��	��0�C�9�#��=VcQ}{%Jΰg�|�2�/�ؾ���:��L��鎚��8{�fP)�Me�ׅ6��T3�f���iA�o�ޯ�^��[�g���1_���*�\���� 	�����#�!����d�ۅ�D�T���3���XV�!��|���*oï�jfHQ�z"赮R*1{��G;�=��\X'cbL��'8$�3Z2M�����&  ����~�m�7�X{ zh���P}�H��G��_���i����3Q[`�n1����஌l�g%�GngZzK��ߎ_�m`�I��߁zջʥ퐳�g)N�����a���t�m�K�ܻl@��d^](�p��������U
�?0F�?��2��Ba�<�.}�^�3[XkA"�?�$�������>�R�`#�ې�C��<����+��l�>��3�6�՞57�fL��� ������9f�J�|��Δ��n�+�ݾ�-�o�e�+�k?u���0�'$�2CK1�[Im��M�q?��^[�	�m�;oҧ��7��g@F���8 �W���iJ��v��тm,=��KWӬO�2����_M�G�Ym�OH�_�@��^N�@��CfG�0�2��mXp���)�W�x9~O�n
 �]�/�Yw�܃DPY��Ņ�N������Qeu(��ͼD�!�+����<h��'�{<Ƒ���Ǒ�
�^�@_HU�Re˺
���[����_M��g7En*;��r@TJ<�E��B��g�L@��-�Q�*�y66䩸b�A��N� xi�F�m��/�L:����_��2T<z�SG|#������0��ƴd#( ��4ϥ�4�jP-��q)�0tor��g��Ofe_�a�4�4���']s�U���BjZNƝs5�5�HRW�V��i^,>RPF�(��˜%ϟ(�h��,c��
��H��	K)L�C��r��Ήֿ@��/�O>:��l�"�
�ߘN������;��0�[���ZA�����=U�+���0�BLX
�����Q0F`'w����X�x .��2I��9
�^9���y�z�#�6�HW�:�n������,�$Ū4��_��b�`�t��9�RU��%�p:`�ؖ�y�[�U�T�A��%�#.�0��I*�t��XA[����e�X�7��'O!x�a�ً�]�<��W{�&[���bڏ �֨�3)�����C���p9��މ���l�o&ǁۆ|�"��m��2d�{k6�5��9���y.Ԕ��P����!@k`���2�C��3e+f���mn[]zyC���n���1Fz��ç2�u=w�Ժ_��1G��4��WD�רg�9�����Ͱ�1��m=� ~%D��g�ZWZT&4�W#�b���K�?�Uе� 9쏶{�b����+�w����ڈM4ݿn+'�X����T���ȇ���svxg����&�0�)�5)�6D��%����$`��$1 �_*`��"�ЩBz�@�j ����FiK�:sEȎL���N�ɹ��j�-��0��[�v�pd�9�@G�[<��3�žh]��1v ?�9���-��>�R"�g���gI?��V����7?n�IҊEJ*�	o�ΑS��Mt� z���?��v)p$�����W���9;w���I�?}üO���p��h��G ��׭A$*��*� 4֕���~���yY��=��\:0�!�=Y=l[L6Ew{�>L��*�<�P�l�S�2_@r�I�9�×��~nxt	���������wN�@�<΅����R<�i88����9�BX�d\��գ�kW:I��t�K���K~�X7ع�L�&0O�9/p�q���ᅏ�������!sC�H�N���HN���%�1c����;�R�&H��I糌������(`��������F�S+���;��g�r#^��u�1J�y[��8S5�sl�S<��bΒ��p5w��@�nN*$�${��c�ˈ��i�XR��O��YfM�f��"���6i5?`��K.�h���oJ��i�w��e����jؕO=hL�O����բ�}Kb�g�rW��6GKC72͇_<�D�o���I���\�d�C����@\n+���$�'��+ ��+W
�YZ� �ٷeĠ���pK̎�H����)���X��5������Ӹ����Z+��*���D�
e>`O�������4�쓊�{O�
�cVιS���P[���)�z�OܐfJY��B�]#�'C�ER����21���tb{z䅉��ad	M[?���W)��
��'o�l�䣊y��?꧖V�^��0N�=B���9�F�X���
��BFhQ����&���i�'�܈G/0��R����o�8��LMk�c(C(����G��X�!��l���riT�؁!/�������v���R;�
OX=���Q	Xb#�Y����$'���g�5�H����#���X��%��@D�Όٵ����j����	���άGp� �HtS�;���p��
*4\PF�!��s�1%�e�����p<ϩ�,Y�����x�U؎�<��l¤�Ɣ�C��]������!�4�(H=���~��1��A.i�`���^gV��)�2
��D�\!2�F
��8A��ܞ�7;\^B�q�f�6^@�tz랉]#��H�`㬭a8�xY6�=\-�V4�띵դ	MYSz��,�F�)�?:A���1
�W�^�C�6C�z�����C6��Y�9ݭ�&y^�=ӦX�q�|ӴԌ�Q�z���Mue�%n�Q-���qj����V!�fa`�c&n�:U�͂L�c��Q'���+�e��b�;�SQz�3��v"�ufB�o��~H���{m�/-�m�i���M�c���ʒy�L9xl�|$���%j�Cؼ�%Y��4�����zX� π�P�����o՘֩60s���@��K�-��OE��)���TA[\��ٙ��}*�������+���񛞑{�&X����YM�f��g���e�V�k>��G�nXJǾ���B��g-o���^�a���&����yfD&!&�{�_/H�q�3+�ׇ>�$H�7�(�ҝ�OU8z��m��o!(�(o赪��g0h.e �N L;`���� �\B��ޏ�`z~����>�j7����,?�l�6Wh�Nl*`V��Ț�3��K^�FfM�� Y�uC���G����?ȥa�w+˯I\�ޫI�LE�hz�ӄ���R���h�8�v��id���'zL�[2si��R��dm�n����)��+�06Og2��'�� 9Je?�X'��J�nѿ�I��O5�a��J|�|"�� �t1|�T��$�k7c)*g��:��!6�C��eN������dEU���{�&L�4�Q~}�$��E��0I�Iߊ����V�����I�8��u���t��99/c_������{F~T���>i�Frvw�
�D�J�A_�9�⮀��#�L�($�{���pkE�����4��O����2���a�=��ĢsP��Ϡ��2䐜�]v�S2!��|��Q���:���^���`�|$	����*#��71��%(�sj_k�vz=����%|*!
���a��fk�p�YN�rÏ�Uܶ��>����MБ~
Ք��8�E��^���IjM�*�Ӊ�-��#Z���Nps�$��I��Fix��߭M����yMи}'�3�����O��Ky�2�k_ݴ�u���ݪ�/ ��LA����P������WA���4|}T�8�[v�Ƚ�24 `�b�0�~Nl-/�J_��J�Vo��䭦c�v�m�s��FXbD�˹�3̤�����czt�Em?e�j�mv��~���yԵtk��U�ޝ���n�i�,�������_�m��f��L�Xy��~~�Qsi[ߖ�[T�}�gY:�ů�@G~���\�E�������rc���DK�(:��8>���̩�{���V��}h!�x9Z��I�K#�Ʉ	v��⯒��w#�w����(B��S2���i�� Qд���#vp�p��n�2m�����?X�I�kȁ���]��!����5�MY�5�~=p�s��O�\]*f�y�%d�Icb�𐲖@�1�(Gc�|�~Oo�*�ҨbN��s?�A_Ɨ�;�\|��_�ȷ�ri����k_�$�Fq��/.�"XA7�o}&[�yi��I���}fA[d�OGL�[�Y��`���o��ު�Q���e�'����K�,I����RXP��Yg�¡��P�K%����u�b��Xإ��i.��~:X�%LTzbs,0`
J��L�b�O��7��+���&�Oe��8c׾EYWM�S�ه;��4cV�Bt�;�t���Ln�j��'�2� ��F��1K�Qu��Z��E�
�g�G��;��nO"�_07{hӖ�!A&s ��O8�9qq� �"��$�ɹ4L7OA�b�k�zu�{,���p�H�0����hs�4�F ������P�h0���� /�
��BOr�^�+vy� (���2'���+��Z_-�e����rw�����,�#=K�ǌ����|H���~��bItG�q��N���I[ÃV�eK�g����p����(<�.vE�ɢg�����֓#6 /ʈ_�g�'��mk�i�Y^�����C���������El?�]�B�(�N�9����/,����wPP��*i�x� C)�A���Bn� ���I*׹�����X�o���w̿-_?�K`]I�JUksK�X�� I�؏g�J$�~���v4�c ���k�o���
�()}��s�
cL�4=	�����ʇY��{J�P��������p]{�=�_+\S�!��3U�U��&ʲѠq�AMz��ڽl��ᐧ�{���e2�z�%��w)���0�Hn���3*�6za��r���n/?�!e���@�m$��a�Zu��y��1*\�R��*E�QL�2�����7�����U-�����ܛ^��_�KhM�3? �%���]�n��^�:G0=�P�{�f���������������'��P�OgJ�ҁ%���0E.��5�ߨ_Y�6D�_�E�v�����I��	�n�N2g�L{��䱯U��?��^0�e=�S�0����c��N`�ѽK:7a�FˣjV��+~����� .J�&��"��� &�7�I����㗛(U������SJx��*�%6�8Q
�l��[�l�%^��z�7�����e �LL�L�r�6�=�f�/0�XE� TR8X�q
��a������cp���ُ��"q3+�b%e>ߢ�ۓ��"�k�[��게W����g����0�m�9��m����H���Fʽ�	C���D1Yw�p�"���EZ���eɌqXh�|��	+7S�[�h���&+[p�5�í�.��f��1��6�����#C�C�Κ4W�-�R�iq�݋�Ȗ��N���0�t���a��N�N�Ͽ���#.7�#���<��иF\�bD�Gc���K�٢H�7�٘:�^4EFc)5�S��M���T�޹����YOdX;�z��]�����w���X�Ff����iR؉/��|�[g��(��.z�*�'���E� �欅�{��\��@q�Y+�PsOn&�n��B�*��BB��Q�P �Xj��s�Vũ���'��r��>�ͱ�a��9�,�MB���Y��D@SKªJ���|&�`�-�j4����TD{/D�`Y��4���>UiC0s��u�1��WCtIЭ����cv���OG���A��؇��f���stA6�iHîaE-�|D�#&L�tu��#�szZ2��w��5r(fz-d&l�C�����'h�\��5��0ϱ�f�>�e�?q�L��P�k�}��`�¦�8vŎ��!��D$�cAM4�\q��愁]��J�7B���D���:�J]]�M��+�/_-��d�Y����UtL���j��Fe�Yk�p[��Я�������G�')
�1Š�����!�>�2Ķ���)7��e'j\�S� eRc<�s6��=̐�KA��S�	b��-�kxi�:cغZ>:�`L LYn���5�	x3:��X2�X�E�#0�ѮJ�l��X�2�O\�q��𗖪�2����:,�u�}�UC��ձ���+Q&9���iP�%��v�-���'4�7y^��ɉ�[I�y���Rl�4t��qC�����	�����Q���{��C�SA�XA�nj��ԕf�K��^�*���'��KT���uW��镭\�X�A��]����|B�',=�)���Q�^i� � �)6��Z�wQBq�՗�_�F��D�������v�G�C��'�(�$�"k~Ta�[1�91���ǋ	~������~�QR삛V���N�K��%���9d#���'��l�����\��e�Θ��&5���~�L.:H���4[�s�}֩��\�x<��(L��G`K�ۛ���udl�,�����W�z���(g�ʟ��_;e�T�����=����,��E� �fPEkJ�ۿoÈ�a��k�צ���μc��xZ��Ab���ꬾ��N����4����d�O�7�	Yͥ�|k�^]�g�ϴ ұ�tí"�!\,݃��Ә�I_�@�:���2{r�9쌯����3T�O�Iz^+�)+�h��9��P[�����"�X�4�^5X[Ϝ�aم�U0㴞�$�^82кw����O�!�WVhE_�<� ����h�Rj���ī���+n����a��h��"��g�R�.�j�s�ȑQ ��c���Օ��<c����G�#�A�Lj�U=Kk�fp��(�[���q�����.�$V毷ؚ��jT%����q�')Ǿ����&��*K�PZ�5���.E&�K�5��������޸p�P���$�}>@A�Z��4��X�!��%~G�[2�˯u	Cn��E1�֭n	��T$鎊��ѧ�G��XxF4��b�M�(r��"� ��x�耜w��Iug�0�R�ʵ�_T�.��G	�2���AiE��T|;��)��$���G"bI1[hVo��"D�F�0�k��馒jC�|D�R¶F�&��UK��5V��l�)���� ��s�]l��ӆ`��^�`i��u���>!˨/��^��l�!?��rt����~���呮Z>}x�R�$�����a�4:mnݷ��mD�֥:o������c��Q�.%Fs��4�R\o3��t^ސ�7��?uNt��.��s�:yx��!g��2]~�';�I�P��߻op�ڸ��s/h�;� ̴m0�^J,��1�6�V��|^W'�
��W-xKp��ո�(�ԣѸIئ�z��������]��ݰ�Ӽg��������R�f�H�s��PR<8�d.XkI?ӫ>poN:.�V$������8w�Yz���d��G���d�'��iꭰ8�c�*:.�J4�~�aU�����ԣɮD�Ҍ �[I��Q� W��U1|��i��/d	h��ax���o�c���'?6ta�4���諪���=U����8�&ʟdܖ�0|�3d}8��@�|�/�t�h�p��c��uJN����Z����`�`���p��LYs�wm�L]މ�� ��f�jԣ���������������W&���ѝJ;ߩ�������s�	� *�+�\�=tdH�&�}�
;S�;��w-[ER� 1T���k��B�e4�,75]�hٚKD�5c��|�3�lUb
QӚd	8ZTE|ja�Ҩ�UƎ�-��>��m��q�n	��h�$�����͔��K�m�H^�Jq�c)���h��D����s	�ae�bT�O�mC�-�!�_�xbqur"��~س���ta6�^����;'���S���n4�Gf�
�ww���57)�j�W�9L��L�-4O7٣��n�KĽ�z�w�QL��l���	�.ɡ˫X*�-�ʢ��|���IWxv L��չpa�8n�ia�M���2}#�C���Y��3*�CW�.s79y��O��Xi�1}��
ణc�Dp��b6�1M�^�:�@7�)3���,�5��_K�gO���K���$����<�}I��ZòP����
��xa]|�%�d39`����u����<�GMJ:o�b3�"�k	8���2�H�:5Z����
�3UT��-(�1�J;$��N�z���(���y��߱[1�����U�r�؜#1�XF'�I5=l�f��gt���Al��:hB��)Ibo9�Mv*6)�߄���f=��!�&;�x���Wf�7a��9-H+1���5��8��+]�L���[��7`[����zGܯ)�5�h�����M�����,�d�j��_���#�{�%oq����䀾z�G�8�άԖ%)=>��^2��3#P߹㼆8���)��ېަҼܞ����*���gc��2�Z��[���9�!����n^�1��[D6���H���+s7HI��L��;�1J�۬��H�v��r'��c�5�N���-[_�ңWe-%���3� ��y^>n�O%�Z3�����˫�d�IkU��G�� ����t��;D�Bn)'r�ި�g��	�A\'K���϶R�u�4y(����}����Z�D�%
�X��M���M~�QS�#�֓�����D���g{TZrO��.�<.�,��<��6��w����3� ��ӹkTp�}�y]�55",���4!v*��dl��hV���(��<�v��ۃvФ$����i_4�$ٖ3���Sa�@��3�����@
�X����Q���W�آև~���C��"N�Cf}L�Y�� �p�L���J*�:���8 ��=��Y,4��/ĺ�c��]S�$|�����1c7_j�B�����ň��� rW�$�� �s ���WA���3?�p��)H
ZO�%��a�E�YP�S\�,��k�hR ��� _���!(��z<|2<}��d��9%��N�h�۩��t����[K8RQ�o��9�:J�w�wj0Dth�GX4�+�(�?���| �vk��3�G�J2�m.�$����1�nF��%y�������xj��R�Z��0+!��m^&�9�ƪl�	꤮�g���T�o����bl���� �n+%k�j���m�z�P�ȑ�B� ��#Y�~�S��ۀVC�ZaN�M��8´~��ηo���X���-�!��Cy�b�]$BU��Ff\�ũ�,F�|N��T9;�U���i~��	�S|�4���bf*��v�n_�C�1��؅�Od٭�4{5:��5����ųW���:��t�b��j��JE�LF�Ry?W���p��w��!Tu}Ob���0?�C��y��Q;�U����6}]��}8�}$���]]~aK���C��M�Ge����gq����Qu�o�l�}E������P��m|+�Ӗ����+y�<�_�h�Kߪ+��wr=Sx5?�I!WO�����	.Q��]:�V�O��x�p�G!j��GF�|Nש�	N�rV�f��Wj��c�w�+�Av5#PP<�
UQ�%�N<T��w�{���^!w �J�N�)G9�ҏ��PC�v���f�U[���k�%{���諡��'%N �@��NZ�k޺��O�~Oͷ��p�2X�TsHJH~ú���`�S&KCÄ+G�j��||8�!'�0C]^g����X�w�M�$i��?E��%8|0)[�3�p�*�~�Ð�Ȟ��[��fq���$P
.q"u��2�aa/�^*��n�O��{�ԕU�\0*��̔��A@.`���������=��m�h�����
_�O��Փ�����?'�>���q�ұw{��ْ��׳��@�����D��͑l���_O_��%m_:����_�`�\w�����*�<��pϓ?�=�(�:�w��N�cL��7f�c
�Y8������i|���5��	ar;5}�NX��{�֓�'��M� �qq��qͧ��'���i��^���-��6A�
�,�m�	um*e&Z`?�r�J�S����3S�o�� }�)lf�K���Y� z���`�/k��J�17.��3,���c�K��q�n�~� ����F����	�R�/M������Cb�k2y��5����%�o0}���@&��c�b:���<Kw�����`6�O0��|>��;6]�7Y�����+|B��9����TG#I^�u`��	� ����d�).�N�)�Z�t|\߹������Sn$P\�V��
9�T��\�F�ɠ�RX���)��լ�T��zrB�q4f�(�M����D�Y��bxL~�����V&U]��X��J���Z�