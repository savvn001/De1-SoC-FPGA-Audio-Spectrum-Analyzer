-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0G3g2bw5TESDXWIoS3WhqEEim0Ww8WmUSW1So4wpX6x98JGi3W47BGb9vM18u8aMOLc59bXf6hsX
9fCIB7zFGNQJjK/nkEEjRWU8Rml1GWEnqWRyPk10BgFLV0Nq7SMQ07ZLZZML885915bOjA40QM93
qr7JCSm/Ixg7zfKs267mG3fOYEKAKXJJmiZ6TF+hEPDyHeIquTwq/gYSDyZ7WRR5c/FMySBJEu3B
w0GE2Lf3naxzcLCi6mM8mNWm+EhymgkL7EIgVKF23JymPxpH/s7k/1MAZkm8HxOGX9XRQsF0wxGO
H+8sKVRBg6HzDA2z/zjmE4BdMqdMQQqdPUo2rA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
ieUMZQI+b4nBTxQQE8/Tj/wfYBEsvY4RpafMUIAigb8B9fkfF7bm9EgZ6om1vU3bAGcmFSpATb4F
KVmRScwlH+424R09U/6qfU2jxo0GmXbhAudxgOJpdwUltXgdaN60tSFSfMB0X4t93VXDevnXRyC9
E44s2YTuUbcLH6lHq1aP2M1GabEDH+AiuGTzzisC8H9Z9JYUmOmGvAmaNsMbYKx1qVgNc92GGl6u
LM1c6KJp1UCR5zc0kpW16UGNLeSs6EdUGjJKM2XeAs9s3K/7WmLxfjNWn81CdzEyMOR3FsWg3j4n
motIbsCDDTCGvgbFzqh6jHZqWvVLq0RGupCu/0LxF8VK7LeyLgZgT4WGJ8RlREi/mXWg8qNT9RXZ
di1bFZDlKgTr2eGJA5sA9gwxfMWZg2k5age7PSlvxDjUQYu53vOoyzC6VgfS4i1v3/MGiAT95BE1
eQbOuzpHVDQ2FXWCQ+w/TZGMHcW/dqN8hntbk0IMnuPorznWeaFlAQv4kp8x8oyY54Y5N0A4F3Dy
5HLjEKF5flLqjM96SdnXePEM4kfFYcLx7EQNpkD4RIvOS0+l9+wcvJmlV6UrrPHrhiBE4WtXealD
fP6aWQvxnBm6k3yy+YHDeoIGedwUAe10oXxjkoPy4saIrWKkhmlNAgr+XnPTetwMdSYnkLTh/pKT
JL8RNLbkNPiehjI3/fAdJFG3BPGszbVHydPRxkfPrHZsljVy1rKfdtitzGUnaoNl4tGCRtWqpfOy
1zbeHT6mYaICBNLDyrtlKpJTG2e/rqhc1m/UyaSSsm+ft9kHd+Arml5wbDTvMx6d/uZ2frJykbEy
Qj7bdaGfstVZF0kTNnKzvTn7gBL1/jkGlfwsDkHzOTA/iUDjgqP+0feSqPH6PkVFY4t1Cc2zhmU9
xX7jZbcBqLNvhVW+OdN8wLxpk8UxRd+p12oQLe4271kY4xpg+yzVWxhu7o3S8weXibpOzjKml2FG
uTxlvUwtsTBGUZVG/n41PWtLNuI1HCVYWLMm8vh7AUtUgSlxxZHYovTpYyCGfMzkF1QpchjnejwC
k9H34uI6h1BTQam5pRTPbNprCNe0JpaE0kZiHAkN3kXkRJP4ZdoqBdrkVnoNoUN5p0WNF/6gIsYT
K3qkDpHP4EfX8/hfFn5qHjo7BCbaqGkYXOiwA79IsC7gArdunOtw8+1QH1dJjz58W1BhDy8/i+JK
6qL1XwbBnErhmAB+nmZVqqGsBkUK8JBgqcbztUEJ5gTip+BL/aMzk+hAS7UUdDXScb7m06Zq9LU3
xYm63ex5FFSA1CQoVcxxltZpONcH87qroNSz4X6CxpX9oJ6ewssyDY3QSoRDtmCerNmnvBwsYh5O
Qc5YYX3Qe0RU+KIoNWsy7uXvOCqkoxhr8G3PEL9j/FtEI+0TWTtB4tMHKK/Uh6hbOewgW8hpKVSj
eiUt3ZKsmPKQsEZYh29xdIfMK3sLZVG0cfdNeo4dQ6/rfHtrpoRgD/tOsAbIRknAGSV0PUkZXNNo
rGB3LzK4lf2q+DhcYZB1KvY0k2gkjSZpafKfCPYuYM+qgX7tXdwVS7qgJ2vTpQV3/39nBl4F6WED
F++P3XoH0vQgnHXg+dpYgAeW9kxwDqwGNQZCbv+T6lMSA0eH4Dnkbts+Lo7wZC6qdIgYYK7DRgbE
QOcei2Jn3V2aJcaOKUwhuVh0byKKtYEFjcgWQxxfTLI1AYwuLms8lmtLEq/4EGWcAtAiME7SBbdc
B4v+3ud8KJ2nqqJNks89YFevX/gHhZnKr2zB6GrL92yQW7ti5LCWWHTSlwJ/bFpb8dXA3JLVg+W2
21gGEOyQFFPx5aLXClUUlGYgf8P0AjpSb4aGoJm9FG97cfGyhuTiQLnOqVRp+EC7deAvoOzrWdbZ
cjM5EBP9e1i/GYjy7XmGOUx475UR7VwqCDRI/MIdG07ckKaBgDEBv4Z9hZcSGygD6vc2c5Bxbuvh
KNq9yKQUPQ+Fwx6Y0jWbZNzrwZuJiIEiJNsiRdokktaFF70S57bBPDeVfPXcUM0nsLlp0VSrOnhr
prEy7D6sU0DhzRTeAK3qdIRC0KDQgHp7o5mdCrS8OBXjL8PZ61s7aNmZFjb7vE0ov8e2OO9dT06m
bCF+a+Wxfjop1G9do2E5Ln8I4ijK/TquIMgvjVXS8zcAKCgYUqoW+HrbRkB6iFjBxVPXr3XjdAYe
IAo8hLn9j5HbaT6yymBaIOCeoE1oqzMG/Z0hsBDMLPaZJwK4wPle5/PbSaelvpFameuEebrkc575
ZAfnKsBN6ZByuVenHGy/p3oIAkgDNnCwvZSEvsPjFINOxvM/r+vtT9x2PjZ2nxrvHTdhY7E6r54H
Ouuy/ZZPEWG1OY6eavtBtL7dALbwK1Cr8JsJ14+JE0Fhvu+NK7nZn8spiuWGE1N8+bds3GK+wbEn
p5NmbM2qlVQZXIR73e4dO0N375ACWWYwsL4ErPHm+qyUcV2+Wt3TrlZC4p6FxIreNytKAUaTqQGU
AqZ6owhQtkiqw2jmcVrLBnlAKSvyYpEZ7JaW2WeHCibZz4HO7ejeVcZWX7CFH4GjPx3Cw9w8Jl/m
MKziLomfyrAUmXHY6AOF9hyafuYq6Xt8vW7wZuP77yyPy/Il7uQV5fAjBdB/SbdrOFOaEXwbevCV
qaHnnP2d7C63EAThNbsWTCEzBBh8VmmNzJWOQ3dDiutj3Je51HLwjiPTLqkzr2cpA2n1xsF1WXIo
ERAf1dEqaT34UcmPQjvbt29BYRlKX5GdPejfuTF2pKLjUfxnSTYojfbUPN8yNML54MAfw4oHsw0Q
2at5/zdhCXAPc1Df0BQjaxUivwnc/EIgfBL868oz2SOqgcmyL9sDh3rBrCsWVaAt0yroaq4F/xkR
yk8EKr4aF6QNLnKz0TTSdIb5lVFl4UYt5/j59IhPKElsQOOGg82xnMqgXRVWrzeVWxFzi7U4CTER
d3O8ZYtgonhyzndvtLauxuYRyqD1BTnLpNj67LTEkCJzyy6ExvLdrHJLlh1ACQgdQyPMRc+K/Lzp
3c1MFID42YNlK1yewrvff/tiXGlow/9kMHoPVqZf6kfQweYa0iywOkC3ELwzBreOP0vRfiFTe7oc
cOLhMC8EK+3bxvN3Sul6E5/Iqbj4+rCZmXTuCc4qEN+szssOvAY7xhdMlR7v+AW0ixCoKmJ2Wy2g
L8Ir52UgYQkhnXrtU6pP1ldHL0QKBmBZS1hUOnaMNV8tJxDRal4e+eQN/UQVAJzSN2mJpDgAqr/K
GcuEXd5uK6/0V2awf06irN9KGt05Y3/GGt3Pujzsz/CQ4a4OIOsodzqyRRBNEfphAcKrWKCij/17
Cen/aW2+8uWkEKbKPkRg5iEB7wPxTHdcDnzAvIVg3/rCYXrcifib3UcXbxOqpzuP1JToSTahEGSD
j1uOBhs3Z5JRJEI5EJj8fvgttpfqEtlK6dSiSWZUqI401JzBjjktAtAeR/kNJmZW7qXJ9rOa45ML
oYXTvmWbPjgnC2jMBz6llyiUgnKI0Eg9j7AB6rtTAon+qs9ca1T1uXeL1QqUQ5K4GSNvYJ+NOAEd
gcSCGZaJdNp0Sd3SHHhfraV+rNu9TQL0Moflgq0ax1h+aFZoLk3Aq02KLDSrLj1h5EA5DtE28qUc
WS1SWIWx1bOqWZKc+YKLmQ0mGtQjiu2j/3/uDlxdLKHdY7/HJhn2prL8J834rvKLX2pOu/BJv38n
pL5lBxp4dgYCP3AUpS8DhdpYiB5aOI6hCPsGXxt66ZwZkd2VO9Kem6C22b7B8idKGPpjHx56BMuQ
0NxsSAA5y4bwch/E6SDKZO0/1TbLXMFH5q2GLr9h1OBI5Rsw8suDLoV8qxLFZTSi/fQEZG/Qokoj
X2azWJUgTPp0pC/nzDgx8d7kjgVytOa5WF8uYmaFlvTZQMudNii1rgkGEA4dyb0CVXmFf/beD5F8
qvu1toNkvq9e7M0Je3phnS4Fgxz6lMKM5TcRvkKpI1pvBq+Yw6I6IyV2VNVa5hHvWgbkwEI0Goa0
3yx2+TEdx8JVEIQkCdCgFWHkffPeVBqCbkid2ih+UpZMuujnp0FAhPaDv/4T5y9YGQLlRFRtbeoS
8J2o+kOyYrgRLKDlevEk2PzDvs7KZrbdS5Su+xpIi3sdIx/NLQuHn/a8Qroa5cjA5YaH6+ImLkUn
mP/DAGrQlJdV7KvdZUlYsLZyCt1fgedzNvE7NRlL9+deyOa8Dx2peWK5BQmvmnBCzxwm+Ua3iP5i
3vS20LdoxvK2DNXf9Om0ZZ1sy2UPJ4h1H4TQG/W9sxPxfDW8tcIwsz+0wJm6Gqh7F6BFi6OdEgvT
ukeTx6VwKt5ItqlgCdbf9Iv3tFusLRX83K5FtYL7i4yxyDXDOrYphh5I7YvcEGYzU/sjswyj7nLa
hYSsYDd4myUynr3sb9JhwrbzSPvV7qkU+OHCrBUGT9V3XbE5okL3dPja3rNLBJ6kJwRxHhAtbEFT
BrXFRPdxFSgSYgxahODEGXDgfJ5C8ArGFenj6/PsWQMDuO/fO/MWwB2BTngpsQ2qekreAtCZ9S9Q
EZTtsOjqeoMK6HcmizJM5tSCrWrALXp0+GLIG1Xb170YCwOg3IBHB6UzAT4D6kNh1vGl1GWxpYYJ
PAYXrpz5D2CmH+hwy5zXNG8PS35ETBQm1+hbu0paxFJ3wA1CGmGnUCENq02CoJgQP9XDP/by9Qvh
+v+/tMiKTCRNmuEpvsvf1vxfaNiHEloQCgzS6LHMTVyTpWh1pz1h7WglNi9D0gny/LME2VyTRGH4
SexJiZgNAkqkzRuaTIhZN+GYdB7iONAs+uHt3gh3UB9lWiRPKMI3c/d4/N5PH5nOQL3sYex/1VCT
Z0siRk+WOgEPmMHQueX8tJ3gEY4ddenwXiGJDf4spSYGEHVPTR5778Xi2f+3IFafp7CkTXpnlYtL
KBzuVQMZKGpV+QAXCLvqD9qhRH//RDlg+KwzMAvcSk3aqAV4y1FhqpYUHNOW6VRU1He2oJvN4j0u
6Vn44t42Yd7um3drIOMseZRYSVBu8+iLd5JikPVHtw9+JjQez+02982duRs72axrPg+uAscMzOiv
F3fB+XXgQnFxxRZjy4tsh5l1slT6Lie+ZKHF3KfT0lEsI/SMw06cM3elkeMc+3Tj34PaFdwPwQ3+
G+Yfmk0GknY+sDFFPZ4tFiHYCPETUZA/8Y3x4oO6U5GXzuH+2XHr5fQ6tTWb2SVWL53rCmBCpS+U
tP861NcTGHeevr/xZ7WIgzLfbgoCxD0Af56bPPorPqLf1uDBhTukn5Uox62YKVEiYWvVkaS1U1P6
85e4Lj0djPDEHQ0UI74LxjI4XMDmCaKJsBHfNA4dvvezfny2Bay43/5WwBvjoR9VJ2QpPW+SiKwi
XfJAGFncO6fVbXP7XW2s41yc0u3qKI1p1YlRCTBgUDALd41xq8puW2wookMsVOiB9tOfv3H5c7jC
m9/tgZdVOXEOMDKwnz6Bhh3NOAZbIBBTSfhGdv6Go6KQ11KzZ7x375XTiyIzfA9B/HLfZhquLI1G
Q72I1cm0k61IZNx/WEVyJqlTa8a1k9S4JGT3u931raZulKYloXTHW5GmRugqCrYSmopjogBWK1MV
0/iW1MD0NOg6PAox6VxIXkfB79J+kF6hnMXO9snjtBzkKqwPhOhEvK0WZpUg4ey4bIAMOPWmXsfm
rUL4MX8m7UwaMweIymuYabZKd7SoWY1GveqIOY0lLHe1IGGzwb2lntcd2sQ/bAJo9j1W96eqvyCX
fIICCi47PBxHs+8YXDFJkGksEpQy87KGUIbiDxcAA3zEB3+F5YnlgdEhAvc5cSNzPYWRvS+NuYQm
pcoXVMUvbgBxkDAACzvDEvCphlet1St/o6HpfH4AMDfp+X0p/CQtmgVE0x0/YmIXbABSEOcWuiL0
Uvq9GthbyMgpDhhy2J3nVauZWe9N7Zyv7T2COdFA70rXWWIt/wg2vkdYvtvW90f8LFkhLhvZ1ndD
m7KojY302wQ2uV+Tdm4dmfr1vs03ZykkRrCy7l5lU/9b8CROSQ7aJNsGMSYPXZfojg3338kZ7FSG
ZQbDTMy8d0uoJDmJmXHs86sVgRek1AciqD9XHF+G39ss+Jvl/Mdm1vWKEGcGW5hv/HUm8Hs/lplj
6nJhdj8orrucdo6M1sv2Zin29tiedNFq2crtLpm7AVSqJcte55SMPRqiLPFGddIhoE8mbW8oaMtI
dHwyV1yVl96O0sdKSCeuHlqD87LgHV61iFGR3Mi60Jjzmqim2kOSnGMWBYBUCDbYQONAYmfJWV5v
qVb7lDHNfh3o99lkMqT6wTPdYjh3xk4O6eyCrb5CkLH824yL09wxZZA9g5yUDADIiQ5tdkGmqxF5
tuyn76YRnVUkw5S4fnhcSGiu/4lDMP1WBURcs4dTIvReBPf3VmOcob1PooyiLoKiaUakrNhMseSa
DEwu/S9CfNvXx+7SZ9i5ThYIZuZRxeWQ4mmXreklgPpzjspXsCholKYmev0Qq2phurebamDVf220
/RZ8VuMMdWo3c/2quzV/MPEWmfTOPnbvwB3CH4ZDe/2XFXWcziot6rdpFPBuG0OvHp7LDoE9pVlt
vfJqz9PDsBjzoj5fP63P8I0UbeidJKaTL4g12d+gw+PtRxCzep68RWrL1FQeA1pA3rTyOYmjmCgO
ZqF4nI4ALHmE1sRkktlPUwAPiT0Q2HePo0Er9SQ28uWve1h8H7LSgAH8z2vAKl+OW6WuK/nouoRd
8dNIVPkuJnr9ocBju8I4UonN6WwFtBe7DfgX/inuGSxMWOgu9iFE+e39JxYSfcLoJZpdWa/3ctQ/
DIsDoINj37LKnfnxMTi/3IWsody4pSzxiS7Exatkoc9ZaWwep/McsJ73pb7w4TBSafReGPkqkXdk
wD8HICYTNQEHZeHkDKlvxfbKO/rBfoIbUcO8m6j3lDvEpryZjBeKoqbYWVGJ6TQMWhJ2b2XvX+DU
hnY9LrmT6Pzhi0vOMcrXcA1lptyFDWOl9rwq6Ykge+qUK2bVb5vZFI5hv/PYywvQh5oSa6oHkwXe
T01VqFuDkTbxcIrmp4ohf8ksG2pQstnkc+9bxmOUPjVPHSRqUm7EGbK+BtAi0QOE3a5CJtCmGelH
IS00fNkcAGo6FJj1Siqx6hDptx6DK6ONG4azM+UktdxJkp66WEytSjRAXgO4vFVLSsq2ptyIo7TN
JLE5L8xukcBZPP3DZF1Op6J/OqwByGsCmvwhgpz8JtGWiUxIUjGpUG1l3mwbBBd9BM5fpofikOB2
zhPg4tgY5JYZHmuwY/+hrF17DZhvNxMOY0PsnDqqUKF7SZKFO2fyoNdXRQUjlCMfe/I6IFthbG8e
NISH4wDVzHGo+dVqbrw7lm5OWXA00SDOTmA88mfTgDAsjmI2XHSk1RMRQlNMS+JJY9Rf+MXp6I7d
TVu237/G2q3g+uTrr7BbwU+gVOVHVWBKkYwZrQs5yyNfZjzO89bCyU315VVCSQfRqymj76LreCAj
LNx33bHgYdDVAZ2xwWb79O5c8BD3w4V5xC0k10No1v4gb3W9rZ2WAbOP+/tJDcVa1HMQODUKlMLi
6ObkOzVL2VrK2K1IZRNfeQ3ywisvIF5xKD9IHwtemqFAbieueaXecda2xfwNld4fvGPC2EOQZsCa
IvP7ecRLWHwfYVhKJWcsB4fRm7FJMlr3b1xx4+k6F2NHEvpOzspV5T5AMK6fTUWxiBiDMKij3WFV
JrdabKqOO571o/mMP0bG+plWgvzUBDt8McilxwoMaM8KMwv0W5vs9aXY/wMzlfBhYozNqzva4h4l
SeJF0TnFlS0kzz3/7dymDVKRbVvtmTJq9NM5xolF/jlE0IfshaPliKYPYVTd9cuAz7fPEHnBOP7e
cRpjznkXmThPu9LQlHtvRbwMkFjR0Hqh1S9swOeUpd8Jf+8Q+4Bjsm/NdWClOjeiAEyYFvdxB7Y9
YAVOFuy4X/PR7klS9M/bYNp8waOl97lcvxrdDrjSTOgPqpcbYQtBNsKXpWGzD16nBzuVrOpAvEP/
tTsKL6OsQ7/Qb7yVKQMPIHHxiSV/mhjOugTYMX7v2xhkgliCJBUs4iBzfU9sh1fYF/eRCEAFtRQm
agw9yL3hlXPNOUcw6Jo4d86NRhi8mGgi3GyV+nGABCYjehEoF5hdbDtFlFCq0T/ZLpL+TkFSlMOj
M74kppR/3HuDp6cQCvwvNeiKqflugqjBf7JicLonBtCg676JjfM5rQRob4dImkCNgPWRfA==
`protect end_protected
