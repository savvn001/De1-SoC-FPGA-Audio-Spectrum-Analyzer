��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�u����(";k���{�d7n�3o��J�I��7���Wa��St��7-B�9!�T��rg�LD���a�)G�~"�ieנeuC�z�{�,��bD�#���)@�(���ME��p4$�M�F�~�����������Od�.`P���?��sQ�Ӗ�Nd'�æ�������o�k�^�L+?¥5q�͹�)Z:"LfP�IG�3?)�ӳ��)�@wV�Lq=I2�o)��
w�o�����5���J��#q��}4��/��C�_>����<�G��-�${TzZ��g|wK���j�U�#!&4���rSr�p
�����Iu�N��v�e�j��`:�{GF�vqPʞw!	��m���V�&(Y}�ʺ�^�H��A}��e��S[m�������8:OXl��+�vW	5/(X'�tO����`K(2Ob�U>z�F ���X����� �v������s`������է��3�ӞO�V�k,�m��V�#�|��;p x�����ѯ�b�F��ouFTA<Ʒ������(�j*�� �nn��M
�7k�lY�f���'��I�3��
n?�
���u@����O�����=��[T���e�z
80�l����R�m��?�~"tHz�ʽ�NQs�r:�H�{��f�e$�}�ׇ��;��=N��,��v�٪��(���Y�����?�Tx��*k��Z?�������9X:���sm��5���EO��}�M��E�pgb��� ��bPd��"��I��~���z6� F�M�H��%�h	3d���Y���� �W��Y�M�����wL��R�n��5]ok���e����� �t�Y�;vq%`���oeTF>GAM�~��D&q.ޚ��G��za����L�6���0n���#�F?�
rą�%���F�p���0�2���-5V�/22|�H�]�`<5|��𼛀P�'!�l���䯄xn�����D���년��l�ډN�D� �&hP3�/4oC[�c��:����d����X�w�z:5��w�3�2��]3�k���_�Y_���h-L(#�tA�c���c��̪�jS���X���`�G9����'`�<��ղ5��.�(���c��>Y� �1#���ØB?��I��x�7����wq	�K�뉧��E]����e�0��HN�B�	s�3���2���T�n4���"���P�0u�b�ƿ��2�趡�~���^����s�`�<�QЊOQ�r��e��b�R?�T��o[}��An����@,�O]t�DG�&�4�w�4xġ�N����������r׹�Mm*�s�}u0�\�L�=��]Fk����Z)Nò�M\�h���r{��
ϒw��W6MԴ��Ӯ?�����(v�ݧkʁ\�8F�q>�v�r����Wc,;S|�7"�`G�&C*N
i��q�`�|�̏KA+�glfl���[���^����"u�/i-ڝ�1n?��O�I�zP��:�������>s���=�O
W��y�����6�2A~��b��B�#C|BU+��]e���`�w��n�v�ٜ�s*/pL~ �0�&��Hص�?1�O{��u����k6�&�˓��A�_y�י�,U��O:)��#�%���D��`���*X_���/�O�N�_:����=��)�I��[Q��/�|AG*!���Ss�U'e�em�IB��':�B�gp���IDuu9�
5��0q^Ds�ۧH�4(i[�Q�s>��R���_���K4�lU�q���A�
�bLp��|o/ZQ3ļW���]1'���������K�|�NC����?�_%;r #+y�V�[��ߴW�[�}TO��?���Ez\;�n���#��+�(�MK�][8��w�^�dB0��Ywr�!`
�*"qH��Ev���5���bS��9r�}��nAX_E��bL;4u�{��Q|�`��^�D$�y�2��V���� �]R]�C�+1�r�1Ήa'C��VF��.���*"�X*���1E���:|���B������'�
ASj�Py�@U�%H>?<h%F��>�F�#��y�D�Z�̀�	�����IP�?�+)K��c�O�o*Z�|F��;Z {��SZ�+��^<=��Yύ��p���y|՞S�~z*]聥7vR-L��%�ڣ����o�S	)9��ہ�|�����R5)o��鼴v= ��%��Zb�ϩ.�U]�q�<%V��̆�.��Z�fY�����O��s�5��Oo�c3�D�agѐ�
]�6�%����L0�|������'��1�D{��Y�&�T!����U��J�L��'߇���X;,��)�[}�3�!8w��`��m���{�*�.�q{3QI��-�=،l۔��!>���sqm�����.�F�Y�,�yT�u5O��٣(tBo!47���uu��b����D�����pɧ�uI�8�v� �ddNҢ�2"TX�އz@kj��0驹%���}	�C��>L��?T�B[q͋t�@<�c+��b+�D���U��:J�_�aM��Qq�wP�'����Z,o+I��~�a�>�m�p�&L"D��`���))�c�Et���N6���p��C'J#�c������7����7��Y(;{�^DM�x*o�>uJ ş�/H����%��ؘn9!ֺ?Ƶ��!���YPDL�ຽ�-��n>�w� �c�g�u"$�>_���42��'��; +���9���^[���2�f����n����E rfT�SXy2�6����%k,庱�E<'�]��1F�_n)�D��9Lk5��� �i%:��e��&t�ӛ��w��3z��02��'�QС�^?��0O�~@|�&��P���6��',$<�ƿ,. /.���@{��e&qH�Fц��5<C�n!�O�zq	V@M�����G��W��6���O�D��ʻ_n9�����C�|k\�Jo?���Yf*�WW7�/�F�Ī5�/|��#]��ft6���Έ�beA����p��&,p:o"
��K�!��L�71<ز���n�\ҦJ��vb�ȝsԂK��g�-��?�_�������]5�.�� �a"�k��X������4]���N��j���"���`���9������&�jE����1�TY�e��҂;&bʑ�ɝP,�SRӗ��g�Wk���ӆe�3�T�͐������|�2a��x��ڠ�E-sb�E*u��z������p	�ՙɼxM�0ݘ1(�c�plc�B�X��Ī�k�,t,��/L-�CB�[��	VHqW�EҮ��n^��.��6�&`);�E���͸�3���n-< wk�ݒo�\��ɹM���'�4�}�6�����K�!�Υxr�@O�&���f�~�lP�`��9��9O@Q�r
���qmrP�:b����eÌ�\g�NG��,.���H+Zf����l�\���M���נ��H\޶�����8M��1(M@FQ~(��˙hBT��-ں�q��B���U�sĎ�G�;����{������������g(�튕Y����T��X>��7��[�}����b��M�d{x�������7lx�3�I�\s/��Y�M��b��4ƀl����&e�W��Xm��h/���%L���@��1`4������o�
ݍ7sް�#���v�*�euCs#%Wa�^Pt�����2]"���Ʉ���4�%6d&L68� j�[:<��<�!ϲh��'��t������Ђr4Ⲓ:*����(j���H�">�ڭ��n�<������ �|�?WI�s$��r�z����z&t��32\?{���K%4 K݅o�cR��9aa��]��K�d^@ny�#�����E܁�D��WA#�Ե),�咉�����0����[��d�LU���4\�q8��,V��#<��dVc��4�Fhx<�C�8
���[�u�eE�$3��d�9��Qի}dm��%TUؕ��p$�';p{{�xc��3�� ��/��:��9'���k�b2�<F]�W�l3vtM��x6��D<"�|]��۩��dT:�kg Zsd�e&�%`)7����X�FȒqh��e#Gތϵ/�I�XR�=��)���hrI��(��|�'��,� ����-��M@��'jF���Z���m�@�֗v-�
SA.�����ƚU)'�� �M�ͰB�H8�Lw;��>�>�(���Z�-e2s��<ot�N��_��Lŝ�t+7|S�lƪ�eڐ
��Gx� F	�u����p2ka��b��P|���>��_������ A1X�Uy��S����
��a/��W�<w���o�ok.�5�$�E�@�(J�)]Ks��ǰ�E<��6���}�Q���~��q5U��ޗ���6���s�7Kd�cVB���B-[}Ҽ�/N����F���;�������_��G��3�IGt�(��}��J.��$:�(�(��y��䁉n�6n���K�=6�x�u�=$Lg��*��D�����II�;��D#��!��f~���n44:rO�0�)��[]�<
�_��W��V++�|�'�l�4I�%/�����[ڦ9kTm����-9�@�&���^�)�6�~3�<���2.�3�Ĝ��H��ʵ�]���ni/V�.���i4M������$'�<[&�(eQ�Qx�*�b,��ݔc9�;����H%j��S1�k	�`̟r�7|�C4�%���CE�\��;}�J��3J8��Ex ���TD���FB�ц;�����܆U��T��k��!jL%?卧�� wM��3���
Zf\9�*}�tP��.��k���N8j�&�Vr�?pä�����Q�y���s��CVH�Tlm߃ޤD�m��(�/~�(�\Y�o\o�e�<SO/�Eᠥ�%�����s9�g���݀�s�g�C�&��f�$����q=J%���`�ݯ��{� P�hM���N$�H
����74jE�fO�������/��6��B�S��]�-&��B�j��W���W~m5�Nr�L�:��t�;Y�=�s�hl3nk7�gnw���Q;̔��-ޠ/��6(\D�ٶ�<:-O�d7�aQ��DA�#W�$��#�+~r�L��E� �?�ԡOa5׎�-@w]�tm�}��8th^��s3A�F����IQ76{.y�<�_�b ��%�{G��m�������ោPum<�+7�U98K�Wq�}U�$)�tګpf�[%,(8�=�!�*�+�4�r��de'�+�lN�0d�p�����R����q���
<�;BL��1����`$,��٨��w��VZj޷�X�xJ�Ք�m>�z��_.2Ҽ"@M{���6Je�)r�_O�/�J��i��g�F��(��U$��� F�[lV�Kw�>O��	�v�6#�V.ŷ�4�x;����n6�y�����a��@8���+����2r��$ <�cIdm�{'k�@�&�W[a/�p��ٖ�Z��Q1M`�[��o�<s��ɍ$p�W)d҆��벞t�Q��3�^�pC:����-���H�W��M7�O6��IY�f�;� ������f��az��ܩ��9/�!I�mx��7�BqtKj@;����ç=�X��7��r���`��#)�#�,�C��$�*
7c�Uv�"�/�bm�C��M�/LÜ�jG�Y�q����s���q� �
f\��J�^��#�v8=���i#���A#����\"�x]ی�0ɤ����	"���^�Az�?"��q����K۽�*ί���3�ZC��{����_���[�8Cd6̨���^��w�q��3 �<x�I�C�v���z�pv��;.����f�#�^�?j�F�7S���!գ�{�Ȱ�,�f'�ZζDQ��{$��5��ׁ�Xg-����cj9�I��Ƙ�WӉ�&�")$��k=��]'/�Q��}�.h5�".�9n�}�_�\տ~�j�H�4�{��tO9'��:��ˠ12��o^��;��<P�O,V���T�nj-�P�v6B�#pp�͖<L�2K	��i��
�����8�����F�?zх�|�*|܏���[F�	s�<`��bG����b����WxSo���e&�RpY��x8BфJ��4x�sh�񛄤k��%����7�gS�9�U(}İ��-2�{{az���Y�]�I��y�"(��;d��{)�U�2�j�<_�gc,]
���r}���
��]��e�Z���z�إϦ"�_�G=5X[��O !���{l�ˏ��	JX�)����ȘŶp�t�kbd���֚��  ,��jQ?�Ҙ8l���K���ez�A��������pV�R���еՊ���-+m���_i)���� �����	�V�J�ՔK%@b�?��m���R�<Kw�� �}��(H�'л�䔳oz�����J��qݴ�2��Lo�~v���հ��1
��9�K���D��֠���+Y��A�Fa0T�8�Z�DD/�N�U?�P?op~�k�F+R�^map6*����I`8�u��V�X�{?�Y��$MG������C���e���{�dߘG8�~c��jJ^�&��4]�T�9Du�����c Y��RA\��ޱâ||��ׁʟ+�'���kx��L����|f���j�-��N����ʰF���z �\�nVP�%G�Q�&'A����/��q�,"M檳��D`���$Q�k�$S�8�pds��\�A�������q�|T�����6�U��"��9��d@H�ڶǔ�����M毽"��1�RM����軩�3�P%���6�\�¼��]t/�u���"}i�jQ���w�R֋�P'm��8c����9���s0$#��j�
���$n�d|�F⑅�^�Wj_:G��;s�	L��!�m�@�z�;�)n��J�51�¬J���W�ׂ� h O���́�M�B�r�2ל5��2��`H-�DȬ���P\�.x#��}�"K��`۶~������]TF724s;{[C�oo�$���d�4������������^�ж���!�����d/l7Ft'=#�U�[����H�w'�."���V�x[��,�!����G|�b_mmp��!;DG}���O��*�$b���$�����Q�[>B��&,�S5�P��=A��%bn�a˷��֧x�K��r�/s�u�W���E3q��Y]�s)�,7���񍑜lw`v��`���jX����Î�} :���{X��L��Z'�ڋ���}����j���`�m��?�=�8\A{�)u�i�Ϻ��̓I����"�8��+��y�T�x8�kcUk��g9	��ƻ����q������>N-�A&��'P���i*����Љ�M�ek~`�M�cu)��[��/��$I�P���[a����M������K��e>���ԯ��6���KVe����V�c�i���@�����d�m����j�H�2�g�&v���0"d�d����7��O�������3�ݎG>i�)�iЦW�sz��ŲaI������7Ӻ�Ew��N}��R x�S�v���cM��$
�yb����d�>�	Tb�n���x�{;U�2R����2�U%}ȩ'���a��s�]��t_ϊ��K�}��K�81f�V������� �B4_�;���������I�Fn�#�D-H����x�����q�Cd\wA�a��a���)C8'd���-Kb8X̦G]��f�0�����b;�������N�X����"So`��O勷	 A����6��$O@�n�q�>�D[�s�U�C�T�M��%��sQrzN���Vq�i��z?��?���1��cd����t�I�9:	�J6����W_�I&R:�?�D���'qW>��n�%#�J���V��'8h�N��N�Y8�Ù��9�b&�6K�
�JOTLp��ڼ.e!
�yB}�2�\fǯ*�.�9�]��B�l��O*��b�D�\XY�s�ۄ���Bܘ;(z���8��S7�G��1 t0D�`T�r $G\�L9Ej�9�Ӵ�u����.���-����f�w�� �)暛��G�����-���ek�%P��:T\�>���6�	�09	F��dϒ$k߯W��M�E�^�����B����	to��
��Q�l톼���}�1o�����K�W�Z�@i}}�JL�FV���Z0�j�p�|g�֜4��k�i������W�G���\!�ж`�AY׸�p�ʇܖ~7N�v�R�d�W����&\$���U��)����L��ԍlb*2~��X����I�Y�Q&��mtv0]��D�`PO]���)8W������h����9�`����c�W'�
�?��>Ghk��*)�2{�|���nG)��L} ��]LJ�-�Pw_�j���A� ��f���{�n�n�'�7����G���u�� ��>�2B��G���
�"�,6 HKN<���l��h��͎7��m�Ǚ��J��Sܗ G�]�K�^�p���� �Q�{��N���+2�/��(�=�l%���2O0��O���õ�/��^���l���6�v�o���7�r���+��-ף	��v�D�خzJ�el��x�`��n>�C�ks�d����"g�R��S#т:����/X�4�i��́�gBM	X���BH�`�6*'�N��]H.��8�LX'oJ�&
>4��|�a=[(LK�=�[2�9������rNg'�|5WV�s�ߐv�8�FL%�QF�ʖ�x��vA��o���m�QM�E��y h�<;5H#ml��>�B��"m:R��q�� ���nI:��Pe�׏d���
ѫC{0��on�DN���º�Wo�N�m������.���D�vr� �Pq1v����֐�DF��+6�]����!��ӼG�+t��I�8km���>�r�1�JsP�w�*�	2��>�B�yh���S
�6��{Pݡt�T|*�u���@��)��s�߄��<s�3���v=MD�v�e�L�ifb�X�P@o���>]IF������e=���M�v��$������@�bJrc ��[�e$��R_�/�!.��$)��������U��ѐ2�s؍/�B�g�F����hJO�P����<���E�g�1�[=f�+���T��*CQ�(04�y',�ɍ�ژ����e�}��r�5�K���h%V,%9�w��c��c�����u
����$0�/��G�j�����D?s�v� Q��Q��x����6�H��M���g��G��"湴��l��i��_�-�2�F�J&?��pޗ�ŉ�:,Xc�z�pygZ}�o/�
y��O�����+cڥ���e�8�:I}�P���n^̲�t0�0ռ�Vl�H�Z���H�)6�|�	[���|�wc'�/� �$g��b�S�Cp<ա���΄�_�GgY�6�l�����J
~��O�����0{
V�gT�������&�G�8��Ta�̬�F�+X�Xs�aR�z%�B�+����g�\26
	�hãP���z���3+$TXǅ����En��ҭ�b����f6�[ n��Ŀ��w>?[4��ƅ:װJ�:�4E�LVhd-Y�����4$���g"瑐��xB���"�1��ϻc�P��C�.���V���W]��4aLG�R��ָ���a��bڳ*�2�����m����ok�-��Gd���=���'.�~HLK󪯕�
����h�Z�/������;ڌ�9o�ƑB�T�M걠j�+�vY$Xtɣ��@��� ���ׂ�(��Ր�4�+%��sh�Q�Õ<�)�����ƽ�dyF���*��!{H�y�L�|����'��xN�����D!�F��8n�d�rY��{���\��-���:��e���s�`[�J�r�wF_�U_�s
�f��OHp��������D�I��:Mk�/H�/����_����4������4�^�Z����S@f��~��EZ�[;M�[�