��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	뎊�ִ�\ymf65�k�{X'|��J � *vc�ș��sV�O��P"|�����G��4�F�?o�7�5���T����n8M x�	X� Kb����a�C��Y	F�F�e�	�eqPH^xI,�tK(����������O&�S����Cv`��n���m
�Bħ���P.X�	���������Up͝q�:��a���k�X'�N1��9Tp���
@�M9�;[����*���Z��a�V"�����!�*j~MVR����tE���A-��-�N\à���A}oI-��O��BY��>���F2A�Zj%A�s�Y[xG��L�OҒ��_����ύ�݀��>5�|�u��Έ=�0�TZ�>����l��ľ��K�jF���`����r�S���2.�~wh�>�:~�Yq����o~�n}�H����c���JCP\v�A�<H�S���݆)�}MW��5٠b"�w7޳�}^(��h�'�~x�u4��j�9W�e�<[��b�pJ�0K{��e%�D����(|�A^�S��_ a[���Js�)�V��]��e���Ҿ&<|�Z�֐�
l���c�V�����m�q�N�ܭ���6�O�qKD����*3��w��~��7�,nGgnǩǢDR�-&�;��vXƬ��v��!�����L��×~�s���߸4�~ҧ��IB���߀���h,���c���^/ߥ}�����z�s��c�N}�5[�qx�H��m�p�� �*B���qK�V�� Z�:h�@��q����>�ïE�W�1{$A�3�&��Y�;� �$>�ѷk�Q�x�Dr1',oq�S�7����3)^�v����zE�gZ��D�٦��J9T�e���m���l`�~�3&��93]�F��쭤��z(4j"����l�٢�l��:Y��j������Pc)�d��5Td#���3Yk��g����_O\��V�O;N4���N`���>�¿����x,���������tT�KQ�Ō�;nG��TI���4�E�˹�b�$D>��%�x��)W�6
E�{y�D��}6����d��$�]�}�u�;؁K��U+�Z-��`�J���16��<�`��E��ev�@З��������x}9�Ae�/�nYM�r/^�L��ex6|W(�ƷLw���7
c@���{�:�r�����B�fa��դb*M� �Mb����D�뵕�N�fab!e�����a.�hD�x�G"� w�G��qc�4w?��&MJt�O�X&M����Et��iK�7��M:���Wxwa���"KM����������|�O��kh>�p�!|�T�'f� =��@[b�*�2}2<���1��l��9l��A����Bǻ滀�Yb�!�X^����J�P�Pa�ԺV�;��<T��8*я��U��8{����S�y��Ǳ�����	.�]���TF�Z�U3�q)�-�I���g�