��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	G&7~�?2[@�x���"|�h{������官��j�܂�����j�إ��i����E� iW��8G�~[�.Cs�+-���D�x�Z��RTY,�t�3-�wi9g�-�ȟ\�m'*�~v�o'�x�k&"�'��-�ү���A��;6��[��K�aF~��������(�ȅ
<������]l�tkWҟU�ށ5�C��W𔨼�h������t��Ji~�1���F�Ł��eS��y��w�
�t^�>�u��x���1���!A��gK�IDhe�9Y6H�?/���I��#T���M�CE�#=l�%[���E tݎRH 4X���[��XGv�.g鮈2%�-R
�4q,�ly���۵.��ɹ���9F�4����-�a���pb�� ��3/��!
�	f3&d0��䈈#���t���&\��IG��
vm�l��w�PQP �No�������π&}h�+�4��0o��� �W��3B���9���9�c1+�	|X�a?�:"ǖ�E���v^q���+�
Zl��Ohu.-&��V;U�����S����[�nѼŇ�3�,�X���&qz�@5jq��&h��C1����9�rn����_Ϥ�=��J��?+���J6|��rd�@��U�Y%�,��w�q2���ĩڳ�Qތ�6���ף�-Q ��_as������Tܨ��5s���8�T��#��	�p�F�{�iN��X���8�w����j+�4�E���Ѐ�����@9�T��(�m��bd�	#����4\Hmi~�d�e!�r��%�y2H��c;�y���"����Fd�[��\?]�"���7��-�Y�i��>�s�����h�ng{��k��c��%`�7�\�d���mY��w�g�x���ȝ���������5�||��b���E��5�����i#k�᫼��/f��Z���@�(.n	%`=�z���$@~�{���Ǜ�S~vSd�dzx�i�C:0L.P�K,x�4/(* ��ƈ~>�C���Uv�Iő��8��͏��x@Iz��W3�G�@����
���z��]�nt�Hn'�r�?��i���cCAg��� 쇧�c��i>ū[g}� ��H��+�d=�A�c`��~��rO ���R�m4�ܨ�%D�����ùd�� ��w8h���ra!�=1)bl�e몱1lF�ȇ�s�,�v|�K-��n�b0�^{�Jm+�%�B�j�wW`1��8ҌG�7��<줨��:#��}�w��P�����rDގ���{��?�"��Q�x+��-��#u�|U��Ό`C�zn��UW���>������r�4r��#�
�^j��:��[k�#t�t~�#��Cr�:�/���L��,���YҴ'+/�p��J��&�EY+���P)X�2 �kf�z:1�5j	����컜�;�>:rv��������t��K�A�83����n�4��������:VS�XDDD�c�x0AN�g_�)P�|,�w ��p�'�	;�nr�H�=vh�?[tv���b
W~���#!�O �U�����?��Q���pv���3a�lee�I�`Ĥ<�r����Ӗ{�Sס���k��qˠ��W��L��o�H����3z�ݢj�XM7$~RFz
䔉g dԃm%�Ó��&�w�j�t� Wp�K�
JO��Y��Q�am���Q�&>���:I"�	��&�'5�!�����En;5�F8J��ǞDd�Ԍ�8.ݍ�:�;�Nض=���la��~���aAE�c��l��+DnO��P�K��O��Z�&+[H5=�`%�c9Ȱ�*L�����4�4G�ޠ� �Ƃѭ���±x��h�ug��IБ�vn��A Q>��L��J�/��X���gi���>j��BX谩{,�-�[fks҅��Z񔀲`��O��F:�5�%f�z���56跮�����o��E�z��c-��,䗚9�Č�+w\^�@_&�[g~�KI��:zB�@U�[Tč����0��&ؾ����T� X�9b�ɕ�O���2Aj�_ӎ�}%NbʋY��P�2�?�,��ש_�����NYC� ;|���-u��� �2������?�	�� �u��hٛ��rw�����Y�$8CP.��>Q��ճ��O�E������\�,�-n�ɜɂS����K>���3�c�i>���HG6�	�=gV"O�ֵ�u F.���X�-��E��։�%>��=e���kg[������`ghb�BoA���-�p-\6�｝����<���]�m25@-B�,9q�����0�Mq�����<��\+��\Ģ4��i�+(����� ����.i�k\~i���L\ ��j������zJ>�;�i/FT��h86�hktOQ�nR��V��+P��?���8Q���~�65V��8�0ݟ7,|��<��e��6�����(%g*%�2M�F�f�^f��Yf�x$~{j��î#ҟ�Aիj�A�Cނ�? ��Z�����Eǲ'��0�#��,vnE�M�{G�YQr��E��Z3'���fp�[�]�v�z�̳���s����_�48��o���ZDJ�)dk�(�p��]MgQuo�w�v|I(a��:��Vι�)o+���/"�)h�G�-�$��6��TsB��a�념��w�����4Qr���o��	���~�Jg>ZTb�Ѩ���Eu'��D��D��}R���t�������O�<��✛{���h�N���H�u�F4��1�Q���Q���G��|�i��Tn�z�jT�u��M��n8���~hȷI��P��qǌ���� CDy�M�>6T�[�ˤ�7�o�0*R$�R�ji\�M�>���r9�t�M�����ieX�2|�Xh���]�](˺��r����*�HV+�FU���'�s ������̿~�7�@��8lw��!$�J�Hez�.J�W�ۀ\g�]
,gn�U�����
�qj!:]/�p��,���P1#��Io_'�P���u��w�`:�uE'�@�j���g���<y�<��n�NJ�����!��>&�>7ðf�H�`��'c�(:'�_�ߓ��#��j�ehL�(c�'��j���
Z��Kr�5�V�Kxb�j3q T��\bZk�[���}����D�h�pF2��V��qSC��9V��J@b�J%�L�	��n$��P�K�5KLb.�9e	D�8�zN���Ҟ��rU�� �:����a!�&�7�$�E�݀���9��� ���Q5!X�[�8jH��4�ot&�z\��z�	%�O"7�E��V�j.�80���pݯ�������o��zN�p� s�����a�$&�4�b����l�h4��k;i�;�{���k����L�́v��Ո�J����p}�yZ�w�VsC	c9p(\���vkZND/�X��9eU[%�cS}7Z�)q��J���aa�0#9+2����	�D/��N�t/��]Ps������U5��GDRU|����2MiHT���''� �����쭷�U5.���`�xn�� R��G���W���:��\Bi�r�պ[~���"d�;53����<PO�#��V4;������1ܓ-����{��~az@�B4�pÿ�y��X	RҘ8�.8~#�9�Ԕ%����t%W�DSa�zK-��*��=����ɚ�0��ې��^>����`���d�cA�!���d�Z���>E�K\�AX����z�B�<I�!\|��]�_YV�E��"�U6��V��6������i�7�Ynl����}��#�C�g�p�R0Z��^���6�T9��cVCd�>�g��5��V�;���ؚ�������~�h:�kMy�~������+7��SCw�@a�I�+�A�{���8����,j�!؊����S�����]��NF��y�Ƹ��:���m���j�#��q�[�6�Ѓ,�
S�C�%4l�Kŀ�G��]*���Kl+�ˌ9��,��G:�>ۤd@�(K��1-@%J�P����6���Ǥ�fQj��h�F-���C.�ݯ�_��seNC��d8+�9i7��(��i�f�P�٫���ݯHn"S�[&��ۡ�k=�s�
��,0"�u�V�+����V���?�u f8��Gݕ�˭�dO2<����]P�|�CY��"����S%a䘻CpusOG'鈄�}<�{���ݦ���id�((�] �q%%��ϼm�� 7�[U4'#<��O�9	`9%���Q�E�S2أ�+�#R�P��7�- ܍ʚ��r�A	ָE�ᚔ|���gF�c�78��Ǐi)�9b��0Vyh�#������7��ڇ���ʑ���D`�- wP��N�`۸�?!�Zf��x��¢(�z
�	ĵ��<eA��^�(���UPb2�d2�d�ע�۠1�bV= �ҷ��Ms綬L��G���K0�l�[ 3�i38��|R2{ML9�G����u-Bҙ,�qR+���7����#�58�v�_e���4�}/7���� #����p�)lf%��buKC6�Y��d=�Yl1},��8A+[�J(�+�E�R;Rl� q���3�-f���֜���~�