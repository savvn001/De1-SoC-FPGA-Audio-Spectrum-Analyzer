-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
c7lHqfr2/BZlZ0Cm0/BVxCRo9SwuCkaSwh/F9B4tmdlIOTdxD0R+nZWBlhv4LGb37YnBXOm6dpyW
g6VbafPxoF+pPsJlEZNIwVAnB1ZHskPHK2nVaejAELdPXOjJzzUsjTlAjA2ef49G18K8QmQrkUfE
togLw5zAou76uXAye9Km5nQW5EScd1HQVfqUBTCgcS/+CaC4d95dWQuFIMCACpd9BWQyOrm+Gs+z
ZTIjtF1+rQeqlwK33nU3NZ2IgpsCLPqvT5s32eb6b8Cxe1HjB82OZTLYq/iA+Lbw17o8h3fFG4oI
sSBQwvCQb7c6DCsexr4kPzmxTowKkXgUBmwCyQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
X7x2j/bm4uC7aKQWMT0XnNRmuMpolLR6X5WhneiIPIMo/hamI+LY/Fle5S0fwsTaOIy99e+lz2V3
yAo2NDO/Dum9k6+ET4gfcz8NAKIXaVKKSzFkKVWVH6l2d2MCniL5IuUJ+uNQuPk3R7gwAGTXl49J
qMnli1UcX+bSYzw3X4y2960P0nvTPgjTZzny7MzWUN60tkpZRH1+p7sGDbmHaja5uHpjp34xc+ui
SrNSx1wBsWQ5F3dNwTin9qzpeELOuzOZSdyuxC9q13ohtdEM2hK1dwPo8OyyamaL3GeTHjtXJCqq
YHLcWN06d2mPIZQGsrck42wjW+MYYRKfhlcmYQKsnKjXB1EsTnChZW/kA1RiIN1fOMx9HIliAe+5
x9vQLrwn4jy6o+v9t44RilgHn44w5stOKRQf5blJXaf6xEmey8DPAIv8+C9KlFEUQcoqF3yB7232
woYOtPry134csMiw9buIas9g4cJYgV0PBpdTdIEDyY/5eivzqQKAhSKCegHFQYKxXbaDry2BpdWr
fVtCmf8LbHp/QkqROMuWH2np4Owd+lw4ACIuhZdcolBFcbDlrLbNsbDSbGIrcNExv4IVhYdbUJtu
o4sJezMD2KhX6rbIbCsG8hgqvS3KrnjH9RlyEtTtjpnspxK9A6YUsM/Qa2vIktPFCD2psJ2bRKC3
6RHWD2tyu+jzHfr0DaOh7vjAsGbkA7SaQx9E7EjGaflPD3nphWTJdVOfXr+k/ATT4/2I1hkmCu99
VO9uW4CmXDqbUmPG04KsCrnPKjLXx1Xr+BSHAEvOepTMqxTuifCM5SSbz6J6kjeb/Y4yMHyinNSH
bv/amdZ9H+VVA32u7H1/xaady/F4JCHBtLGWnzK55+Tcs49fMZwYCaqVnyRwu1dmJ7EnAzKFJ/Yk
aXKhSOPmfG/+S6zDGmTIWP8uTC1P6mvlnpuy2Xj4eTU6IS3WBb8gzp+BBvvOcGyeOHQr/mumnrvf
WrMbHkDVHXcBzn6bUSJCTQouP1Jk9EdNxmtPvi35NH2a6zlOwNIqkvMgIy1joT5SRSmvtSnMcfPi
byTVqWWw+GE9g2mK9ApO9ZQCK04kWfVo+hEJOSKt0GqLt2JS+UG3qSYCa1zNBG1GtlmqP6bGFT43
s9nWZS8V0tAeCd7Kuq5aapGh3Of7MvCCk9YToRbeO2POt+p0G1mfnIHapx/gQfpOYgu5RvfGorJ3
bqUhPXrMZojrhXqUKjaUJrCryMvUs3V5EJAFOpNPzCUC0/CxViT9daJEycDk9IQmuj65FKjazstl
vDrpehUQRlzQUqTTTnZqkVlM23PGY44wrCgTpcd7XAZrwo471Rprs59LCeWh6p/zOPqnHtwbFEFn
XCj0eJPRxt2dYIvORCjrVaDPUDTY0sckyttgATpqAeX7WDGdTzf49WsM/ziXhmxJrEQgioaZU+eZ
6dmS3cjVlH3Zs4Ck0mGLx+HywiOpRQJeGDGdcHFoFSWbPu4AbXOh9RzSI393dMIY72dB71Beva3j
5d2bzJxSJxR9/OHmyqWi1jQrggFvGodohY+fERxNHL4FVvv2kn+GJOB+l1KjqMy2NpoOefSgDHWp
Dt16AoEvmrYmcM9ZBhidhXq7iM7+fqxuuWq+pCHM/hnZA1aI5Z6mHRvyT9U7P8IkZ0/VdazqZl8l
G6qZtYe6wSddJJkunCbM6g0kmdHUZhUI8nglSG3cIYphowhkYQY/eoWPps8byOi8yyOuOU74Ma2L
aKfwd9xGCa56l5AjZW+oLle01N/GEibZ+NC4KF0bQMaNprNYyPUdt4OvNJuQwcltMRTOB/eC2lUo
RcFAIm09tulqu4J7iwpvIkG/sjVoEYOBgH2uX3u5y3lGaohzvgcUyYHusno/rz9PQSoi48/6QfDu
SuLD357ZPVPkTmpTvxDAGo7M9cf0OP+thJAsi+tJH4/WKhKA0VTgoAM0pdfnSNhEbo7dduAFMAW4
ScLPCsRck8a/dS5x75WlgcwKpF4DAXJsPKhReBL8MO3OQYJAxIp8/Z75ViK6Sqpf7DMy/ii+aVzb
F2TSdPOTVwBzZQY7b3jYfO3XZ2IHmQ3c+rHwZN0SUBHoqcuZNsI6OjdaH6JcAfw7DUA00n5bI6Or
YDkTKPeTw0GKdjhndA56QGGVoXPwyu5inRlOd4Q+UcgYNBuf1NCpWO98tVLyGgSv/qcyO0vSFQYc
rWFD2lWcGTTlRQ1LFRKh+0FAvp+F1wMV/fug6c1EfGlnO/fIu/wcS/p+zw652CAAuoQMUZgYpP1o
QOVRkV//yoQ1cVdHIbYKA/J40dCBZRnuoAWLoHezLAlsY81UtZeB7YrbxHgd9g/pq1QJW5o+VpLm
9aNGOrcIlXo0dCf1nMJnFz8kpdJmya/cIoheQ2qhgkE2V7xbPVxV24+Jxig7F+uv/LgBaRodDB9e
wRVpHKcVK5HORMHIWHNkvCZDKCvJhsonro7REqjmzaBDstvKy91T7OGLu4kDFihI4NBzryFQR8Eq
jCsBtid18PqsTidNXEtw/F1Pj+2ONArLlGzwiaa+ZB+wLDIWnFtAyt3Q3FNSY7I9Q89HXwlKXiNl
f+w2eB0VMJLw/uJA/NLdSG3/pNucl+nJO7wfP2civSwXtri+okMqfHqDogMWATxaq/miIDZnnpAg
K9Tji4Z5nHYG5KtIoOH7GsxW+DL/7Vxmbh1erNloZd1+wlDJpXBvFdEjdtI8KcPtvY58zBz3E+54
OfbkpcYAV7pKPgqP/+fXnfgKdB+IaRHAKlpkuPvmCnjBq18PzbF0oRfOuxoQLtvcuudAzn/65CPp
29EoYdZu58egBO7xqnSJmQ7jTjUg83NgLSJCvBs8EisMoM4E1Cx6yziqZNXFIcAMmnwo8tuuRGm+
lL3T1clJ8vR/6zjVPT4yawdBnQ7hkH597vc7u4eGFL62GMaY7cF01eOm2fWxzqxi1msPNd37f7q4
OutJ9BTeBKDuxYkJK/sJfXpond7QX7mFhLUjchGzZ4rRgq8PAqdeOdEdxFtwobzQPExfzdtH8kVK
dJErQ7kdZqWwz5N6apwrUk+B2WNa2tzV8U5/BtNDZXrujqUaAhRHcJC8+CUfNxQ/BuJb2ampaW+f
Y+Sfljs7TOWXTKmWldsWVnMkQg7rHfjqbsJcC3Z4PLT9nOD+hqisAKsTmqT103osBwaKOqXl8wIt
1h4EVoL5c3H9z+dCVI8tbvlvGwbWje+QMfex671/JJBe/GXXsK0iB/A4ygw3MlS9Sv9CahtXitx1
o29TosFR8kiz5e0WGnTSJCa77pTBazVib7SKzyBcTLD+8yLmGQSONWCqmuo2VMA1364w8JnxaOXS
4E5PD7/KlNfU91izElyA9Kv3iHqbWPcU6Pdz+Sx3EuaR+EhLkszPWRUjlNiiQGJGsvEqWbTP9a2P
d1MHH2ucb1vQyiXzWo9P+tB07hfczVy4rad3xI37NpKpPhtBIT3fQiNg+J/4L9PFP1/Q6d+FMDhA
inhNGEyIhlFuXmkEuZa/qWPYpR0QaXhnHs2ZAxpJG6ITdGETfwJLjBcE9CPc49zfilV5rywpkvA5
Mzp4p5NUTloRPKCE5T9tCj+pkt6nOfTY6+7a0WBT33iPff5fPz/0C2qL97Ma4oMaCfIOPdlEOQzG
GH/8QITbSC8IJRu02w+IdQ4trhq0pywXsUARfUDa01FAV2SVkMtcz4jgEI3zkUIuly4H4uqXVAtu
qlrUCTnRqvHwZSiB+V3k0Jp8mk02155pNYITUXyDZochGdcf0/OzdD8aUyBQ8dVx67zlSpVK2Hfs
gQvTiUw5Gu0U6ZTBh88XPTpMJAqc4cE/obfMi9jCDodmFkM46dPV5cjrWSpFbVylCwd2vSqh69Op
Zs6tCZEnm+KMaRqygPnPJpQtfKzseHlhUxjbsfk+EL2b17gr8KJdXNpx4nGsa60rT/nz11rALkxa
eQwsRfqqoUXjfLlupPIaC0KGpWNTZPCZuVvgNEoKj4k7x8K2ftx+1pG1YtqO4iNEjOqPzBMZJYVs
WSKpoYz7jzA4BU+0V4hFekU5SIEi2Wb43hYCA/9N54gvQmW5lupDuVxChYqJpzvgySV4CofVcF7p
PwgKTIsw9cCUMeliiFLd1jf/CxCimKxqZadqnedXp+giZ0k6gutP1mS3W4R8ummWhvJJQsVDBkTS
EkAAoBrxPci/ZiT6P4u2OuaYKk36HAz9cOYglO/e8jMJMkpf1OOt/7zdOUKNz+2PdCfNCqcNbqE+
APNqbZ0LNpaWjsF3WbRjGpDTRpjzU50SL5sWc1zoeuwWXSN2FbzuftsRDz5plh/7DFtGEY6bcArP
E5NyMfy5pIpDArMLZNHZ3tDXq0eSj86lPog747MKDAxIyKiXUAM+RnmT/JksH0XW0jPLe/0MGsT8
DusnqUMgZFXEGPakW1kuBn2FZpzKdOEJ1Mhz6pe7q3yULoZp9iGZcLxijYRsMgmIEoaWZcrlmdwb
+aUklz/XxGNmWGn2CL1VkNqHxPPholjaaRZ2Jdz9UJjzrnYABgWOHqJcl0flSQTbrXJRZg2nQlvh
FevYDE/8A1XdnrUPfO0oIdcNc6zml1XR9lNNj3GI1qaIuyqMz75kDDmm0omeixY5UXKCOgRbTKCB
IMxq/OerGEiGLHoZAQOKlgnfWXSFqo8IR5LsLTbE1/3hcd5zGZlklWCgElMHad3jUl5AIbdFJjrb
nqWmNRDgnJ2+TNC6+AUG1n06ZGQN/X2G8Y6BJxb8FM8vII80rmqaaylHO+Xv5d3WneLkFGuvTdSr
wBOSiA+FcjseHZTiiLhc4nQgCdwM2VqTkFDsGIZZpArNnl4bA0cBruLJna8SXBbusBCdxhQ097XM
7jZ5MMGf5Ez2HTohHPar7QjAuzARmT3P0ciIjwhGuG2d9aJXf88oGQYwxHS+3p2AD3Y2B15V9qHl
7NycN5ccXIdqd5DQejH4VvinVcBB+nclrS9dS6lxcDfOqcUkfd+A6UdVD1+cm1I/8Ug8/nCwHepr
dEWESS/6+smyeEUEJ+PTwcra01OOFg7j6FjdQqEbUB9l8dLI5fcz9PYlM7jI7jf1G8Z2fc7XbFdT
AkQuy00GqMTOJeLSmhzvSR45h5eYmzOSMWTifjMrjkF2plH6wG8CSV6vj1vhcEz8sL5PjMaWpoUm
Hw2y65nDGp+1FCBByZAigvRrnETweZGxqbj8v7IH/7oFK4ep7MTLe8hpTIzZHElPQqM+HXnLbAWU
0Jh/VGa4fv/E3mYE1Phg7PezX0ZopBchqbbkNgLlm+hTvk/+xRZdP8SX3p9oquRIw1qHdbYslujt
Ti646Rj9MvHsAmNZSAGFKOmJM9IB+YDo2H2EncJ+jtySy7NUGEJua68VPMFhTrJI63TJKNlrDoRX
2DCCqg04yp8MkPbNhX/a2ercAIREf0Y1bTM+mI58CJbkn3wnrA2g5sySC/KGliw6/XJYi6DvhgLy
L3y7lbMMUB6piQUUBJ5usg+54lLtwIx71M+7PcW6yEG2AuxwSnOVGq4q0oXrIfVUOK0JBENMUjqr
Z2+8ILc2/F5t4c72gh1GCXxzrTBPOQEel6FFnKp5vlwYw6KIt8ZtMVWR4Ieyc+ooo4M/NO7S6KCD
VF1k+DDTL6L2CTPYgVMuTQULMD7jwE07r/r/cdHWSDEu9s5dVHhZtJpoWWrsWxWwOOji2MIvhBV/
o0rT5S44/VhBvSVScaSXoXn+T7WYyz70d5vI76jDimUgFDgfKqRzfxkVx5v22EOE0GZjy7X9aK0v
nhEZtYFPFzBphi7cn+e6OU+uAVlekB7hRtbDRLUU6aG0xhCsgowSQPouyOC2P8BrTFg1jSPiasyt
32dLi1s/c4Jc1aZsejqG3/E5otygufDWOnv5/1Ko5M8Gab1/HbVtGgpDQirLLG4SIkkfc4+bRstA
cf7iBqRZdW5NL8MoBoIW16E6IbHcyYzMqC6mRRUZoRs8P5GLwyxHWxU5z2vzlN+xbHBR4MfKWCxc
TL+Nwf/irCAF+4VYKAPvZyQ7fed2XO78GsujJrYmAGnpRos2lVBrS2ZuyfR210AKN1Hrfqxad6i+
2yJn2R6kZ1i3769VogKFVkMBffSgEhJ137FD6k3h1SWTLwVAfVzaqwVul5SS+KaT5jsqw0s5MI7y
ws66zN9cWaDEeH0sqmHidV9spW8jafjqXqWJED+vzunQBOprfzvaMiqCM00Qq+hsGmpS16iY3Bee
28IjdqyYepiwusHfb1iNvc/7aGLrpCkI+yIAks0jRWWVibJygq8AWdopnkQp2DV2N2MhbWBcN29Y
NOBJimJ7riFrl2igIg3xWmX5TILX1WD88HfQGxf5oy9G5UFbWWrzUuvFYC2wSkooc+Kf4IiuxGRl
oMi6aaUenAJ6p3htM0nsONOyZ6RbggXPfaP/ZFd9E9H8kGR2uIa/E+d8TmR7fi0PS22DgbMvJCgX
tcixXYs6dDDWw5m6xO5Lj0ORGscmDKChiX5bOV/jEVfc0eiyByb5egZDQBYTQN+jV7bCyrHs6Goe
m/QldXt0ggcBLUyzatomr0yK4OPldt3cpbthTBxgyTRCGyyODFFEhbiXmAhjNfQKoDNoZZXMLLi8
30mhehOhGdkHRX/NKw3HnbEEUxBigpBjG8kMJRUb60oZTxsT+4RqkMVwluOZLbUFz02FEKA8qOEw
iqDEoBxW1fbvcsKZL/1upW1DFRnx1Rc/R4ASpSz9JrkWJWikyzJMdQGO43EP0z3ozZE0BwvQYSJb
ZFOboK9aDa7nZS6ScN6drDJ4vR9wwfIV/E3XA0aPkPOuVSAg2KMNzE/n/cwc0VHpXV8EzW88Wr6F
b/utAInOCFNZIPmcS8q1PN9ng3QIUSg/WYY3cNFwI13ZEWGUU67AhpnPZqcbzWQTgS1LCZ9pcKCg
Urc5ysy1qVcWzT1HJ/t8rGlT6fb7AtimdhMgmKtITCMmkBpCLL49isnytExZj+e28lcvv6FSL1Yl
ImpfY6Wra5bVVpJUbnymhfSIwEwE+0KtuMzN9JLvCf46smXBz9oiUD169spZqmu3WAaDcdJxn598
W1haJZpVvSxbBocYTlqrNL41XOMWBEkvBIx50A1BGJokBG8n2xucNLmH4rUeA27Vwc4T6IzJrgN4
+cnsddVsxZZKHh/sHsEmY09IzkAwClEWpgcp0uunsBTMTzh2F4n1ibofuVx+fEYMV4mAIG8hjP0o
1fEWCyKYER5VhIdgJbEy24bf+uXi1dlXpYrPKona62WTTlTHaZ9Yim9gv5H8j9EndhYofLCl1kJY
mRzHjImDSDhZIHDmSWWOO4LIaC7xTRqWFYfoFaufettiSFtLtK59VTYFW67mV0iInpRor9Ep1Uql
IoiKoAvy5eMNez3XMd0lG6qADgHLCZMafOlCWLnvJSIE0uVtsTVxBsy9fRB25UVZcmq60rSooW+J
USfV+GdkYpihzwoJAjdMx9SkEs7EOUssToUK1hqwI8Qfax6ikn0f8xbyDvnasL+myevtud2J7QxO
CcK4t+I6fmBs/f+fdvWm/tjuc/rLT30wZLU42pZGyogsKzRYQjWx3bsb+IgDGO+NtIQwH7MQBySt
vbBTzo+1itk++Zda5JwM/Hl0RNT75azWc48Ol5oYpEOkEMqeGFvWqBn9543j2kKQAFBtRUj510tL
apqtFZ31TNB9uR3y7H97gHRzGokt/U4902a3/n6xXnN6SqpmH7+TyHT/ezVLnVRLOtpzROoV+rVZ
WGwqbkXp1mXjI4w8oW+liOsGDW4vhZytArQyvEBg/KYzRVLoEFQRpQ5aWYwBwWeqdrnuLED96CwV
gGN5caRDl3I1K3LnSIvaXagQSrxso7KzYzybEVEyvEwoOFFXh/jBK3AvvoUjcPwU7uHkL3czsZws
H44TmjAk9jxxHrnEzFSTHL3QqEt4G3ZToNO0IlPziv6SuoVTB9s7Auhgr/tr1BWPZVGb7FP0TIrp
djPvNmppvrULi/Vd+s4hhisXJsHxheX9xYA9F1+5Gd5lPGwhKklUylHUdhv70IL/ZfLey2nC8wsl
EY2iSgJ1MRb5LZhGql2bsKXeiUPGyRmN5LS3yTMpj7OBgiJHLcqL6YyklAGsutWKrAEVT9yXlhYE
uoHjYzIdpL0QCnedVD8kOViXTMVK5i5pX0lHha4Aq63TD0Hw3tOcYMMVzoMPbRXh7sv12+6CiVY3
9lYghvKweBCKQdEfIvyHoEhEVqqG40w7Qmbhig0kj6c9SSDwqKNRxEQKuHXMLZsmjYqAqjhLFgf4
IQY+PbebqCjv3ngzmAztcbvuRq4vJmX89xDA1NaWTiPfJKVADMrFtbpTI9djBA3eWkdNHgczKtLo
RqjuxM3yLM5RSZK6bKQxbK9UP8A+g8KlnHmSQtbp8KJDGhNQpsecBaNhFAsYoCG/dBdJDfIVeUtp
kM4fXwEbtACustCKUoBx6CNxAcDoZm8DNfr192FyXkgpoxFJWK4aJFtHUbDiIT6sDj9U66Hm5suF
L3y6tc3jlCiUoJcWFvW/lSbIDd7M86htcEMCjvSqBdykjjMPWbLNXMYHJk1YySwWPg4JZ8leSKwb
83dMnUR3htFMJFfOeuiLXfYWhpb99TyexgrasVbT8mTj9g5IpHRVFeBk8yBZsu1ARI7qpS73wrEd
RfHmj8HkZKhRTUNOdwJrAzwgUTtAU/P4ZlZDMzrLZEGQyedFZNYewpkR+WTQp/GDowK2rzbqMPm0
YT0yFjtdqn2z3fNH7rLveqH4jLZgn0eqsyZ/J3kNhY3kVI+wVKW4S15vrWF7m5VJ/SYbFK5rttK9
0yqRI+bPtH7bUt9qZMhp2wVFDMEq0ryYbzHNVeTVuz7aZ8LxEzLVmXJj5/AVNo02tSR934TyG/pt
YTNGn/lTRB5a3/L+wJQWBRW6h4A5VSH5Z/OCHC5VB2fvg/m0TEKRtlafQcsLgHcZbkBUY6KRbLGU
OoScBFeZFO5hlghuegG4yZx75rfEyAZJ11IDZhccQtII8uvGNH4joyEfOLOYLkY4Icqad5w5Sru+
FlwNynZWqPGviXT7tlLgP7kJ5iXHuoL65p1oP+PCFmevTLK3SN8QCuXL+fAAl0b2whcyknVJ226m
JuTd7w4EL/M43HjEh6YFuBuJTYje4lq10yyQydNCxFZk8ftxt9KRMwYSiZVnRpBilH/Ckbn6GtuH
2vUe8hixUqriEt5jpEnNRUrGAfv9gZDMjwZ/OTmMeixfsBM0ffhCYrCHZXlg6v5xyba6WssaAEGX
bE1PPjcb+SsSSSKlar5br8ggCiPan0vjWVb3A/Vt0847+QLNBrumVOE+LzGF1WvJQZIeBNHl1NHQ
d7w2S0h5ZfBnGinqzSO8iaTAdhsMYyESMrxCuMwHYKEyGFuO6baVW4xSpnafccsbTvd1UBHDWpgb
UZd5SGHA79nh6jz4tVfiVRSaj8zrlcthHDxMU8dyQhjMFIwopcX8cy4LOuVl3aaYhzpKUV97Xu/w
IWc7S05ovsUye2nUvH4Wxz4aZwPF5ak8j24XFlQPhPGg7vXVrhKPbx9BZMkOLcQg/UbR27HJwSwf
WReGDWZPhk5bEqoJD2+xkzKdHB4aYJcVBptKYt6tJ5uSj2lK4aSTBvoHIW8JGsokFz9oleJIx4LR
WPBvixPAxLMFdI4qhd38lCRPaT9yJad34OFHPxtiwgQBFQIg9Vv93jktJGFLhODi2UOti8v9Vl6X
vHkVWE00SLJFkWgpCDuHAkvcWiDkAwvpqtEgbateeE8KzeEARDKaJ/s0ynwKPvKg70y73zRQPByc
FK0mmaEelkfs5HtZCGga4CVvNgeBINnvmCLr9ufEC7gAF4fVspOqDrYc7f+EiGImxVwL4pROqKA1
zGN1wTaifR46B3AqXEr1WqGHamcMfrkx+tvq4AcXcqNs4DLDTi5LqIGiEq5b6ZXwG4uvgioKA1mU
VWuhvAu5Qvg5RIkWw8+wrMMHCGoA0fk0OZIa2AnDjgRHLVTv9CwKt/UOEFWLgtBUAaiPw7ajMJ8C
T2Us0aOs22bKDmH1dx/ynlbqbvtyBVFQUPQtNw5dgnLYa+lfH+k9GwH0xfJbP+NUZRYuPBWXQHN+
VnpT96uCggdxTQjJW9zcEjvLZTaJbhRufkzRq7B7SYjZ5tZDpfaXLRhArfZf/dy08YnZLXJa5HSG
A0ZXr1I3VZr420T9AZayWKg84a3tjkgZ+ALrmaC43JYxAmrxqmh8MW/LnwVidte5cXhplJ2+Fx2/
jvkPmzx+OnnIRVvaTxZC8OkGmw/Ldec4ewwwFkyfNVlVcH7jxDIM49Q4CUTy7jvZ5w156PvUkPqx
XrjafbNQKD3zdo0d/lrkQ8WX5QkuNzhUycULZwQen6ZU5/tl0FlkS3hmCEMF0C4Ni22T1hBNbvtf
0xXDIhUTcFoPc+M6MwTuQ9tsgdugG8GT8Mtg0dOeq9Dgatksi4JPXWsoYiiVTlHYXhqgA3uSoRO2
nyRP6DGDD0fvK7UxeP+H1h9exC129TGaKlQYBJ98oIl/xK+EzzGysogaAsTlOJ6rvnZ24smYSoRQ
UaM47V/wH6UdxxREaJ/m5Ph0wf9GSOypliGMY+M6Gnr5YO0mUDwIx5DmhEGDU7edz6V1MlwrZPwE
BjIjol01Wa7cR1kGMSeifUsHGVNcEa1FqheTHe0wUpIf8rLPDfTw66YgSYxUMAZFm2crj2M4Tx6u
clTwSPbJ9PHosVX8egssXAa1wnUJP6QMQ0GheSu4+tHLv9DIuP4K5zspUiLKlbGgUCHU+9uiZ1Hm
lizJeRuruT5O0T8/s73N6Kilt6kiFqpGJRhO9TqK8d6TSGhn3bHdAkLGl5rIz4ZNee/r/ceQzeE6
1v+OptedlyB+vBO4hbUxqf4cpowk4OfrdApaOsbyVPQqnwds1axzpC+Hxul0eHirF7QNwSgOhygu
611VcKA3vCk9QcVusoY7cdI3OsQG4T9lJ5dHIAcj4bqTbid83AnP+K3X0NiYvjbq6+/peqSo849H
0KhVDiPlMBWRK4Gi3E1VqXiCWkUwVE7aeCa0B5Gb4Jpt5chQAYg3LjWvpFxXEObi+ZFuPf+1RT5c
uNP7POtQ+W3MTEInN9CfMi8gSLN2K4bkaVBb/bQQ
`protect end_protected
