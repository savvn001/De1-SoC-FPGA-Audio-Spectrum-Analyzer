��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���� n;�7�Ov��@a"��3S�(����=�[�\l�|�$W��5'f�vWtX���>#ߏ�|ǔ��k�q|m��1}Ps��S�{ܢ^XMK!�_�����ľ�У��J\{9К�h��]/-��]�37{W'�1yΤ���נּ=�m.'c�Z��a6�+'�WX����qg�Ȑ8��Paȏ�8;��Uk��x/ȶd��gNc�M�]bE����p�B���rďe�Q
M��r=@�����C�3�U���mnd>��+VD|I\�)������ʺ�P��?�"�"}��6�,�m�ǏN����X�d���-\�����1�PP��f� Bi����t�#�b��@J��Z�m^�"D��G�R���$m��J��y�ho�/Jt�B�<j����`W(��{�C�vV�ͳ�2axA@��lb�����6��Ҭ7!ٹr�$�f��w�t�o��U���Y�N��u8�^Q���|2��P�K��g��e��_Y%�ߧ{�زX^�A(#�3vc6�(�@zsd����ݫ�4v��B�i��T����I��9��mdR��c{��T�/��P���]��:��A�s�=,�4�&#-;��a0���óT���;�Wt�|���0f�����x�o�G�yRCr�#����[j�󪠗Ҳ˫��3�TV"�N�<�P�?��5֮DU�ëtd7���4�(݂�R5���G�����[3I.�'P�Ӽ��έ/���A�}̢o��Ưjt�m�	�9��		�� �`�ԇ��L��_� ����99�7̏,J�̚~���LB5�Y�y,u@�@�13�R:o��\��]�^��˷�@��x�5�!�֗���_6S��K��fE�Z��+�aZ�	#�aP�8@iuP�S��F�T\��)}�vF�X �2����K�c���T�w�b�0���L��u�C���0��$��ǣf���"U��pc������X���ȡ�K���,в�8}�a�EMo�xzt:%���\Z����
�p��P�����i��D�=$�9g(\��ԩ���,��'��I����5}�s�S��D�PH���R��]5�-g�*���F���r.5Utvcz��q,꫓���3[��͕
x%x��0��[�����l��_Ub�脄%dT��N�v�i�<Eޢ;�BV��%/Qx7��fy�z�St�Y7���z��o��m��rXɊ�AW�;Y �a{V�,���8g���+�OC�%���ODo�@�B �Ϯ%��L{�ßI�'X��l�Wa֟��8D@������>��S���V8��"��(]0�پl��VV��Y�m�����Т�H�|m�J!��p7'�=��IP�]i���k}{�k0�,�<�1���!�Q�=7���)vf����,�>PN��V�	�+Nh|4�!�fMȘ�S����6-$�᎟��\�/�����X�����w9���.�avzF>6�2�ۤq�2�Ks���2O��Hb�
��x�Z�K��m��ir�Z�[V���Һg����!	��@K�W0�f�c&��i�b�z��!sѻ����C���6mv�Gp��|@R�(r�\:��Q����˹0�٘+����T�*����o���փS�M�क���8�\Z���)�o��ʕ}F I�&�j����b0;�So���,9�$�EǏ`[`��D��M
����W���ؾQ
~�ZHR)�G$
����+V��bE�A'�I^^�Y\�)�����~�Ur�u9�~��B���Q�P�¦�l�7_ic��o{2|�H�	���P\��[����4v3P�ל�8N�b{���N�����=L7B���P2�����9.E<���;��ȞZvЎ,l�ա&�).�-���@NOxA�j�8v#�9�$%���}�����a�0a��	 R�ߏ�Xj���@�&���>4T����?�I[��&߶cf��]	��M�I~#DH���\�hܲ���[���U�a,&���p�K4ɞ�FH��Ӿ�
��w��a�$ϙ ��O�l�S�����L�=�܇�]� �S���0��[�ĝL��� JU��ofH�&��[�^6���|�!Z�r>��D� 7/S�<�=s��V���)�J^�ݘy�%�w�o�꽨��yӿW�k�V�g��2����o�{�aϙ'��|H�?p�~>���wV��c �-����hPL]t���y�!<p�/a�"a}�L���zS~����
։ˉP�Z�v�l��G�m��|��(:HF��*�g`�,t=���8��
zQ�o�g���N��� �W���C^�@[�[��#������زEM���庶\������Q1�m��v��G�@灳&���H�\��������$���Q�������Z���	���չC��SUɿ7#v���(A����(ͧ4ܮW%w�d�A6��o�C�*��R��!NS��YV����o4�X�Xa[Khv+BjnS�t�7�^��J|dJ�&[P��X|�S��?̬9lV*+Io�����TӍxi�E9L5���DX�V�u���Ol���T/�����V��MP�(f:
����M0u����}�`1�%+����G���a�z��?�?����U�W��!xqp)V�������1mҊgn{hg=�_����;�B�����?�t���(X�]D�!�׹)<hV"��~#��r�S�`!ќ�I(iu4'�0Ce<[g��(RE7�_o ����X&0�ז�)^bR�I��w{Չ���q���Mʒ�܎Q�j�I�ۆ��#!¢"-�_�B�66�sM���$����ER��2�X"�# _M`��;��h�a�$���N�ϲ/)���j�����Z�'d��'=��l��v��ߓ�G�b!��C{�,e��k�z�h�X��-hp���j��W� ��V�(:)'���S$`�o���,(=N�r���<h�pq��N�����*���x1鳟��~P�)j�� ��_���������)�0dbphQ��*sL�Jpc�a�Y6���Ӵ�6�ܰt�{�\�� ]o��P˧��s��nI荜͚���9f�c-���?D���D����eǶp��)f�:kX��+o�@j��+֤��uA��풹ȷ�)�i����;�#z��;���d*V|A���i�,���ҕ��{���*�悟����Ƭ�#�,�2�"��5[�M�Ҷ[=w)�T7w��_�G�'�\�}W��Vw���0~�k�1���1+��ݽ��`�Nq�4�;��e�� X�L;EU,���a+�ڱ��\b�˝)�1�s�k{���{�7�Ɩ�읗|����*s����T�	g0�v���\6]&��RE��qvEjf���:A�f�����E>�q]Q�]��`��j^���ev�r���e=.�i�P+�k�V�a'LVE�a�l76u�,�yt��a�ݬ5�rp�W%-8Ɯ�i�{�r��,�j��3h��}f�e���y�s���r�E
�,_T|��1'�-���?A&�ZKB�Gy��7�8-��k�}��!j�����a�P��+؉5�Y]ǹ���37� z�CJO/s�
;���/��ށ��jP����A��)mG���АT3q��C�U�����ʎ2��?4�{-s8��o�$�#��å0|��ff�tխ_��*i�%*���K�P�t~�;�8��)NǮ L�jȚ�&��w�yP��k� ����X�Kf��e�	�K�5IY�}��śb��~���I��kg=��ӢZI�B8�.A�/���)�}\�ϱR��|ϠU��q��1W��ă[d�Q�{����8�n�5�g>(���*h[�	�3�G�� �s��������	�{o��.J�q���[�k���vY�Ϧ�e(�͉5���M�pxy?c�ֱ9�h��ק���>7�S��Y��w;��;�Ǯ�C��]�aoj�G��K�B��{zu�uz����:�-d}�H�#�5�[h���zҴiQ��}t���2����M�����c�Q&�?��K_x�$,7iY|�Q��1�]v�/"YR�i\?=X�n�� G}��o�2�y���E&Bv�J��;:�_�ZΘ;V�]�`S���>IU�{��i!�E�k�y�y�