-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Adpsb3HFHD4YYIzYHCJrRdYfU+jVWSlt5ViZ8haL96+zwJ1ZipF7Y/iecj3Fr0Aum5NqV+uCbfdA
PHDqX6MqPCzNnu9kiaGZGTj2NyibA6iSok/G32U9YL0QssLpsNT+P/EMEjI1KeRxbAIydocklKGp
eEIkl5DIgJy7qzb9NLQ+WveU7eGUC0IhPMb8anrOapmtuvebUg6R9WHGwXzRQuMvZIifzNRvsWNS
pxpvN0+5OY5qpEc4cW8F7q4vNVyiOyFmMxvjJgmid0CDH1zgpXTaw9HMufzkYodvfvZ/2saTHITR
EUpyZTkpd5V6tePUqlCXiKVdnnc5L3YtmAD+oQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
cS9+pCiBJGwHtltP7Wt5As89CPK6ALkf3GIzuaahFS3WMKALtZAzWM6RS+HqS9+t0G6JAQGOShZV
O+gpKnACae4LmaQErjupbkgOWmoCXe6lfKrYbx0dUMkjt5aV9HbCy8Af24MzujTuXUXJRxzOLETL
4eJdr0tJkD9a1DcFDrtI3vwMIFckmKDik4wv6tR7WRCeSI8tS67vXhEKID95ISFOg6KzNM3waoQZ
pucpAWZrzqTVQvyRmVRtolp4np02HD5kqKr8DA+i2KDaVAOhkVYyCSk/DhbSUPe6jwt8wnBfwz75
NjYzs56S1tJVPslA5Qg0yKj8t+od3faFKi3SSyIF8PYNANABycEn1Ani95o5dAnhc7KDOOBRTQG0
8wBhFDf9MIfyr2oZ14W1ESNKf2SxK7nKt63xPDuh6X+zNCiNF6XyaFK0cKXYXMtVb+YnqfqpAcyA
r4VMLEKuovsJIPpubTtcpxTsfETQBeDw3buvSPIeCma6tqiRasYX3SUCKvDEbz+RA60ig1eBattT
FiCgQpE+vQ+oxdKzl0mn3JImRBcA3iaJxBcRf1euQeDCNh654gz3NXb68TBAr0c1cpxtOjHLwkY4
8djrwvn8rsSAepcXkApCb2UWqvCUSVXE+aSZb+X+4NmkoogZKiGppKq9OOI7RvfhVERE26wXA/T8
20KfMVnIaFF/pn0jtCK+uxTcOjhgQFc33VlhXqW/J2PGjK7bZhbYi2PSEIBfYEWLvxyWBLUsv8U/
0nbyx1mqK0fVVFPsuENOuK9dmnW9ZcnDCwCHtl78a+kGhJKC4EwbYgkWy9u25CYXLkThbV9qQd1n
L6diWI3X8DujW1mi18ZZTIX2rEtpJfWEsroEWph7vIyuiqk5yHuMn0rcKWfn1xAsXHGBGQsjgMIF
3TFQd7luwfc7yin9fGNpo4pTdx2FyYSJ1zrnJmFbfGIqT6qnOBI6DNsL3g13CaYKb85Bqm0fKE+t
XpsWCEaPSNTQ7DUORaqQ5v2x2T4T6YTfqOpIUnAJYcUP5x9jimSXSym/yCl9zC5TAa09N9j2J8cU
GyUnCHNPH6iOi6/NHr9s+KVBeT/5E5tqqN2GAlB95nIg8Pprzx/GTnDmhmm6CXaMOXLg14cdyfSS
Ph+zJ1Vh9+arX2qka74jGOLU9La1sqKqUY+11BrAx2VgPPGsiDdVEPKS7PF8ENkxxIc2D//pb8dO
b7CZse0Lz52yIL8o/NpHdvSI00W5ENkfKoGsmrgfbqFButANgJXoHirLEks9/0riH9Yk0pxi3fNH
0SbhWqZDcb+vFgRjs0V7fG5XBed+4NOtH0V/87lUQlXT3jm6mMgl1xumE6HXZ/esneK+YygbUh5O
vYnpYbAeoAZFSNqf3/4tAsU+D22TPTIEHCIFWstNUm3UfIQiNN3SxR/4IcfoPNcPd5n/kYtn/d5q
PIsjSBwPncOuJehktFo+bdzOFyWeenhT9ymvYJmqsZuzKTUprKgWxRJ+/wbwmR8PAb4wb5yeqiwR
h6QvEu73CAgO4umhP5GOwcMVJozmUDKLq6/VIFv3uFQ1oe7UDWyGCX/jgEVrG1ob4SZ2qhXWSq7/
LKEVGKYjuQDqvUj4K01nUzUQY+oaISsubq6RfcFv7P0cHL4mwVJ3NLbenW73w1d3TiJtmRwheyeF
QUdmoAEBRqcOv9xO9kWNhUjPiCcz9bJa9WOD86NhBVRl+Yl/6LkQnlmeHMkMZNbISOu7jRS/4Ilm
TuY3bL4cvc1OQ4+D0+H8ZdnpvENasjWffL0TWCjpjvHZ+78ZqEaQGKKfwgZWWW3iKEaCycyexy/3
Wa81cw9Nb/2TBaoXKBaOrG1jRvVs3098qsvUkxTxETOq8ORTQ+/5NjU1CWA8qQnxCRzCGLokkHZ2
T2561745N0dz1D+I9q/iFTwX9sc++SsIwla2x/WUFUg02WnMdiWs2D/ky9euOicPL6lE4CetdybN
+nNbVK57GiY0hwhW8XgISr9JfUoryGXB/rw5SszA4kJ4kJjnXv1hqo98yn/uGZ7YXerHV5uQG9AF
t3zyF+IhoLdv8/gibFa8uKpC8SXrMs7EXU5XI4zgIuPcmscHi+ZoFomWfCvwO1OXpH0p80mPA8ST
YpyBZNCWu7x+uU78jaZs7Op6+XZ7hzTxdxsbwz5RqdXmeNRVMqXsrlNd7gEviHx6uACNcuVvsoh4
RMKmgyaiVXSau3WYmHbf9/QMoP2DW6e69iSkPTTT9eQVwyhqU2sUHQPwevMjQmP/MdEL/3nK2sbz
7PY0Fe/PLpR7mNZriM5sUT1WT+aSdRhrJyJr3cnh82mH0YsI0KcGH/FIQwj35WTlp3aa+/o8WCCv
0O9KyUINm5QP/PjANgSsLTBo0P3+F0JTCq5BCUuUmg5+XyWOYLEqsQ18KMPdfZfain4JO4IScOSd
7gzQ2mVggikfFGzabXWLAVcLdsPdAldDcX78qYMlw1Zn2W+tingeX0Jhi5Ax1pV2tR/+XwTEbDFc
apemi8+TZ+/7X9yjCLPRF2Fi+nxOAm6I0B3ToRmFGWLUUTufvFir+X7NgfxqDUKzkRV4Sj7sszx1
U/5kEiK6gkqJuDHn42WJvQAJ5RU+vM0ccrC508xh04O1CBc3XDy5ayeGjgXWkQpxExkzJ5kLhgvf
8NeZJZzwPpVQxnTHU0szg3RVis/PXTo2W3Evhjrrlw+o487fTreNro5lCpDmQCi3YtpMUrDmbHqd
qSSWfw4TVGoYUAif3dE6LppvuBJLi4S81U0AqAXLAz/TuOafQMWurXYnPyJqC7Fu+sEJKndxMCJz
y4rI8SJ/7GyXlVwWILJJiWtl1ZK3R/PwkdWJBEM/pbRXTKSzAhwC1SJE1h1nFuLv0GvgZz6nzZs7
MmT8BQ/2wZiStsA+axJcwIpCD+xWpXoPduzybP868sOPkMfjpISZfbC+Sg1x0zKh7gCwz1DT8lSe
DyiUTdpqTpiKGGmIUrpfLMQdN0ec0q4BOFq8DoYj/sj6tDRFeT6Rq+7B4k/ZnJSpzlVnEDCkQjuv
X55lkuPRBhyevII5YWIRKihdHgynNtacsiX5dFGC6iPE4RzubHKF0yVsHdeXXA3Kjuk19Bn0z+Nz
aYstnCT8Mb5DX7PhsVtrju4nZR37yY1yuu8oE4Nh7MWSoAGqsczBF+375H7HxUesIu5z3/ZGiWSm
7n0vUeYTcMyNWN1VQkhTRFjUS8sxaMveKlF8y7MTJ95UDYuTDadEuAg6coLuocT3uWYKTZOdQBsP
D8t6aTfb37JSyhAxSBAp8MRTwFp7Pn27el0M4zXFCWHX6d22lToqM/0t/6tbH7MXwMobEjdjEbhq
QY2FAeZdoXVpDUEbpXFilNm5cabylEbmNqGHXwb2J4yrZHhojv+ZB4KOZFuTodxKNI8wTGRQJq3T
wXJjz+IRkrSRRj1oHmDoGpGoFJUDODNOyi319TczPtzUn81hWxNlPcSIeGjoOkyYvc5u8L4B4lwh
V+AlSiNYCz7oEIUSLINjNxoc9i9vkRi5rw8qgzToSxw7lsHhbeqQMdeT1bSsmcDEkkeY4OYbcbtG
ZOCh2wmH/H28hG/uisoWrLuABqPTV/8EH4vFChj6MgY0mqjinxowhtCUWqwTrX9hJFf2UthoCMSB
wnh8Ii68bnHMv17itsPrLQY6vki0c+PQmEinuI46hOOOt2qwPExIv778LSRJ7zAOAzvWl4x3LiX1
05ok+hyWUj/ZRZ4hiRamW31fs45nv+gD3DsOpAtrzfjR5cw/kIpzky7kgYIK0N0K/oq9XT7VHDi1
Xf+oACmEREW62CDmTK6KOb0Z0g5hTjaBghdM4W1C6ZRZks8KgaCqd8xbRTRBfheVUy5zivW+NtHl
xuF8XKbYCZPfm+N7hR3TjnRRUmIRLlcqKgEZLDKOANcJfKt3HoC67B8T8Z2DSvTaKUP0epbmQrJR
zx25MLE+4lWKxx4cOMrNv5CyBfoH+XJBUJbdjEbcF2JzJNw+YHGCkomsfSRrQqdlIUankYlmR3px
HkKJZpy1UYbGBMuY+RqbnBV3i3QeK5L6eS9ohrvKClAbOmdhcZja3JOXwe7yqWhnCEQies1wtyPc
0lpaqnGy5+YCXXTmO1/FEuPRKMN1bQO0nWa3eQJW8zES3kSx8jHJxMVeRQinUcTA9CLBkVMtTpJ6
rccE7weaYSlgszUfsvAOsVmkm6WMC4HPyDKW0Lm3fenPw3UOe3l8ErU+YoMiMSvcO68WklOrzi/M
mWhjZlUs9qmwjYla7y2oWlXc1+UyrkoPLm46GR3ysn1DjFtV9Obw73SJlvgtF5ZGPvZmP1pDvsP2
Bu/csj7cr1W8PR7SeU5YqpxAGyYzJl9cQZ1Mu1Dvuu4OdvMdlNpZrvvykAwa+W0ZoqlMAtGfzW6Y
nd44KA8GtvFbNUPEGdLkPajZJkatw/9RnuGQpHj5COgdYiFiBp+YevZLWn2e+qR7xFs6fnLk5tPH
yRVopkHrMmjm4wLsikW0Z0eUSzYippBKnj/YzKbUR/FNfaRmlA6OiR9InV9nCLDv6lSA6CMLLUhB
nklYZbBHKasa2WVryyOZ14A0uT4U4aIa78J4fvIV7LHAlVewhCzKzXdB9/xfmkBNO/kvfzwrxOxa
+DQqx1ZtBTAlpq3fSnnVGawhKRynzdoqga0PujtcmaML9IDKvckySPe06JuRnwOe9JJmR0rd+0Mr
HnLmisKwKcNBYRQybXOqt/y1F0Oy+ZfCPltlwiZA1L8vHexlgP6rRWqNr/79F9aA9U1OvR4qdne5
Ch4XOY4UWHAtOrETEX7Ff9ASV+GLsNd6Vd7l+yIb3a7bmWL2/Fr+bpgowk5Luk4zNOFHWgmpDqEr
4XNgm4VJo3HzZ4y5nJ3HSrxCRyIViI0Idljb0HxWuSuw0kFyA16oMU9FxZFMHfBxiGwYcria5SFV
Ec5Tqg7q2WjPf7H4HOCWMBb899J/Auz/X29vlt6RhEV6In/IAt1LT4y4GZikbHE7isPykIEuI9Zh
Mw8x6dyUYWKOBj4rrgjH7YMb9LcqyNN8iSttlFawnbSItB6vkO7mBYhJmDiU3Iz4qkFHJc08i/vE
BcPo/BUX3KMeU2QypC3aJvRC7qJB3aCQqtZx4UCCzIJe7NPIReWyjXywGySrY+F/HX70y9Yqx0Lc
QmxleNDewH3NW6I6n5HLJMk+4LmFjHC4wr+6HFL5c0rPBedGqYNW6eUMuNuw7LXE+eFR6QbrkPBc
LTS0BVNGec7uamZ3r7JQq1z5zyZFQ8EmdB5rnvYW5xvS6dT/sLXmdM/laAhLYo7iUDJUyTc57q3N
7m8GzB9u7PUdmiuZiTkuy0TkFTVw82oWK1liCYTLfnC9m8w1VnWwh8lHiseQ0Oat2LV3nnoU7cUP
KkvRCI/c3Yfu4+BfOnIejzj4K/i/GpTO82VeIc3J/vAs86KkmY8pLyROA93TXJoSPJgVjtRNZUqf
w4akzGclheuzKVps9k0l8EePtLtq5ovacICb8c5gSajFDvdEPUcYjzSuOF6ZHhPhuuUufVo8E4JE
0u9Wm28B9V9957WVEKyFlfrkkq44CqJr0XiTilzV90l6+XK0Fcdv6+61WI4Z+SfVGCp+kUeaGunS
WVTNbfL6czJ+8tgTGeNcPaFNLCXykxHhzOTVisoQGO5h0CLLNh5LmE0p6HQDYyxx6DKkLYmxaSwZ
PvxWIqm+LTipCDDg5ZvQx1EOyhL8kTobSasB6AOiuEiRxd6rnCtAI5zGOlogdqIAT93C3W6tBHw2
d3/rtg1S8b6JgfAuDi9lgMqFfQaUgS/9PyEUiQH5TnQFlmhkXRW+R9b0aLk4eGNITssW4wdv9pOr
kmAUmg1xAlzIzi4KYrdaxPQvjN/9xA4xD1tj4X8/nO17TZ1T/yKlZuk0R+J1xwCnQPPDgdoSQS0Y
YHZLtx1moaooZuJPwLmN9BTRjD6ARDCe1DC0JnuqkZUhnMp7IbIfAHdGEqtVUe7BPp0ji84j7BC6
Hhhwmt05Hu2FtSjmqosaaRTOla8SCJu7GXy66S1EJ0pmL30Rh4TCj8YxYg88OU66SOGP81ptCbQy
p8ojYV/Ba0laSHHtCkRVfN2MKhG1wDUd8lzPmTN3bDeqmgmEGI79b75nyoZwWvpnKGVeCJ03EQUW
5v6/AngyNbePorNmw45wCS/SfrDDQRu5a2aASHmx12foPtHjodQT7lYJ+Vk/0jhJkBsS1ax2cDep
XbixnWF2Cp+4CBVG4R1DZKurqVthrDiVCxfPCjFC0bBLuseci4LhqeAMbxS7+rkHlvHtljgCpndt
s4BUi//pjTGsFeiftCj71oA2mfX0zMEACyhtqUOGQ8wdINRLzwFaufBZ8EJJP8w0mr717UJkXIKK
X+RYIEEmhdx3sl6+5+H0mK8O7YOueZ4NxGnFNIPjK6yioCkR29o1i5NbHi23H5lyCN7wfqkSNMDo
EAFaE11eSGp3sja7iaxV8GmfQBX8D8DMcrqvLKJNlzCOcA0MP1F5Mj6mbHYq3LQy1OqqCD3Cy0q7
zFkMohrhUvoy67Ob63wv15uoJpBrYp/d8WT22mZdarmxuM7lXJONM9BZid1C4oD7MDMqzflSI1e6
cTEzAdjv8mv2jqgwhqv2soIXvyGEEChhUzdcJBZ9jb4iaEh4x4W6ILnbjqYB0DOzz74bHLnl01hi
lJQpq0Ne9D06TYOVRTGZbQmkjGbmBWOctSRoWXClhSvqE7beUYX2ueSk0QaNX1urScEG9R6y7YKv
zqJcsvPPmJMZ0r/vsTPcwqQIqQ2kmIp7JboR+GgVJSh9CH+Q3wI5Xzjwtc/4c8Jd5cDV75uLRT02
as1as2mQoK+CbvwAjgp3ZBhtb53MxAg+qE6N2xPmLiGMKukddoa86omLQXHNlGBhTI5EkDD1wJkw
K4WGHehpfBdI1RP44bb9SazTIoeE7i4lDpFuounJYRj6t/E+riycqdg+VDLJPgv0R4akr2RtvUHI
QMxV+QDpHUJMDdbEFBSoQq9ZTnIz/zHjgDOh49nSwBDnY/9ITDtnePzKBRROq/Cr4B+LtU2qpJf2
NPXfNQSu5nub4avZb1rtgGaCjiC+Qd48EXBlsjiEjjXsU6qAo/CRjBlvNLwOOVI0EAYjGpGkqYk0
t1GMFdO9XuiqwTTSGVaALy2tTmx51rpGAzLouOR9YQeztBncaB7gOSRunt5xW0Vpci/AfeLljDKx
BhJ2Ljk4IWk2Ql2ftcFVfbXzq/QPfX7lZ9amv5xhyS62kYwLXN8pF4cDZmmT2PxfITIF3htvFcpg
YiZDhysd5ITAfR6mhZ3mya6hLGsjhKV557j+TFCEVBCmmyzXR8pkurX8cS9npWUbbHC482ib63Tj
zbty++jWmOCfSBXc9EKJgig3K9ZZlhyLLPF+xEYR1NcC6hHxGsByw6q0sWXNlF5kF9naSJ9X/bFW
rcjuqJCTPm2kMrQfwLjY/qc9U9Hnby1rUYfuonLWeiuwskTVBjn/vyICsU4hgV9baXrR+Ep8njiy
RkFdM3YYG1k/6Lzqaz55WIW+BLswTYl51/vMt1+gL9w/0gi2Q9AvWjW7jZ0ppuiOYA9koGJUohNS
tvJt3374q/0piW7C0Yx3GBo67f41nWD69YewJ5/EL97lZwqqtX/m3S6E4ENDWuvsly23CBKp89oC
YPLFGK46S3XZzTNVcdhf6tpobSm3NXDyGgCQN50YxnA4IF2U/xMn+MPLxlbLFCCxCN++EJc/YVH+
5PirsNQE9vWirNixOcyAAlRvSeRzekw4Pm+RCb48J8nkDz4B1jrG51ogLar7H2xBF4bXUx8gdcUU
db8g6WzAXQNrQYa9xe8PdqBRNcxpIrSteLedXSofyJ3HFaxCMO3L30x7WI87Ekbfd+mK/7v690m8
Re7QQUe5G/8xivuVvH6p/BZa5MHO5Jr6OyOhqp00nT1bR9c2wzbeWyYlVlBTnW96WHD0D5Qb/LCC
yg3Pcx6VRxzsYp57PRsH2V4hz5TDIZfTqgOT9IlYKG28gypt9lCFa/vmg0tyxNhjkUuED8NM/vVT
hXT7w5MxKy7q/KygqunR6957lIlEMWIXhUUdqxQt0wo5hRlZhRHFKgJ72QoRIzYcx/rf4+xmmzgF
LMdOzUWSUo1sA3VQEOPKKzb1bO39kpWiE5rQQ2lwTGQzZSpT2tC2Cldg96A1s1E5VXCGrxOzwxZQ
UVeWdwPhmVibLaq+WjI/dNfBbKQttWBGkxSSkQ5ZQLDVpno45y4s7qAdymtK866rCKDoMO8d+ndX
YBkfeXwO0uFqlyQw78yy3eG0a384yqj30EGfubhQZxjtwEW8ccbdId291JMwKtWUmwSk+1D33nmD
hwfnlqRajTmv+Y99Em4P+p5GyD3qLWluxnSYSBMlWKmoAze6f+IkFKT/Hcb9bwgtKaD6hP/YJJS+
PJZ1Tq9KhzcrWGToQ0AoUPkQYltropEV/oPWf9PLi0zpcUbs26GbYkiwb3CdSxEyyWmvMtuXuFas
GGlCA/RBB3FdGxtVeRkSPoxmges1kltoBu/emvqWpKkAld3PMA4E3jkYGZL1hhIJia7H8gTmP0BF
J8GzLMQ0DdzEsqfRYbU9OukbbD1a//zRCrEgP9cIILb0KDbTD4z9fWQSLiQTeFCuEUz528ehnQXo
BbdNmRHFLGqgsy9nEizysyxJG26skdP7AhFTQFfq2azzbkBecu9EPGSu3nUsNAoYMW1/qoB4GLHU
2qrPDzc7QHCNLrKwUMWz9CG7slbFUbA75CrPIEnqympbh+Ots6VBGP7wFzQyWFfdWGcIH0vUnV8o
i6hjZw9rIfszBoq2UssGSZjiJm3BC8uf1DFi07hAn+7vMedJHeGcanBQ/OS2U2n5V8MyYkDrcvQc
LhyOYAwUs0O7OoZt3LamNf7053jFgO30FXznGS0EiAaSBz+r86dRAgw1wyrxwYvaZLViqssUwbN0
dt32nDcY+C9TnTP0nidlryl7EWbxnTasWJqGi/P/tUgcr+5TxOpQJzVdmfDu44KB96pPL7+deh9K
1Wj/nsWhM8UQaMUpIQpec/PAXlCFpYUsaSuKwJU86Jf0CA92oGgVYTEtwXVfAJeOVieEyW9/c/pV
NBQoMBvK/tsA7N4RPQkEarnfOlUlhkdTxK/LIETPH3LJCc9lO70fbN0eg1MPu2FrRmuU8tgxjz7H
7CxPXye3oFrEYr2Ej8bsqZopF84tRLg1rQMyAQfxNSnQMXoAr9VrFxFziJgdVxSme4VH22EUNga5
tfNyeH75cRp1odXqXD7RR9iu6aleYtbr47xlAf0mtABYp4er0+Y7vtUg8nbEnVZRRrr5vSLbIWBz
5vvmyi+ehTxwo6luwcFctg+SHdhveYNnw97KcOprqjkmLZTwsczKnFRpwzJbykpl9rwWe9jTeG8+
DOU6ayp01gOHM4EgRx3zmIi3XUnrws04UIomLGj7IiU+JWezGmlF8qVXtEKv+qmYgDjUDnLGJUVV
ob2QGhqQ6BwEBCJ2aMHlA2RBsyT9cqqOYgONdlsM00SR1Vp3aqB96g5mOrT+BOh4XiHcTEJTobGI
CoH73Lh8mmXZO18dnDvZ48PPUpoLjfPSAW6784tQ6xYEQVWlacluXtGedEdA/sJDqnUTwBYZ4Fns
vjQhsZ6E9cODi17HLXGCB531BQlMT0l/5JjtVUiTsaPHqKraYEhiFYnVbCp808E2IULckQgfJ2pK
ZuFdrzAtnksxdnc0wza6lMVGeH9f+Kv4ymLzL128w9fe+jD3+q0RqYmYMsEufkKhrKhy+JVHo4PV
nW1/AHClqPiQ8AxKaUl+3X18s4TTgIaceT92+p25lTTuUj2SH4gEvlPH1DiQgqAxxlxWM8+NQ9Dn
kj2yWc6vsPMWOQbuXQycx3mfMc85CVMst20ui74rGaEACA+MjB9ngBoufVxYmveqby3DASS/lgn/
0mfjszUMcjP49Ezvvpt+5xGWf1TbLIt9ny8ZSBU3wkwIccpFM+KHDm+kpoq/NF6OeSgPyn3jBcaQ
98fyvU7ByRYGXd3YLCxrbpVqDqRa2pbJ5TLixVis49AiDjjZitboYqcbjRBPWUaaHp5kjSlMN7Os
xTQ2loR2nYpAB4Ih16eAI4uOFGARjaFiq4Xt0gt7Jgk0XrRDsWMiXRggo/0YE/O3V0gyIq/Gbyww
lRzhO3Ho2ruP64VZXTqkRRcuiktnjvTq3ac2PQLCjFDJTuvekuVYc2rssocbTwZuOy1Rp6opqDMW
ml1cxXyJBFHOzO4dSx6T8GqZpRsZlc4vwFEIjZi0r2IPnx/Fr/HxkUKAcxpzm5/mjpxU+QKNYBsL
10oNzFOWn2VNX5ZpUh4frDN21glYyN/A8kUNo0ai6UyEGb3e01mLvG274Nq0tIQVupm6K0V5cEp2
f+qGdXcR4Ydy+utUZOs5DA+VNrexRQ9xawJLGRju2bzICwl4Gyow2PkwZ4ZlpzroiNvfVgyOZSdZ
wjbs58h3lFEbp4rsek5zlhBw0ycM85CyY3cFkCs5rtZnZufDKrCRiEf1tmnuqVARErfnFE0rEhKI
gNAkjprNjsnmY7Pesj7+WWMbBtD9+ukNUROI8zThanh5tnjmn6B/Rp1Zzd2bShIefLyijrp7Crm5
OKhKwB4cyRmIdnU/DBxhy0LBsRxzC9So6VEBktnqs0UuvVyMkDThzY3OrN/ov/+rAck1XsfwSX09
717XJI2m+rYszN3nlwjafW5z/bYGbBWtwJWcCPkDyFhqptIn7JZfEA+Fp2uHE1xkCDnM6gCRT9Xm
pVr3CSwoUQmJ4f7wNfGQFc5x0fWIrexuNFj9SISMtd0c4e/rEgF3vE/9pMv90VaI0TCEgDpkxBr2
CGHGn9hmr9HEAyWCxAAjHu1Ws/ymeP68Dg3iDsu+Jy4qzOsppJC6yFDFr0rUdka9Xn8vVKawe7Zt
wPwwSLg561Ayo64mRvZ0GQjAtL+GXLG5yiYw7ZHlYFKXB/IZeixqtOxLErpOJ6MKGqsbKUBthvPu
okJMQNuwut6Lwqr+BoElk+iQg+hD83Qex2FE436xRx+YjMf+Om66XOfAeUUPZS/ZUbMsfQ+akAt4
RMgbcR53d/NCdWZ5k8UJt4CR2nCAKHroJgCR2NXKPMAAPq11LRA5LRCBBQvtfbjlMlFCMioibz3G
BWG3yMuRmJcFNTjtrps9TldCOrcuJS2pj0OdPKY19LZkCl/Mks3pi4rX7HZTvRkjYaEH2OCm/bys
olxodGet5/wGeMnd7lc0Hen0o+6M+RrZjSeXDJ/STwiJIpEIcUlzrjFGBkX/SEmDO4xq7bnOeGmt
sxfT4EBCX+DMhBAoIb8u//+t5rsPrqrtaYUaPrKlr/IzTBTADO0kBqyDGwMc0h6ZItMS383d0hSs
2mkAyWkQYGMu3JqwRSU8C3yIHVxTx/qefwgQkn15zJa/2SxMrXgnhgwy+r1AYNVuSrmCD3RqparC
OzcqC+xv+cB+DDu74t2Yke3lyRqpm0ao7QIq3G6uaCe2AauZuz9bRumwUtKWX7bHUXYe0P+Mam5g
FpkUUqJUO9R/pxZby5gsvcOPF3KDFySiIEVQ9Dr7U2QlW/GMA5VRHskrRChmSOdeXgdLvmeuNwAq
V35PqmAKg7ZruX8Cx8O8iGVR0DC5eV1XBEfd0zeO1GA9fIi4qNo+e8k0QSctn4jCUzEbAyOr+E7q
0yjkprR9Y54KbYnI97v2RzBoF/DMoBIyMQlai5sopT0pZkXpYePyPep/zWYWi5JWJJ4ZiQ5IOtGl
ZRA3l6LfD1Zi09/5YXj5j0UEC8Rt7dUspPJts9K9mCsaf0xhR7oBdjmXzDQX7Z43OsRLUduMOs5k
cdIfIqFQBVUUyQgNuZ42T3VAFuiBEuIZ1aF5/duVi/ULRO5g8w/cGyX67y0IX4QGhwC3wI3Z+z92
Myz9U3eFiYB9FY2ROWbWajg1jVppAKYf2ck/Kszd9Yw4WAs82XUFaEo3T2rXPVKylCO+rp9FkxOI
cii2/BubELk2VENDyQ1Miz+sSMi8dQ7YeY9sjNJpYDwte9rLW39HvYHTN0BPJ13WZ1jtkC6tDiUl
7rKG44hvQ65KeylHsu0mAVte91GIiiubE2s6nyur+snc+OVLV/QaawaOzfuVV//40gXw2zOQULaB
mZj8TB/ZLwOAMUZE4LxeYH4Rv8+kLB0aBj5g7gIVJ0alDo1FZt3Og71cpbbiuMVb86PQMSfwXgVu
3gMYDbpfvdCbptCu4cyblZU9++heQc/feTVX5YPwwYxZlOgaXXa1oIG7/PgT6US+1+uw5T9/1LyB
9LYr++Xprg4dutS1n+4ctHhPxHH5oxwuePWM06HTDgBOoyzTENo+4rmL2FM5O4+TAL9PMhYXnl4K
jHpf5iORuh9B5dvtGzXOACBiBbqhiPNi0JyJdWtom4dZvXmm6iguAhncZ+QJQz66yGAZs3+GUjpN
lBKQeQqd4HduonXrYp2Qx3th3/+gpar5r/jK5S1TDj7gLu8T64SugERDWZ+cvr93KZcQFcQhaoC1
nL6J/ydJbyar+Z1ogPcTVMyAqNnpTXdi5fxhD9SlZzd+u3krlDEDDCtyI6LITWWkI1NO25tLiV2I
TNXL3HXTSwkm+XG8ry3bXmZzVoBXEHz0dAG1aTH/p9qUBn0HO1Jdxx/9e3QDudIrjnQmEWkJwLS1
2nG574x9bs+D5rafjJ2eZeW8wGkKI1gaDWve4LKm1Req4JJD+H3kznjSjLsiXUMS23sXOxWxqzc9
UXY1YzfepGtYf/aaMGhUFgy6ARbtsstUryRsvJjMLPLWDDj3Mqz28ZwZ3ACfQwpIEbrnh2Eog0tL
xoKKJMTXQXQZEaT/75WwSSwfTKj6CI3UPqUzYPHceSKSUqaNDO0HCUfoS8mDlKNnjSniMyJnYk2D
lFu7HRjidDfwczSxOAAxMGDrvA+HbUEzMugOwzhjuV7T6kkqwhZ+2Oz4jXQftJppB8mF2RIQ4Om1
jNX7nTrBibw1KlrwOotoegUryeybmvZpnhn86hepqTrSs07bsapi3fw+zcLY6eAO96zRiq6Zk/wR
PIQa4s2/eGn7DcUSjO9GB/FbnIuS4rKXCvWmf2S91TiNt0Xpdl3cWrtvl5TcsRRIC7qSlBfpbOkR
7Jp7wqXzmIUm+U9rRtPyH6pnB53rKQzm6t3JyEWjh+hrGRM6yPfGjfCrBp42/sTC6BaGV1i5ppK5
j/CzK7HRurW2PKtFwRxStxFXWYVTTxsUMiFxjAuzZRptcQyXtrZaN+cZwPe2iSIc01nH0KcHaqoU
zVOs+bgjJfidF7CeNbCO7qVLK+zHFK2wVkUrOoZOCq6wf1EQXxAKn/qN6Jp8Bmt9PenSJ10N/7nC
IvSKFG1JUqAqS1+qJ4bbI9nv0qrIiZMq/P+faslcD9IKuErD/M3VdWkAmX04HUk7R3ZuPj3oksMd
BfAk8w2JW09vBFDLGEJPEkhQYIRfQ8naC0/317agaNivvdtuWCKresmH0cOCdveYQPzd+hGCZHYk
/r50CDt3zATfbtncWxLxfPaO8QlZqu+OxAl8NoKUfPMcubPvSHyreJytSNH+Qg3mseZqO8tmUv9I
TN97cwvOlv3c02e8wCmL0wtNmVimh/QYM6KfZmGvodwjzutYCb6u+4s8JnCN1HWnGKvGRA7411BD
BD5xBQwtL3kLzdeU0W2nbjjDFTbsgVz+cai90PtBE9vMezp2DkvIZVGWiqIcMxexExc72jv7ZePb
YYuSHIoxuXYPkXU2+1JOZfaeSoB4SteEv/kfJMMM/6L3+SKsHy9EPA7R9IZtc53sHukIl5Nkd+sJ
bhiyC1qkZN/uk8Mkji13JuDyPdRtgsixBvRxFYJTnhytxGMkrVEnJvR9pljQN6M3mSUoGV9liKa+
//n5gpP9eWPpJWoBdulmBn5Sa8Uf5Wbjw+nucHV28M0CiZh7nrfnLi1NgpMwjVezKrJUZ9jpbADU
cj93uQ74VI3jeLhW8d9NeFiorEz/mCb05S5z6tEEPkqBL4J29YdnEGUWsj54LEEkjvmim5lr5xQY
xQI7V0x5FxUTx0UEEEzlRvcQm3PSK5D6D+Qfhe0Gfs4kqlBqG3mmniuNhQpQkb/Beo9yu1JAFvIm
hUB2KDFmYzYSjvPG8eXqdYrl8vyJHaKwB6h/XEFTZSAeA4vP6PTcbyX1I6EaAinuCzy8tcorA2Yt
1muQ4lNIz8kJ0Y+rUTuwvmpfLJvNg64Vb//3ISu2dA0TtaDltaH7xL6Zyi91hu9eVCp9FwuoDsJu
pj6fUcPXqd2LZMfE0T6XSbeYTPxVgzoynmc97EFxkXWUW7QX3AWjqvzXiZx/ZtPds5Du047ZyEJF
dUsEE/GXtdeBvx3P/blcbOO9ZRtndWXxfK6h74o0KKgmuyLYAVRSAffq7xIvTN04twU3PKma5s9B
LQ9s5BZECQPiQlQ1rZ17m4QhAyXlKfCurJPtRfI9cO4027QWWbLnns600zTBfkspJMd66cBpEilj
lQBcn2yTDjr7ulvrkvfwlA2OV9GfrSUU23m+LINBFU2e/bJ5SfmkHcRS6/gZb29uVs+9AMA3VOty
419JD0CPrLUuX6g+/Y9qZj75kWO6seGbfNUueOAluNgkZDGNLM6d53sx96JJssZQ3AkhCmkhFK1h
rMD+XqT8vcxdh3h75huqgD42Gnjd10qIRny9R0mX9xtQN+ZEK55HhMfzR1U0d43dG6h35tjSgSgr
kPv3k1PIiTqHof0NZmxMJigGeud3F4E/HM2QuDYSJJz7qhwszyjkJKbDVNmFG+K1zT8scaQ6KHLe
vD7ja6H3xpaqHdeJJ+pzLFwlx5Jx2LgHEALMmJllnebdlQIghNWn5N2X+Do5QlpSMWmEzz3yCs4S
FLY1OFzeXLIP6M1R/yiqi9QsqlR6FB9xHMyvwOcsNJDyYSaIAFvxDtFpF2kA0JY3Xdsn2PP/l1V2
RU0ivfyE8ZoKreQ7E9NbyQJhaoER7mxIjLGFxyI/fRmfZQ+kzU5NrJGFBr3iJ0Jk1wFndxtd3GK9
8oBR5Bq2e+2zcwZmWdx1zSt0N504Oe9WD3sniz9WQnq1IpvA0EitvYwT6WhI831VE6IvckVRQ0Ct
Ohl918Hkc1sr6ih7T7y947/v6zA9ladlJmviEAX50Ah1bE9eJD6jNVC0Cxr5RZhMM+o4+f4HU7HU
pclqZqIYLBtsoPXRJ09jg3qB5oCPzrGCDS1J/nb6ghNUD8gPyT2XNkjHpd7tBGjr9nb/xIOE9xIn
68ArgxUec0mnZILmEbdn5sCeUO0El1xwE29euvNo3F2XowXjT8mFC0t5oxeqQvckdmsVoxdt1CLi
I/N2XwsCgiYMfPTsjAVonuh1J4S1dPXcpWKjMWHlqxB2zvWUWAFkKt8fWCgo2eHf+wIAEjMsxx2l
IuJ4Xdxq67fnO4USHCuTRiac4Ad+sQD+M2WsenRGrRk5DrMhVVnthKkD236c79bbIAQi3EeVPH0t
piUZiN2D1qrdw9weMxQfm91JMSppq8ZkuEY5WvqvI6hXEp/KoumpwvVN5L1DY8fs6pwr0AvQjnX9
+X6QoPGyF1l4aawr7BIEn+oSxyhezra5WjSVqoWJcGzzq/3NdUjJtsNq3Tf3d32i+do8afGWegMC
uqa3m3/Tb+n+6eurfP6aNYlHqVu0zRBTE6mYydivi8B+lZn9jEJW/TKOIpPnUCn5tMPneaUauItb
w6CDL2mQXxzPhTxEMFupksFspPzbc5yMKSm4PEZS+E9wRKeA0MTWaBX++oEmJINnCoHjuDsuZiFP
v/p6v+7nOJPDkht8CXoNC20IDDLPWKLw4jrNfrebBKlONorQom+fso4/SPvxTqNh6Vo8ywXpER7P
nCPZgx/VgAbpUTwrzZPkOuX3QZ62tZdGJkQZHkO/BU4Rj+aaInEBReXNPttiDDrSjb06JxTv88Ox
onmPhDKhWylU2AudMjdEM8IQSwE4zhBtHdyZkcLekDwx+QpjTC9kmoywUBMLihlm9G/JMaPFRGAb
UgqHyzr2/cxu5dtgzWnDtiuhxK+oMpFBt9hjIVh63IFK+uMoaQDBLn7Epfsgs2lL0du0giJfLJk+
67VeiQOf3ZVgGa030osCOG7QFTjg9hIPFPG9quE334N2NZfmRy8gFB8+1ZuHnyGVvEUXRFcHqI0Y
u9vQH4swV11DnKcPLHULaDct/o6IS+IkiJSk/r844oMR2R2oeT7UafvLMDAZINJF+qTfaN7/9tJH
PMvoVUMLV6JP2K6uL65atS9XeJQDe5fGNpVzIg0HaudNG9X7oeOZK9BfB0Ls94307bBV4+3j+IMJ
ZlrySe+N5MwZlX1z7qSqX8z43RJ6b1eIEifq9r/1ME9v1ZuxfkvqpdSzNks1jugRvi8BRfC5CYhB
OdPJUqZy7V2MXK6S10j5lKMIpAnAp3T5klijVYFXPpSY6VLHFOPkhu5KA71e4yzuPu+t3yRENROT
jskZAPCs4UdV4xLwzcnGFr+oCDOBF6hKa/iyyLys4zXkQjbaEdSdC/TIR/jThyrlNKwvPNKYFHsv
yTKQ/rQ49Ev+j5xZaZIYu2hgmTIqwAZQxdKr1CE8FrJFvp9mFLXHrHiqc2XAPiTBJm8WvlaydATi
9ajYn+cTCnULl+6zF+z/ePd5z8Em82jQ3S975LlUpF3gqn7s7sg5zKf7ImU9lAaCfLNtnEWFJbpa
el5eYHkXsyOum/+HFAr5rf1oJfaS9qmBDFoALz3cEWB+3ZR9EopSQ+NDDZfqP0ZDot3NypU8wfS7
X5zxhMCvcTnavdOKaxOEkIwQJ1LMDl54AR9NaMXdErvVPSnY5c0a1sH8nBwUol1trfeNuffpq+Nm
BKvX15GP9iPlmwd4wHoLsBMeX0VCLzLHTGGoFFgpznajGx0uAC/gqhSfcRILA59pvbBigvwyLb6l
Os8KP2eF94K+YxornabkiAO4ooRRbNq31gWX9VpSvrvIA9+Ch+WyxwHHem3MjCsf++VrfK7W0GNX
n/FZA5ckSORN7EqA01Uqd2N0+h9JsQ9E2mEJMdQ4JAg9/WkiHyM0cqynDKHc+1SdLdQ7AkYuCABW
cwo/PMpCnxVPyuhuVQTV7Qcu0yjvwOEu5AV9R7tlujz2/uB9iI1c9TwQk7PIWBHrCMJlGjLWeAZe
6fnpSUh7bPLObVKdaiZVzyu+BdBQS7L/WlLyPI5eTlE5NS7Qt3jmgAFmsmaP2GOlVKIiwyBRN6OO
jkT6UZg9EYUvyxhJP9/SePwM7C1y90Kao7pzSczzSNg5n86AzfTsP+hfvcJiKMiBsIFtulwpyHdr
svMAwlReeFPaMqFY5y/Rw+5TYPyMD9xxzaOfKbA9hi7DphfNeAISL/rkJMW+rkB7xt1MTPp7OR+6
L99Ja05xxzmg5f4yL5Y+I6YvVKyUc65iatTG1iXRc1xzbkpyPsyD7rl/ctGGND1AOFqflnvNHkF9
6PuZXXRDKluvas2QyvdjL3rYLtdgyggEZpPrAEfZNBpqyD8mFbtbhiK8xLTjDn5ezRI5XX3cwqOa
FX9SiHQYUcM6UIJmhND/F025wH1LElnG16HrKUduyac3Gcf2N+8H3XHpMFSOrLOXn5fUYYHbcnmS
12i2pChgFb3GaErzWDaifFRFdG6n6MJmJHX7GCqDC4Ap3oKw7mpGafrukdn32cJMK/HaEUApXG4U
QnPGSFTR7qTCtLUV4HueHll4rzyfypLELjdY/AzDxWquP652C/4HcxJAWNcxPwWeeFudZ16YebDy
VAwNTkXV3s/snVYNbUk+MOIap9dMqsWSiXASmNUDZ7D35rEvf8/7LoxhaVAEfxCV7aQahZ8BkFpd
K+NefoGkiwE2vlm/xLhuD0i9Gsd6IIELnVcqn4J+jj/dmFaAIHpWySKFZg9X
`protect end_protected
