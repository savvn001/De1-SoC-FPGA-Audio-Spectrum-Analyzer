-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hk/2ABlcnPksLV4nkmNwi0Vy5viiCeknEPWRxkrV9/68chFi4m7fFHb89xZpwVej4Y8FVyR4pZgB
9uKnn2BZjytR43SYvl3lujMveE0zu1m29s17Z0ISaU6kCIXGSxdhSWQucGM6TVrAla0kNE4S48LU
IVm276LMf5gqvcfipWQdpNz8degOlolWY3wvJ0DhzLI2Rj5Gj1gA+/f7tNR2YOiM9z+C1FvPd4G5
vGzEa0PYqXx8WihraoH42MevcLxAyoTHXgdl4cPR2HzElVP4TWieRtHlb+nAveYYepqzPKCysDwv
pJQwX5ORWDAW6UKOw4qGQobORGbqcn3TQjP+9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
MtXgzJtyJbBIFWi+sjoKbh4+16kPFNDU8v1p8hGHpDhOGyOVrH2R6lMklYcZcPKB051j8Ww8GA2L
6kM6PuzuH8ngQd87tzaZNbli6gyvzxPHeE5LbAGUJCayHHYTsnxhqXHNxtWtaCHUDtcCUfPOyW0W
rUQwPCiRS40flUXo2qq2umPBRPW4Cj8lx2lKKbT+kirEAI1a66xvtSDtrG0/FWJFZnlvQ3+FLArm
GDUIdDZBjK31SG2zD3c0dcDQlmq7WroLutvvaN3w6laOaKLy97ug6MayU2+f1s2v9910zjMyPjQQ
t3peJhXD5yziqjS5nt0CR44waVjez1VFMrphvQAlw7Ltx5+sw6lVLHf0OCs2MT5WqB6afRwulgoU
vFXzQ25ErMUstFd0KAipaZvF0Nli1kGS3U9RW5+4UFzCOkkIQwI2/wssB/Q8/X922r5ssjbX3jJ1
RosZoncI2INduSqR0ur3iQOCn2pxmHMNrVGYihO97DnJjZbWN97B+jKl9Sk8ZBRZgCdUZmIXJG07
nA2FB7c93kNY2b6fgdcC6b47/TRFubmWDAKrYr9Za9dIYU7DC8qHmjsdrqKA6MvD8Mh53LbwWhX7
PwS1ZgCzAMW760AK4Fn+Xz/WVoghjNP6wHcLjIN+9iDjAVt2l6Jq2fv26Q11PcAUfzqLZefKZy7C
Wkb3Ls+I5jW0EtKQfeVzqcz5cexhcAb4CfFd128fHeWUZHOqdf047gYj4ZSXIPU5gvWs7Sy40bZ6
6O6uo3lZeeklW705VVfN2dQMlqH/VjzZSXZFAOEE1JkNr7guSyn7UOpirhB78n9sesCmfrALAQ6j
oap8Gu6hmfp5BWSDNXUuNHZA85bvMteB8e7LCBB3lz+3Sists5422T02gB2QBnmrbSe4uHjtyXHY
Et1FRiMlBh1WwvZ38HorfR01GdrcHBl8pswU0DXU+IsDNxJoRDdoQro1bEIECEJ3MOgEEu/tZ5C2
aeIyHw1fs0KzDsRBFiDeGwaZMEEHbFUxMDJVdBPKDnz3Tn2/sDVq7uxYhnIRpTBZsph9c0NNeDL3
m79AMB22qs1wuqdnarmQwf87Z3klKXkqSO56Uxz7mVcidF/Ev9RFbKg6MFjXv4Ghi5rFND9v5Gxy
rJRFWFs7essDFeG963PscBo7vJP4VOe/bUgXTgC1duMbc40S3zR+7tWwYgvdyjMEV6t4UjCkCoFE
PmPYQ6NntNzvkOCy3gkLhuSQTbYzdlCc3xUaU2HXkmYefZdF5LAjUHy1K7LkycDC5vRFOYq5v9xl
fRMfgBcPnKyq26OiYqTuUMG+i+S96Yjy+ITXGTWXiWXX94uSTODzlH8RL7OGBDOfJc5JlxnFnsWL
IS2mF3VKBOTxG30d84l8uIVEkNzR85BgtEjKoiRhd3WEixlLmhMI3wZW7DVAVludYsEYzjzqfPj5
0xDniUUAUZGRoKmRYOAX8nBSq2WiwjIgrjhnmr29/hW6+krKxB1opaOKN2i3hb7hxjCyBlOdqUzi
tBVLnFjOJtvj5U6qE6wUrdR348qJWZghQQZL8H/KFHcRAE930na+9KfyPeRyS1g8mzAfSfTTGLwc
uni+6TYOzC3H7XG7N3/y1vMxGfLtGmaILizDcUXc4K0zf2ZRHVfhGflRncm4Otv8uLCCtJiYmph4
pBb+I33arJZTh/6v+JUZX52mC7GvX1lhUHzYa4Yb4EmoRT4JJAOzrJXoagG0AaoDD9cNZnnBdYCh
uYIzqEykHAMxK9rXK0EugqFNRMXLmSnzvVhxYX0lqDHI8I8tRaz08IqmZEouFiNMiYhG10dF4H0b
IricjrToPNS+7Kk3XFF/JtqhemxO5VJRpIvtVpjaI1vrAzlXlV2PFt7RbsgcsoNYiaXl6Y7nqJWh
sAA9LDhgK4YXFo+bmGzDn2nbS/PTsNUgqo9PcL9oEHvOii+FobnD/26jerPeiXZxm0BuDwqQ+qo+
G7TMclAUbnluXV1A/a0FigMirC7a1B9/fme1vI7Obcgeybhe4cwpBzd14wSmIIFe2HDdLRHaXbNv
JiDmiCWNn7tGnABIBuACuKzEM7X7XpKNHlslnCjt8jp3pvrUm+hF8RJE/92qetl2qdts+66luM7y
eOpzcmFjFhO01DFY/dx2YneLgjZA+2tGCU85j/igYBbYzQnawPJqRKdVRdtbjHjp70L1G7yROkM3
0Usp5PqtE/X0ZD6yr/2vWSaccU4TnvH3ubc978xvj77eo14np+HIYCdH+/xugVm1zJF9KJVbug3M
3fN+eIAg6MQAz8LxhjH1bL8gnTWduQ9D4J/u3W0sV3OmY1V4qe1692HXB7pexPV24QEUyc3fYaVG
Wj70XmVrUDUF5a7UQj/672umqnAt7rnRWcRjAXM9krFcSaOdoBgg+KPsnPL2gTClq/PQqH2VO1CQ
k+chjhTbbl8oaDVTwBXiAcjvUNVgfvOKpmKgwGvg1MjTEIXe/wOPiFL0xOLoa9WOV7mmU/60bqpT
kW+iAexR1NGfPt03ZEAYV+Z91e3xLp4+Btk55zuLUZF0+uY+q5nLa5jBRGJa57/nSw98MbTWqbbU
1/ttAs06mH4pIulNbBZfdYnn6qZ+Ms3A3Pd6/QdA5Fi4JLIfp5gsLC0LtIKLyQDTAhf1w8TVfdU6
2BGuKhufR1jpuW/a4I+464BVLXNp2LA/ldTvzY6cQEFz4TGtBvdhdHmgCRGwTEgR6A3vBw9sD7WO
2SIiqymwmCf5oDVeNibpqUNrGYpfN2MD3ThmGUwN2aREUh8agO3i8+Oc6Xcupa9JFm/KDVAUpchj
ldhqdEtPr6UgqBL1RS8SgHE5GP4Wt3m3qyVnFgR6Bnigb8xWrQFymmbD/Q5dqo1V3XIYSPgh78WN
0lCZALLNYwwgKd48yyD/HSyQRdk9JDzxktwhOvizgEv716BSRW7T8lmXY0pZ0Ch06rgZr5dg6K+o
o4Jf0I3rb4HRAJJoz2V1r7tZvNhoBSyZc8TIZdQtf/jfLSajqJQdd/D9ah/WwkyoD4NSobwf21mZ
cye5Ev+vj8/UO/CPHLDKT3GQrhukbQY23rJ8wK+jVQnLi0nmrXPI85pOAIOrDQrOQ+7x/Y2SKudb
rj/auRM/2Bkk5BdliHVy4/fo4/Row+A6yFG+NpPZewAYcg8VYoXZIqKeKddqU8l9xknTTLsrr6Am
iBuY8hu8dN1g/pBtZstT2glUZF2uUwR/BS4EEOGEC7UV+8RFpC2ZWk+fjy5TG5IJUutnUABwjd6O
Bc22/1yoa2/ajpZ9AW/HnTPek1JQ7D91snXGT99RZ5uAawRF5/2WW5MVqUy5/vJm7vhD0/N3xtMl
+cPjg3BRlq5S72kjGUy5+GQs0TNJrqKOIp/Ho9g0flM5esr06K7NI31TavG6Al+sZPfMzZvr4ktL
6rGDn4rydTDhF4CAtb6InbFQ9w27yBreKHi4qxuWozA7S5c/4eNz2hHBn6S45shW6g0OD4HJ08Sz
uEtRJkroB3m7iUKgJaygTsPabhmajossxDTi/KWB1Qyoozj/1Uebs34z+X8r8o+Br9yZV2djYrtR
qYGcC/QleW1vttjYMmdFIJLycR5iHMFxD52CQ8gwXAlxOWDNDoUEzEk9jJV7HOCuXn2xlLZ6PzAt
TeKOLMx4scdP13L3Ds7cRI5oYTuOzJlbKvbI/RCI84EhTMMd2B48GB0fqmXLHur8YdDGERCHc35x
Ld+bkIhb9Ea6d8ykd2mxpmSkScXdyL424HAcfr/Q9AF+qrjn9VgkgpeEP41gd6gKEAlMISHmsLJj
cW/VSuK5ri0Lzw3F+a4dIoLFBAECLFmFjCjLJwi6D+F93gGG54xnFLMs6FSHoO/NHkMLWBo7fgt7
EMDLL4hsKIP13voIwQ1dTzYLZXWCMf1vrgNFdGt4fC5VGTelhSQwxBWT1Wgktkdq/JBq1lMeU61n
9/uBUeQ0tYQR7+WDh1A1h3E7dRQRYbxWMlwL2WER8iA+XguLKIsQovpducC/xw8TN7d3QREZddod
KnCpAJ5CmKAXiiDvv0XjBYjDTSokbJDcQKTnj55dYVu65MeM418ObZMFC85lJ2P8ren3UNXfK0cz
grPAB9vteoUlKeU9hOOaxQAKMtgdXOOTozNPGeA6dXs36CyQNuV5uXCuulwczuCc09Xz+O0dOd1R
s8fKf4jHY3iSjz0wR53qyrYiifgiJ1x5JcZuUoZqO2B0/9UoBieF0diQzS4iCQo92OVQr9evMBie
k2SRvlZgB6xl34EhFwgy1cP/wL2S/2rlP2aQM5J/ZgCxSvxXbfRKeY8xSPiwG39QvNfIfnCXhbH7
oouimy8oeqq4DH6ht+fO6xSWz0n+DmrvB9/uF8xelUxYYwfSHDNTpd0QiOxYwbF7qoWba2jQ8exe
zUdt5Hq4yV38AW+zru8X9Cy8EPE7+JynDX8tjaJMxir0BUUnFsszCXmkFGLc9z7WlJLyUt3BSg4m
OTA3posWMjr/fhDJu3145d9SOW+iXR3kqPSi4fpPSQxyJKfgAodQ2AdUq2WF8z/cq/fbgbUj2LP2
afnO6xRGg3uU9UjAcKSlhTHEutxFGQ/eCCAab8SxzBj5mqofOmes7UXA6SBsH0t/ZswTZyKYzwga
s5L3J3JaCdEcbOE7N9cErt1mELBgJ1YIyrUFxTvPM+9LK1YVPblNosQ/J6VLfz87cog1YEgSwl39
GibZDQy9L1QART7WtKC8dJUBEuUsl6DAumF5AZzd1WbNsvYfOGOczlLBUxU9NDpyFRArwoYjVL5H
hLApCr2sNmbAgoVnp/FhAEpGfJKCTVt7OKPpUboa+nwXWitotTchYchDsheTVPD6wpGIIeeXv7wp
B9FaBd2DkBuJ2BhlTBsOjyUBwFk79i6oKs0xErCLZFy6VzpfcfEnHjKFXlyQV0pSOYjtZRpqY7VE
57ChprKpqBmqqgfxh+GSt4Y7Oq8cxfONifbJZR8FRxEa+8mgzACMVq9Rv20rrx3QC+uucH1UL/9a
vlRmswKYmZLx++yYTtIYQDs043DSRknRBgRqHP65ll8qjtBgoirKiy1CZgYqQYop5DPIEX9Bo3ZL
U1PcaYVNKGIugxECja14v9yPwERUxDHZGFjSKFI1WSKC9RXsaoHaV4z9lDzlPtfxoepSeteoGQmF
23ldnE4Zr0oGxGA0KXQiGXyrx/bvH4PZR6V9WxiHwK2/Iq18DN4uM1aQCvqFdx6Fqm0Nwp0IbxYJ
XNC10r6IVrbOLcu6Of0dx2M0iLbt8UiDlTmHYWyeRXQ77Lwo4xQw+09wEvD2bPP2ilDw+n35Iyd2
UBHI2azCiBSAS7lbqCAGDMNP4NIO3f8/9uk8kd4L6443MMAiLTV0pDbuHoAny7dqFda4uSV5xv1b
6au7reQWFV4LHeXLt3jHGVmqQOc5X2SzGu4/ubctFlixxNn9/39vxzFqB3BJQfLaEurdIh2WOU7G
c3yiz1olKxfWOQ5unu7Tmy8zW/qq6vREiE5GDP+lhodwCv+aIDeJGmSaQIDcBeKYaOp0qzNo1GX3
7dk00uMO7yqW+vOf7Uq+559pzAUYovGvRRDkaDdHV5MMxuHQsMVRAixSyluW+UdreL52d9TsncE2
IJRVu/0ReQkia1nkXyuYRNaQH0UB/IOoBPbcYZlnBpg+j1ge2yakwrAlKd8e0XakWxuuNcAm1uoX
kHJE2bsU6zvqagmBnrqAbkGWbIojvuzz21oFTeUyeojFnNJlL1Q4y/7wBVm0kf/e7YBDWSi4lUot
YmCjWdrpKvh1+tTkGTTiGvDd/rrY6TJ0EwWjoSORQUhM+VVpOHKxOWOKj7w0lw+9QbTNtZqelsVH
44ylm0inHanIZ9h9N+JrNK7EKagln29VxqLBq7z6muQrP0/0V0bpHKnTsqK4c/7XEgfOdPvbcgVR
oQjPewUjbry6kjG2sSftJbip6eQPh9y4/rdhahte5DtlqwO6iciEqfFRPVW2uoJnrmNzMa678AKv
RG1CcBXJLpMNJEDbFcuWSAXjZdKwG4O/QDx34ry1ZwwS/p0Y6L5ZT6a+4Mc10X2wQ+5Chn/MwBQ/
IRVBvr79QniGP3vOb0x39+P1IsYwNFwQJPlNuMA1n4i/8FLXVhh3ujen1U0mFvwxlMI/WAeYprCB
F7vR6Dv4QrDddumU4fOPMeO1qRp3TrS+TYbqoUQA4A6k5Ju8kEBxAba2aMXQL40yJByEl52lR0x8
mzntgn0NdRsHhPJzab+The9yU/kILlYXh4k/3sYeCZNZ7l6vuLzpz1b/4Y6lPfQ5nuOlot4DprAN
ZLniCG4F+x4kWMzRFDlRM+EHA8vk9JP1UtcX1ZeRJuqGLJQTHc1mpuzSOV0j1XSEVGRUDHA0U7q9
eTZhDPIBio/5buL+7Mvto7inKJUeEqQ+ZTzYilPrCHdqXdn+1j8TCVNm2vQkscqh6diOdVXo8GuZ
gjN38ZwyGK/ia8vOE6seSs1fDM37oTtXGQuBzrIsd/1LBs29d8S25fElpQi7M0P+VALailvkYc1N
+EgKc6I7HjG/zkXGe8x7kLnuTVqUTjOAee4pgAzvzjH8P+u5OtFl2cMjOPTexyaaJN42HxjRmfDg
Y009+afaJjk9V/ZLpks/zb84rOLVbCvuC3ncUmAwbQWMRI9ifo54o1L8Bs3y11u/Lqg6tqbKKAjA
gtDdnf/0YreOrnHhfEEsPD4TQM82rpi3OTGDIeFyLtZhl9L8N2a13UThyUjNZq7h3WT6AlxCnH8J
ZqYr+uNIbcpXmW9R5kxYk0lYwWODEUYE9/7Zj+DrNyWixKyhIfycxMO/MUOn+kZnmQdX6u/sJQqE
a9CKGUgZfxPebR3dyvHNgrzJZCu51Xkba43+BcC25kZun37OSBkIJVMIuSZclnZWqTMKnHdNu0/M
iYTAXS17hb8N8JVmHFxW4MTu9TSDyJdsvU52e6SVUZFSqgwE86wAMrtlVBNiH5K9RspDIxHwnEHw
VVauQM9ua/q9xJ53p/g5eNkAE3sNh06a4fFRbsku9ZAiRhdqsxH/WYizkLCSJ/LEvMjGBrtTjV9S
9hDUnxIbvZyf3/VoYjDog/WMlmePaayn1CHdLO3I+hy9/Ktgp3bf3ggQcuDiyb8od7quiRT2nK3H
Og85tvdq1oV+r1GtbXopt6SjA46lDxdmjqg7niwwrQQ1Xc+yOdxiNeXta8b+oRtHL/IDOliXlIaX
afsSb+xRsvcqBckKSy25QY/ufpx38GiC6n8EQkJlAZ/WdaWXQclWAGlTzCuSRMoU0dVrDlij8DCc
50ySnSQQUS2djn5cnPTXxclyhlRbq52h8YkuiDh9vb5i15AxF6PbiGELpgb90Tz21FrJ0RYgUK6/
0NVmtbWhjc28wrx4PXGSwT65IahmGeTU/zQYBXmjYr4riL19wCS1Trh8FUSSZD5mNNjhqdyMmkgH
bYwmrz+06w0BFGF7vjfIPJRzXcsJ1RsHA3w/Ur/eEEOVkT8u98FbG73o0D8atlwv1bh5UIl21kH9
4HSOfuKtDybiZbOZb/ZKYj9Wkdp9+oY6SnsqAvkCVpWMk+hNtKX3ZdGl9Ezvid/LKxLgFdkd7M3P
u+yBoBoB4jdGlX2qoJ9OOcDLm535QcuxIjQhKNHFuJmL1dEwu4fWmWpzqznoOuvrNBIcFT7CZUei
BlmZhFHza72lMZZva35rEW6/vPHCMJmlAoRsrUkbvzEG/pwGouXTmM1TMehjh0mN0K5Zy6+UtTWh
RV3llKWP2qiFVoxGwMg+v5TzBSpVjAnck2slleqvyPBgG+KlPT/UCgBnTOehJeAoBl7YONJezjgU
TAwv0MkFvSeCv7Gs1f4SQZZFgtOVbXQaNKA138KfP/LNfbHzTwpK1bObqoD5S2vsBjTa9c61QU2V
OUqWxMAMQwnv2Qe4Le1rEjOQz0V7xqd9ont2gMt7ik/Q5bCb3j/+Aq2DyhWAXrdZQcpUbY9bbYZf
QuDifgUDSgfoIEdx2VCQGcnOAfT43SPh8v4S5oCBPhquVn5kPKL02puCzdu8k/EnFDTP5Rj/EhiY
vqUoko7yiWkZ+ozo2Cr15Ihyh4T3pzWZUITKXOaIIdk6AwyMioJcIXTTjns3U2BDE3/JQ3daN114
gFQv2oEjAxoHQHK6YnZjx1oP+tdrM7rR7JhlhOAvG4IxMIkCTrnyG0hjvbgY82fQhIYqahZKTwjm
ZA6p+gs7ROH8P0kzcqWQm+y0MGJbSr9HDbFOaDSvWhYYzExPNRdKNeDlm7xphnC1LJeEHqPe4BtF
wh28aaY91dvwzCGr14C3rfEwCJylVMIbTNOQxCCjHgq/jrLRQTfqaB79EdfYELhI+oVV4edu4EA9
GA9mXgebnPidhPllDAonflhObTp+mfZiUvbZXbcILi2Tdh30V0hVNVPNMNjKpKIXMBpiW9WKSwOa
LMgWrQtUxWJ2yxzP/5y0xWflC1wdJogD7WsPxGMGEqRmuogSQHl3lHOMwk+EborCp9u6x1mVE6E/
Zbx7MXztthQgBGsmYNT5dGYvS2NWPbzfRlsjO4Q5jr+TrodtCF0zSuijEewdUwd7vTHhrcugM4W/
u74JUUw7fzBVpOVb6/br4K8v9lxgM/gEQXTW4HApjjPCOuaJjZDiadb6lHFhe+88CRWZNAzfAbUr
7qhg2CbCm4vkovVSawDpGeu9Cwhqo/yokaZtI+BhygycZGA39j2nq8rEjR7jhwIDTzBUozuPuO6C
lsuvf0wd5ee+q2WxtvUKVgVZQo2c9KfEJK2PmrdVspz33es74rJFsBHN3zWxy31ogf9wE95TXFgQ
CaZYyKB2ewM71pREr57lG/clTDIZRar69ej4B5ITQFJnqisN6tR5lvBT3FlSYwuC8sZUGRCwhWPZ
EJMaky+2l0PTVjAI1eBbvt93/rknO71jtDd5XVvR0GiIYXt5ok6TR34Y++NQXI8dxrBLNOkcpuvf
8MyRQuq8OW0bCKg+3NqXqN12mDcRqSRBUr89pjSehzlLVj3nYE0xuVcPrdtVIe4KU9kPN9b3Yltt
TKKBQikazzkRjIkt8Uju9uY0AxCW0alrYP6/a/+ipJhIelAFuyfsKs9tH7d3MRDnTgQtncbMm/Gi
254LtlHIn4V0rCmWnV9iQXq3HFYYG54pELxYuFOHjJyXHRsccmQUzOSLLxzdj8fU9i1D2heSPjw5
oAT/7dK27sHFpP6LF0L4XZBtG0whBquPlXB1Ec0l1/pzwbCU2ce6/GW3myfNbXduOy7F+uG0gCTo
xUN883row7UKidZKbyoHlZLl5Yh3EGVmV79ouRJjoN9BQx6Yqdi+bzjq8xiiZKxg8nrg8VNNagie
Z0pqToKmDz+em4ABOcD4iMPUhH9ilG/0ExDQDfD6zvRoAGG6Rbr0D4feCcOARHf0Qv7AXzcmnBzY
WrBr8xgrK4KljcDCZ5BmLGPOituy/cRgHsdHafvP1VDtxWIzcN+DZu46bIlL3luye5HniTqtS/G0
j6uSSjMACO83QsrRGiHPVykteoypvEjkuimHMKTwgSjzN9bKu25lYDqip0wKGS4tZRfJ7lQrqfev
ZWFQTUbq+mzRfmSkI9hyQ2j9+FiTlN5/mVkOnW65sqBtKNAuHBU7r/9M0shiINBsl9UNqo4GAwGf
MRiiNUlM7wzvqw+Vr7C51gG7mBmSxvTDSy/maDC1xFp9Ht4QAeI+cl79lvUah/7s2dAkuqymaIgo
W3htE++njhh2QlCRsy3KDhaWM/OpHsrUt34MuudAjsdBsABBodsnZAc+8GXkIubNUmkylo2NgOBf
O0Zsk3SPBbWA6WY06eHv1CILy0cqOaKLoms6K9I6BgYx91cIHx7XeE7N9rA5K00LDfQXDQI3HA5N
j6880jQnF4tOIIX+IpzNRMzyXrTaBkafCjT/YoY2q6YgykMzu+t9tY2XUgaC4uXgPzE925my/0kH
5URqx0r/qEQtuGnlcWOLtYC2XJ6eH5Ox5k/jrJBvHkh5AAQ6j8N4Wa+hk9xtlTEZx0AwdoBxGRX9
zXjJDkYp+uTsdnFwr0vsd3fhxpUaEfnPnfP/mslml6DDFopvnMr5crRq9gOYPRIIxXyF9YIsNqX3
wZkJzhJQuW/lL6E85CI4yM0/8zNvr63o0+1G4btpiOHyb+mvKjlzCliCdsg5sVMD56cAjRbS/ZyG
rYL7UIOGUqdONE5EqPv0V8E09aGYE0FLHOmJMV/E37lUEzGjeOw+27LIm2jqW9IRApjyHvZwasEi
/+0wIOAXeBImc8fBkkJbtsae+DewZtKuv76T2/fWJ4thNM+nFpiD2xNR+mZscxem4Q2XmzdmC2Ee
XacU03HvJTM/b4uayl7TizWXZYqKz9Sl+S1qfPS/5APSylXgmzthi2wQAvydhNzupdGrZW2RLBbH
b54f9f4bqkvQIRR6OrHIUPF1HykSeq/Wl4/1+OZI2mXRTRhR1wcZq3Y86nn8xbFYg1Xn1kbVgZRI
NbTPhkpGiOp0xj2Y+l2xQHEp/n4H3pU5HEPIpnwHKOZpSmUQIe0aToBKFQSUK6mr6K0OCSwApd65
XQk7JvOLiSXHE6ygDvuDn26ty9bk8LjlocZQwteEumiqsUAnb1QOHVIE8Mwne/0VMn2nhL4CrgVu
5C31jFnEDxCvxyeX7ANSarxwqEdtx5VNYgbtzUKMT+YbUDz91BUH6XF1qBykr9fPc5a8PIbRAsMQ
yYy4Sz7X50kNvrxWnLR23droj28SCSSjQ3lHPKfvK2FnCmEhWX6e+FgqB81rqKDuZx5s/BiwoLV+
Nr1A6wsRkGGEnIqpG5bZcwtDlH2NroADZ0a+CIcCwg8tyccT3dbLFY9yWU/V9FRGBa/5Fb7yeyCW
GyQV/SkmYoxo/aFEXy6NwmF8Eu3TUC2BonuyNHchpdbClGgchyAau7Zttfkc6pORr3sGabLaEPKp
Op1iKd/5CyhZn6sANg4gSJlrEJM60ZYUf6WaWJegsDAqOpLzvujayf4odraOK3W/w41Rf8p1GD1C
9wSXVsBxmxdkSiXHJrARJpHeukGTiuBgNZ+YQ2hfnI8tf7EknmHphVUew+62pyIMGqKZU9P9RRXh
gptHZIuWJsGtQG+SsyoERmHO86+PphQOskxgnN4H1vEfPH0Vwol8SDA/qrzg2N6VE++uwf8pc0xY
HIFWZvM3DB4VqUalWmckl65uz66jHzAu2l3qWqnPz9vBClBzN3u+TC4lB0gSUFUIRdUktzKd0AEk
80VXf41ySwLfcwKmH8WGAnQbynWny8Jbeqqit6zz6Rc4SnrLxQ01BlEVOS7zagGazykYDrQefzM+
E1df695r5/W5fvnewAlNSd1jdEahG4xPD+8+sJhsOKx3sc39Ucyfe3/CNVkdtMCgYeQFklLi8ynT
HOwHluY9WNExNXhsygdkVcGw3KpbjBIWgulXKtUv4jt9Wh/2pNVOWbb9QbwRPBr2ezpDRKHSBkvg
b2pg08pZE7ke3Zu4QRN+ZudjEw4MoLSXap/sO0xC5Ug1iYM0FZ580wDMNGpdaFDcLN+4+gKFzA0K
sLphPte/nS7jjH6jbfwFtWRwGsfkjzLbtnu4qQhW1JZFoS/16J9p/Gg4wdwFxc/pyXDY4WjWtE5s
6hHsfYCBCt5YiYQORoGSRefM+y7923tdOWlL4KbA156jZ65MRRZh1cc4uxNc5qyFrf9Y6zggwrca
nFBi5XR93O5LQwswjW0BCoNSXkKYyC+FHRSUXzdRijjysXEXqtkoyGIXEHuCd31rnpzbE/cfQ6XX
Kv3QhtoPIn66ofhtya6J/bZ5c62g6Bdkcdtq/wstOm+65s46Ma77vItMc3q2/6y2QGzDTR5RwKmW
ioS5szE0NFFXSyur/x/3iRc1+cNHHvY6HS4vw8s0CDU/sivqOUgCz0kTNgaaCRG7QQBgZvCqWCtd
8ourfu96fxbicz4lJBjvduihZZ+GXm5l4LOcOcURQm/3dmWItvH299RHBnu98LSetWMgV+mHPhas
FAxYGV8bGTxMTBtfAUzx3M3f5O/oJlQ2bBvcC4Fye8dom31ebCDCj6zSv9hoPkFzqiAzhg8i6Iq7
Zwv7lC7e6ux7Eh84tkJt6cWN88kbX+p3SKIiEb0NqBtI52tURA5Xg6/8T1dQQ0fWKhnnVzFNeTgY
ABBwt+Yb+9X3J2bFx2pdLMNZqEsL92vUvlQSGGE7sgnPBBzojKIH9zSoNdREO57QKUWgElnZBfXm
LfTxkkO8d7zcgyaIK2yfkRD9Jla4oT8VB/vx71iUOAz0I2D8iGQZa7g1y1TkYArcNkD8jLbou9Gx
juiY1hm36A1LS0yS4sF1/U0BQ8aaUMOj34sjYiHVf4gtBDbPSdC85a+MZfbWqjMW8w/8Rm6b0kmO
0P1SK6YpMlbAGElRCb5zqb/gUJHtb/Rn8btQlXwifquMF+MH8LVtl9che7JnmK+HdtYutpy7hbuP
/FibmGVnmcmVMeJAUi+8CfojVN5ReO8GE7/Nm7tW5JUri1fWaA+G5F+YcVTKNGRXNlfWTyqvkISq
MDBxv+ig5z9igKaNnreLcvnpAo+/fjcAMtcw6EOn26qM3VIlVhNud3dyYLoG+41lKeCN5HZrCmcA
uQPuZYglcXucFeFVJFi/2UWQyTBq6V0Rk1fZimqHqWcCS9rxxPsNsq91PLBqindhFhKZwCAJ8v0t
xSUYlDP2J74Q2mMbb0RBPO6R4CpBSEaT4eKM8h7OHEG8inbSkooPef00qP4M7IC2MHYiqMvZ8J5c
Qk4wkrrFXHdBe1cm0ch2GDgwR81DZw92neUldleNQPcjKlRy3aPTu2M+y1sbNMiECjRHUrOUPvRy
PFhr7V4tx+bTWW0l2PSNTfTA+OCo3+dStqj/lFZKrHOHJrk3Xz2Bz7kpGX6TUX0HEPrNcSQ4yrUp
+OYm9/WeZCMVewvErk44PQDI83hUbJzoGDwKhFtO9RePp/Ixs4tpwXAmEAzVRDSs7vhZ5vjQyJ6L
wz360QPvmyoVZjd2RyZkktlWtSrY1gbkj2zxgnL68HiRmtaEAQbM52V9r0bdf/3TboOD9BBKy+uv
F5G0StAzFB4K+eTwBXzJIerDzRVulzVGVwGgOqCkzL0cqZwi0UwfNwdDxaLqbD8ZdVYjpN+HkRCG
EeAVErV95jZgbZGaD7jJ2IaOoCpdBimjoQpk3V4CppX6eF+cM17lt7kC7cSID0+4O9FyMhoJMzFE
pWZRR4Xntj8qF2AYRw93j7CsK9T6Lm++b3NAq8gWceZSGbxDlL72ZHADz4wshLV2/OGnKp0zaN2x
K7CuQepi0jlgX+XEa3PBYCDEnNjkxRI2fIhiM5nQ1No+nfaxVijhDLThTOaQ9A79CxR/rT3x25wQ
WuicpID5D837D3d8nV0M/oWEBHgqAhWaAejtaRvwklkEiXxgNLwCJlx2Cc8900kezA9VRwJt5G4U
q1QievMwlsaEmuG8qiFcN9avZQFn7IQrdbRZa1dE06n/MwOPikEIsKNgCCZQI4UGUmiHdUgnHfk4
gFYi3SqQNyvWi/YoIbaN/cBGPG0xJBfk4UUDJMsZUlHQrdZq8jDN3chXL7rZO91fcuzf+m1GfuDS
S069gLDM68ApWyRs+JzqP4EN8Jx/5iRvxZW9++xhH5SXjtvz3bBgRLqKAkPedRqytzmfVx7Ke2LH
uougP7Conl/urtueqXO2jbKMxMKG8c11RhP9MEMSammreqKGa5UNiFGcWDcJRMzOgknHoV8qv4kd
RKhlSyF73gvEpQH73grghBuEHTkmxMboeCpxjXof10jkSr3co2s9jkaHJcxmsXqA/EffXKvd3Iia
zjtetiVWNUGhhnvo7N9gts2VA7KQ+NjmWYdRnJQKxB2/fDhifmG+/+Cr9hT2RD93YBYS3BE72T3C
og7ZgtwZ5yhxVPPQbJjZmPj8VBvtgaWsFQireWtStThjdafr5sXDLYiLYJvr5aN7XdNDVeMRitvk
pl8NENjBemERvW7nlor8+gCcDpXCJ96PKOltLuNIAdXO/6lneID34axFyrWsi/nMGD5+VOxvWh2n
L7f8l0xlW6q76izwGbIjsOlhFCXpUUR4hiV5dRJzrxA80ZtwJUK0lnWGcd+RewUTF5DqpakE0p1k
V17z02eFpe0y61fE1EZgulULSicx0kodxkYoRbkCU7TDuu+/7ghgVzQQ0Cs/I+y1etsmSOJevxTs
N66MUOwR64dQgm65xw4da3uQC4gvweP/lnkV8z25DuNm7Pb5tr+/09Bk6abXv9chpFD5lKYvRIOd
pIVtJ1Lf4P1zVE6uTUTjC+cxUW+r4HvjuRfu5Y/wxlwH3qUNCOJCe+3OMkcfAWrGEZqXCeG3yvci
ppR0ldmOK8gsnXEhcFCKwBMEFcodhk0HC/93D/5gu99CSusKvVlbUQd2SCmOrtB06D2L/OgsXWfd
Jolh5dErt6y7dwaQpyGN6mSLHJz7u8+Egg0enWQt7tCMth/FSZxEVNJqUCCvSpKO28BfoDtpMn7Z
WPztdmZ2O4WDdEMT403SOVB7Dt9gMzuJQXjBeSOdxQ3Z3wb1D4pX3nqUFfPkfP5RQvvYUnL9ueVw
a+wMDJDlUcYzPDV87ocgiK6gKIVcNWjYKlulOTQIxB7RpTqwRGwRwiXo8jfgy9hI2jVKqgyonJ2v
70OXISLtDAf1RQxRFcv8bExxOUq15vwGhmdgvF+l08oFqj2bNN59+Ow435ivosjVdayEaAG+STXb
GXfaRfaOjuZe0EQcRhhWFz0MrFEKAPkE3ZqJqI40qCQD8xWhz6cDLK2MIobsetsWmAhekBuMoy6x
7hCBBpGl0KZHjZwAnuMGNLWZyrZ3uOzKwotpPylIBGfS7/4whqNrcOs3E7UxxpIhUcJcIDZQi1K0
GvSghsQV+Gj/LtZ61EnmmY+1pMExnM66lNoNnNBLo0HB+ddGZPyFDLlK5mGN7tyTsDsA4wJMrg/4
BaPxygztoTaWl3cNAQ/exhzRlX37yXkvRlCh2Ub1SFx6LKIImGzy4PgKcU7Q1r3JUR4JiezaxtQk
U3OHhYMUTFUM4y/DVaJDuczqtrD5E3XQD/ECGcMTwwQ6hrwHr87GibDt8k+JVQET8Ly8dPFjXiaq
jeojwOKTSoKf/7nXRe5bGYxK+fnwIsHLiH0/89ljvG6WLAUgVUEZjhreUZUaz/2V3J+iFJwkOShV
v5Zbe+POfDxM9/WqeY50UYgoXRLjOzMOyUAHVj6F5NQsTOlhfwHK7V2ro0XDLEr54BveRhyQjcvo
hr1Wynq6HJdxaPQBQLNSrf07XqY+fKV98dFNEPXxER8gmYKPyudioxyYp6eYih4pOpQnEShFXdnv
UwCoSnG5NnWOE79dKXWg8RBuVdKbtjHE+k6ym7udn7OXGQ3UE4+aliltCbmX3Wgs0woCTXTeG2qs
GUlT6kd3eXRLcGr9okerh8zIa0d961S6A3Na89BrWw3v+wAu53/B6GwqV30GTcsqO3za3JK3gZ/4
3LFjx+xGDirpHgbyEbze5Dvypyy+jiKeS1I13a4rR314urQxXz3pAx7Sff4CuONDEjNp+PoPTQUK
xJ0fbWd3vmvdPMlcQOmS/FW9JaxPCgjLelFo2/EcCrbrPmrM/h5n4Y60tTKPW3eCCyhjge8ZzQQC
vRdDlegtWYPxSr7Y7XMqvCXWjk7fz6/zgaH9Bg/XXogO5ROJtMRNMlQDYCwXv/c0voBjIxHdNshD
s8877V5jeMtO1uR860MhQdj51hUFi125rYFIYCacAruWv0Jel6bs+Mx8SB2602TpAuuV0Apg0EvW
sY1S80m9UuRMS35yZlC3v5VshczE08mu5HWVhDe0OOMJTf1S1r4pan4souLtv86xUjeL/vGheTpc
0CMkAljMl8mG0vRRKOmYG2ERxK3Pd5xKDGwaBt1hrnIvXta/dAciyyfoHABxvrtdA2GEh06U4XiB
IACXXAtRPCqFzQR+UzqgHz+1lmMO9X90mtgYSIMm9SsRbEV8N60D0Nzsyt98C/2jIst7ytsCIrOa
poSCkJxoCI3UDTc1bmxQo2fBydoOCbJk+RfIEZtE1kRkk0qeYUuS8zhQzz1bCuMiafeGBVR77QXY
ho144wS9W1JTUx+srMsOv9itzYpu5wHHa6dngEUJZxDulW5egAGZdrD1h6kZ58E0at3fydg0ByGn
oeoe3czYcxKCKGptJAZGcEwr6QLLGWMO1wOw9u6W+tf1h90b0piUADRPnyARd08Xi3l62rM5VgK+
LvMS4UV/nZY2ox6CYF93oZLidRRU/cuo0X5RIA6Eq8bh2FZROnxr2N48JQygOZ+1FgsONLfOm6lU
6+k2wVf9iWD8eVLBbvEJLKOrguEFST55PX5l4jSGVOQe0r1QZJEFZvy+15SG6cZ5NNGoLqV2IpSD
6T9y8brIMDTHyqtACROnQmXhwqtAdz27i59yVhnqfXaaChP+IWB6Zwe/eH4UC7ruEwNcIxOmplfZ
jc7awRR4nzZsrvMa5DonbHGmUQ5enQ+VKZikpOlIwmNoZ5DHvHcxqwJZnsPaRG9Qg9Y97Y6u8Wkz
hnjUDEsM2ih1GxYp7tiDrR97X92Sze63zjrRLyqx/73tdbe7NqGWozgEbQuk4QJCMGeLX5PNU0Om
IQdBGY9I6f2eK9+7KwTiq11/5D62P1tIsBOGHVG25yCoQC4GUqiVFzvu1uka1Zz/62oNy0Yg1mYs
zq3ZDGjis1Q4ac7dKv5QabCR1Y9AIhugFo2RaY7uGdPk5vvS5iGPs6aI7daJwLTBEAYdmvOgQS93
R101uav0KRyAxzv0pi+TjMZfj8CfKzW6ZDG70ofefb4gQO8CFPGgUsUl8xTDm/cifApHxrnA2G2r
3ib2RRP8JS3wH+zFHcSmHlzWoImBzWYRwX5/j7Ywom+NlK4900FsRpiG6b1QqeNXE6Ls8Cv6+dzH
Xkv4TL8Y741LEvHoxgb8UgJGFO2OC4SneYyNnjilLOOtmhuAs49sVxumw5mt119O/BdhdRJwN06t
UNPea49OTF7V2FLRJrSJha4i/HwuItPtPHFoNaoLzvHxLc3pAAdvxG8Vm/dGwuutB9NkXgYdHIC5
8EtYDYmyGe46J5tgUBC2mrUzWH0s77kUkho2TLG7Yv5tVURAgrL4Zvunl9I4HG5tGbbEkNWHWJg+
mjcjw2JM4EyGEpWUAQaQmlXGFrpAc1j4l8Bd89qLV7lLe2HHG+cq4oiNaXAk65uiXpc0sqdMh0xW
7JyMHW5Qa6NnEna1i8VJSc2IEaeMOrSiAWk/xG/UVVua5VbtBn1kaiXlq83ix71gT8PTd7psWWTy
y3qmT/vtEwxE4CdIphPqpHoH95jDiVkpFIurZCiU1qtDv15IVsh4RU45AKpBG7Gd2w58SKYRaWrX
W48YX0LXTe5Sa5G4e6H1NzgUkVx7PgipW9tY5sv/vjAfUBy7UUeqRtWY2wl8TEFGDB6O92ESZAze
LlyvM7WzXpaE1g685bNZl5/9ICHt3AsPRxPhzimvxg4/r3CrCTqioO9GG8WmrDimjvV5oyS6sid2
T1diAeW6uGCMXI/O5OkxZtYb7kqA2cCiEd0Mvg0hr8bzhdsIPZn10EZKhzb3wsgcvBqkO2EqcS7Q
oaZvNKgMvMHbGzQbnCMgB4HteVM33O3XCeGU9ryBbVzoFqegE8j3Xe1pmC8KVwnwrHqoe0+Jm1Jp
Ci/h1y/gxQUNCqbbpyMuhB7KF2SZLjKCTcUEBYOwni74UQ3OpBC8yi2ovmxP4rItYPSgCn+oY0N8
ja0z/JaUqtdJEtGS0O4WsJuH4mL6bLUfA1UKQHbwpGGYdz1Ifir83wo+V2+68MMhBgJq/j+XZQ49
x5MAwBMaZtUNpc1ifxvv8I8vc0CBKfiuY+tc3U3lg6znWPqeYg3BspuBxrUQAzOT4z1MRdKLYOpx
FA400dRTbNCwhFsPt/JjHsuky7jKxjmRI0VG9hH5LMS6A/jgUdWaHn/pDhO8Rv1vkgalImYsOHSA
cBqUXZcQnCGRCvo0OKqpCcgRSQesdJ6JZfMmPJkwpaCjqMNVSdua5MDO+b0S8Oeh9cXxEOXJC0p2
ZwLrHBNTQIvLD3L1OJFldGE76k74a5rT8lAbN84QWD+/ACosHm30a2ak+dqJwDlsXAaZjva6HqMG
Fa/Pql9GJhVcma0LJ3qWUMID1jcferFRVGSC3GFzyMM8qxCWPMuTYAUyRKA5iTYR/oywPCgZVtlH
/0bmI3IspSXU7P2iAdcp8sjVmvW1DH0+oruEb59SGrQbwOjBPZr1pdhOPSXttJoMHVF4fVaPicF5
4x7+xDTJ23AUeHhHkbz9ZMBotwl9io69fU3gIk+z+ytupFcfGWmvVedf623NkKAXg8WhY5TEidI5
Trh/ZATj5a/h8YCDMSB21BKGxr/HnDXGvzSfmZwjfppkLlcmflP1kbzMiuhYvgMbfyYVLOfV1aR9
gCXpbnjkeeklSKTQSPSoYZx8CMsi/ZVp3Nlhi6Qgj+wAu8tuKW/eR0ifr8TDb3KSZWG5Wdiekx9E
4WMamzLMvf7+RB83bQRuQlxLvnVr1pTkZH6lzwtaDyzhfOar966OjwbMgpP9JZiNCpWNaYwuFN/w
H76WUqHcbpolyUKseUjgd3Z7FkSrQHHO39mJoGk5scrVJpXP1gTdngm2YZlDnwqyVvUpdYYH1JC7
fAf3bQX5RSs2QRxttdG6ZtgVjprbl6Q4etRdqGHsD6AQoCJuEb0rAgUhwbotThrKp+a1FmbcmIxc
5/m5+Q/hzzMdfDL7vDFiXsRADPe2IdFJkCIXVoKwYM95waTCOy8V5R0MBXS3FxpPNNn3FhR+aA75
2huyALTx+2G8ziKD6KcKnMGWXHbr43GDMvopF+5Xr4ttNK6idQ/gK8JNzhfgs8s0Tn9feDovsbAh
wCsMwe2Jkn2mpjbD3Akp2XXy/Eibq1CtxkXlT6m5Q5izDXYcWbV7OjrETxeRmzMKD+eW3CFo5eAb
FG0I9yOACK9mHPKamUOKO3Fl2+RkAFF2m+27cvq4WJMM0Cx6ZmXeLotEt1QsWnjC+i5yetKYQr9p
NlR58BIXJu9DuRlzfAvLNYYhB7XORk2gsILGJRlmmf+mU2CTz3tV1yw0rZv/d+e+wXjkK2wtq7KU
P+Vyn0375POIFf0Jmd9HJYABoV2JAi6sKBU+YsDt8/A4eAGwngw/BhXQ5pFwXjTtNQuby3cQg2dv
n17cd8PiVWZKJXRex8+p8BuCB9YySzKTlTg0WSACw9RqOz8lXkCbf9i7+Dcpu+vCnStXHh3XKeof
q/kTA49wOpzQ+UYjFKhOnNLUC4iRX1c1skwvfV3kyyY7KMK2CBGM6hAlYS6xhi/7uJVl71Xphp4N
ftKwJAGnk66voVHkond7ItS/wmhiPO71y3MhhcU3RGmID0IE8/PJZTAQF64BPUG2IFo89DNdu5O8
5DcdXIfJvk7K8adcmd1TfAGH053YZcZO8rMqUBm2fRxcHF2zwk3PtUGGfVg6nPZhzKvR/oq5/pa4
62rHjBcgWqRo00k0t3NniBZpP3eDM2iXNTy42qOScUZH+iLfj7C4zCU8wNsa33d1jGx1kOP257m2
/JtsGipFMf0eMnpD7abpAA9ANwl5rc3lJKJVqc37k+55ICa6inc3/xDwIzB8z32+QYfNNayoBYMJ
SqcWgCP1OgZUIy2Gqc45YPegP/8KMEE/SnVLmVHFZhVK+aXen7K4e68hQcuovxtqdXMxv77gar6L
wnpG1SRBOk393UFbcY2BReypL18O6kOqupESirP70N1L44Ev35fev8n8kiE3PLL4CXLaGnoRQfuB
VHAebfW5zUlnsDR9q3Nk2fEd36mWMrRtus0rt/RHf1lMNcpP+JgwQfDg+6ZJ3f9NironihXwhJCs
YNXCmJwCUFtvV82GliNLfAEyCJnv/7Icalg/MDVk0oXUERfHTQ3ABpQGhTA80js16tKJxypl4iwn
WkK0AJobHmdPBJL9iAT2binGKnrErWL+fiFt7an2x6BX4qr3gs1rsdbuiS/g6f+s5DfQr+JEUeNi
5texuSYTm8311pSV2uXqpdHw4DaIMSF5t02ZDBIKyyjJpdBldDXHdAYXkCvyroh1f1nJL3z+mWnt
Suw7YiASV6t+nu8lL9Dtgc2PWt5gSQg9y8Zdc1iSAZT/EQNngoD4SesKHJoC9OQ7uCOzr3YjfXD8
+wMvbUSGNUOJNUd3rls7bS2Y7alsavwuVx5YsyP73zwyBcwu4cRuYoK7MzMQZfDl1SWcwuIiwTjm
nzv0B/z4XZTlxv4WMPO4RZ4KtbL05b0nUvrlGx2wzNWVW13Ao8Uk6P63jJay9i2JzZ95G+duYjW2
4cdcU3/7awoHLeKCKuhkyPRzjWjNA6DEzHRUHUiYX8iysOSDDKJ2UPYQpCCbOELj8yYBlNmkyN6X
qG9Y6t/NUY8z//3XsHpKZJYQZb51PqSA45Kfa3Jn0oUePXqg+PRVvtUywfxHMtSlE3zhLHxt5MHC
rZ1GlCUEKOoqaYZUDIOHgUDD47PaxRY8n24aV8IUy4dd+sDroDL8YFn7li+6q/gAe7XKcutgUFom
0AqG2DIXny9XnO0IZPGuWYojMyQber6Zp6/6EhncjXLNklglMimSbvaPR8di+XGSv5bsbgepxCMa
9GKMiRfeCYd5Zw+Xuzww3nZXj50aWi/wprrShPVg2+PsoLhp3/HgUDv81IU+ZczzNyMzVZ75uDYh
2bjoh/Z7p8IPJxuAm6+2wNB9DY52oesT12P/BymyJMBj8A+hul+06thlnKRU2AnNstQVfItz53Kq
bw1Ri22r97u7ONa8l5HNUv5YuPDtQxAvDDJCmmkIEeEe6A77OhR9p5uNxRqao3TvGx9KFKLiitq9
4/f3QLSmOSaDwNja/Xtq8JqFrBbOGG/GFuTADHPWgiIioKjYdqyBlGXyt3gV/wtiZr3HhFZMsCAh
j6rZ+1ikIOmdNFt+Efg1tWkntnhVyFjh0fma3cflgPH8uoA0IT5mxy/+Df5uJpWNGjCY8ygQf9T9
jQIL3s6OfDHWyuZEBUMwLXctZcnanbRh4XQzEZHzWc+7R4lBr+UOzk1Suj7P5+Vdo0xbclKk1xHm
+dYu+p8Pls/NbM7xBWD05LUDclfIzqjeUvt1n3gwMi+5JcSIadSDrZN6LTbx02xGjMtg6gSuGAml
MthgM8FllZeus8m1EEjZ1Wnenu4a4un4ajl4ONQsO9WilbBi1p4toqxWF8dMYEcN27Z8eC3FeJ4w
Dpi/nZ49lYUU4bdETVsJwR12H1yciVg95+XpZqqQSFHGhuBJDXZtFMN6fNoGHpbxGfNvGpb8wd+n
oX8F+cxgUsq+HSg1tl/Ap94MCjV/U2N4xpwM5dghggecBlHZm0s1XNtnW2wwqC1SwOfnMBayX4SE
TmhG/XzTd6iKUfgL3QBvr55UeA6O16aXwTnslg39Vi92630Z/mSKF3QPmcwngqkn+bngnRi0XGXJ
+5/raqZPSt3PU+BXp0jJS9ZdhYxV2oIOLOqbOiU61crRu0lWOZsHwTVIjd1Ja4IcH2k2UEbZecM7
SqsFVwvkGTIrRoQrPsqMJLhhnyPzVMGHY0TPEWBxfFExM3YYjDEXV4sRSDMFDawFg8YQIvnk9EMA
InYuhlXJ6mr9T3gycRDtBXSRLtM66y9ZMGFAndwYA/1ksTP4DTan9mwQIdQlGCj7mZqt4GT1ElGG
D6OyUO6NIvr0/w7Fre42436elp0KL5DV7jHIKAO9wqP6pDAM7hZaHsJJ3la5el6+2jfxs06l0Ix0
wwVwxFWJweRy4ZC6ile4Zeha+2N60jR9FC42hkh/uJQxRQK22vciGyFemGt19cXb3TrvCDHtORu+
U271RICEfzHcykNYBLzxIiXkkGY60sU8nTsYnuzm8fx6pjEOFDV0/XfHMHcwHWZ+CZ6tV0GCOWoo
pPxN+RhT/UfybEDqQLySuKv/OSD55YxwzebuQWlaGXHS5aROA4yMzp87XBPEEAyZeQGASl899pXg
VWXK12IrqkN+uZxBKppzA5emXfdZFGSQLsWezMMBZD3Xv1TfbxX9MOffHdcTYzPV3/3QluhXX9Dp
v+oXwN3x07+6nPKIR4YgrlWPEunvi27pfcRAJST9LoHF2EHwwbGGJiDcczj4fmSij9iGtb/0AzOb
NHY9gYWgB14q10aopmwBTJf22L8Sz2dpfRMBsQxwiCz6VannSavaAxpBQ74KsH6bkNZAypwCbaP6
NPjpcEpiH1XU3YA5Q6vbuE0gv4SXHx3GuKR9PalkANM334baGidqNNy9aBFs2b6SR6B8mqoph/8F
1bnMeoOWIYLjqhPkuzAVLzkwkch4GHxuqVb+nJmmwggC/dFbNNIlZVnzkBYIwp+EFgkb5zbnPfiA
m9VuBdzzl8Z4L73NkM/7Sw9ybXVdsggpQw1QgKbJINbsYlnzjl65/ASOMVF1kRcej1aa7o5M+DlK
5shpF402nqW7H9xPV9z07ytDMdJYVuCelrkHgR4eVCe8ObWF7BNEQ+y7RQ6X5Vbl6m7RcuyyCNGq
ysvlyQ5JUIs4qIhA6qpBjag3H4tEruInEkwnn8Q2ciYtx+ZGrJFckPIt2qr3OYxPg0HLs+BEoicS
IrWKnM4t7xcQ7ouwLBzm7RRPxxKX1fJPCAA0DVrMCyfWJA2ib4HTOH2o82UgyeBoK/+wR/ejYJff
MIccvwhqJk0cmDJCQT+t63yTyyohTfytYxS5WMYbWa373f3G2z4HgT7eFO5U4RQk36XQq3iFsfYG
x8vwLmixIWx9YxomKXN61m3ZJUdYLeeH9tWTHp+EpQabwt5HIVOK6lNSq1+KN9KmAv1oZVV1nKfR
RcBFzgpoE0Fg6lTzH+7SzHGxfR+y2VhD9YAJO0vMXYrL6gVzTL34pTpxiH/IbzV8SmGsmMn3EJLS
KEY/UAUizmw6PiRY9LhmDFBQ2/tkWz22M32w0AB+EhK5Kw353kNPlybQyuZtrLz9Rtq9i8ekVCcW
nFCz3uSuMAO/YTACOnP0TKZcTbeyTlKko0qkHbIzPm2WE4F8LBJ5z35Uo3hp9Jar2G5N7eV/3vZK
PWrKhuqmOQwW/LdTJe5MGaKCGHG0scB/I2HGX308hJUd2R4fpjhS5wMj0bzOvTHlOzoQ3n3/Dqjd
NYuUi/ygw3p/to4lPoX0lZFxT+sac5+H7qOtmb8cgeFxVi8nI/LnF1z985gJQasObBO9KLMcFXWk
YjUumBqvvFPuGG0GnP7NXR7ky8wzCLCd10Z2slsp+YC0+UJhE3gQfMCEQEZZtGtHXfqk2H7APMh+
kDaZlvdQ72HvNiRZ5bU5/vFpPzzZ9bAbaks4GjtpUKEjAhm1l7OmYYtq8tIOVf6f91BcKIbtT6AP
j8B1y7QrPEBljyDerZH0mnazTWYEF9CekfMcOA9j2WMuOYsd7Jqsigj6rzrvLzUrzj3XVZK/fKEa
Qq6mVtfNJHN/fzQLn9LuG0Nxnv1uOH5THeMUY2dQn1z7XptKeKFzZGiA1uolDkT7u12TFewISzql
qXuUQZmRjcvHiUIERAWkGPE7lNvQRMqZtlKS469VF73FURpLiS614+KDyN04FQq5GtVnEIUIFYBN
G7P6KeshR9DvxTOGwss6ELOdakgQiTwXOpo2Dw5d92Ms/1EHjwPXqZBVULRKr3K07FDFW1cMyY7P
+dadiGUZMZF5WE+ElsKh5Vwj9PeHIAcCVEbWxm5LOqDn7Jai0O7cMwLY1VUp4aOUDjzPqm7K15W8
pzMCr4uNEGTew7Cf+ce+A+5KZsrWygXopsSqKm0sOV65SJCUkssw1Eat4fr6GG49DmJ+iGGThG3m
BXFhDTcLIvlarpAukHR4qXby7HOKA272UDWjMXHCHw55HAZaXsGbisDfVF8OXz1vO+DYK8m6+ild
qAxTjD6QCRw+ap7qv7JnYtPeLZMZ86rmzEQ1rb4Zl/JXdq6gxJtRFExH4IZXN0chxxj+cvJmSZPL
lXSHAJWF0akRVROW1Fh3S3qJrfttD4DpW8284STY63+IS3GQsL2dqU2reb1CS1V/X4CRmGCI2VyD
OBh/Jr7buJK5IeXRYJU5TG4GImNql4aJdzX+S5jSQ0MAx3hdTRZV3/lGT+WdO2TSUrcBQL2YclsH
wo3tBNIAJtQBxKcxN+lbC9iWDRkU/CyugX83bC7/2UlWla2cEKsr9VwSbKCRr12LVt2/blKGFAad
o/5ryX9p4OAdV+RgGNv8GBn1XqIduK+IUZ+vsB2xoO9C6RVokbrwiAg4D9/Fvls6TGXflV2FBEbX
ScC/YMVv1f2DwKjvh1OzJYZwm06I4Gsb0WFM4v6AaTpdiaSRaY4KIWf4PCjb1jIRwr0anvOqyZcf
C2WeUMOimsYC6HzfXrtEMEXljtKw2mZChuVyB4MItSB6rgrfxOFsEkKNnY4d2SSX4WEy3m79Em4A
18hxvsb/+aujgbYWDFSjsi5dfhbUYL0hkR38CJpwZwEFYdDkWVbEvBdDRjGeVILt/pWzWh8MVGnA
NVJjb30uFKoH/+mTzrEhNFHemzgFEs1Qy6cZOIF1zYAGTGG+DZ76D4PokUqOJFiyqhDFl6yIwEni
kXHggRQIcvmQgbeLGTnzW80hu9gtK5NU6pRCG8KewxJn/7mvHhWkAE8DnMPH6M5AwRHF7OMMujjB
HVRWsTcxUD2bpH6/w8L1n4d0VwkRORzVjK0XJHhKUtMtYEg0601tdrtb0qWgDuHuZyixJZ+KDg/O
9GN5IypOYqcCHD7hdkHCMoxmBum1WtEio4dIRXr/E985IhH+f8qyNM5Ds1KGgaDZcpxkRScEfZbG
hmVpMQg3gZZcGLm7lmPwDQUTSbp1D6kVqyagP1DR2ic9FvH0/PD6UmG2HXlF0OhZw+1hWGQnhEIF
Jpba5q10I2FSobXdhRBl3ZEaXpAkAncyST4Sx6P9ukGVPV2FUnyCjXiwtmyC+f6e9vwdHiw2SNhj
FJ3pYBc2rdtJLDWTTmj7DeTAB9tiHBZ7Xj/sGrLw+Aqan+05/6J3G4ib7RDCOGCTQfX7D/e/fXo/
qmDRJBmJ/DdOrhx7gVSOomJLGOK/Nzuj7cJuaf2b30Q+2SIcTZFePK/z0Yf3bahat/r5V2HNxeoR
NYV+7O+QqABYhNqGaurD00gVOsJJmGnd2p6z5581t3PHx9GvDiDvZnSOls42BtFaihWMmq2TzZ6K
3KzWpjmsAr6AzUAcTtBKAFnJUdh6X97Pg3MCO6CZMFWOt81aETgXY2BZavQOjwwnPJ7Yl03N800Y
KOqBTJRL3hQVa/B+ayesgTiGfwJnLLWWkvgXy9fpQ6VDnBUq8qoKXkMr9HmwPgi8BL53dG9uQU4q
nbkgJ6vlQM0Y0ocEUikefphdLznHG2TRFka0pZny6XGD10BLpM7gd0eARZCSnAKu0tmI81XyWcmv
YR7c8QfAHTE2+rTXIZzzDDksu59uwTOyn9nH15Ldz+CqYBmVLYhgko01gvLnKvaluJmOYydAwdRI
QQ47svUZBizESHRaOUcvVvys2oQPc0F6pidMNGPIK4XqawSvKACfvyJkHy6E7+uX1sEMtdNGAa8j
u+XA54vn3aPjotC+6C6KojXeWP+mhxhudFUEnFoGqunA46K6bVwClYrW0xCuWKiRqDQUGatPcnHq
eg7QB9Zwic4yVkIvYFteooMdMpIMX2RswSu8x/PCXTBR7e7THKSyEDVR1niVZT4Dsz4SD3Z9PsWY
w8rRdXc/3d8iz/83Chab5c07tiFsNDf6Xj3qH20bVLbx+LWEzGoN6eKuikYl4qVSO9ItGmwZlEMa
+Xi4HmxMsyUXv+42ey6vKkgB5mj8c82nJ4ccbRyUM06dcLbNbsSySbWC+dhvE/TpSWbsAbhE8Ibd
RuWHyUzAnnKza8q0HXrj4+DH+ONFHzQRE5XX8w4o7nuOxLLLDYTT5UQtBGnhDsJjbzkT2u4W4u+d
pm1idvFXCc9sxJryT+toKcZB/d6HDCYIOiQVPjm9zMRMm09vrHtwf8IBcYEEpUBSxqPmcp3NoMgO
dZ6th2GILl1lGPEIH1EWzUaEC/Uva6uiWfWDjNZd+Sd1IW4QPTjgG4LXsMHNrx2a8MxVxJnbidO9
0p9xSe+Ue+iDoasYkVYv6sZL33+5rBpS+Q4nCYSuW4Obeo4Gc3HVYKk6FVAWBCocLsMbXN/dQ4G4
vAzFZ8TBLKuXTDnSOANzV7HpiXQBWvJdBTxWDCvPMBiGlCsnOliJ/Fxy+x5Y2EejfOZSO1cEHGXd
E/lfUuGhzD/ZxFbljxWfQfywg70t3LzWu6qckbOvjDwZazZW1BI1Wd3MmbRERWH7mUsQHYmCpNKa
9YZNApMQEBz6bEgkf+O3Kfe9SJnWNhuVDJjhOLfMFFacq4/gC0YdWEdlJKnQhwLBJ25mNpGyRRia
KYjWbHGNj9uDvm51+wOfM2YAQZUyZU3gLX3gSTv+Vjti8oU30/N0SqEjivxP/r65We1siIlevGVj
bg1EHlqgDL7um7c+xW9vYa0ECKvE7+4fSZAjaXO6qp8oZXIezAsryiavhYstuj3GoeIhLAYPaRWF
sTXFlr48JlPehvF8QE5cFNYhrqQt2O1vo70hCNA+0vOYs148kGK7nh5+V7asmDLf1m76MQ2L9UMJ
+XB5E2qLX942PpxEjQewT+LDBF19cMJCMwI9CNowNHYpm8BCLWKUMOkIZlgKWg2cvUG79UpVObS/
BddhT0yA08uQwD9KIz6V4mchp/7NUsHt7y6xNYVBFiGxPN3iWn8dFBq2vizxIy8Y4mT60nAuA0Yi
+0hxjSC/bazMzsluj45UypizAtw77EoMcjAFztctrnYkcv28BxmM2jdjQxTL96D3JAN/9z71h0WD
E0oHOiNBcuCQiFimaI0KEv9PXzdkV6+aJY07vcM7eyBdEYJhw8rC9hYZqd5WCaVCD0oMo3PELPlK
lFpCZuF9ywJvFQAkXnT+PjeM00a49Z/MZ2Nut54KyOYoLvA5z/E+q2hGTyWajfuA04kpWYk6wBWL
0Be/mVNdf2t9SETkEVowlYfsVzw1eGwzr3AKVrWxqIbbgY3D2mL3SZxG2Bgt2C3ya6xpKuplLIF2
zk4lx3ki9tG6Fn+J3etl1yv+KXn5B/AC2wcd8fBpiVOM4eTYyPyvog1c/NvrHtTbcVmDok3hA6Ve
pSAglJlTma/2dQ+ikyNZVIT/1RsAPFfMciYzGp6RqhIJFQyCUTxwNTgbr01k3IZnC5pg7KlEKJH6
CaSEdx9BCt8nIV8KXhLNWE50gqNgPSTHvH7V8YIUoRccAeEcNMglTh1ajITemY4gSusXSqFbwIwo
iYofbgDNWx4vrIn5Pyq9ztgS1yuhoka0cTpHPMQPozyEars+KiVUaTntx5bH0OuCR2oFAuXNs1A+
nuaG+YCOsHG9a8+OmwpLV1POO5AQ8Nmz7tE+eHWnRGF0uIVt5EGzwo7oukCpX6h/q2RMmPrFNmsn
W2PlTf31x5Ao4aC1oaiG13hbG/XWzAPuGYpASUPvpLCctavHxGvNBnDONJwW3btEsT7ZTVMjfqij
WZ5eTSQuEoQURRCoNF2k8Mm+u6jArBSHV+xItR8uJtvFObJy5xvVxceCRoJATbnuGUekhjDY+GY8
xmGFREDpi55tYet9R6lmUd+06hmv0db99chYQedsk7yScllVCTjyEhIr1sxyqbyzM71Qcqig6HeE
xHH+8pTPZ9EOa3fo/ahcCjsRmYUs9XZaZ+kHF9QvxRuqSV3LPW59w4SVnmlbIt2AK48r4lke9icp
RClAnjbFIrWBMDnLFIpJ+fbkQ76QpX1DVnDHYg4zxPlRSG4xR74xHda0cV6a2/pRgea1uYK27p4i
wDfDel/5p/QKgDSzBFwAVrUIQDyITXOxbkr44Jbe/QiKvXcCFveD/VCi537xLt9St9XfnU1x4XjZ
gZb22Usox5MGPassoww0jls3ktzgyks26ukA/WBPh/ux9+ZOjdRaqMTIjRib8EpcvRSMm94EIYOR
+DV73HXZ81NwW7TwFA2U58mysRRAuyK3uW6WYsWR9Ym6i+Nk4Vde4G34W4Mx7wcFqgToUmme5a9I
VM8Q//Cb52Nw6yGg/dFmwF84x+SNjaWqUNDcSo2afaiEmvc/EcajOOJL6tmVB6RdO+egI9/mSH78
Cf0ohYH/vhj5WZRKCVHzh0jHEJa5zh65qoOp7sVT83qLrD8hSo825v2xP6LwlmkqFmQEDZk8qyJs
sTm1+/GPd9m7htmcw0XNKUKrLYZRGSXi4JSb3klemywTNyntTCdou7bGVvfhPy4F5r6bBg+QLw2o
jlbMP6B6mEmo9InMDAgKfJTnDtUv6bsyKJo05+QDH9Es2gCzhdP70Y+wndldLq0cMHX9tWaQwX4h
FOiy2rD/X2tJTW4ovawz84R9rx/hL7//bR+65rQZvpyJhJoCg255F76OHNeE5tif68pDYNioEaug
JafarnHO+lFof0YcDWzT2KVR8dGuECtH2VYLURgSQUS/bSVFm6+j4AHPKH5e/nCWQbK7RwFGxZnB
/1g84lzDkpRhU2JtyP5ri5OyYT3zWtE9nLcuavuTgChYf3KSP3FS8R/AORn98lvYaW7dfcImkD1Z
PK1KTObAu+BTf2eQ9DrC2R7adXoimMD7Gs0PnVP1raXqraOxbQGa65v6TwgeP31ZUuhgzqox73Ot
sSeCMJiVGdCFbmgND3yxVLkfQFda+yCRtecFdhd0EGCpudM79yZUnSEVIdf8RXxB2h03DUdmlSAh
3MMxiCGOe3moljmIM5E8SBpJaW8qk4ndt3HbLzqw/DWDqtfWzXMPHJ/Vd75dwCTITuF7/JV4B2ki
Y4MoKAcTRPedOYSIBKNqHQAEBnZKQe22Mxe0sADTZcagW8hu62btTB3tM9LcdzGepCvIqPO81g2h
ywcHH/pUdMepnIasIGbcOqsT4sZK73Kg61skW9hkeQrI9DVsAXP9wp/ZJCWE+sRAgZB+wZP2lw5o
FpbWf0uuZ4LM2Zqw48tO0xUe/fz0mC1mhpz9d4cnjOjvNcw6BiKh3w51I/Ff/UmFLS0jWY4cQY57
rZIbRkkzR1rBTxsviGbexnWs8dKZbTT9a+kh/bK6HDGegYqq9aIaAMzmZ88iYtRJawmAVisTafla
uaQMAFQDQ1qjQnFbCnUxy/rv7WEY2etbtP3G383q2hiPOgDSuDcfAYs3OMUUVSylBSTvnYnLBNcJ
uT26D5RiF35zxQJuxTkCQEF24cSubV9R7Bq+238HcnghADfkhMAuYKLs3j2XTihXyDEtlpo0Treu
R23KkMKmVzEUMz0ejwGXa/L/Y93+lT0PixKaVGmKjcuQ2+icnOj1pzSwclhJYVvKpkEwaQIEtifD
vKlXKIyaql3qdr35/kOXThEcwLQX22tU7JW0BFk+dc0UlCygThdvisuv+CR53KPNsE3JAOzDCE0E
89t2r3klInlJ2L578hgFraidkAvwauoo+0rFEBEBU0uGXpmYHNhIZpvXEiAJCmYfD53yRDS+mGJK
ViGCjRCJsEIC+QNSrhfkmDejZfozMX/y8n9fRuvoZRkv28FP8HoBvgzQ1K6cNVvWoXeV1WS8HAeD
TYXpzGX3qeW7+9gZyUO31rozse8EiWHbf/lUh5Xp9Al7dOindArBKk/40pr5WKCguUyXlM+eZlmz
/Wvvk0+Tzud2s0fabADxpy/ZvQ4orskFkSTV+ezAgrnAS2VWJY1KjNTAFgxqDPhWuPR879pKNcRm
G3gJHwp+5g8f36hhBNFe54RMWzgXaOhxb/bCv9dB0t/NNrjgsZ56WroTa9s64SoCXwEj4y9Y6YHY
tCZ0tn/nXMFCuRxvuEtejXV7xizOB554Z+q/VTcrMxzKn/vLqR0ewjP7sfgL+XdzC8IoI+ahvmuN
pYEqKXjR8jtcgPsWqISPy8UKLrMvnY5ewo8N0yT2OA9aZL+7lYxgiD5v5bd5ce25qWizIgHdPq7S
H+sCB7Vy8CXzdwkdYscgEcdf7yOqXzZ3d8A1NivD6jTcxotMqoOB1PKGS7k9iKHdJ/XqwzUpZqzN
NUYeTFBEQLDBeVNghM4aIx7I65J8LoR6FMyTd4x+fjHw9p1JiTLGyJnsEq5lXIkFYPksDXZSoBA+
ddSShurMfzefxPS0CMDcll0ZD1eIXMNZmBXlKBonSScZaTbmZVQtaHmo5JSSczI/Wm2ueY+MLHku
u2o3aj2qbHkldlfVuS6Z2Wv9dLqmrw6MdhrmIKcJw+3CwOEoeJSvp2YWw35khJvlQd0+WyWC0jFI
4hUelbHBI8LUChaGlf+ZZk7DVqQQqK4ESwAQDniLdRH5ZnNnsm3RLwEsIBbMThXZ2GPDZ/vl6qvq
ZWK5TsvuS+MjR9yihD15cgxYNBI+EOjGNM3KGCYsxOHd0mi2Yg+MfjyGQ8mD56RH1IMVcwE5mJbA
HAbaAPFMJi5JGDkyFoCDKyoAKXsTsFvnp3ikPSBtZyAPIS+tBOG7IEpfVmCaf5UnZG19uXXvgzH+
8VHltkcj7fdWNgj6kjQKk2x499w5k6fESRnS9h/e6rpRURKYnoREaCeKPzsO+/aV2GO/2zj/ilH3
BMFsUDx2Nwj0nmIctxBIh6DmfV5EQYmWnZYwBduJM3h0mD07A5mvHEDR6D82vUNBhT8HsiIrBoUO
3Vf4vtEBVDK3PJzI/1f2szsk/+ANz1w7PEbvI1vwgUGlng4wFXXwgE3JtCrVHBVGP+CRWaJ6Tdss
8vWc9ybtmd2Ky9UOcpLFGaeE17Hjp+N9baneIkuoVniMVy8n7SRwWrYcshA6M+Ag5fiAMSI4IYjH
PM2MPjqBPF4Z/0wG1qF8n/8vkRBLvNKePLwwsI6kXo9lnESDxjFHb5dbB2t4g/7RX7tl3nJ4T2fe
sF6RYZ1GX4S0s/YJGfON5snowTzqdzJCYmLZM8gs4iguUMR0GFzImC9WT/IM8zZH+ZEk7EUS2ktF
u2ANI2FoNr0A09wXW4mXtyHNzj2YXJiXEME4q3nWizFWz1OaeZZgL4l1i0QD3SQx2bxfLkCK6yp/
Etamhi9sou1KHFWagZu3KnyreMOxhMmat9+rwy9LJzrKOeSnzlkYq1penhaN1QJb70vep6nURIQi
x0QGltnJzl3rwNd6R2+lCJAHVQXkfGH3bgLc/uOC4QBIl0gF3CKDeqXwei1OCnL6uakf2F1ZFVNs
nz3JPK7pf2wzF/ACCcD3PDYGqx2+aX98bXBmOK3N4ot6ypqQ0sigarpzmJ7mmPgcvVrSq7eAeo0r
djFa1ASK0AbwZtzbHugcaPipyetNEXvvfm00LcZfu8ZauW/imS4H4GqrpiVv2l0FovhU0UwkI0Vd
2dJhSBXlUpmj9BK2eMqNniRmDYVK56j1FGVx+wswADAF3MbFxaSJm9vlScwZJoHERPuirz63OvAr
5pdKfmeg5PcBOrMVdpmudljnMlzDO1ITKvU9F6QpL+cEpa5SPpF45Cev6R4M6q/R+NKsmBDZ2mu/
3xpSUwwynTCaTToyrF2Mg16MQvR8eNmu4e0tknTHHIP7dZbxgHVCn6bHU1GeooL0Tyc2dPKhu/Si
77MaUFwY+jqLyGWLHTG92sndDdoczi30XuFPDAlhk8mcQmUyu29n4xli8yMPd3X1X4XwD2wRQSGP
1pbT4K1VMYRi14iyJksMXLPTdp3JgVaoqnzFx/r0Bq18a8uVa+3FzpGG5SKgOcYGSjvGQx6tz+B6
SrqSerwO3bV1nGbHZbavhhBgBq/dbq8Jp1Ht4IsJubJXvFmbCfeDdnXqPz5ZYSymfc2hADYjthyM
e6l9OwE89rGIDdWm0OoyQROOkNtx1yI9Wbp/5MHcjE9r31Lkb1pyfVN0Vv7HTcp3ProMHV84S7EU
sgnCsK0E6pa+847/RXD2lqXufRMRxVieNY9s9TonAeAnDURxhhjh/GjgzIPy0mgRK/UEC1e9/6yG
p6fLVp+J8WhSNU6DZabvCJEO3z+n+VZoCUX6wRlWCRdTNhvQpzrTZ4qP98MY9QPPak72lHgyF5ll
AGCCU373AswNXYB/iS1Zmd2QjR1AQKD1w7MT+JycHYNNyfcOZLHYRh+2qAhMSv1KYt00RgCAstMS
P6E204Ml318Y+t6EcbwmvDVi1eXhxhpswP2DKPRtFTUo5hxx17VTn9Vr01M65qHQ/vmA3oeKvM+O
eh3EM+eejlwYKTb02uGI6B4ZCJWt7jc7gFoZtDBBFB+hIW4uT/doBtRLBZGKh4uc3j7ja2c7br2B
tMqA9+RDLWtCGKyVpo6ms749zG2jS8iIriuBdMfa9zcWtiDJWfPKkhIYsMleWqtrPvPB74aJ6QGk
H/ulbMRchY70gNV5q3iG+Xe8/f6GMjjKnQzTdxFyYZzcx3HwqmMSSC+T77lT4zvJNX3uI8VabKVf
2wGXtvZTRMquYiKyU0IrUHjksy4gyl/Hkpq4HYxDmuIEdW/hCq+TCV4hFzL32QO946+bSWv8GVfa
qEs5uPSmkwVOW4VNy7I9jxCcbJ7i4CgpYcX3Y7n7w3b5i+YfArwNIbzR2RbYlj8PGTkkIhGu2ykv
CXHcpMjiQET3E65708mvFOYqeg/Ol75fAmVspJ7tppm+0s/8aQJge+uYJPgtIKd+o1u1KjA+GWO9
xgtmz5b/J0WRAy/ZRNa4K7G8eQ+4Zfx1nA0kjgR2X7uSf0CpczYoD2ic4TsafBD9tBuQPQEus4iz
97kHyFr751ixJQxpDnQxk4YlHaiBKaKpk7hlopImynzcWGL/oexj6Tm4ZVO7YL/rqJYGOj+xovEC
gOCcJx/kuTF5EzGt09LGv0Xbdzb6Imnbe9VblAJi0923HPcMQpVQV4xosGpipMYwa2l9UqWya9TY
202+A9Tl5+ez+Ymw7ay5tlgsXsgHpoTecNWgizKg3bEEXyPSbg7U5umUmJ1KxZGOVgQftE5aEqXG
ClqFpby/g66lb6V/oQffWu1/n+Zq8FSRm4qSP583rXRrn8Wr1eL3pUOn1uxrpk+Ad7WHNNX+U2Hw
C9eGcKzmD72nN93/HuehZP/VdoWWBNvPisOACt+MyP6STPYut/sK2Z2sQqleXYQGeacBOOlOl+zl
dM9Uk8WrWk8z6NcWH8uCF9o4gjdyZnoBI+7IfNzyJI2Nx2DiI+Qc4RC0pxMGmVtuEiojWAj4T+iH
u1GpnytANQLVDEmDj0VE0txYKMFx+R7pHKBK5V0uq5q2u5SmFibCFgo5CgHZknMDjhEpVpldcOoK
5kUAIdBDL/Q6QYQtvU6I6tDwUWymHv6fd3BQlRjzNjuW6mF4MjnYLRPfKnlvIY2LL9TOMsfvf29J
npj0L7F6NsRxBG2GGIT9K1JfFXbQMQxUIKml1R/hR8V82E1eO67L0LUZCMDmmkjua6utXrSFr/pw
6houX5veog1J3wf1bBnz8l/ppl2OLsHT01CHD6PhH9/VVrQI+gVXs6VbL0BX730kTs1pzdR4w4+2
9apENmOQtX6CXlSytTrEUY8tuK6R0nvcuXay7TyC42gDCXp7FJaY1c8egK/heJJQBSigUmRZ5Mka
MCpCcoykOYgXKNOH3PqrYS2y4+vGRHwZ3UEtl2mlYsVYEpczMV3lDXx5NoGQBGQXMoirJOHFbQXX
rUy5EgSlyIu7ZPjtkqwApI897nhv6FfTL2UvGih8RY1oBF+0k5zAae8v1qQbXzbyyasKYAlRU1on
N/0YaxqwyBobdh93LsZs/2HVD2PkE5QI1JuIZtQNuWDUXi8CzN4VuN7X0T+UcmkKDy5g0fjFhJ7w
wc/bVn/zZWHNW/DF3+s2F6rPwJfx/wsWqSsQkQGb3ScXhRQ+ESkVy33xgDkAjDAg3uAiGnPa7RLZ
p549+cEcLywv/ZWRIbDc4yYYAUK6rMyrjcZZETyDU/xVh+2dRprTMnbRuIWnxOpxtrRc0ZmI9ZTL
PeGN6s3oyvHerny8JetgPceofsKBnZ/jsHTulCVphZTgemzqAYaNu1H9Nsy8cnDS/1RjAoYO2waS
ka3HiyY3QVlu9YEgop+BJMOWYRmYUDWp2gq6JYVxkkDkJ7CoUbVxxPBTFTH/FkiJn5/KTlGGi7wU
9433Z1tVKURfiN0nMdFv+6mjky0ayekyTRZhk9pUDXUhM3QJmIblgl83Grj3wO4Mxac80ILQXHgr
wB4TL6h4mkvAzyxWw8os+VWgP04ad4XmgDuAU2zB7Gz4tygpUVTXLgp/yVWwmvqIsrsnrXpdsJ1/
/1eBar9uzmrTe9kQ0YR9qUzqM6rZZNumkCd4wqQAEyK2XLp8I6pc5kolz42z2inSDc8T9MK+lku3
//PO/MjMNwKmUkzUHmS/c291CYLeWpFNzGO0id2pdbRX8Ppn7J3zmA83VpbpddctjhRE4QIkUXG0
HqKo/aX2aZ7Rasr5dboAsMyzR3HnpYJLoPYg1E2AKL09m1CjGibIaYUiSNiabtUuuN2923bIJ5X0
0YHA3CCxVWszTI5uFFNVUwCUuXrc0HG4+IqxkT6p7IH4QQRVf6205wJy9ZRPOnu0Or7QmYuXfC4y
LVOzUCWZSMsvx8oXmrQ+QRBp185YnTCezUHatpJpxnkM48UwdPcUlByto5h8RYlKGKiK8XCT4wJk
dBCnbFfrW1aANa3q/zzJbKoFQJvYXj9rZzqO1ZBsElFbvwZPLhtVOa0T19xfEvlrZCixHUI4eyA1
PEroDT/blzAqz39DONgms9SdQ3yR11UruxANNvH2+zzRUqBuhUYYbJu52u8Tr7OvSv5dMp0q/2TE
dCsnJu2CvAVNAIliUlmKUpOKEBKjD3DguGZXHFqucdya1wPeuH4JAi5g3SEsKEJAdqAoLqQLvUkd
IFYj5Qmr98dtp3nO1v38LAfovky9mZ4RhnU0JLisaf45uUcMrMHuO1bmIermtAelkzH8g4rFE62O
JxWcQSySOZ1uKrRMwn+5hmxnPzfxHfXmMsKz7NzJK/UKulZQYsKe6ctOZG7QnsPAt3+xcRPGr5A/
LIrd7U2B4S2klBW/NHqMRa3rVuM3yQxyzdLpkb2J3eGLmk3jYPFiM2Be1mun4DWu+O7ozESN4YLN
nxyGmXbY2zjD44B4tN/Nz8ARkYJ56O8IMgAwbFZV6ocEaNwSKURJERhbwExv8hjssKpbZnxFLVhC
lYVyahA1vyf2W++31r6kAkw9WPTxDyQWH0wVfPXSAJ+8A1xVdmpghbScMCJHCF9YHq4ewA8ry/mS
4abcZAA+tVB3ajQWMyJbQHPKL3i2dnWKkNfMeTnImqzw021fH/AYYLz0HrCkyhLSRgIySspiL6XE
LMDD8jcL4Tlo7RzowtK18x6dBGInfD5tGASZRtdp3gMEaB0GwOQS5Y+i4Vh8i5Ds95QEuEOnHtXb
HzhZUfP1R2LcRcGk6P7xOVs0ni8Y5Rfyrj+flpcZBF03Op5nkHRy4zCjfUcqG69xiAdQ0zWUn+KQ
fmZUCC6a1/h8x5eJGhk2Lc2A7lQb1/ZqilHEmgT6sihfjIHGX/qFVfhQYM2kb1A+/QLKISPgg5on
3EtfWz/H5zX3bQ2aXYu47aylCayQYNgNbgqtyyvg8QTtLB25PPsjNUJNfMbNRPuPGC4y8l+z67tu
jHfLSznqRG7tkDrfByKWbasYDQ+rafefJJqSrusevwzfac4GBnmZe1v26IID+LPQyBlf5vvqmPFG
fqgR3AvQdzVldcDo9tKR0y7CasqZctgwUasiUHOM549C3gvxYsyzooGYWDga1DgJQpEgkYmvpyR6
jro0Uo4fJ25nlPjHCj//x1bdRmv9A+hOj3gKZdz9iPfGRX5QNB8RBgNrnXjaKs+Lm5+kIL4m8QRI
PBlsnQre3k4at/2WGb9deblrjWkr5uFIF6psNsczm5Hub1JxDCeRa9qs9Pwh+Y5pihAh50oKcEnR
BwvNHmCC5xLeZ3K91Ac1q0IL64Gheq3hO7QhmoF6WWAzHec/l+4U6kyx1OFIWoQJQcyoRp0utkG3
DPP3uod9rhblExm2iiagKzevEO8FSZd4Fu2YYExtU9cz/YcCNJOUi35+u4OrEZgScswixyk8L2uV
AOBlFqp3zfr5ubHimHJ9MDHGtcKkMyOgV1dZOvdx27JfiWvbhKa7b9t+NI3UjDW0cTGa6o2oC6kA
gZnkn+WcBz0aH0lrcGf0qPS9vSe0hEc8VFuqwohs+fNl/loLMnP4Qiu4+97V1b2A8WDL1YvTmnAk
5At8zRKi8eTEd62yzbTdGjVqgwpYJk66VdYK9aU+8jx33PvoroJvEWNxejxH5Ya4bkXxN4ePaHjq
/FuOrYPx826MDHlMuXbysqLSZ6EI5zUYCcbNY2n28hS5wgUjsvf76hchOGJoEHI4VAof2XZWLD4a
aOeKtBjDhtAEsnnkJ0w7TdLyPszpZfyqPOpjWYAGOPjx9SGR51iPaAX4LO10AWVb86NpCv2+P3Hx
0n4FhY1qf/3H0vhyBU8YY86ZVyLn2373UTidbqwOYZfqr0zfvQgYhWvews6SFQ2Zcf++Q+Ad4aJT
Ms4Rl/wWgkysCj6gPPNzbUwjD+OEhYHUVetnWckN3eVkCKe3VG76ziSOYY/jNTzmnza/cp4AdoOE
F6SUOIYqR0EtxBU3ASIAuBop7lBxLpt/SZswEYTEki2gSRZHNerrygQkRLmddIoGuvVpDC2Z8zEI
LDw8saR0Biwc1WDi5sv0K95SAPpBUfwzuL7F6qXNol/PyhDFNH0KO06MDrInaIXRAjFdTT97EBbl
OXGqrM2IwTRu0YYg7qS1s20syknRmJvboc7DlC1+MDlnd7nfFNDcyyqqYo+hrin8qi9P7XgAXowc
Z21TmjPfJXGVUgEWbf74Ub9ydfCBfFZ4DbDKxkpyMJGSEHcm+52QX24r3e8ET25lv8uhsMwTD4zg
RnVu06ndM72JqAU70xsZaHt8njOdxy6w8YhP/KqNZ3x7gzj577eEFdI5txu/zBCXfueMg6EqBV4g
pP84BStIqPVYc+1UtZjxdTTsvOcwJstuBMV0Ol7I0IqQ/khuuyWYx4C9ufaZ2Mhlkvyl2U1VuT5X
wpumhvc5u1wmWD94IImNSf9umzpeDy50vSDiecl7u8ZJ2kBMjqyUMJyuJMe98cLqdZR7oAtv/P76
Qx+ZrikNgohJzl9S7pnyZzl6tD7QfZVykoG0R50qKbVCcxXc9n2WL4JdcEfAsfNU6hG1xgwN74rH
+fYnxC24LdowI3h4SUurcPPqbdQZZXbrgMP9YS98minx61MwCzA7e7vkf3OgfaiHm4qe/c4wcxiv
FE/u8Z2mgkF74gkw6GPLLtqYXIjGyLes9I+c0WWdg9rUX7bof71vG2AjHNiEmQvD1SMXeNdpvFAh
DI7Ai4q7e2f1d0PxzW1cYORpoDsLojGPeoS3QmSm3SLK1z5A5QZtUggz7OaUYuhfmICfk/3eMraD
Jw5FBTrkSJMCHeo6g5HOfjjWPRGHf2j8XHip9Aw9xDWGQIHmedNfnkf44f5Scph9c7kZ3094Ee5V
3gXLu54tyI99qwVcmZRvynICsB/5Yh3jRZEba6x6fLToUIOTTCMF4k7Es6emuEEJgiO3aeUNX+Zn
vt7PXKKOmlirU64B/mfIOC0ZzjrwuTfDNuruX0CsrUlCxyha6gZaWwq66Jvnw8h7cwyvYlOZjELJ
HSii5imra82/I/0Rv1MpwCNCTDJNHH3iHDZfzCpRHWd0mOq+yAAiXqvBAo3phwhXmJBDmIYF6UJW
02OpOi1Q2IrPMxXStP6jngr2C3DTdLmsf7huLfwDCdFVfbn0+oZZuTycmUkc5dz7RRH27r4TSqNX
4aHLuwPXDrnrdc+vbCLoDSPZe+X1G3/XXl+Em9zlNaV5gCZkbBo/4DIIRwDf8qaBoBK8nBeQe0Px
6Mopx4FGoyniN64dMbi4gsWKYWrwzJ2i6XbELez5+cP5HJzLFnl+XUbh9aOHTu8wY+G5Siy4aGWf
clI0uHhkxZ9CzLRvckfxWdIRceBVrBpJEV5XrZiY/OhLaLe8rgBiN3qRTrOJaCRnNZt1SyYaV2cm
/8uNjh+vLuHxaQxwdXiVegJ9rh4Z1ytzvMcDGrA5bTZ0a11K09ZrIz8OhkD/vrRQFn8lNZ8oKzfC
nkpM8uF2dCK7oLnw+Ivt3qDWP/rKjFhx6PciKnZJwFREESnXyCA6/sYTJ42/f68EhHfZIKOCiK1S
Pu65Kq+EsKI2FiG2PadEKMKl0AlgP2qrZJ9GACrW+Kfmct5Mp8PrMsXczmuH+ckbp33iqsZ0TcwD
Cd2G0SMSgRLSKXNYRAr2feXxvCep1WtjiY1OR9V3cmj/H0eCPe/TeofqLPjLB2IGpXA2GPvR087+
SDgyuGyaZx4gQf0q65LH6Mi/TdKB6+XDWQq9LnyPsnJLthx2IFiFu8n5TdFtBsi0/PHqynf/0D6N
4txl102Q1HD8ic07GFt63Q/KbBZwRs8ACI7biRjgCC/20o+ESd762EmCL3f6rTjDx/wL2a0rl7ET
/O8xSe6098ErHZad1Uj7iYp0TyB3Xa89Jo6WaavW0Cz/o/yde1arfQFe8meId9rFb7ANazCowVWY
+pOUJVDCBb+Moxgu8YbFKpq5Wfx6hBA9onSPnvEs9+l+8Ju/OxmPGt5eotZ52Y2NHK2ourbTTYTG
/x4QdJSBo1ccePgF2m14Y+m99ML0hOTSJMp7A0EmnZVwhL4ZxzjwtCJIkpLPi/G8HGV9diJ1jCTF
C2aZVKVcbj8YNOu1a3SMdEdT5VrlsrliD8gg+kLYJ38/AuoFG7jKOuAB8XRjIpbIT8WEPRcahnWs
AzVh3JlMQYcweVPO9DAjiun+6FrNtua7Dz3YGVMxykrp5nIC1TUmhqW4cOg+Q9XeFVrbOyXjb8xz
sbh84PYv2/cCqDPB/f3sKV1WOEKGg6CMYqGB6hIKf4up0Eq8lKi7EjaQRvVY/OxfDiUTuDvf1eD1
tJFr55vVAt3T9tgeoB6Rdx0k5YuoceaVdzzrkT9lyDA1u1s6TSXvh4mT0YWoLZAk6yX/q0BJGnq3
sSc0hSVGQlx+AeoWoXdH82HQn9uWkrVKCF/V3CDMxaOLz6TdSP1otk6mme/C6cpvFG8K/EQhGgF6
4dnzLRzlK56cMZ09tdwi9H3M/QdeqFsBJ8bjrIBLNIZA9ISgd7Rpm/ROeiClpq79tS/1FhxAUVoU
gW9OJditjQE2bcyb0FW+cpXYacmDaBNFHmVndbfQMDnuOM9N3GMnfD433frrcD9Ct5a9j786cXC0
OnIyp36e9zrhjO4sCQ5hEw8e1m2NXZFUCMg9cQw8BDkw06nOxl/bzwRmMEdlcD/SRwFbWLIzN6uw
XVqbxAbIuHGRifmqUwkatsyDqIg/+RgTqIw2ZZyQIXxqSIuWDHaKnCQMGwjrOM5f1xGZsG7aEncW
xT9kpjE33fWquC11Wt0jilPoEvwC8S/ocIjd0b5b7E2bwQWQcFqdPg5aJvhtvBCRD89OvWKWDnZH
3s1RkryQo66ELt9KYNYOINFovZifA2qwAE/ELdwfqb27Laeuq1c0x8bK5g/D7IcXMTdxJhmMNRw9
RN90fbj65RoOAt1+DBp1xIzr7vj9RS7PLCV13eAxik8iX8qtDkj1ClqbJuTW+6oiyQlTsNcIMWDe
zfPHJsZ/ANO5h7PuChZtkHn84y1u1lm97FTWYv7HzbyBHxy6FgAq67dZLYIcgk5F5G/4fA+DOukM
VjbEh9ESXlZA3pewDdinSlm5FcG7c/ofCYubESLtYZ3VUsRvt5BoMeDBX8O1r+h/IErieHPaCoSl
8rgr7UwaTyfxt6Vd8Z5g2Rn0cI/V4TY20rx9Zf9n1qUczF1L4WFL3mHmjIsHtxvgvY4+05hSYErG
DQWEvSQ3qOPiiQg5DazL5dLDz503kk9hPb84vf3FQT5EkRD5iRCTWl6fl/bMg5PZqeZLBaZYN0Cr
sWGRTt426xZH9C5jXTSGmmrRlwK77xo42kW892Qw4uXO699Vrtvt7sEiH54HIa9iOYPMuBIsFR2f
aT5OdqIM7scqNGros/mE7tBLMtC5NsqJI0ZFs7WsGE4RNKCqf7DSeuDFmNlL6BoN5iV5WctYCtiB
zs5mwlynBeqCk+T7nAOSBWhwktYBfpCIVWX+dqpt0Bjv1TpqWr9D3AYr1W4FXpS40U1tgncxw4x7
0JprbFXU0cG+z+HBWSlFJKy6ANJA7Mxenwal8HOfV7uFvWUZArxYTEteckNqPJmMRqfKw5rId5/L
Dl0SsX0no63JcoZuYuhGzWpAefnZ4w41Lszzyb3Q8rQFI90nuDe36cNF5pw04gBSlvGLj1uxTpeH
4XbhnFuhTwW9/COYUt+qrKE5waenGnzbGJEee2aFQyzukrFw8NmHB/xW6OxEqgfRsxp4NnMNVsOU
QfCLZ276SiKs9xnFkh061MBcIv/QSV1ucYQaF2p1apiPgPh3avdqA9EUkw3MkdgN5SrLJDdpwntb
k7JXlLGeXchqAruz+RohcNdLcsQSsVELQcEP2EG6mBEm+JFgdNxFOGGU1wauMqwMTmvrC4xK7x9m
jHffbT2T6wEpAGte3G6QjNA8l9twdulhCwK6ZZzY0bTfe1R+lnKYdffv6OVYu6kJZxZaHjHBupum
y4ThMvwl53ummGRATWp8rOsCa/acvrkGpUD4kmNFgY1sDh0AmPWx8gX16xsOTtRsVhKQDsGjnynp
zawdsjmupu/m82pbCK3SG4MQaMYby0OZoPX+FL8fpGvVlfH4nCJyUc8xu0dSYRl16VOI8CoQAx26
hmpw8uIIIR0s2hdrDKw6HNYiA2wlLVPG803NGG9qTa4EK1wYXedFbTI0UO1t+lO6QiXFqWOT/57U
5Eld2P1jn8lZ2GlJ3iimje7x8fahiy5pckIl3S3FIyrn6Lv29QmPM7Zv4OwTu258stmN6TD2Acvt
YWx4NZt8+Y18syfMSIhUcOGaAMmi8i+V0Rc2cF4MCdwY4qVUy0DMNNxAy41QtoxtmMM/LUhgWOqf
7HlK3Woa4MboZ4Tuj4Y42iIThKMjlAdjoOAnXrdaDPSB/fwlJPaIdo/xUxsYsjeLMTiOw1tE3ESL
/rgshXqrPNGFgLPSmXZrI6Lj6hSMIBICuVYLNLSeuC3z/H/12HgB4gbull0OLfnG5SgOehBC6lSx
HIiKDmXi3pg4P/v4lsmR8wY4xWVOFNSIeIaPbt9rPlYDsro8ehii4TVQx4GM1+VXVrXyRvYg4fby
2BYf67ERfUOzlo4XnBeWCMLboLOw+/8zH/mNPtZXUSAUjucWpU1gIUnVycUMiih1msVt7Y+dH1Qx
0gayqYqoOiaz1wufbawwRhfn8PgYIiyqgfAB9fWDT2yGBYcJ3vLKOMKbGXMEPa6xmBlYH8GPs+p8
FGruO81wRuHMHlv4WIgo6UF09yUHvtQPIwf/+nokzspqH8I8YJ8Qm833SnSAnQtmlqkP8kQbANpy
SCV2q7H+eMyFZeVxD5aXw8sXBSgYEjKVDW7ub6C4CJ1a6Ku4U6koHlTpKTCRebtZ/5Y9CO3AjJKT
mc8F3y/GETeBowdnNVv43QyjSXvH98OTz+utKF6+hxCb+jxY7BgaS3sjDgDwbUGd+oX+aX3Jl5Zi
XswPvK/y2NSX36cSUvRosPcGvSsJU9WnkDssp8QY2L6CqmyXLPZ+DHkuBsCFwNtpWXf111bpaFuX
EgeXA0RasqsKJ7/T3pFW9NfFN9tPTtmcUfBLpz5/MghWorX9/zsOZxmm7oyvMQup4bwyCglXzLv6
fd4kGnpmAcqT7B5MNuHctrtT9qZdA0+9sstaP/MjOGhDrAB3AtOS81oUtGCFmJmUA1u+rQnuVFJR
NKIhMrHqaOkv8YqTTglXCjVdTyFChRm+WN5xTp1zO0KAPI+Bds1TDVfkTixUZeTpJUQnoKtXZ1x5
jvlCfCuw8hu94tOFyUjOL3PWggwyi35iat5O+vfobzWmaPbrxWoGNRD3XcSEfBgEuspnFbyW+WyA
Pyr931aW2FllL6H+hB2Sso04IVUduFeJGPmH7QFfK7GZv7M55+kdKmg9y+o34TP7I+V+z+gz9rzD
K2zMx2SUcJBzd2y6bQma4W8CiK+ToKaLKUVV2N+sM/LECcWGt1beZN+q+Bxw7JPRq5whrX8rmK7l
RS3+pmHIXbbcpWQ5ehXQjTVDgUbYP+bgeVN7Im13QSfEgFWqMhjHChqJ/iNW9bmM7yFeNjx0ClBr
nGBvCQ0SZb/5u6hsz1BAkVOd7cPnxq+zmyHInZ0GF91qD3OBhNNR4bLMb1C5xSrMP1xV6cSAOdsX
uNijTkH4BV9j11145NfGa04aUYQI+1sZhwYNOhPnaxVwTr1ghu+zljHfaJSyDQbI/J8PcAT2wpKY
8etDH/l1J3ZIn3U2d2uHcsYosCYnPUm4UwncwOA7nYpbLbTAW+nV8i2vQrJpjqSBNvfc2fleJegm
Kz2vQ4aUF5RK6fx6iSAuf/rSReT9GSjCUUt45gjDiFCXvJH6yhPW4VcdR4EHDFfriauOwpU49SRI
wyIvWFbGMFPwBFzfU0XE2EmPzOTiWoiJna7jCOFF9YLAr0foK6S/6hxef/hD+Xn+dz/dSWGh7cK3
tXH/SlbkdGvpMtz0o3QjgCrhXrqq+dQENA44d0dTROfnV2TbSgo9tmFQkRDLcMaQhcrL0ooGXWWT
AMZKmD672SQ818H2qHdwBioZpfuDaJyOXv1gGNwqyjjmJjLm+tly1o0CMwkoAqkIAZTUi73iug1R
g4XeDrTvY7Tug5a53HQwjEccLdaJaFUlzzVJPyGDYIKnnbOdIFKzHRaC4YWuGW8L/cuNHkIgupYt
bnQ8YuskfbkWkhBHAlUkCLb2WqOGJzkWNWOluFszPh+/hvxO6NjAQR8poQ7/Lxgn1UZIiZWRrklb
dl3Mh80xxlpNGzG1Sx+aIliSBfYTDfFYR9rY5vwEnyII9Vbmas//I2/SEv6kaEDzJbgPovjDZOJ2
1IPdQAnB3+Y0g/3CLlEjws5MkPCuyTdlh1gGQzyAiOY8uq/fTl1rppEY6l2WVOYgGYjvbhL/l19r
8qeswEAP1o1S5Vms5VGrAmZI40ULC7qgy1WROEly8pUMaMYAoNFhdV1Hg0yXlzejZEj+hAxf9ZNM
K9ZOP3tQyJsjxor4wspFR7jw9R0oTFd6Xe0QrwuACgvo839CrPYIc0FiSZ44Vb0JJ6cN2dNG9Nv/
nTwPpV6zZhghEy4u0GxMGluw7pqUwMVyiDsDOVsmGg0sx7GnPTSnkMDCh3CWkMeynVrcyPgS6l7D
8sfpKEMalIkkfF4BCvWbTLwDmbvc0AqrN7zO9VHHzg1LAazRMM3zAiBGx35wQ+KAH++1SZxjwh01
rd/VafWBGgxcppg6NAmsyCZOamm02PndQUi8mxAHsNk+WIQXWoF7LSLDkHwThmRBdk9a4h/eXpEk
W/cu2PSx3FjwnATAnnbhJ/RGmBsHro9Dqwm6eK8teBA/8tWi2a8ijem/WFFDiz9ziOJ12zxvhLt4
oH6948cyqcR9K5HNGexf+RQ58vNAdlRALsJeAdQPoY3EREjtx3pzkcaZcDx2WoyxALXsljDou6h8
Ue0W8Cd8dZ0OeOasTJHzbdP6wA4KdNjxRmOdadX1tfamNaxHBbCsH4ZB2YsJVT2cuAJ1mk5KPP4h
NTHeaExqUOHLcGVPzYQJ5SoIyuWMN8H2iNqGLu9DSJvPgMOUGPmxSdCdH3mOpsEyiUAgEtt9Loyf
4zK3gJX1s31s0EaO+7rz86I021GlS588hFx8NX4d2osmuVN7K5miJKVf0DjE7laAYkYcrf7fNmtv
ltLcPS+LMXC3MVl+/cWAc5/OS7OpFvCjxnamQYN3b5zW/PVWBQ7+deM4XpW4mQgarF04mYn6C1QN
Sz8+rMIqcaYnkYmOeReLZBrb7ftizw2P/z9DTbG4pZn7w/3d/6o64UKGvoQJf/L+xBLEedkkdNHQ
axMs+c5ySnEfJsnzaAPVDJtTqov8cFCk/PtsbH1K5361kQMeNRTYNAahoAMCUyoMRMZ8rLmXCZ4F
2M0zBWEe5nnXv3K0ywjpOmgYhlxgnPx8Mk60Vv7UNHiiGScrqqFfv6JK8C4RkyLrcL+jmaV6mFz8
fyQ3QVt4NdxUMlTlJJCWOGrOkbrfbyhEFUzZP47F3ReLnwDH3oMte/KrQDUI4c2nlOY/frlDYals
iTTjJB4dYo6E2Po++jTGa6zvsXf7Cu0ubvtD7B0z1j8ZcszF5IBka+DGI84vBrpCLXqnwjdaH0V/
fHJ47aZAZCXA3ZP2dskbOS60STDBQPkqmkayeH3uVORhNYNoPhStoGwuEHzcg4NNhCi9/zUXdlTc
cCiTEPWAOoFFOnTbSSaK0YA/Yc443TDxm8WQ0njcKF+0IQNZ/Iv9+UEnxXOpwLfs3FQdaTJ4kYv1
+9vbQkElI4+C0rEP3GaTa7jJLmMpQmQb8cUfw0i+ngKoBkbbBXV2GmksAsEICYTBdPmJdRBq3HVV
tJE6ep4Ob+kW7AceMV0Pb/6GHsnVv74cTCXWXI2oHWmUoHFW82v+5H+yzWyxRq7ShlVJ+qKdSTBu
VMQNvVb+Q1S4onqoncqXi06v/WNe7LDHlqZy180R+rRXYx1DzR/PQwEA+Ebjym3G877zlVXsTaJ6
dEA+wM2vyeGA2SO7b8YVQ8pD6WMvCSivqchZcINAYu94y47KzUFFj/5SXD+LRTiHmz3UMtQU8q3S
OYP0qAzDeK+9qn7WL9A9ueAZYSfInT7LaDuB92N/tdYcwL/ENCWuPrqZc8KVC+gYxxqzNOTQgJUm
/qsx1Zs8lSAuk04b/vqXUgvlo3uY9MnWOoFQ8lzkluCmqrepQrT0T15Q9jp3rJYjL5aJX740NTNp
UhulnzwqtUdSWnMuUYqzXv/M2xgs/yk7T5n4k5uStDyMU/dqXVkGwlsT22zwVi/FyI3zeNdApD/6
B5/Z5fyNCHtI6mTqhaqwOEz+0K9kv6qZxOuvqDsr1V3eQaGJre5N5uE8FYdhOUkKoFt2E8oUicdJ
UJD0NWthKD23sMkwboO5qOcBojeY31hpKhc3LUXsDkjZcf4Fi04mBfYunEaK8jPsGgwb7ayhPRqO
iHEjGyqQcR+RXDICEzU1UGUen9GyZmuxiim7IH3WdLCw5UtnKEk8/wcVPwX8+7A88K2SCr5zFFK8
5jSzJvq61q5JqyA7wIGVNesWzxKo8OEd+O5lokANPhruv3euc8NLDAf+ciPEkFJiH5vlzTTkdb3n
p/O2pJ4GH1YNYXX87Sv7W4y6IZ5L5osms7GeQlogrwdG9US7HJhVEcuJZi1W0DHYi5KaU7UQc82+
eHd5ORerFpf/6ENsbtZZ+/9jATVpuMLKlF2H7jsnEM68oXqoYdgS3TkNu8bQWEBjAK/N6w1bHWfP
WxcUhZos804LpRYSq2f1awOEbDUXDqZWKSZeNHylDKv/V1o1CiaiySSbxjn4Sh/GRONvqEwWBWJ/
m0BrLuNWMqc/UgX6FYTDCHDuZGn/V9c4ot9gFg0huV+IHMScw8a+4gYIpzf1EAxSb2evCVRbg2K/
H3IwCdqVKA2qFf6/MAHyymrzfH4qNwBVBqi2BAmzpZl1mBzChxgAW8cxZhOainGsvKDYaeZ7EBdP
enQOQHwVu6+Brp5Us72d3lfiJ8zSn0XOKjt6B+nhC/iQrfcGxCRx78cTVCOZiOPsPWlArjd3gJWz
99zp+RHDGMhOxRuXlC58baYOOdg12GJfaNwnCi+EMPJHVV8hStwTsFt+mrbInZdAlTTxHJNKefZH
+/X20YHF9dVBTHiYKf6ulLQDUZLyuBL+Dq/TpavYQWqvYEYtwQnS/NBmQyG10K+Gk3MLsQkOlAI4
hL2fvhqntHuvY1eyhuY7s9ewFNimfkAnnLZ0XnWX/GgCPghOThlyl23HexsVdCMsq+6DB0IJbF+J
1fpBOqJcuynlnliDCH9JjnHhjMLi0Gyn17M3Mc8y4ftxTiH+Oy55wYdGcma22HVhfKLRN9/iIA7H
BkJ0KCiPRriQfCiakuAp15koQSDTOkH3b9DXzWf7XqcZSAq1Vt0X578PzqI3URtJDF91a2vj+kNw
aKzboXo125gOvNfIU/WPQreM3DMi5Jxeb6i46QVskEgFDaQadE7yhl+rfRATV9OoVlmdMci0uj+3
ALengcVzfvsJojEY+8v6RQFijoOG1ao+IBzGw15jQUCUbUoPMT0iRloI0wlVeWwq5fNSc0D3pJ0S
TbE1WN+UJ5EkLBoJb7CW1uMxmabgqPTBLHbEF/ljcnB6T/NIfsIuTVRna3lIa7ka+syPHrhbr++B
CFbGKWXZ+vcnuy3eieIgzj1xYu1qBWHkSL4aUlYr50otQM/mQQvBjsCrzakKzEwvjw0Egs5ke/8K
fN1jICj1bdYV80MBiRY6Url+jirWNjNDFM8U8HWQdasauoSZWR5Ozxkk7pzX5cbEHs/OBLQaecoF
KNV5F4k+j2yBfPoWqqNKGBUNPgJMqWP9QGuyBByDKDy9YSgrs2bW9BPwSmqASY25LRLoPfa4LB+n
OXM+hZaW9Z2UB95r3vOOXr7jDQDyXhsjrSHBAdVemrVx/WmdpibZMw3tYiz07hm48Cp1URYURB3N
F3DK8I8wKeqOaVTdHSj0KI0JsUXgO7USDylKa9UaDLKjR0Z+X+j1cPBk1CU8xB0ezNE9AIUoD02/
eHu5IUjBQAq1rW3J5l094/QHbTgBfYjJnVjyaN1cuQpNlTWkW87CemvA+8j69NuZoaI1bgUbLv7E
ApMgUwsSzrxZt02OOUUUBszBLIWV9J3FonQlJM51CHC8GgDtxHt5UYHs9l17k5ZmC/xorWUg4s1h
nh3hH146toTkYS3dxPaL/QXcy1JHcKU5MlYPDsRkoBrkUunksAhV/2bdBUHAwTbC1syYyU/go0Or
wk1RNWIaf9uimr7g/pbZrTOz3J1SiyOQ1DNWgarwZwNp8R0YupiPZ8EQjemMZ0I1Dme7Izm7yiAm
KHD1KLdpgUnNhPjjMq9cUsMKC4x3HiWpFjYVcihO+bNHjdq+5xldMy1BwQBGsW9Htm2oJijNS4zi
C5dz5JBo85/GXSIg56sqC1FIi3LJq+GV1bwH/wbx9sqOapKdWgDtSpcNyI/cy0end6SJq/9tDh7P
K5s9Ki+20HhBKcpB+4Rl7OQD3Yc//+uEyk8hA/t6G0JMkB8FUacuJ9qJ8b7sX5PTmj8lBsHUH8Ya
8oZ7U+bb7sr19zA8XtsWNYfsHc9hsMpvtGci2CLMV+FjKsRvNDQGsMK6e6RAg5kc/mHjiTYluZTZ
bhg4oY0TUGI0OJSmXsIWthSsNnVTiqZi6TLjiFPH/ncNj5w5mbUK4WqDhyqVtEc8pPYSfHIX225o
FISkM6TrCFa9xNzqT5zTdbEukp0dhkwZQKyckeyB47LbTbN19RkZyR7ZXkiA+zUq0TMQxA46Tkj+
5+P/wZcfpAwrcjHcYUnJXn/EMubhokkKapfCZKLqAQSmnTLqEXtKAwuYYEie3y7q/LPkvzBX64zE
7/mIfB6Xk7And48Of1B522FEF6hLbGxpo6xqU2Dl/nFRh+BHatcBdXLXMxvxDwNe/VSABtzniAKa
z883RvCvks/l/azJtcMikJqFLnbZ5a9otkNYZR3VRE8TPVpRZat0MD9FyP0BLiD4giFlOptKNpoY
yBYCiILiS4vRLBL5A/9vE/bjAiCz/q30L9+dFOnTH/SerXWwbiuzzXgYgwBh9vXJVnF/tx1Ohdh5
sBB5bm66Z//0FOazIInqsjjPbOey/FCNwWbNJFOlNb7Kn98nNvqpUYx/OgqhGCzPuhwoksqjXzaX
CRX7xeI3YcOmQMJuXJqYmN0tS/ianKV8yhiQ1VJh+CTwtuNHeUSdBUWUmKSPRLHGpSn2wtVOTePN
4jd18n+qwZQ2GZUAcYVHS6MHlFuhdRaQa6/07w/J7WqW4nR7gdo5hVFwEaOCRzLmQgg7wGhNoGpF
Wz0d54uepezYgJDeZ6VdLo4Ks8a/+lTSQS5ZtlbxQSHv0tOzxF2Q18aeecsrXd5U8ITxMyurg1So
ZNR58P/8mD07TRZlVz6YSuVzdR3DNmCX8a2R1EQ0WMh+LiIN06y91nNEqTyYJzWUewpgATJqmqR/
yyTkDWdtrWq52mcBGim70ALLC/HFpMgZ6Ki+CHX4Ih10G8hs3/Up/h2DhKw04vtwjUFVEZ2VS0cI
eIU/6XChbeaqG6qnvFyySm36SMwPkUBhxM5zap6vHGA6ObTlcaCQZ0dWIlnjyMOTrBM7Ihcno+ef
VaT0FZUbNU7MKkKUZEKBE6jykmZpQtWRX5hgypxmrJkaRE11urdodcUsvw7yqb14UJSBZ9wht5mN
+K7jfOL2Wc9lJgXSG5gguBznNWRGMWHFQ6obOzFG4NFr1M0i1ucFTujkOkok9zYeGaxFWrjv+UHy
PZrbohjtIppv8AL4toi6fQNlVcmx0LjBbYKW9KYItCAuY5N5pQlm9VLxdsZdS1as/+t1FLCzJUdC
OopQ1r8J7h4O33Tr2UrMpgiOluGrzlBltDIrLVbFG0sD0wfIXIbXHChWYrkS3fnJ89vWikYf84M1
4QdP8+2YBLgWru+aDbWbmkI3VZWxThwv9IvU+HhLuGNi6Q449FPne9zXbqOWCigBxX7hZAtRQQtj
HVy3hRS5jjhCBfmcs4lPIOuI/scn+KP5/fssRTk/sa4HmYtQE22EKx+Ej7DykqTGE9WeDrlj2tCV
uxC10LNKCyQpVLgni+LLgpF/SJ2JX8ygY/Nv6VZX8tdiDhPwH8IRTSKevQM6owuLFoFLhcj8CiFp
Coc6wdbBRlu/0nrIXCuZOD2uWkbcQsE8nRSSfkyT9YYtFdh8W6R5tqJUopiBA4AHb7BMmxdedyCE
4RpfyOmSlGURO/F/DIpn4xJ2SlT8oOcuj+etNC4zN0ydLRDDVliqy8JhGblWy+iATtkK0kEC6TJy
qDeXT82IyzcPAvtTsmbmwp/q5Cqdg8aMyiaRZ4+cjwH+pKmviQT822T2DONDTvhScZGkDdUHjHQI
O7q+LD1zEktuTjv4BGM2v2Wj3EnJxiqyr7YO2sJM23byh+JB62nnVv89gyg35+4xnUPB/J1uHFLH
w604dn0RL4Y5dLfy3guicYknZhB+rQg8vHOxO/jbrzM/YHDURnUa43/Q9/Mctwn8gef2X76lxmsQ
d/qrrVIkeVINXoWxrevk5Zz3AImEgMrd0U2vUGMEOSLvV6bfVkYIGCYMkb7O2/g31MQO4fY2TtM5
7DZQj86UvNfFyAAnmjEpRWzRjqoRP4+ThiiZ8HUt87EBLFAxV6cOfrM3FTSjQvUhwNMhh+s3bAXs
QkiMSwQsNFZHWkiUiszsFCjS5OCCDDRJlwpLl/8mXBCvHtu0uq0XDDuRX/UayiJSs4xgZG3HNDxe
KGBlB++VMpUjH2Wg8baEqjUXhV5Pe40sSrSeN2az8wXqpv5ERRReuO+9QnuznmDAXOjdb/uOdYk4
hFPDeMUUeohvuR3Yuzw62B5JfpGI4KuNKYPhnZNeranQBHAFjx9YXWEG57nJwteLxiKst6GunVXk
49YMb91M3hKxYXGh/LsaMx96bersAqZhhwaJnSfx1R2NKkCooVzBFXzv7Czirka3WgmZO8SWmqfF
FBFHtwFB71Q7xZqPENR2oqWKw4nnk06xxbuIPKvp/rsFFpxsfpm38D3A6oikFmkmz50z81omS/er
r0KdWd+p8VOakjv1Qrx2Rj8dd8m0LYz+KN4B3iz5AD31bEu85Jc5mgmOjgAg754J3krsqSvBhmU/
D9uiMAXvNJu5PuGf3ICPqSVTvMq33Gx5ZQ5tMhZt9kRRf6UGP30zOzwBsHl1A9gKphzPm3Iadv/8
u9NpMR/5wpuwMTDvsTh/GWbMoUKu25i2arks4ykyjB6fFLQOPAitpqPuaCHdtOAGn0Rg7UeX6U0q
SZiyFqJkKr50Sn4XE6npK1gAjamaVg+VcvQQEMtaRe07WtF87+AVRYRyxLIChob19fUxC0TpHqBL
8tfm9nTfq+KO1N66uZYXdXIM7vIlB7uyJyx7xqL4/qluxFdx8XJZ4np1eysRneffEnmAU+7Ha61K
l22KftW9Gs6x7YLGKSGboH3CGG0nf/pn5k1/6S1lZHLVNc+K0bbZwQSS63jKdnz3m/USpf63EOYG
Q89YW7iyrFKRBd0gBWvYGJZCAJL6QcN1NuSgSyXkKGtZUdoZ80dIMaEGGuxQKThcCkAesa8toaae
a4hu6VKytb6KQcKr+VfJeqLxURm5ggFmriFAaPsDBf+VtV2yFIJVKPN5fojqPOGYt00v87kVDJCu
hODs3WBPR+e77yHD97+flM97s5h2+pkMPkbaB8Hp+fw00NcSiVRQzoPNZuiQZZjh85kwFzAMn856
QRp4SXwe9CKXIhOBFosG3VaDBQt++i3kwx6OJXma4u6hWqpsBZW2FHC06++GBphFGHZqa36+A6k7
eVZx6Pb6acbrQjdqYMtelrStcmOi7TIF7onFjrhS6KQcgCH9DwJkL7zB1TJA6xjQbnaxazunBkdq
4YWYlV5UDNKA608QXAnr87ioSNyPA5M4uFjbtcrNK8U1nE1FUftZdGcNLAFcxdGyPuRV9XD6kXdf
vbE0ALmQv9ejflemKX16zjKTOISeRZo6/Ct/N+x0ar6dEpSgFwbn3Z6vAGzNEwEiUMMKVQZ+Aj/Q
wpqWwGFhiJF2UCsnHW8ZipZi31w0BzzYWKeKmyGohSroWeGIz5ABOkFj2QkIDR0OwkzN2wXqy/op
W4JsyThZ4DyPG444aLW7+LtMddLvCtZFXjsc8TQiNiYiZ8tYY8tpBJ93GpvjLng6B5wDSkFYv4Oi
61k/W4b3Cc6asWU41Mg30dvB41s0FSJf3jnwHa0/d8B7PXEQYfQ4dv9AwpGfmTopesDy7N9rwmxA
Cp0uKLOU72E2Cu728mWxQXEkDTBnzONVpdg6hTX9TBL98nnwHeTFihCq2omJdNSX6FMblP6PzQwq
sduLsXp+O1oWTHXOAx+tu0EaFSvNmMfOX4/AbjOqVL+s6IeKXh9OAMDgJ/5iesfdnS0x3GGR7a/O
EPd3rbnOSfIbdghQlczGPd6oejvBQ3cX8Qp5ng820TOsaEVmgwhwFBusSYmDi6KgxmtwgeF9HG1R
zxiZK0qC2/AP9bWb8+SWIYnaAt5+f+xHQnoZJzhcfC12Wct2V6e0cY0VQlI/6JZlKYeUUjGpoO0c
vQk1o4MaoG6dDzbbtBhgm0iZAIbqmTVyi9/I/YbxtRforeA4EKvamn74X7Ed3VyMDGZIh9XqmTWK
AqRajkq3YfEJh/4pwzcBlBFK0jmK560jSb1d9e40RJYKIPtfqVjdWjeHdKzbZsg9v6jzZdQ2SJK7
9oj3TtuFOspbKZBRZU9cJdj6y7XtlsaMMpSHQ6XcfvtH6N048TVwHLB4ox4Q1FhnvVgujPp48d06
iol2Q3ApT1QqqRbKVcMnYPXuJUq+lRsAiUh2T/i8TZyhvDLT9nZi5gLe2mazO9J8xdtLYAQHFfFn
OqT2v5PtjUbGSmLbqCygV1bVvY9tDTw3PpDuuW+Fv0q0ynC2UDju72DTUX4zPVz9kcDymfQh22qi
m/sByybQH7C9JRtefa5NUD/v0QKNA/+MvMcDSvy7xYmUKD7SbD9legcnM6+mV8bqkFpTSCxF9BYB
si8cnhNyQn1KZYo9aqwB+lzh+NX4eDmqFaDbTITP876zi9WFAGsyYIMJeT48udqwTxdN/794q3io
c/PawlFYU1F3WmKrAGDdaKpOCKg6n15cxIiN/2Tjvc91kzbeMfdw9bYarP/U8/JwKN4fssl/2kvD
vHf7str/kgrMG2g+crte9/oBQkyNyfMIinIuZBz4/K3mxTNbYL96HwbamWsQ35t6T0+0SuJ6br7J
MG0IKS/fEtlcsedo1B026hO0ccZAiWuMGzpqF7hyKqy45OT6XRBAqQsp4yVdwTHfR5TJX4St0d4B
q/zMLRNZxSQ+sHbZNVVHMoZxEroCMPI6IwMyaVXCaM/P45JY+6WaSeYmsxR3tgTmVD6U5sUBqYkZ
O9H1w9gRtKwrIhgP0M2FHMAuzDfralSFO68oBGdr+q0HredHv7HR5yb0tAwxKM916Q142KzTV+2/
jk3Xfv+aBNC+Ja/YmOFUGKQZ26a+pR4TVafZYIRGDCq5hOZluNnjw5I0LuspE+zJTbHPPhJvCiZF
dXplrEiAJflLGdLejiKPg97FMzEu+JiLB0D9DoqynRiBwmRa38ucaAyUNrp0TJUrqUMvdly2t2Z5
8OdtEsOn/2vPBtIqS/Mr5zD+4RfQle4vZb4GWPbO7lEDrA/1lGStFvtkAWWaWRyLjyMKmkl8rV5F
E0/3CzRG6rPiHJSujXPDH7gDiFXno2C2FlAx8U9hYKFDZ1TA4wx8/sx5JHq6O0UcMdJ+WjGnt9TY
ecllNvqKQzKJgOIUaiMYxUiZT/+bVbejmnfklzhd2ccHgGZoJ4NXirs8PVcXKAHrwS6+j2ubcvfA
Jl+LOf14lFZoduMEvdVzXH74vBYp624gQNIYc5yoMapLK5Xj2H++cB5T5Kvd50HQudp3iGE+OSLx
lqP8cthDTxPG1vNaMmaLPZ9MkqGBONBM3VqJh7kAEmwMh+hLKNpseafdVF/ffVwkvGyDsVw87jzq
Ffwg1gODt1kXp5BHjHSWZ9FuLQi2QBm/n3e/7gG//QN70mvLOPm9opQKkHWu4u5TaTplNo7R/frQ
GBWt0MTzRQTFvvmfmrmYfBVv3qWm0MGZF+1HTlgJLqwxAy+nRWB7FMHYsNY7mfLC2Gcv4vCH6D+7
IujZAjDDxoli+pnmBZ+EolboplbdbXwRVxbJMr4PHYbm6ZP/+K9c3yrqFwp3JiNmiVg7aQeYN2gU
wF5W8/UCW1qsvodiu0ZxY7xDf8dK4C03OVXkzKvp9hLRmL4rUPHR5biyxsaKewRQbZc1opyfntvf
gR7KU9hkAXnPgDYF8OuG08Vg5GamXGcYOaT4rarJ+5azxk8mSIemLhgfiUYiWnzKgKLET0cSB7aX
VQqO7ifTRiF7zmdnI1tX+tF26AlkscRi5GA+o7nbteuzjnH8LbCWbDh+3LA/9zv6P4bYMnDbcU5P
g+nPdrXZ3fD/WoRiyLa0meohijxULO+oBzvMviWPJSH7wjtBQJSlcYWk82mzJomoW+IpeXft0D+x
765YLHOkaA1xfv+VvPpGJf5M95OJcT+28Eb/QOeVnoZ25KYDNBTXwFNaGU3EGlGzpxjpIvPyxLuT
x3ONn2tgSCq5IdX7D7jnFW6Uh+7kGH9DSEoy203ypt7eqy8OP6Nnz40m/uWg3Gh7Qjo5u8yHlYzs
aERNr/mhTA8B4wgPoPo26Z3eRbS/j8xDs1cahaAX4ogvcos6evZbTls63uywCE1Mud5CnO9id9fe
wAjKukxzbWkGptij+Xg43HCd044k10G5ZpSYszF8NscD29/fd14+btWDzb9NCHFVl+XfqdsFl1yB
FJm+kRNyjLO+dEFt6hgXEfcdusDGOf2scMrXXYIbhI0o2dvB2eNekBg2BqhItxlWZ2MUQjKMf7N/
dkJcNDLbAI8wwenf1OLg/UqpzwTCCjhdCj/Z7T1LdWQuqM/bMtJCzuQSNKp3K5cUyv38h0oZagNt
FHgH7RRULh7SEE7W6xRaYlOC3xBFomCVwtfO/smv9TcJ314zgmmHo5sbryeRtDf5MYO2AltrJKWY
64hIBq72h0lItb5AeVYbSxw8c79dcfSNIqHoHvh9SgtN3wnaHG83IQzIQZTQrt8vCzVvT4ZaJD0V
8z33Fm9ZzTtpMXjYIMCVAyThu2pVELcaEhko1ghLKbwDjmx6lbUuHL76GHMhOkUhI8ByNGxRJ8p0
FN4TPpsTyPr1qk/Kth2ujaXmH07eoIf9gi7sf2QilHQMwUrCG0EMMLoDT992L1ydUxRqDnhQhY48
Q/1bwSYCBpZArBuepsJYVeC//lchNMEk05FgBpcRpEzpa3e6DqT/1GmwmcfoGpIIuDlwzpOA8xsl
Pid9o5zgp7UsfIaWE7/Nvfn9r9yTgOBbRtossfgb6zhYo/7rDzKMrhM3sRbuaxq8zk9ktvHCL3A5
5i18ZBBQwowz5J7Lk/q7p0FLU2tjI2Ohab0XiTfJpmv1dVdkU8ocON4OEcJwdphIQOEzJl80mZJ4
scE0sDn9OCGRicX1zYLSnWcc9WOncw8oEsXY88T+7bR8i2RO2dA+ii4eCFFk3Es6lbfFclgyNXfa
x37lGV0yUEl1n10Ypr0QVxDI3G7jAc+Oao2CPwyPg302WHryll0530BPN20LyvfMC6qWsA7wWyiZ
mC1jBZne9vlIloX8/MtdFGIjkVe8f3fZQrCOgpYSCxVox1LjfmxpiSh+WQu6pnQ/h9ZhayJ/Uq9i
h7ZicExgg1bkJB1CEWuCTp4U8jL4tjd6IPKb8SZNDoxKl2eYBzuVLc0Py8eL8M1wKds1cWogXOrD
hvHpZrLnB5ALmRQHIngC19lV/y3OV4zkkCf680MuDdBtxPT95nvZH6v/OWYOMuzdlNCPHxUb1GmA
o6Q2/1R/bla6xUI/UCNUY/bPRkEyI50afc1D4cAboeshsu1kayZc+DJ5LJcUFvpV8eLicqfAqyha
Ll27r8gTjP/QIGG2lmEIcBC6IbNORgGbjp8YKp7pj3S4YRYl6avvncnS6rppSJVXxKEXxasyE5YT
tPLVcxO4JkWpTkA+Ah2dhN3K4Hg/JTOy8EUaZn1XvQQMOfMQEY01GAsZRrDTtuk9cl4VkohFRmBS
tExbmSddUaM/bNhpl0ctsGDw8VgsSoWCC+X03NZTDEuKKMrd9EPg/w5U6yVHiZhzVXE+5AcxpTPy
2uycYhdBRzVSPg98YBczGkaNnuSmccr/ENPMZo/aWsVRC+AAlVklUJQvhDDikZvGl6FAHji6eWM1
p8yEehfkgqiGN7F/KKdwXV2tltDKrYmUmdorp/5vT8TX4p2oq/m8pLxtHF5aYfCVTTbwZI8MTmOx
nHfNvmBSrq5b/qhF24QA87UYpxSWU8Vg3cnNwY1aJJ2aBVTlfG/HBVVwFt/QWoV0ka3wo3+9tV/Y
pFNOuYFYb/GTZY9nixRFmvaM6fokpItQXezTW2ZWacM/UPFTueTIzZTlgNgtW5TSM5XBD7JPDi2M
+X0yrEj82hBbHk6+aL3q73Kvke1+WY28linwpOpYVLpGUY6VSVML9/rg6SKQ8yN6LPZ9pCshM/NY
e5GtiTlMyTyp14Dh4SUyV2tq5IDQjrvhqT44upOoDFKjkfem9r0BaZjVt+0E0S4OJog/tsCJeqza
L9b42KgRn5xU8HncZ9NSeb07TN3pZgiKRwBo+mbDMzvVgvZFK4eVN64Ct9+pKdNvuehFi/M797IP
MGHQAKevpyrfdIiu4ncx23NP/Khmt9T0EWY1IxrM6nnbz/eZbvosvI51UzoRkEy7OaF7woHV6vN3
0JIAOZzMvkOpOYQRfkV2FjJXwBqv9Ka+B+kjf27sznJeLPDRRD8dbadPQY+cx5w5cNfGOtXvVULP
aqxPN6xZlfHBdxdheEPIAFDdYhIXWNEgYblxw/tgk0Frkyc+s1XL7bhbMiOgndDJOj/r+PuPt0xI
2enOmFBEZasUMzc/HZRbi1lAM8kXwWbD0WF7wIEsKef8sDYiAV6hVO5Se2Bl8Yn4Ej2KAAQ3kc7D
BNwZKw+7g8PrpJBYpdorRV0UXmgWERao6Rn9Z4EPTbn2OFbrgDAKM8bAFXaOUFgj6xkqJa78L+wL
QhQ1AxzgpzddnuKFHlCwc+/p7FhA/dC1ud2Nq3BNb91Hz29/SBa5wC/FAxM7YWhJWp/mi3VuKMtz
99dKEfmYVbziBvSYzOqI+rAHXfK0PGEuEQNMHrypBdrGOO54R0bb9FbifceVtvum8h7qJiQcqw6E
MM2h7CJUmVU0W3PFQ3qYwh7lcz5CVO+eqJjSHLoHqkb7bIkLrs1fUL40WB/XAmW7u0o4ByLOPs/J
6VH1vmk0Hi40If3gyaPzy3FvrdFxIQOKgmueRk8ykpBkgVKnNlnxhtRpD5+KjgaTHjroTVU4P09h
sVt/FWsi7awMuht4VAbb3MymiKBaJ/ocBqvk4WiVOZ+QdvKrHODIRSdUFv35w02odlH42h+BsYhv
aVuKzArjIpPIzNm4qES97326QwJfndcgsbEtsojVT1e7RvJczq5HFcPoK8A0wnfH0T+/2XA3mjN6
xkGN1ebRIuOuThzmP513ap9PmPqiY2Uf2y1EOLuuO4tTwtiS4DNka6/HxxF04AnnbGTI1AuG8NgM
W1lanRmccMDdY69yTt7E2IaqwTlQM9ZtGFLwofg/acJM+u+pvclWUhAec0C/Swq3+L7QsdoXtaoa
l2dMncyibrLhC+EToqzYjy7oUI0wSlQwmFmol1bh4traUCIrlcQPrbIYYxyYO634wnxz0vhcDEPw
h2JAM9zpQl2AX4lfKyK8pAezt/Wffi7NtG+MWMVulNEpexmHJlCXA2a1cl9QCGVYMoHR29YyzY1z
Nn2ws4s2SnFNlnjXJdT0B7K01jQAiuLRWzWZew2MiWEEq009vaFs8h+fG6bohfeo7smphOICbPep
5hlex0zqY2LsYsIE11Qu0aqMSl+q3o4X4fs8moDbfUYARXqMUY2DmYzr9SyB05nUH1017b4IbqJV
JWFNtHuAimXbh4XZ2pKwOziBrv/Lpk1DO5AkDVlt4DeEodrw0iEnImx1Y3e3Bft33SiP38JIiEnx
ph8IBmtNaz68piuMcGvqa0bMPpngMK7HENCrPU1hKijAQLfemWX96FoKE7Q8C1JjSJF4damFfqn0
AejpzfEbsTqBKLs4kHnXYKHMiAmvwHUHEgMu8BKa48bf+aKDThJp1ttTP775yjhEbYGeXz+0IKgK
A1Mrn3FTqfYwULfhiJhMiQKGqRbvn4tBnUZnSwcdTRZfYr0HAvA5oyGwemlGsoepG5U4ASUOW70B
s5ehYsdDZrdP6bvf47RZxMsMdSvQPB+YdTjCBzWq6JWWODESQfPmi+qZrKtIAHZVAT0622JLxP5J
SvLKQFo6TGYEiL5e7vVmp4gFSR/PIbkdkea8ViAnLdfAsz2i7uoGUoDqbIfcuQPLR9JbhEEjaZwT
/y9MH8faAgecpwN5Y0kCBnSaeqCozcbz2B/FuB9c6dShkwyq3jRLHsL3EWk6CPKh5jPBXHNnihD3
QXNzOZV9511jNQIXD15AdMYU8LIZmqRSMvIS+xuzrFr5lUZsmpv+aoOn8D0LHZhrqXUylzPsc+AB
AEvP2fj/tAckzx4Y5Lus7/a6B0guuZrrI+GibzGQwaV7/PI2kFQZA/D7iklPrfRe5iQpuAlAemOU
9Ze8I1523DRosWvMVjJypahaqIbhztAazOeUnb0OcsCg+zSadrZQ2LZnNQyG06k4evEQNAdXE/oP
ZBMRIAIBDixcWujCj6Wg8rglNw1ESaUvnUvUR48bQLmK1CtH6FyW3J5xYH2U4eDDOMJXWH/x6Oyi
TUocDG6ydzKvoFSuYjCtdSDdb16UFNvFgYP/9hvSz/+RawXX2J+4sJpjUy38XcTP9GYt3RforQNE
a5gdmRqiqCR+KFwW1T33tRgHCAROst4+H/vTzxgPmRUsDPvACPOfFZ0Ptr51LqWAoFndvJGzILzk
UYBfXDiaN0vmuRQtaFFSRBUNre7t5jeH91Qyzu9t9DUKFDsvzYZ8bbPkBPRHYPt1K69WgoFe/1wP
HHxCxpIHudbUB1NF6tQmVHagZLVm3VHfiYBY140mjhABMKro1Y60R0NKro4yZvndI6M2g5IEpJXv
CoSS/E3Zd4ph5tIaMvbBvIj1aprlr+TKsL1pbHC3flUQdMqoMuDLIWrX/DQNTqajRJS2D1yiHe+4
ckDVK5y5aik7byAG83vgjwseQGhNDVK8g061W4QmewTxIEVJifcLMe5PQxM8pe861sqL2RiFKpcA
fEhm7elHTOHMSsdyi5uyXNiMRmnzmmj0HFKRGQZTTj6CMscUuP8Rsvaj5oxpXGWRMpP7adf54ipD
sh/kcsHzxPfWzP2cXzNHkPE4smDOz9M9YjY06249FVqjxXMPXumAaUZdzGOXGLV5S7kRhgCUgFwp
F1vI8JOSnIzit4bBDXV5ft7Usvh+I54+v6lU8Qs9LH/tVZGsUDJbyRFMYl/mWJSCzs9w6qZMRU+X
5DPjn+R4D448VzNYrHBTtUIefSpIXSDMtZCYFvI2G99BR4g+V1mxqdR0/cKb9TLWW202mklaR/pP
yxtk/1KpONZjplkCD3qk9PP5TAAv5rQjsy5kEBG801cSyh2ubDnkFfWurrQHjg9QcUt1kUT+kPST
ReRIRCvKuyMXGjSLHzsRxiYDFRGhFEpTc8hNWoo2z9irzZ0q9xaEs3pJj9FiLOgWUtNGVRJ3Bt9R
WAlcX9xwB6WSQvtZtjVmv/HPlRWs5Ur4feNUBGUtjuJ4Xg6Kus8PnoYP8lzBsVz0giAWkoz2gbdW
JN+/bgg/x5Q2SCExtkUOB2NVOjiOTNULUtzfvBVY2Pv6b/xvhdjwOAtVlaMbbJR8QLnOpJq0cLj9
zoMQSmtd3H7nbfMtizNNcS4zx5XxjUpiNoh/RQ0Fj8J41hfvmi5qoYjGAMxhleeTfBEue17oUQa1
2BPNFyJ7SdA5hkUMSDGKz7MT7sukOJ4NjN1HXr/6EyDjT3bSFm2UC7ptiddsyS7OJmsqiCm0nKrk
rEiaiop92dTiFmFbQ7+npf8Yfo7/UPZ6sS4mJtE7F0JhhvUuWPRjd332tOQQ+/WBWEO3XEavXj+z
MMN5+jTivUwYh9X+jSJBZe6xLZAPu5pDgl+0NWRNjbDjsNi2czSv2aUdnfNMcXsJrFlVgnSSUyo0
X2m+oxzexD1i3XtFIUMai8/oNpYgkm01z9zmy9eX5bJsvpO91ksRe1zCEhhzEtP2GpN8xIIv5Ode
77FwEMDKsjEu94mpfIv2moXYViZP378O1Fhj5H+xjdBDFRrsMzY3fD03hpl1XhnxzyD0j8gvEHKi
RcbhZ4+M8bt/Mq5SMBGM8WlVaRuftoV68+ZbZnXBZZsZO0ulIxQa5pDSqcaAIeyjY7f22/H0cG21
Grm5IcCAOx/q32CRmsFlvT7arjEDp6QnYl/akT5Z2TEj4LSuUtzzYlDsB8lYUc4eCjF74KOfkvH7
iy2M+tcWiDTjsWCkPCb9c2v+HfazSJoCeWwlFV89gZ8IIvlPvDg1Te3GOI7TjWAzgaroTekxTr65
+sWqMpxXg3ATdZ27B5YyT81lxt7+C13XiSGWBEiKmdN3yARiDEOFzLqob0Xerv+AxgG4B2rmITKW
D3JqEYgsaOx4DCHR7L9mAlGDwdIB/xWvpntHHpUmb2V0ol4MDsntLypi5C2a17umnQDdQ+j1z5FX
+tBjxG0IvF+yX8azOJEli3I9R0Es3DPsUEjHDyGvYitdyFlX8Fi7OpL8IJPr34hgswhCdsoxBjDb
ljx2hLWNWbzLu098oEYrePZLjYy2EHjRFPk7fB4GBEjJ0YY8tHJKzsqyCu3E9E7tsak9u1SqcQnw
vULZ2RxkftlHGkd/OfHcvcI9ZIbSo+Uyptv2fKwyLI5LKqWPnvtFjBJUqlJmhRTCE3k7T7p9pdzf
Yg6V+V43xLxlia2ByAF76lhtFanWaMOPPXButZbhjfj6Eye74b+WpKlPh8pXGchdNMQq3ycKCBKd
9vGoAxcCFzRyZS1eSAfLqwUI1JJBPXDPGXmKEj/7Vs9oQodkfrVgGqSV8uY+Jn84rmfRUTBvEuqc
ukC/28gdK0PVm5rHS9fbINDrbWiiPSX0TFbsqzMOi4iNxwhRvkv+gD+OlMQ6MQYN8Ha+Rj7rZeVP
TrgDs7NnO+WQEWwiJ2YxbeM2mXYuquiBR27TgawcE+Re4hdcrSyHSx//a+raFoNCxU5FFkJEJ2JU
0JNwiL4vXsbpZpTSUr7lOOPlj7IiMpexb74x056s2/PqQjrxSWDFcumokBTEN2u95SSKhVOX514g
7rWyYGwDWz1i0LbilJ1yE7uduC/gkyq06UVinDq1rdT9gwpuv3hostWQYddVNJ4V5LPzmTAGIQQo
AZcFD09FDwQALyI8ijGH5hgsBNHEqfGl6DFOIHWby3PshFW62baJ9moGm9U6jOVhKf00xEMB7BQA
xdhdCgsCVeHeCoDNsYoJX+kvs+0gEs8QmaaXNE3BSgg1dh3zSia5/r97dlpifJBi30m5bhO1nN2j
FswksOYqM2PhmI0xcw9kF7apr/x1F9GEy97+k+6n5F61y1wsiGIAJFs6la80ST0W7P3tCIlhLMHT
GKfghpIWY/OaGqQOI4t1uwLqoLe0akv4TSBd1ZOgrf/Y2XMNy8c6mm5yNJzWKerHbsGiugmOdL2W
CRnbILV8SH6UtldVVpzVSP6j692jR1lUSt76xQdnYA80myNAVApYMF8xkfX1mDDxU8N8ZC/+OUdY
BSCw35PsfgxcXaJDXwvGZtExpS5bCYYlFxGHthfn67xrNS+rvvkA0ZjlsFOgRinWkspkoPh0tyqR
mvxvxD2F5PP3FpVY8YkGoK3LVv/1A/agu5ekr0AzgGXU/RWEcEaqtJ3JjQDRMuTd1FJ5swTINFQD
pe/Jz9IzrgWNyBR93zXj/Wj6v5Ko48CubBrY+irqEOWYLsBAKTdlIIWec2EjHiayPDJXc4rcyOlP
JNOz460ioDmizIGqOvJ1Vzx84bEBW+XHTWdzqeVe5OGqgTTAcKdvvBKnFeWLGZpKZaYAIg/IOGNH
8pSEkYglBQIjccxGksmNVAwGBkYaAI22wn3c/+VTlEh605UCAfzRgXMMcWzlc+3sRd4ePb8Aa1dw
rwpMjw546STb1aAFoZQl1UldXs59erPJx+zSgtupHmGWsJUHe0nmT6WnEJdrnYxXb9+oEtnF9/Ht
jG9lAt2haEj5QVCRTkLDgZPvVRLTX7q7lzDgj0vkwtryKhfJXZhNH6gbhBSDELqscA+ltth4Rz3a
w513H381gray8pg83CQLDj+psWypntSPfPryf9FY2SrDSO4Itq+0FTOPV6A+b6V6YH2PbhkLPh12
0A+qD3TOyIW4QXNG4lZDjDpepLK91vB3G37uZQLSG2rmM5Ce/IVf3gXsXRj+aiWlGWGPA59Fosef
TmsD9ElRJyLdYQBOPyKJ5KfTQPMB7hFMIhVMJiJouYZkPrvnE/kFXpdKUFi3EEeZOGE3H5U8U4Jv
6KxdFcEa82ornUJgkN9M1s99U0N9hSn3EFYDulyBJXyi1dQ8PvCDddqG+6yPmD45kkv2hNtS9+hP
6nQVyQuV5AzFrNyLJ8A4T/MU8+acrN+MUvirjfWD5/4hSCrXuWlHAgnOI7fNlSOKh9jI4y2Y442P
rJlcRj86kofCdIeTqaTbcfyDCs85shZe0j8WtGht1YCb8Hr7Upc7NH8T4cAP8NXnVuC93MF3akxa
E4F8sHetsJyRZaWo7zkAlTAIJstIHG9/uQ/EqOGTVtju1ZvZePWPOVdp/FBpLsBQrKqEMmDmBN33
2Jh7NWn3SRcZEIgCzZypOv1DcaZNNfT7k5wtLFvRw82pqwK8hcXeNj9cdYFTTnrZa2aM2rjDL7RA
vJhdrvTpzXcuroaU1RKN7rh4rY/r2SmfP50rClxapfRZDaqeJTEeraKVr+/hBWre3s/r4eIJoZG5
0ziT2Kz98AT3yl6edEXUolYggMK9VO6DCSYESIXNjQxkW2mu9rRiJ+PfLu1A87FoBqYSmgGa5wNV
dK6XGlNQ7hryPB6Roeal93BZGVw/rvfDIMz1mP7fkdRgK9eLcxbJY9aAQZBFzmnrdZth2RBW/fdI
Q19i5374L3br7agHOMrgBOi6lhqfI9/sdl+tm1XUdu3WxSS+ka8Br68Q+BBi/LmDvvslVxKFud1k
bGMInz/qgw4jCg4G0+BQF5kf9vxzWg63LssHld0P1Dv+xIRgIp1VPbpdvR9kTwwMe/yIDsYNj8k3
Ii/uTTLDOL1YYz7RsNTGqUulDeS3C1DlmY4J/85IHIyus7R4G4INaSaiacUoXzbdn9SvzvgAAGSk
LomCTnNs38s3zBnRMBONQnbJugoQrUpXX4vBYObnycuk1fkEmY4DaVQgEugqq0IJoGYFmcEpUoOp
bO1HYcIcIucB2IjhwJfRrGR0EpVf/W/eaPfbXTXWOrC5C+MMYIAjtj3mD7D8fec7DZpyxPpuMh03
wK1MAvlpp+Sp5qjaKrvMElhYvfcG4x2dphl31CKOudTqt7IqsOKGrKf+xqVllkZeGvqy12CxisZN
gXyefbR6th5jDS4hedoRusi2FuVU6i4fmmWjlNzVvHne+tmUHDBy5/+5UXTLqJcky36+kDqSOXp4
43Wjy3Gd9a0QY2xPWZHrtCe2n92K6ZnS1FFPUnC2bADf1ZVIHu5Z4rATLfsZ5d5+rhhlnsxx2/pR
/+CQ4Jm9iwnkod1rhdzXior2cVItHh8ul31xEt9VJZ/OWWUUZK3iT5AhW8t8SvKEv46qjtKV8n9N
rL/FbqyaZSW/Xg1OikHpE1tP+utLeFshKnIy0SAsHZJhEH9L88UNh83l0XgNn1C1AEwsbS0uEBcI
pRjbQI6Hs38we3KWhEVhCNFLb1W9TLkQiqfqco9hITWcHChbRpGFwfVOcNehRHvydwJABUwEX10w
p8XwJTGDvJ9rZReeHORQe6gx75cPwEPk8mk7kHkU0G7NdgY2eAQHpcxBbEMmdUf1GpPe9sZcsNtU
9VnAj3M0vl2RZD8KZUKqf8vqExGOQgrX+wa7yndl0lz5+yvQNFrmNIw6ldgcfruJNLJ5YkwHvv+2
nEiIp/0y/UZe9dK+DJRgFImGaXpVAs9jk+ZG1lhzdDEweJxDLHttJTt/iqHamvmXNt4T20Akx0bI
y3b0NbBOhsmP4vQJZzABhHC0vQ0z8FQdtcvdnJB4FxzGXa4TbcOZaBNNsA2ukfgwfdaiPUBDBLIq
jUzTcQkyPujiT5vVssQpeV42Nl7mqADuFf+8KmGMDZPdrEESmedVmPAFLMwLb9866AArz3WT4dZo
MS/qPHKvDK9uupeo9m2zpaQymDUhXoIF2+ff8JbBogNu/XpKzUGXeLmlADlIR2YOZ4rXiyWNGs2K
XDu68E4E0JM4qkECMqZonkSqBN6b1g4+D0CqSvitVLLkYlHs2+AY4y6ed7DKgcY/QxWNYRwMmdmm
9OJPr2cth0J3QUS2LBASLhp9xW0/j6j03s09qPYWAUzIobuSTL1O4qPyC23YsLNN4kdiku05pckq
7zT0tBpxDBxbZ5ChjHnuYM56XwFX/prM8KvdNzUNHrIzfct/KwaQdG/hXFYSdRkoGZVf90zPuhXn
k8GT5Mo9DJv/4Ocj/jPy8wukBcXCGEs8xB5txbizX96jJmTF36Nu2Js20CLQFa6EtLIp8DbsZdBx
qvPngqMmiQ0ZOeBwcs3q4iHmL2pCLfGSbBpg7Ex8p7la/OFsESFy+BvfBogqIBQFcxK3GtweYGk3
2qGXi/+ttp/KUxBleeY36CsOUjrMFOHbqJ9axcehCXD1kyI2VjLv7CLvVIrnc1OO98jRuPnjuBR2
mxntsnn/PKR79W6Uz4sKENgjVl/FsD+hX00QxHiI2kujYl60FCVdsrthd+XGEIcgBoTEod5yKmoc
4MEAWgU27f5O/x2tE2WwoZXHijdx5K2ic7gR8QqmVL+3PHngITRL45q9MWSxgNIV20hEyX05bH11
+2ddXiAPrYhGDkKJY0OJ9y8rQcMo0X/7K9ZTUcui+zR4lbJT7ybH2MzoDyw9inEruDSYnCzGNPYP
7udWzEjjlUk/NG9yXku3EANPe78taEsoHveCojZ3fu3ZkFVrNIq0sjHvmuROcMROrHvT6EHK8xb4
sLcycYw8DQkHJwwIsFRCbneTxjA/pTLIoip0XOvUbZATynNsdP/HIrftRnTq4DlB6yxAr+Ql5/29
Thr3guxjMkQE22D9MWJhYQu2Kv+/4oWY8ljAZcm2gMQDfkANaGYG4JY299QNCa2ccV/ijMoQPFNZ
zPDShhRdNrD4bamErfmJmSl+pu12EVcv6i82+74y9mTzfDnwn43SlJdDuQ5Shon5CmhbR/oZWAUV
8GulhRxTSL/Yle3Eb2qWoKEhxMik6yLHmK4UkOJ1x/Q/r6lXx/CwtDTplZR7h5WW3MMmg8vWDO+c
rBAdoMTBf5VN6YxIiirtuomypHVvat60gogHTKFw67RWFuYMwptTDdKW41XpCsCAGrh9cDBuoDrS
xVgKI5Papd/NaiShoGcg9iTE5e6jyoSPUW7beOuZ+bHY5+045jkZ9Hc4Ic8T0bgKnbTcaEhKuNGT
3tX1zqplP0dd2pyDkhIg6rpiEY1Iv+IT+aOcrv9C0UtmL5u3S2PgvCj7FRleeG9JFMUTm/BO08ic
gTi8PnTWowafs+J3DwyjY5PGO2+5dcpb1R/WQrKAZGIogRUfuwiZ4RUqkrIjTGf6cBsynCcqmnRr
NDNR0ba4GXtXOAIdRgQ3ET3NKiulnUoKZot98qda6OQtvOPFPuHBmeMJAPWfH0cKoYBj2h+SsZ7R
LR69661WKHtD6PPIsME/NIpBaEW3LESPj64tBgCG5rJ5aOFceNhxqJpaNcayKiqlT5UJrXaqEac4
cx/6U+UTkPaoadMCEWl3amQnN5Nie4efeLLee8BUPlMXyfLYXUto7XHEuimZSt/Pwe7ZVGrEMOdp
tPa+z30z9crqFd6hB6Gnmxd11W2X3VeOO6Gn4svLMHtTaehwD8ISjYCFEEEqrpOqRfH4fzjNXzp8
L35AoeEOoNNjXHHwGfyMBPna+XpNhTJiDANBYYu2w7NbcdfqxG2+Li8wh76D+5xBiMNS4tk3VKYi
wOcLFpEF1pUNrb2pL8vSgMsEtHIPc72GYTyL8IHJ08ozvFe6Xcj/BvbH/jSUyaheq2H6pFMSYU8N
vHfapg74vq8J/F3G2s1Y0bGSyC6GhLg64xd1NvBOpmJ3RqCS3X5eAonoYg4Rs6MmSak/CeGJGbI+
Kik7YBnwAsrLlQaTSPdN9W5vSMG9LnWjfi//Oc+kVKU/sW5xb3wKYkpHy+2nmC97Rg/oqBHQF/77
3VckviF82xSBmd4HwMVxfhug8LOOH1LBaQEyS2FHkzNRBPUmAw8F9V7oTUptqwwatRtwTGGmnC26
S09LYUAURQo4FIqvTQYDE7gE12qCHPprNv+e8LaYEPkYoH8QVQkUd3LnQQ2BM7a3Sm3XK4oj6gkY
5hYR97kMYfXsAC6/CiMOA+GYQ3IzAC9A7lpuJdnux9QYL9ccyJt6PyR+r+lxp/shHro1Kbg6SkdU
t9N/RbWYHux6CNyNp2KTYa2OVtLIooPrh6BbVMSdZ0Ma3a+PfWdotIrNKAP3J1t+SIUkMt6Z2v2R
e8ZtF3fXE8KO5H+xmoojyo2SO43PcGLC4qvAsyBTyvAojsORPVZKU8ZUzKa1MALg9XmVlSNH83KQ
aJmGNo8N4lhmbh++VsRXXVp5M2OIsvlugf9IYeVzDcp7QlzhEoWdovezITHwVMOJv+Hqgg0TePup
K2JvikFxsyBfY1U3V/Ou6zjbA6hp9fU72Fj5hzhCex6IIXAqLWp45ctwJkKrGQTe8NS4Mh7PBJN4
VDXcrLL3xjt8XPO7SWsJ6MJYD+TRii3fS8Ys8tY9YOw1T+TT8dJA8f5QFAkwIgAkANMppN8HHHec
34Ild1GmDej6MVtG8UF2SE6rwW+9pDm3i299GGRoGadkpw79YcMxr9zp0R/mEMdGyOz/aPCIFvcz
0bRbHwbjTgsA48CqkNaexvk2+kJJnbIzP+5q0gv0bBVs0S1Bm8X6CiwguB9CJlX1fgG5zZIjf76g
Kj+SzAXQnRSENc4gsfwTr7qvkDDZIVgH8uZnY2s8G+TcSBbt8ASnXoJuqwiydBRgp9UA43losrDb
BTtPE/OmuGRB2za0nMQ680HE3wYEhBt0tGqgXx9BuGbPUVB0k+6xhkN2H7x/3RNwxKc7Xmpbt0Q3
NnfJIerhTSIs+CbHlAdg4lojA8xMaVK7dbfmVzRIlZ8eVCtvd6LReSbLU8Jav1QI6f0/bRe3Dec7
QHjaZQJRaYdN7aGz9MEcqGNH1y4cdVIXgjOZKB1nuV7HZDMQHWpJABPTvnj1jQ4DYRlHYiTRcs+Y
tbvZhHVIK8a5iG7xsc5C/zV1COcXMQoj9gBxUI6bJ6eQ/ds9ro+cmbZQL9rT4cE1sgzo6UHRWck8
HM5HNlqXr1mMzgfnu7pRbbh6zBebPfh1EPOpaiM3/Bq4x6ur8FXejaJ57chUz1iN7ZKhCzFtfd6C
WseahkdUn2tB25sBm+wafKyQRU8RTcDGXuyeuJsW90R02ZG2IXpmPxka65guFFEVTDVqvQ9aiIux
g649FLmhhyGEGjYMyfQ4M2+CaHxF69fDTJLowtdEdr5upk1ZQhkvmAMZMPaZAjlwpEtnNROB1hts
nVgN7JXrasz/oXLot5kSaKVBE8fWnxZRf4Q/GZi0CORjJM7hziPSmTvlR+O8gaPN/escXuuaGpSa
lB4mvJ4PdOBvCJqcICwtWGaPa/FuzC5/eu85ZKRBGiZ8IW0K0lrPEfmkwhGq7HAOfjABg7GxCSUK
LRoGv/RJ9u+MgdyKpmR2QrFCBIbq6ZsDXsnHFAKYww9Lfb0E5an3dwOv7l2n5MrLXcSxSwpzUoa5
JxJOCnqRxeGygp/EIbLpQuCdJl6FQr+GNMPrMG+2ZHk6lyKOHv25eYhjXqSOs6wd1pbYKPJaJcMk
2yRsnexEdU5wjnobrZGdC7KWsz8AZwZSUh1gNYiayjhSkCWVMzSJEZ9vwzIOaa12QZH+z62ho8vr
gZn1fnHAx0HmqPWcA0UuUr6WNV81l/BR94Cx1avqx52HwRrAkrYgVtBhIY+TsCCxQbtEJnvRZLSI
j+o4qhklik5xpa5xiFCs0x8mtxYPdHanFVQcm1ZJeLeEYUr9gV67JSQEKWQW3Be3w1YVrcvuOR0b
M9mAMzUon+hKs7jKFBKyhpKWI8/WmcRgwHdQ/B8KoeJ4xKxfUyjj4jLzfZhWWIWgSXU87pzOMngB
GBXun8lwjtMu2abFP2Eqj3QhXNCPvvkSEsQyA8OyCls7q5o1uFyBrQikHLstA1dN58ljrjxt6yet
YDXM/FNkNBPvMsgGmW/4HJI7Sbhyf4l2RG77naAnMFbojdnxrXUIHYoyhtVF7hi2ybNVO8wqFHq+
72Xzya+vy7lyMWSYbqAagw9HK20i1ofS32x7VXces0VuiRGBP4THJtbYol6alI15JVvedGb7TUbb
XXERoZXc8beiFtx+ItCJ7HfMhjAXnHhtdOZJdqe8xXlgD03P9gvFqNOcuHLrMMGx/lwxwe0moGkO
d6mKremfB9XIU3okEjQ/xQ71xtmtgpOsPl44bqoV4oguzUSWKtjJwqb0argXY/sdNu7idy8sXNd2
3/FHf2VuXhsKH0ZVdJgvzaW2y4Rhzc5CCMzHpnOciWXujMyqFoBhauHhSetvLhRroMR/stwJa15e
vyBvZCh4Afl/Fns8xXb3RwJpHmfVKI+l1x21tSpcervVKU3FyIaVIuWQq/kigUAbh75/HD6jqvV1
9VWRwSBjdnQSaB6RvcVM6WVY35nwDV0KYZA7b2LvwOKhVdFfLGL6QLf/q9xYxf71tqW4FjGFjhOi
p+KqJBpje6h0uj8qXTF1N7goMqmjcoAyrw/BrTnF5jOrZtgRWN29cMCm3IHrcYTAYVBwSFDJcPNM
50Rehb9iP4tvrj/5eN0sh7NBWnvFRbYRl5mxhrRpLv7e0rxr6Ey1O8PGPcvTr9NPNpxJ4Zj30y4g
p1g1tA9dRurlu8WG9in0ctKCN5U9gj26luZtk74UJR9JX6c1suwm2SzgESnWcYAq7/8L4nj/83Tj
JwbmT/WOkTNm4CCAGVRjFb4CsyTlTNyr1QyEgyRf9GljnYfP1kjJavzn9XezDD02OkQLL2/XM7Bq
hs0ssjIXLhNmEpIsWCU7/hwh43HBJHzMNA2BOAgeEm2aU15h5L7fOT6bkkCYE3vO/2U2HsbpVMFo
FleZwZ9Owsel07LXEEjNuYKjQavmMCNeVAr50EwtNI1RRPSCba6TPrbDKTHrpQwKEmJaKjq+Nhmf
LZJbW+e9UqGBGlJyuc+WX1NE6OtonfhB7h2o8uuWqRmiq8eEG0I4Vi0AlN56YzjtoVH0300pZd8M
MxXix29vuxOVczTaU2fiUSOm4C3PpOTZHLe8R+RnUsphofGX0by+13yqZUInxROUH3T5t8ulYHbL
opzvcXb4kuAxH6HHmm0SU92Os7vITgfAFrEFTiQOWeviR5cGR+F9/yN2lp0OmxeLkYN6grVzTiEd
aakDrHrO7tBumNxfNbmB2huVBI9e8CsVmwxGxuDi0RNiD4LsvA1a6yinSK7wE9meodSAXtaKn07k
JEYgwbtt7e2X0gEmqiFjAJK4pKzAD8KkuEXwyByt5gQ48AvgXEN6TnKEtkza7SND7PtdmS43b51t
zFXSWZXAsCkd0Fftwq1bQl0BaR0+ZBFSUF25KS8LGyyxwqYgrbLg8718Sbo2B3ysl1UEFV7PF6G9
qHd+WCQ34WXMOgRBYAms3qOOUnCDBNL4wBK84Qo9xzH1eo2ASGw9wIbJu0a1u3Vx1SENBX5EB3Hi
nlx2JxJIeGxghTrIAQRFHVvK5c4OlQm1V32lyQdVSmHI32nn22lIHSXzvVBB85W+wIxel1YirnGO
f9WfWMNP6XmJfRUXRKMqfcQVZr8A2d30GLi2ZYyop1FC85lZ2PGT/P6RTW5uCNvepIFtU52UENCD
BwHoZd5j8ShM+v19QNNa7ZqrWuzryzNg/sjvWkzjH4ysikaqUfYVKcHC8ee+itvgjeSYCklozpzp
3oN4zV0RZGgXVNLoM2/FdD/YNleR5oS0bgWJkBzPuxNuSX1Ba9WRSDUAo3b/za9pBO+0NUHvTpZW
TAYp5luZDg+TEwKTDVAz6NThYSq+EaqYOXNKXig/IMuoLpq9wmfukoeGNmhISw+fJQdA7eqOVG+J
WdL0rjiMAAeAfwMJjCvjN6bD4Zp1QUR/4mFtpoYZ4c9iwNRlBAj14cCQuYHgnVpEoxmM1dqsm+xM
Bo3lEwlHLqSSheKExwrShAFWPO5vEAVeihnWp1Qkz00gP/rN9Y/JQLidF+oTYCXRry7dIop0xwxd
/0aYOvMgTznbAsqfSqXhqr615vjbui0bN6WWhP6VN/ymRnAX/FzO4re+lEW5Dia3STvhz6fwdww1
5Ih+AaK1UZwhCDnF7Q9WGMmL9vwNna5/l9uH1DZt69fpdXwJKczN+yuvev4JAJ30gW9S5wf0InbE
rKqM1ItpnTSKMv53ElIgxw9l3HzO2DXGKFR6TDcdDTOBxSGT9vXNqbu/VVB2+hsPKxaTViMRlPUQ
CHrNhYCNuFbYW4VXjXwffczT04p2afdqzXWRnej/WmEmyxWRAD6m+tNZoXSo32/e1tiqjm3Mtnbc
cqc97Tr7ScN2LeVoWWsO1dYVvRGTo6tRxwq8JBQFHSpo0IlbCINJRgq15C/59/wxTPmNyebBqdHj
9LzC42AmmdFQ/c1U6slxfqqm63JeE7q5tAeQyEcQ+xAe2bFhsyYrOmLrQXl6X8QmbDEmWtBKUMxF
6CzfoxYqYv/2/gZVJQkPH6G5aiX9VkLF2sKxCZhTUv2zywT8c0fYSCOqMjs+uOhRn26p1zXKJnuZ
QbVpriZPKlzp1JBcdxlVstIJhn853U3EVvBFGhemjigYOVW75sD7MDetN0KJzn684BqCpMyq7hEi
e/An9OL00THiQ1BhGCS5c7gKl1Iww8O4opWyiJq+4+eVTGpPSUsEhshLf8qFWHH0C5eegaHZ0wJw
Qmr3LBL1AOfOF0wwdVXHkbr3T8Q0iSCc2amfA90ADNpBC47p9u0nTZ2y11t9GF6lTtTfuZssrbgQ
rjktqE0t6i8A8C3VsCPtPIt6y9ywW8tYHlDyvWSrgq2Sdyxqhbt91/JOPfe0mNCRjhRZ94lvx3jI
9i8DXae4YHuCI7RPLDimfk/2HMckU3clFv3vCPwEDlJsHdm3GrA/WVVehli2jCjxqqIjmdJKYYnf
Zo3C15Fu8zIqTvc9nUiU8qorQ3I8fpow2+6bmVBoDSLPk4CrxM77cSA2b8EDD5hguQSrb1VBlrPn
N5X8ZSkvBQEXGJE12CgAjpnYHJ8FfUN/R+0sxr2/Z6A85aXQZt2UXBHoC54uDtLzCuguGhpVr5Hw
nN6LJTLGlSvjxAWMH0gA4/TiBYFz7BU34lZqubt+MPmjUAOuXadNdLeQhWysDNTcC7hQUps5R/LV
Jro/sdeznVY+tKFn6IvOhPn8V6cp5S8H+KEOfIoqcEGvELBRydqSjcJUA/tsDeIDu5gQb+yRUm+0
HP2ELh0SBcacINNsucinnhh0VALbMjdkJWCZvcKqJNE6wi8bYYiHYVthaQbqVSE2Qn6azTl2z4Mg
Vp3B0iJMuprIKzFca8KX8ZAhCwIuHrD9/cNeSAnOwE+JT1yYBmHJq+fLhQtYRJS4XuoRAK6A+tUe
Cqw0GmwQDOCN+F/cbcgCbdA9woxUGw3JyvGFys0UJvMmiDqqJpnwDirUY85ErekDhnVzDLdFquva
Bz2PHAvmtpd/qwdZXz0BRcCRwJo2Nny4wV6eeetIx++4jTlFrFWaWSPQE//Lx1h9d7lgz31ucAyo
jVOTXc1xtro7CYSGtKa+gG22V6rFRW6NVBa9Mdd2gvJDzXenqOqm5PFvIOn2VvdSsYRoVeLdsoL9
EF4H26uKJES9SNNSttY7UOCoef0gTSua9s+1okKKLsTg4r5GuXIogGSvuEq8pHUSYE2ePS8+B/t5
WByjRu1p2y723tIFbEQzzYm16CqaHm8stjCgPq3zXFivmTL4LAXbrskCg1DoqjxNJD1GQnh/oici
JLj5OfrkC/rdP5GNkDlmifCiK/Dl4oxey773iwDa+TSfNCl7fcbzio9CeO7P20vzhcXw2fHRtV7l
wVA+HSPEyZyW93vcT0VJDnmyQFcqwxEnQyE+Elhrf4Ot2padNWWvoulhCkaKo5t5UROVDcobLpNP
cTj4mooAKIm44jBBU4edfk0+oejnX3wcfu7O8Vsg+POJ0a25IGbYhsKPpYJbNPxHdzrD4rgpQUK5
/e/u6X28t2/JDeYUz8UR03Pz4QEraM8ViMjjSWjwbPiXE9rt1KEtCq3/kTYTt1n8Wynzc/8wSWMy
IH2J69auypI2s7/bpyZwfweLaEgTfsYl1/ev6bVYPeH7xVJ1Ii4I0lkrm2O8L/JJkbfUfQv/H/Zq
0LEVWkYZk1w/i40NtuL6+TvxAAFs2JhcJ7FrQLVIUYuGsQ2FtDS5qhkesTcSmMrXQMWZjUTFiVoA
cSQXAVZ7SuvJzBtT44WYmwNrrlRPy1uXMKnVaQq5K/IxgfLwhWW2Z4A3E4CGL+0ldH3Oske0KKmR
oNUuwoIPbcc/rUeejdmXULTeo772Wn4l3JLqVJ8pfoHI7ogbHtlQYL485sC0gplFC7WnofE6UcC+
b8gTZcswlc0iB7ajUI8RWep3kO82SwY4wn7KTCzXPIG9T6lcWlNyinvVz3KxpIS1CjwPkmnlOGW2
TqN/xED24WPuju9CZf1VktyM+6ZGabxeVM77uUovd9sdF7q06Tqnd28OK9o7EK/K1MGN+sEZhSfC
fwf1hgilMwbAuembVxtR0vi3gDzILDTtauWfi4nHoVAedVKVSfsq/izmHrGFRJxAH7oOlbDvYA/M
WA8gCiINQvSsEJfsWMFEbhGWlaHph6fqX5Tri7ehw3BAH/zrkgLe8ysAEwy+2OMHohNCIfBS/nap
FE+AxG5kfPWTS6lfBeWiJiyGwfxXGnlHXzT5Kvha2StbtDUI51BxU0DzZuc2+xQPWh2uEGChZILE
ng6a0GoCD/t0sDDD+fVCUYUb0zSWDFC4Gymq4v7Y383R136MvF0bPSAecY11BN/8ENNR4Mn7tfXQ
2kaj2BF7P7We8md2Yq68FXKXv49kIo5MT1O3dHcgEzEMlF6nfWJRpFtK0pEojnpqEwoizr52Rhb3
IjQL5PAL6A/z7sImmdIx/F1kzODlWrrSpUonD5mxhf3Pf6n7mvm83xo5dzRCo8UWicTrKtn+y0+f
Rrcur2jRZUeSgf6p2dNwcAAW5Xk/xL4EFJRx28uF7VrcsIfYjaQyvYAxh/ErSxBqXmBr6+FdTQeE
9C4Zc5ikx/sPQrIDp9EMX7P8AwzZbcHRNorsPn3wE5FDjCrrbwuFtvrLf/g93dZcMNRQgV4HuKHD
g2ugjcj5d+iz4mCxmKL5NlHpH6MVilG8aSuu0jS4eVRbpSC68DpoWKm071WYWzk3wCpGfAVsbeCU
ZpXMEMi5qJ7FAv7Q44Kqt9Q8PSxV0Q7boL3RMmIgy+gHK2I9GjDc8cDF1+7fslu5+MIDcHtC9Gnj
BIAygGN+3pvATk4M8PeuHLe+GSNta6v1YItZg/AMI+e3TiV72crOg+gaxsI8igkxyDFiNMSpuzPE
0KlFYxXWhAdTMajnjqi1soH0cGCgj2nLapo6fGD0u7pQV+M6t7nfzd117lb+PR9yjoNbBk9jKVSa
tXb162QZ89i08oZm1viwfdziKPu3i3PhfN9/4MRkr3FM8LhjEgZHapMEWOsr9tGNE0GTLsRGeIUV
TtfNFKrz8zIXXGhI+klctBYb0NJj+qui6cC4RP6Fankh51Y7zWD8hH+zc7qvWlVUkm/JQ7r3CzNV
JXb9PENC8S+QMSA5Hi86xaqG6W9t4dFfjiiY6FhF4PTDGDTw26f6gcqe2zMPdhfXOj86FXTrCy19
/u9nQfj77olrjXIw/U5Rb6vv4JDnRcZg8CuQxosMwvOVvd3DMOvISK26xmOmlYr9y/a90cbKlq5g
+aOSV/0gyH8D1Oq066Eg8p7QIQrLRhpDtduRyqtkTGvG+r+emmCbaAN1ZuyqI5d+pEX/wqoH+vp8
wuwa+qgLx2hQILu8Q+14lg2GwOR+hESy28ZivFV7wRVcCFraSK9Tbg41/Nq0ed6t6zf3s/0eZtGm
xFKhBXUmYlTO9QZdsOegr27pDfves1gZWs33Cr+brRqZOysyGAIMDKNu11GDIYpdSBmBeYLgajoE
4ikeFTvhc6VfhQuGVjYOmL97V5iycar3QEeVzSeKR98NIBAuRH9NYxHDIny5V82tBhfhkmYUGwow
Rah68UHJV8jRF6J2/l9oWEWVXDWLbDUjmlMCalSQlKh4cYzrJ5/baG3hmPimeafVCVuzVxL7rVrG
vcGxv7thXFVvGNk17QI7YLvf8HgRiKppvUkyzYj/Bwgnw8f+lW5an+o3fkkVHDnGChXwQ5AIbpIq
K6ABfSuIt9XKoyl9tUFAw3AnnMNSTNnGPFE5v4EeJI7+ofgmheIb8jBB+VYKzole1WfGa8ZQjuU9
GNRi2x9rKuy55pTMichSR9fTuo440/s4T/avy9HJFuVvtOTiWeyO5Q8hSXow5KEAH+vgUt8IuPAY
zUGLIDqrCgxYbrDEuS84nsAGObGb6N4w/01VqgAZaY8Ii45bzuntb0wyEwFiRmaozlo6A8+xsYMC
Tl1aJP9az7Tf+zmz7V5zbwMVt/oAq9LRAd2HOcLb2YJ4FKO5ejoCiE/VhukgwokOQzH6HocXJNLc
dKMrF733oQ78evKpORyAHoGlarZgStfofhsEE0kIFmbZpxBI1LyX/ttJHeQb7e5qVh3+h/8qaWHZ
SZXp66hUflYwfWH5HxpioiQJNFGQF/mNHhyl7Bul0uSXp/YdCfxJ8z7i5k0zEKjQA0m41C9XbYxH
LSIcn9ohxjgqO77TccJiBWAzGE2J5DqIf5HKdBBOfrMeKIg5Yr8n1VdwptBK9OhLvE23Ziy10zNI
DtoO/aCbKEcrA96gRwFWUYYOVo3dacyVtUliK663ugWpQSKj/06/AhIP0l6+3YdixY5aFqRSLKsD
fpfHqUqbxMMrufrKdsj9aI7E0fOesk5lW6L6IxaVtbz/zGkVqawUJy8c7x2A0QJWtBrvc/8IHxjW
YcJsgYJ25dCUq/eINd7qTToaZXGKAculdyxc6b4OMasXz5r+s+DeTCrsqSOqhTzSbrruDlY5EBlm
NXmnlsBPC69w6lV815aL/i+a+TKtla+DChbbDLyOI/IqiTpc77rwr99/TlJhRbJoNz0u0SjoI6TW
1y/4Co/Ud1puPSPJcVNXC998Yrv7U5sYOdrtnF8D8rl6WjbNxrM4qk1WTrC9/8Bxkvl4oI6DYTuE
cBT4R7yCuUvVjcNsgcAbONsZXVrYo/+3bnukQTqoKwxyoY+vluIrCZy3fvchsr/S1KhoLoyYQGfk
UjiiQKo7URnhLl5piQ54j63KqmPXuCq780/0ykI34NzI/EQWlQ5PN01kVd2vUAh5hHUWd7eWUpHT
oIK4jmec+7w83IXmu59lhk5aOI76gWj2+61OGPVK12gilDizK1fGFd89zbnrat84+aw0SwfIpnM0
x15iO15SKRxSEuuEqdlDl6DAFrfXzGepsMMuXlD6flE8yGhOSVG8LDWPJ7qiiDQBT3bLcRlIsbDQ
fifqooI5gwpXq0UGW961DK0WY2e5LUV7a7BzmqwvOxHSg/Pvs7V0LtSY/IxqdCzjmjGcqoFbBmAe
rlV4amlMAf2ARBF7uNIMY9pICbC+KULe/AynU60lRBd7crkp5tHOFzlnb02dvq4tWn37L7j/HCoS
tV/Qiv8tFxgIa+sEiU8bna1oKLrqP6s7lKXxbq2gKA4gfi2mgQsEO+oMADK51JAEK2xFX/CUY/VC
yQuA1mr+SZFhkETzHEM6pXu9tqJNybAWuI4X9Z5oa00YRAj+BZiJHIulT7ZOlC4eqL+ryK/ZfM2u
ME5N+bVJ+4VdkHEAORizzwy5ZIe4NluEz/XV5+iE5jvUhI5kc3jmk0a7ewI17MMKDcJEuccDeZb7
Nti0YslvOiSkPwMJnosPCnUpjiBG3mncdI+0aZHVht2gfokTlYxP8TwDvWrpeZbrfJfQ6+pgmoor
XSHh3JrYGvV3g/PFCZnMjeWbpOvkbz6JlckeS+5nNKxg3q2CAvb/hDj6qMJbF249gbQTFxmbJmtP
Ng7eOgPRXp9YWz0bIOBa4sAwgtUXsLhpy1LSIc+ydz/fZ6fN7Koyel77J9kRXnk8+oDdxqDt+X5x
yBS9K9VK1xEaIo45YHt6sUkxPLpyrBfzvWxf6i1GS5z7sWZjF+67sBk4UFBAJP+v9KxmtmpnRdS/
MgvhMLAmQEwSMb+ww77HGm/Faj89hDai8ykgRA9l4eeBoHkmMYzN3Ln7aoypnGf/BB0ShN2lrRyS
RDYteW/IZVnLvPDDNjE30sFBE4YXt5KHqEh4Zc7W135m1CSmWs/+yF6xyuqg9DXKl1Eyk+bVx9Uh
qT6uuhigZ/OIHFlu5W3RAVgYn2r6m5oF4l+IXX8bAAjHkoBMyAkWDIkRtELRO3Ze3EnXOCgbXW14
nbxP1Qg+3+2aW0NHjnATdu4uDOFUKffd3LW3k5HbaSGNarOCsVxF0+6f5kYLt5bDPZHtI9KJw3GQ
kFbeFUJEkTZbEezXStOnUrOii4pZaHBYyA6v30N84WAMpdriIw7DG7QBMGyPrIm38+P8FfgZKkOM
wW5uNZPbzep0XfPyJVBdgHZO0Rmv+0KODDfnTggKdQUbC5MBgF+0pnnxpOPLQR7eaXnXC8opkCxI
ALQt7DbiAZRXj6IOFfuAGv+54VjRb16LgJbNRZpfbJU83/xqCqyjwBJJfu+TiK+d+5+vz9R5sjCa
VvcfyWXx9eT1us65u/+pUYXhKcQehDsXNg2Tip8A8F92FqOHP50M5tdO6URzhVBfXoYbVPHoRaES
DCDJuyjXd9NyEI3BXeC1+PZGhzcRv9nnglRXw/qCZWP9HWHnG5MhJIFyZ66ThqcHBLQqJlrtBfG0
gCi1YIz2lPLwhnu15WgxUinGIemkKbaozaHxPoiOSMRgQXzXlz6Isj7UGQu/p5B6csi3wfy+oDrf
ad/idSzUlIbD4WvhOW9Liy/Co0a80C5v7J61kRDmSTSlaOD8u/pKxYU49AAmjOf2+C8KNOfjAofS
5lmwHnI9ov4dpWuIztb3F+8SHDZn8XEYVoX27TbATgv1PcS3iH0EV7l8TYCDvxHKLRYgyopirTDm
4WwApL+q7ZR9+LMOrpL4Cuhxb/Z5PqpBzqL7yaAzhYdDf77BW7PFVGA+KlxHDDHbLDZ1b5U9oYnK
eF3AteNAuZJaz86H+J4GpiV8HVIzpkutH3DniGosrng6DMSNViUaObYpVpTrovMnAeMf2TdDVg4o
OyooaJ1pcgVvT9yK4x+PRDqFr5Tx1ajZo60iadizqyBPChNmrObEtopfx83hGXiefLgdHTMYhwLs
kEx2EARW0q/pTEUL1NZymiEfZbvTyzZZKquI+J/JdgKLyhiDxlAjQnHK4UoTMUQhbiWSRe4VYP/a
Gw8NiCEMtAOod8r7WHu75MwWL3ng0ST3nblqwNDiA8BKYFvwkGmgWwHMSgRRcutsE+4zYs5vq8H9
Fk+j5pM1T2W2xc4enCKRcad2QMQTUiY1dLcCYgKAUpxUZfG2jrJSPM0ymDYffYLmAe0Mz1XNf/i4
UCisSDRmYFX1kb3JAAz9CTMXv7+uugBrBvtmk/1z3gWrO4hFmrwD0eqIR0S3WA7zrPyjJSYWEKTZ
y4TtGoyjS2v81tfzMMGPakGHKjv5HiIV7sNgVpVUWMLx9gOLBVkA8C3uoYe8yhyQxmzNSyAST7g3
l+1GeMrIUWRpNstbYTJHIf3xOaFTPVfpeYl1FZGOExH9drU67skK2zbJkMyATIwQKXtFGI45iy1w
SnVMbDsBkFU++1cITQzL8etCfGf2mWOgC6hPgYe6tZ0iVcIKQHJk4Y/sFcvhL6CB+7mp51xWXXkD
msYN3UKDu1B+zd7fD/fUIUM5PMB1cDLqG4sGEcMvVD+1ZqT8jMf+6IYuUCepFkyeliTJJ6fGghr6
vm7QEusp0HDbmYp/qhazNxIRwUXgnggk24Gi/Vi4l5Ys4tFEObelGS38utBl7lku35utOoF48qyC
CGsbZQrtGsctSTNYM+sVkzJ3x9rLI5yhYSY33F9IfS/iQ0GFOizS/u2PZcQJYHj3Zx5y1Ypqy0u+
KHpht55+6K9u2AF0qZHwCT4ObXvUjkluv+T65nj36HnS/OY42M7v8/GlEbTwNpkJ8nQ9kPBRkfG4
4EcTPsOWwMXh58Ix2PYb6hfPYU0yA/2oVhtbVSjrQj7hKop1JDsrI3r2T3H5gHr5bgvrJSP96BwK
m3BA3TwJH7i82SGI+Zykx5VVrshndK2S7luQ5v4pbZeE5sxdftS6EPYVYN10zSRNe/o4Pym560Ut
KGT4z3q5EvCMjU+j/M6tvzGvXi3NC0tOTeGFtJkiBmHaGchnAiBLtRXSDbVoqNFoOaPDW3wVdnUP
2gxCJtLmUeeHE0WGEBReLNhInbpAT6NpMwpuq4cGitJI7NyCYgT0OSZUGu951LeI8uxyTt+DWmsu
SdA41vFPj9O843nNIYG8pbNWH+C2wJvQh4h0AdK4gV97/Xf8zr3OH94mwktJ2OOGUKj2/hdWafbE
TFL8PT0SkrfUHBwiqYUDeH8/U9mlXMl6HXzDU19nE8ZCKIBiTf71guLZuuQx8QrtAtYpSTFH8a/R
t6C1zUZIWWM4FvfNDtlkfOF+xXEAlKVklDUBHCBRGyxYyiFb1aTnTGxQ6F+snWiCcg5v9eAdmucK
RnApNOrYWUYQi/89c9CmQc9WOxMl+9I13/nxQBYf4p0dpc/+Wo8Z961dIYNuV2ABwaIC1sCtE6Ku
SdQjXaGXmdTV5YDBXxc9qrD146p6cIpADosNhPB2hOZ1NeWGw5hIdzF+BzeyrXv+8lDXKg9R/qjy
KbZxTSxfFztWQuR7uMeyRtx/fQ6Oju84GYTVo0eXXj8b2GpbEzb1rvXJ8ZLgNJVtWVl3cErDAasi
7Whh92yxhMO8dJPlSUZjFTIB/B3EDigi9DYeeSdV6aYSefkFlRMc+69io2/7uKW/o0kbSmYc+EVj
VxdVpduH7cH6inDFNyjKQsRLt4uTpdQduE4XczbP74kt8nTSg7d5erDKAjnDNAsplnfyB00698ib
pbqxqzV1h9z59oZfxW7Rdc1O0MnKCkWmv59gvxedW7xwZhcanfL7z/bayk/McJxstigIhcaMjzGk
6sCGf2n58ujrHtCp9bpwQC8o72JxgFBWbURK64jYCfMz0t1yMAtZ2TyPJBRXsrbJVe8E56/JeGDE
R7QAf/pQSylnfwV8h2LPAcfqpR2EgZEAjgieDZDUuKw+wTtkA7cSAOw9Jn4XXinsgxMSjCP0NsXr
H5ClagqZMT9Oj0eWi5C4gQLLAPf4VWXxp8EEyPbJS2Z2MIVYR4QTxrAtZXSadLcOl/mL/D4zes7u
HgeBeW3potL+f3hBCo7i7NAWw89lEM9AT/KjHWIpSnWX3Q90Br+3f1+gfJBNbHiwSGFYSx5vIjES
IUQnt/cuZrfvDdkbbOyuXYJZ89f1TN95et7huSVUVyWaPPcGaCeHUxludWCj5GCfkde2QjUGqShq
a7wiunh2NBODyRhOG/cvdjAm9GPfbNXDEZsQa2k3tmlBHXzMAXxTv0h68M4ZmEkxeyHT86amXuli
mBShiHGwpQOtxLF9TR/LXKusZg4G9t3SXnOYrLse9xs3eyf+tI655RfDN8LEm9v6LZRSgPyt4SpD
MUyhjTue/4b4zwBe6iAebbGXwSUA8416uCWR8NI19qHOWnYFUSCvJs63wfpAC4tpbPkedLJA4hHE
+4FiBeuyKHOAzARCicBiG9nIt5aCmUUqqrbfCCMwvYxoFqZZPjIc0X5qj1C+Rnj8Y1I7aJaFw3mI
Wraoi/C9bUgXwrwq2MT5y5CKzFUgsag2uQERVGEm9YeBl7UPOkh8UrxabZkmsWdsiGyAd/ceTgp2
DpD+NyUu4aXQlJL89nhcrSj4LlCxD3BForMhG20z/tSIjzLj7HDR2ejv3075F5lwutsOMgKWiCbk
Ir9d5ozVwuFYS2xNVJomou4vocCszQqkT4CfftGuIt7IJoMzG6BUSbyWVirly9rfCpc1mmVRl+FF
p7w+Vw9Hhw7rsaBOf4iYdFB3dzF2ugOHBiMsr7PXACcVZKywqZZvSJxCnbPT+37Z2jWowBt55j4Y
yPMm3elg0Cnegvt3z4Xd03pnXOpB6CeW/pzPOaJkvyFd9L2ca03ElR9eKajwhO9WyA0oqIFO7FIo
7iT18AkRcvT3Mycq3hLtvtY7/WvVMzE4SiBqo+d2yZyCE/fzyiDVzWoEQglBW9WFEtffgzzvgCuY
vMe5jcurqRMVAuV15kLokhnLoXmZBXQ3g6ZhujQ4kfajmumOPy7JqJ5J2B3fD5qckmgxmgLJXCPw
HKaWR7x1uhUzQIvh6l5ae5TmRz9asnlbwNKxEmGrsViN57S+4+b8lUBYZw7Qh9iAMoPDVRbsXvXF
aFntVQ4Dd/GGcPab3g6mbhFkn778vYWY2RLTAIMSyDVGm2APCxA2wv7ZTP1+dDrJ8RLOLfuVUO5+
qoW4ORRiye4zoOTMdkv90iAhg2X6FapKAxmtFgOrdmcaZUXalqbw9oGO9gPQU45vYAzIeE4EpOkw
L33SanCoQgrZmHJLBWS32/16rPv79Zf4SdF2bQveZB4D78fiWhgIAUTKBPbFPNBWrMCmd2NrPut8
46jEMbQ3vTEb+qPAs64lRqlrddjX/ag5rz5lL3KiB6zJ/U9uOXTGrXZzrT0sHTXPJqHz02XAuK4D
ky0U4nsrEjDbpg7B1YKC/d13j/Q/ZxlQKJhvDwXF2BQzNBio9zoGInJLSlwrthyq0SQIKD7f2qKj
3nd9baxB39fr1WpI7LfnwnEIbVdAM5Nitdmluc3UCcbToBW+bL4FszGeZwxSvfvQ4PRMzz7NtWXG
ryX2jBAiCPiwhqw/mrm2rE4iAwG2YsUFHDttpp/A8vZlgkWaYjnCu/sfrwUK3PtuUmrMeu0sKMZc
CVvjWBNVnqn0bjo6Gb8qboH7av9F5baMNELawXiMUrK2oK2VPiatwkYAwgds0wi4IfMG5zPaL8WP
r+ZYiSg5DrX89jMzy23zVy0fw7tq/mCa4yZV/f9Nadi1u+/as/21xZzeea0BVv5/XS3kfccS4RUd
2FtzEsLjCqoIdrru1pB1qzrIM03bYVOaqyMErdeyEZ20ty2WIp+RhNR75+Fn0JqE64jpPEwveZW+
jmiITR40YAMdXXVU0rspDyEDMS2Qj1yiaRu5keIENi66HbwzrexTJcL+Vww/tUoBoVomCNwPAZUJ
OtNVNRioAXgKSn4aE7WNd9yBJHcosfsgkzoYiJCROwRqj35KIP43013tWqiHhcxbXqrrja/wHlYy
APUqenP7twO/iDhaY+FzO7YkFwlrUZQ17uzeDcVVJVmALJqJPH+iSEXB2Hq/7EQ+asHYFQuflQgs
lFzs1/+2q1Cto9oNz5dgXFo2nL7FJAx3usiMkeCBuNNaZIyALUL+1GEI++mEx4gOkYW7VIRaVjXP
bXb62bO12vnsy6m7tPiI7GwA7nCkGoT0REa9gm4Jqf6pCD1FfxZtKfTvC/XM5OvfrRLAlXqgc6ev
pLXgbZDOzEnaWjx4LfTTh0EGxEVktmJ0QvxVUvOExhcy/LV9vW7SPYYDU9x2V/Fh3S9QfdMxJq2T
AGX44NowWua0kl/9jn5Chk+VjgarHErSzkRLIA5ygRMeQ6dkGU4hEkOtDJ+4s9C8acD/oTcBS+Ue
7t8CoKAtIRCLqo0gVqVyvzHv9CI1hC/o2n4Ydd1QSZvcgptfJh6i9AaULHaCSI6vQy5hdlSir6Ps
hLfCkCzFu3GQEKbjAgV7VdtcJWYOY6a6wszcvU9OeGRx1+pit6PkIPgEPux3OKXfOurkQbXhYeLB
S3GJruagVtUTWfcKxgCpUvfRn2J7w6zcjC3UYayEhhY1tiobAISR2silhr0/LWCPT8V/pDO281sE
C3w5vo0A9jyysKhA9jGEn2sZmbe0OnhMDxHwoapfli+rPRc1kHoJn2KEgbM3P18DhCjyc89wvfxe
n6uKNRflkpM5JrHfWU9L8dZMCmKWcCymPmInhRlDr93ypRXzmYkaF6D7lxw1Ooq6UyGXRjx37eEh
CSHDIHRQIaVAxjbUJ7QQL5nw1lPS2+aqxW9OjsNcyyUGdCDJk06UDrEcspSNkS0lrUakLuyry7zK
aDDmJhu/lGPDiWCFRIiXqPf0BxMsdKNfSxnGbsSvKuhNoaclt9vJ0ooTuUJyX0nKHWzV8tl4WpFo
S9FSDf29EYSIpfsVZ7qJKqnmqI4bAMs7b0NMR+sJOxJ3j6VbrWJ+911/gM8RSnAc6Nwhz0PEbbWL
nMWXRrLTu0HQ2Sohlbcd134nYiluxt0cmHsmcCPycYGfPC2lli/d5AcT9iWK0re22Yu4k7f6mZAh
IFkziDJCVFYRwR4JbpwFZOTzYrVBrPTToYsn1USz11wmvLKVKjv2CkHmYsdIdx/4c0vq2UvFtaf8
Yyas/gR1oyD1VrDWrYY0HlKP+nKlvsasst7HTR9UmFADoR37a5cqaAsLFzSR70inCOyRd+ZzTuy4
tcVFyBYIlzmJslrLd42GnCvh/nR84gXXfItZ7ZjXtI5orq0Catc8dllKahVrhuDMDSzlhwT/mGZ/
Kqvw6J2B4j21R+ARYNVtlJkQ72r5d1xiEwoXxXNlCgqhed+E73KtEM55bZAhM7qOccBvGKjfPwZ8
zGaRjpL2nlniRP0BVcvY5y3e8kpmcuRIj6z4s79N5qV1o7FeDp1iI/sQ2tfjR8AV0TUg24TjXhfW
CNlMJtBW+gNXBKzRvOoyp/pgEIPya8F+gpDcAvNX7Ic5d8pPfoDh+nj1PLc6ze1sKpyNr3HIjM+q
Bpol6lg4GM8mztxmE1m6Z/3EXhzBbh4UQgjj+++VavVQ/+1Ex0ll4IeJggdV24Rq/RVt3ndOY6Ek
2PdrVoF6fU1OQD4tTwRqyfLfLQJ95fWPyMzb2NFS/rS+RN/lm4CoWaNP2PJ1UAwrCdZsyL6Bj1BX
fiw90VyJLPA/p2Zja0FpuvNqIFL7sn42ydXxd/YROUovRHjw0m0LmkOqll7e3ryrUA9Exfazcujo
qLLtyw984RDbGBtfuVc+IlNWc2SZR+TTBcWqfloI5qgbI6FIH6rCa8QQzO5p/ar7Swn1/ZfEWs6F
tYghPY9sTDUlYGlJkQJxNPgyquopdpJRdHOsz5oFzLgqRYDlTn4zIPVWXDM75p361BeCOXT8tZnS
RwK5dZSjCIEPY0MeIIvJJ1K1j+uMv7hLZaDPBXJNmPU/ehXTYY+vCsvoKCCFsLTyPYRngw10ZTId
0SKb45rUOkH5vVnxgZ/3ECI5vYcYvwi0bnbBwEQsACdp/+FDyy7QmJuSO5dCthRCiIe73kCiLWd6
FJIO/yi4t55Bo+uuw3z/RUQYHgfef1HP/KqPO4zn0htioBczWD5tZXBJwjGQ+aBw+r7+8YcMx5JY
1FB5sSxe1naBhnMg0j9OHpzlFe5fObPvF8XQu8JpVCQYtoQB7dGPQN1W/q5w4f9DOfeA+tDcfcf+
WoEHjzRcFDN9PFDYjVxR9e76PIaOFcIP33TTKckTUpvwGjsrmF49FG1NiQj0CvaanCGSkMySqnQ4
LJlPMWy3iA81CuOJftPQ/Dxso5FC2sNSNfEZx7vwPQO4gPAUSHmTqFU7BSRY61aSTeoOY0T7YZ1C
y8ldcpXjS0X/jMtev6ealXdYAoXccHTWsxbv20LMxTvnPvlwawsWAkifjs9vETHwLrUOH8ul4lpr
4OruKqykfTmdyX+mN6sgUKCR/4HOCalTqQRiHC7dWOt+/yKnYvb9fxOH41wNJjza0Q/fybVOzXdg
7q1ZZI8Dlc0KDLBv6xPyStFf3+mg4BJO1n5ILvizrm43QPmD2AEVuDYktwRpGD7yu3uvjjwXAcJi
sLFjcs6L+SrWMSez6cuWj0Jc/+LIs4K/WXpOuhCOPapQ8JeqcgvzEq9iWu9i8yrzjoA5GFsHdh2X
rPRh/ddhE+RSSaNsMF7LMzhGfjDW3jOFTEzg11/Zx8pS3uWWiV5fkFpa3PvmiQWL/ZmjseukROfc
xASu1GxM6MHkEZPvTZT1HRzbD42B4tiFFApYk1guDWcBQpexE0sOCEPl/3rNJkyktDbKslPOc8Op
k6zfZHwREpUZtFpP/dsSioBfTNQkTkW+0Wpi66NSCY76JY0MtSy7zDhNgkfVZTwMEPcyp0FFyMrC
I72xJt6xLRfaRAR86z9eRmQ9aUQcF7tqCYHWDS6vqAS/FQ/PjXtbXP02KUUKdANx0M8TdvAcqZ4r
rGxA/SBRIM9NEMpCHazHFbmbMsYHSw4oqOjWWTjbEF7hivPI1PIr1S1KGLQY+EgOnGgPpaZpRvou
ciywvPQT78MoXuGEA9Cw+fPq3lfADCx4+fkG+PK+FtBIOOomiCZEisgUhgGfstY+1uTBV0EzijRw
J3tP2JFhDKtE6Duym/LmhLsrmls3/YmXN16kXzHk+jBq6oNWGq4pEetqO1UmnygYl0a2u0zxLPCe
x+sq96ihS+tf5xMGQaz5aGvHRArH6lwDxhmxYoioWFyg9fFu+qs9FdEK1IT5fwKIST4eItO1PK0U
2w0Qg1kmv5QvmO5ea5swbb5HhzIBJzuxmR9DCG6/c4NPU5+EM90BHgoJzXctdwvZk53H7KzGeqlb
ksWEoR+fUXDr5fuloBznn+X9bClkWdERdvIqMkIJi029I0FAvyfA8PLMEZbFKZNWHyoVocLKz/W6
Efj7K24aebV+ZVred9DeVOH8OqjsagHM2YPfd/c4BZ4UWjL450lvUbnSKAbBLK2k2YeIiCSWZbEn
i9mDGDTibJ+DsPc+t0LNIkvj/2RKOE02RyoBGDRoueEEPG3bCI+mKNuFFvEXKpzW66nhhaSp79ms
xT3dMK1C2xUJXTdGUVHh6aXT/2CWo1Qv/6VreIEnMt/1Fs+ZPVKhmCrKPcFLWBRbQ5K4p3qd2urI
ec82M0j4FMNT+LMCzINtZ/jsf27C/d0AaaXwzBpqOHojso/T+GV/NgY/w2AZ9rMQ6OWvKAkv9y/N
ZRrkMToWSFlz9SWEOhB14Y5YdXEpiyEcgT17cX8FI8vYEE1oaIYRpproCFFSVqAPsOu3Nn7pcaFy
Fg1ngoBuvqiMLCTOxN/vZ3408SQXtpuPYtTa7xLLN0MxtCmmXXrVDhMumI17nkhqutegCxnPLWrv
PuyT5L7MEfuQI0Tlbcd9uKXXV5PABr81IhQfvfgJpsV2UZa5ePMq28GdaErKzcrBNoK0NfsbtROy
7gvLOYS5yhy7FZFSZCLDhCixU5BUMbaidPfSKq7KYUwIGITWuhN63h4nIBOuRyDF7nzARR6LiQNX
Yv62SXJEDm9/u2jBhEXCSBRl+PTqs2EzTD7zlT7KXAB/sqWHIPPUNx9GCWwUvIDLUcoIvhT77+/y
JZPCIsAu+RLjA+p6YtqLfZ9+6Jgma35LW9xL1FJI80ez4EwOLNTCnwdmr+pbPFF9wTDKAtByKb5P
1FqbfUq2N+3BgMKuErlwiRL1ypZIq+ZmMv9qq9b6HUGQTzLwN24j+GlI/UsqjfatW8gFj5CsscQR
fVUAWgqmFOAblBdBMVv4rY3NKrb9ozli2OF2NUYQ6SfUzPkxxwLrOdXZJ5ZI2s9C4y8KRZ80KXyL
rP4wvqUSXk+jHWmqBig6dDgRcgB0Oxq9nKrt9+olreKMvZ83mS4KYJmO/8fDnu022ocF45x3Dce9
Top5jR+nkgYhxTpQH7IbqTuQlqc+gE3nAe+m+cWv8obD/xHUMMX5McVPVrnACJXtAWOiR6Qond7s
bu0rNS1qmFUZ6CcsDNT7CHtPQgDiP30IXF7yp6M4bi+7fCGdH0Hi3ys+rpkcD73OVe44VlOdeALJ
dDXVeCvYfTPm2TsD3O3gM1NR7w4Hiv2Qd309duozwNebjWb9nxdDqRdyO8d6Yy/8FmNrnrdvjVoH
tQPrBzNHGSWwZa4v7EaI1xWAqIRgfS3fcYho/4TmYg0gtAVERDbXbPRfebsJzFYLeYikm65rLZze
REKJQJE4mh3A/gxOWw0frnlHGF+pJNHZdhwuXssqgGfQ1AUujnqE0mu7w1JwetY5GhpB3MAhNm2O
fm2QUlFh4HjNDFI+DUKMWAYmkugyaQTjq2QVMLLvvM3mQ2APRrZzBX5RQhDpy5on68ls/+VowP+z
/2/V212DITcBjhkxAStKBcvWlP6CJCitVvgw5+YEsl7DN1OwdSWFkaj3WkaeycOKx6PIz98pNCoF
/ravq6DE9U/XDR6gWxYM81Fsy5cSE52rdAoi5lwbbh+KS8cwGvlHEmYjjh2ScprV2hXoTBeX3w9r
2cd3eobmlUSs4mj1GdEuKrAIC76xXiT6tIc0HTzGhpMo8VQY+hZv4XNlZQjlKL2KpPoVxw03RVoJ
G8s3g5awJtZ8HGIOFI939FVDDxyB1xQ9sHX/iVgOCaTfx8kAIXbfXjXTDdsX0rkYEI4jVG+WGLmG
+RbENZSuwPIrfzNHqsVNXYxwpM8NgSB2zun5u1/R4aEukDqhIcFkq48YVWOcmtD4m0U9eSiFPYPR
FEB7nHfxaXELWo20eHGOrvZENTTGdWONuDTWK9cjVl45XfBJ9TDUBLxmHNEXhcaHxAG1HMOEqLIG
zBJn7R/G7j1DNVtMxJeN2fe2zDWIZKjHxOua42zxszbb5WES85Ac7NS7ERF08ydY4/NeauzT1mSZ
cM2UDKre3ulwuVlCs6zWk2Qs+jBRW8f329C88rJ35PTY62TEy8sy/whYCcPLecpKsc4uA32EZT6k
EHOjUraABfahEO1P6Wf66ZprS3prnC0ToEHTIDy2zUP62793DHZm8pYCZ3Kfl184LtkQZMFetGdr
ugTd9gZy15TzBFac2o51gCLynxcz/BJZJSCoSxdpdmueK6YHBQed0WMobOS+lw2qZiSbI4bG6HFL
/s6V4qJVt12qabaHOj+Vae4KSZEKUN+luxpER0rWqJxj0jTWZzimaxMWH/kK05WjZW3Fe7Hv4X5c
EB/oKVK5VJhedKKxstMzlhTpL3T9ATLLebgeg/D1kcQ35/LAtKCoBUHHaJEL9YoeFCvsFTIbjst8
WVcoYdF0+3BBa12FZroLS1WnzkCeIQ3Pv5r9CI1MHJsyTl4I7koPHFpeolvyEjZXKQs7bAuOcwD7
F1v0HxOyQxRQpexQtXpeYiJ08u5DpUmsnWLHPg2DnGXAcOj+0FZEWwM7Aw7glezMsNzpAG1XWgfF
A5MZ+BBURHv6X7MxqEv8gMnxDbxT8mdziYg4wKn7zqKlZ2P1SXl8yA5D6gBvwP2K3mwezLz/2p/c
nyXooT7Pdzymt8yYyJ2PG0Acanev5yV15AMoiVxgrU9PFMZ81d//6CsnP0mV0RuaqtIPVoG9/l6m
KUMzlSQopArkc5XfdpEKqjW1cI0LptEhTNzZmGFACA+NhQFzP6oZUbyk400mcKMmssl5InrC7CT4
4dyy03WtBDxY6oesviYHbHyKw1ziVSfXJPJVRhJzTNIHIHoy44TBJWYzM051nVgXfteAqMIYwuk8
mBYi7g6BDM+B+zYTdv5WhrOyOjZ7sj33GgRa9pfW2Em0z65BhuRrEL1DCUxpXZMQLNqhyB3mQGCH
rcM58mNA/rFtP8nZkUW7BLHXrSUw0UOg3d8H7B/OIQLw47b3d+7c91PDXjjgXizym5uNgiHOsibq
vFQ09GkPj00UuWinChhW4WH7yh92zdJybLup+BBpiFydsaZOqKXTGkf9O0IX+Pcm+06GnXtzr9IU
7EEZw+6hBQGCDPndbLtU1DMGmCRL/RSH7Pi49/Um0RQWBGMEZkUrHAj/myO5MPGDXJfQaWJTUQNn
XE77kvUKbS3ByHxj5d9AM9RTLxCo70jfhyMWOdiMEaB2eHbklUeP05Ai5FOQhgzMijxvmV8O/DCX
/jHbYvxstArHw2Qq9/8EwNNHKTgC4Vn0Qs9paDgEIH0djAU9fxD4exhu1y56Nh7yytbG5BQJdZWa
oOWkvm2BQZuGYk37OFotuLQMZe/E5lkOXbFnDlzAiaiwZ+pxHDixDi1IYiIap+BFjQgtskEBm+iC
Zh1uZ+QLT97eKpHEV60Je1dpdAxDtkKhwjpelCPWlZpU2qQVfC0Dcs9m0GmLYVSfG9BMhOqL+2+m
WWcBvVXrYHFzD9F4KkSm9kJaZNghrkD9UMgPwGU3rtYa1oifyl117FPfqYACMithi3sNe/T3TFLx
DEG64CxFCA3gouoDlJNNWNqVFJSM1gKetsa76dsC9x7E0SQ/o0DW7LtVOxDXwBcTsKbDyWuHqLQg
TWPHi4lI7naaFqD5M86QENO0trXapO9U/rPiZM1N8n2F3Zc3YLvqag6WkuZINYnFrg2BMRQtywzi
vU4FsV5lejwxCLRqZroieJ4EZ8ip+qbEyqkdy5406+OFKLKNbo1JWLngWH9sSCC2w69hlUjwQpfE
frXN8ptLfQr7TOV7YjX3qKrs5QP0vgzfZFPaMhitBqf78xgKejiWA8wigpfIZVvKBbl/0bWVsmmQ
zDCrHb/Lx1v5voV8DtEMrulE+UBCFm9SiPhRstWj9F9AzibM+vvPffXeCAeLXyCby7PzwLFpsr14
sFAO0XN3zr8j4AizKBbpSixqBW0YtUZ/ufypYAzGPaYUtD345HgpUK3MsSNkxUyuFVSUtitXzIIW
qYoYfV74kQjs1UEpqAuW5a7pZU859LZGOfmS0MC21tOctvuNj020yYmjSCuccuZ5iwJkhUrrWdGF
p9gZR9SkB5jQHjqqppivi1FRMMtVt/m+3qw9WsDIQVvzr92S7DPWGhSnRepd9Uz63FJpcacGVAtL
I7RropcMZpkLXCEJtymHQ6RWowRDzZdeKwQqOwv7ylaa7b7qkpo4VwhxiStPSck14Z91ozPm/o+C
trp6KGwcrinmKUeqKKKoCn6qbMkXwBCNxPH4pi/aB0dZzHmt0iFE6H0aCd+IwAD2EYFrdYZpiWn3
/m8u1uozUaW0/9v/tEbe9S/1tKV/2Elu82QSNdGwQ7nMhL9Q8IAsXKChkJYhXOEs+XNsZMVYNIhN
8UDtMktUEZHaAtBHCPjQQwAX44bazsbsoTPaKnOPL95ZTxttfNdGP5CO1pE5H7HF/3s3u/Ptf7GS
OPvlL7MxqPAv3h98td53SCBHJVNWV09/BJbRUtXqz7xdcYmz1wXp9rnRn1GNQ/U0DZ7vvo+LxqIB
xizoFqxqWX17t9J/HaOXJ2AAn6bNq8iLOVgd4odRmlTWCaYAlEHk17OJrJpwcmO7iZ62thJUQv70
yjO5EJiu0EOFJ55F/z+HtZX9XbMJYaeBBqWKD2XGtqreYTUarQ5aFzHPzL7AQFYMTcyVxR0VIv92
d4+etfLzva6avjusYRzdYYox+Jks7q/Bah5BSny6YuFfyY6tRYaBaBcP2kVTbDFvD/8k113RYV0f
Bg/qssN6UgLQAcGsCVaq1X3GlQre03Yb/ILQdqaki9QgrpCdllXzm6fUF5a/o1m4U1BfRFR4CN57
zwUyx7MsXIjNdc+lzR8PaAr19NiWyiuEGRM5jppfDvdokIauk+7SNR0AwTXr0ybSO3uAmuujSese
ARXYqt570uY5f2xqsDkLPYg/DDIxByy/bYchlFiznGT2Pnq+4ve2eccQ9Y9my6Lx4QQl8RVhSKKd
krATfxExMZVfXERxFfKHS9tglAuH47WNrbiFWxtdrJctgBYZ0p56LDZKxeZVBiInylhpytyX0+gy
XbT3ieWnciPNhRETRHOCUb9LZnz0WNWMzFop9Dz7w6tEXO/hCrCGmJ87ZuqM4dt/bT8NAKs43eCx
Kcqu8x9kG/6xM15sq0JpCPZDPDb/gm06DgAiHDmrUCXaIEwdFxiNj8C1IXGq74FOpjyw8tAJ/laY
xDOfcWoL+kDHPtbwaVqYT2x1FS7FTlQhQRZVrjsL2TpW35jNvPSNuDQMMDALfm7jDnRdoFc49F6Z
wqdn8K9x5WURBOPJKc+T9yZVP5W1JhWkR+i8lgMZl44Ip5BMFOh6NoByDpkjHOTBl9y46IHxMiOL
Dq/10tE8v+v4//ZcmjRHkzwkaMDjyp1UmAU6YJ+sCJYP+pI98rV6ZoR/KXszJ5FNLud6KmgKWsN4
+9P7tJlbhxYIhBujeJTGu1wC2qogxgKT5GVsH8y5JSnAnbjBHAGwKr2gfwbJ5y/6sHYCOqgxnyhG
44aeyYtQkq4xlZsw5YiK6Q8qmur12GRcQqn44ezv4Yv5qM7mL5m7GxLDxXgAOLPmzsCgnvTdd89L
/rsxLDNMnSH0J4Goh9kL+HX9HdomdTGByPz8EWATBmH8C+C7DDgAyvtpMoIlkb59jIdjxF+rnzHS
GofoVzDG9+KtSekC8vtP+FgmY2DhXhtYYlA4yc5mrnNgh8sg9Cd0sBsim3IRV/KoufcRyGdLakJL
U/0z4ETKgWaZkdZf8svVkbZlfUGj8q0rkp5slqwybolKTA5okQfHLsSx+WsOVN1F0c/puDrpnD5F
TJliHkiyB7x2uzpMdtgnCwKa0VZA0iibwB4dfZvqOkUDUOCPeNndqaPxajPZCQ8dnoaPP16Ft0Ss
JgJHe06tfq576c0QeI/bqYFsGbKCV/rxpquA7CsGF66InXA+tblpVOWfcelZS3TkPtmbmtjH+cEW
A0HsTmDm2xLuDUtIUdSA1xI1dCdejcoag7zyqMxqv8/jrdwavf9stQbdmLXCmWKhW64yYteQhgRD
DadL8DlT1kqe2QhZYoVT0cXYu279Y+MYzgSkgikO1lyKANIspMfDSsmaQN0ecofZR3Bps78oH1o3
H37GvzNxX8GJgTDuSj8iQ1ezxeP9FqoPxuf7AlG0FLCYAMAIYKy0rE3AycQ8vmstc6YHreML29ox
4g6ujhNNlqruVnuQSHSArkqU0wwUuvqDQHs8rSGHYioBw6okUU0uGrFTqFk0uA8kOp2JVP3x6eEI
pjemxWubfKO+kuyLfFW6ngyv9WCBaSXgfYRMsy4FDfr4f/0kLGJipRQNGVOiZWULqbVH0svc2SBs
tyBB3ljquz6MsNZjp+nOOtuJ0qrL7ilUMrojj1SMFO1SL32XKkOMpAgPT2UklYn/ZCtuOpj+kcWT
KBJgBRHhFTBf0XzMx/RKbo9LD3bB2x04jS/nxIAO6ZY8hsuqPauEWjvIFTUKynnuMUhxrBNw8uM3
4hJs80hLFpidiMWJU9Twcw3GwStKrSjBvM6FtsHEcBfvBtNZJgOioNqLSdVroVReXGIyBYFxnFvM
41gWHNS40AOzdfNmfUho3nNRBrqM3IfYvi/Os/5PpOiJ9zxnpJoDuOAD4Z0NfcOqFC6hHhUuWOG3
Guo+qDa52+WICdywabWqlOKzRkKpGw9WjNrCtE5xTenH8oc5udLTxTfJo5qu1VhWvtFvgOhh+158
1DGTqFMShyEFkbFC00fuWpNE4QSz/QByue1042DH3GCiy2mVRKOF0WcBvAkCl42OhDVS26jdH3oK
BqQc5UdczQAZSXEKDaREebdk6O2xueEbv0nG6CsSGluSIkoumvIs23B3CAnicPA3aYdmfjMKJW4Z
ctl70255KJpFIT08pV0dXX4w8q9SSNCCfUB6f6usC89HtqzGs8I2EVM3GJVCut950K09rDvJY41f
w98/qLZO6mElShNvBkTGHIOk4y/HPM0dclbrZBRxD8ob7FoSz18ljSyuSO+54bHs02AehYD97hlr
jl98WJYCvlH1FgfgDUM8G81Ij9fZ/rFbitJc+I26bgwlJ1+bjZjHJccIq8cjCuMukcjXakhYEg34
FYLfDgrcIRdqmrXYJjCmlQDNuPqFXAxNQOTsEMi9RpCaF87XUVfJar0Po8ABLeS38f/C1ZaJ7ixU
l/Qg/l7W4j3m8w8wviC7uEPv4MAnWSkFHVKtznJeCU2FuIAvlH/wCL4v/G2umZRLojrZLbsDjb0w
UkpByZcLQBnY16mzpK46r8256Vqsen8jEv1mDOeBBMviQXKah7h6QzlXUat7IuEsK88KlylAsyyc
LwQI7m+ertpYgHpuGFyD83nbsuJ5l3loldauFaEUh2esPVO6JgKj5w4azTofIZCK5NtxFj+i3wJh
Vd433+/dA1TkM1jUhettzhvQVEUiZQhHvtdQHsku7kOzCnSgskJ7l1XejGZAgmzmEAs9bQf1VNnF
j1x+Aof9KOhIvtqFn3TI9jkaDHsiOwaK+hF+wrH02aCPvAYtf8JqUeMN74fiFXY+yjJKAFw6fDIt
jShwbuBnDlEC1k9l4HI1PKKYi8usN/tR3ejVDbdUs7enH2HEBy098cht/x4NqtGOQKvgdVtxf8HT
T9Kg2pfwQ9GS3BXq3zemutms39lwnMxhGcpKtMF0S2f2mMAe2a5Av4epUamo4Yi40kcTO+0gvs4X
ZhYqPSMuXEriXCJEQecnNQG9NpsqQJWcFEi8W/aSbdDl67Ov0slWvpEpH5gB32C7jDzboQ1YVs3C
Wk7GGQrr3cdE7X9q3lPrAMfE3VSTh/yi5vW63xQ1XcOGVgjQCKq8uLVCVOc3NE//ABGLTpZs8Y1y
1PWNP5Nklc+1Q2Y4rO3upComxL6ZZ9VNvwIpImwkG7mNDEgFJzKQK1yGrBKhHLA7m3pLCkNL6XW6
sTWOHQHCPAO9dIq5qRmLwiLB1WgOqYICKNOIvDCdGTmBWm+fToNuNKDdjR4im/bcQLSaTHcAroug
F7ueidvkzuTdYfDwoS7coDyQLASFas0goKfHQ4FkF0FggJuaMLzd3sWgauNbvL/FwU443vnZD6Np
TggewSQ486zhQnWpMrtg9XhReljibWUvlBQjg9TOoYp+vPPLjMiYN5V937dCr3Y9bF5i0VGAzu1y
xOLXh0e6LKWZBt3mPyknZUd4BnqyVd5ni3kVYTKmpnWg+n3aqr5dgJBr3fuXz99z+OwsVXdxyfND
aid9kJSe8EyLbXXy25DjcrK0WN2oAZHxiK//fgUW25oP0D+S2b50vh5ZOlrZAhgZy2OpZSustxxH
iJoxs7qCO5ir0PzOWcddQbNgeSvKD+ruEFKupeiXRvyv2A/a55nNJL0jJXToKxJ//Jf6+OCXrxY/
S52fo2WHUyHxgpEWug0F88T2qREZDsQx/sBMucWGN+iud2b5//xF0AaO7woPaQwa+V4qSbhKBFPi
glv4O+jt5bgnjp8v26gCWTIo2FmZvqV72fUIT+KaRGCETIEUN/mLMAAnxOg/pOMbHmQGQnOoMGPJ
dsE3CF6Tvdws/SF1mhLeZL1r8mXjbDYn2TLUIIj1gazW+XdjjXhVhnt3s1xLEcKtu6AUIWkqwyk3
m7TBO4jCrlR6sfUw9XTMF5ioig8qW6qP9HbLB4Wa/r3NdicX7nxm0YcE04JdKhhEknyp3oKVvVtj
q728RIvrHf2imyXcOVMUK6KT+s944GRPq9TyMduJbOywetB8X9/I4qhjmW4wBgT2oJssxhlxH8UP
dGy7uBRCbb7Rg2giMLqou1gpJ/6xvu61PLTXwt8cxAkgvwgOX5Kj7kcIYrGV3Y22klpUFxD7rMcb
Ity9UKZAxkQCv90XBEMgeq7FoVzWfi3szVT7gVnuGLSpsw5KLj8JN6dzWP05w39vUZemHRo6CPwZ
KrUMpqQJ8fZASBCUDtTluLD1ewudetOEnlKOegLnknUdQIAEru4nTfbs7yt9y4nFugsJWWv99aZp
NTFB8f32hUYQIyFBXtxUx+FLulCCsYdGygcGoiDr61pC9AjCBK+NizQAocgfhgTL1oBpeW+BHJmK
CS7oG60TELU56LRB/nU/LNg9mcg3DKQ9ZCh/9lPqU3ea1pRgpdbiY86p6SrDztyJWHj8HxIIYWvU
Nk7jCniKh4/nT2IaBPoZlCHc9k43IeLmPpm3l2UlbuAT6LK1Y4dvnJgu4h7Vls+NHcRxXNN7XHwq
H85L1nbA79NrdMV6pg440KrTUvcCSyFy8ski2cRv4RUBg89W9ttmvgF+69dzpD5AFvRlCQzFvxVg
vX+pjADKvGnUaOPL+hUWV864I8I9LAzu1PCc1JN8peJ9GCjgrzXux2Pz61O2x7Ic3tifA5GbbYVk
7MUasW22SyG0Qpz/3PyI6wHD6VjjtHjjj6m2pFYxZwNdFqWzsWt8h6Y4xfm8GoYNQB2cvbLypeNb
PRmc4YsXS0+Vf1JsDnzaskso6lzITb7wFFYcmy1HF7U4Y33FQ1MKRtoi/6IEmOg/uVFPBDB8ZsJ1
J/YNxxM4YZtKA+A042FYKAoDgJr00AD1LrPo8jnYB7/+sfthg/IXUC5y1SoRuBGFYR9WR6DT+wxO
cru1yUfDq8fj4YoIosVAC7Nu0sBDwXaqQNfKAD9cAxGetzvN15S4yutDAErPo4jGOUrnYwNtRbVb
PEjV6PJzkoGDCKdEmzvOL5+0xl9vOxGqB302d5GItIhn5wsXhllh7MrDKxnAKz2bcqGOKKghKAeB
U9YHfMTk4jFG9EEdDBZf74yArAPFBbkYrDEgqm6DaszRLLl++eqsTrt8mFvSRa2gF6HP4wY3LGXs
/uVnxaI2cBW6/j1rh6zk2YIPHoLnnSOljf1IJ6lbVUtDHs2W9HR70ZHL7CwP2OBWsjF72aEf27vR
OqRBgb+sqV39+xa8qz0SYipOtS/pjrIXbcsoPJwd7mBTBVNylmZRaKYlTWg4NayFkrcL9natMArZ
PHf1afiEDBDiEc8tpPzf6IOjN63qMhQ1k9DAdl/eDQG4PfL0O7FZPRuMCYtxDNxfO8fVfNdX5Yz1
LIMbjp+Ro0/rvoANRhFKhdpKlsa+/8EQ6/FGFiCTFrv5wyd+8zGxSIuttVW9M+tjeJmu0gQtjt0M
scTiHkNolvwGCaWAPLvPtSnJ/iWoatbTDLjt2+pKehVhyLhrHr16eejx9lrdUgmaYGMGZnqf7WDf
6Fq+sNFjyu/odetiWwNLdKlPh5DUdqd+I3oxogZVLdtWxUXQ4L2v2q5C42ViK4Q3oSofUXdgwKGP
ihC/NNsJQrLOJwcHi3dxEgXj1nmmV1PivTFq1ujgwIZ6lnMe8c4Ne6wFBvzQ5nEa/vq80tL79Vmp
ZH5ZttgvAqRbXE18nP4Z8Omz9mah53WjBX07kiLVL8nXNRN64EdRyOcUrnTwXlPwG4QijjanA3/0
IkLFxDqoPsA2ziBAeN5BDVQlZXaTna6w0i306x2Gpq0Rx0DNc1vpBucifzua9kOGA6GICaIZ153H
bhAwtO3RWzI1oR6NpCdsVd0269Nhev1R6++kmA3DioB7387AyNz5V+UV1xEx1juvrzwbeablKKRY
rg278CzpZott3fjyrnuNLudQdNGcb04COr3QNjpGe0rhfx6YyVtH6OX/SyMbCpOQRr5D8b0A9BBe
5HISOnYh2r4O3+l0x8lGmGz2njMo3TgUVMSJWcUSlm1uqXOnBiFoqIUlqX13r3zMoC83Gsxl6r75
SALaa/o2LD3Gf6UJ364iBhyTPsE0L43R8BZnc5fWB3UZIiJT1XqYemP6TA/OsOFMhroi4dZgvpXG
nWWMoQY8V3bgGQmnPQGkpDBErFNqVRXk6aA0J3OI5rUFDTzHHibd8KMJdNofzjYKg8tZmmBRWeGM
/e2z+JYzEZBO5zMe9EzshNoSOqEovkGLins+vb6A/rv++Mw2mJLghG6R7A5JSfCTpOPq6GjIJfHB
OLoX1X0brKMgSdYlxOY84FR29ywQ9J6EGD9knByxlR0i3+xM4Vrm8lM0sWqaPt7KEOqWq6OahB5r
FgyqcOHhht3pQRO0mlP4/pOj4v3xx2K5maZAQUXXtlp3HP/R/X40i+6UIcA3rmfG+BJYkiA7ZkbR
gmJ0q8sz2a0ADF5tS7jV0hQDXpTGSi9fMT+v7aXjkbxdxco3TwHh/SUFE5or8G3LsANHADxI4iUh
HXNXSsizyH4Lwqb5CUGupmj3q+T4F7r1+AI+gY5lgR/3Had+OvPFRg01EbRABWqv4jIPygjSlHgv
M25SKyA+Z4BtNkKzHZ5yHFyATdi3gEs4J5wY3R1e5XE2vlbi1hDgLYjP+gXO1hr+99Z48c0WSbCb
zwIGwf0gPC/cSVhGn0MzxhKqKWCXfUQYst3Iwzpe3bvCQ/4FsJyIE/JTl5Tsfd2j8Gm/WqaGBvXR
f2QR3bs2drq+IVECHho8xhr0+RjouaU3ounlBnkuVI8Y+p/RkYBmcVkM6kOfOEk3Pq+3qLw03ONt
JdebUBXFdkRYXQvYCPq3FGfWQzSa38ZDtetxjUUyt5dOjtNA80sRy4/2ckrEKz3eTTlw/A8AVCcn
5pwXRV2cB8fUfX41J/DfHk5Kae/okdsD3T888rw/OJldtzegmU9FMhUrzgJl1KcUkEcBkA/ziyJ0
2+H41KtBXvszrBHlngL1j/JYFkWcqfFDRj3LBHlDL12x+D3sPYzCKIcZUPc2oDhSwg4t9XYhR+YZ
Yfpnx/G/bJmJs3NfvKL340YJC2IFtMonqA42a5AoT4RY8QjogBoiG1d3eYSqw+UAlMj629eIBJvd
3LqiN44n8JXsSUvivBeZmUqdv+A/zz5VHQ0KnLYC8uq6rt1jflZcULaUzzQ1s9cHOf0sC+nzHazC
nX2M1hxF/4qsw/2YbavcgwiDqugw775Od77eBg7QgYUNGMyjqeBPHGNheLwOJZcd180EsJemgqNY
lDd2Qjl+4JTozcYHegsHeAmmTHzGCY50AG6KWUNWEye+mNsRlk5YSoeSfZdwgBvvmUNkTUQ0wRVN
qWggW1xADa1pDisjiUpLSwMpCZR25hFHVDepltu+XdogaN6L/K7ZONAbTsVBXI1XCUKou9jvGCEe
k4nJi1sKn9hqDWx3qHK/ie9WtQ5w39CnHP0ULS3a5PjO6KtRoCfGsJCCWEmf9KkuGsKFgMvnyELl
NN6yCe6H7iJ8l4dlkvj1ip7WioTgHzgI86lerHVgeK1IONEp9kJoGDNJvhvKJ7bmdVCaZt2K7W8Q
uW+CzH2zX9QgH99ze8a0YI3OtvPn1/9MJy8Eqm2TJjjtBVRN7Kk7uEP2lEVS5DpfpQ61OvEjeTpj
o6XFiQrmDhsMmG/8WeK/gI2ZTg2L2B5vHp7tr+fqEDW/NNGThNKaCa06EkbZAz/kMTmRAoMl1SrY
snpePU0kfCJkbJ+ntO7nffJQ4PUpOoA6A+tNm2GYVBi0p+kOEbBDtH4/k77McHocZbc+7kOs2uf+
5I8IGDS1xgFqEIwDgbElekvkL9n7DTslddq02GpTAs1l/13DHZNzX6t28jULGXMChm23/BWTZ+ih
JQFhDWxIJcajd4INjB+68g/I5WsBHIhp823XmIMXPBwlqykozrdLS9tOCbbtzcyowbimKXQ6uAHT
jQ2E2dLvQzyUaWTqBvJh1A9RqGKkHQEAucgEXnwTfzHcwysPjt0nfPMJbSaCq3Z4Yj+fKTB8wFLI
c8LVln4WmCAWVxGLqpMDrezKl9MjKqDAkB/VZbvMeQjh0AMcvOi87KJJgyWPYUghcWyjrqXj7m1P
BXOCyNX+7w5Mq+j0F8G0pCYelfoj/XQHOuUf5N8HB8G9RJ+0l2rVM9wFrlHdzH5YqYudrw+Zu1os
okcAVvl0NMX22/NLUSVsrOtUXoax7ErdRgfUXo9BeAGJKBdYz7S19k4b7Qq4YTl1b8BPHZ4hC1Ai
fQvRWYviS3PVfhYtrfP5PYk8MRILo/xUjb9jDAVcJsN0AedaEhGjy9BXbGlsGJSKw39Ozo1GE+b7
WsLrjZT5UecJFeOWlPQDHH7uVupKqqzNbb8LnJNhTaRgebeKK94HNAF8Mae/eKBzTcQvbvckX+va
f+ds2sHahAdRPClIn8oWrH9oZP4bkRyanUlgZD6VXpykk2mNHkUcrBovyg==
`protect end_protected
