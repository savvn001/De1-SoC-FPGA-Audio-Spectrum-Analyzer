-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
noGR3YBTMRrG6p+BnlrmL64s8rSDKkmT8ClMP6wX+iX3N0MecQjbLZhzDpKRU4SXqoZvbIYu9M/U
zdsw0UxzpT1UEQGWa2cW8HKWeBPz9Pp0mEpoKixLdy1giQYbrZJd5D4p8i2jdDqf6AwEkcthlogZ
iEZuzfQOaN8DrqbqF8P9S8SRr+1POM0nk4ksG5iTcv6j9IDZo2qCBwEABCMVJnPLtyH2Izkgrq24
mbe10kXHwoORuOSXXcQd6wGb6p4uszAiSRluaPbQ7BitXVhIS9yE2mj1HHnkyil/TlT8NOzVFXwp
4O6uADZBMzGJEAB4hdVXxaZ/fwjC4V8EV2ANwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
TPZc6hbc9HpE9IBEPosGsi0D4mTy68RD5Sp9Ekieo4DSWOs3rZr+oZ8uuPWR4W7e5MpZNWlWUXZK
5WlIQ3qK524OilzTcc/0f83WXAUU+fweSwfy+5V1R9Zl6cnH7o/cDt8Io+BjWfLvxHjmmbXMal9C
KUwLa6hw/qLf5pOm+mJZWRH1CEIaI3VJTkAF5wRHv7UMWKHnbTaTSJa4qeR0HvhILR/mFQtqNzYo
WKSYo8r72miD1xfbZpDeX5YZ+Yf006DaqbUoa8sxA+3tSVKkZ17PC2HcZE2mmSYq46xPv9yFuQHr
kgQGyTJQFCkvgTdU1upLtS1sUUccOXW72QXmWZXk0Nab3qZhIYNawj82d4fUPwC1NoTKqk65hbw1
PTw7satHdN6Hg3AfNrHrCjEG8TNhuHoi2K275WHvsglXFOtOKW5N6REZslpVEaVckKS+cTJkTR4T
3K3fEYy9JnnVJbjS0aBeNuCT071FIurDwS7vtZLDBT2z+F2Jy3m/Wcyj+LNkc+VQni0YxjFmMWm4
n3lAmgWFEqSWAB5LYAgz1++9L6eUcoFnjzWILfSV1DBb96wHPHGX75pImQis4CBbyJJOYOnuCWgC
Zea/HeFhPPIpGoaQ3fo46FkcpSaFq41vBZQ6BBt0cXfJcD6o3TM8fImYcMRvE7TRhWgWRI7dMqF8
rPAOt6jVG0jCQMvCNtYslc26YOj0Fcz2vbCC5iQjaMOkHgIFLgoyNY2lVy2mTqhWZO4xWpJYML43
U+1uXMGOEE60oJl85MrA9/fYDgFIzf8xiH6UMxYLrk2RHjxBlHw+6cU5fEbI37InLy/Hz9jNRqk/
mTLCsrnnzGmtJHr+SqR8sNqk0X2/XbXj3cOSyDSrU/RrhEeh68ggk1QT/Mjh3ItyXDNTByh/orEg
0Xia6f+tfN40aubfT0TIMZltCMxmGjj3Iv+M08BymK2dAoUrhdnUXO0Hdp2HYO1bS5nfpQN5Bvhz
b/bN4kKQwW0bXgxChiLk94sJBS07144HGSXosrtZ4el3gXdQMQqiB8mqrRWzyOsYhVZfXmPwv/Og
JL/EbBmbLPTGLdMmI48Y6yYuky3q9pJ2ueHDnz5bMa1pHyJSW4p7osbLzaMFDKxYs0R6oIJ9W2uy
sGYym8McopJGHZ9lBChaB5esXF9jE5zqcfGSBN/emy/BAHB/j/g6RBo0xNReRQ5FDdPjkNqtbxAA
bVvnt2RSPjVmEB0nXMKUTZH1xS6IN6VEW7HPMZ8tlz5c5I9q3Ja0Y2Fj1cgiFNuv4s1WbH0HLPyw
yAT4eogXckYfhzeJfwg/ZsQ+DveNVA3W2x8UyZcQM3KsbKCuHBNpTad3y1hafqU9Td0Cq/MvY/p5
GizX7kYkzbR1QplsTijW4828AlNdWJejVad0lj85/qBPX4acF6zRGnToe452jDDzUYuN07KWqumB
RvXnZMPsKdw2wY7sqyO8gEn2yKMoi0f0kAOzmGLsdZDVm2Lq3vwjGSwvyRNWejPpWhRmUQ6EUvrv
+kelUWjkJh8PMepF4aBqaNquPIw24VKiQavfrpnIz/MhSK+NV1Syb3SryetKVxZlYmPZdq8zQHRO
jPZprZZsa23YWm00d5I334PzrZMMdVgA367yRlMK++iiv0s3v3qc1OrD4Eindy9tTG3TG5fh9nTe
ahfuSDBVr+tlD7E1yEPSEeQ+ki1rrVFN00Al2dgiqwniJ58kGm2GXBpoI9PVTksZLW1hCEkARTxr
iEhzEqMj3loHIL4T31SEWpXMZvfvfE6TehcTLMF3qxFNjzGV0naTLeWcF4HS94hRQt13JDyZv6LZ
j8u8OmncjArejxWGUc+4qa/sfreYtj6QxJ0itSif1cz8xqIruGQwYHyLk/5pq653X7XTnf6Anmcy
y9duKFcCoGBUNdPHfcn8g7aSfzhcfZTwpfQ+uSysQifXUCuG3Lm0Jw0FjffuuobZFIYIA1ifWEKv
STPOueeCwCLFitrka9YpmNURnEGmgPgJSfmALM6MPeUw54AWokhCq32gb3+k3uPQTDczFDv/D/yk
A2Z467RiGx3PT1xUZAPRzU0JRM+RmIkUGP3RHN+yIlQhuVi+C2CPZ6JKElwSw5JgtluWUQOcx0Wk
LVrTRESvx+Mrm9iM2nwSlyppxhA9JAlAZhMeRGVoPqo80P5Uw10++YViq5TCiZMg7FO4rybW7MQT
a8g7W8uwG7Dgit84Y8cPkE/NcF4JjrpUkoOr2nfyF6c4yOQDsh24ZSbGcxS8T8lyjy8GrGijUswX
Eec2aCNSztzSu8s+1ctVcMW1iFMK6E3Ob84ajg+JMpVkXonKpzFeH5C9sawbM7pMs02/LKqPb5o4
/hXnJ9ei97SPs4RggonCD9QXjnIPphrvJDUHyTJss107v7lvd9wcrcpmeI8MUGfpqAK9dsIWKmyl
02KVbLnw/7mCcOkmrCqGYcJoh4NVFMd0qrWG1n91FZvAZZpCOYnv4AJIZ2XU160f/Ym9Y/jN3/TJ
HsLJuPpAfsOC+lVCMHHCE1v8UNz4F2+fFMGT+r1Hfimpf04HzzNOpMFg3PyRUHzQDsUjjf7LDkOP
ZIYny8K/SZVJl6N+EGXYvxLEnQyOdm/zKRfrNce2o5b6FtPKNfYelzMxnOQwWWGTlgIMJlw8DJYR
k2p2Pi8YnNr8/GJtcrLYNU7TWZgLvB1WOZ+z666sPZXbcCY3Jca9yNBKDJ23APz1v0y+WdoExf+q
A95/24lFk1R8CYZFqkd0kUmnbNK+dXJyil5ZNYq3c6jAxA0hx0JHkyvEctNKSNytHkCV7k/yy8nc
O7N5DtNi0AViBxgwV8RSbmTB96Xrt+cH2VpiwlYU8YCXggOPqtJKDoVkmzBxLN+e5ocOUpqxoLbn
uGFF2xjXe3CNcfXJ71RXCrOOuf53WLSKtI7h9UMiUQnqE1Fd6FfXWCn5mLnjlHS5r3Tj8kDIxTeI
2tJTQ427XuIo5cF0RpvAdmF/bywTi4G60CnAZ1hFy7sVK4WEN3U2B2PFqYE/FJC4HAsm1Mi9Lvty
QUS7DQLAFIG9M/W/2ZdtAm6CklSdibmMP/0Ojyn2VmpS/+Z2pVU8IhtpP8p+yM7XMXzjaBCsLTbE
xO44BgZKXPFuvNC4VLoQKrtTefSwj2UD/KqGojb1gfnzFiv0fzPikD3ZJYp13lLrtSLwaGtximd2
irero7n2bnIPIBsdkREodt6v0ZNqNUO4lFbsdZW0/FtjKCpweKGqp1fb+BFc7i8a1u1r0nbaYgIZ
5tA07qeW0WoFrrjwDWiBkSrT0Xw5C6kfmcmnZSIu8znc39MSR7FH1e6Xt8bHzfV/FlP+DzWVLPac
V9CDrxZZ2H5Bq9SN5eu66dI56uWaYbtwDSKdzMDqe2SG2b6dK88KELN2bxFEvducPFx/HsWHKTe/
4KNCqbK6+6S/SKVqyElVxigi56Wj0tC67++DCaIvR/h3pXX12ztugyxhrjSSGynMYx26MqZD5u2x
/8tJZr0t77Wi7XREtZNbs3gbleE8GXLVB1Wyl3vOTJASVpeL5n5PqX92eqo8JFLti7F8C2+XaavB
oWkz1+PhI/+QCUG+UBQQXHEdQtl/6brK7PUJ0RTwEufrHpFNb/Mu2v0dyR2Aa3/GNLSOESY3hetI
TtVKfYftTnq/hSblgsrQHJtJRUYrJtb38O3IFuFAA/P8ZYZHrqjc7iFzok3JR22M/3IoMcaoo264
uihGYQnAHm3GmI8tWoodHWqaeMAZoHFwgxzE2N9rAhQWGUDJZn89ELhQIzRiDVyaKxZrcnL8UpvQ
/QNxZ4eLDEd9Oqp02DsF2EiBxj455lhFaqvHeFxdkF289g1dusykfuahJ3rXzGxhHJQ54KiHC0ui
VP0uMk9jh8xh9KE6yoskOQE6iDn8kPGh8qleYJ04g3vI03IvGlMmJRziJnX0oQCMcg2QFO03YWRV
oyX97IrRiIcWQSEURuF/6r8ddeJNKMK8U4jj+4Clr+IFJ8CpCHttEAWGZ+Odbr7yh7DHc7hdCdI7
69luFNpXReL2EXkyGyFA8JLQrP1eoHKVZm0mvngwzuv0JFY/aGMP0MjdboIFw0zv/NUB9QPg98S4
PSFTNVxvUQC24NhtQQeSoadetr3HXoStU5aGTvJZA+K0wJ3G/yYXr+18JGzdhRUxGoZJ4u0ZigrZ
dcSNuTMqyMejqwUK8bOdtjEUC45tFkerV5Unxr80WcGYzwPzt/1nUkFMnMvlZgZRhJ/Oo65ZTDqt
e3jdYtK0kBIn1NS750bFV95Z7xfG887YwGzH/4HBI+EKeOrBO11F9EkpMZ3nwxODLNxYROUVbyjB
P4WoTfCOGc8oYEa3q9y+b/cs1jGoyqwC9vJrF77UYw5DOouQHcVzxoNV5y123+Z4tlrgm1TK0Gqr
zR0+qloLpck9tNHYJQ7lXZyirRbilGQm6rBJ0EYoprq4cN9DIq9dhHvFFRpV0xeMuGf1LfkzDO4u
IUCd09S6kIN9xDNrFC7KQYak0ehIi2B0wkhdHz99gRNRzKpPZnesDvF6j/omN3xcIME3/3MTvEtZ
8qh35oeHTUc86+ePw5QEb1eQdwMbgi+AI5h5rUnf2oJgnGk6cK52bTb1WJIWdi0sb5K+XKJO7VUA
jBVpRiye8rH12So8+9P/oISd9hAloP0nruYhCq/JWiBPj82wU15Uo7g1Z/zg2mM4UFCAoYw7Q09d
e+8lxbs+s7etPAuTkjJQPCPvF4lcehi+h3Q46ox+hz3Y1BrKvd9rieFUUCATLWuBGB7V+apdtW1C
S0E6iSZsRMGJ8l4sFE5CJ30mtn5NW2qGVSMmY0wtmZtfxkhgwmdSvSV7mx1l2EDn4xj9MljA/95h
lX90cAnu/5HRnt/DSQloAp0/FtFbXAfj9peADJrSeKbIpI/cq/iydqlSbiQhgn3jZtijL2JM0cGj
ZNvROJTEzOpN5Xql+5mzoARMx1BiqPURY/+0/+68z4n4zJmTQ47AwN6x6k7JZSWhVZoex/6RZTP+
GBcSgFN4vMnt1jyWkBTPp4EuVVOQ3D75JFPLIkGvlxMXNpMqwL3ZVKZ4ur93i5HUlqs5FSzhLD6j
Bt8JialHwdZ18I7cqwHNjzsvZIeVtJSs507Pr4VbGZp3BDbU2aBH2umPc9iBnk69OFzZ7Xezuck2
hK742Z7ABBc7aKKRzWTwj3wdvyCp+9I9ypcjRnHvgJqex3oPKDbhTXBRAShKRQktqlI8GK/XfDbP
DdHhfJGQrBQp0ufRuLVkVusfhcVLkFeGq1noB2v67dr6Wgv/a+gWRrFSQ6GR4+NGfnMK5oegJKk3
FYbjv6k3OGrqdFBrpJWywnbXgWoiV6c1nmJq/s6cmtP0Mn6lRd5z9pvjcPnjzMhE0PvWiuR/X4kI
/wJZX90gPKGtULr293WrvjiVnylFjm2b6spKiXFMUtUq2xVx6chqugYSkRp0X0Np1ubBKQ2kzc6O
VvAaK6OpADtk7u3mkeR1LVWBAk6UcKo0VAvkLo7i3xynach1iAXDIhgIAVtZ4fyyUilZo9X6Iek8
7L9tuZFefptrAFQtID4pBSBi4AV40O2YSW0mFfjnYHDnbtOXVgi6PKSGhRv1n2GO9SU66r+ppjZ/
+HSCglSO7AwZbp8LjzOeSmHqbh/MhazwgtrRfWfcEf7jrl5VgfZwtHw2I9hIf0EAC+s/wrXAN9V1
5xpgVoCj9XFv1zmgfb9MrbxuypLNrFkLyDfeew1zY1D8zwaDyAfRbLZPcO/UMCEW1MjCIxMxl9yP
3lYqA8V67AtQ+XG2xapPkp4uaL6T+Q1WiX8H02o4nCtzhp/h8zjAiBw48CjNz9xTqncc03YjkCTX
9CwsyLD3bQVHbIAXLPaLxMIYqqP0W2VEtYKgTR1DS8K2tsJJLZBwUVJNxKi8tozJkSOTUQr3LJKb
3WAq02taYrGv2lZ7fP2NVDZDLHqQlpc3LNsKZ0y8uYWIV9AufKbZ82SIpNbvMFCryiRVL8+WWwlH
WPj6Ci76LYtKoII1IUWQvRirMBd8OqrH4oh1B5YXv7sD4lgvCxCWRTwg71WoviTiJ3Y8ZkmUquua
w/NLYcbJhxajPW+2eewOByYcS107eC3jYZm3dTb3iRUCIIwFIqPrFVOaqRFgKMQkAC9mxw4MXABB
FA4NE953596dMMKxz283MV9zcUEU47C41V6pUfND2KTq0XLocKitcmUwr1YEEidocXJsVXdGAXOB
PK+80kHz1NqFNtemggmQZcFrhtM3BsJ+0vKv5RV4hTpwUkLdUeSLM+KlA/X+1OYjzGaST1ydhh2u
wcUJZ7k+vOtjJ0MPev8Fl2OYmiCnOlMxaAyrINHNWHsH2o3jfjoftWitxEttbQSvlZpCYPIs32th
KJv3x6uAgrIL3Ce0KpK7TRGzGDqVfymjfDIYLv5M7M8/oYhXmcmB8AREnp/m+JcCoTrhHG7CG0vO
woIKHFgeL0+hgoGIa1EECHenwNiWuZfoi3jJTwdtm4fYdjrQ5jzXmhlmQsOPk1sn/CAXow8Ielib
dItVTuHVHVJ4fll6cV4l2kIgCDlZSjk5MN9LHHjxYOUGssFIOiBiBEcZXNibt2wj5CYNoT99KgYl
zm5QKhwASdBHXM/5rVXdvgv70xX169tdMRKfE73UhxHlH6BtGmQDwd9buQyStuY3bC7g6OR47AGG
Yn7mBEHb3AQI9K+N8daeRbWyqN2AuCS35mSeAhTzt4Qjx0lMxVnT1I6fWu9XDH40CD22UnwfibL5
w+UHM+vOXzre+IdJg1Il+C3PDi+aX9kwhL7Vg1Io08KU+w7Gr9vcUpcAAJbHBDDzyDf2VG3R1Nmr
OpPWBU7zMT87nvbvfcfgoOQvjmAkeEWhsE5djBMd7MGBBUkSVBGkxCpohlMIzrcj9UvY3uZi3LOh
YsdIYHqL2egAWoMMsA1C3SHcsE0FHD5TW+beRkmjrnkHbrcs1QXpHjl/wUVOH2A+TjR+/xaVMrLG
hVLbW0O3oENDWYK3OrICMdnCjWVK+H5+21fJh+y8E9UqZz3zXy21OGmobEra8CdtDQ8HE/t4hLNx
LXC1wmn9JD5xEAEAdanAKhvwctppf3eOuvT8eOPfBp9dCmne05fuTocKe5tSPTJZIPIvyRv11jqL
8BI46PsrKBAzHK0hZIt55nDzRGFVmJhe96L5QZlgVcmvZ9Bci+vPWsV1BZiSvD6jTsAkgzXE1a2a
4jApt3QnusdWMHXbRHaLMIdtA34HgIrHW+S2KtHkCUeEL3vR0qhVFA3EgznixFk33DfKhWPmPyDk
mb7FwuDKDv45lIRjO6I4w6Ojlh7H34qvrxywZFTr9JK/c5wUwxirO+2CoIILy7wCkdr12wPhopXV
71oIpvSnQ/R6RfOTByisbUH3yDpH45qRhOFKeK0C4JMJdR1WkXw75pkDQml7TVXVImbpKaFTbuPW
CMhicfy551ouK04qTvKwQbmDwlRM/FANmpMaRDN0txz3hWSxDH67WdhHGL1qb1UU8DA5pMq9jJzt
9hUm5QwG1NPjatoY3mwZNOoyOcNkwp4tgI4PRRr9+1w0WS9gIRYfx8zA3LxZXVvJaE51iL3fL7wD
fP2j39sEWOuEK0ojxYurDekv7gc4ZdSw1HxqVGdfNX6e5mN5P923l++Hk2GL7dFJT+VaqpsWrzZh
5qsCWgE3bW/Ej9So3nnudeq6IqMmhZfpF6vQZxN2h2MYmHmVuIrjmvwfpoPzJ0N0Yqi1A/GD1Z7z
bHvVEYu/MJ6EjJNObmdXqWRHiwyAMcoJQHWynaownFfIuia9GgHg+ecFoR4uoNHPJwZivUNfQhMK
gDM5DkfdconYyI0+mfBaHRBmW3jUz9OkBX8mdP257q4P35kzlXKGWH0Jy1wy3PVCXYS0NY/L9Mxu
42uDC3YV9l+ITzXoARKP1ynOQ4I7iSYFOeDe3IXqeEFPSI+wCEgouwLCBL1GER12YceK5brNP7W6
Wr4FOivwEgBnQ/FGpQzXjmi0E+yGx6Y3peIne4hlXj4JnBh1A0BDoyNvs/Fl3cnT+xJeEjzeusIm
a+rMV1jL8fY5E3T3ZA6HLN0jnEemy8K/9asgqBdpd20jy7/XloSmpXK6dCM70G9LQTLMY6c2knaP
W5RiSreNbRayxqQKBkQk4F3uYLCDBa7Fy+C8TdVBYWDF7JPpJ0UR0DhzrewkyRNn6tkBpVJkFIiR
AYRBKFI5AHJoIuPxnukyRCCy0KShTB8eD6lb5RItP7VqNYsfV5T16y7yNHDZssXogllnd9FL3zHq
ArG6m+Jy9IlQTKXI3ab0cQMBHsvAHMh6NeDUVLV2EQt6LA/lR3udAoOjBg==
`protect end_protected
