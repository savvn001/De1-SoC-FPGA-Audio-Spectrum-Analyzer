��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl9���RA���n� K9SX`�/�V�7��hm�4'0w2��	{tkF��QfRV�ٰ�R$=����Ƹ�9:sC�0�W^����(�os�-�8�OD����Y�/s��;�C3��� �ɞ��I�3)��J=$=��0q{������>�v�ߖ��}�]��ˁl%8��i�:v^��<%�o���#-F�_���*�p@�b���?~]�V���_�,�|�d�cooJ�%�x�xB�^s�mg/b�]�1NW7���v`������쀊�ӥŻǰ�0~ݿeR���9��+qy�,xcq�	��$,��ƥ7�/�suV�Y��7z�4�	MB!xx�Y�\�b�+cMf��N�g�u�.�8��b-9�q&X�s���9�V�st������ uE]�'�@P�eJf���+ǣv��<m�&�,�
����[��֫��JHE�g3m�ww�~g$�`���#ej[V�Q�@e�hin2K4�������uRJa^X����"6�a�Զ���!�_<(���^#���e>9:N@'A�P�1�`���:l}�/����
�ٜ�R�;����~��2hH�3��>�Y�P$B��y^q4���1�����@���n-�SIJ`�"h}��
tۤE��V���&��򐐙ƿ��m��GIf�f{����aǲ?�7�vc�K�2�%?���j��W�}&ݿ��&��8�
[����Q��+JG�86ް��o*�<.M��yDT~M,�t�>��K�,\��@=�e�I���9��Es�A���3��#w�vy���p�G����9~�ޜS�+���_�"مY{:�\ AB�̋^GD���f]$�rg(ٗtMW^�#��CGL�:+sl�ا�
r����:"z�d��%d�a�g��%]�� ޑ��L�4i���t��ʠ(K��.�[����Y0��P�����z(0�I[5���#�'��A��`��2��m�xW��_T�K��'���ԥ�A��O-f^�aч>�d=�d>�~�u��3zf����#MU@���Yڷze�<?Ot���-�1j��̯́2z׼��T�]5G���ϩ�<�[�53Цb�y��;�neWPTƁkN������?��̞�8n�|~��h��r/A,ģ��O�J�����4[�{�J�����Pꐵ��j� ��#L����4w�75ng�_�⟹�}AQ���|²!7�b���}��u0_�J�洉�x���:���
:��k'�u�F��"�Y��زy�����,��oek�Z��೬�v�0h��x�b���mLP����㢬�xI�ﲱ)aPf��j���F��r�C�b�i� V0ޒn�VC;����t��Z�T��k3TZ��B=��D-u�6<�6��D��B^��Ej�LN��oO:]sq+�:�MP@�MN5ث/��R �*r���Yح|��?�u���ԅ��.��_;m��)�T�i,! �����-s����m�p&kR��/�6'Y\���	����)j7�:��`��<�ή� w�"h�-�mB4Ѩ��E,���U��"�O@�vO˽�R�Y�+����!u[��>
�P�,Fp�5&��#5���`F��d���˛=Re��	L��vΐw\�x˗H�遙��|�`�V�'1�b�N�}U+O �NiF�����$�[p���78�����j�(����:#�c|����$���|�>|������ǟ�:��ѥul4Aw�MJ�[����;m��?��=�q
�I��/��F-Щ��!V?��F�=�5��D�p,����-��w��P��>ٷG�[~H=᠟�q�v�����/�P�"	/|q+�{��@�+_~����)l��lIȼ����<�h|���$�_<��R�P�]��b��6�C0�6��)Lm�ҥ�|���R����f��̹?�4(�K���%`�ܘj�N�ˬ��p��PZ&���9�!V�D�7Bo*;H��K�S�/�V^G��N��a恍3;͔�o]z��r���g����9;����{���fvR~�Ua��?����6'�7���KN��S{��=��.����̍T7~�~���W�3��O�),Vhv�Q��� ~gqo`H/n�:�}�YO�kUJ_bA���0�'^k0W�D%�mh�֔�W2�$J� �wz|�3�+3D�����Z#��o��E�鳱��m�4n��6�?"�8#���ǽ��$�)��V�hO�����U���v0����� 0�+C�N�a�xs�s	unb8;����꽈a�����N=�Qr��i	�=َ]0�FqU��q�ۆW�N�sC^5��[�]'fp|�������^[����!�j�� \�}�Q��Y�3���Ubmu~D�����+KG�/E�%�U>���:�-�Ȉϸd�Hd�=D���dx��%gt�N��!�A�Տ��3�=��n�h�>>S|��nЫ��́I����؉��YeA<>e�sE�@�e HS��7�B���b��q�����7�iF�V�+(�C��fz}D���?y�Y���:v�N[X�A����@�տ�	�͘5�0�*�H�H�"Sp�Y��X�;u7�ڡ�3�+�����If&ҡ�'��M[�*p[�!�@;�U@����I,iV4��k&�N�K��|���";���m���	�mE�W/�ZU����cx�w��rzc?�F���|���Ќ&�㢇	�M�J��i����r�&�� ��a�^��)���k��H;k���Y&��������{�`W��
*��)��!"�%����=B��7vmI%�9������+��2�ʓ{�������3�f):���ǌmV_C2�p\\�S4��T�Y�<���jb9�鿤S|�iO�
m���,K\�Ojyo�jX�C$1U��B�G�;cR��y4̓�ߺ��I�!��ڹ �z����O����;��'�Y���#������i.Y?A��ju��"�$!͟���R�0�*%C����=j3�-�#
��1s]��U���ʠbZN-y,�S�$���_���&��/�+&�Y��!�D�|�i�jB����N[H�Zu����*KBH���Z��#��[���v�$� h<����w�tݓ� �X�����P~��ʚ�ZU@t�Ϩ�����{��\�r?����I���BZ��sko��gC;��[ݰ�Z�j�'0o�2D�;�`��#X�wIE2���w�=���}����/�kvu�,�I�#w#�C�����	i.���i�vKѸ2P|��gs���T���)��F���/( _�фF���P�~	u���ݠ�7�v.k�ѐh�
~Y��I:]������I��)'�w�5�ptA���^��Q�؍�D�J�ŔE0a��xK�w�6w�*�����3o�ʍ�Uh�2�B��H���;�����J��R�SY��U�@j�;�1�w�f"�%���74�ˬ�*)�I�_��?�E1�������L_�8��>c���=�T��^�O���������:.� nUE�^�1�O�����h �H����� Y�%���^&�/S���2�VE�W��/^� W���ZLiUP
X����1��->*��$�n$���T�����I|�z���R,��4��'�1�<��2,:+Pq#�M��Qr�040�|Jz��³OP�*�`z��߷Z�^�c��L���(v�k�2�ְjY&t#γ\�PޮHɇ��(��18R&�[d������b,�Ϧ=P�ӥ��8�3P��X{��n��]�]m������@��ݣ�\ܮ���	�ķ@�+��G��iA��8�d!�����2���}B>��~W�������-���������R��[�ٿѭծڮ ��ҿ�	{���a<�P�>
J&@ς@����	��L@��^OΝ�vO:�DgaS*޲��2gQ���m�揭�QV����e��x�}�e�)"��ݴ��v�!��F��0.���T�87�����.���dBm� %z���f�^|x�8Q��܄q�'>�-�	j�6�Q:�ǵ��@��&�k�
������ް��i�&����b�m�D��L��[�hȯ��ѷ��ds��v�{[��4��S��+�ӂ�[�9@�M����E,֕�h���� ���re A�0�t@�]A��}���\\zǹ�_9#2Z�5���ׂj�ٿw;r�9�iZ}"���H@�՗�L�r���k��MI���Ir��S��xu0b+)�)�
\`2���������s�d/e���n�ds,&�?�����ً����!�o��J:�w|`��"�m�l���C�ccU���"%���u�\�����0���#�N �m�rfo"k�?sl�����A��#&2	�PH�!7g?O�0���Nkh6����K~g����Bl�d��zK ����NBX��Y�ב��Sk���7��l���3n�g&�����l��a�哱�0[\M?�{�����Ԫ(@(��hT"�eW0��~C�Ȇ���H�0��8eˆ��^~�"h���M�!�k+��_�_���vFy��b�'���ء�Z&�&�'���cpCCi���.fH˹]�����;n�,��~Ub���7.k|x>�<��9^v��IO�uA��ޥ�\���9�ʾ7&�u��BS=���1hϒ:�B�����Uj�(c�Z�%H�T��T� 4�Zz�Q�}��?*���(��8y&I?���~u��{�mf\!�[�.�C�0=���Ā1�b$:.D~�;T�:(-�ɤ��h͚��դ�
����k����}r�?	x�ݔ�f���x�f��6���@�.�^g���pȸ�!��r]�l�OĚv>��0�E�A��0�M0R"����]���F�)~ir�Y	(�x��Or&��O�"Z�0|�q;�<@�΃�B�-.��)-�'j�]��<����=Pu�e�gf➺[��-�F�����џ���@�Ļ���Evl>9������7��$�J={m�vy��^ʚ���ye�Ip���@�p�=������L]O,Q2�.f�8&���Xs0�ٗ���t�]�z�@���F��l�H@�3��:��F/|��*lx�-�������	&S��Ҋ+K����8@���[�ϐ��~���e�g-�X�t��W���e�_|�+O}Fr(�t�s@�ۃ�O3K(�/^HQoA���*��m��q�<4D6��^���;{��uIk���7;�.`_�<��B��Ʒ�H��.��ٯ��jz����2�?���1�G�۸AH��.f�h){v�v�I.���B�KM�k{Ĕ���^c8���S��$��!� ��g����Q�5�[R�B���5C�s�>8�	Ԕ�b�`X��q�.y�������X v�x�~k����wGT�h^^?�;��圅��/����j҅f2��������i�	�/���v|�f싏'-(��݌�1�s�%�iY��[z;��&� q�U�^Is��n��\�}��}^�7\������\0m�����Uu)�5V�7g&O�U�2��!���Z*49�����ڡZ�W��f9����>�,�#G��s�p|F��~�Q��Q����ӛ����K��,ja{ǧ������q���%�y!L���uko�,��-��Q���b��9��/K�5�}��R���Z?J����@b�?��0jT��d��RG�F�1�9���3�V8D����J������|A�{#��S��S����]�_��K�L����<�f�G}iy�{ �.O�ء@	5k��ކR�L͇�i$aۧYMb�ΎEcE
����c�}Zg
�N��O���tU�H�`��"�;C�a�a��_"��-T�l�үNDO���?"�����SN3F�y����݈A��i�5�d�
a	
2�X���W�yD)�����3W ��P�ڭA��/Vy ��VLڥʨ���þ
T�Ս3g�t�:+���=]۾�7?)�Iٜ.�p�P��|~;�@����tF��^Nr��3f�m�[�$׷��׼>[���ER]p��d*��H�"ר�fjr~�>5���lz	�����!	}�o1�'�+�W�O��\n`$��E�����"yE��^2�QRk9^K��Y�?kY�īG�'ȃ�-�=��.�02���{�׷}�D�7�=���]��5��|	Bc��K;qÜ(8�����b�S�)4�ϡ	|���A�Jq�^:@��3�l�"�{�/�4FJ���!&�pŵ�m�����ӳ��̮<L9�-�|R_��#}cv60�(��t���R�;S�y��$2����]#����v,�n��eX�%����L���}�d��y=ZAVrG�DK�t\z �ڨ�v����:�����t�0 ���p��躾I��Lo�z#�wo���h��uN�ewf���¨��XC|�^(��4���X5X��i�k�����b�9n ��pW�q-�M��u�2.��-Ɲ����* ��������<)��dEQ�C�ũh�L�u��)p�"〬l�#��B圄!	�6$4����a�*~![�m[Y�2����qT��3�G}�٧���gY=���*���������p%���,2��L�s<Ε�t�߯vHbq�
��)���#*��n��ؤ��{��W_�-m[�#��t?2-��}A���	�&q��畈R��#�	S�5-*d���袕#V&(�����ٔ���l!X�h�PI�"9�R9B9��_k��}Ĳ��~�$�����n�ҾO�O.��f���]�~2ˢۧ�Ѵ��0�y�G�`����n�JZp/s���,�5<�4�\.&�I|M9��;x��4�مT�� <L��$�0��x���T:�
�&S'z�t���M�4�j}������#ss<���i�U����xZ�	�B_[����[pBFJ=ߗs��k�_�
t�(<� �i�Y� ?È~)��������
^O���ꋤ>����$���> y�5��l
8J� �.IC��rE �{6e�o�9��G
=���>N-�cL�mx�I�w�<�T�639��Ϩ����e
c-�%�ך3�T�s��$�pw��R�>����3!�eĩ��� ����O�U�ɂk߬�
�[��Q��xlO
-�+q���v�krSz�`���5��p�gB��q����J������T�P��� �}(1�Iָ���*�s�?M~�ٳЫ�n�����{c"�5E�Q9�����%;"g�8�	��/o���l+ǡׂ ��c��h0vm;/��Kyr9T��BA�N�%�����)e��Uj�M:��;����H��Xlβ�&���"��x=՘���*��,Η �<��ǼJ7��-�aף���M��E�J�=d������s.5sK�^:h7�ئ��1"��p��X';Q�h��He<c�ʣ��{h(�V�9��럯�I�DL�m�� 1������IK^��o��[��O�\nqDQ�?0ƌ�⠈�i$������䨔R��"�%{��Z�u��2>o=������ҍ��׸��0s�磭���D��⬶>���;��I������������w��`?��+TgLs�k�:!�::=m��A�!�M4���xźU���֔^�Ȼ��H(}��G"�A��*�J�4��^`e$�ȃe���O(�G ���_������7r��P������,��X�����AGT6Tl+��%���W�"�f���S���zY'\�O�GFPs��/���������T�LP�E`K��w��c<���&��θ;��$���	Q8_�_Ɇ~�v�@O��O���ϑܼ��Q��(��=ʗ��#���ЙK%�T@������i^b�n6#��
}~�½8���6�FiKP�����7�_qGd3�W�l;�ȇ
�Ϥ����R���m�� ������������:����L��>�.ka�!�H7ʬOt��c����,8�"�K��/��C�м�B�lJP'��:�_3���ʹZ�`�d�1ԓ�WP_�h��y4�a �]:lF��C�۞t*���[��"�2��6iI����/t[��_۩�oM�65�Aye����w�a�>Q )��V��2WB���������.���7�(G!���mn��� �1����O.���_;���;jJ�k)V��G\��_�{�s4��`���+|�_�����:�"N�ɋ葭�EK��ǳ;���j��UGe"�m��}��`�o��ζHV�f���U�n�_�m`>wN�*��:Ao��&f���B"Rx�p̥�;*�ev�4FM\h/,�*e/6
��φ;Y�<D�]"�Fxt���	K�t�r>跔��!?�[i�?�d>�f
��r�����d���1T�7���iV6���y�tf�_Y���Oޯy0�hVv�Lb\���I/��� �Q1��7���~X�Щ�.��(.o;���T�z�_��b"�h/��I���-���Q�h�c�=����ʕ� �A�b%[�;J�zO���j5��:�IR�@#�و���z=�4uR���s����z�(�?�����ܓ��K'������-���2tW�.��xW�,�)4{�L������ d�����e�b]�.]�8�r)�(�к���͊����ƿ����yqw�vi���fj�?��(�C���f\Q�d�Q��.���d�lg�,U"��Ӹ�� C`��cgz�w�*���j+Dȶ�X�a ��p�7As7�e?�+�9/�M!s/�!�[�a�����L���[�}'���I���nֹ~J̐,��-M`�,D���Q�7��1-�B��Yn�ǵس��?�LH�n�c���
c�׭)g�r�I�c�s
�dM����5����bpMs�+Ɩ4ET#Fو稁�+/{QX����y:��ێ�-��r��B�J�3#�%�����l;+��Gr~����~�.�J�,vV�����3n�(�-[s�,�e�,���e'F���A�ME�ܜY����{�O�e��Ql)|�����N�㵾{Ҡ�GAo��:�eM�ȉ�2�ӻ-K`�m�Bn�H��_���ŖD���՞32�-'��0i�`�Qk�b�$H8�6΄C��o�vm�2�R����}�J��������G,�رܡ�H�-y�L��Dv��ـ����Ɋb�&��R�]�R
��wz�b�˅���I\�y��>�$Gpd#k�]���./#�ԏ;U��>��w�ѼͰ+�� I�{8�u�I��k���/�� ��u�.�g-G����<KT��*�K�9f�gj%�MpG��g?L�G|���=�Z�h���Ez���U"GtV^;h�a%
�儏�\�Kz$0����|������|;�a׵EՒ������)�\Q	��G�[�d&g�{�b�>��|�I��&O��@��'ɾ�U���yg����PZ[�D{S��G�IT�Kɤi�@æ��ڙ ��g�	읥�ڃ�nWZW�m�k���+�e���"�� �μy����_���p��Xة�푂�R���m���$��8cB݂�'�I���0�\P��N#�xp�F�M6⮽f�gs�U��+Tc4Mҧ:��x0~���#�z�a�We���*�v�@}pG熔��%I�)��@ �"���������jQbN��Q�>L{����}'Y���?qA�Y�U��l�#d_�K�ړå���&�Qtj�J��_Vb9t�q�p+r���9�����-
J!���r����� �I��k77�9�H�����c;f�\���[!y��Qd�}lZ6pY�	2{�(e�Deޱ%�p߇��d�h�z�%~�l/b-QN��� ��TEX���f'&(P���6b�O�Q�w�Z���H���cbSm����,o��:�"j��9�vS�Bf�F��mm�B�%ƭ�9��6�R��jR][{0�5HR�!�a�x]�dh*�,X\�p�uuo�k�,�hH�i������}�\ I����cB������}]�v0��XR'��4�<�$��M2�@�|��ƷԴ�Q�ZG��J[B[�Sk�g]g "A5A��U�' ;0��j�E��%�M�*I��LQm|�q�������J���V햓gk��`tI����ǝ<x3.�bG)[��@J���ʱ;jJ�@�^Ěw��~r���z�9��h�V/"������y�͔!��;e�d�(|�.,�s�͗�Y��-���Q���)��i�%�3���8���Ro���1+��ҏ�G�ݐ�|]��Ϣ�G���㗈��F�IG�*J��ʇ��0�y���f�jԙ�?����b�Mξ<]��>� ҙ�{���iD�7�&t��m�BW��a�=�=�:7@���*\z��~k��T��ND��mD��"������J�@(=�Q��{�v����A�e!���*��EN7�����G�Z��G��ц���
�r ?�V��)�5���u"hM�d{l��?t$����7�M;*>,���@P�ԩk�y�E 5^:m!&�8(k�<8�����NlӐ�� ��V��e���^����C2-	��Y��Y���{cI�+٧4=&�!�㒾�W���u�O�ձm1����~�1Ć�x8J6qqd�Q_{���ˏ��i�^�J��a�P%`f���jF�z~'KP}H5��%�ί`M�z��e^}��?/�,�M{���^����-o�Hhs«��F�h6����B���|�\t�uK�ԛMܱ;��T�A��	�R}�(q�3	����TR�t!�'T�@���,���`�)�EM�b����Nf���nbZ�YB?�l�Y<�O�k+��~�����+���\&�	��VA�m#hfj��U�/3/Z����da��4��&Ш��ё>]��t�Z՝d<���ܲ�O�P�u!�G8�NB�x`G���"�$�5��o�Ӓ�u}���B3.�)[��<sճ��8*�z�Z�m����2��N�����L/����0�������-I,M���iV�ff�oW�ťu���l��y��
�~����:JV�BBh@�a�ס��g��gh1O{��-�����޾GJ��0�G�bRƹ)�2�-­zd�߆^ZO�^Q�d��8}����$���p8� ���,����]:�cO���Ϋ��m#T%4�=�f�����$����}6�}L ��`	�iI�Uq�F�
�f���\�K��%����É����gv.��W����g/�����m�3�K�f]k�HdՓdA�ϰ��$5���k����}�Z!}���B:��g��a�宨��E��[[nbٕ�rw�OC!]C|���hY���A��]���8�{ő�D��͸�eN4!:���$�p\�KqMf��:F�c3[3�mܮ%�KC%�!a#�8��A�)C�����_�����1/֘N�.����N{��s�[����65�4	��~��1���U�*;|eo/�Ա�x�g�#S�B�ͺH���7�m~�k�-!��/۞x��怞��T���8�����(5EvY�3�:�O2s+
�	(�����}��X�(�GA���v=���:�����'�MV�K�<�T
пű��O��I�!��pe�z�I�'����,��VEB��E����qF��ӁK��Ի�+SR�y՚;{���kA�GrUq�F,�l!��Bl���*�݉�!K)���;H�"�[��V�����bb\�w�� ���e��C�8ʭވ��Uv��5p��֞�͠|в�&�����C�ȼU�`P3�Q�╌QJ�U2��8��
G�����+�|8�قzsO����/�^�S}��Q�ٱvG���k����f�X�)�d\4?��v)K�l�_K���b$L/b��^L����I��l:��{�u�k�
5���|� �3�]%A��2`�/ѶTE�a����Qd���T��$~(����L�Gp�Z��z��e<D��O��Q��]��q�!O5�V�*Sw�E@F=v�O
�*�W|F�ë����֥��cxBI5�}�������*r��Z��2d�Oқl%�#H2w�u/	�@2m[�7LL�%��T���f�n�0�J��� �y���<�9na�k^=�{ݒJ!l'��A�H
�j����0���C������u���}��nQ�[�`���]��/!t��<��T:��r�8���=z���P��-/`}���ԣ�TAmm-�*�n5�}h�[秩n����_y!���K�������.�y��Mn��_��Խt�¢�ȱ�R�����*)�`j��3_վ��
 q���R-h
O����L3�ޱ��}"v�I`B�#/��A�uMi�~04S9����x���\X�D"w��*mgT%�}�R$'I,�k�G�Αx��ä:V�'��U{�ۧYE�c�&r������J�=�_vn_	�PL��$Q��j������b�څ?` ���j��0�^W�QSs��-���x�((��km9֭�Xl
�gM�ly�)���/�\�B!DRDi����O`����8��m��@�.���X⠬  ����O.����jѰ��Dc+m?��J^�y���ڤ`¥K�:��F9�^�ѵp0�m����gk8UmZb]�q���^)�������6Ch��C�h��t݀K�����+=���j�|�	U'k��̌�BZ�ީ�i��A|���0���?�0c��� ~�n�k���~�jVT��'(i�ОQ�#���J>H`}Od�e8r��O`]�x�!�0Ӏ����¿"�����o��ZSy���)X`��]�n�nt�A.�=:�6u�^�d����2�]`�*����s�b!�$_y�A��,���K���`#�>g���ڰ
���Oy�*�2j8_�.���\_j9 �C
2��L�h%$5�V=�&��Y�nC���(`�|p��u�TpP�_W�o]C��,=����(��R����s ��w�]0�d�{]�eGO6�Y�^~ߖ�֕ �a��.;�_�Z2��FѦ�\Jґ$�|�	����
'Uxp���'��:����4��)��E|�(*�bWg�׊�Sv��⠵&j��N9v�S�آ�OY�FW ��/���0�;�M=Ռ�'�U�i��SC:�$���,��;+�i(��e��s��0�@�<��x�#�*�G��g�Ol�Yljv��#��r_����3y�鮛��=ց`�_/'�ъI��J�9wx�ߖ���"i���e<`Q��Օ/��2�����k/�K��l�w���:|Ӈ�nq���� &c/cQ��d����vb��X�&f��U��٪������;>/à���Z;N�D���b��a/;U!)���i���pD ˁRz{*�IQ�<(�J,�kvdp7��<�y���U��B�"��3=ryyb)� ���n���(a;�5���dC��S2<c�c`zN�J�9]�zh�N#��]�:E	��"<�ˉ�K�l��O��%��揪9�Műv�l��%&!ۈHv>�Ɏp�vc>Z�'������M=�+�ki�װ�￝��v4.ϨֵS_� ��0�د=�^ao�8�g�~��"��hʌ���7rG߹7�َA��f�\�Q��ު9/Ӽ���5�*��Z������c�4�"��R���Q.rt.��\r�I��ۋ���C�ݧ���%������9�Ge��߄�'O��uu�]���"�**�Ч]�9�pʍ���#��+����a��@��n��"L����߾�/n���H�u�|jpR�
),�	�Kd���1��e�1�zX��8R��>��7.��a�w5�;Ỹ�t�^p{��`t��������}�g��#�EH�|���Y`��í�7I%�W!m�<��!cl�q�Ր�7LG��L̼�)`;�oll�
m���m�B�>ד҂���=ZM!��>���vŻ��6r��j0�����M��CL�$��8�_+F}>������eM/���*\�&�S��@����J}�L�e��}�O��mB�N�e�G��ב�;V+�h�'�P�d(WF����H�V�9m�>:�'�??���Gܺ����|F7ߜ����%uB�۷����#�D�ꪭ�l*t[�G���������L���U7_K�c��eB���֤���P�0�_��oz���\�p��}�i����&6�T���9u;����Xf|��`Y���?&�����o�ME`w$�7���E*��b�O�B�c��lM*�ڻ#'={t�%�|�2)җ,k5�����NG�-_L�<m��o9���,!}�e���FФ��cۼ�خm7dWzD;��k�`�bƍb�/�s�&-b�{����42 �L:	}���1W��P��(i�!_u�o�9�!���LU蘍(�`�� �=L�9���r�8 ��K�>ӽ9�oMvG��}����ш��4�G��:789?u���]�L���H{3Gw��Nd��$�bH�z���8�����������B�Y��+\x8[~��㥃ǈ粶�@Y��Rt�yO������,��W����7�DL[���1�����(�'΃�d�)��Ou�'8�2P�c��y�̊�Y}kxz�e�ބ�+Mg�}��8D[� }`��# ��\����_ձ�D>��c�7`��V�UԩV$� ���z�΢
�	"�6F�%����^%���[�ōI������u��j��_�)�����{���!X��/	S����4�VeM����G�|��_�rSL�Z'����b�uɩ2Y�"�Ig2"a���
�A��d��5v�~2��ee��X�F)R/�h=��d1�ٽ�t}i�od�#,b���]F�h��> Yތm��X�ӝ[	������%��7�B���`b[6���3��=K �
�Wwݙ a��qr��8ٶ��x�1L
�2���l�v���-���@t�-�U{Նr�>y8G��I���X:xV���ڨn��rǍo��ױ-/��ff�94ޜY�+M��m����v����.���Pf؆!a	�����BX�|�PLg�Ye��$��ɉw;�#C��&m��]�ӯ��'s��~��<��/iU~�E�Ѭ{{+�t���� joRaj<cc��b �B�(�Gr)��a�U)l+�\'�C��#*�d�=֟��nd�-��u,��El��8u��;�xj��!3���&%*ՂfM5��2N�; ��2U�ţ��RޭS`�$�!�gvۼ-�包T?��G��N�}ɉ��5S�/�R44@�gz=�)N=	�Պ�;���%��18��ad,z�蜎0t�#m)+o�ɭi�)��I'� ���+%; L�X�tQ�I�A�؉RG#�N�=}����H �'�h��p�0zu�x�P�g��h�W�ہt��.Rb���	~�S�@������3!� �[vؿ[ۢ��&���N���f�K4��i��pd��Te_4��!�������@X\*�z~��K@�j��/�7G�#����O��qPp kHd$Ż�fl��W@kv��et��y�j�RYs��͹��������ݝ2��&��ʷ6 Q-��07��>�J�/��B��yMy�Z��A�q�Kvc/Jm玲Luu"���>ډ��a�-?F���`QT�Cb�{z[�B�$�
;`5~t)�%���Щ��&!��`��8�n5��yMO�s����F�lK�	��$�H��b�d�<�y�E[���Dǫ���o�?jy���h/RP>�8���0���-���
���Ao$�d��Lhf��§>��9~��Bn292/�֛S��$�sS�^�ͬGB�b��4u�V�i=J�q�Js�|W�v�
B �:[�)��Bo5�;ԯ������s���@p��C�a��6?,�B�\�)BS�����&���7��T;[}�3ͷP���o�n���u�B��"�}C7J+V�ky6fy�b���q��5�z�ȷ\B�F"\.�VT�K����r+��J�R�Z��@�i�޸@

���]a�[X]��,Zso `aw��~$2�͉:��{Sc�Ԍ�$q�p�P�c��%���5�$�'��cV!hxT�G�WS>s��Z�C��ߐkꉐId��z��mD���X�chw'��F~�\��PƟ�X���f�Q��'��OЩ��ā�U.--�	=��i��������V��-ӽ�����C�+f.Y�@��ݖ78��pH�����%B�N;$ފ'Vo 3[F��7(gGM�=m�Ԥ'wA���E�b��~���*��'-�T���:��&By�t���dI�)�F����f(��T�ǌ(�e������%l��?d��p�8k"M}��A�.����O��[+���>��۱>���+U�"��ϥ��*0��������W�rb�2wm�im<��=Nz�����	��;�.g�MA�h��;��0M��_�V�s��g�]�J�V�taXd�b���׈A�&��,���_�X�+e��H��7�F;E.I�=YDŬ&P�p���ϱYi¸�
�΢��C�0Svm�l�ͨ4痁�԰�m� nCi9�=�T�ug�&��m��ф�v���p����/�OmG1�	�������8u�-t�R} �3ccx* ���Z���jA$D�,���g6H1L��*˛�-*V=ă�������1>py�4A�l�@-h�J�\	Iz���-��J[F�6�_��3A.����-vk'�x�Հ!dE�se�[P����, �U��"
+�����H�4��� �</B�B7�H��Me�[��!F�"�f[lW�&Y����ye!��X�T5:g%XDU_��'&������N�P���QΖ�m�г�������}��c__[�]�����i_}����K��tPsi�ek�����j?��P���{>r_`�U9�"8��s8��;��j���6����kE���d���Lw���SB�G�"tZ�_�NqƑ�/������#���D�]f����rX�B����-;cyQ�� @\\��m�Rl�Bۿ�q�h�
�þ�"+�>��|�̀s1ǩ���a�n�8ŷXC��R���.m�i[����E���L+*U�������2���u{�-�$h�-N�R{�:}N|%^����5���ld7t��c�Bbyu\B���3Y���<�D��}�)-�9")��������l����{���  ��n6;n��!_��h��Lu+�4���~�03=,N��7�ܩ�����R����_��/���i2~�zr��IO��A�h����]��#Y���{�J���\1V�����(m���&������� n�=������n�`��x'3׌3��'��к�]�J�o��/�:r�;�TS�;{�)��m�D�7����K��0ƁP���(,;E.�2O�N��ݮVf���!�HܥZ߆�����Ws*�5f�s�����&�<Y��M�A ٷ�!>��V��3�x��%���v�_%C��8�NG D�OZ�g��X��)it��������*�3[�|+�7����<tǙP͜W ��l�$���t�:U�J�"~��{�L���G̦�.7��G� ѩ2;;8԰v����C6)�Pg0 �"��{�GlO{�II���q�BF�$C�*��)mo[z:��W8w��$#4Xkv~�I�|Ώ�l����̜ec��<�qQ���p#�oi���_��"�%��'*�	!&~�}p�yvn���l��~�ʤ[k��Ye켺��ޒ�Sx.��¤A�@�?�
�Ĕ0�e45��=��zԞ~Jh	��kHfa�v
�U��y�]��S�"��)�MA,��6�k����U�L9�.8e��=`���Ԫ��Zj�3�n���x�����Խ������.��~��A��!���=K�fOJ�/�����<Ķ����n�a�d��_6#�(3���)L�}��T.��!�ֿ�N����ў������bI��LN�F�4��.�x�ۻ��S��}m�,��:�ȁM����/_�c�'�ƭ�pY�*M*������8|�)��3J���Uw,9s'{rg��D��u��x$�]�G���u;s�ꘛ��h{�N��*�Z���7�53J��C�9<�]�V<�P?����)��ڞ%]
��B-:S���s-���f�0��  CVyݶ#�@�@M�b�:o8���虌o�k��]>R@�VM�o�9��!fT��H���A�{+��8�h�yz��s<�R�ڤ3>��[�U��+��kqI���򦱻b���L�,�36��k��׾�V
�?SC70���n��������j�:WJ��f_�*�r�m_"��O�b��9mt��<M.~����c�)��.^�7�� ��,u쬡o�(�D�Z7�d�^p���)Ƀ��$&�8��ry+\(ϋ���|�r���7f>���U@����Tl�^�%�yX~�e��D���{$w�#>��Û�~[D�X.�X��:������7�9�J�@�Vou`j�$�5���?5�#�|{Gy��~�%�{>����KzwR�ǰ5�#�-��KA���ᆗ>iN�ŬI�/�7#"7�>�-#F��鴩�$�6!�#���|��p�X[}%Y�Q ɾ|>����Q�za�I��;�+jop����W��[4�),�����ID/�U}K�wu�=Џ�/����]�%ۻ��yj�[�{2eTr��[E�<NVǑd�@-�d�QT�{s�A��5%,��3�
KuLc������P�����Y��6>VͅmR�:����`�|Z�����S 
�Kw3;{l�>�@W (��u'�~��qqɖ�0���H.w���ܨy���Ջg��+|ߛ_�5�r�4:ؚ�5r��=a,��i�'��*t$Ĳ�:2�@�9닟\�n���+���+11��+��89m�[����mzp�ΩXyW�Ru�P�7�eyĕ��f�Ln��f��)�¶�����Yp�rX��y.�=壴�G>?`�%��G����;���-��F�\Y0+���骩*�l�U�R?b?�&�J���2�cQ��&��<��h)��Nn�d�C�KG�D��~�oTc�8��"�1�)(�D7➿Q����fAs)��{>x^	�\���$��m_Dn,�/�u�5����[[5U�1Ղ�%0�$V���^l;w���($�4�,�R���|U7�}�ȼ����\<n`x�9���%�J{i&�>�M'�
�_o��u�c��V&(z�3�`M����A��w���Q]����������4�_@c|����2��
sE�}��mޠf�����U�q�M�!xG��e-.��ŔE!7p�R jX��"K�a0���M�e1�M�����ӛ���5��n�Pྖz�������N����u,�F|i�����#Q����{�#���r�����y������5ߓ٨�+(  D�h��~E�ȓt�*ɴ���+���r�^���� 5����Fڜ��~��I��X��!���k���KJ�^c��CNe}���Er|-WDb�6����pn�q�?W�T���F�	���)[�Dz׊C�e���Ц9 �r���_
�.i�K��t�kn	qœ�[�� ��*�^���=6l�j�v�=����P�FH���ح��z�}���D��87[A0��T����eC#�bL�|{�(�rT)�d=I-�DY�z�W��nR���U��V����W�s�ڍ�6׼�������QG)E������+tcJ�eķGº�F
$�h{HB65��=,s������]tj>NDD����[�2E�d_��Rk��+|N1�����Z%���~7Պ|�p7����K�l��S'���)�
G~�0f���t�<��v�׺:�< B�:^aowwV)I�OyOq�1�yη��_%�1��1O�5������zC#�ôՔ�:�����)�ֻ�0z]V{�+�AyC�X���G
 �
����ܽ�� �;>;է�g����mX����J�,�{עf&�#r�x�D�dV���p���`�a+���B�ᔤ;��O�]
�t�V�+��W�`�F�y��F�<5C��O��s4�;b^N�����g���%��:u���~��5��ؠ�[�I�\��\�|�ϫ><��V�"����c�L�"�T��8que�)�"	e�E��5�Q�Yɍ�Yw�<�Y�/�g�y6��>�q6'(���4�c���@��?Ю���x-T�=˸�#(��@�ֵ����Hb1���i8���p/v̉�hT��Ԇ-�\�<_�{�?)UR����e퇼���z��I$|���� �cd�V�^R%g���e�Hc�K����������AHȐ�t7��x	�C?�Lna��E-˃F|]�,�:z�}I��=��O�������^���k�rd����g��B����X��egm��_�x��N=F~zn�0����1��,�Z�$�}Ǩ�s�Bϭ��x)�6Z����5�CVXDzɇ[n�A����"�#02^Y�v6�������'a��v	�&�A��c���̈́�!{����}�2�J��M��Y"��3,��n���G�ٚ\ɽB�,m�&�ȃyr�bM���n{.}3��}0;�-M��<��`�q�q���[_m�i~t�G��#dR�W�I�����I���#��41�S����}�u�o�Lb@758l�ߚ�il$� �@�h;���D���������a�� u�)<�Nz��i����˶fd��F>��&p�Ș�x3�xl���-�V�sr
I<?(m/��,�+�>���n�ު�&����-:K���]�ޙ�m���p�j(
a����Ĥ����j�]�����'����zk�PN u��r\S�0r/�=�ȵ!�	�CZa.��"���G���M�ut����o̬U�=QFf���$��C��%��/�����_�k�ھ]���ɬ�i=z�8U� 7j�[�[a���m5�T�{9�h��T�#��|��`XBz�ӄ�'��x�a�E�h�ꊤ:A����Y��q�XmC��:B�Uyr��i;�(���!瞫4�-����`��NO�4T��l��[o�(�W#�m7\��Us�55����Ϛq�xv�K�U{���ȿ�|���Pz��EwG-)H�G:�K����\�
� =K��aYH�h�]i��b���4^M��H��x8^e���4KM(�8+�3H<���}�@~�������B��{�����5�2�(�ǔ�Rk�K'�m�`�E���Y���3�A�9#��*�J�J�2S>0{�O��p�ڋ,S���C��8�*��}�� �[���W��Q��'bspկ�0��]ߤw�e�"<��
i4�`,e��u}�ac�eG������~3��ڰ7�J�`�M��h��+�Lu��?�@x$�^3db�ν�8&�+�Yܭ�Z|����TZX�=H�6�id^��s=��r5����߃¡ޗs62-ß�\!Zf�no��M'Xy�0�d���V4��Rl�m��1E���/�JI�VN�&=
���M���m;}[v�d�N�I���`3�&��L%M����~��;x4��4o�	}�q�AU�p���eI�8��FS�(��-��#t���Ѹ���{�$�5ZT� ���&��J�Ɔ B��ŴA{ƚ {��*G�����Y���|��܅>�F��
X
�%�|��ך�1B�@���:�O��u��N�Ҭ}_�"�1V�~h�SJS�.=wY{�a��mIuxj7��42j�ǐS2�[�k��̮=�����$���F� xw���F���-Of��s�)��<EH�J=	�<8.Һ�l(@�����n��d�"��@��2���UXqI6���O���_&oT	<_���)��4:���o����6!$��F�J�U1(���P'/=��Q�i�� b�h���\�`}�R�7�Vz�b$��dCې����2}J��p���&�¬#+��v��-�`��k�Vrj��҄�H����O��2Dt0��X}��J�]���UNo��C����>��2�T��M��y6����j[J!\�]Jk]�f1��"��ۂ�����&����8�]ܪƚ��습X|�"��!�(�nݳ�(k<q{F�V'© ��$�=���m���ǈ8�	�I<��&�|�q�/��^���6&Ń����m��AZk��i�Ӝ���
���r�"�M<[��WH��w���D
��J�-��edt�$�gP�C�����:�U���M��X ](�HF���?�oU��t��{�2��Z�,�&����Um�n�ro(-z�F���i`X�l�Ŋ��L@�v���l�߽b�1yH:>-W��C��M� ��!�-�����jq��&�KwD��#}ܦ.�QEI��<x���_
s�i�f����eɫ �����<�����?���nH�&ͪTZ��ѽi��g$��ۻ�F�7��Z��<�	�^��f~jݕ�)۴U?\?U��a���) s���:I*~_3oG.F81>��$����0p�Ϯ���懗�,Y�$.$�� �<D�ܑ��:`���'�[&����7�����tj�{��/��0�G��,�hO�UR}s�^�����+�N��3!��Bu��bب������ٛW�/5�j�`Qs'�.
�8ey��bN��aư�D.���C��2	V)3�[iٚ@߷~Ff���3����&<'���Ų�|����'j;�Y
��u��cK�O2!.ID�^����Մ0�-;�P�� �X��.G�������C8KH���7t��,i�ݝ*�I)p���)j<�n�:����l&J`:-����^����1+ȏ�y� 徨Im�B�1�w7��
À@�{#�uTL-���b�`�[d_s��.��Cl����qc(�⟌������i���f��J{�����M�h���"�k���&�h���4����e��q����%=y��"LX�b�"�&)��f��� k �(��=�e2��p`��-82��Z8;��[��Y}�I�˩������6��{	��%+�M����	i\DEG�&��X���N�Ǣ��6���
�8���h*3jg�����-�n�i�<Q �+��=찗�N�	�����EAp��p�������������_���'8^l��g,qB��̄��J��w���F��^��v́_���0���A�*61#�-�H� 0"pB�X�'��*�6BP+��_L���Aa�<�gz�i�t��fN<���V�<��j����9U��[�&	��2���Hsf�q拂�6�l�G��D�ӫC����u3=|���B',t�P�ڞ/������R^L� �l�k <9fD�)�|�2d�vI�y�����������(p�S���K�=N��EԔ 	��ݵr�(��Q��k𹠦��)oػ |�K����,�9�t�	����O�pd���{�p�%N�R3�t:+i�lKeN��5z�2�r��G�}oͷ"^P>�*a�_��P�A�t}�9��dh;�E�\è�%���N��
��9�x)�ˊ��Vg���z:�Y�F�u��
Ӕ�3ș�v��e��_yX����D�M�!�)":U';8-If<Ժ��ec�bGm�px��:��<���:�V�mO*�j�I��_LI�
�\�$����a,�\��Ir���ߺ,������
��9�^�4:1�;�tJ��b�/�N1O��J!�\5�q�7��4�Z��5��n��ȓ7��*�J�1.S��Rh|MlT}�
�.�Աԫr�@��l�G�Ԁ�|F U�.!��  �X����)!����$�[����0�9�e��s ���@5�Mz���T� ��9Ș�'�t���Ad���D�����޹+'����w����b�!r�s5Of�vc麖��H�p���o2��l�o���e�V;�W΃`B^:,�9��s�:ʒ�{KM�����,>4��y��Ӕ

��*-�]�v�_qW��4�)��:���ݷ�����*^���y�m��w �)J~|P�l��1��P���VWqC��b�N��e���|
����]�v�AV�#;��!u\�Ӹ�4�B��m~�")m��,��i�,��Ɲ3y�P(��� Q�+Fڼ��[�����Kp,�LAɔ��-�x���{}�TTs.R�yK@����β��L+��=��J���_s}�@��+��S@F
�5'M���h���]WH�b�g���d�o����aT�׆5�T T���rRv,7C[@t�:2M�>���Z��)�!�m��@\�Җ24����	��f�թ��M�yz���Q�p������������ʴ��|xD��`���0v�1��R����n0GJ����H~ھ�n1S#��q7���9g��[�zl����fa�}��,Bb��m�q^�s����o9��8f�X|�����k�,LJ�j��
Yp�8�E��Lhge桛h`�Nj/�}(r��ůC�a?PCF�.4� _�`����į	~W��/�� �I��"_�@��h�ǽe��&O�)���+���g��ҩB�7Ǩ�L(�۽�^�����9l�v����f:nO1�|�Ag<9��cTI�Bl�p���.d��$d$[,���?�ƽ,�^����b�1{~�w(\U,��x��>�怑�0�jY����F�)C�ȷ��U��w��B��EE���t^��S��cʉ�h��|&��f�^S�(�lT����q�{3���rB�f	��,�Tk��n�ڶ
5L�o\�å��b8s#�4?0��D�JuL��vH��� �]��]��~
t�m_!����6 ��<�yY7����c�D?7�/�1�����O�0'��w���ـ��A9j�!�`�L��ݘ��W�$��GC��2�ci_�&/}z��OA��g�La?�ĭ�@�e�k�\�+�|1�o.���B���'��P�i�/󤂃�����}��S�q)_A�;��콬�~S9��Is��o@Y��V�л,zXi�Cg79��A=l� i:�PC��e_�cdDMV*a ,�s4@MI��;_B��+��ċ�с�G���]�<��f����֑#m�b�蹒/� -"��}����PKp�.�<������`f!(Hn3���л�k�ˬOd�.���۔��t��7�c;����z[#��M�Og����Ek��D�������o~\�+6���;jWq]���c=N҇=�rqҌK"���Z���Q�@���!�E���d���&��D��\�<��,}��E�R��P>��ؤ�a�H=�m9E��I�vt4
�<w���h��.�Yۖ��(��,Ly��;j���+y�� ��Dr`���n�����l��F	.��K�%�F��\�l�2�+������-.�{:"�s�Ĵ�%���n��{k���Ρ/����.�~{{QA�z��a��u�F`���f˩Sl�>�Ud�N�{R�8-]j�v�f�_.c�>	^C�B��S��������%?&A�Y��Ц�sa�׍�@O:C�qU��&ߤ��̠�8��ٚ�*o���
�
&�\ ti��h��j��W�^��~2��AXg�Xч�^كSOS4��^W��WF��W�iE�E�	�ME�Sݚ���)�;r>�M�($\��-�3Q��ל���>�'������?�ݞ&�(�5a�X3`}��ث��I�� Bh�����b�߇�+���9jؚ�Z3����<��|�� �*�|S���xrm_�?c�9�����+0f_+�+���4��	�+�P�������[��'�Q��E*(�m(1��Sw���ā��Z��1&�Ah�e#o��O,�-�d��Y/,����oK^ʬ0���$�^�ӡ�d@���-~9�R#���-�K{\E�� ?��zY�;�o�#����(u�%_�u.�㺩TA��Z���jF�&nq"ɇk�)
�y�@[����I���q�>��8��/�[!��ޘG�ʝo��!�_�g�n#~��䵴����Ԋ�8ϊ������Mv�n��m"�n�7z��vDx��Ln;���4��-{ۦ��ٿv����M�P�s�-Bp�=��M>z[\��P@H:6���:p��^}���ù�Y~��~���C=��'�S��g���p��Ѹ��a�uj&�]^����zQ��M#� c�Ikj5��*o�	��L��Ў�s�5��7����ʴy��P���՚�{΍$�Ⱥo�� ��欶Q�.��2;�����.�>����.��$7�����S���0.
I��hT�߀]FSL9��{�|�/g�PC���vf�(<C���.�iZ�;�dh������)Y�v��'A�U�U�L�3���y<��Jm���˘�o�f�����%� �@�����j鄝�>���X%����4S-Z 929*�ib��+��� p�������+q��Qm�d%���O��[� U���	���#������3q8�-��|�r�5U�xZ�:tB�M��>[
�O�Yu��ģ�o��u���M��r��{v�>83s8�Rw�����X���LՆ�����O��-s�P18ݶyl Ҝ}���zm��*;�$���7H�T�!���O�l`�`�-� Q3}��7 �F�]z�%��z�6��6̅��`c� ����G�'�'�z ]��PX�o^뎽ЬQ�yJvt�g�'0 ���*-�9Vq.�i槔�_:���uh�tL��$�/����wo���:��a�bx���<�\�H`)�ݙ�a�H��~Xj��]��/��u>[���!�� �0����a!��*�M���gX�1Zt�Ɂώ�A"��쭛Y뎤cjډ�Z�o���K<i��G}���B��w���8۩%9�YB�]�?`�E�AM�P]>
Ҝ�s}w�+B�4��'�M�k��Ǟf��Vb����Z�e�I#�}9zpt����w�b� �5�������/:���}��M�'>�����U\��]�\N�����D-vE��e\ru� Dw*��w��)&D�13�I��p�1Ga��>Xfz��e�$j �\���{F�oS�ژԙ�%X���O��pw������猊�3�Ǘ�J'���L���'7q���ހ�e{Fu��L�k�v*Cp�DW3r���k�7A���S`�����R���/����t�ˌ�*Z�hDm��q���n�R<�9�;�1����+s�-m&G~�,�+ݙ��r1D���yt[��-"+��C���qi��@�^R�:a�$P�'S5˱ݚ�n�F��;	�c�/H���~y�G��1k>Gے��ʲ���Q�AT��ea��;�vЈ2�"t�*�4n0�`F� }z�Kg:q~�Ȫ%� �#�:mj�T�����|N*�JS:�\c&�y��w�Ҁܩ���3<[��]���jL�jt�	�0��c��h��!jj��]�w�T�t!-� B��p�5��ʶ<*cQ�N�I�N�	���[jb䮐�3��f�@�4�;n.��K_,Vp��9#������)�Ӎ�Sϊ#�*�C̗T8���O��\�ǽ�=��/W��y�d~����������sų���c
ǂ7��3�8d�U���Ԙ|�Ղ��k��#��g�}�{���1T7��$:z�uAv�eMe�Mn���U.�
�_��I����Cݙ 	q*��
�Q���@x���P��<\���eIs�"}�e�"��t��_�v�F��t��'xxⓚC�}���}Ϋk�Tڙ�0����TF��q�'Y��A)� '���yv2_Ou��^�Vm��m��)7a�ؿ�<�f�Ò�<8hB���"IN���[��F^c�.G���<�8�'������,L�$&5��svXG{�\1w���]��=Pͩ_?�W[m�����DC���!��?�b̩@s%�6mf�1Nm~�n��F��Ӏ������l��EaX5�960�*|k�����{����V3�&=೺�O
��C��B���z���-.����md5��������M����z��R�ΒMrR#�=@i�^�yQ�΃����q�vA��@����zg	W�:k�Z�Shd�kY]�i| �p��1���V[�&J6m�$��+Ժ@ YA�{��g{�{�h�%sWy.�(������|���O�|ܱ�A�����ǣ`�����B���C9z1&��|,<��3�y�'ʳ��D��F�tWs��b�_j�0~~waې'�z�`�lg��� 0�'{q�1iu���o7|��;[-�	���L�_!o�^)o	G�KD9���AFB%'&���d�5ٴY��䳶��
l� ��!� �)�?][5��O
Lȳ��!�: ��1���AƢ��/��>90�y�e0>� U�{��l1d���C�ŧw��5�.ڍJ��,>:v�٣��0	j�]Kp�℉�C��z� j/U2� '�&3�v�4��F;��%}��2&֓������Z'�@��x���rl���� �=�q�Ƭ��Hk�$��x��Y `/��R��@���y�Cn��emN��b�։.:�E�*M�ze�2b �.	����M�N����U= �#B=>�#=�+�P���u`���#���أ�2�t6���zBz)�F3���NWh��+	@��8�UpYeA��*�}�FK
�Έ:���x.�m���{�esٓ��H�����OE��9�Q���úH�hN�,�*{咔�wYL.�(M�D���x\��߮�l]�MI�ڦ�I�z�$�*�h̵�Hk�&�t#0*g�j�^41du��Q��$T�y:_Ҁ���D�/O�׽j곸T�XH\~_�7��{P%njO�⤭(2�S��Z��Z$xǓ-��0���G����H�[+�ɢ��t�Zh��2f)?x�Q*{�qȔ�a�iZR�Z�pZ����t��,_ǘ"Q�4PU��[�q�W�[����LS$��+���e�����S4_�U�(��BcExy���a��#��Y7 ��Y �K��BWx ��e[F���	���c��iy�c�������OQп�c�@)yқ d��9���9^������@������H����UW��g�/�#b����5?Ge���c$	�>r1�=�/���;Ȓk�Ƙ�}Sm�(��2�Z|��:�<J+c���=�xM��o+��8�5@��2r�ŞM�RGw)%�;4�鰀��-Y0�\� b����Pk�Ōu�4�k�cC�"s��ϓ et�	�XU�� �l�.Чf�Cy��ʿ^���+C�M�;%�}N�n��$J�L6�c��Z�QP�8쳊<v���3��m��t���-�S�h�%�\#�8�-v ��t��O4�)�[�C-	~�`Bt�Q�b�A�;�����F�n�V�Zzno3M�2)���?��E,�m�����"��-j��!?0��Φ�*3u��4R�A�y�=?p�ǂn�u�S�m� �h�L���a�!��B�T�݇z�OJ�f>�p���3�ʳg�B��lm��^���x!*����G����&�G�2"��5����jJ�`h�����_��N���pUđ,�Yڿ��^B�Kg�U�(�<ہYd�~��P��k��Y��A"��ＰX^0�j�!����\�t8�>��5ό� $�0_�J����z{U��e�qwۚ�N�vl��rc��Uc��n�~e�-!~�-�ig��P�H��Ɛ��K��V�u%\�z�=|zt��������N����ta�ª���x���A�Љ�]N� �-�ѫ},�K-��'G��D��p���mJ�xJ���� ���O��5w�-t�4욽q0��-�����Y�:ˁt[��_ԛ����R!A�X��=V�4��:�m ��"��s>�iM
ׯ�Ic��W^�ު�+���a��7�w�ֲ[ߚ;��?��*�B O������b7z�y������鹿��c��σvr�\S!I�����eR����-�vs:ٛ#��H~y"~U�(�(� ��F0���p��l,îϜ���;1I�k`�C�}صW�se�.Z��|��X��GG�c�ڇ� :��DX;�]�b��`B>��K��Fj�-c/���ǍN`C-�%E��� ��.+��[�Υ4!iڕ��O9�[�2B�;m�_�3��o��D�0����u��R���l;v�nG�|q�	�F�ׇ**댼&��D}%� :jFt��R�3�yD��.�3үO������dօlZ,-@��b��ay<.k_ڂe)׊V��ZíM{w7�
S	$ʿ�%M�Ì!���ڰm���n�3VR	wv��O:��)���x���jb"Zo����
�>�d|�C�ѣ,�j �ugǌ�kf��Bk�}Mߨ��@����hw��G
x��G��Jg�����}}� 2m��`�~��z�K�(�N�3*K�pif���Cow�nR�5�JHs4B�夤��'UA�~�7����$�D�]њV�q�i���}��p�<�y4m����`�w���?n�졕iW��l� ����}�V�3V
��q��=���I�z�R�k�2) ?�e��b.L��|kx��E	.��켰�4f>+	[�,9����P9���~NT5$�%�>j3�b�����6����q0Xan����rE�9�,Y��
�҃3	2�Ύ������b�>`�[FX��3qa�ɾ���.����iL0�(��$���A���=�z�P�Dd�⬾q��7�>�����}��֘|#Rd�����񸹏��n'���,S�#�&���� &�h&���go�&�A���4�3��B\^i�x�ok>d�ߨ��X��;Ђ*�~Z��R]���O^�G%�?�jAe�z����&<Ґ$�ud�9��ˤ�����D8�|�֗ ����,���AM�
e�~�f��]U�L8VCU�(	��c��A���Q�O�*W~��o�`��>ɂ�X����A?t�L��`$�F��Ʃo�Ls�Q���:X��N83��ݲ���Ά�y��|'K��4��	�B�ʩ�.���;�1�k��t��XR~�+`cA��TʺC����z �5m2���C�p�]��ץ݌�Z��2���Im�p#�]�n+���?��$����҃�i���ia�����.���\u��Q��hd�el����
S�����ȡ�����eYp�|�T�qD4%ȇ'��3��-�g�y@X0������@�Ա�#Z���/�3Bg��a��4}������l��5�Ro���i�Bq��|�����V���N�tx�	2����7Gw���ټ�%��EøL�2	E	+&NfJ@�u��q��,�����R�<w��:�+�r�9�)�	��|��ٷL�ۗ��^�`�nQ�K?��xv�W�j���Z}���@�<�{_	f?�Iw����I׌}-�����O����L����d4�W����$M�?\_9�նN�pջz�c���2����ߡiZ�� ��£*O�fQ�/�#J�m>��TY�J�L-1gN�g��\��CQ�����L���S�
ȥ�$���d���)�O �x���L䧕�KS�|:�?��פ�T}�{E�&��K��JE�x�����Y�d�E-�;�����g=�@��dl��ngp
�UT�YTVy��)������K&x��8;<$u˿�*�0��?}V�4`f�z����ɟ��+���A���c���/[Õ>�L�/
��5O�@&6`.�6�9J	��O�蛃*ϰ�c�JL�Wd_�t3ē����4���>���X~�q(��K!V��vP;l���`ی��l}�SW���:�)q�fo)��"7_4�5ȶ�W��!#iD��t'��O��6v
�2Mh��҂ʯ��dI�~�������_���0~T�t�M���
KZ���`Qg+�	�$�Q�Se���m��o���fy�%?����������~��i�L�.�d$��c�&n;���Д���Hő�d�1ɨ��G�)��/0���9��u�r�ޚ�Zk)�i�A�8��g�CO��"5�F!Ʈ���+L����)�t������s�؇�po��Ǭ������S.4�Y��B :!'�c*���ؓ_��x_ %}Χ��7�	Q.�!�W�@����U_D�B�wA��6�gK�;�p�x{v��H��b d��k��(n덿��a��7�������d*W�a��>�+�]o4ȁ�6�uY�� �3���g��il�pg3g8�H,놯9^BS��W��Hu�������b��o�ke��H2���Uȩ`�e՜����
g���ƴ8���Z�:jL<1��r��\~��!IB��C0I�gx��n��"Č�n?}�����-:�`���.�j�F�qԼ92�ns�d��]/�y}H-�R!�e:ɒ��-nj�Ui��AgOc��M� ̗^��vt6<iճ(��1�ĢM�D��$	�ER���T��u�ʙ�@c�0[���"�A�,R��񍗵�өa�ʹU;U�q=�gOrS�8籕ׂbA�e�_�M�*(i�U��lk�V�r�2� K,Uk�(џ���N�<Ç^e�V�� �?N�����`1�e��4�tf�?��3���I#?#����MR7�L�r� q��l�Z�;�Q�u)E��ɏ{ejF��_'!g�lWJ	y ����:���gV���?H=�J�<w#�{�~{�;/�c�#L_�O�s"W���{�p��n�g�Y��u_��{���r�g�f�yO���f�������áiW�����|���+�L_���TZe.��O��f�I��L�Y��oc�No�a@�� #���Z��YM�7%Hһ�H�p����Y���6{}+�Y�$6J~%#�� J��k��֕Z������'�=�16����h�/!G^�yb��B���w©��Bbu&��R����ֲj\ƾ�[d�V�ͤ�9���.��t\��I�x�]%I��#8�Yv��3ճ���|R�q�$�4}��z7tW���y��� �u���=\L�d��c�o�n��#���)��qZgny�?4��i��C	�Ye�u
[)]X�I���`�o���ǀ�;chX5�e�&� /��������SdU�
1v�C���kO_QU�	Op<`�#Zu��&�gN��C��_��,V�L�!�@�����_�3y�U�銾WG�\iΆ�3C+�˟��ߚ��|}��yI��`��Z{���2��ԗ�Y_V������ԋ�L���?aH�{[�ݶ507�="�Ը,���j��6����A�?�}�e�#�����2�#g���Iq�4�l��U詎�:�bl�Q�ዚ��s�	������h�X�#^+p���d=��Ԉ�ϝVf�x9I�� u����[׺�ӯ��x��4��;����b���y?����;�f�O����b�yƻjƘ<����Dv��
I�c!�y	nv���2��K@0_���~���9��?/b��,>���
x���G`���^�^�p��#�p{a����F��׋L���KE��׍u<���XY�b6_Z���R���%P�3cn8p��ҕ"��co������������V�_]$�[~�1'ɰH�^�%�o`�#�����h�O�����_�b��)Pv�+�U���+�oX�&:)�G
z��޿���l�,#�ܓ�_�l�t�l7�`�K3,Z��mLX1\�)L9Ǳ�"��d��#��񡣘��)���$�3=#s�	�� ��3�Dz�v�X��GQʔ�qZ����!�7����M��M'*�˗�3r��W q����λ�(y5��y�!#�5���-�_TI2��	�
M {ck؞_���`�k�,��Q��a7'4�5���t�s�Λ���M8Ή�À[�)�U=��ݻ�x}���(���(�����@�#@�	�"f!w��lf���٬�:\��:}�N��1v�7�y�B�k?�FՓ`� �C�]�@�2_`��.���ؕ0;3�;�Z��m���W2��(��o{~]�T���E��)2z�!E�1�r5��N#3��&A�q�"M��Y��6����
�m��M!��V!O���Q5�n�Ѧ����+����	�֒Wz�"��yȠ��8��H|ױȷ�Q�!Rç;���}d		��M��L9��׏������U��|B���Yw����pG�դ����27bm���s_��˓{"��KA�w�6�u�����
Q�J�'|f��/� �>IA�B%��6#��ym�(�JYD��7�#�J�3�ߟQ@�Q�5�%�	��4VTR�#*�R ��
�Мc$��ɟ�����h�La	F��@bT�;|�0��:�y�+ct�R/.Ŕ��m1E��b$�gWݠ��/bm1`�Ña����b��m� p%�%{P�7�C�+Z$2��̵��v��@�]�Zy�#�Z)s�[,��g��q�05V;��5-pDYh[��^�&����➁1l�h�R�Y�(r|�b��}��$t	���� ��z�s?F�0Q�y�`��ǭ;@ ��7�6��#�� ��o9�J�_j��9]�2��P,|(�F�4�<#���u�rJ:T�����~��c�!����3�UY�Tfjj�۱,'R�b�������#���6K,�0��86�2�)4-yf��`�0Q����<ip$�嬠�нc�_���Set?2�0�Q�$�tI��,��'�9O�n�ap���8�r#�f>�ma��cM�`��s7@���Ь#��yh���"�c� h�yDZV�O��e��L-Rm�F������j��Q�fO�:��h�m 6 w�Y�r�]r��Ȋ��C�Գzӏ�fe��soU�Qc����/�myCTo�c��
�Bb /��A�'r��cmb9�Ks�jK�d"��om��]�DjE��׏�G�^X���_�N]���M j�o�7� ��8�,$* �Pb�c�W�vef���g�*�T2p�n��w��
A���T�l	�6}��͉�t�Gp5�z��N����翏R�{쳁�5ITTK{���:;�[Y�`����p�'�:^d�CȢ�S�y"�	�ʱ�t���V�L���Ї�(��������� �;�J�-@�k��υu!�f�q�������[��t$���y�bJ-
 �ڃp�l =���~�-%E����Rkh���QPQ�z���	�l�s�]���ϋ�`�+,ψ�з���^q�[=< ��&���$�T:��[7���op�Jv��m��1�"Q�J� �t�F�U�Н�����{�vC�x�N���̤<i�ӫy^.{���"��޶�ڞf)(NuueO˱�*\¹��J�J�B�3���)gT=^hc�PF=�Mn�����?�5�*V�	�1� %θ�؎��B��,�,oA�� �e��H�n���Td��4� ��.J@����c�|�>4�q��\et5��|6wU{"t���IZC��X���ܔ�qЃ��5�ޕCW������eiNY��"Z�_��h��>�]��yo^ܜn�G��}�J.����`Lv����ӹj����Ҩ�:�c4�����[&��P.�B�y�u���)���$�89XnHx{�����@����x� x<mEP�[1��2"͖Λ��uYaN2��^F��b�9������bj��"�Gqm�?�P: j��˟7�{FC�P�]b���Oi5����'M��>5�����z@���䷊Z�<�b�g�`<�tMX�j�FNzQr-`���NeT�8T�������U�ڂ�I�&:�9l��;>�s5�c���#1Gx���b�|�֞b�L0{9�����5�f�H��b$_�edy2�W��:Ң	�XY��0$?5�k2��g�ou�E���� �q>�ⳙ=$�!#?!�Yp��5o���c�Gx=�m}��x����}�x]RR-j�#Ɠ�Md7�W�6�+'�d}8WG|�&����%B:3���l�J�d�l������~Я%kƃ���^�sb�Y9P�c\��ʗC���|��B{���o΃��q˰�/�5�A)��a^ਵ��>bJ��h��p¢�a�>���d���uұo�?��d[��ϙ���f��z  *d�c�3��r��.v�5�5w6�c���'�BQbנH�6��4
�b���_4n��8z@���5�ڃ���J,>4W � ����@�6�~¢7B/��"[�������x���?��k�����
]q�O�����2L�}>�yY�}�
~y?�=���Őzc�ؠ�Eӯ�����I�VІ�¥Q��'C�fMb�|1Zd7Gw�x���?�ִu��x�ֱ�a���0�z��58����B�Hld�:_h�.���Վq� ��bFBo�{i���c��4����E7�Y�a��S�M�4�l��-g)n��롨��P���-ZJ/��F��%l�1�;_=i=,X9�s�.5�A&+�eh�|��y��0���8�x�������fē*�8�pL��+��m�H��(pb���]��0�h�E�ŀ`v
����E|�7��i��歽$�(|��3�^i׎��t�w�4�,��t����V�w�!&�r-�K����^_���Q�c�ӽ;�`�b�iǑq�ij%� ���2h�=O�eڳ��}��P�Z{ꎟ2
;*�B觕-��[h=5���s���e���	k�p/ �^����~ۢΫo��b.�b�~ ���z�֟1I���d��o	��.`��6�'����DŉY��� IBb�d��P�D)���YJ�Q���Mɯ�=��~��f���B���8�����[u��'�_ѱ[�%H�4�A��EJ� �-��l�uH$�풴���~rp&�-t��,�+~��݋�*��37e�1�-���j�G{^b�hE�d;]S�������Xb� T@�1�	��|L�H8�d&��������c����(:���,�G�b|��4������+�V�D�����o���b�7��|��3qߤ?�gT� �H��ˌ�E����CIc2i+�]�<Ѕ�9����7}���ȷ�B�!�sZ@ ��o����TI5��3(�f��[t}j{@����t~����֖�u�܀у�������߆x V$���,�q272�g� I2��≭H�ݲ�ο9�u�3�|Y1�W&O[ek�Y�7F�^���\.q;|��-��`#Xz������ �$(;�����v�f��@��켕�ZeO��o}���e�3)���~�+~/#[����~��I}(�l��t�4�q��IM(������5s{����׾-~���%Y��S�m������ �f�E�{0��g�J�ċ��}$��? ��v��^i<$���#�W'JOe���&�s����R{��3��l�~�x�Ē;�xn��?w���N/|�o�(q��2��?���i�=�Lta�.'�m�D=8��<�����nҩ)�n�73W��58��/Ų5����c��A2|cr��nG�1�-|�#g�~X��[2�dL9��s��ҹ-\���ZT��$���w�A�=��h�3���rNӻ��r�ԍ�I�J�݇��^�gU��޳v���V������!�ޮ��QX$]��0�^�Mkm9�͏�C��ٷ�}���b��>��H'���	dP)�T�&k�J�$��X
]��9؈��W����q��s�� ����.�.AK�AS��]V
��R[��o(P�$^��t��s�+^?�ą��X�A
K�����7�c��I7�0��s���V�
����f�v�"�)h[=��W���E�F�t�&�lR��nJo'}Bo�U��vX���#�o˻{!�k\b��c>�1��'A��~�ϓ��f��(e*cs��ϝ�4�����HQ��K0@҃���SK��'�!�כ��rA���=D�<��*�bvH*�N�%VY���ͷ�o����U� �SH�¤;�
��2���
��4�Ne{�i�=�ʆeN*��6:����`���;u���9R���MϏ��ϊ��D5�.>��؁�x���B�"�u����g�!�=Q�Ǒ�Lt::�M�}gǇ�7٭�"��"�Y�f�6��c��;w_�	��i��L܍k��CZ�OR��ҳ�+�c7�Y2o%�\���� ����y���kc:yϗ�<�6��������o��q��>�5���U�Z~%�t^�[�(b����*�e�B�9��_H�3a�����^�o�=�`���C��%�Q��	�N���h��zߎSX]�zq��)�I3Nψyӱ /[����|�h� ���|�|*��l�M_�@�h2��!<��X8��W���F
� ��dE���`���	6�BH�xQ�bR�5��������Ѳb��J3�fM3�J*H=㦄E�2�4(+	���)]p��%f;߮�O%��E�3�$�,�z����N4�M�o�N��wm�ԯOn���S��MZH��eМ����ӆ
y^���=� �.�#'���8A�<�Ϥ��D��%g�v3���b	�C�FK:���iUb2�#)pNs��
��&Wђs�i𝋶4;��+Ǳ�OG�x����GxIM��nƹdv���{HV�%�[?�v�0�Ƚ�������,�7CNxߍ�!��J����aZ��ğ� �`R
�=t��F�G��e7����G�x�_�P�=��j����F ����o��������ͫa���G�$��=Rh���}"x[
2?>�>���h��������t�K(�7L�<T�00������$9'����C�nL1�w��P��4o�q��B	>DE>�4b�@M{eC�)�]t�Q�u���EZ�d�{��ۉu���vM���[S��@���T�(׈�4%�:|��)�3���{�#s�V�a��K� ȋ���_�K���E�e��h���o��v/��(n�]u}#�<�
ۢ�#��`qƠ�s�fC�jc%��0��[�eL��e�Pկ�j3�7+8h��w�D�!
X{�}��IƐ�1R�\Q8q�]4��h�tEE|��'H�]M$�,�2��w� F�.����f���u��7�	�A"�_m}�D��2�R�]DN<�.`!`�@'����hEa��MJ��7d�Gb����W��\�>u�uv_�k�_T������Yұ�G����D��)갨��z~��VN��-~��M�^i����I��̷%�3��dwd�j��nZ�Љ57A5�\��Q#�&�"�mVD��]����UNgG?�Y��o�������0]��Ԛ���d{H����.Y�T
˪ţ<߄G�dxc������kx�Ggv���I3�wX�`#é�(�l���>�2��#9��#c�`|J�ʕ/{��0B#UW��1�y$���n`�W�����'��OqS���1��X��.QQ|�)G~���0/P_���{֌>�*�A��ax�w�����S�'� 뫲�&c'�߭E�L�D��G�<.$c�v��pl9:��Щ?�%3�K]hV�_BKЍ�Oth7��#̡��r=d�����ߨ$d���M�ud?٨֑�x�`���K�����x7%�HU\�<>aQ�!$soK�`��̒g�I{ �5�< �&��2d�e�8f����܅�[��g��Z�`���P�`j��Ӣ۽[�wj�n%�!���/�=�)Ab�y�J�{Ղ��Ƅ��q��Q(���X��ڀk�qP?3"��\(:�$��kD^��/[YW3�M9GFh��j��ܓ&�[�2�
�}w>�
҈Vf����TtV�9��߹}�����zѭU��C�}2�æ�1�B��KY���� Z�3��Dt��Y�1>v&8د�9�Q9d����+g��ir��p��l�nu��
%�ڡ5BY��O�%M�D �d�RaxZ�P��>��,��)?��=�m�EҜZ��ݾ��,���X��	��'R�$���c� ��k���Ϋ�6h�{��s�p�s/��I�5���_������zi�E��PX�2e�J�&w�XO}�ϓQ��@q�m��.U�ߟ�3f�'tV�%T�[~+��«���Q;�����7GJb�dW �k���;����P֔���:oA����O�����/8�@s��	{�C0�"G�� V_'P���b�#�	Ϊ�'u��w(A��x���{1�/��X���ڼ���k>ר�d7vTd�N������ܶ�3���I�Ǚj�팮M�=./`������Ș�2}��l���g���`����<�Srs5�+�\���^M�z1P�=��n�"2V��W�M&�o�ԾJ�~O�[wդ�4��Թ�E���Wx����V֏q9���y�ҩЎH��j8c�{����f9���ڃbm�s��5�=�1�=�B���2&��������x�-��C ���ۚ٣��������I���c�}QIWq�n��n��/���h�Z�S	�_L�2����F��+�J>Xu��m�rW>�EJ>2Sc�P����jq^��C�j�=4������nX2���3l*���x*I�����n6U�ɹV7�p���`lJm���^Z/��
{�$.�w#]�]\H��J
�ޙ�TUV䧴f�ܴ`w�1p�*��E1�xF�L$���îB�_�ăL��w��:ʢ��I���|��%|��:�ju�vW''×�p:{b�6�I%D��8Ğ��6⏒Zj�ڎf]%�;aآ�D�� D؏���X.�a���>F3�IS���t�D�[�2�5�������!8ΰ��Rf���S���.��Axh��4Rt�����nơɤokl���ھ.��@� 2��DaA3q����nݑ�)?7���X0dڷ]]���wu�Ɣ��MiJ�#�bѐf�/YB!ǭ�-�<�+����U���}��ykda0�L�Z�+Pp�z�g�8Z_�\j�?�D/Oj��X}�1�85w���g��:��%42R�Rb�\{� A*�%I�	���kk�Ȅ49�j�\Pk���_��p��$�r�޻?#*������W���E=�yg ��6�`S��˗��)Io�#Y{˪�P�]���뢊��].����\�6�C��ۤ&���Y���������h�YFV_�l�f��q\|����3!������$a��tiI���1���t|�_
��Ӏ'�2���Y(ӭ#
����Λ�����4�Շ�?6"��X����Y����lY�^x'���w�䪷K֑�ѭ��s)
�V2t`{�<�(��z'���?A/!�`�g�*��p	�d��:dd�6�4�0K��.I���XFW�(Msޡ�>�zPC�u`]e��gP�
���Mo��;��aT�!�E���t���F,�#I �/M~�2g˚ ��e�S����b�/	uP:���hj�J�]�׆�b��ŷ�e�I��P}�w>���T{�v�h�)C�΂����1i����#�6�Y,_B�2R���tk�ʋ�y-��� �/�	�j�r>����I��x�6���M�T�>F'M��H�Yu/���kS��zf!�0�ǰ1�r�&��G���jUJ"��z����pl���v7Yl�!t�K�<ӓ�5i�
�}����[ T�0Q��b�[(��ҽ����X��Hm�?�� �5']XT���CB��Q����&����,9%� �C!�R��V�ڽc���1$�#J����|QsT8��Ò^}M�֏��R�z�*���T58�(�~�U��L��>�ue��'�z*(� ���N�A8+d,\𧸔���ʺ�ffM�����߶��y�U�Uk-�z�p�iL,h�,�Nwٿ��?��p�R<p3F�ӱƓֆ\],��쨫6:0����+�Ƞ������:ñ�}��g�$te�^���˃Od����f(x��gk oU�8�U�0]�i�0�Y7���A���]s�h���9��^�[�?/�4�a���04"�iвh>���Y�J�I����4w��^��o/�1.�G/ɀ�a�2%�O[�����?k.�^US1��U2�9�}bR�}�D�"�nR'a��8���T�7�1��y���e�<��$�U��<3E����P��3x���N�����&̝T����B����!�yBA��H`rFwl��M�[5 wH5�ץ��<���#�E_/s����d��# M%��f�k>�@k2\	�A���i�#	���kH�Ԗz*s�P&e�((Q�ɔ4;|��n��٫/�-#�gG/��gs��u�\���g��eK��j����yЁ|w��c�"y�P���<��"ݍy�+��sK�p���G�������cwg~�	�1e����l�׈�^� �9��S4�:��W���E����RZ�M�=�
�B�����ӯW"�S?\	e��OT�:�+�����+B�r�ߐ�Cx�*���v�+�v���L+�2<��@��^��E=���J�X��!��
����>T�]���yR��������Q��C�õb*������%��&�k����߾����o��5���U���f��]tB{���⍭���#�R���AL��V�kG�E�G?���d��"|;� �\li�5�W��H�����i�L9�Y����R�"�?9!��|�2;�ٞ~1T���=!͜�.�!H�������;�t�o=��m�\ZHw���$��?��`nٛ��Ɛ��M����b0�N�}ʍ�k�&@F���UVr�_��}����I���W=d9�����f�.�'�2'}i4�J�<��}��HhڃE!S~'�Q �W'��W��Ĩ���M�$_H#��}\�q��b���r�?�F:j|
 )���]��#e��ƈ���p3!�~���k��R��E�%\^�I��jtj�==��8��} y)Zv�����G66f0�N�0�aY�_�4������ӓȈ�*6\��6j��'q�K("�y��w���H���3!딜y�6"�p��݀qŖ�0/�"6�������v����������5$E\�{�m/W�N�H'+�m9!��ш�Wh���jG���RI1�i߱�-�:!�=�o�3�h��y��Lz��|�O:� m�zEt6;d�A�sЙW���&B�f�K�)�#;�UI��$�7��g��5���}ڸ�$��86С�K�B�J�om^���X���&Q�#�L\/a�.��4�6�0\A�nR�h�jn�OA]s�xr�Ԥ�l ����Ga�>���Uj�h�s����nvX��]��R+D�v?v�k�D�?�u�-;��w1��`)�O��Yb��Χ
5"V%}h~i���ߝ0�\k|��_��Z��5�<�.N=s&[ ��ZD��p��S��N{�C�JU%��X���xm�m�+�N�@!7x�P��+�A�{�w�-�֬�?�� �B��]h��h� |g�i�#��1�޳{k�<��\R#�w��f��g��<1*��&��bU���X��+�7c>������v[;���tU�b`#�k�K\Q(�H����ξi��?�ܕ)���d�fg�mw>WE.L ڶ�+N 7��OU<N�D��]
���tA͌3��#vib;�&�I���d��b�t��|���x��5����b�/Q�E�|���	O	��'RU[��EV�z�N3���N��_�saZ����r�_����$9���h0�y��¯M-d��H+��-KEB�����0�;�J�6����",	>Q������V��^,��k�m��b�� ,2�G{N��r!Xrl~����b1������y�����(pi3��UO�P��zJGɨE�o���3��z���������}�j�/�/���Z��A_~��ŞI�&�b$5kO���D��?6U��q|�"�����a���a�G�86�rO�RJ���9�ZXi�x�\���Rf×��g�d�ˌ1�[�I-��W�ȶ\���X10LKY��ߓ�M���X�*�)N�m��F-0(��nua�6���CFY��п<�`3���'��Bo$o��p$"�!eK��c�^TVYnӽ��i�^�TM�5c�Is>{5�cb�j����y����a�|��p\�`��Ȍ_��YB�|�A.�+wB9I�|F^t���1M1�J:A%̀W���[�'y�����D�
ɴ��}LT-]]�L�����T��C�|��H������P!U��L�L1�����X\�+ŉ�s'}3Ĉ�lf�k|㔭��,�]G���_8���	>��������j�j�K��m]�0^\��!�z~�P��@#N�i2I��Jgk��/����e�� O)�<z�@����^�g������� �4����shEn���h14��-jk�v�$E���@ȚI\B�IaJ�e�y�w+��T�52�0��hZ$�q̡5ɺ�ի���'N�W��5ۯ�(�Ẉ�����x����Q��")B�	1`d�+��oB��lRq�=�Q<�.�y*���ǛX��`GL��%��j,N8���㯿Dm�~���?��%3��7�`�Bؐ���N�'�0	rv�����y��C��(ME�y�t���0��1uC�ΰ�+�:�GP�S`v,�(�y�|�@o�R�PJBB$�w����_��*�SǱ�D��Tb�M"ພ��<Ȱ��˔���MgdV>&q+�;�`���E`?��E4�K�++��{��j~�~D2�	����v�$&�O���ю�>�]�$]����9����K�e���a�� s��5�G}r��jO������A0�O��4��Ȍ�:3X^?� rd��خ�D+t����x촨D%�u�]Z�4�;8����6���Fˡ]�,�WrT6=�!�c�k��LD�y������:6+�)�=^���ܓ�d�]P��К�����F�$k�f	8\�㭷is$��r�F��,!�<�N�}��qI@�/��Ԛm5��j�e	�I(�������� �	-'n�����d!����e1#����4�qj9��\b1p�j}��*��^/5��X�$��:[|o3b�� g����rP6�²MMb
�K��=���C�+�ϸ��JިȥTG����+�8\^���Zr�7��	��t��̜a��	Xy�X���m1ܙ���`!I�2le���=<���F�r�����U��a����YIxo��w]��_�te����ꀭ�X���~Tgi�rk�]����o��c����rK_YxX}gqW�Y����/Ϙ ��55o���t�"�L��&5��ؒ�E	��@]����A��6�vA�Ge���=0)�m�~_�2g�d���ܲ��SI�ε�D�cM��������h`�X(T1)���_\jquG�R�]�t[�ͭ�d)I�`�~�r�`���}�C�H�1��DF�p��!xG�r����A7�}�̡T���#�f�@������s�;A`W]��|ĉ��G.�����xz�|���՘��%��X��!���P�x�z-#�V6�q�M2�-�`F�%�A1����
9!��KӼ>�$�/��dc��A��_,��i�*�η�=�;�zF�����D[.�O���|�K���K���Y�:�2]��nj 15B���ͻ�b���#3��^���{�����|���?.�]��y��3�:fI�|_��L�B<|rC�W�@�i�[7��Gx��0������v��C���M�b��V�ߜ��G�(g����F��Bl43 ���fC��+<^�$*�
���2p����B�558D_�m�:������m	���>O�8���e.�vo}by\�R�/;b�h�]�e�]s:fϥ����@ҭ�'��~� ���4���!��Nv$V#��;F��������3�8��:�,���}�E��Ue7���:3�y_��")o� �YF!C�g�>�4�F-��^���[���D���W�T�+�����F�݆3��b�3a��Ǽe͐����$���������m�m�ϟ�G.�VI���98η*�>%4�Z�^�R�����@iC�xW���G�~�u�*�߬&�����
����^>t�3��\�Y#��˽����>6\dSٵH3vE	�U/b�a	���	v�%���H�l4ᝡ�VL>�l�b)�Y����$.Zt<D�	e'�t -��5
:����y��d����w*~������x� ����ρ9����@�G�L3Kۥ?���d�蔷#� &�yf��W���S}�4�4j9R�>mu�<0����>�\J�	8J��/}�+Ipb@�-�,�z+�b��ra�<|/�U�M:��R*	�Xۊ��Y�i��n�/���O�1�2p�����H���9����@Sl�A�}���OU��b�!�=k���H6�q:訝�<O�ܵ����}t���`]2�/P� �$�f9?"��0�ZĞg<�;��c�lڰ���J�v��u]$F<��,4��:�;K/�Qǣ5 ���A>�d���`��3-�4�A淍�Y���7A�6��>�^ ���g󈁦��3i�k�h��,�Q�P˘/���S�r+]�߇o��̀��X�w�Di��-+IH�]�Ֆ�#������J��|���:�R��xP
%z~���~*����`�m4����� )��S�׼q�P��͛��c{����1�EJ[�#�u~�hx�~Yv����?z�o�_�b{n�\⺰����u�4�"��{��lP���	�����)�K���èL�-����`��<1��SX	L�-9ͨ]��0�X��ꥁ��q��'0����ê�UƏ���-��Q���j�}�h��h�q*��
���3(xN�ثz���X΄�z}ĕ|�i�
�"���kʐ���/��*{ .���jT� ��S��$PXALڠ�����7��Fh*2]Tد����ᾶ<]�M�9R���9��.<>������4B��C�_ܾ�b�L������ʗ�7Z�������;EU�Z�@��'���5����m�,:΢�ţ=R�A��� 6���5��Ó#�Uo	���N�<n���,	�Zue3�%Q�K����{�42��_�L�7�u.��Ä���h���r-59�(�R.s������=��U�/�:B�y���Ď��^�A$@�^�>�d��O�x��qUM�)��A�զ�����T�o�w��Y3���x\o��A� �4r��e;���za���
#�'k�S2n0 ��b�0���qR<>}w�iH_Un�M����R���?��D�ۭ,xT��B[�s�u]�kM�,�.��i⒡�Kt.�[�	�x��d� ���q�<O�Ņ�.�w��&3��Z&<?S�Q��\i�vJ��}!��8A!�4����f�T)���c.A��2d�����n�܋��9��'<^){��I�~S[v��S��U�o��1���`x�U�	�of����}�y�%ͣ���ؠ.�g����~�������~}�,П�E���ݰOu0�|$�|#�?
+7Є$cR�ZtU���X��G��ۑM�	�e�d:��^�� �u��&7�R(�������4�Cɦ��T�rd6�季�È�y�:C_!bDF�1�X�0|j�����'+���ʮ�ef�!_�u���Q��{��5b&꼳�m��JM?�$��R\E2Vaɕ玻�V�
��7ݦ\�p��0Rۖ:N�"o��y����P]p�C�>Wq5��RrW�M7��a��G4�t�hL�b' ��#{5.�Pt�V�_�?X@���&V�����%��NY{F�Sq��#S!��q�/5���鳔M�8QO�R-/�?ȕQH�Bb5%�f�^+�y���F]���d:�;���w¦�O�$�&��k��[��&A�������n�䐤!%��V��Lq̌���ڥU �=q�A��{���������9�`_�
��u��J���A �5����L_��-���g�Uz��Nk~����GSO`���'�����A�Xb�!����mwY�Ŭ;m�׬ԫP�F٪p�}a����U� _�6�`�Y^��N����� �dUxZ^�0O�Ȟ��U��l�0B濃Kt��`��Z��8St�����b���"%�	$�c%�ā��q����D��=N�Ԑ,��ꨥ3�c���L�q3u����DS����xo�����)3���8�-�B����e�����Z�P�\�C��-��g���[95j���}�>��,ōA]�8�B��:��Pw%�pd�.�eI��������q�~N� g��	�L����!�q�4��^DÆ*{3�B����bf&4 �2�$ W_(��h����I���2mhO�ȖhX��NG�=|P�v�-F�r�=C�F�@�cuk��V���B�ѯ~2�"�8/�rFV��G�U�_'��'����e8�X�Eq���H�z�۸1��;��@�-C�m~\��
�Tȁ�,	���}����w�e.y��#��Q��"�k����-�_�=�A�o��=�\����cӚ��X��O-�/���(Q�W&�<L�:���*�?{��U(�>l�s���#y�ዧڊtG�q�h�L�(�HWY��i�1������V�v�w�/|W���h�.��غ��¾�3#��l�N�$tS���0�~��$/b�,��8竰w`O�4����W��:*�KV)5]�Q�rM��JjW:��>DWna� k��r{�a���?h��Q#�谽S��9�"�?��wHJ�u������ʰ�$pQ�ɏ���6y�'���Ƒը(`5�2u��YNK�~�q��	���i5�qU�AZh;�zRC���^��㴳�z�2�>�A㉵7���c��j�n�QM��X)���g%)T!��H�b�@9$�{�v9�����ڶW�����R�k/I{*�TOl�ƕg����pf|eXr���
0�d�p���.���$e�8v�_}��SĘ�dJgCL;5w�V| ��^/+�x���L�NE�Sdp��"=��n���� �+̣ ��S�#5�V��������ThK#@�,��>�[�^�z��F�rhٝ:M5TAN@��c�2�@"a��!��E�Κ������%�l�}��+Sf�����j�z[�Õ[#�$h躀j��׾]�d�M�V5H pa����5.k��5���1��4A�`���V���(t�*��D��bb�h�3�#�a3A��`NB㨫,M��n�7q�^����l�%Q���m����f�-;vɏ�:j������'��3���5�!v�=��,"��&��c�^:@�>��{�����ޗ�^���|I�yr�<{�P�����M|�<��F�"'��=�2p�����B��MA�����:��!}��AS�;dj��@E�u�����H(a��H�9^���sA��/R���B]G�ZQ�/q�E�].ʖ���;y8d����X������ �t�	�#��h���	�30��z�A�>�~�s�
�E�3;����g��@d�"䐏B��1O'|">�D�����Jw�ei<�
T^_�\$[�&�ψ�f"ֲ���h�(�{>��������D~����~�IԙH�t#0�	�*����L�����^QE�j����l���6�P�R��RAsNgSve�K�8yV���;�8���w���pz�F�6g?1.��;&uY#���PR�]��w��<H�7%��R�w�w���F���)�UMߒ��=L}Z�����s/Ic�h��XQ�@�߈�'��/6wd(�L)�|�-���f-.ݓŌW�ؓ���%B����%�@����lX�5 �����g����ڤ,m���r̚���̃6���Jg���1ԟZca�Mk[�*$��Ro^E�Gإ����[�"��LS�w�֦��hWY?���1b���������N� hf$X !�nV'��&�g�E����-�z�7D/�B�:��^y�}כ���Z�\7�@=���x/�FkP�$���k�
���� >��� 
�tCO1lǭ���Q8��	�)��:{S�2�����OF?p�r�i>��.:�UdgN���9��s�Mh9��
�OL"� mM"!���g�O< ��~Ә��/U����N�C�R�~a�.�7���\��v�F>�M�<��(��a�{�)2�^k���m~����w�q�w�N��h��M��ߵ)�\�F�����b:2?��T� J��?��Ok�o�����*س�=i >e���&��l-��0�aҾk���$�'\� �jk=뚒B������mH-"�TZ�I�H�@~�����?q��
󶭓��CE8ڥ�qa���^�f��t`x��r����V��w��R�C;b��s�wf���rj$�,2b�=�k��-��,p��Ӄ�8���d��&8�F2�a�S)@Lz.!�@���(����j�X�4|C1�q�����cXA���0�{iR��d���"�f��pW�#m�g�2q�es$��z�K���ZMp渇MECH0��sJ�H�!�`����%�H��j�[�\�x�\|��1�g�Vڼ���ή���w!� ��Q����uP��ڍ���TR�g�:�n���l�S�]i�2�qmƚ��\�*�zF�d���Z7�i�.+;g峳��'@"�����J
\[������k<W����٣C�[1Z��`�z��>���W�֜���n�2���u����32$1�-��)�6UXSRg�[g�ޘ�d�Q�Г"��]U:FL���I����hz$(�h��,:���l>���/y�B/#�����4^�E�eҠ;���@�qG٥��ɚ�,����"�������^}]6�ھ�
P���#�8��=h�a�I�U*��ԅw*�O��܊d%C�s\�������a�t8�k��Gٰ�H�p�q�֊��|)���N���L�\'<X�Ƙ�V6��>>�qF�w�p�n����~+�D١N��w�x������|T�=��tt"w]V���V2�Z{���XIu�B��Ӿ����cq�8��I�rV7Xc+u�n��TOU����5�g�;;#������vԬ"��p�$��2�!��E���IQH��X�Z$��S8��+#+�F���md�F E~~˥:�hf���P�}(����w��HK+����m�.&ƨd�S�<��i�֗԰�
uL��Z�+���J���f~�?���R�@]�:�O�I���#t���A� ���B_���L�U��Q�g�ht8�d�}�l�<���}�G���4���s��^�H�o?8����o�?�Y� Q����X�몂��d�F��^�*����YJ?84Lt]P�����������Ŝ�!�ʋ.s����(��nB+�P�%�s�"�r �ɬ�t��N�"8�Z�&��,�x��^�vm�@�^ی�W������O��y�''^h�I��'�� |���u߯	�M&霛+��P���O͜5r��mAd�N���bn�eP9[6��>���y���0�	s�������[�"���@1�)n'o8�2�e�G�F��յTx��	>>�`@J^��r�Oim��׸�&^�.�Z:�
XuK�s��QP�UF29��/M�C��G�۲64���o��%]���M^\���Ѥ+�QR9쀄��x��C�*�+��:�$�'\Ɔ�]��6E���?��T��Mg
yj�d��b��0���M_�D߻�GL=��f��a��}��D��7�} ����5�F��&^��l��S��Lt��U8�LBJ���V���t�B����aȮ4�uuF���o��K��`B��M&���/����<r�%-�k�,L�*Êgc%���!��_v���Av�"zZ����V��n!:��v��ro�����Z�p�i��cr��7"����P揀5奓::'�G0}<��!�W�=��ϩRP�pY��V0-�����#|y
��v�4��m�%c7#�NW�J�PlDE�7�\�z ��O���H�Z�����Yt99!8.�ں�[��Ӊ�nb$���1p�D���1X5�to�P��uB��@����]m�
7繘�]Z_�JcAL�l@�	v*v�W"`�n�|�թ��楙�n���K��F�+"c$� V�/݊�ܾ����������G?Cq �U���d��\�_Qâ�*��5�ĳE�)���F1͚r�3ݰ�(��Q�h�WU�:���dB�8��!����v�kd6�9g$3�n�A��`�)_��0�$kPs�4�#
��A�j��w�[|��x�Ǌ�������B���Y���}2�_*ۄ����W�k�I��|��nf�ӱX��1-Kb�p�֋*݋�����̮t��d��pn�y���v�U͊���h�uW9DA!���,�B��� ���4sQ�t��SM0Q �����e�O$�˅���9�[l�w'��Z��V�����eFp����@�a�"�"��Ȍ��D9�[.!�Z�R'���Q3\ޅ���m+��2��3GoJ���5���o���i�&��(�t�,p�ױҢFF|����(�:*Da�r2��}���	3�8�|m��4B�0�fc����A�tL�ՋCi&��cG�w*�3QgB��s�.��OZ�h�@��I�X�TɸJs1�k��Ń��m����l໮����p<�7�P�,|��}#tp8j���琕j� � ��V�ct�+�����*t�p�Y���a���\?�XN�5�U�J�B���Kmq	���XH���_R�'\�mE>� A�	WK�o��FLw��z��1C]�$��5P+�����:;�!��ɃY��Fx>Ԛ�od���U��i��ZqC��U�2x1w�`g�"� �q�} �;Yܨj�~ ��;G�c�ߜ��	���a��Q�Hi~t[h��!��W��:k�F��s;]3.diڜ�j�X��yag:z~���P}Ո=�p_R�V���e�C#(��?����G�|<9\C.Z����î�D�,	��[�s4�In�#<��K-�7޻$��lz|ЊhͰ�|ۢ�f�4�K���L�Ł�;32N��/���4$@zpw{�a4������G����]��h���ѕ��&XB���6j8���f��x4F��<R��^$x�Sf��r7䑸=�
��I�7��K=�|���<�{�,���ٻz�|�^���مxezC�"�IhĐ4r����'�O9�\�CX	Vnz�?Ë���*ݺ�yo�v&e�܀�ܘ�g������_�pE~�^���m6u禨7��������
!]�M��+����ݿ��Y�g�C�h��$�J��cu�~���KP����iG�k�*�	)�]��#斞��4�iP��V���?�����5D[_&e�En��a��˅"�q:���:��E�I�I�53�����DyӐE��5lC�_ۗ��M�b,�?H�D�[J�-���\�'�� ��9���S�1β�2|�i�d(���~ ��U�ǒJ�t�Eά&�޿I��8R�8D�}=�+!Pz�&���/��3!�{VwQ���J�����2��S���� ŉ:,//�7�)�
�S��)�"m�4n2@m���7�V�W�I�$�q�Au�s��\aF8j�5n{�,E6�w��7�|��'`� �-��$*t0M)���P@g���5�(����ruōwK�݂}l_<�6�&��s��>X��\��ޞ�J�~�,����kj��j�����W ����Umw�s��ɹ2�ބ>�vm��c�&;?ɭ�߭j�� ���#"��5�sË
�}Z��n�-��(��iP-c�#�I�Ĝۛ���*w�iCQ�ëMr��ﲀE�D���as�յrE��<x9r5��;�pK+H3�9�D�n�8`q�<-����}.�v,��m]M!��SYq$� ��tcݖ���3<��?�pڄ�+���с��DZ�!�?W͇2�Pi^`���-�����������A�'��[a��k�p����O;�d̨}�� �;�M��m� �9�K�,���+��TTY�+u핂��>;U��t0bӦ��"�Ƞ���)��	�F���6��1�ד��K�)�n�@P�� P�9+}߶ ��Z߄-H�����D2.�[R�#�%{}�bk3Y_h�(�}R��X�>.�4N�T���r ���6W��4���4J��#��I;wZ�����'�1�؈-�w�s��D�\=�<f׵B8�S����0fXH)3��h4t��{0z2%����%EȪT��/W~�ܶй�:
����h/��C֮*�xË��I4P����$���L�� ���/SU
|�ڋ��P�#�YAn���ȟ>$"(E���5�OK�a���i��$�FO�:rT����L�i;��\	�3�*�9T3��5�6�n��/�.}�ܪ�i9��l��e�"ü���WҚH�2�AVj$@��n�JS��8q1���a������]�(a��X�7�.��O���t���7�AQK�ӾZWA 7v�_�^?�-��H�V5��5R�>"������?Ҥ{��L�y}��>{
��31]��#7$N�빩�/$Ni;ܒm!�`��h��յt��}�,�~�����������po`��*�������)��sW��������.'����w�����g��C
~�* �ώ�`4�G�ɻ�����2ۓ(��U����@��,`��Hh�itC����
0Z���+����kÑ���VD"�-k��8�F��`��|WM�N瘤�'�<T�tqQqעpK��^��N�����8����~뙖��k�w�<�溿+-�ϋ9�\��%��=Lh%�-X�JW�q)lX��?S&\����E�껇e�I��t�Go��]���Dѐ3,�V�y��1Va���]Y�`Q%{h�9v�9��G���I���\��u��0��c�ev/�3�'�ro�U�1��P�^ˈ�\��
�b��C�Q?������E1�< �����ޯ��k���Ǜrj�T٬�XI
���3ɶ#65x�Ц��T-{�a؄-�w��7_�fe��KO���Yt&�[�e��[�VV����<Ud�������I��΂�\v�A����3D�.�
��s�#�
rI���J�)�a���Id�_lJ}Oy�����'�r��<�j	������^�B��e�zm��F�	@i�k��q��V���`�L�r0x#�nssʙ`ȫƤ��j���ۍQ��{����K��b��?C��%c���w<.I�l&㹪O�Xi��{T��Cy3�Y�b���=��_��vn1J�8�`���e9�P�9�r�s���� ��>
Ҥ?{&��<�b�T�k�'���e�nZT����E����p�
Y0�,#;���2/�.pu���^7�뙝�ȋ�Jq�W�bk}ߢ���GM�7���:�+�3�E�X!���V�2V �{&�"]�VG���z�X1H��E���geҘw?���Ig�2a�S�;��胗d���%��BY��1aW�]y��͸�:dbk��җ�뤒�'VR�R��Bɸ�"s1�]��7�7�*$�$y0���4sj�p�{�Ѡ�T�>���d�����6��qvQ{��8wU����q��.{��k�Kz�.�KӞ|������9(b��`��WR(��7����e�'xY.zv�}���[?E������_&YJV������(Et��c�v�kxPm��zm���f ǰ��7��@m�萉'Y?�j��J�(C�0�C�2�-[����JEđ���5�k���~��$�鹏�K(]�߉�X9u���>�m�f4~������@�ʘ�/.������{��z���Q/�1k��NaZ�����&�(��b�GME�G��Є�M��F�߿�
̮�Oq��5X,�漕��ʝm��]o�C�$ጮ*]:Nh"UQ��N���S�)��\񞶯�N�2}��9;-�l�\��K�޳4���0�48��*�d��Dz�FJÈ����W��<&���R�,[wt5%h�� ��'��A�zg��5M�7i	�{g���]l�]���3xbʍ��1��iiੰ]H��N4I�!s���
^՞C"q�~~ggk=z�"$�+c��uL����o��=�r���Į��[t��Bpq�:V�_��@L�u�������?���X�x[�WZq�����x~O5	�ސ7��zB��/� J~�� b�/[Lj��IJ^8���MWl�ɭM� m�{g�� /���$5%hN4.��V����	��^2ͫ�"92��~5�%�fqC�_���A+��̂��ғ����~�G\!�q�߀#Nj|q��_����z!c�UQ'�U��H� ��Ҙ��*�uK��-ʨ�5�.;�]��]e��,u*�`#���±b��t���ŐkE��Ԇi}U�#C�Si�c��+���i����~�~��g����vA
��P�&��v0��0gK���dx!��$C��f��MWw5f5���
	��Oر��	qt�9p��Wi��t	^��J�abV�z�ⱪi'!����+!<�,|�J@K�n�+.|�} �h��ӹ�N���iH���$)İ�?y_8������ި�Q� AI4f(�>q���}�X
L{4���0��=��ޗ[J쮭.��g?�V�M�Ga��9[�V��w�1�=�o�E*���v��!���'vQ{�46�Tv��%�nH�	c#+������4�V�E�0V��F���,��#�����>m���<��wE�$����K_+���$�؎���y�l��tO��&��5`uP��8h��d�$��x��2����%�F�X�1G�oR�� '�ї��"�n���M�Vݱ��X�w(�%ta��w���
�a��j�cm�@�D�`��V�=>�:�3jvތ�ߪ\?�n���	x��[9���?�g�\�T�>��
�;�
r,� ��@�w��\IOܕ*��4nW��_Qg��%�b͆	��/t��L�M�u?g��S1hm3;=�\��&Wu�|[֋�}��%4��՚��u読,�0� �% UA 	��)WP��2��Q���NSx˶2|�b^����W�R4�ͧ�%��V���a�Y C���������F_/��S(U�pΣ��Gpb��y'��>+x0�!��X�V=d8�����H�E.��Ǘ��Ys���^��!nj��){��Ȩ���Μ��g�`Qb[1���W9}+/��E�9%w0�z^�=�-�B7��9<d౺��U�M��Uz�����W�Q�i�v /l���ф'�p:�P�Ի��p%���Q\<����Z�e�!t!�fS06��" omٝ��P7�[\x� �T�+t{Y@�m %LC�q3�^% ��dX���+�~lq����b�!K���'O�~|'�=s��Й!�r~ ;��k8*5x@}r��a6���rХ�E�d��~I����ڬ�;_^��·`ג͊]A�{�w��ؾt��Z���H<COhҳ�̀m��#�����g�����mG�(��"e��{>���Ԍ�X��8����ȍ�����,�7Z ��F��s]d�xUȧ'^ShV���؎
���ξ�x�4[����k.�f��V^�*W䵐�I�M)�D��.F��o^�rDc��<_�xZ�9w� ���y/������=�"��hE�o]B>�|#ۯ��m1��6r�y�$���ֈ��9�^�v�r�c�&v����.��ک���t;�����0��ӄy g� 	,ߠ�P��zPO$q���Mm���H8I`��d��	x�#osPL��P���o�z5�փ���hd�wd�ilJ.eG�R�Z�`4��B�F��>���rGQ�Ɇ�D�%�Y��4�{,�8*�U?3���G
������5��k� .bL�$M�������?�=eȅ<bx� -�S�!#��ᕞE�Y�y�1��O[�l1k���T ���cz���bY1��3���]*����������+� �ǥ���V|@�ӗ��xHٹf{�p�s,��K��\<͵�%y�z_Y>�\�h�, 47q�zD���N��`{u��4��mb��h孱~P�&�b�4��A��Q��TS�v�����W��bqE��1&�� ���E�s�Z����zT�5G��V6�M�'���C�x;O�8��=-;vz%4�	C-hg��D��Odh_RF�W{|�;h}L9s�%-����H������ _����DƓ�z�B��t��c�RY%սw�&��}�쀻	ܠj�';i;{U3V�� � {�)łPS5��;��� �]c��Qg��1�l�+H�9r>y]0n�Aݼ6v����y�?S5Z��֎p�M�R�ưhS�����tV+��]ۜJ���֓E�aNA��'/�ɪC䡅���B;�X#�0�=�:�:d��q˹f��S�I�ɒ��Q]JMӁ�Tŀ�L*�7æ�]0Ͷb�SE�l�X��i8c��Z�)`z4�6�� l2���-"�+�`\ϊ�
~RQ;���U'�6�E5l4B�Ur�x���A��Ӧ�G�:�6 R
���ׇ(���Ȥ��_��S��Zv��{!�K�.�偯OBE_������ڧ��}]��GqYR
@�1�hCE���{��D�|T�1�6:j3rB�ɷmWV��8(R|X�:(s�������$n�=?m�=5�T����H)�)��)�sJE0ډ����(��&ߵ�'�h�q�h�>.�h�;"1�C�0#�Z�lC����dJ��M�^���3ݜ��b�k�������0��1��A��WH�c�N;�������l5�q���GS˻5;�ǟ
�喟��P�	f�����&�W�wϮ&�<�k�.�<��E�E�L�Vfi�L�>��YHo�Ʒ�ܦ��2]�ܐ�L������bc�u���g^`Ha�ku\�>�@Z�c�^��P�D/�'�t���b�B��4k��y���ւ��t�Y�!jw$Y�}�9�^������ʚ��*�A���x���E	�:[�"]��@ݵ����ﵒ��4��:���;�����,�STw�Q���q�0��!j��>�0�
��Z����,\�} ��UZ��G�L��g�bi��b~�h�n?6��p��Z���z�M�c�w�zS �7�K1�xk���ʨ�7��Zk�+
�挻�d��"����!�"♣Ӣ�]2p�h�6# k��pJ4-Q��7�7�Uu���)�>�×R������7�¹Q���T6��9�Q��p�>$��?��W���,���|L�7�\KG���
����#Ń�z�f R�s�/�YynΆTz1�L�o_�
��=:TZb g�mn�Q�Q�ٽPW��y _�LVt{�z@0tC������$HM��A�����Uhi�������^�V_Ai'�J�^H�?]���~"�|z?��M���y����+}�ݱss4a�� ��Y�����BV�`��o|��	ZYwp���g��t��a"�� *���a���L���H��ҧ���Hѓ&)���,,��7G�
m�և)��V�@����\�dؾ��5���\�b���
�iξ �z�*ՙ���٠K HP�2�L��e��UW����+���d�[�]�9�{�����7�ۡ���;�\ۙTo`�Hsj����QPr�����O!0~�/�E�ౕ��Ҽ�
MۭUi�`P8�i�l<|ފf.�����!y��r�3�~��B. �v��ũ�G8��%t�-�t��]7�A1���v�+$���;S�h�XB]1�fׇ׊��X2�[L{����$�n�{��:��5]���m���~P`�p�z���V:f�6��p'���c�o���k5}ĉ75�i�+o�R��˕�8+l��*��4���F	I�]�M��]=����>x2�HL�1e����V�ȴH!�Ō�]onn
���^Dn����KQtƉM�u�����]�o�ۧ�H�pBd�j�)t"��`{�����J�-�� 3;%n%�!ݐ~�@[�a����*���&�u}`R5��ui������g[T����۟>��������o� �l�
�r5�B)���|3�W(����+0;8�<�I
�|K�~i�JL�F_��ɭ��
[�:e�Fi/�?�:����PӋA����2��,:�a������bڥJ� ba��D[��J�C\���!b�(�"��j#��U��OO�)$1�XY�b��:<��+���{0BIi�,���W�d+-B�������H��
���'T���^�~�y�h�����E]|����ЛrOL���Q&	��;H����C�dp0l�C8����;��D��a����>�Լx���$�c��FQ�9��d{�5R2j���Nv��>��9������ֈ�gTs;SW	�5P�߄ZO��Bȵķ����}"t<��;ۏ�U����t����!���g�ּca��;��pb�r��u�z3�n�b�86�j�O�j�����c��	� ���t�)�G�q��7����Jw+䳅k^F�}>��T��ҽ�҈K���u"��lv۬���X���A���Hk��rey��w��+���Z:�b�J�Vak���M+y�l$u�,?��t�z�El��@E��i�>e��ʊ��Y�K�{��z�1p�()\͒fʭ��J�ռu�A�f2|��&"����K�qz�!�5�h~sĜ��z����]=`��H��/�ė��,�c�q+͸��y��l}��g�-��MY�|m����0{�r��j�����x����HB����<�_k�g�o��p�S�u~��a[�72+�U�\"�u"^�h��8)u3����p�{O���KJ��uz0C��N��eW�|ys��
+HK�yI!�-XH�p	a�}V��h���9�z�m�B򌹽(A<��}�b�c}+$������-�9a�L����4bq�A}W�����,��4�����K��7��c��it��(v �ڧ�3ݏ ^����
���Q��k�A��F��a)�����I�
siI-ά��jK�ӢN6%��֮x�z���S:�cV�"��ˇ�)u�	?LK��u`�,�!���0�u�g��uY�8�:޸�-S��ت�R؏L� ~�na�]U���Z��o:���}�˭
��/�8�ݠ]�F��su���)�:U�`���K���Ԣ��k�Hto����xփ�k���x���u<<`^♡ré����.;;������3�}�ա����me�P1$Y��) �]Y�JR�VEϯ>[���y��P�x;���`s��(��2��B���W?�a�"�h�^�+儧���bvn�y�J��2@�+y��og:Tn��t���$��%]�%�	�L��P�9����qm�>rV�9z�F�w�{'N� {����@��+c�K0�;�Ǭ��� �C���j�8L���7��k�0������j���_�����az�4�*���k�(o�P4Er��!N�X̚k��h
��~	�1��ʐ�,���(�q�9�yNN �A���\`H��%�ٮ�1�^��oG�9�h��fl6� �Թ>�=q� KWA��X����0c�a��x��Z���O����i�cNq�T�+�F�צ�5`:���!՝d���րnﰪ�)<���'P�S�n�]�67�X�T,ĩ�����v�p�����5ï �˗j�sF�ȳ/��x�����1�0k� �۹
m�n�{�n5�A0��*x"�4��7i������������{�u��T^����2g�UK���:�aZ��Uin�'������gS�"�~?���Ǚy�J��M6�����ڡ�����G^T>N�p���?��n��ؤMr ���5K�~��^��$�!�-M1�i��nK�t���)Me��6���-Z���TQν]a5���-�n��`k5$���1*t���.�*�Ϫ:j�#)py�8���>Z��C�[a(��ء�b!�sr,J��L��i�����L.�	�D�V����=o]��?v]�N}�y��1H�a�8޼�^�ԙ./��{�A��Yd짒������<�is(����=�sj��g0P*dٟ����r���i�g5���@|��Fygť�4��^F�	*ڃ�.T3#"BС��e�i]�����ǥ�أ��%�Pk���0S�ڥ3��z�@my�雇ҷI՝oD:���0�ϖU6�����s)5*'^	/S�i@
EU�2#��/��0A��!���[p�Y�rl�Q$��%w�֢�#8(��8Q��*lf&�Ĉ����/)+�7T�|����O^g�ҹ����ϔ�Mv�o��
��,��ٸog0J�D*~�nhP��"�Dl��oz��L�1A��l҅�
[3��.���7u�5�Z�X*d�s~3X�ѧo��Xu�O+gl�g����`B5$S�E���K�(w��%���4+�h�[_��R���b%f^�l���^�q�h��R��^�TR�� 4��?�z;�̘�ʫ�'������Ї�'0�=L�e�����`��e����lQc��� ��5�qlV�}
�cŶPU��W�/�="���+���U[�u��z�d�P#����q�k�@di����2TNUu�?s�O�mzedB7�̙ݛ'j.�H��Ȓ�gN���VQ�:L<�P��ܓmY/^�8g�[�$-���t@��aaN� ��� ��dwwo��ћA�׏�/��)�eU�I�^{<[�8,Ւ����ѭ4�!i�����$1<�Ő\\c ��)i��z���oS���f��ԉ�$��vD�ݵ@W&�̊�X�< )oX�ȕ��Vm��0��C�q���r��Jy�,�x4�?��=>;ya����$��^� �n�JA��;Q�[�0�:%F���!ʞM<�+9\��v��4Ȍ1���4�;A�3ť�sx�E֢L����U.h�I�֍x��w�~
���L�#�� ̌���U�m0���q��f&�j�4_\Pr����q8ʐO��{�G͈!|�^C��|���?��9z��Q���)~�w&�����/��s�����s���2QI�%������W���%��Tܓ�
n�%��_�uP�sE� �\��-�v��U6`:��녑�}��iڠ��0(-B����<7xZ ��b�&Ҧj����}<��ZTS���zZY�n�&�m��R�c-����#��F~m�`�x�hN�ߠ ӣ�}y�����|*��i�4N�><T�`\qR̝q��H~E�'�7d[e���en1妆AC�ڤ�-�5��@�b2���'@v����߉w�dLa�-(�gL��$jK����ā�����G��?�r�����}�Xa@J�; �T�Om��]T[���<<�wM6�����d0���}���ɧK�[���Lڢ���1q�]��G���{����`F)�J������*-�W��^���X�!r���U҄5Q?d�r��L��R#_|P��E��0.ۊ�{ԥU0�HO�rA4�H��o�̟��/{ҍ�p��K�����$�S5�h�e6=h�c�fv���������6�{Ǵ]v�F�a���= P3����4�߯�P��?�X�2��#8V,���#G�.�3^Ž�,�MMsT'���@�ɼ��*���%�#3�Ϙ�}�%��ue��buQ3;�����fψd���uZ8TgGN���� }~n�4�x����7K�-��aG���s��ڙ:����>^�v����D�STR��,/p �� ��YS���*�H�a�<�	R�/�7!��x;w�'�9��Ңv��搞�^BJ!�@���?H�A�����o�������$ 6y��3��eF�д�o~�t##	��1�7�ײgH�sV�&��0ҍvO:'+8���Y�cioo���:�!ğ67����G��to���j�8����|�SѼF� ���W;	��g����g�:y�.<�f#-��L�����N��G[����K;E�*z�ZC�Q<Wk���J/�L�.�4R~|C�}�Ҧr#9ъ&I� ����o�yu!ټ}f�x����(3S�$u��<�(lʉ��:�v�V_3�+�2�%�E�*k\p�3����`d��,�m@j4�+�฾v��RBT	ʹ�/7�*�^^�6����h�_�ٺ6��������A��1�d������D4GS��(!�7ᠸCx��dH����r12�A2��:�.���xB�M]�֋,)�(��o%𝋀�)���N,,�0ju�a�Y��N8c9���˓��	&D��u�Y�;bK�N,?=�����V�/�y�ۧc.���TZ�K�9} �Up���c���Wʾ3Cs	*�ӧ��Q?i��`5�2?�Lb�)5G�J��o4НuN�X�6��5q��z�^�����I�g�HLM�P)"��􁷚��*W�:���Xӵd�w�` T瞐���ș�hP����Hv"�eǞ��,�!Ӌ:�v�O����.|\!J$;O�K;�*;1u�1��EM聕I_\��5h¢ ~�Ҟ�ai o��-�R���X��
B+K�v6�E���u�t+3+>a�2�)Ff�$zޡ, ׈�E���aP�����U�j5���'[����K�!���qp�2��h�b���,ƭq6͑���u��Jc�/�N/�ui�塪�'0
����b�gw����o�64o?�&�H�����R�YI8L7Wuq�U,�5YSY���,�Ϫ�K�����>ӳG�fԧ�$-wLP�qR�<�.��r�U���E�|�W�i��QY�ݱJ)	1�bT��-3��#,I}}�0�#p>�N+1p�yA?��-5e~���7X��b���9;)��_�1���Ja�(�
`��7�YN�.9FEb?~�pё�>'�V�0N3$Ø�= }���;�i�OEz1�W��d���a6Bڪ�J�� E�-��g��R�M��S��	e\�C���4d+�[��3WW�4��^ �5 , }����SY���WlW�(����o:�HX�ӫ��%��J��G?�d{|b���ʾI̐S� 0�Φ��.�-ߢD���G����q	�X��^�*I��Y�u1c�g�J���sz�.4s��u5XN�cX�3��/��P�_�j洱����ۻ4�*���}�������P�J�䤨�IΏk*�Ҏn�����9% �hx:�����A`���Dg�����;ϩ�/E����9[�D+��p>��a��������7�V�L%�ad���^�SCf!f�TK�l������y���@�#����y�փ�2_@v�=�-N��i���p>r#>ٺJ <�oVF�|gaI�:�:��UA��8_��K|��{Ln��u��ԡ�Î�/) ;��a=�Uz� ��q|��.��%,�ӓ�ٓ���X^@�akh+a���A"�E����D�{�|�_����e�Ud
M�<n�>�2o}�������⊒��ե�����NU`�<���6nuf [�#���L �=��޵XL�?`���{Q�%�/�N��?Wz?&��
��
��R��;=�;uh	0֙�O���1�5��M
6�+�զ�1��	s�r�u��[V�D�9������s�,a`��0v�Y��,�<b�����MDZ
�P��ا"!���t�,��2�k�q�V9,�h���v��!��A��c�a���=���H#�� 2_�*T��6,������E�F�g�u��e��\0�:���/�����	�:3D�
�`!$�o���~�ǜ�m�����s,y!�lޭ��.!o���&�U7���c���,����۷�u�ڿ

A�l���S�v�;�Y���k`+�c�k��,�>Һ��8Mu��?��W�n��ɚ��gc��|�k8X��ͬ?������34��CR0Z�X��̛Bt)���ķ��r�
���FZ 4}�΍`Ƭ2�vpt7mN���ӱJ�e�!�Z�܏Q�L'Oŗ����vb���gC�4:�0����`Hk��|G���1q������x��vL1e�P~�6uao�u[�A[�[T��V��ޅ�����q)�}�.��/�1j3�S4�������U,E�-c�����]�)c�q�&�S$��K'40�P6rN������"��*x���G��ӻ�Q.m2�3�|�1&���9�j�.��'Հ���jƅu7���2j�E��rT��5�|�%\��������u+���%��E5 C�{zs�"l��\�D�-�:e&��d�X6�l�������oSD�c_Ţ�4^x�0�qI�7���t��Ld֠\(P��(��p�'c�G�d?���	%��d�n�@{�B��c�9������w1�lQ7����ss_l��C�X4T�U&M�=xވ�z�a-6܁k��E�W:����\t�~mC�+h����}S��4�5wx(
F[��CYɨ�"tv\�{-���zȳ��Ζpp�֔!.h�(�'����)�=�W:�/���Y���#�e����W-�Ҫo��C��0���.�Bn���'�}+�gF�\T�=$;;��錅���彮+	�W���O%l2m���U]c2�t�R�_��6+�	��P���}v����I���"�[�g��j^�R ��i��qE�LG?�|��m�Cx`(d��Z��=Q wؽ��upNy�􄮶�l��#�D%�YJ�Wt��#��w`��?B�������E�ygD�)0�j1��9Q�2�$n���h�Y-�0�.�� 9"L�ŭ�a��Ԗ���F�:ڐ�[��\X���ɷּζ9���9M�{c���^��ݱj�9��j�D[��E���羭�Ks4�{nwC=u��ms�r��ډqx���t�W7s�i*~���Z����~	#h������6��s1Ϊo_ב���C5ۼeI �<A���~@GyR�f��Ǜ���t�?5�/���ٽx(,�?WW`4t3y*��C�	,�t$C��=
���/Fl��x͚��:��Տ�գv���2��������NS���Y����-��=�ze��	1xG�X5eԶ>���]��(g��m�,�:�_�
���Bctz�w�R�8}<-�	-�3D��rN�H�}�x���p,?B�'���3ų�)�v�S��<v�����13��;���Q�쥮����?v��]��N����V,0�=��d�p�Y$�������D>��
����<��y�^��0�2P���BBv��BJI��T�l��2� C$$4��<����jj-�=���@�9��@��=eEө��leЏ�:���E��>G󨭱�G�5�Y��Fݛ��n��=��G,i����|�-)S	H�7(�j�ɳ�l�n-� e���ʾR/6B�d�(	�-<���;�\fg��c4�$}��a�US�qbg����z�����9͘=�##i�5�5�Y��S=���Y;�^G�ڮp;���Y���)or]s_R��d����s\ T��{P�Nȃ��'�-~b�1�$V"d/�t}��͕ O����إܫ����0{�|u���>��]���|*�hSd�ǻP�Y���n��Zר9N�|i�c�T��9����<�o�E䰃�x���?;V�NNv�����`�%��p,�gְ���)!�#;�5�w*]�v�HA����@������p�IX���'�W^�˻F�Ͳ����1���hv��է����j�dψ������9r�4մ��&��������(����뻳��W��C�Ä 6�_zX�d�0���H��� T��R�[9����o�<�9`�/��]A����Lr�+��coiH�6�,��9���a�b��:"�Mv�	?7|������Z�F�F��R��{�6��yۅ���9r����@�%M��&�d� j�KWZe����j6##�]=j��<31ބ)F����� h�.��$��}'�OÎf�yU�� ����Gߋ���mI���R���r��C�I�)�&Tj��;Ju�X��Q���qG��w{��m\��[����t*�U^m��Gy�v`�w��
\�v�8����֝�!�H��rr�!z���������J��t��GF�q(�G��%b�N��G��$���Ԁ��9X��]��EgJ�!.�U ��Ɂ�c�`�U����ů�ݿn��GSof)/����"#�2~,&�N�o�9�Ca�OH��1��Z����d����	��z�C���(��6i���u�����oSH��,��ҕ0F8	gh���QCGxP�3��4�N��7kO���B��pg��uB|��&��� �/��gi��h���Q����s�[��A�x���FI�Z�ۙ�.�}$��2�vW�h_D����c\�˾�g&)�l�,��;��3H�7��~F���� ��a�g�̿������z��)
s���QƧ`�D��{�f;���ySmS�Pc��&<W�kA�HU�S�ā�KdY���<�d���>�|d���'��4��c���I;ُWX��
��GEee0�V5��u;���j8� ��s)��j!Ʊ��p#�3�eB�r�A]ē7`�'����J�,FB�6����t{���+ ��,,����s�q#�&�v7�W�o�v�Y)ˋ����-)3,*���a#�{o&�6�j������� s
�V!!^�7����Y��T�A
[�HT\|����;�] �ڟ�Y���cc�\ګFcF���e�}��YDSt@ �'W�>e���(ތ���Vf3���ݮ�r�����Yj�:�;�T^^���Y���Y\�:�^�=o.��W51$�]���W��A���������H�����QN��k�#S6C^6z�/�ZZ%�mu��"-Ô<s���C�-�MBv�ϐ5!�+���l��v�,���&W���H0���Z��vƕZ_Ј�w���E
.CK wZJ	ʌ�ڸ\�#��X���Af��Jm��pD�Z�r�R��o�ȥ�R6�m��r��J����Q*R�'�� -����1��Eک��ky�6N�2����b���p+v�F;�\}s�g|������b�(�@��k�M*�)��N��[^tޫ\�wZ�`��c�Q�� ;�.��v�s�O�\�"F��7rP��(�3%����u,�b�訬���<����/H�<��K��R�,��3n%A�>��y�<�N�YI�|d���qF'|П/>�y~�.�h׬|^�-���|�������/YKs,�V|i�+��Og.��թ� #����wJ��)�7��5ߨ�*N�p�q�.ͩ�>>��*��!��xk#�,8cݫK�+$`�����|�mQ	����x�`��e}𛇯�Q���{[���a����]� ;τ�4�e*�2a9�JW�| [	:H/L�MQ�9h'!Gd�\�9ގ�ts����M!��V[�X"�aujy
�OT�X�u�M˽yJ��	��vx�[YP�Hr
є���@i�EWm���ĒG,��%@׺�f����t�$���O������WL ���J;�}V\ �օ`��6�~mm%Dg��v|>ه LXr�a��%�6��Ad�6�?U�y#�,����e��v5����8'��Y"X��$��9��M�V
B���N�M��k���x5��cl'űU�8��Ϗ)F���.�n��'W�e��-r�4�T��z��6���U03]έHTZ	i�x�=�x��N!4�*V�ue�P���~��F6���@^gpҹ�?�^�`�ړMq@T�S��G�T�g(��[�b�N$��8K�2
�����Oݵv~K�?�滖��j����Ѿ,V�WҜ �m#N�k���������F�8i:J3��銩����.���.��R�	�����:�k�1���xm+������&R-F���1�9(5<��������g7.��,�YqW1!��싖{tG1�A�xt�adu;��׈�9?��H�j<�Zq����L'��2^�f`�'.�i������L��(�yA��L���ס�����h��&	�ow�������f�u����q�Um�Rc'(Q/������e����
 �hYh0G�CÁ���m�b��I�bJ�	$��C�3r!�Sv�u���{���T�\x���67��.�E֨]�`h�&8P�U)���}\XS��{v>%5xV}�i��@��	)�Ì�dpP��FJ?�d%
C�s2�� 3�o�I�(��a�L��q�ƣ�?��Fln��["��E�<��Vm6�o��^�'^�9A���������S	�b1��F���ȃ����6�����U.�~\Vv��Q��V�}�k�γ���i���)���6]Y�*��o��� ������{�oe�@{M�쭧��+p�(�	�NO���tZR`x����Ww?��v�r��������o�����R�/:PF�<YX��!�
�$���86��I���g~��q+�k�|͖�)�P�ͼo(�"!d�5(����` �'}�������b=����R�޹o4��	�,�:���`k�u�`�'��c�DXL87%�~W�VG��k����ڱ�[j��-/�B ��X���-�ǻ.����%�A�}@�x�ck4�G�n���H}�.�y�T!+0Y�v[n��7����R�)��,�B��.wi��*v!�0����)F9*�D{Z�6�Z"�q<�V=ݕR���:J�q����<Q�WXa/��/z��PA����M��tjr�k-�+?�HT��&��,m�r��Ȯ
�1?�0R�*lJm�(�Z�恕q�x�.��,���e��[���Hլy4�̢�]�G��V�iAg��vD
�������x�/� �끤��6¾�I�smJ��T�h�<�A絋0��x��GP�Χ�!�P�<�M��G����4�54�+�*�aՐ��`3�Fj����L�ՊG��e�6'�x�lGe�3Oy���\�>%{�r�-]�a��ͬF��JR��ApG�>��Jk�{�����\�LQYR�N?����E�����WV��
}�}��t����L���׃*��C�X���ݓ��c�
��JT{?u;7�F����Fr8�|�Y��³�]�!��yY�jp�� �
BK��i�<./�e���.D��!k,�
����
,���׶��{�g��##:��?�=���OT8z�R>b�}���֕��Dɳ��(�eo��j{�@�"5��-п�	G�K�C�5mw]��!+|�պ'���e]�O�O=�Ly�]��yi+�˃����5�.�-U>6�_]�Rm���=���}n��(��5�B��Г7�ʃ��}E�=��vş:����UU�%���?Dӗs��3���j��?�n(�ԘXC9R��n�)�$�kn3%�?�i���"�l�yp`Bg���,�A�Ĩ�I��n���E�*�����������2w=�����?β� ѥ���^ʒt�)��̀^�N�" m�ٌ��G0��������c%:���)�Hl���|��֟��z��b
a���c��Řq���>��OZ�@^JI��5��>�H ՛M�^j3�e�.�Y�G�>^K$��i�T}�^pEQV�p7�S�o���O�k��Q��Û� ��dP=DK�ZG|��?L�@���~�	�? ���'u�� ��8�ED�~#PF�G6)�R��kƙIڵǀ����`3Y�r�BLP ��d]��������t��Q�mT�a�Z��Z�Rb߈UI���l�����a�Z
���i"0��_R'(�� 
��Ud��G&�~�����8Ͼ��6*�xd�['"�Vvx�? F)*����
����E�t�kJ��ք�5�S�o��oO�y	��H��b�؍�9>|i�S	�l��lD[����Y����I0��?�BEn,L� ��9�Sm�pQ��Y��Ƥ��CHi�	[I-T��/̓�G�i�C���^��l��Anw��|���Pb�E^Qrb	���hB��d,���]�,l��z4�](���2EJb7�Z�`f�0�ڏG�f�*&�jP�؆��N�D`�[���9 }��ͮ<n�y֟�ފtV�3@��Z)o�s_��;;�FBFl�dΔ��?2�)e�i�+�T��G+s�"�yZg�P���lQ�\��*���� @��.�K����6�v98!#�503���xD��oX�3�%�P�`H�;�{n��H��q��);V`W�"��3��T�qkrݒ�8h^���Q~��i;�֢�!fϛ���0�l�'�5��q�6��(�}�ǭ\�&D�q���_:����G�3���Q$O����������r���٩��cw%�VE���T�r%B�����q��x���!O/��g[%��&I(&�8�e"�U>�ǢM/��S�P>"uc7�"�-<��L��>�����1��ë1c�Q�	;�C��/��ф%o�:�h��ZRV���)��۽
�B���A�s�ll�\L6�^����=�ǵp��p�'���-��y0Kߵ%��~s�T����k�4v�m����U�Q+��dx��Yka��_,GP���ѕ��<�؅~7Ԏ}�鬊�q���$�O���!��4V��@p$@f���9�t���$Wenª{��������h��L;�bC�q�l�q�gӿҹ���^ e��8�19]6����Dȃ����S������-�^��B���"�G��@�=pQBks��J�l�	�㲭�zgdtP��)2�-��������:m�}z�]�B�+�����aM�H8�
���<.�T�7F���^nB�]lC,�#�G&��f$gK?���k9:�=��($ۢM��Ã(�?��%��iV�uH��ۧT�IĪ%�- � ��?��~ƛ��5Wx�6�䬂��.���h�3=h���89���Ђ<>�b��z��_o����3��w湁�i�z����,G{2��@�IM�^a��Zg��b��y��O�[��8���A���vf���k��w�'���-Qk�H��Sg��	|��qӜ�������M����fR({�h���	e���_&�\?:��}�)	W��� �e��Ѳ<���]3��@��r�j.��(�d��jÝ������E�Q8��y��x�z�f���7wy����CE���*�v��c�N�P�f����F�<v�o�@߉p=#�\�2���o\͖x��hJW����C��O܀}_E#����x�cZ�o�e}ke1�%�Y��� �w���}@�Qт�т�S�7��qQ|QȽ��:v�2�������С���G����vKN�� H���L�����zCL[��v���H׏&<�0�I�1Et��(b
X�[�ȗ��U6y<[ZW�i�s�@k)��e{�{�ũ�Ty�o�2���O�O���.�k�i!J�R^��ʞy�]�ؙ/�?��[�qv��V�$��e')D��i`�K�c�=-q�J�eT���n��f�Q`�mm��W��C�"?ѕ�նR ���i��j�n&K�.�Jx��$��C2�^����&.�&-F&�K'G�����&1����n�n�:�H��c/�3�An�D�p��G�)�i�I��j��NX�ٲ�I��sLJY�U7�7ErU
+5����R(:Y4L��@�q����ktK�9i�3��yB�s�.���s�uqx�h�(L�!kIp�'�(��sW5`n?~��$Cn���:=D���F$�J�BE_ܘ��&�297��cvݫ�����XÒ?��,d��z#��3{��ږ�� +��G)H�c����[�:����&��g�@�"�$��s�|������7��\ރ�~�9�׋|Ol�A�Q��.�Ťf1�PD5�jP��3�ܟ	�2��;ި6Gd���.�G�{���3S�w�gT�����!')Y�nTm/�C�45L9� 0�}����++NS�W���e�Y����כ<��\{���Ta�Ҥ���Ah �����3J��W�9�g`#��H��W�F&&�D<��t �z1�E����4��#s5��)F������3> �������aw��Yo��8��?�}�~��hK�����"�P��L�<49Kݥ��d�Y�x��l�HD��Y�TbH��B'D(��F��!D/+�>T6�)�vŉ���;��d&Z�K�RdGV�=H)�7���s4*B>�D�}�i��������j9����2o?FIf��&px+Z�Y�Qu��_* ��8��T�U�)�ˮ	$b�/�����x�[�(0KxvC�Ը�K%�3%R����X�5j	��b��Z@қ���%��OdKC*����!,�0���4�Ie	���Tr�̺cDZ�����Iň�4G��#J[v�q �&�:�������3��!�#���N�3�ó�Y&n���N<^���"�f���j�Y.�8�7ӨF'��:��-#QjS'�dm�0Ҟ��L����>�*~����	�'}���-	���k���|y�� ��S�[y�����C�:d���8O�?ܥP�hQ3<�
;��\����G_��S'�^��+Ѥ��py�֬��{[qD�ݱ������r����`_���r��b�c��r�bHYj��,|���G[<OX)��.�n��#9X�����3��B���YvyQ_K�c�Df�B3ĝ���:GOtF���/	�8����*D8dR�;����>U�xa,������(�������P�~R�Ͷ��Z�.�,>�\�n5}���t� ��zG�㟷Ty��;R����.�S�Xz�kU� U�cVS5�V���%e�Չ�.L�N=����}��D;�y��Uu`��"��cP�˔@��|�wǣO+R��LqU�Èf�~`�Uo �3u���z�"Y
�l��]��$���WM����6LL���G���6�ЖBW���dz�gn���4��fQ��fdY�	f���Qިe��o�N��`N�W����j�ꎞѥ��!x>>�Bmg�+g+�1#�B���N�։g������\���X��Q4#O]�d��㺌�~�y�@G_A�
\`A.L=<sӏ��Qz��X��BgE��I)M�Uur�����4 ��2X/�Po��)F�/��h�D�!#��-}������@�e�UY�=�R-�0���[5<A�e_K���?q���:�|�{b��"�k6���B��T�T�-D&���B�E�/��6�����g/=��m��e@]�1�n��Ӽ��+��	�k��H�8ʉ�k�/Сؗ#���ѯزm[r9_�Q��	Af���N7;dI�q��&w����L��^�hH���!�����m�F5���f��k�i��^���1D.\O�r/#����8r}��u	��6T*�f�ױ��.\��0��**@��b�j���]��"P��Xï4�]�沨T���+�Ҟ�P��f��7v0Hs��)o�E&6�p!g]�WD��V6z�]�U�(A׮�5��������V�idRk�ho�ρ�>�>|f�wH��q��z@[6�ӆ�)J�k�����g\-���{
�	���_J٥�S�A�7�x���Ѕ7��'�@Rꇦ��:OWu�Ñ�ے#"uG�2���(/�d�̹T�$iwb�@����|k�'9��,���#����� ���^�s�-��*t�:���ޑ�cSFO�`���p�˼�IH�L��
����Eç)��}k�n�u���;Z�� k5%S�#�QXv���8ݫt��N�NU�P�ų�LЃ��꾁��H�E���lx��Jz�N��o��ؖ���+����}P$�.1C��>�6���ga\�Gt����d[��F��RWuv�;�y�lTK�HW06`5���n���߅뇺��6���A�*#R�ŉ���Z���U�E�C�����N�H�O	()�@�ۛ��̻(��#�	��g�WS�Pȯ�'��u2`jV�=��V#��x��;�yk��;�¾�7A�W�Xa���	��N�m�v�K����z��L��Ͽ���-�Ҝn�`�TKc/���9`�4�i����⹢�93,F^�������A7I�Ew>����^z�=�_R8��-^z%�疉E�U�� �zU�p�<e!�����Bǯ:G�j�z�N
Zw #/�\ofZ�,8�3r��{; ��H��7�����t�q�=?s�O�#h�@(�\��r
�q�t�|>���;c:7]o]?�qA)�5�G�C�ޝ����Θ+CH�.����o�y�r)k�xɥ2X��灤g��.!�j��&�ˀ�>�z�|r�2ͯ �����B�l���ah��Zn�{�1��0�Y;Zr1a#�p�l�߬l���˗);�p����I��a|�������s;��sSc��P�ľS}�[�&�&�LO66葎�7"ho�穡����������>j8E���>�̥�ȿ��FN�Ȉh��`vtp�m�}1},s�>�5%�0���Y�\b��N�z�INu�L�ԋ���)��}k�RzJ{\<��B
����DK;��ѳ����m��������ˣ�5�C ���V����\e�����g\���aMe*��з��ߖ%��J���+��%#��s��}-7����x�.�N��6�7�����ܫة]��Y)�z�����+�����:~�w�Y(x3�y��Q��J{]��q�G��n�#C;^��!%�|�~�w��������i�Ăk��n?�����c�Q��{��?ϻ\DX��q#�Tϼϕ��Q��	ƖER0��A����3w�0]#/����m,�1tjUM��}��"ɴg����1�$a$�RQVf�@��.m�L��a4�'p+�U��w�ċ�2���~�%ڛ��t���O{h[�0!k�%�� ���[�c�6"aa?����'tjUnY�w*8/��e��Y��|���D�aM]�A�nb M�����}���,N��:��1nX�z�j���Л�d ���g��::�K�����錀K�*Ph�7q^F�W��)�?=f�@Q��X��6������E&H��	�,t���zȱ����p�&���Ԛ槿���1ln�tJ���$s��Y��a}�j�]�?��i\�ġ�^�,�4N��`���ï�&��
�w����Q�p����+��G�i:�>e��|3-���	g�3.��I\)!��wûD�b!��ƗV�6���x�h*OHIB��7�#mRƪ�3I����LL��ȬxT�&������i��j�.���N�y��tds�̹�TE^h��01k��6#���:H�^2,�)`�i�u
��4��h
��(��8b)�>�o��曨|XXWPq�^�n*6߀ܷآZ��L���f"زr�"���\�(���S ����Nk:_�U�/F`0z%-�xwW�^��ɣ�*CL�z[G�k'��K�N��>�Z�Y�lo��������̰�񚏺� l��l!��Ŵb���5XUj.��i��5c��v���Jnj9C䊡�LW�TJ���&K^�;�����,��|�r��u��o��7��ڠ 1tn�r�c)?܇7uz�H��e�X�/�h*���\ٶu�x�Q�|�	=�'F�G�4;
���0@��l1��4il	.%˅%E,Lg�r���+B�J�h���)c�^�Do.����949(w�Ea�l�_�)�:q�.���g�^g���u�F��J��.K,c!�[Գu��~\zxE��F��"��=���JL9S���!��%���'�@��6�Y���at�ሑ�/��ˮ���m��(KB�]#�Т�\u+3�F�AScE�'����c������r0���+�IjށRE>��N"�Pά+M˼�eu�|�#��i��1��\�Cʺ��&��X3������R�J�������!�e�`���A/;�6�U�]�Ϧ(��Og�ߦ;�o_�I�K�p��7 7��?T� �,��p�X�jHd	z�g�% {���\����x��1eQ�vTP����~�_�|*��7#�y7��O��}����Nj�喝oi�Q�i�lh
������[��6;k���j�p��ԧ�,�kl�n��<"�_cW%��������~s'~Zύ �v�ϟ��D2U"#�W�wҩ��Ц��+&8�"��b���'[?�M���3��l��F$�߾ �rv��;�u�ډ�I���P/�ˋߊU¸뗞�����}/��~O�NӾ���v�1����G�������� O���Pe�|b1I;�ǿ�1�r��ث1�ي^����6��T/{�*�֞�&�g����5���3���F>W���[3��rCIN��$��� �w�I�@ݘW�פ���d�v1dC��� Ď/���9�J����L�b���ԛ�ta.�@�N�2��y)m;4C+���B��~.E�Q߮371��2)�6�6��%�>��qU�&t}7���t�ַ����"̍�j�e>����A{:qgD1ହbm1?���j�����Otvά�^у�������j�+����j;*����{�@�Y�d�},0Y��7�YE��b��Ũ>�m�j�j�a��u\������s9��ے��Z�ߡ?����ȼ�ׁ����,	=�X��3�l�u���u�e�]C"2�������Ny�O�U��Y��nZn�����G� ~<�Uј��8�$@�]N��g�F�(�^'�n4���O��A �/F�y[C؅�ӈߎ�Ͱ���.�O�-�c}Rx2��ϥ��wG�����-���W�έI���U�f�rZ2�$����(�nwFJ;��7Q��B]i�����o��gWS>5��5[�>|ҀH2ݼ�C�<���߰п���Z�EIb pm>K�;�Ϭ�k5ƽ%,W@H:�<��9ے�StH'E�%<+nE�9��!���k��NM@J�Q��H���K51�C�:��<���%�q�`�V���$�y����=L�Q���\uBa��n��(.�n��]��N7���ʃ����=tBn���,�B�m��R�V�H#���d�f�A�(r��K�Y��	@
X�ݑ~������X��(4�Y{f��H�!��MY�]8!�m�s����(C��8��i� ��8O��
 �Ih@���F��s��Rm��+��1��-XW�Nۨ�
��$5��^k#H�ݫD�,\��)<�A�	��j���Q���eC�v(>�-X�~'��Ě�(��DKb|B�˕��ä�A����
$-�';�yw�Cp�v����5�2tJz��#�:�(t�?�S���{�N�൦��7>1��P�]|�c;P3O�2�	4���*~�|�S�a9�AEy��w%
�b6J)W����qѴ�W�8���+!��y���1����v�� {\�&���b�<Pl1��iWL�2�\���p��m| {��>�P���|�)�>��n4=�(Y�>�z��Z�e����.e6w�&>	��=ܾ��th4ZC���
�u��%�b�k�����kzK�O
�Ѱ��U�z�	+������go�����^bια�D���@�25����ә�=9%�dE@�C�����o+ɠ_"h��UJ���r@��^�9�ڧ��4O�o�j����~�0�˱<�\]�QrD����s���]�I���V�a �?}کd���w����n1��^�C�wA�<�|��(���=�L�����c�ߥe��q���y�F;��e��Uا���s�P���[��%�����J�r8T&�А6t.t��~љ W�����(A=�E~�]-�R3�5,�,���v��#�V#4��R�E�p�	�?�����7�$��Wt��k���I&[U��	��V�J�W�?Vf�����b P�f�J���#ui�%�����Ķ,�	pIF����L;�ll�;�D�G�����՗���YP�cp�zN�~7���?��@ut��Y�������/�WZ�k���)��Rz�Q.�/�gw� i+�^C���J�c��De��B�����9��ac���&�T�d�D���{P�M��vr�>u~x�����YT1�	Q�_5=���e��C��|#��~6p�D8 	�����άru���F�}��f4+���^2e�
2uW�����n��C��m���S�Σ��6�a,_�s�����@U"<g�eG���2�����F`f�����j¥���G���4�	�x���k�~�"r�wa�$i<z�t�L' �%՗�4^�z�MG��5;e���:-�r�r�%V�����o}d��t��2��?)q��m-�pmx�,�D\�M���/#^וD����Ұ�s4��tMy˝|�Ɯ�uK�9�fU{	�&�`��b��O}b4Ȫվƙ�� w6+V��ajY�w�MG��eJ=��]ʫ�O�?�N���ǋ��9��}��Ed ���>��A��3��`F�{ԥ
?�zY|�qM�7����N*�P|�Qc�
�����\gkVg	"D�ԉ�$+�e��Xg�>|��͜�B0�M�D��6/�=G.Ct���.pt@ڞE.�'yd1�A-9O2^�E�SHs h����p�3�_-�����jĘ����;�"����R�����o�NѱgA��޻���q�,U�~H�<kB��3VoUo3����(I�Q1݉��rb�ʠ$yR���z%Y�]�>�)��҄����a���ɨ���w�F�iv3�Œ0j �(��ȼ���q��뿇@y�վ��M_�mw�v�V0B:��� �Y�-H��N��H�"�qawY��7n�t�Y�9<��k=�#�G�����Q]�e0�4נe(x�è�d�BJⰾ��c�JFm1�i/����u���%��.ʥy�r�����L"��IdO�^��k
�{_ݥí
cz)Ԙ��[�??c�g��;#tέtT�T���a#R~�	����3�����#*.��N�
l}���J�ai-CRݟ2]k�f���n_�ZF�(��y����l�`�8�4�[_J��)'g�����a>j[��
�TL&�{�zH+��~]KOG�"�h䛲t��p2Y�S��I����s<�S'};��2�����K�P��,6�#M��8��W�����k
��L��#�y3��'��FX���S��I���S!�A�(~1��nNfi���L��f�O��*�na(p�@��[y��7�[���OZ�{ �Nн���W}�=$�,C���	��I�?C%(����$=ب�6:-�O�G�"T�d(�a��JA>rb����z���Ys	=��'��8��>�[v�݈!}:~�c���a �\{�������ǌ��Ϲ���HS���y��ih��<��.sg8�ny
"��fDGu�}�@ʙ�I���rX��i.ϩ�f%��:�N`�@$�߻�(�����T��&��m�S�J�J�]j��y���Yy-��P ����/҇�z�v-WJ�+kc��gT�'��d!����(g|�Fڅ�Xq�Y庖0��������/g��Ҿ�K�Z����$�A�v�]5?ws�B��cE����͇X��測��=��`�S�s�� Z��{��KN7��?�"�NZ֟2����k:�x:����'�*�+g.%�%�jt����ɪ�����^0y�7�	&r��֞t�/SVɴeL=/[<X�S$̃�>ۙʮ�֒?+�J�/���Z|R�zr�& 	�%�D1�1���(�It��}�܉����%p�KX6>�@oX������G� ܉f�C��m=�m�.�x��o�:�7I�*�����L��40I�5�������NdU��P"�:�@�&�A#�i8�1��Ty�Ex��"r��U�0/�ъ���M�_ub�w��A8�����՟Q��/]�S�WtݪИ��?�z��@�4���r������7,v�&�M��߰>S@|�\s|�t���x:3?}�uOP������e_�q���E��U-'MM`���3���m�j�
��l
�B��p8�������Z��1k&�0�f�0(~,l�^�R�<KW�o%f2DZx/�?X�[B����NZ�	K�x�l4QuA��0CU�L�v� Orb��']ܭ�,t#�J���'��\%�#}�}�5��ɾ�5���w�MF�JBv��O#�4��,Z�_��������� ����	>�<K�A
�L�އ�y��』�6�������Q����z�p�&Ʉ�gb/E�m�_pG��>:��dv"��c��I�G&U1R�*_���f'd%�Z��Q�&��ua��DQT�=��B/̆(�/��>��Um�OL�ְ|;��Ǆ�`a�L2�7ރ���T'�z(���ѱ�*?q�42��FW�*��Y�����&�OY�j�y���S�q�(u�N2���B6Ovr��q����W����
�#�"qGnzH�4p1LQ�=�Z��^)2�5Z1�oa�3_�ՍR!	�~�k�_�!�����;K�&([�I�e(��D�=9kז�����s#�����$�p����v�[&5O� Z�Dwz���aqy�b3��k�uwL®k�=Z��TF�Z��=�O����s�t�"3�|��i'oə��J�'NN��;�Z�we�����Q��΅��[(�l�6�iK�!�c �g��V	-|����7��c�j�~`� ,����TC���'2KR��J'�X�a�۵����/8*�ǚ7r[� <x�Jfl��2r�%�L��<�;�7���
5���,��'u�X>��U��7����;��R"\�³{@]�?!�1�O�Ғ��K~�R���%��)�</v۸(<�\��8��Z�Z��Z������y��&��!^�K�š����N�BK�b�o�����o|��'X��!�L���3�?N��hhZ��ځ��eQ�L�t�_�3�&%���~i�t���>��ܼ�H�Su^�EeB��71�ǥL��̖K��SG�/���{ȾZ23�h����S;��<̝m�&�G[KVI��P��*����y�5!��>���sZyΆQ$=Dݼr�$S�CUdԂ}Z�㳟��r O�v�*Y� =�] �8p�Q����rI��G�ݒKl.�O�~�G����O���@�B��n�`�NG�o E��u<�!3��t|��l�j\��>W�#�%��:6ƶ�1/�d��߰��h�K����5������A�Õ�ش!֖�/tг+R�~DL��z铠�o�NIh�U[�.F�?�ӌD@���p�3�aM��=ֵ���7���08q�)]�W�.��ёs�*ނ���_�	����^��G��C8x���s�԰a�(_��Y��{)��,��T(�d��K���ï�ǿ"qIAbyT���t%UM�/Ng�3�l�^��Y�`���$+�4Fh�:#h�5J�z�`��H��hMUͬ=��_A���Z�{�a�v �A�l)�����	�Š�Xŉ�U�����e,D�<��5��oN���e�XX���k��nX2�i�����hȫ���ܞV�3���!A`�@�z�62��X����%���^��wW(e�-�|9f+=}�HpT�׽kwJT�S��S�c��tOb�E�\"� �m�j��<�@����} VAT�ޛ��dO��w����"�\�ϫ�ةnJe&&�d�)�<=�G��\h*Tŝ�Mz'��_������T��s��S4.�qo	\"T�!(��uBޔ|�E5M�z�� �MM=E�E��+FK������I��Q�;���Mm�h2��v�t���v��?�m��QnkO*�����~���6͹ � �D��1]�Ȗa���<��y� S����r�H`���L��@ ��`�kpL!%��g�:����Js�7Ϗ���I�tG�Ne}!}�x��@OM۞�����}� -b�C��t+�W��2�p��ڥ_%
�Yê*�&�Y:�fn�`h�36�&m��z[����n�k�<c���UE
�h��]v�����y0&{�sA~�z恸3�S���\��I���\J��r��a -�uټ� ;����'#(��^��Ԗb�N3ތH��y�5��8ꙵ�X���%��nz�OZ�3r\H}�M�ak0\Ss�=�1Q/�u:J?H�-VE�� ٽvN:�'0���&\w��p�BCM�?i�� �{��i�C�ZT٧c^������
[�������p���U��J��.�o�4�ϓ��4�%:�0�y�H�O@�z�k+>�e=d#��&�n#� �^�b�������ȿ�d�$���m��u �	�P 00��?Z8 �ނ�'΅���Zd�1��.+�C%����@E��cL�r5!>@�ڑK�	�Q�(,�H�8��I�hZ`��f��(��KLK�`�c$�Q�23c>�!�u�6��"QEAMD�^]���R�EO_�Mĺ�X�A� ��w�̤=�q�c5I��hN����ʥ��W,۪��F'�X^���5�������$:��)�O����=��VT�\���t?�����6�߱X%J���uܛXƗ��,*�7��-b�������*��8sI�T��X=-�@�� �	o`�t^_\���=��$�_8�� ����h���\�L�s�t�l����d/�!��I�
��x��x_3�{���X�b5�6�"7�]��h��b�!��P����%�볌�����.�kec���Oc�Jbz0M�T��!���1j;��#�R큏�,���f� �I�zj}۶Z�� ?5�IJ�H͂/t"�K�� �b(����m�V����I;-{���aq��]�n�&%�_��"�9<!��	��/�������m�������DHct#���r�^/=>�J��oHH�H9~I���2m����U���¢���)}�u�c}}㝄N�[�k���jGSp�h	��0�S�$S��6%R�<�.�8�sEJ/%y�7�~�By��#A�Rd�N��3�Y��iHﰵ�
��W�o�]�9o�/�[^]�h$S[#�/�~�
v�fS�+��s��뮷=��_^�f��CˢE+E�"\��X���&!
�(=W U�z��}�n��AsucS�A ��\�C�N��1���eyK'M_iu�2?�����Ie������ذ�Ō�)��o���jd1��iؕpc0����7�9�jØ9U�@��1{���!z�vB۳�(K�*��	�B6v�uE��.m{�"ܲ��^5����{J͡��W4�J3"�����Ҕ������@\BMz\w�) ԱAC�{̠zc��b.�j<P�ѣ*���I�d>ݳ�r���������
����b]���	�d�NT�M��`B��XH¿��G����iq/�&���g!��Qop��_?�'^Ր�.e�J�8����
������	�C����A��GMhۀ�w�~�4��5�0�]:��;ݾ���m�S��bm2	D��X�wL���r�c����2A��qǧ4�%��T���o�}p[�� 8G�J��{��}�׺���?̚*f{��ui���YYֳ� ��՜h�_@PlA1ԑ/�;,;��D[J��|-@��Sn���JlM�s���iq�=n�G0u�@�O�{�G�	���I�C[7YE�~���{*щ)��L��mv�rc:5%��z�9���v�T�_�I;�yd"Mg�#)Ί�� �2D�U�ղT�����=�&����ₗH�97tt� �(�I(����GE�d�˽F`�xZ;4e���4~�*������F-�jԏkؿ�\ �ʹr��e�X�3�Plb�A,-�Ա�:�w'����ȈY�������k	�x���}A�@o'�.*�����MC�!�R������X����h�ΣT�eF(r�ڄ� h���/����WR��'�jc��caQ���i�L�l�Y8@���u�VV��)J��(���d�����̹&<���TTW��9�a�,���{A�=O��]C�$`b{;���ac����(k��`%�6��'�v�����'z�}*�Ri�հ��"����~)߿�C�.Z�����_h%[aW��q_�H�B�Rb*�5Q�qfL�(u��o6�|I_��9�;Zb"���֘�1b��^C���O���j*���-���S�{���/F�9�<�M�~��g��ޞ?{4��^oS@�}�4dcI7L��5�$�LE���"���f�b؉w;�+|T�T��#��zH�I̕jG_o��t���Bma@�kQ��W�A��IX��0pymN= �u4�ߙ~SW�|�Rܞzٍ�����ErŁ�C��i�ͥ(P2�|�4��@����`�%���j�,g}����{''3�|�W��hO[�����,s���2�m}����5,�,����l}W��9Ro�74ٗ�5�E�d�=��i���޼�c٫0�B�,��E8v�pk�]��ƈKnܟt_!�{_�f�:��|ߪ���
�26A���?�9�#���㘎6�&��y��`�.1����]�!�C�
	{5��¦;=�ɩL������F��R��qYv�82���ix�	�q�Gc��y�`���B.G2ـ8S��X r��_���̆hk� �x�F�u�"�}"�]L����MG*��l'Z1�[�v�vJG�'��C�op�I �/�yPm{x�Fg�{�L���S�<����Y�ɼ������@��[A�B{��:l��6��+�'ZfҤ;����l��m�[�/U#�J~�|X9����Hqp�q�+���u��j���N6����t�_P@;��F�dT�ՃuA�*8��;�	���ULT���q=�2֛��ㆤU$̩PS����$Qr�@��x��!���uv��
��v��w�U�I���(��<>�a$;}�up�z��*Y�-J�����_F���`���]��
<�?���v���&k.�L0c�%��b������^��7��>��3\�����I�� n��1�"3�1:2�����
G�z���1~U1�m&+� �&�!@������N���MƋ��Q���ۧ���7�k��L�#���`�|�&:�rؒZ$g59=��Z2���UL[��pK�c����]���
���A>hz����{�z��33a~ ��ON=��P'�2ɍ>�8g(�dV������Iђ�G ����
x�p6L

��:Ң��MX��	9i�߼*��� Җ���>�v��v��\=�ʓaQ�V��@�ߪ�|7[�ρ��%��Fc#��T�Cv���
l�0UL�ܣ��]������<㲀�F-��$�U�_՚5Sb���Z⌎u�"��e���s�+n�G�1��Tbf'h:ꢮ�Z1�&�? \���P�{0RE]@��G*zۻ3Y�X)��$ 8�!T-C�{�[!lz�}岼����{\��c�������䒿Ku�a�����w#T�G�j�ػ�O�c+��F�B�LܳQ���֗[k�K����p�p��hq���K��7@�N)uyW�v$���vfL=W��������B���/��Q�f�gVut��p�_�1��N�~{`uJ�)U`�j�mY�}W]����P�j��]TB3W��z���}�mig�������M��}]�Q����\����= &�ڕ��
����+/���m%�E5�@I��ք��r��cN��@�!A�u�v�x�c�b$��
j��bq���CG�g���U����甹��T+Y"�$^_|���ԣ��nb�0���D/�ՙB��&yF�4�KJ� Kʞ�����4oW�ۤ o*���z�?��׳��J�����+�h]�u�:A0��g*�]�p,�\�7: ���|����:��4�k~������	��'n�$T�= ����uh��)�P�߸4ت�HX�Ռ�0]�T�F�N�Z���2/	�Kh�h��V��_R�,+�4_؋�6ũy�CL}G�`��4�ˬ���U�m�p���m�F�@�L>��2���U^�>p"�&����vT�LvY�d����f%����d߻ٟ[���!ӂr&M7s��y���+�va�IӒ2��ي)��$����e}#	�O�����"&��uukШV
l�p2��&��f��e�5�\�3L�P`|j�&������
XO����e |�����#.��v0�5�z�A�mj�<�%B�����?r�PC i-�y~3
vY,�<��
�v���6|�r�]g&s,���@[EA�Y!L�tKD����b%��Y:�YXr�QϤ��d0�aa�k������t�V�W�}�*e�y�E�_��]�I�\������3���� 뼊�q��2��4i�o��Y%_��OTܩJ�~X8+YƠ�K�}D�*�Catb��GH�1al����K�M.���U��ȟ�{��-^ˀLme@E�(Gv|�6���*W�՞�׏2�O���/���1�>��9ϲ����WeUsB����v�]�`C�k��'�,�������{u�^ǥ�b:Ԣ��if&c��Eg%���@����
Ъ���9,Nq��W�f-a����a�Z�Uj�K6�rcx騑<#p�q�;��G��g_�緬,�=���y�W	D�Y�nZ�g;Ԯ���!�ʂ.6���ޔ�����R�)l/��&9`����!��XD��ۀ��\�*� u����@Q�L3�aG(f{VĬO�~)�_����y9=5�m�)X{K�1��OK����P�Y3�_o�D%8B��⡟�5|=��!�-��d�_ ��z�_wF�Y�k��Q��2�QB�da[���;����6�S�a����B�Cic�s����YWt�6~��!ħV��Sx�9����������9o2�j��%bH������7�PK�(��8mT���Y1�V���rxZ���|��_��}@쵎
h~�з˞+~�ံw�3��7x��hU�ꖼ̸�d��v��i2ӥ�����=�7�Ӑ?�9p� �)����G��V�a�f�t��٥�H�ǎ��BU��Ֆ��-�B-�}�ú����Q�^�<q}�ۢ0Ʈ2`f�#Gę���?�D-�w���Nl��0Z��;��yz~,��g�i\I�IA{��NU�o���r�D��}��.����'��v8���z
�H��b
�;M����[�U(CzI�Ftt9CM�~9l��s#%�fb�<��aϐ�
��#��s�Cn���ND�@{Z��e���V�0]��O��܊0��!M�(x�U��x�A�,��mU>O�8<y�ˏV p��t���d�kt��;B�SĦ��̨MS�����	E�����A���bD���tĢ����ցE��)w�-����6@��}�����`Ų�^�B��:i �X�](�)�ka��?�2v�ܚJz�����j"�0Zi#���NЉ3��ؠkt�-����|М�*��bI�˂J��7��c	���+�P²z}��N}��l0C�g"/,<�p�k�΋C�@���R�o�)FZZ=����BM��-
:��4�X�5�ߝ�:�!�C΃���֕)à������zz��Зew����L�:l�6�G��a��Ռ'( ��>p�^2ن�[)?JD�	�������6<5]�Š�Bp�? �F�6�����}L�@B���*�(c|ƁM��ϙ���å��K�}��ѵ�~(�;6�8��$�2/�x|h���Zmn�W�����(�;|��Q��B"��a�Q���o�rG95В�O,?vWW@��#]��Ri�]�
��� =("j�~��*�4΍xx��mZ.'y��ܵ!:�����_\P���XF�� ���4��Hຢz�����'�u�9�k�G��F���8�K�Q����|A�U�&|�w����&�V�0���I��^�ER?Z��,�)����B�0�N�
5�V,��-�$�͍�o=���j��OIw��-&��̔dC�W�[B�7�����?џ��O�Nʈ�rZne���\ ���� �S&�!��XP��/]�aM&�ۊ�1�X��o�$�-<_g�?�;�}6���u�9��G�Oat=��D���Ob��?2�	�t��
��6WM8�6�J�J�_{�JeQ���7�Ħ;����JU!˚�mj�WY0�!��\��D�?Ru�9*�8����rÜ��l-�X��uQ��L������r�G��yL~1s։s�"��v'q��' ˩���x����yz�����_6!�����Rj-�̫�?~j��g�~�ڵ����J�Z���y���'�'�T�����BGı�8[�|}�@`>���v}�4��@�W�	EU��ɱ�:�L�ʨ%�Qp���ˆD�*"|73�PVډ�6�O����a9�94��B��L%*����-b���fr�Ϋ%p���4��{ �~�_�#��h(H���Y��?���Ǳµ&���Щ��T>�~��\���#���)�5moߓ�%-O ��T�g��@�LfT�)�PXya����k6���/}���GC������@jS�t0�T���/���b�*�f�\ �w)V�v��+�?R��,Y��'0O��mxBp3��C�\[ae,�
�`�G�s�/>t�EʢR�~
���RO��#�5�LA��Ĕ%-�3
XjP���a#3�	)it��ͷ�$#9XW�ء :����]���/�&2nm��5�H�,=f5�a�
�J&����[�NW��2��C��n��
�~����F�I�֍��bJwA����:������;vy�rUl����s)8�A���]L��$?�7��	3�i��mհt9t�E���Bw�{1Ǟ�`�����N�6!��6gE~?�с�5��<㝛���[�ߖ0��iG�H����~�n�@i�S�ٯ���"s��{���Xdg"ʰˣn�Hѻ1� �gz�l����X㎕���]�g)����=e芘��n�� �D(�S�^���p.����<7h���z�	��غ�"P2��S�o͑@ד�3�	ga��x(׶D�/J�D�a�a|���r7��ѱНb���q揆�N�z��α��42�)� ,'?b�>k�f�a����{��Ј�2zXC༝����	3��"�x�� 8�3J2.Q���*�Y�'�I���>�!��z�-��"�F�E1ʎK��6R���gi怜[֬8�\���:�ruGr���ч�
i�=�rs�j2�.�C"��`	<�Wf!�*�����7��Jq�
����S!ń�.��'��%4�c4��vh䃎*�6F�]�����y�E�H���F�ҿ�e��PXN�g��vWB?�4�`�os$��Z�� �{��zai&M�Z�R�F�jK0��T�TRZ/�tX_�M����N��٦�\a��&(��	�5�c��NCYp��O<�h���$^�Z��ÿY�����C��VʞR�����W��-;pl���[ޤ�T�ҏwց�.���ˁ4.z$���mNrd�D]�T�Ȯ;�#����DkF��b6ަ���J���'����C��p��s��폰e]���5|�sT����j�M�i!��f�T���$cQ��.n�S���#7s�d��Ķ��1���H4���E=���WM8g-f0�#�K�*;������]ޝiW�T�>yGM6��;�(j=\�=�o�JGv�C�_,��� 1�t�q��p.�H��eRD�=�?������"76雥�c,���O��?Cc�CW�>�K���4�"r����v3���f�B�%j@Ǿ8��p��c��͵���kh����A=/�a$���u��/���cO��+�о>���g97w��_�D!!�Fz��ab���<�{p
0��|`:�?�`�L+!C4/ʡ���1�mF@f���?=��ll�f��n�W�#�S2Z�r��?���f��WI�1��B�=��S����G���In�%�%�t�+k�1�}�A��VQZ��+��I�(��������%9��6��}F �%���1y�HT���a�e�9�,�!.-iu��v&�8.s�
G��Q��J�X�w�2�'��}Lu��uε�o����+SU>�Ȋx�~!d8T��G��	�s֤*3˹q˕�04R�9|M�,M^��T*$���:��QUP�x��w���%Ş�A�M�Wd��vA$���.��Rx
���0�TM�VfmX ��<r¹^E��&G�O����Xe(3���8�i6M�s�
�c�0�8�Bg�z&&<�P`f�&�W��f7T�*h.�>]`��9;�1�p`s�k��˥|��+�X����j�5!���;n�HY�Q���ԃ���D�-Q�t��uqDf��N�S9�|Yf��F�٣��N���b뢉t�o��xz��U��j�`�4��S�i���J�$gF��Î/���.EU�~�~�!��N&�!�85̳ٟ&@Wƛ�$��?����u�C\k�)�x%,�2K�@�ԗh�3#=˭�z�����A%y-E�C�����^hZ҇�g�����jL���.�s#$��_�]4�F�8	���7x�9#/�G�ۀ���&���]x���wm� �t`r����(���9�H^��G�?������i"�����_ ��-ժ[T�!�G���rñB�Ħn���z�+E�@��A�,�cx��;Ӓ1�'���i�u�c��O��$�=��h�s��&XD^�[£k�8ddY
�3��4@!�oJ�R�0������L�{L_G<mn)��-71�l��@u���
[�DYyvo�T���W,�Nŀۡ9�9 �g�1� �e��{���:��7�E���~B�������-U?�k�8��s�նO��]x���Dc��r[���J|9�b!��]E?��_���-H�cr���@$���c>��|��M��1�N�Nd��<��!amq��'+�K�T���!�1���d�w�K�;�М��e�0	n]<�KoÛ��)������쬾>�V�.�{8��P��"aЦ��Nw�:���<�sŕ�n�����d��w"�^̕dL�RB��Z|��d�'�x�/��GEG�TTJj�e�����:r���wI�d�-����^.>tƃ��L�X�aDW_3���~�q���e�+�Ơh������}�3y`�E�*?@�Q���)���!$�:4^JuX���Qg�By�*�0���\�����f��"{}��j�j�!�����b<-�P���M|�~<J]�,yx����̅�9xx|���V ��h}��V7����
��^�+����*�9�@:�N�3'�j.�q�:<5*�0�eJ F�^��=��@v�H#w�ù�NlH(��\�����=-����>�@ᵎ���G�n���������E��a��S�_����h(*ۡ�S��N"�=t ��{L���!�j�+`O��1��/��E�_��Ub���B2Q&��e����V#�+[iJۛ�3,�@^��{%W<��9QqH?�8�K��4���r�o��anȤx���
������O/fL����v���s��!���t���j
�Gn�F$��#�%LQ Ǜ"�	���6;���n��ъ����)��\�����( N�̲� ]�;U+dT ��%��'��i6�5��P�N"�Q�|j(�m��ò�<�qnC%�`���lb���_F��R��{Z�W �G�7�2�I�R�|����U�*�_���{rv��8RB��K�VE-����fs�&���Yd^���{���[�oH��;<NY��/|Y5(,&h��=�ȍκ�0T3��(����ԗ\��Rp�S��v�tM���\����tkґ)�EWb�O�K83&9F���A�֚v�,�U�V�4�Ԯ���(�:�P�q6�p�}R���fMMx�;XG�'��I�5�T!u}X��2)�t�f��U&��+��W�HU�%_z����_���9b�,�+��e}���_�hޞ��KG��_��[+V3�Ҿ���������a��6�/
p��&Z��Bv�[�:��Y��c2�Eӝ��:N~K�嘛��?��:�#��G��։�s�����>f��W(�����O�&+��V*���+���i>
��wACIMzdI��.wV=4"�X ��d��Ⱦ�����p� `2�[(Ȏet��>h�d9a�S@��<�E�(��3��oE��8�\(��:�<TIG�km��x�W�����#���=19����2{︤��W7�+Ƿ�]�Ue � ?�؜ݏ��¢ȱX�����D|S)/.|���'���؃�Ƙ��5�/�ǫ��U�:)�"�vP�[oxIp���@,�UX��g�<�-b�uw�����ȶ�Q8�]��`�w)�?����Z��4"��ך�@7���<���� ��Sߌ� ߧa�Qs��s�M+��nU� ��n���]w��=�����{u�0V�A�Å�bP��)�*�O�[p"&#���Q���O��B.��ZC���Y�o�V,I_Z��|dc��݊�F@��L�*8��S�E�s��Ԥ�6�����u��WZ��o;&�
@ú�L�p�dG�t���_Ǣ+�[SƑ�]���o���$V]jяޱ���u!)��|��� �4PD��t�S�-w��(��#TK5�j~>�/���q�A�]�Կ�
��W��A���uPPE�o��;I�A��:���)x�h��&Ѕ-v�VR�*S�g�D�Y*�٫Tn������"Ct�tZW��1�� �G�Ҿ;F����궘D��E!3������0|PA.Kg}��ԙ}VtD����}?������С���i�;v�c�b�i@j&u��Il�o���7x�y��oH�W��4�@�.������7�� � ��� ��#ʀH��5�BN�w�Q����������º��H!ac�skh�3�/���h��)��`ٻ�@Yrl?(q�A��#�����!аa)n쑫���fCˏ�u�Rª�,�*����j�*Fs`�}���8�f�!��/��@bi�9:���F�Vi���+z�VW�Q�����'[F�ā$�sͿMC��T�zE��t��6T8�܌x[�R�b���R�Q^gx�RE�Ԫ��m�[�K���?�� wDɧ�ڶ��?מgX��h��9�{���ň֥k7�������D�.�'�f�3G�ٙ��5��~XϠ<�RT�81��`RF�^�c;���1WWd��F�����WA>�� 6渜;?��P˯A�ԗf)�U�S�ug{fu�)y!���k�����G�]��\E������9���t�=L�^(ق�m=���`�}x��B�u5D�������mµaD>�5��bݘ�W�Q?�bc�@u�%�:�-�gn�ZCLVe9�����A,dU�Ҫ�O�Lu����y1L+�4]I4PגA��2!�׎ǅU�O-;��)X{=p�f�<������y�T.>A���\����e����C��t��5 �h�[��D��y��>� R�N�d�Q~�[�p��:h"���L��4<�5�����!Ϛ+�F��4V�U�R����Y��v5�wd���froks/�q3{��y۲e~\����7;@ʕiC9�NЫ�.�s��a71)n�;��чb֏�>3xr=���|P"5*=�! n,�<am�:�(Ĳ�&[��{/�s�}�G�.�Q&�������&�Ҫ������+Ӳ�x��7���&z��C���@,�	�����Nu\An ��UB�|��y����?�.��U'�m����qa��w�fC�N�>�{�BVƄ_���i?Il �iI-�!�.�Zc�6q���B�c�U57,����ׂ�b7�w�|���7s,�\����FHQ*x�����y��,�<`1��5Ī��a�^�e�_0U��+<@������I�H�Cy��L����YpXQ4X�o��B�ye^+	=���Ī�呐�V(�Ьo�]�� ��E���Uv?�*��_3�X7�ğ~�Z�aN�[��4����X5����0܈'?��+��]��{�m`�@ڛ)�_L�1J5��V�9u`ŖlUt��z'�u[\l��F�g��Q��*p⟃h�|j�z	C1�BHߵ�6O|�5�R��Ni���$؃�S�
�kw	�2q�����f�`�-�+=�KPؕ;�i"LȎW�HS��<�*���׬
$�ɴ>m���*fe���U]Zد���Bν�����V(d���G�H-�����g���4�
b�>�V此�eZ�m��_���*M��g��9]���zZ궋��}EP��C�{97�q���Ӡ�}8��>Æ�a|j�ɽ��';{�a}1��1���:O�)N��|n|mT2L�������z������+#��G�.Ѕ/��q5u�i��p^��A�f�g�K�̡�D��z�Q����H�(2�]�M�;ָj��B�HS:Q�u��aZ��<�]{e��y��A ��`�d\�H�`���(;�;��k�����=�벗��F���Ҿ�WZ�Qq�\��a\�� ��Zg,S�RSu<H���i���T�<D�/�<B��\3@��K������H���/y�ǫ1ˑ�JQM�Τ�N s�T��厭NLóitBk��$�^�em��	��2TH��^�Q��V�Zwg�.�I�Gl�L��o�Ay��#����K ��M�d���ȅk9tؾulv;�]���a�c��zS/�}�ԡK�x7@��r{�e	�Z.8G��N	
�6'��ci��B�SUz�DX���c�&h���~�T��<�C������f.p���+�Ox��*×�% �cyq��6�<�#G�_�3l~`B1��E�cA?RgIYP�Zʈ]}h>W(�b��釔ż��lg�E+��n�e@D�U�֐��ffVb�atֺk�Cf��4qP��)`vyfwH��D��uX��%�0�w��P���\�)�J�w����\�TD��tD��:6cc�.�?�W���,^�X�����=����s3x��*��uM���)���3�t��,hZ0KGnr��߀�4.e���+Mp�?�7�b:�K����̊�r%�)V[Q��'�tz2|r44ؙ�˔ڌ��� �"b�<(���	�S)�*S�9Z��J�2��n�V8�z�hK�j'�I�_�ar�t)����r�Ѯfoc_:�o�����T_��m�'3>Q���L�m��qR��H�͂�E���<��њ��M�|V�X1ݦs���)dTټ[c+���?�,����x2`7�$ �����A��R���Cy�b��Y�T����o�w�6ȸQ��W�_`� \��	��82���,���o���=ud��s�S�"��Q6u����\I�1 �vL������uVs��!#$'�c ����GH���(��ö���Q��#�����)���>�	a��� ���"���I�Fp��e����4cl�(��ǒ��&�0��w<.	���yN��G�ɜ	a�#g^l @xM\Ϻk��P5a���I-�L@�������pu���C������	�r0ّ�j�4W'mK0����1n�0��&ҽd^�I��h�V��3�_��P_�=r�7�G<c��zi[ܯ4�?*���ٗ�REh'n7��I���{���E���ğ���ĩ�_E��1j�9�l��xT�0��I�2c���j�r�e�kA8�dڐ���=�'��ر
��OM��3��^�� ��H"��3�2N*���6�^��-Z*���Q��}���ٌ>�#��;�t�F��X�~,��s�����o����٥C�7���*ieؒF�Ǳ�ę��3�R��4�P�d���q/�g}Qӯ�N�	6��I8
���l�M�}��s��g��X������#����[Ğh�]�c�
L��7U�G[]��5��QY��"��w�\�Q,�P�u�(Ku'&l;�Mє��xO�~����N����E��+`XA&2(�]�Ğ�4�:vl�Q��������u�"�a��z �6?�����a۱���nD�XaI��zn����dś���8t�:va�{��)Ȼ������n��3((��>^��ta�/Լ^F pg��wiT�5r:�^�s�*�Q<{fM�8 ))\-��RS�v�GG�?LJa�RC�M����r�Fp�8`�g.7/�=:S^�?M��CW�Ge���jL��ӊ.�h�7b�R��}A�hg=s�x�n��PS����s�m5�4Y�c�`�/�ս�/�1U��yJDH_xEU��*�G�.��pVq����h�)�5o>��P��E�����1��ujs�M�Ci�E���}`�9���V���q�\t��@J�y>|;��g����,�m�TǷ�g)�@G�Z��]���,���B�������2���m�@Si�j�=M�h`���Ϗx+a�PU,��W2eQPr#5�?��jV�O�<,v�n�i$9��Y��9����$zc��o'7��>�B��\}%���Q��m�w^��?<����S2"��0ye���i�="��%X���B���?�D��ǔۀYm����PN�z���)�L�f΀1(����Ѓ���y�A�����0>��=E���X�-�[���Td�����I����;�[� A�Lq�7���R����G�C�Ϛt]i��M6�AQ'��"�z�����1��1�S�w��}�����6i�pr��݈-�I�4��F�6��0��s�mܡcqu�H,�(8z�K�h<���fTҋf�J �՞!�ǃ
�n��ᢤ
�g�<�K"q���K��6�3H�?��7��Q���W�6f���m1��K;�����I�#��`]VL���4�TV��ۧ_�|��!��Ɗ��(f?s�%':��K���M�C �xT6�������3��2GE/���14hW0�ِ�Ұ/��Ò끟�� �6�hMT��o�(��_^��X�M��>x88�d��}{�"s��ď�c��܈t'N����4��"�Z�E�G�v������"<#��b�5~v����v��H�d��'P�۫Vű�W����,�����Q����f���r��'����vN`�cl#*'�T��yF��&m��7KD�S�}n+0�Xց����>��-J�����C�pc�n�v.w�bX{v*��\�úS��4����r�w}"]޿�L`�BM����5�����a-J�HPv�-H�d�0����$j� ���<���Fӆ�ڲ^E-�;��7�/3Cy�W��.�,�^�A@3CIg1V�9J?X�&0(�1�]\��.mZP�1Ώ)�$}�I���'���9��yd1���.���N^�Aԩ1ط�ߛ?k�.�!����m�N+�E<��j���R���ɨ$Z��y���?�����q�C����n��Is0g��B�ԩ: �G~��D����+���c� �}�I�-�s��?�P��{�0 ���;����Tx�c�^n5���VT��C���dd����*�0�����2ڴs���p��3{)�˦s� ���1���ۀ�oq�	��]7�������-��G<�'�N��S�U�iHE~F9������<+��#�x�ak�ᓓ�I٧��Z~����$��)���g�J>�ގcS3�̰�L���1�Q	Խ����
�����7db�M�ݐ�so/m�u(t�� ��������;a���
W��BhJ��&��}/͠���B�ȉ�u��_���S�h>�����?��
gy��.:|{��yX�ݵ1㘤
����`Fe;���8r� �]��3�M���oe���%�u2YX�C��]�ő�T�K��Ħ�f���TS�H��2���"���|j��'�ߞg$N��y�{5�z�i��-���b�[�# ��m���=J�rp\]>�h��hW��0�nI�|��r���O�H<�9]�O���\�����"�l�)c�����_�H�j}�\h[�}�3����䝬"�,�{���j�!A�����q������3��(_Y��(�g�{l=��|}BrҰ�6\܇͏	U�g9���0��o@�����������Ɣne,fZÚw��}���0���p�����9�j �@e�o���JS)�C+L7�!��w��A�D�t�X�v��Bmr�w齕����=H�y�n|�'p�<:��-� �a��w������GX�m��5�����~����o�F�.�W��E�T]���<x����R=u;*��S�M6'�ߗ�Y5,q��k���;}N���﷾�,�{���?�Қ9l�w��%�}$�?���:�2��P��|Va;\if��ӑ
G%S��G��^�e���<eiS���߫$~oi#�YqC$�6�M�G�`Ұ��ZE�Z�*������������${ ���K(;#V[o���4Rk��l#$`Z�g�#Hk�ƮM �T^Q�"���2�J�EIE�i�l���i���su��~$��	4�*�2�,2$%!)�d#��0)��#&�lT�q�_�ZԐ���^��xQd��ۼ�]sي�����S���b/�b�O��yj��w3��mR�`M��a�w]Z�<��곘�?��S��=�mS�w�a��B\�vŖhZ�kX�P��ƕ7�����Bn���
�եE��~�\e+
V�zX�2��	767������	�2{N	U�@�p��:�g�L�':�a�f�O��11��<~Q��E�����	��M� `纵��-Ag� h�4@Ԅ�^���:H�{�x[�&��а����\�zZ��qx"�Z^Y^P��9�_J%��J5|&��X����P�'X�U.�!��YuUD_��I�lC���<:�� W�6rE!�[;�*D��2�M�{���&5+��9�jJ���#�C��#�����z�o{���w���vm��,�7C�w�Ͻ��0���K_�,m�@4&���'�̂7�p�'A[�������i=*�S�F�"������G�����F��KG#(�s@Z`��6��7�8����Ju��*���[���#Y�k��.V>�+k��)�3��~L��2'd4�6����Ej¨�\�g�>�j���'������2E����Q������J���Mf�ml�Z�a����$A U��.*&�����&[!nbk��d�znp�ZM�/Rŭ�(¡�^������{��@49��9e��:6� ��*�����Pp�{�W��p$"�wG�?Pk�-7Q�P5���2q���匐@J�n��Ң�W�vӱE��-�x�L:��B�x�q��}�)�`,x�����I�Y����p��)٧��`h�����9�Ed�4�{�����-�lh.�o�J] d�r�9T��)G���8��I�I�W�=,�h�ve���6'D��HH3��ֶ͔�� ��a���U�M��+չ�.��_��o�H(�@�ݔ��K+��:d#��y�<�eJ�4���^�/=�܎,q�t�K�e��'4��'`��з	`A�������)�k	�[C�4d��������-e	�E��5�w�'�:R�{��W�������@�+�)�y9u��Ȝ�}�p��- O:m�x�T�qk��%p�
o̴��.K��(��it�x6���hº�Ɣ��'�m�ʹ:�����;?���Wk,���F��3��J��4�E�0���0:H�(�����j��!/��h��<��,p������sb�.s\�t�-���,�/�Zh/��2C)���2��O%
]����������Wj��z5��f�5�|9��z3.�%��\�e]WX0�b^�8�Hi�:F�B͖0î���S�M8�1��蘼��.�m5�&�
��F������$�@�x3��U��e<
��Q�I]��\���I�S����xW��u�f�Skc�0�L0��YO������D������Y7"avz��r����8F�ĝʢg��2�j���^�����I�*���\t!X$��h�d��
K˕�܍`S]����:̰�ތ�7����N$y%��|��5=�Z���|��'���};��sŏ�(�H�7�[`�?��tr"�K2���6�n�Ю�hPL�6W�2ɊS�*� ��&T��<�'.u��:����K��h";ۅ�K������HKݒT�4�r)Hw�ݎݑ��G�$!ht�����cC���!?s+څ������kg3�u����Ec��5���O�i���I���	�=X;Y%��z�O��2H f{u�#�ދ���*c��I�� �+�4��m�z�N/�,Z�S��@/�V�-S.�м*[��c=΁O};6Ca軕E���d
f�zo��Ʀb:���c�%�weȍ�8�B.��R��N����i�.�,��q	���*��d<Gkn�[�����U�)�5YfV�4�:gY�VF
�l'�E.]�=|�Me�9uFcW��W�;Ci坧����>4
�'����
�i�D*Γ$���?�P�N�FɕWr-�������ѧĥ���
G\w����:�m�&iO�l�B���9�jO=D��&H��i<G������̂���Ah�~�UX�:�I�JUr���Qd��sݽ�{�k���1<u8�r�-��XC�^]��:�	A�م\~F��vn�{��� .�����q���ʦ�Q`��z��l���yҷ�I���=Q:~r�_f:�Ӟt}1G ?%�����/5�Ɯ�e�!�h��%�f�ǬM�햑<rO�|�JW>��2G��U~V�V�r�{}{���	�Z D/1�N�*��-v�Z"����Ö&Q�6���������([�d;�W�ysZaT�Gh^W�S�tS>�/#l1D;�v��˞��o�!��^�j�_N�Sb̄X��ʐ]�	ʘ���q����ڥ���w�C#����>�&	�E��˭�g��e�S�tȑ�� ���ד�b��&��Z��)9�Ī�, �0��oՄ����mu*�V�<0_ �X#��F���O��KC��և-aǮ�׼��1�/��v���G<��-��K<�o�35�<�_1ʤܾG�0<�lT�������P_t0���u�D��������B��闵<�Ө#n��4""����B���4*'eO ���b�K!�;��cTW�g~�m�5>C��T���d9��Kٶ��hQ�~+�w���\�d{;���:"}������&�����9߱�Puc����9TRu�Rj�6�t�����j+�E��l��5�h,~w� O����i�,���(���kj*��O�x]����KS�����x��d�xns�B����9�7PHBd��}0��+���*�EfX;@��h`J��E�a��,g�t'�b��:���/�$J�m��X�n6�;��'���~n6*��;Ȓ']�U�-�.=���CB$�Q�f����5�3ρ�e"F�8��-�AزZ�wa+��w3;
}�\0 q�,fW�����1�"r���Ƹ�m�q������S�ɈP��L��׿9��p�!��:�ǓJK4�°�S"�/�9~���bqT��ƍ���MN	މ���$��� O�݅Nжh�d����fb'½h��Pv�!<aT��`oz1���uԪ���AMV�n�[���1<(If�)�;:��R����T��we�Q������t�v'����2�Z��1<�po�N�o��w'hAm��c������L=���j
o��w�F�ڠ�e��Gw�*���\	��6�2��ԃ1�=6~K��$�$�6��n�0i��iA�)���懢�.����/y�5�؄O���"�_l��h���I�M��SG_�kDmˡ:��&��$.���l�D@�"#�����:�)�"��T�6����.�-�a�9� u�L�#͸�/�.6P��~�4����<���-O�5:)*�ݨ���Jc�N+3y�-�ǋ|X!5�7^<#��Z1��{���Ya}w#j����4#AI��$/���h$�\SW��5h�2x�[������)-[��Ph�b��|~�{��.#;u��L�i�ޅ�Ԝm�c[!jehf��+�����\�_�\�O��ż�@i�p��c
^��#g�I�^힂�zP��@�7��?��6��?��*��~%Ϛ��L1\j�4�?�9�]:?ʏא�6���SrWN������S.�>�҃��e�q��a��&�I/Ԇ�e�H��R4�@����aDa��]L��@���͍e�}}w�JH���)J���{櫍*%Ϩ��X5���SI��4/�������}a�����;���A�8�T/������%=Y26����]ݕ�Uu�|�"���B���Sб9ա+6bK/����A����,��=>���
,Ψ~��q�����u���iL��KyJ������_�jN�E_���k����7���زwS�z�KH0\d��#�[#��Mu8¡��y�^�,��X��_��)7��֍Y�8Կ @܆����݃DZ!e}b�>	��MpPH*R�M2�H`/A��J���#+-R{�����G-�.$��_~�oR_�ۤ�{4�	'l��N���Ȯ3}�"��4L�-�����et7}У�t<�/,��!�&R��4����� �����5�vA��=���5d�ґb3G7��#�-�5!.o�E�3&��Lu�KY���u��<��p�< ��@I�7K���0z+�VNT
pxer�
�uP����'��_�<�͈X��H�%ʲb\�bp�f6,͒��,n�w&�q�;�Q�W�L�^ҝ��n��FS#�9�ӿ���L���4������De�����~ڳӈ�,�f����T��ꢄ.�w���2"o��Q����[M�T��z��)��^;��/so��N  ���䓵��.�q�_�B�v�95�������v4�D�m��/��� �6��E���|^HY0�!����Jc�U�&�i
{�I^b��L\��ȹ��/�P�N���O�]��jZ[I�59Р���4C�Sv�5a��0��x�ٯ���U����o�.�T�0Ҥ��~?�����z��^+�]�s�2�,F���;A��%�\~m�L7����H;�Ċ�s�n2G`��!�ي�.�ל�Y��V�%���̴q�F]���І; ��N�[%v��﹣v�O�n�n
��g(
��q;8�v��X+�4)2t�&�J�լ
���P�d��:%��͆��1�JKI�o:cYɪ�I?J����ˏ���ǳ��J�k��~�}���R���K��_��#��]	�*�}��̓n�����P�}��Iy�n�O&�f������c �XAO;�i��J)_��#��6�m�D�*0�E�T��}YV�� ^V�\h��@��_@�'�D0�v:�9��./;��4=E����9�EA��usv�"�A�'��ʪQ�0�'fy�8G�E{[��O${�I��;ꈟ�;a��]Ŝ��ؘ����Q�b���]��q�P
��Qk�R�����hqA��ڷ��~F(P,�����#�`��(@�6��깹�U= #sa�E�,����@�	] {*���:��� ��lH�;o�\ s��]�|�+I��̸�^�2�?�;hs��)�E��b�Ju	a��y�0#&U��*���O��(:jMM"-�UY/H�ܰTp&�9?���㗅�%;�]6��Vz�y�;���c�o������>�Yq���`A߯��nx��ןVX%������2��R�C��,�t�L:�Q��3Shp�&�q�!��^���k�MN�ψ�:�㏗K8��M ����X�tB����������UDS��/����8�>IZ*�A��,�;[�Ӯ�I$8b$x�s���IlEI
t�~���+��\��i�O���15@�n����n�
��&'��Yg��4�kv�;߹E��"{����B�E�
˸��d�ض��f� ĥ�^_z���Y��;�x־xc:��,�ʁ�x)p�S�v��x�u�����ܙ=ENE(t$hY�w����T.�{z�H^��C��{�5��Y��KO�C����Ƽ7��Y,�	Gn��.��V�B�[@��[-���TWST�lM���Si���`�Y���sX�����	���{�8qm1���r��SB��*��7US���	� ���/�	It�A��&�u�)t�Us�{I��!��vMО/I�C��W�Q���:��f����;^7o�s�;�{�4�wf���B�N��.�:tx�!�۸P�O2s��O5�q�X�{u��c7w��ma��KTenZQ}��k����%�7�]P #���:�]��0�F?� ���x�
"����v3mpG��b?��.��x`>������d6��"���P;��/%������E`����+�b�����ų\*b'��<�r�4,+��dKP�(��S��9��#�؁d��j���@�>w����H��p��, ~���{#!��v=:-(yo?�d��x4}﨑!���a��f#t�/	� ;?�$����ߺFj���N;�e�AD�Rs�2�wy&��P��<̜���)�����%r����;�A$"{zA�
�C�9�G5,�A���Ɏ+��w&G�ŷ�� �A3<2s�A:7 ��;������ӥ7�z[(Y7����#�76�r�d�"簓g����nZ�B-r�5��J%�+&�Q���;�#>�]�&�����1�C���B��(�T՝��'�+��e�Ih��
�x�1�mU��ߟ��b��&��T4^�U���VVeY�:x�|4����$ 0%̴	��8�ӝ;�0HbF�\+�'
$��k�4X2�����t�vt\�S��$=��b�J��yU��Z�K�"�^c������\���3<�*y������U�pV��	�2�Г�J����!����_VA�N�<!�AYB���P���d���F[ݫq�wc&s>�`�	o�q}�(gݣˎ�t�i�:���G���1���U�:D:��a)�s�t�띥�Kb�(U4^�
%�w0U��]'���英�W�E�Ls��e��'��S_�՛�\_���K^��n䗹��~��O��&�\n��e�@��\T��׶-� MZ��9�Ι
���gN�ab��T�]e�5��+X\�yS��TnLZrms�Wm)Jr�nu�%�.3������x����'��}"tw1�?[�ج˭�jbB����X3BA��4�R~R�&�Z�w'�Y!%#��8����1d���� �,7����?���h{�� �����ȿ���� 8����'��4Zp��i"�k��١��wN}B������4t3/C	Ձޟ�	�7�x*�����2Z�u�k��m(�*NQr�v��[$`63�?�L/�ʧ�R!*����џ�St�К��t[�cF�u�!Z�>>N���2m��A�������E�����'!r~w�R��u!��/Qw��1�f�v6],����]	�0.��T��B/_���B������+��!5�l~j~�0���D�K����Q2bF��;�rw�풫_|c˟)�u��Z�;�Tj�J;���dd�%�ꪫ�syum>�� �^�GO�<�F7��AZT�ٗ"�����&>�:=*�ƣt�G�S��t�`M�\��tث|3[h(�����,��l7�O�'��2��B�tJu4?B���+�1���%��dVtxQa��ʐ�%� \��%���I���HYha�=��]n���3�Eÿ%�zZX��*�:as�V��FR�A��j��Ebʼ�:�Ǒ(~��6��1���e�	��j��^�T)�aZ0��P'�,b�<.Pݯ1��@a�䍧>?α��k�IP����d%�*��M���<F����P���g}��<�J�[�!��$;!yϙ%3�8�ֿ��a./������M��ԾpT���;x$�8��M�Yj��*��
H*A{r��
	#r��m���Y�����T/�}ڋ��N�9hDu�}�`��~9�I5��;J�UK�@0���ɔ<=U��Wc�Gji\�����Y2
�,����ѯ5t+1��
���;�}^#Y�S�)@���/
����f���8��Xb���pUn1��n��y�91���z=������u�U�#�W�<�
��~��5��i���-3�8��ԙW��]Q	���T��O��
�U
�Z	*�]���7 � ��Yк�FX&ܚ���y05��R���2Ms������!/�D�wY�We��@3�3]��^�<-��e$�v�t+��F�c�q]7�8��	`*(���PLC�����;�i%E�M���d��PR[=�>���P�e�$pP��� pԭw1^�������Iw�}���OQ�K��02��x@�N���� y5V~ե?"T�d
�b�����7��{�vƢO;qWQ2�F[q�ͅ����빏�K��B�k�4�����.03 �S�Te�Ӕ�'�5G�աT���<H׍�����B(\�� �i�����g��{9�$ri�ܖU�:�f�j���@r0[��$l� $�#����*�(� ��L*�H�����jz��D4��.�X�S�l�||Û�����~��	mЉJ-k�͊��q5S�x�d��^�|��N��SB�^��P�X�&kM�$�`<=���P�+�'�����~i��"&S�;�ia>�������R:�� j���bx5kuRl �}.���C4��
����Y��2��������ו��D˯A�*+ݯe�QcDH-��b@�Mhj^��O�./]m6:�n���Fc�P �ӖD��p�(5ER҆�'�as]�:�G2��cW3��O��5�=N���vqRY2-�'b*�������Vp��s�#����B k�z��U�Z�,��=�@�~B0�έG����&2;�{XCM ��~ە�K��ƍ���U��0#In�cթ;,"�jAh�p�1[����^c��m����_}Qr�̤Ƕl���+��VO�|�b��|��vp4��Z��F�z�'L0�P�I�E�K�����vq�r���V�
��_����a�;�w��mpd�,��m�z�JS=�n$�F�],��/V�@CL�v��D|�N ���l�8u�M�y�u�Lyǜ��A���Q��2|��e�����2	�%b���erKb�����>G��O��A)��9��3l�z���)]4�׏[�i~�ߔZ�"��+9F������$އza��/D�s?l;kЎBq�<nb�.|����?��'\��y|��u����OFL��3^���xo���+���j���Cd��Z;{�&���9��Z�~0���s\-�
?��ѡE�m*]	^���d�4:��1??����k���k��%H�Ve��Ya8`�7�O u�i���n�c��.o�GJ�G��fF�࿑�P#��L��9��4��U�9�\ꒃ��R��?:�yˀ��3cu�|m��󶯃a��t�>x拏���Y��Ep3vjX*��<H���pA���+_����>��L�~9��@i����@�:�?��cm?�D;*7���$q4x����`�= �Y4?縎2<��~k[��opM�Rg��x:]��p\�¸�����tt\^J�g2�f$�ʯ_V}#�05;`�~]�H�#���[�#Zt�qUN
 ��^ v�bgLD�&�Ɩ���!�;1>M�/S��*|9T�l�<����H�2R���N�T�;#2�b� �K.o�+__�=n?�������=�T��q���2o��H3^��S ;8�$��uh��H��Z�dv1
��+�+Β:ҁM@�>d��'��ʙkj�B�|�s��('�q8�����;[�A�lѢ�C&c:'[*(��:T���-[t�"�Z��k����$�V�b�5O���	�����oP�:����h�)�#B�V�}a�]a�39�r� �J����LZD�5�6��?�`���N�KK�O?"�Ў��\`S(6�����67�`x~�:��/
	|A4�S�)����|�ƭL�S��1>#�V���5�Xnt>B��~��z��S�bgQ["^�ә�s�����Zޚ^l�Ew|�VV�e��W��)�ڒP�E%wɗ�7���}r��k1C�Q�W��gY��O���P����X��5?��5}���l:#0C\+0,��T����Fn8|ͼ1?ّABg妀[G�]�q:�l�����i�� y`*Q��t�o���U��۷
��Q��җM_(��*��v���=�"ʟφ��pS�v�Q�I�5���	�d����{�G"�,"�c���1��>3^\QJX�:���,�X툯`s�n�
�'Xʸ�;(0��pV1>e��l��@}U:�H�D'22F+�|~p|mU�D��\J,Y\'���A�o*���6��*�g�Oۘ���*�~C��+�?b����C����� �`6��u��J��Y2���@��1��KS#���YX*Aɗ'��Y�9H;��W�d%��d�iE��gj�>��@T[u� �Mj?<���N��!��ڹ�%n�7U����aC��\���_��u��f�q5j���y`��C#ץDHb���Fu�CS�)l�}SӲ+��%�<G�5� �������,��X�&8B<5����>N#�s>X�e���qU*�j���t�~�)��O��n���,r����:�"�ʽ�X���V8l7~����C�J1�1�2��U��\��{�;(��B#�#�Ӱ����, v��M�\2t�u�UriG�����8��in�P���������
����U���]E���D�b�CYX�"�zM��l�];���9>�=��*�,�L9/���O0pս��O��`��[lK.U&�4E�{���y��1��sdrؖz�׹�o����,�o~e�r.�����Q~�ɫ�}�/n���y/����>�H�<B.�W��h��J�P�\mx��ߑ��/��J���F%����� �4��d��f�v|��j=h��E��>�Xz*<��1h6�ל�b���G�)�J={�� m/���'��d��Ҩ�Cj�d:|���ܠ����\��3�����/Y��̪�p��]���ڼd��y�9H��7�Z�(È0t��/���JTFIO��Ԛ�u�	�Ty�x$���0m!J�&�����`�Q�!��e���lr_�����f�f�~ecR�T��l��|��T'��6I������3lP�F�P.��5���q1�a|����~>#�V��ܐ�
�;�k��ŝAm�A�1��4W7�7U��W�hy_ ���wN5ʖ� �E��{k���)��G�G,�æ�d�tdpJ̓�g����;.�e�r���g������9�m�P(vE�k��[�!'���ze���,�tP��|&���k��dod���D�_]'f��~Zt���?%�m���}���4�"UX^��W��P�ꔀ�Y����/�u���S�U,h�1�Z��n���З��Ȉ
�T����Tc�ŖTae^DV �8.4��%��$�a�bD��'�sQ6���m��]�9E�sĵ(�X[2畠�CĦ�U�oM��^�*�Y�7���]^������5$�e����ɋ������PXj���"aۈ��3;���g�����lT�������i5sר%�^�TSϞ�� �[-�������{E�e��Vbo04d-���+:0�"�
�	J�r��c%# �� �W����XMN�;Ҩ�{���,���	=-=�&��6�`��kE�]�z�k0펇((�ԕ�Ӏ�����~����C*@��/�NC��k|d�����Եh�>]"���u�c<c�K� e�`Bי�
�c��B"���W�8��P�n���+| ���Y8I��9rȷ+>mh�[�~+�[��I��K�\^�8*,(�{��_�8	��Oz�$����Pv��<z��Fh*i�/J˪�R���^Ӳ"�/�^gk���z���=��ٽ�C�Eu'�.�����K�_�~>RW���Z�v]�4'~C!�gN��l�x�{��h�E8�AI�1�,%d�솲��MXV:s����P8{=�G#ϥe�^�~4�Pz�MX㙀 ď��5�nZ4�V]��F�:��檑z�4�XW�D).q>GREwN+8��6�_�N���3���Ӓ�&�iI���Xi�q	҇��������\��i���>NB���f8�8�����b�a˔'�7����[7�5���e����`�(Ǉ�{��#�0�ܪcK������I}E ������c�4���kWx�_�Oe��U�K�j�e���a�_���yn�:�C7�Q�0껒��v���8ҩD����Y�zVY�u_�>�@�	�rBBZ���b��,#�4���-�=�n1FB�v?'q��e�5;5>�⢶�c��"����m�s���C����k��1�fռ������+~��V�V�.�R��l�6��~�.�FkV��cnE�ػ�}d+��!�ۻJ���6�'�n���	�١��#��_�O�@�#a��3Gn�Q�Z[H�Q��M2 9�!�]�/rPNvw�pŷ3M6�ਂQ:�"L�`��,Ϧ���s������}����ϯ��*K�o;��OU}P�9|c/�����kr�6��HN��P"������V�'d�XH��2�t��?�`���Ě�P�]	ڷ�^Vv���
Q"��/�So�U��^�-+��1uMeA�n[��c�