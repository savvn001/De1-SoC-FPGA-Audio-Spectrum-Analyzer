��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��YlU8�U-d�y�پ6w�����g�?kB��3�qa�اj����h���g]-N���0�S=T	[{Bp6�H��3?h�%�C��\��������͑>���������Gk�x���0���G�&�L�sv�ﱯ�
M~h�ѥb��L�\	��N��i�壖6�H��H��D�2V7�Xs�� s�U���GC)C$sTS�*D�:�M����D9��O�DT�¬saT
=yA��	uň�FМ����
L{�����3�g%�&l���6R��L5���b�^ֺ8�����VVlޝ'T�mV�Z�?0�Pƀ����K�NrOc���j��4q��F�3�����]���^V��r��3kB&�f�^�n�G���c���h��s�,�J��ԑ��̒mБc�e.�-ʿ��;�*0��ϸ�}*�W� �	u�$�9��9�m΋�3X{��Lƒ� �Aܜ-��ɑ�$��| ��f��g�=ۺ�e6d��'�C^�xq=�j�toRJ�7\�]�Ӯ���Y��;��OX��`+a�#\|�,�Pe�%q��w�ˈE���ϥ�AD��{���\�L�݈>�GteD��1�{�_�ҲL�D_���9���أ1����{��֠�r"n6��m�3��յ�*MiVu����֋ǣ�4E���cr��>�ZD��f�OH�:�8闉�ՏK�8i�z!�Rj�Ղ	�Г��!/�����c�(�CW9r_2[��jCy�dR@�z��+����&+�S7�R��KԬy}�ja�[ҟe��~f�U^JTq�t@A|�܁��	�g-LV��ws9�k��ω+���31��*Z�_᫖��޻�k�ItM���	~���ˬ �|���v�g��4��k	̀v�Qd���Ȼ��+t:�mx���?���`�0���u�ɿ/{�<!Q��я����Ȯ&y��,E� �ˢ���M��R��_�X�ֆ2"��sm�RM���M޼0�/��K�I$��۬B�n)C%�%wF���|}��I/�_P���\ ���{-e1�%{�{45_�b_�΁'sS�9�HG~AJ���]�1'�I(>8sX����?*��� �NO��'˲9r��Ɨ���j�޶Q�'�v��L?�.!��9 �==k��3{ɳ�	!N�>މ{�I��ƻ��!� �Ҽ^���ʴ�UU�Ze�#��N�S�=<f���!R�*u�BȺ�aK5��!H��M����~b��}�D�����[���/᡻i�04�H�Rg���퍐>47&P���wfFBZy!�e��i�eg�&z�?2�泙L�6̵y
�"dB6��Z: ��E�_n�~��P��V���r��Cw�:&Y�]���������Aٌ�A��������Щ�db��8�>U�a�d_x:x�%��B�cN��Јz$<~��bw��qd.eGN�[�N�%Tȇ��S�f���Ӊ�skQ��81�a�ڍ�^�,�uYY���J[��mDvo�v�iu��8�#�������c��O��^��6�D��:	������I�ʄ<����+��I5,ap7E�>z��v�Y8n���@d���,�~�5R_�BK���`{7�S���*�^4�nh�a��w$�0�c�b88��OA{V揣��e݄��Sy���PO������[2[���:�]Ҥ>0d��M_�,*��}}a�vƝ�Dck�% �=(��:䔊�$���Z��q��� ��p7wp�����ٴ�Y":�b�rƥJq��
m���n�א������nV�S�hN��?�A�i��4
y;���b]�uX܍e^�W�wˋ:��[=aֽ��qy����''U������>��Лx,�`�]Uʑ����8/	�	Zs��m�;-�\e�}��4���7qf�`w_6S�u�CO��.	�Y��U-��T��k-�Q�xyp'�vH��E���j�M�g�k@θ9�^{Jb&|�3��Pn�As{U���pXe��b�Ĳ��r2��i�p5���	�w�խO�f*��B�3J"��a��+d�̘|��?��c)э`�tV"�l�g�� �Ҙ�U�u�B� �ӖxG_��O9X'���\��x���FҰ����ɉ8!��|D~�ZK��[Ʃ���[����|��E��H�c)�+��c �XPA k"p]zNܖM���g�.�C��z�*h�i���t��TlB���ͥb�>e�����"�3���Q��
Y>x�Q���@9r�\�q�/�oc�V�oT����V�0� YM��C�;5��@*Y2�bP��.j,x��?�CXr��Y�%�G����{,���0�ۓ�Ɔ$�1���婲�;��2�5��+/bR R%�-W�3����vv��~B�)�rR�M�`YL�81��[-)�zݭW����~�F��4JM�����ȐcBF�/�3��r�m�a]~;$�0E�M�Hy��SZ��
݋а쪘���&l�ބ|�& u�wy��L�R\-�8��c9`��/O�d�m���z	~�iTs���:��p��żZQ��V�%�#.�����'v�-=��?��c��|R�j�Ҿ��2!Z@��[2��l���CM7
�lb��8��b���L[D���(�ډ�z9�+���9����*�]X�;U���g��H|���c�8V���n}�i�i�����>�vuG��:��}ΰy���\Ђ��d%���G��YG�#8�
��c}vk.�q[��:�]���2��*+����?�N��Aa�Zϖ#oE�d�LMZ�z�f��/��{u(܏Wg�R�H�x�����oX@�a��OvW�ɀ�eν,9�g�x�McCB�B8�`��5�hI�B'�zp%Hi'PWb���x��\���(QȖ.Ȫ���L�\�Հ�$��%�[���q�t��}~���g�Z����ㇶl��Mߨ�"�BQ����N�:`�$��
j;��Iu�c����ֿl��Q�d�)z��%��b�,Ӕ��+� ��E^��Yԭ��<U-\;r�v�?Q�ļ��}Zf�>�g�X@�̧tD������OǴ�i�	���rU�yh�KFJP�V�������P@� ƀa��[
���Y��[,u���Ҝ�}�Z`ѥm�"U>&�;.� ��vX1����Ϙf1֮��ң�ѓ�|�ǀr����y�=4�T��E��c	��Y����x����׌ٙ����HtcM�%&�I�-av̝��[�C�b�CM��l|��Z�2�4?���Y���F6�ns�!?�&��Z�k��W��;��,S'�a����&y��K+�{ƌ�+��I�eo^|ѡ���g��k�{f�as�"j�h�%Y?NF���TY�9@q�$�?����C.�gMH� |�-�z4�e��T ��q��E%98vN3dI��%�F��Ǟ��b�nRw��l�<�Q�}tF�X��۞��e�4�p�b������MB
:Y��<!5u	vZ�xB����2��tif��v�W�Ç�XaI��i�I8�R�~���P:���	�x���t�Dn���"Y5��bI�GǙ,`�Z�֍�Ց�Z0e9^x�*�oƉ'�Ԇ��ؖ�c�Fݧ�����F%T�.�	�&��H�$��<�����@�F���Ģ�g���! ����|������.��T4�7%�A�a1	�%+�7�uo�W��t���m�@�I]��!
�{����jM�� i�f�D�F岡Xu�x����0�H�� ���ӧ�i������*��EI^��D�;�"�Jz;N�yr�řĉ{o���������4����"��A����K�.���/0�w$�wYa�qz}Mxfky!�~Oxy�>����.�Uk��-\݉�Ej���{��^�6�M5�K��f~�v{��xmT����:1)9�]N�[��оqzJ�s0#C�ڵ��Z������?�gY 0l~�e6�7�����CbR)��{�Wڨx�z�h�_�Q�è!�W4壌76b ���k���A��,+�~�T��]P��n��qB���A���qtC��uU))rF�-"8�e�Rd�5L�����JT+Q��w��<��_��6(�����\o��Z���|ip1�X}��\D������ ��z�1|)٣���#w�/��1nz5פ)�����t�G���0��/�iM͎��V]�%���<x�-�dL+�]w�G�S�6�晒Y����2f�9�dt�"�̀��[�n��̖+�uM�*@��_�f�q��A��H�� ��j�P�Q}n���)��a�<{:Fb��}��Sh� c��+K�K�#����WJz�R;>���c�V�qKF�������x��1!|)�(w8�0F8�Վ��r��]�����З�u6 �r�e��x[��[���J��j�*����Qm�o��]�:El�ku�0_8?���*rl�󦀺O��X��+�v��K�a��Q�š;�L�.k���8�b�_����X[��q:e2o�fQV�7�o�+�O�ה���Tɺp5��c�,��g|3�xÀn����(�p��X�82ϗ���:۞1R-4���O��!��oъfڌ��V,���Hו�a�d7$<��-V�VTl�N�MK;��y�Z)��������Q�i��u��Ce?ޟJr�ml�YG�ȃ���@k$��y�-ۓ)M����E�H�O���R��$�̾ *v��R������V���`��{~>���]�Ka��=��u���7݊��>�����X�u�U[�b]KS�w��N�Z_YI����)��x��#��[<jɟ0�0>C��@�2�������K=��fKZ������_������'��È��������In�|�������[�y�5�F~[��{a�}M̚md�[8^�ݛq� #.��X�G|fM(=�����q.F܏�^�oo���u�]!���%�lfŮ��o����/i:'I!}E	�u�<<�& ,��L�X��؊-ߊ��/���]�46�h(ʡ�vi'�
7�^U����¬��Im�Q�%���Eq[Ꙃ�#}j����g���GD��HH�~�*�W[��`�$�gdQ�[k>���ً��K�>⦍wF�`��hz�7~�)�R��:/�n�y���7��$��h�������ұ�4�#��'QJQ��v�>r��[[�O��%ZB��h�S)�� 1�𒌵�I�d�e���l+!Q�A�T˨�-��쇨�q@|Sֵl�X���r�I��E�<~oxRR���˜�䲾��
�K�['g�6��ysc�¤Kdz�f9��]M�A�@��*x�m��e�q������K�x�o+s�SZ�����~��4�B4�x6I�MM-�U�}����jen�l�U�P����Eg��� �Xy�誽�ڼk�'T�V>���n�n84/c�f)Y�`%�#0����������aP�e#I���� |���Ǩww������ve��6��_9M����I5���}R�����E،��h��O:6�督7֌�� ��g}�8�xv�<�H0Y�>Z�8/�+g� �m	�Y�}�N�����z�ˋ�?�'spj������,�} k�ҝc3�������QA�:��L(5�.���-�a_��I�����x�)�w��E<ϴU�܂7H�g��Byͣ֬b`b��27�φ�JHӘ^�,���H)g�z@�o��0]��n�N1!8;G,����G��X���m����Ck�e�/��$������\*�b��+4݂�}�?�K�g�\Y)�S<���������wH�	B�S�ʹЙ1�X�8Mq�ox]�f���n]�K|�]�֕�`l�:	"Ot�Pg��wo��[�+�q����׃{\�0�M�}
��M�?���zޥ�]��fC"PC|l�:7�`��d�~��LT����6�byJ�xw�/�P��v�F���~aП4�3��!Hי|!��u�03R�o�;��v��"�?R�&��$̗i&	�RM���uQ�5�|X�5��7b����&0~������� Z.��	��Vh��+a��D�7	ٔC�+���u�R~��fΧ���Y�͂��1x`_?*���Se7��Ϯ]h�S�������h~��K���!�U��<�UN���AuP{����x���Oy)� ��:++�YS_iL�֬y`�|M�2��|�m��x��&8N��x�Я���ɲF�E g�2��G�m`���G!>S�d��}-��f2T�����V��s��n��"��k�>v�� f-���cʊ�!�!�Qg���� �X�w��=R�w�"8��蜮�mw�2�����wK�=eu̋+N�_�8��Q�
�^�2rr��S��G]�Vo����%�D'w�5Ԧ�O*qq�{�Ț�u�"Ls&*ʤ/�3p�%Cyq�S�@��I�˸��tRӝ��c�s�-ܼ�!���up�íZ��Y9�Ix��p���X��(2�8��XA�S� ���bc#�p6�꒴I���P혷n���[ls˿���V*�ѫ���1�w$�
O��6��/؁g�����i��r�b�TΗ�	q��4�1"D��)��B�7o�����v��!ݲ�M����v��&6�2� $c�I�
����@K7u�ز��� ���<�/����?c�EEpC�l�T����1
Һ��^H��MQ2=j�J���yu]����tXd�#������V{�	����;�iI+������$�a�������Mp�V�6��݌�&�I8е�;�:���y*{T����7���`�B�p
ʮ-*���fZw�+�g���3�b�g�zd�����eE�eβ����}�W�˦m�k��J���q��D�M�/�d*��ù$*7V�O�#Gi
�g�<(�V2��V�i�7+y&�t��[��MՃ��;�H�3���X�0)-ʫ��J]{4��/�'s��Y�hKj�f��5���2 �M~�cىr���X�+�h��Bq�/j�1s�`�`��8D�uݡH��ú�i��Z&e��ۦ������*��f��0�"ai>o*��)�(������ePY��l/�4bL#�;F�.s�|s�:�
��O2ëDw��wq�9�����leUg���_/}y(s������m��T{=��X�.���W&���T�m�A�9�5|e��
cJ6o�5]���Y!���
y�p��Qٿyg���PK����;k�b��{������g�]�Q��80_�0nU��T\�0�_ �`���!��Cȇ�<��܅�U��/x���e��f!�&�='����f;��E<C�l`��V����H��0���jowģ'd��]��]�,6M/��"/R�C��D=BW��f�P��wOStN����U����(@#
�����CnH��E��*+8;��Yt��i�V������NA�[��#&����酋!Yo�ŝx��A7\"������b�x��4!�}+=i�1�&��Tc�Q-��������\�J;�Y��]�Ζ��16b@:~���ģar����$�鯖�C��tW�W��?�|�����u�3:�.P�$|�<��Ye�q�8�C/���8�MC=aNc�m�̱a5�����?��)߷W�ߩ<�a�G�M4t��.�"�t���2�ǚwZw�d��)m��`�ZΧ�w��y��$�� �#j��!�!�߃��>�iִ7'�̸��(����'�6m�`�!�6]l?4���3�}-荏�F(���6.%!���^v1�>�I(����5h��6��2�wȃl�Dd'+�mW�Q>����`c��j���؍��ӆ�;c�2��Kk�8Wn��|n)^���܁��i��do�" ����H\�r;���oz��R�@��k[���� 4�ЬԼ�)_I[� �Oԃ37| 	ɏ�v�R�$pyǘڸ�b8s0�޷ʂ�p�����w�J/�<���rh)��FUX�XfJƫ��m�6z�Y�L�����'8���o�$L�"HmӨ*��pO����]۸��o�G��NXؕӬ��ZUG�`<��e��H�u���ۦ[�5�� '��V>!(�ނk�¸�����6�>��~8 �Si�mAs��Xn�}e �q�cfvc��)����n���[Ԭ����������o��H�bר���l]A�����O�n��x�`.���v70�E>��8,�7TuB�l�F(��㉕L��H00Dqr�5G�f8�Brⱳ9�A2x;��lG���
�)� %d���f��Rn�vu�>�0�	]�=�DI��c��@~D�e1�C\�&��n���MC݁:6Zrx��� �{��_��:`�dơy ��>�2��6U��+�vpJUF�b�y���O��V9;�7X�H_����/�����6F6�߼!�j<�E�(|^�����t�%��D�����:�/T���E�g�ǣ|�a*�����w����g��x]�������9Y�����Lڡ}��	w8J
�^�ϒdkR���M^�>޵�}�߂��]K��?E�����^�J�����^=Ԃ�6S$�PL����j�O���}w�`i�ӭ ��;g��K�a�1�ϫ\���'���[S6��.��Q{+a���^��󤓾��!`�p�X���g��z��aфo4�i,�k���A�3X���z���]�0�����G�n�#)��;o����Zl��O�b|��3��g�HQmHpҿ��I���*��/�~J��9C,UP�Z*�,���3��W��ϒɣ�x�k~�#�uǆ�߅�t+�� #��@}�'���z�q/E�N�mb|ݤ	��S�*��N�$(�M����ȡ�fٻ5�r,�+��0*X�i,#ߣ1���J�t�H��9���mƌ;�V��m*��5�g�����-6���c=���o������� e̠̒���A^x�,D�8f��[�|UU����Z�ʩ��N����5�{�D��|���̋��<�0�z=ˑ;ZP��w�8��Ӷ|����.�FȜh�b�͊�����m�]��@�9Q��Ŋ���ۈ*1 ��F����U����t�,5��($���W\��Gw�Z�8Q=%�@�ЊX�4 t���o.z{J͒ӈ�N�s��g��Of����6�B�pG��r�w��R�����2�z�x{n� �-�{b����6�3?%?��ηt\	�y�p�:|�F�C��6�v*dJe8e!�jx.�s���=z��OL�|�B�[��^>��G��u��sm��~v����'���/�M�N��~gS�W�����+����&�����,��,�ޔU���	���� �-(EAѢ�S�0�%y��ĝI�c�#����1׉�����K%Q�<k�Ro������= �c�<�s����h)��V]�?ڋ�57�S��q��X��1Q#G@S؉��o�Ev'<�N�>J���7�Dahf��@ƄkV?��Ym�)�,l��R��9x�q���]/�)+iPzcY�m'�x�O�}�6<*�����j4�<���g�؄!����#ham��#��~f��/�lt���D��ˎ�Ϥ�-�pJ�1����PQ����D�ǩ���J��.�Q��������6�&�.�~]<��e6��Ds/�~!�<y�N�"�[���tY#�Qs��Oሟ�X�5ś�ˎSicr�����ů�Kg?�$��!��i�0���� �N`���_�K�ĚY��s�F���ωR�'\S�2���EC�T���QA�����(r(�c�N������<��j��	�[q{�QLw���}o��T5 c��s߈�rІ"�P�7�ľ����UX�N�B׈u�� �9F�&�@N~��3`�^�ܶ�Px�4r�4������T�P��E;whn^i������f*����)�l۩�3<�	�1�g�On���� ��ʓ,����C�ғp���Jl�T�M�)��
�x��ɴ���D��)��
�������B׌�����DS��V�%�*�/�j�;-{+,�6�F��rsB̧��Jl.�?Ѥ�m+��� I�/03�5�0�<#�P:�m ��L2�Kߔ@6�m0x.�%��S{���d�"駚��@l�O�3��c�ڎKP��M�%��B��UT�u�h �Y}'b>U[��r�: �Ө4�|נU��
�_�� ���X/�"?���"�j�5�8�,�H�n�Y�����?\?I�jJ�
{���0���WH��;��:���;�Ԁ�W��V�猥1�ȟl�8��o�&(�4;��:�������0K���;RY��.�e�CDٴRwe%��}���}8K�E��n��˨�V_����6D���h�����T2�����H�����r���4056�u���RC��#�5,V� M��d��KW0ݦ�!�>���C?�):-71�%1�QdRc9��L�W��xF��~	ƁϦ3�!3�e���^�9������IL��쬧?-5�U�D�V��ؓ���t�aK�\����9���; Q�d#�=1V(��9P�F�פ�葉\H�
m.F�Z�ԍ�Hq�,v9��g`�������8�q������+vN�<�T�B��Od��n��D�����_)-��U���me�^�K
�m|��1m��%��7��5�\=(�(�U�,��K��m1��y2�]m�i{J���?�J�7d���u-�\D=
�r��L�3�u��zͿO�K������(كL����݌��(O��txGs�ݫ��]­D.��։�M{ Y��Z����F������L�㙟`]8�i^;2���Q�'��G&V�����1�K|}�.��LvA��}Fx��hצ��m�U��!gy�1�u82l���^�o L�t����G������^L4消��	����y��}F�\�:���:#+Gey��{`Y���g�96�4���?Қ�������-t`o,S���b���wy;(u��+��|3H����`�v�h<fb��d6E�!oQ5��z������Ϻ��}@�iۮ�)�@m����=�
I��?��n���S�D�nx��)�R���?���d�ͼ���"txM#J��O_d#�\Wƃ�#
�iq�\
'�!�Q5y� �E�+y�=��f8�a�Ѱ#�Nc��Dq޾�����0?/:�&�y_�n�΍���x��F/@�̉��R��sg�u�����Jj؄�q�jŌ�#1l{�	W6�WA
�<�%[��l���Nt���*t��?��x��Oe��d��[��o(R�ep Q�U-x�m/%�z�=��߇��bn:�|'w������(��u�ZK��1V��ڈ<�<� P�t|V��X]
�k,�X��l���ߕ��q���lWȇ��U`����y����&�:�'Nâym��p�]U����bA�t��9:獌6���6���K�N��D�f�{���s<����5K����g�%  v��/|		�<�\�t�fc�2n(mh��bz�G��`7U�xѱ(hW��
 ���[%���lˬ�bۮuرWߍ�!����E�?��#�HwWa��~�i-�B���c�-�γ�4���*�n�ڥ���x�b�׻� kh�C���{&3�?o�-��s�j�^��O�x1!�I�BŔ��t'fV��*q���]`w�힇�6���6K�&:���b�'��9W����[*(��lt���`�.M���G��J�q o���h5�}x�@���󤏅�:��"ى��m8J#G������wA�m֥'l�������� �yEAx0;�Y� �j8�`�SˠӔ�FT���e6�a�Ք?E���y(y��PA��h�]\��r-���ؿ�����3f�a���q�:��-��|'2�k>�w�pC�p�,F��/�M����xP_���hI��@�tL2�z>�~Y��-�Ke�7�����B�?��Y���.�ɱ�x:��V���di���O[���������Sm��ν�o�x[��en���\eH�ᛢc8��§��n/*+#��zE�B�^>�I�)7��m��C� �8ߴ%���0��%}���jKY��5�W��[:�����t����z��B��Y%z�l��Bf1�5�ڝ����h���p�����EEt�8"��H��:Y�e�%�]����= ~��eʅ���/AC(<�i���*�mh����!�[��Ӯ���g�W�#�am�$��������q�m�vI�NW �UN�j;&�n4���={��L?�a�f`c⠓z�S���O�"	���O�����O>�n^H�"�o�y�G!���Ibi��}:�y5���r�����')��6�iۖ�7o�a�U�)�������`SYN��Q���$��Q���"�(�bE`.Y3R�c��i80��Γj�X jr�a��=�؂rоu�9��	w��N�YU�)��xӅdf�Ў����\��W"��=}q������u�o��(Z��F~�]S����0}��kV���)  s�im�I��,�����V+�������xd�zag�V��k�c��6"!u�urҏ�e���H�&'�#{{�mo�����c|���^dĐ�A�Ao��~��d�i'g]�[�X�.Q@��W�Q2B�!�K!F>�8���r�>��7��*�}c.`�|��dlb;j��2�._5]1��:��~9�u�Uf�Px�h�%��S��d��rH��Ycմs�f6$�pǏ�c��K�tQ�ܱw�EX=C���s 2%��Pc[��G�*�o{<�����*^�v�T���{�bF�D<��T���k88��s�~s��p�Y^
A�u�l�N��i�о�Z�4E(�7��!����.9����E=4�������F�T����I�3��NH�K��!��ӈ��8�hbo6/�����i�"�>������љSl�qx����	�ZE��NgA.Z��&k��]�u���(I�{�r����F���6;�'��Bs�E<�o�78��.%Ո�\A���)Rk�\��Jŉ��"2��Qv�t�Ԥ�A�Q����>@ȝ���ͦ
N.z۠'��ݹ��r- �Zo�}�����I�V9R��+L�O��6��nZ5�lɸ:�<��?�K��<�o�A虞�$�J�9 ���E$�؝��l��m�5�-�1� �	�����	�B�M�/���Uc�K����>�w��0�r@�x���^^%���lRٌ�C����gR���'��ܙ��iv~SzѪ��e�u(��'�XCͱ�ʰ��b��ע��2�����,ʀ8��.D��}���(X��> ��&\��0�i�c)�0U�*!/�}j�J�GS�L;�ށ3BG�t0#�ެ�R ���L�`����z^'ZKC2!�U�q�M�c���e�ը��C�#I���01�z�����(�d��O9�yZr]�� ��4���o�ux�T�w�����X�_\�7K2���xC0czŮBv�5~B7��b,.6�c�SΒ����&�0���-�f�n��WL�ՕI�8w'��Tp�E�w���ʥSm?C��J���_4�L��)������H/�s
�0�)��d�q_�{�F\�����wyJ���Ќ.0B�.����h�ǯ N�,���"���4��	��Q���F�����e�V�`Q�ք���{X�%���Z�{̬��+��a�'9�x^���z��B����(F���tR+�����_�CS+J��d.��Ss�۽u����"+�|�k��,&�Q��@�ĺ��t��H�H̘�6��3p)�E4[Y��m��}��o����R�n�Y�����.G�c� 8�Y��ψxB�"�FUO��J��s99�����2�32i]w��ߠ����[��cL��!�u&FJ"������|O��V�yw�|7�k��̮N�݇��NC� @ҥv����G���ҝ��=M���HHX���)M�"�T�ō��-Ќa�{8��P}%y��X���9�@_��wY�E�9��Z�.⡍��3K5QAD�Q�%����r�?�Zp����hvޢ�2��%�J�ˈ��l2;���(́h�Τm�zmOP�9�,��yEaD4		ߍ��!U�W�׷��xU�>��..#(��궾�xw~)M\��va{�T�E~Dm� S��W�� ns�^�O���|c���Yٰ^�@���A����\�⺽�\���ʧ`"�'��ٸ�M:�-�8[���UJ�]��铈�کTp�M� lS8*@�t|Gy�G��%ԊBg-�(�����r�U�L��
����+�-ɳ7E�~�O4����� (�v���;#�4��X�G�Oe*��	�k��W���m'0��'c�Qr��*�	��iĪ��_16#�zSrq�3-$P��$>q�'t�R/�V��;y�����A�P�_�Q\.���m:�d��X%�z�iV�!��J�v ���U��-P�";+�Ĕ�o�2E�J�4���oޥa��aI3���p�;Ӂ	ҫUW`�[��u+�.A�+C��"&�nr���%r�qѵ����� �?rZ����1x!&��,��O%���q�qJk`
����&�	�{:cv�J���ѣ~���ueÀ��)1���k�n���501��8D�L)��h ��՗�=�SN�><�̀a�H�졹44�5�Jv[�a�Z��,����8a ��q�ZM{7U��1�ꕱ}�o#]m!��TiT).��-���h�R�����s�\��)��R{)`��S�]r��ı5�iso@,}ўQ��@�������&?�Kol�v��3�h*�E�͛�� RP�us�5��=a�ےk�<
X���E��r������J��h��ާ����э��2�G�TEެ������]������pY�L����c93��R�M}Vn�����[͕��X�ʲj�e�:_*��+V\��ڧՅ~�'I�R�3�Te_�n��.���AÇ������VZ�G��n*]�%��vxf[��&�*��g��a̹���;�}BUM��Lz���%D�)�h�x`g0�P��K:�u��Z�~����:��Kv�G4����"C[�7�)�� ��g{��`tI���KD#�����Uϊ��*��fR2��s��Yd���}��KT�5��1\e@�.:t���]�X�PG��\B�N�<�����Pq�Z���s�J[1IĸZ5 0��ѧ���[��X�e�� C&z%ZR��XE����� ��!pe���z&��
�a��{9>��^O(���Y���@@��w��߱�+�ם���Gfoc̊�<���w���+UNB����g)r��m!#���ӂL�,��/�߷f�ћأ�"f��=v��3�n�U*GV��]�F�L�=��O$r4%W:�+-��fO�ޗ^��C��Kԩ�ɖp<�=#U��ɨŮ��z��%���i�o�u��~;��uA���i���N���
6o�B��;�A=7��E�vs��|@�պ�;=?h=�qYSY�*��Ǆ��뇐��⤖;�����an`�TL�Q����uo�M����A��)iˢ�9��>��/�S]{�/x��[-�T����γ�p4��T�3�T�j��>5NyI1P�8n��%X�.l��3��������³lZd��+2�}Ɏ�)�*Y2�������}Y��9�R~W��c���]p�e��h�$Gڑ��Z�ӏ��Z�P�Uon#>i%O��N&���Xw�~o_�m��z�29��"f�n�3Z�2H��}$����Y���%!Ĳ����y=�J�{�hw��z����ᯥ������)����%����5���KPoff�P#[5����� �&<�sIp0�� �u�(��
��n&yC�F|�Ds��UFP͇�\��b��cXԘzea��PF��nqvך�wuҔ�Y�Y�OC�X��AN�/�n(�r�~ ��+wC\I�3�Pnܔ{��v,����)����z����A��yeC�h�婾דAf��07�>SҘ���O�8/�6�
���4�w��΁>F�����<Q���oĻF2$-T��^j��S2�$�0ed��a쁛I�ۘ�?�t7Ȏ]3�����[�v@�$�풞��Z��X<�=�τ�SC�Q��.W}gC�R�ԛ��݂}��k�hkciX���v������ ��Z�2���ƈVqص9��;`��>u.���I1hgq2��9�a���)�w�)͹{d8x��UP ��H��a/x��ܽCN@��pЙ61�=�er�e���GL�,Z��}���A8���1E�1�\��1�2�*3��� /׋Ԋ3l�9	T=.	{�]S �d��+�8M�X
:�%��q�8N�q����� 5=�فB�g���.��|�Wt�5[�z~
�Ș�@���S�R|b[�����,�Z������cε�G�� ��̲H�|a�U�vj)���H��̀f��Eܙ�BZ�{hk��ކ����Y�w����D�7�+�;Xx��Jo-���mi��hM�b�>�g��\�`/�
���N��#��G�R�b2y�I;���B�����cp�䖬��Q��¦��#y&��r0]�vb�S��AL�Z׋�H���������#�M��P�V����y�\��*E��e	(8�ϵ����G��� ��&�f�YPן�N�Ϣ��!3�����Τˆ�-�WC4��Ǩ��2�6�����NS��W��3FxN�r���Y�ݜ��3Fsӟ��,�{%c|^=B��Hp�>��r��a8r����$ӏ��S�*��jqV���ln�mOz���E�5�	�"���c~��B�(��]?�{^8سs�Rn�#�>�$i�00 ��5�����>6ږ���S���-��;�/\���vev`��q�>|�8<���#�b	a&�0q�M�w ��H��Sc�<�o��9��^��ͪa���yE�-v�K���lI�5��Jջ���b/E�3�Q���c�:�1E�a~�3,�YPc���`����lƊo�{07r�ej�#(/�̷�.�.�IZ`��,�8G�h	��w�^��{�5�	�����~��%�V��\!V`%��&.5��<m���5|�i��0|�:��XR��1���mə�I'�����t;{F��]�hw��n�w�#>��a��Ȭ��ß�4����TU�lI����D��}�> �>:�Bo�*�cq������a��Ih0ȫ��Jb�'�Lz�n�ߎ�_d��#�l��^vwqPPG���E:��t���zهz��;W�pR4yG��I��0�q�L؊�& 5q�s�EͪY�dk���]-P�=sH��(�AQIɡK���Wɳ�=p4����?K�	~�4�l��b�t������:A�yw1,��ŒMߖ޲�=ݖ����7_�#v��]ٍ6_�������$�yCǌ�,(�H Wg��z�,D�&�֍K>~;�
���ϧ�ds
�|�O���6KnIts��Ɏ{^��7Y����9b3������$Q�v�\?W��Z�T��%���|96s7!'�^�����%�b��[�ceu��8���1� f
�H�X��]7J՛Y�P�6E���u��9s��W���`R9,�KB�W��q�Iq�G��rq�	�.�eZ�X+&[�����4��~�Ԙy�;���䕻�99Z�]V�8H �7�����2t��H]����2����?���q�R.��+�
b��Ko�ʕ$����9�T�)�_	�i�j4!�?��c�������� 7�	�V��-����,g1�i�g!9�e� �0���d�
�@B��o�N��4/k(�,ԭI�q�^0\�:f��"�f��b�ʀs�ײ$��T&N�Z5��u4���s���U��*���F-�9�ö�c]\��?�j�����=�U]���6���60��Ј/��n�����,�[#�9��fZ����-���r �J�9*�i"�S�>w������Ӎ7àʋ�ě�B7����<��DVk(t_qI:�a�������d dD��W�ҟ�i���KLPR�gw���(�
�o�o�k�#�\��*p{6�y����=����H@<9.O��T���=��q����-0M�F`mPڗ���YR%c.C����0�Ab��C66�`��[v�3�X�]�7N�a�������h�0�i�d������vs��%0 fM��cF*�j��PMlE� ��
�#Q���2?X�� =�T�(��؇.e��uۦ���v�E����J6�|#8��_��G!��ỿ�m���*�����%�%:�q�����[N�I�5�3���5����Tu\��Uߞ�k�J}�0�g�w��o� ���?�m��F8�ڶ��O�f���M;Z��x�O�#C��G�L��R�^��>�U��)��G�_���c�CP�a�������_�P��:#���w�Ĭ��f����ݰ6c��s�D��q|���g�bP��u���x��@I���q0j���z*(3}���Od�����y��ܞZ4��;i�
��/�;������2���iW��5���� Rohe^g�Ar���.2���O�z���Kr�X���~p�&Z�� ;�=h,��fl�"Y�����I�����ܮ*�i]�B��g��uD,�	���B�>Q��?�G�_90�_�(�6��I�0������ڲ!2�}��.ʤɠR�R�=@G�{b:���Ծ ��K�n���Z�&�L���	���TB���ʤ�\����j(�u�c� 5�?j��-���Ѹcce���*�%�ϋD$��8�$�����-���O��m���t�
K����짘��|�x]���G��q�U�vS�7�~M�0�^�HJ ��a�����+yv����q��֜��G�PҺ�J��`H`�q��{B��� ϶!9��c'��c��6�����?�a��^y��ޠK����dNQ���oyZk��_;_�I>� ӕe���z���[4й7��x�)�ke�����kUO����s4�Oa�M��i:adb�����eg[��|)�zV�$I���x�.fx���+嘥���vD�F9�3H�������ۚ�����?Z	%�
�]P2;���A�RF��D�]}U+�H+�z��g�i�4�H�Y��'UyD�������?�n���ː�;��:$#�:�asO<�b��l`c�_�8m[�o���l�1�7��C{ٴ�Ȭ�{Vz4�ŴKESP|�t�v}_������s0��� N����~����3q%ys��N�����T3�#����M��(�N�V�*`��&f�X������Ǻ���w\��Z`o�-dOB~�]'yBΪ�f
ĥ�[�������
�d�|~5�����}���D�1JՇ����u5}V�~R3�6�¿����p�/w&mQ�ͬ(k�]fg�v"Z �`���
��N������n�M��*���ڢ�>�?N����]x�K=�R��Ne�,�E�Β~_��:���R��ڕ�s���4�5�P�$/̩ZC[̊�^��RRI�li�W��&O���px��jS.��=/�)���/�	
 �ܝ�l���
����B��8�Ab����H���oO�6�vx��e��Wթ=O���e��ܱ�j�ɲ�~WRȵpqӭ�U�W�T���h��%o���p빧K~�t�RO��l����;]�M^��D�{"�$#�ӏ~|�C5����r��;dKZ�^�-c�1����8nSg�>�BN�V�~/���ƌ���5q�;+�/89� ��߿;��U	a\,�������<��T��^s��c�
L�u�B���256�'��G����?Q-���b�����3���%C��V@���,���3��&j:�>ܬ�f	$�5�m�U�o`�kWݎ9��_Watn������h���90q��>��U@T��0�I6A�7_\Ս����+C��3I��C�8+(��!�����P� ��(l�|�{�1����&}�:>
�9>��>˶�zߔ�P���{`v�#��阙��T��}f�Y�����v�[�{��hI{ _q��0��ǣ��3��Oy6��txl��Oќ����y�_���Y�#\&Mb1�2T;�J��A��MyГf�>g�HpN�{��dHK���6�u�U�ݦ߽�S�G8�`���E�1/�����+��Uo{αj=��#ViBJ64U���&��n���5�	�>��DQ�I�*TCt���_�_hA�V�%�G�H�.�3��q+�I�H�Sr��A�^Ȯ��V��,JTW�jz ��-d�>>I{̝J����CrI���mjڬ�@!��C)����0A��Dہ�L;��3F��n��ZWP��>JI�p��[�����V�f�6>�q��H�P�_�9�W����z	��,��H��ݒ�����2X
Y1���um��|!�sEM�4��"���)�a�	�Sp5����l���Fjӫ�Oj9n���0�B������B�DR��i�l�i������Q�%�����AF���1��z2�fg� ��^E_���Ȋ�!���\}�ɸ� U$�+��jb��%}��,p�6�W^����nc���X:a`��g艾,�TU|0��sdu����%�?OF�3UK�p�@�qP�۩h�V^�[�G��[�,ˇk�͇���CX`>��%�FnQUQ��h�&7�o�>te�y�7e-I>���X�-��M�0��͂c�^��0�E:�?�C���N��)d�3��u�Bx���	.Y*�de��SZ	ZԴ�$iھ;sAH���(hʫ�	���7���| ��`��v�ކ��2R�9��^�^�����ƺ�8x.`�Z���9���\=��c(4�X���驎E��6�,b���l�K��1�-�V^�l��2���ۀ����/���3v�������yTn�V���3��/Ab ���U�`��?�)벣��Ȋ�Y�-��;̡#> @G�coz�� ��h�<Z�5"8�����-���C���S>]�uH?/^١OuQF�	&��#��G)'f���X@c��Ա��py[[�Tj�0r1�ͣH�Ӂ]dا���e�K����i��,AT�*�2�ǝ�MI�g�w_��Ir��aRqsAd�S릱Hȝ���f��x�#/U8u����K�jw�υ/�'ۘ�@��D�r�֕��W<�������!;� �k�D���Og���uˬ��Z��릱�P��E�
F
��:����]R�����,�B�%"B(�k �ƨ�0�+����W��,�.��G���5�A;R���*�Ca��x` �������ʏ	FH�>F��3��Bg����S4˩�8,�(�07�77�_��V��74
�=����R��+��L��Ul�]�q��C0�	,���!�_h���ơ�O��˴q�p���F��Z���+�~�I{�K9�3�X���R�$�'uPp�{��^�p�&��]�!M!b�4��ȲF���K��Y	o@�6%�qA�n%x�o��'���K�jW	�7���w�� d�/�.V1c�r�J��c
�R����:��7��ۈQ��ޠ�/��b�b~`t�+�ַ����L�Ka����W�E7ui)�*�RabXCe.�����O#��6�p��G{H�]]:]�������'`w��K-"!���Vk�9���S.=�s��~�,��Jv����_��y�~՞ �/A�1�(��9dfT��Z��[R�ܤ�`l^Th5=�=\"��d�!L����u��^�����,�@,�m��V,'q���qD]��5
#Yį��G��ʨ��:��bÉI��󑆮ºU�}.��9[��`���:��A�Mf�hQ����܃�==�4?�<�L�Bڲ��٠���pj�!bƍ�m.�$87^K/)4�=�R��u���y���<1S�ʼQ�V�������Q�M�"8$�V8"�'`�I�%X�ٳK��Y�%��_C�|�wX��r�ҥ��[�K���=S�%6@�~zq�m  ��}��F�
i��M��ժe,�)F�$�!����^��Q�|��).*#���*D�;�۵�MWn.��̎��>�sڙ��>�us029ă�b���c��_ς	o�-^�ȵթv	cW�f�+��>t�X]���|�[l2��C�x ϯ�e~-ÒuRP���N��-6;�h����I����r�|��>Qߏ~�{����C��3[�-id;�0ݺ�={��#�
g��Z,�Ǯ���'/=}��%���IG������vz�/�>���|�*<%��3
�*�L�6�;��_�鞰��#>e�bv�/�Ty���>����J��#<�A�D��+ꋩC�Ģ�^��u5��t2F�aA�['��'��-�"��v�q�k�Im�/�S�a��Fe��JF]6dn���o�=2~-��� U���s�L��asX��+͚�2mw�/�>��W�e<7��sA�H] ��[euB#^w��� ��2C:��B��I+��d�Ӏ��N��r|F�S\��p��D7�+���z�m2)[<b)��`~�l��_����۝~WKK/
��A������d�`��t����ٙ��Ied����+���aǤ�V�k^�:�(�f@:��Tm��d��Nw�1�>�����X���ol���Q�a�ې�F��O�$NЭ�AZ%j����|����t萖A�GY��4���t{����� ��h��%6������
�����"�Se_�)�����l��<'	]}���s���ߎ�B�V�^�ex��ΨS9�^F���{�mЦ1 �<Xb�zNq�x�E��d�S�������W�ÑC��lzߧ�-�րA�)B�H��);���U�=İ2��^.��t��&��5����I0.-O꼵1�%�������k!NyW'm�,��Q��������{Im]%��x\M=��oL��HM���oV7�m��������q��Kl��z���yuH�|ֵ��������G���N���w>�Ÿ�̅�as�����s�T�!����W�t�K�*y<vUS뼕��7Һ����`D/��g3@gC�l��S�t�2�YMr�	��ɉ
�HsDL�b�GY b�S�ͷ��(���i�V�c���l\n���7�M;�Ù�����+�2���
@����ޢ��#wfߴQ��U�D�dD��T�)
�6&*gp�~��dI�������m���̒h�4��$4�<�7�-x�`I��AHVG0: �,�S��d�I#S�������վ��R���3��\� �I��$_��w�8���?�$�g�;5R���K0��r���ܛD�)�)�zk�OCn���:�������X�w)�y��rʆ_RI��a��R	��_�u��F�JLt��_`�pH(ֵ+�	�.A�E�Ŷ�1{���[�`� �:Svk��a�R�p��i*yr�$��E�% Ɍ� ��O�HJ���K'�D(���1zuD.�����~���	� �r��u�`"@��f}<P�7V���h%5��]X �(��I��M�L�l��_��hZk;w�TP��|Vb�l�I�,R*����q��~��v��<�)�z�_c�m��ek�o�-���8�3�`=��=Ѕz}5ŶI�D��{����V���~�*_�=���Z1$�-0'9{�BŬ�@U�,��.nQL"'�˙w�GD���Mx��w"b� 9� �=�n��9��!	��۪��$� *6Q���,?��%�7]�z�s!�!�{���i�$�4�7.h�4t��%�4�F��JR�c̛�CN{��zxU���G�sN�`8���?QK;��m�X$^
J��C��:�-��� ��ж��$O�E05m]Ǯ������_g�&��Wb�IgZC����4[���)���碿����3�}�s&��1'J�|g?�*j?Ʒ�yQ>5�����J؍�q�Ӹ�ό�⒏i�n�x�;�[����t��1/H� ~�Zt��CK*X��}'c��Ѓ�YR�PcO��/4�fx�N�D�"�@�-_!�0���p0�`#����H��&V���ݫ܃��C f��Z��(^���>͌���_��R�Y��ZP)�&e��<y����`b?%]�I~1O�X�6�}4D�y!��HFj�kg04�ص5 ~k,0?�16��^�o��T(y�n���#�p
s��m������)"\l�`'11#*Q�^X���ޏ�l���P�r���k��U:B%���@���YC��h�iCB�c0 d7Qm�"�x��]�L���g#��[�|�Q:Y��0�F�Y�|�Dp�&��q��T�A�e��<��k>�	��L�*�3���6����աFg�"��k��U��;�]�E�0������zP�{uښ4*]���Οg�3E�ru/���%5vk9l�i9��I��̂Q`a����´[a�uE�Ɨe�p�oٛ%�R��BE�k���0��)��&������j��yh{����qL�r�_�D#Ѽ���i,H��k�q�E�a� ��*$,�#Y��؃������5����<��K��u���k�4� h\�X���$e�ګ�hs�<��*�L��u���J1;�yOh���A��]y���!\�UUd"(���A�Lę�~s�Wm�bv���.b�ul2�
��@E2�qO^�������Lu���a?P�lp*_�����!�k�[/�[�S���	�U���Rq��DN ��J[3���b7���P����ď�<{�*�{����9mv�ަ��	Ŏ���Zh���/&,4�$!��~|<�q1-�����Y%�[Q|B������k���5uY*�?P�v�H� �d?H\x���.f��u����Q� �yφ?�����V�V�!��ݠ���.̜	� ���D�^��k����:�jȞ�,(E����,�}InE9�����s/�q�a/�޻׌��oV�YO���J�'�.�9�,��]�����9���c�8Y�ē#K��	S�H�8���~����Y���@7JB:`����K}�J��N���5���,v�����ǯ�h����*L�){L��~�Üٱ<�]0&5�gz�N��R������Ն411�u�8=ㄑ�('ֳ|�&���ۥ�%�����ĥ/;�{�[�e�����)�����r۴@�꾨�����f���k�dN��[�t��wbq��>a�EL� }Rd>���|A�o_���9��p����(��T�/T*�=����i�yon}TBĕ��`Mhd�K�Z{k�l��YX������(�G&6�����[�屓�W�#�v��%��PA$�{Wdh����n���(�Q��˸7:�ZDMa�@�N�n�4U׾��;��#�P�ȑ�wtfwҥ:r(� ��Ά���>_���LW�|��Y÷�fZ��-v��3�Q'������"(����T b��4M�?`�.��@Vv'xU��:t�B��Z�k�P���Ҏ�����,6�����5�m`�彌Mw3���*q�dA�/�y�{�����	f�n�K֤A��Ye&�L!��_/Ұ�H��j���(VX�l�A&|l�T��+�#�;_��.��Z$�V��*Kh�o��"�:.y<�.z�޼��HqK�(���XّJ��4}�D����S�L1Q���;����	ݘ��L� J�-�)���Q0���ڟ�����=��$��3�n�����%7ÿ̶κ� ˮ�>���]��3�(�**�VA���#6q��}D
m�=�р�/2/��^�ãX��nȬ�n�&(����C�]��q��M���w���J����o��س$��9,*�ݼ���4�a��;'�F{��zvʄ��C����'�D~��O����0��MKe�����m���E�2y�q��'q�<B�Xԥp�`;�D����7#�dK�x+l���t����⭀�
gq"�y��SˎL�TsL"� �I/��X��^�Cr�R���ۓνKV;�ѥ���4�u����#~����j�������g�_P����R<w����g�L�o�:�M�*�e�.ك�D(�"`q�-�;�$��m��1Z�:�Ͳ��������Ђ���P	����\�H�݇�:I��4����A����0��r%:�Ѕ+i��U���f�l�YF:E eo�*�X+�!���; �H��s�������]�-���e�เElg~"�_�C��T�O�ؿ޽�P�g��\��b� ��63��q�G���۠k�bv�?��K~�:(�ƀ2*�b�Q��I��!���u��WW����,�W��#���� �b������޿��hkW"A����0%�!ʗ��pZ�٩��#b�߀�����p{Oy\�&��xcB���g��6�:��&A�K
Y]�
jXG������Ђ�����(�)/�Y�;�И�o��(�$�� E�4]�49jj^˴�K+ѫ�\�ff�;�ƿd'sc�"����!Nw�{�&��n�ܟODm,|~�;�ES�������4�5e&�:�R��� V,�~���'W��J"���۟"��V�~\g���1�#s��jI�̩a�����~"�N�1(t!=�d6I����^�܊`H�u����{�w����o�m��Q�|x8
�2A\{YB!M����j��߫�\9夕���G�a"�u�P���3���F��Wc���x�>�MN�%�� ��em��ʖ ��ggs��[��t9^1]��e�i��)v�5%X�J�E���%�����ٯ ��<�yɏgю%�Z���+hkhӌ��z�Bi]�c�t�)���t�P�ظ���`X�߲C�w&�*=M��D���ڠt���'�^���f��)��[S��1�� ���ݬ �7T��[l��a0�ec�W�^[������,������AK˼�,>9)����n�h��{�;$��'�㗆K�HI7�:>{D�B�
���5�_�9��w!_}�~I���8�w� �{Ϊ
��%��U���=E�r�q�j%޷�&��l����pÛ%�S/s��]�+�>K��z{���I�l���F�����=3+x(X�ѤL���������Q�nSmL�XH�Z4|�&t_s�2��t�@0�G�н�H��B�@��#jXũC����ɍ=�:Or������5k5_8�*��b���#�(W�P��|Z�Wa���� Q��ԛ���7��]����X�wnoA_��=�E��>Z���<7F4B�Yt1ڨ��o�K]����謘��s8%]�PV�[��n(�A���L�D�5��YZ�(/��G���77.����\��.G�B�A`}�����Lj݃u/��l�莖;�-�
��mV*w���W(0l#̒c �P��#��CqT�$������j ����m����"�O~L'7��?<�&�����8)[��3�*�V�y���Ĺ4a�0_f���ކx�e6lҤ���ՍA��A8SyD��)ro(�z O)�jޠJ�2����,��֩}�Ɏj>H����T�Q�7s���)D��.Č�_�:����r���������U@�nt��%�Q�iƟtb��M��=��F`�$�i^B���p��V����_o(�I�~#]���E���5#Cx�6����sC��j�Ι��o�h=6
$g��P�{ *��]���K��S6�M��`У0�Skc���Ѡ2��D�F�tI�d�>s�d�/e%��8�s��X��g��3���6ڕ���v�/�2�'��P��������{4祖>�ja�1����wH�kT�U|c]I�
$�ʐ��Ϻr:����7�������M�5�J�i�ƕw��B�������`�@�%�U2�0���u(�e�0#'��S��A]A�ۏ�X���w�b�>!�f����N�4���{d|����;lq9��Z�I��g���)��a�]��8%$cC�'�F5���QՈl>�v��7:<.�«l�7�� ����6+mԄը^�����!���T�n#�2C���@�Y��O�S��)>6t�"��׬S�WkqDQB�v�G�����t8�N��:�K���<�c�Q����Y�Y��)ї�RS[q��b���e��n���
AG�Q�7R�^�&�#�b��l��V��7�k����_�d�g9w΄��甧�$�0��;���`LUH�TT�Z(��6'�]��ܴVٝ�n����
_}����?�w@*�m�s�ZtH}2�lk�l����(1��\{>�Е��G��<\aB����,�[X'��#+���\�6h�l�"�(�-ɳ��7A�{�w�"�E9.
'�ׅ�{	u@hɊ;\���8Ԉ�"zptٚ@���w4�Q'��G�����y2�bu���<�@.�]�Oc@��D�,����H4˘�:�A�=D�=�Z�󑉲&_�G�,�wn���g��̷�^���|��,�%�/�׸���6�ά	�g�ۓ<da'F+N�	���dV^����+���=
���37�-�C:�]�UYƘ�/M����n���"<Z��"��e]�5kXc2
��Ì ��EB]��cY�]:��=��dM��BD�^����]�B��C {�s�՝�̼+N����b0�V�^2g���T�/��kt0����n�((܁ext��^��Q/�p��`A}$��0����1��3a��J��u�������+!�GzPVd�K��6�����I��"���#������:�E��&�Dv�&�C�ۜ�h7�mB´׫�\��ˡ Zh3��y��w����9��T�(��l�-���}�o��^ٻ��,���7As�Uf������ՀN��^�r9�3���%����Cꇎ{e��}���&`�#g��Ru;#���/�ڭ�L��ebxM�B�t��H��u�b����e�ӊ��^��� 	��:�Lx���uh��l`8.!�1~�GL�nu��љ�I6�K�E��G���-b4S��.3�t+j�d��H��ʄ'�>�%��K�ݛ�^���R�J�pҗ�HĻ�яi� U�5�j6M��]Ʀ\���Il�Wˑ^�'Ɏ+�h�a3��b�*���AT�C�*&�٣�h�?*|ţ(����W �;�_ȱmK$��i�e�`�,�Ta(��:eP����}��RM��^?dDy�W�^�4x�n}5jx�Đ��9�e�񚧹����,�h�`���e�*Z�jr\a �06�bu}b�(����Ζc�U@gBF��5X�$����;'Oi�mg1�����
V�|n��$G+�IF��Ȋ|ܼ� �ovr*/E��y�ѷ�4���W��Ԕ6�S�ِ��2,��p�W�n[r���0ռ��a�a��t�8p�E(�e���b�f��M��8�����;7!o��&���V~V?�S2�m��@���k	��0B��Co�-�\N*��f��\��oY�҉AF�U����:�����$�@~�'�`�n�?��j�m��I�@-��D
e k�q�FT�Z��ct+��9|��K�]��7�[2�?!,���(J
��[pLZ;����|}^�#���]nUkܓKY��TY�0�p�p�Ι��Ѩ]�w ����}ƭ��|*c.?� �����k�4�+�!<k�?��Ǣ�c��i���_�?���*�=`�J��|JJ�ԛ�� �[�@C�)\My*=�N@ey��;�Bx�5��P��\�\��bq�9��o������j�nazĐ�]`ǖ��A��L��P�o����dDt�^���7WT��ܐ�y&~io��=����)3j��gsޖ`I�u�5�4�D�|wκ�G9�@Đ��tڌ�YwNO���nu��2��p��:3�R�zq��9�-�#E*	܄Cw�T,�6B�2��zU�5�&�=��;��.�ص����x'�9�!LW'��No� .֩.�F|f�S���<�͢�(� X�򧫫|U�S%HDٰp��m�*f����na��_�z�p� �T}<*�قM��OI���*V�X�pDݹ#y�"���M���3�Bk�Χ�N0��y��������V�g����#�p��G��,J�;�Lv�D�z;i�nj�5�~��T�= =b���fڬ�b��ž>�Ͻx�{�r�:����ܡ�YM^�I[m/��.y�Ch�SZ1s�؁X�'��kW1vg*nō�}���(�G��>>�	��Q�����4��*�H�0\B$�p�,�B�C���,�ٺk���K	�S:��Qy�2��=���.��;a��� xF[���_����?m0H�魣��"�D�B�~��~�Ԁ�K��j���}Ax}M��I��/�<?>��eur���<>S�xZ`�a���0��g݆�9b��0ߌ��?f�v/�v+UWt��3��ظ�\>��r}`����ˏY���׳&���@�?/��Q�Q�8` �]$Fd]��Py�Uug�&)�G�i1-���G� b��ۚbA�V)��^�1�$"�&�;콄��U�|C���}PŨM��(�ac��$_����������2�P<��/��@)���~	P�ŠX�PL�{j�MA��������.Y]��Q����qI�rl �`=k�(�a7O�:˩�2y����x��q�V-t�	�������Z�����Y���5�MfP�_��gD�ً��k��PZJ�v�,�	��8C�-�l�c*�Kސjw�rBa���aC�6G�I,	>�)%�P�3څ�;ot4š������KV"�J�9
]i�NIb.<���h��K� K���]|��')vI���o	m)��vb!��ho8*Yc�-*}��ʥP���&��\��)�d��U)�9�镜�z��� ➧'=���<Z�x�����n������,rPU�v�~�D�b���7�ɨb����Ϲ;�o1�|�d$���;�R�?6��ޱ�6�A�&Й�`J �U�:`%�r�!x/��&�D������ϫ.���ޒNF� �+�P�>�i0v�~��p�.�*d|�g�l"�u�Ka��޾�����rM�͊���R�梒D6T���^����lJ�a��M�y��(��Ɔ����R� �R6}���S�����^P��c�pT���	�
t.������rcJ?�tѲg5g�X�>kd���-�7���� 绘~���������h�2�iO�=�g4��'&'��D��凥L���\��]���_�m���V�٪F��?Ǜ�F������utz�ݑ�˜r�t����f������gOCSV��-r���Oe�
ٲD��,�(?}�I�ܧ�C��Z��O����*c&��>	ƙ^��!^M��z"b�2JN�=�A�+�j}�uj��sP5����&t����+�L��V �S��?
|����w���Y����h�R��~�Wc�_��ԀI�G�LR7�M����_��C�E�ԣ���&�� �`���g*�V��^�1>�4,�J,⼃�vpf�Vq��ߞ�s4:���L����.��uM�2�E����3�����q �O�k�|�f[ �,�#��vMYr����O$_3J��2��yE�2F�>��p��3�� ��h���bEI�3WSm�Br��zF�I7�c@�b+fʞ�4��%$R%'�N
���,3ۼ�_�lB�)�-+���4��Q��H	g=��T�����x���!!Zt=�la\��C�$V��Q�����ٱɼ�]j�4�	:����MTCx������k�#&u���|���C#�*�%�����'Nne��P����4�mw6��8�\=!�4�qnu�㺾�f�_�zV����6����N�G�f�q�����;	����z�S?DJ՗�������h7M?Nʁ81si�2��>C'd���Q�0�ɼ��+�gK��9GD�������[X��J��6�oջ`�f�:Z3\Yx������k�^+ә���c���=ѿ�A��_��kW@����v~��w�ܗ�����H;kټv�_��$�!���Far�D�41	�0��:g)�o������r�K�w>��B�6�yw��l~!��C">-K=?�?��S���n���ԍ����	tn�X{"\�v/��R������|ք���Y3�"Ā�2�)/���U�[wN��������Ԣ����W��9p&#jU��^�I!θ3����Ew��Z&鳒�M��b���Tn�ee5�-����=�{�������m�pD�@�П̿Y��S�� �lV�M���T��>�jDbO_j;"���2#:Qg*��3R�X��n,�o)7�kg�Y�a\��V��;1��4��o�������Y��S��~ճ�r��q�׌�EѺ��*j�gv�К�`c��߱�:r�tT�i1$Hb����z�z���3"��J�#Y�|����o����b��ٴ1�`y�����p�1��r�2z�(ku��SVZ�ȏ�g�����x���|�V#`HC5�#�}�ʵ�g���Y�ŝ/�Z�'�oI"f�E�'=��}�U����p�=pO�v����c�<�{��w5��H8ĀW�~������P_��(��ՙ�\d����0����6��������l~��8�H(��p^*V�3/���t�0��E��i��j�*b�^�p&�hC}�x�x�~o �N��D��;K)��ڔ��H7�w��� ����P�!���'P"�E҉Qv%Q3�'}*�*�(�Ӥ������rX%f��,/��X<*5�~o��عJ��fpWG����ܽ,]a=&{�/����~���B���� i�X]�bB����݉cg���̃ޱƇw/�.��o흠��qJP�lōU��?����SB_��:?-&@�C=A,U�+x�!��:H��1	J�<�V^�}4M�zӁ3�ܧ�s"�C�JnR℮]�\���V�c�W=:�n��8<Q|sMҨ$�h����H�z�#a�Z�4<TCSҠx��O:�|9Ɇ�W%]��d$p,��0���=�K|�W���#bs��O�d�Y��aG�yO��Vt��*�.��A��a�Wqb�x0k�f3�3�R>����� \��$\V���狄}g5N7]����㛨��o�������^~�mM��^���5����5���t]=�������d�ě9�Z-}�D��T�V���z�>�-���F�P�N�ys fZ�w9�Z� �D����sr�]cۅ37�����7/�m\��E�~���y7��܌V��m��+�Q�{r[��e�li,9�y�^ud|����E�;�s�6�mS��h�Qq5H�u�Η�(:=H,�vɼ�v�/�e�Z���v��6X��h���le�PxM���M��gXʁW�
�$FXy݀��m����k�w/�Ku5��#���e`2�x���5����0~gHU���D�}&�l��V����^�ez}�y�≮8D�$���NgI��Os�%/�So�E�/�V뺁P�m��	�S�]�?��5���B���[Ly�6Yꧤ��e�7��)�g�V�;#Ų���ve�V�-�ףV��2�@�t�2��@G��CO"H0kh�Ra�oM�4.���/����e�#{�������Z�
��n���ɤаk����pXΛ��j�,lvK������Lz^_������� Pܺ�g�Lz��j�s`P��R��OJߙ����������_�a��_�s��t�؜�_�u���L���]�3j��]͈��W�;89�HQ�vz%���
RH�z�𲱚>��*]�n(�>�o4Ce�Ks%��p�Fۋ,� .g�^p��D���s'L����JF��p��E�M@��7����i'���#�^�+;�9X��h�Q��-��xÑGo�4�6����������(7K����97�2�kA���"���^��ܳp�_c)��0�+6�w|Ql[06zh�W��b�S�T������w۷X�D�� i��nN������U+#'�F	�O/��u=�n�S�T�o-n�d���&qg|s��cu�}���#�7)e�<_ovH���-i>�5&Y��?Apһ����޳��4�VS�G����n`)�ЯU�REE�R
��|��[�ӮB����h�< uG3������|��-1.=���U����rg`�n�Kbߝ��/�e�\�>P	��֨H�%��aP�8��i����TW��T5x+�����"v�*�f��;X���|���ޥ=��}�����<���q������̶���6���M\?7~i��T�dx {s]I��mP�O��<�7 ��|��G"]:���!2u�#��5PY&�Q��`��%�,�,���w�$a7M�#d~9'q���"� ����c���è'���Q�t�D�?��k��/�Z��C#$�Y���k|5gjOw���C������6�ʺ?At������G�v��l�Q[�8E�±�� o ���Έ8���g��}0n̸KLRw)�P�6'�^=W�._���|h��M��`·�y�fx5��^|Je��;���Qי����CLg)�����D��6��x�{�*�H�FE�VqeD�Įa��%�U6�pp���w�f��Z�]��FEs��g̦�y��f ���rm��i4EH�ȤrG<���1����G�wt����_��NHpX"�~���1����m�@qу��EG2D�*I%�
�Ѳ��FJI���㖩�<bF���/�
}�<�klI#��E��;��=���kNI^��عJ���p�̴��rc�[�[��H�e �F<�\���H��cp�a�w�VX�֑z K�v��Rm[��S�v�����8Q�C�]G�fV��/����aB�6A�At�&�y i8�j�h���p�:�*l�,�Y���e{?�&�P�\� �➃|��D���R}#��ͯ��¶�
�١�65���w�� �3��e�jt�Q�&%� �A�o��/��̜*��FlXP.X_h)�}���'�WB��=I��T7�?�0��)P (�Լ�:�����Y�n��`�V���]����-z�M8��y��������~�W8,6�5mrS�5�*�/��w�9v�֘�Ky� �HWJn��Ba��x�T��T��<�x�>	e8���;��{R=���Y0BM-��͠$RF�l��$����IO���*�.%�<���s�͇��/��M��ƪk�ٯ�N�A��6��ƾJ��p�+�Ɏ��#+�k�̨�0X;ѥ'����2@c"UD���!�/��C�ج�٣�;��K��r�'~�j�U��S����L�R"W�?n�����M�%X�i�����%����U�,��ywʋ.,�s3��M��ȵ���a����>_�^s��B|^���B�훕U��#��psEUݥ��CY7�����盧מC}e���k��L�7��?m�ސܼuFP�˛VY�J��a�`��7���\�7����zpĿ��,3	m�����6�t6#4��.[L\���Y�8]�c������g�Ly��ۀ�q�IL?ժ��9�����(%������u���z����H�����۩Gr�O���@��*��-&lE�Qe+Po�q�Q�Y I���A�&OJ�`�p�kP?EjGG,��#!�:P��`��9��	��`*�A��§y����v.��?��r�{��?
E�r�q<�U�}�I��:���2�i�m:n�1�4ܮ�'&s9pu� k�K����a�7��$��7�+���m 8�
��������QP�~����Ƅ���S��%�C��*4�E*�9Ӏ8!A�g��߶��B镆-��Hv�����3�51;h���"f:ƨ%k��&�y�f��F�|�2S|�K���:�p�E��M�)�V�q��"��7:V7{P���b���G/�=��s�)M�^�Co�uOM�����pK0k��E���o�ge����m�_k-�4��@�p�IC���}��9��Z��~���
lz�sFRf�Z|�{!w���g� ���[)c�}�jv/��ŉ�:EP�T�Z�1�	"�W��7��@Vc�Æ�[� ��G�15"$A0(�7@I&�t����.�L��zj�/����*�Q.C,_�ufbc�A�+��Z��Ŏ��ވ���V^mjl���E;�n������6����b�FX�܀P�Y���	e��xU�r�*�y�(�e��û�^x�6.#��0�WlٖH��!Puv��8�q��W����S^.O�x �ތT��&���B�M1�hqoɖ�CW�eJ��;�����Sm-�Qx�`��?�=�oc�`��p��H"0�S�W���Ӛ\�����=f=���gx7�]/z��"���}�<���)iҎ i��kP��M$�*Y�vyN�|�$���p�g7F�~d���f)��K?��zF��>l�W�&�6j#���DC����S����<��C2xi�.�?I[�c� �\m
�1jo1�@xep���A���᪢��`;#�_�c0~���$�8���B%GX���" +q�-��[O�:�?����I�����H��VγUf�BrI�6[�?v�˶c~��B���ѹ�`�r��-�#o�v��H��iV�4#Ў��J����͖�~9j��_�V�a�����쩏})�a�(�Q��!�UGƣL��֪V��^�q[�D�J �S&�oM^�%� �4KYd������o2�Ω�Zsa
~ !�����f&�ń�C&����M��, ���Q����ٗNkuw�F��]Pڅ��bb��Vf�n:�u4�i�>�+�R^p��]#Ёc]AF)�B�C˒�||l>.DJvk���z����C�P<V�9V�']�Z��2i���{���G��{]M/��k���%��Ĩ��)@Wp�f�ƪ���� ag^�¿�'\3�A�&;�Φ��@��������KKN����1�nV�ˠ�M&���)O�Ҭ ���B���g� �� ��`%j�+�W�ոE��i���qF>����ߟ�s�g�A��_0��'J/ǰP�aV(��|�ֆ�q���׬shCW��H�����4t��;P���=0�2W=|l�j �]e�T �)�}�����Q�|-�7���`�n�o�k_�Kw�=�ɨ,MP;��!Ǭӳ����Wq[g�I��<k�w�U�y0Y����'=kZ�Oj�n�!���[R��.p\n� ŦZѤ�>���rM.�a���g��#�w�����J�)�
��Z����AZ^4��D���5?S�Nnт�b�B4�B9���`��������� ���$f�<w�v�'�&<o9�fј���5^	���`]h�A7
.��eU������#�����
���\���o2�h�2�#���ͽ.�����'AC���l��:8�����k��%o��� �߂��1}�a9��5Xۘ\+`�!�Qْh��t晼S��w�U%̍\�8=��mˑXV��f�GHS�#�yp�#����j �$��A�U�Qk�h�����=��9���~���Ƭ;�%�VH�1�;�6V:c�++"4~��0�l3��;���M�_0���Kt�)=z|Y	����u�(���I��!���wB���&95�	�i��]��{ϧ��<I�ޤ�{𼣣��r�lN��V����@�l�4a�y���^ZÛ�_niJ��du`�} H�5�s(S�u+1�k U����m1�A�nEVV�<? yG��P������ֳ2�^	�\Kd�Ne._��5?*�q�����N�I����������l������n����z�38�a}�P��,aˊ3k\4<��,XNU|�B�ٙ��m�����b�:�M�w}����_D7���E=�y��\k��:�oPw�3h@��~?�"����fӶ�A�(D�������5Y�c:]MږT�@�������>��-��>M���3�M��+/[���_>�+r���7�[���	��w��J�հx�jo@�|qh�v����%�.��~��m�fƠj!u�����,���Sɣ�5����1�T��H�!u?3:>0�����1�w�Q��� �Z��M��Gup��˄$���_�2d�'�c�S��{,[�C���d�-5P��XV�9�+Z�_�c����WZ����g��W��Tn���t�^7|Бz��p�o�0�c`V0�q�å�K�ym��C@,����I�y!�7�(�}���C?�؏=T���o�M�>z��'��NE�$�m�Z s+��
~�D6>OC$<#\*�� �i���A�a"Tż��n���Ʋ���`%E#�����$�%؎�#�
��;^�����L�fh�A��ˡ�n�W�����
O��Ae7�T��l̘o'����+z�
`�_&|��s���`��~|�އ��]�um�i�\c��m��^��6p�kF-1r@j��c.Ri��Ex��^�@�]>l����&%q=���;�n͝���"���݇ ���f]4C�+��p*�O���!}Ԑ}ø��P%@���q����������Ul�c�3���Aiz�q kG�)!�6Y�u�#{���r���6�<����W�E�3��h�bώ@�R��[vJ��p�Z�K|�ma	`RJ���샮����r=�ܷ�UC���=��R��}�.g��D��FN�B��|���i��+�>��2�ؽ�VK;(%l�V�P�7��ԝi�![Q/۪?��y`���r�:��BiޡN�SdW����9m\+ںpf5[S�Hzi���/�TjEl���xڛ*�p@���l��hlE0L�����H��tF��߿��M.k,0��Gٔ{��ޢ���p�%����n+:1!��ֱ=���i���"_z2}���`�B�z������u���H�����l�tf�&��HtH�Iz��j�]�W\Az	nO"/!��G��Ju����F�0U�/�5R���4���LD�,��+B�zq��7�c�F����ѿڣd��E�2���9�nX�O��� ~�b��}�bS� ��B[c8�$�N۬uq&�+��q��8�2��D>H�%22���ǑA0��L��<'�y�}�꺂b��?S`�����������$�ܭ�m<�����q,3����5�q�w��Te����oI��/ކ�S��A�����t�����%Ygb2���BtC�kk�q(+�i||�|��M&��jp�-_���$�78�uP|����
?O��-�,@Z$nߒHJׯk�R}8�{�?D��[�Efy�{]%�g��R�R)Q��^ͺ*�v�i��%J��P��ު���[m��
�%3d{jk�)�O"g5ͥ}=m�f�g��a��HG��=c��nH���P�3��� ��Qf.=:�Q�b� �C	��b���5������S^j�o�Ni ���^����h�m�̊�_���6�v��}��r��W�����oo�lS���(�c./t���2FA�4��	���r�1ZD��ymU�*�Zy%�||3�R���ԓ�-�T��;F������#����8@Ee�+�$	9�^v�΄=�����2�CHs��bW��2�/?<����3��v0p[�>�F�LSF2���N���S�
b�����A���@i��n�$kҺ��_�3�M��3���6���֠8�*�gEk�,��ʦ�y{Np�
�wT�,S0�1ks�q�&�y�8�_��Zm�oJ/���]��=�Zm̥<d.7}Y�	;v�A�� �!�Q�y�R��Ɗ�\���I�}�aҵvq���]pRc �|��Q��!KC|�~j�U��2�łr��l����#u�J	���7߽�h<���Ć%���]�ԃ�δVz1�%������|!h�88�� չ$��a�|8V[�AV�)0��~+.4{w&�ȫm��o�:��vGM���X��Fz�l�7K��ҽ=�����Sԍ����2�}yڽE�I��GM��=�-�}�ia)��v�/���ռ���z5�'�ր�9�2ͽ��v��:oD�ydI�áK��0���6B�-]-_�����.�q���?#�2�(�~����t���o*�;���(�;�a��UƃF_�h[f`���f�j�G�k��.�5h@4��k����"�r��==�%t������d{X9|*�`wx�I/��ɿI1]����@�r]A�g�,��J��C0'�����?'C���V�d�(�_U�Dӧw�RB2E	�U�B t'�7%��{e/��^.��U;Aͅ��2�
,��E���W���\b�竟�f�G4{Y�}���C�����|�V��������г��`bi���J.�����R��� �tW�s��X�D�P�9��G���/#A$W����Q�M�B�pD�����O�p��o"P�D�$��E��CI�^����6�փ(�61cU�2�n�����"�O��G%��^�y�D�g�S��s}Z�Vؒ����Uǀ.3���.�&X���9׼�x'�(��p0��ڊA x��ƽ�E�%Ȅ�cO�u$5x�}M��o�c�,!x���g�mۨ���0x�OS7�՗�E<��p
�naо����`V�q��)E��[��4�b4�[}���)��cp�?`���w0�p�&o=C?��3�l"�L�rľ��LC���"���S�)Q�|~w"ԩ�i;��g�'3M Y��ۖV}��z�i�sI��$����j�����Ȓ�w$k�)�%���7D���b)A-���qZ��8X0ܳ+�o
K�=
�Xc^j9��a(�;���qq7_C��%	�?�$�d�d�sŲ��O�!���MP|k�d*n��p�V6�D<�;4�7&h�/�u)8��C�}���?� ��q�_����C_
\t�:��[a�6�)U(�^�7�1s�I�,�:�����駔��Ck�\�(fNi�4�
&���5�U�ǫ�k��1�[H9zI�9�ר�׏��T?�b(�E]�
t)�1�
�=�� ����Ŋٔ��X�E��/^�r�94
93q��[29�cl�q���P3�.f��osc�	_N�CVG��\�'a�7|>Em��|�������k���^;�\��z��t�R��pK��aM$�7���3��5`��B�����2��-,�q���d�r9J�
7����^5�a�L��-&�)�_=������y��>�Yl�=mVnkP.��fE�!���r���qe������W�Z��1�lC	�g��K�'�s��~�S�ff�z�7��r��ښR&AA��1�[��?~J��I;��^崽�x^�zDW�d��ATLt�e�����V�r���D���0��3��@��O�dЪu�Z%u�ݭ�ڟ�]�N�´����So*^���&8ٶ��E9/��"���N��CU�n�O��&E��X"�9U��I/�R�v_�|�O<j�|�2=Znr���\z�؏��]$5�Ő��C6%�G���F�n�_�瀕�/O���G�����MU&�!���w�7@^1�)գ�m���Kɮ�QgB�|�k�1�c4�e:�1�'��S@iA^�Xݴ>�2!�XKtE�y��Y��2#�ȤR��d��[59��!��P���}M�2��/r��?��O�(��4��i�����Bi~�nzf3�N��ڼ1�i8�V`b�x��!)MUr�r b���.��@�j��#3gO��_9�X��F�!@3fAz,$�Z�)��a�\���=I>�� �}�R���hDP1��ƍ�6�#���dg�f���M���S������&�Y�b�W�[���Έ��V7s��<��d|hL��^[�6W�a��6�ڐ��u/��
-R��+i��/}���&ϙ��� ��t�Ӣ�y��S��l�C$"ϡP ���S�h���=9)��o҂��h�T hS~v����q�OJ̻��~��;k�?��K��a��9l���b9��P'L�
�O�|�'/�Vw��T��a�Uq{Jo|ZW�n��q��ڸ87�i2ve�.c��hT3�?1|D��s�yq��e�Fl'1w|[Y��$�x��Ƒ(����~��,n����0/�1�d�s�!I��$��G�ԥ�53l5�&���[q���W��Ø��=�����1q7?��W�(\_���F��{Dap&�V.��x��r��qJ�f�O��ϰ��z���0S\R��T�G �SU��Ur.��6�'M���p/4���M<�]X1��jqK��Y�G?zB,�V���5�Fy�a�Y��RQK|�t��p@/5��ƪ�R����NM�L�Lh��.ӎ���43.�1�O�^�ν0F����;J����C���:.��)�l�E�V�(��df��M�1
̯�;� ��l�H��|����j!Hx��h�h��Z��BP��_',
my�x_/Ö��3�]�?�➮�W�ml�(��������(N�x�AR�H}���x��Ou����i]�d��F Q'�*�F�"�٥�!��cMf�=����CN�K�D�Y�Orn?!
X6$ׂc�����Ȃ���m���Ks<սI���;s0��otKK��Jڲ���|D[�����J'��g@�+Dj���C��lǬ�dє��k"X�q����`�5f��ǹ�qD���⎦쯂{�. U��x/#������||���ǣ����5绞6�M��I�A�&����C̭��8�����WW��w50�����"`[DV߮����������ưG�x�����z
i8Z%`TX�}j�+�o�� �1P�N��%��yQ�N��Ow:)�m�����
Kx����&4oR!,֬7��Un}�j��Y
g���	\'�+xn�]B��w�L���D(hk I߁�z �Z������{fHܠC�oؗnm��[��	�.���~Ta��x���o쬑7�1�����ޝeKE#{ZY�g%�{�RW �!�Y�z%���b��8�sKS�l�J E����B�3N�*4Iȉ|���F�@+XՌ�_1�N+��Ӽ���n��\�oۣQ�c��.�|M��p���gʙ']_����%�ݫ����VÐ�mY��0q>~"����7�6�t����^��,�����orv_t��O�Bz�&��!���@%��498�w���<�5 �CHTB�Ȯ���ѡ*�^�[�^�:\i�#�I1�!�l�:u�':۬�v0����l N6 W-n�ejY4���ϫѐ@��w���ٽyIXE��
p��a��aË|�Ny`a��|U�CC�����@�$��.�\N���x��ZQ�Y!����璴��.1[�=�?,H��4K�~�T)�o=e��J�+nuޓ�9��w����&0���v��b3
%%S}�m�P���U�����Fx򈑬#���_�6�HN':�	��	��H�X@��_�$B�~!�o~���y��ml 4�Z�s����[��G���@sk���9��u�^�-Ic��4�m������e�+�K)���ƾfR}o�$�av؃���M,\n�<�s_����$ģ ���dP;{�ω+���v��j�+��E�n],�Ԛ���jb虎��РE�9�Pg�,fR=��V�ؠ�c�BA����a��'���M
�.ŇF�}����'cy�S>��>�d��� ��1���R{��p���k��bA_㽻��XY_�s#$����4��f�S�u|߷�]������H;	FZ�j���j��������S�7��oO��4��*-���{�[���c� t�BN�]�$�r4���T�=��}��5H� Sum�P7�� ���+1�~��8���cn������[�KU��f%wH.4��ʮ�͊��Ǧ�d�Eu�e�_�nvt{M����W�٘n��ߡp���]����r��c8(r��x6+3�ܓ�lVS ��/`;��9@�NC#H/ ��w�x-O�/�^�f�$a[�!�|�Y!@󈳡uU!奙��)L�WVۆq��(�N���g�����8�Z�V��ŻA�A��^��Q�骫l����\ߦ<���(g�n�3{�����@zs?�\��C�!`3yړ:4�U#k��:^�G��w��H�C�J�����!�9˺ZV�`,�mX�����P���l���GP50�Ղq�P\~�={�)��e���d�5r�B+�Ėv��V�����d��L2�Nޛ�����]6ޚC���H��X5��@��Wqj�/"�اFnNjo��
bXdwЁ/�d����<���~�D����Vȷ0��M�c��d�E�|M	m{�USQq:��v5A��&on��n�T����Q�r��:�CE��ܷ�X�ܢO�8s�hNS�/CƭB��T��C\?!�����0R�L���5����qo��!w����)܆�a!�����"qͅ@ ���?f�G�e�T<Yh�yKz;%+u��N�W-����s��� 0a�S%�	��z=�g3�I5j�:��O�� Z�(r��$*>���l��8��"���I[��3��,�7�n�i��<��h�L�o��D>���(5�q�=�2���[��I��Z3G^A�.��5š,�xܵ�K��I�8�w��F]/�d��AS�\��soŤ�&j��	8�(�u��8'n�/�1�p(��eO>��4���Fg@I�3����?�K:#$�,�RZ�D��S�O�<M��<�Ҿ��-Hv�b޳��z�e�x\I�<������+ss�@L�,yE��v�;�w-��?jtD�c�k������Ŀ��� �/���<����<@�sʤ���85yK��9��nj��)U\�� ��>��c�lw�O��L�磓��ְ�yom��γSd��Q�z��Y���sl�J-d��6 u��?kqʊ�B����A	WK�
�nD���m��\=��k�/�d� �5�,+�^9��>P7*#=��zRܴ��@N��@�0yu�c��u�/��9��[g��s��tR�,e-Z��+O*���-�_��"�;�=l�ϾX��|Ug�t\���Vji�x�B~q��
6��4�4I(w�=�"��*�(֪�D�e�J�Xx��~���r����e�Tx�5'�șr�Kgʙ�����)��vssބc��/�X��fA��er��i�*�}?[L�����	�=�S4�ƴ&�e��|q!�;;��c��Vq?P���K�#q>�˃�y����
�C,^�� ������#��n%NR"�Jh=-ˢ�vea�\Z%Ty��4���d�)EK�S�ϷT�Ô�졾��ҩ̝E�����g����>_F7�!9�g�ȴ�` я��񴋇�(!3��`��B��ϸ��M=���AU�J�+���j��f=��?�|*���>ՙ>��a�n��>	ᗘ�¹��B�8Ve�L�i��+OS	҉A�z)�Fvr�F�ɷ��լuu��V��~.ل�������XE�|k�Z�C�)\><"/�MH+�q�=:o�>��#�pl���4��Q�	�-.Z�~3|�乕F� ��l�Ds���W@I��A�F�`Ý}V-�U"ݬ�.����p	�3L[���o.~;����3(����� ,�L�������IO��:=���$Kt9%���_��l�ς�6	�t���9��_�t�����#���CEj �*�]�����]51h��� �Z���0�@ܠ@���d]��7���������`,����u�H���U�΅J1�	�N�s�.� ���p�L�Y�Xf�9���1궏3-=��E�pD�o)�(#��2�a�"01m�z2�j�WHN�v5Ё����X�1�K{�M��7��i��b�J2Q�҄�N=��'|XlB��E��19�Hƾ�g-�u1z����̑��;Bk�sv��3J� �y�k5%��/�I�~��7����x-e��{��|d "b},�W��T��螸_P���<��������� ]�_�c�6)�`1�93�魠�R�U��:�����F|#-eH����h7�Gɏ@~Pd��ʅ�b���6s'F_��~��d��!�%���&������xDk)�п�Q��`ch�*�	y#>G��O�r��MnZ�߅�5B�+h�,��wc��ߕ��y��yT����� ҽ.�֘]'W�"Jj:����/�V���0�/����F!_t���v�`��h����"I6�^ �}?��f�l�x����h��	�Rg��ŗcl}[��.q'�jM�X�-�!��?x�c�_'����X3r��+�܀-��	��q�.��?�����5��y�]PL���%���	_�֨�z�<�Qʣ���:���Q` �8z��|�S�W�|+Ԝ��?#�[��{�3�䘲F�	M~��Փq����L��H!Y��ÀVe|�˄ÙБ����o`�|��E�\=��}έ�Y���m:�;+ qz6�@�Z�-2��$3�bG�HI�t� �Q��szT8
f]>L�1�<l����Է������J,%�;�b��L�
fL�d����S1�F�I�9|e��� _G|�k0-����%*�?��.�M��H�����Z��u4�ȉ��	�w<��.�^��V �ڔQ*r3��ֈ$�1o3��ݯU1�Ͱq���H��vt&�}I3�5��sD1��'�|�7Vb1�A��}���  �X� �%߂`�<۔�M1��*��?,�ry�q@g�X��>Fv>�M����Ew]��x��+2|��l;P�������<��JQ:�S�zW-9|��?1�`E1T/]�7��(v�NemgfU{���Ms]F�sks��$i��d�&����:ۜ���M�W��	�^r�O�Q�h��v��t�Qs�o��\լG9zg�N���z@"y
%C�7����Ʃ1����)BD	uܕf�����jV2�������^R��g�\����Կ+ {L�*'+"de�,I���)Qà�c�`�,�+�C�����]O�5ƻ�Y�?��R%ȲHR�����NF\����s���3ǺEt�!@0w��9�1�DN�M3���ļ��ˈT�X��X'EW����U����1&�l����1V�'{�0�B��+��"C��<
�
f�\zcJ�c��̋�Ŧ��iU�����YI$=� nH��c�q��<_���J/$�Nr�`�[ ?v��5Yf�� )z������(���C�V��!	%{sN�t��'H�L��X���)�Y=�Y�,4N���zLnHpϐAdP�~��̈́�g�X�Z�F~ǖ{��@�=�j��q�����F�Й�*qXؤ�j,��Y���(�#�)fO�PM��\�㭤�X���@�,��#��4
L��r�>��3O]�T}���&q*���{oz��H]a>� ��E}-f��1�0eVG�eո��B��ߎ��4W��xF�Mv��Y�U90ϗ�a�@�8DFc�������>S�1�� �q�-cH�� �ͮ�-NI�/Uԝ��>ɢg���C�$UUd�
|!�㡌m�a�ڮ}���Bߌ����<�`�J��?N�W�?I>��jAҎ�#Y!Q�]�ZR�n���T��Ir+�eT[V�ŧ�{G�p�Ǳ~�0\y�¦���<�ۣ'��At$N�������|����Pf�C8��3g�yIj��)pd/�3n�Q?��ܴ��>�ǫ��7�M�y�ۖ����[<W�C;��l�nIT�%����ǭ6���+�>M����5,�ˋ��A��m�ٶ��@ �	V�S����5՘���L�����]�kV(��
����d}9l��	�JVL<dL| ں�*	��U嵞������[��o������U�M�~9*�����7;�<�.�?:.Jኬ4��D��P����Ȩ̈ C]vAb����r,V��y@.C;/n��C��//�*�U=:�Ë�̖߯���M��[�����QX5�l=!q��i�]���d�bLו�Rl3�zd8�J�g��u�tco�K�69�'.d9��@��Id�F���A��ֱ�������ĒC?�t��Vg�����aEa)�9�Y#^5���9n�7�O$�Ҵf�l/�¾A����a�UO$�6�n�k�e�!%�Դ�y߫}t�I2*I�b}����	�(�P�e�},�#�N�%��|���ŵ�+���.y�	"�1�Df���6�x,)���;�ڰ-���� x�Zn#�՗k��f���x_`�Ӣ4zfq�5y��}jgA#[�e�'V���c�{�	D�6"��?��mɫJ3q�����fb�ɨ��Q-X�HN�3���Z��>�k]�1�^�Ɨ�Ă��1�c��.KT�s��"D�T�p��G�)yg����y}%��w/Sa�w~�};ق���G�c�b=��ڇ���8}�c��JXr�1��`�V�Ďh2Lv���L�+�����b]�~1�~�u49:�Q�)08:�k�H�)�/��&�j�%}6qQZ��c���Qrys67E�|r���9Km�=hP��椯�d.;���@l2��m�M�5!��(�	��J��RS⽾��6��#�댑[�S2{�M�n[?�I\�M�QkECx�]��2W��a������.��Wl���^��5З\�Q��4�Ϟ��?,��c��τ�Q$OX�8	��3�fM��9LP�r?��.�[Y2�|$�I�]>��b�����|T���M`>�֜�ZB��9T�^��w�E�����T`�΢YK;���ڀ��H����gC�t�� �9C�N`L�6���3�j����=kI->��5WE���a�(?_nOȬ��$B(A��l&���eT��[Mj�>~��!��k��-���T;j܋C��Vu��;��xs�h��63�2�'�Z�܈�����P�V��]*�ś�����%�76�}��kX�����At��_�) ~KSnM�VnŮ�fpO,m����xvޛޞ�K[�������4�
����*(5b���3��D?��&�
�P4iR���;_!��-���oAt#�Ƣ0�ä�EN�8 ������Dgk�j_z��=J�-���c��)?�ɭ��ޡy]�rDӲA6��L�~�L���FO�Ѷ��ȥ��#g`�r�L�:�>��Xj������
Í���g_ �ek?��>�<J���oʭ/�;�Ob�ăA�1i�����K	���H��*D,�+��2�\�	�,W`n:/E��Ĝj��S[�+x*~K��"��2B�uJqjMAh)D	�v�	W�p�vOG}�c��S�2��zL�A���I��{$*N���[��$�M(���S	/�z}�c_�Ӌ�"#1C��A�m�H?[���%�{�ē0O}Z\���[�O�ݎ赮�t�)��Tt���	�9W��1��c��;��#�Z��2no�����Kvcoj��`I���x�E-�k�	�D�n���7	�j%aM���X���ۦ"\��{���� �	��^R�m�t�]����hREU��IVRI��Q�t�T�̺9&h��v��`8�YMŠ�s�� ��{�|��hÃGQt��L0���g�ف#N6ZX-����Ɂ��J�%��.Ԩ�I"mZ�j�Sg��.b�!8)�!�e���!�d����2J�+����TbE�M���I5Z2]��[0�Ck���R�O�^0��$�/�kWO��TO�ehh#�l�:#�q����A��)��5�Q����~ f�#�І*�h��`$J��2Pc)(:LɪiL8�I3��a{�K� �e�|Yf���cB	�zc��R�w��w���/v�''<�zI��Q���E���abL�܂J�I��<��La���ڐ�*y�"w��Pl~<e((m��R�m|�B5 K�A�jj��nr�O�ڳ�#Q��̰�_�&S�	��҆�ˮS��-�Ke����3nzIu�����87.�Khe�+��7�B�����k,x��^�c���'���	�>���g��j��GD�k,pe�y�ϰ��	��.���u�_���V�}4��QЋ�?*Q�4���������F�m���_�[�)�nǜ)$���iE��� �-�>��u���`�2��Z��?U���^�����(��>���`uA�������*xqK�`U2,����t��F�i?�&�Օ;��Z�s����j�8D�2��'4����Py�a�[���x�4��t��B5C�E&���q���'�?��v�IKnD:��8�o����q��
T?G_aɁT����-���V	7��2�d����S�`�9�>�Q�m�k�q�[-�g��?v������&p�.방�����]�ܛ � ������n�ؼ,�^�����< -��J�(�i�E�'vWf��	��B�<�Պ���W����n�)q`Q&��#Icnj��fq�d��F�K\���/��H7����Ң��E�3a�5+3��A���kw��eiW��H�a����)T|�㜱/����2Ya��!��_���~%�>	~8%u�x�f��sfYc�p�Y*�Y��� ��ϐ����!h���Yu)*(�0��(��+��4I������c9��2wx[���l,!����s�5�u[���b}��J �0�-{{�ܬ���i(ct����G��Ww�8#���zW�+�F���!�4B5+S�%Y�W_�u�(�x)��@�)"�9�i|�h���y�h��B��hЗ�vr��o����([�5v��[�»�Ru�R�W�DLN��E����o�/f�w����t��0�_`��z#'��l�lõū7\*����`���bI��.���}F���Q�������"B�D�g�j}��FB�fA!
z%
ǳu#��P~�����Z�r5w�9Јh��a-{��E4 ZxZ��{��"�@��֡|��7B)rD����I�0v s���B���#�`��v}��q�GD �ߑ����d�h[�<N����#��O븹�iX
�!gf]r|�q"=�D^$�ΰ:vp��J#"��`��o��}��i�8*�!�H;�����]��w�����gG�g*��XXN�����G7��q��Ʌ�eX�Bfn��L�$c�d�逵Ц�Ys@����]X'Z���# s��8������[uNz�`���}��������io���D�4ƲX��Y��h���@��B�y������[�l��Ŭ�C"�r \�����γ�e�>���Z�q�tf����\eQs���XX��)�hbYK�Ѷ���\,+�G�:����\�Έ�]�/�~$�����R3���_�BL���!�*Diq6��۫ޢi��go= f�h����M���}!S(n�[�*f�q��B��ֶ��mo3�i�s��B���I�b�D�.Z��$��,��n���I��ycD��Z5�Q4�j�d/�����I����
�H� ��Jt�Z@�4U���L�<A�&<d'kW��k@�:�\�3�j��1����� %��K�O���5J��S-�o'�o���O�c�s��)8\�ݥ{P��g��K_�Wr�"�sТW�Ʈ�x�\P�-@,�a����m�p��Um]ɣ/���8Jg+XI��6�7�l�\O�)�%}^faT7���t��S������ȸw��~�)T�������Mt}��Ci��NH�_9Ű�~��r�c���Uo���/�e�/�/]$0�(0��HR���m�cDx�lǉ�t�:�.�*܌f6R�O�bV(ng��"�nV�%�*�+D��䷊���l�h��d�=�E������!��ai��X�^�߅���W�d�ـ(X�OI~I�j1G���1|��q��0�1hw���q��d��3��;���c�pE�?c>'��S��%�*3�L�bs&q͓҉16B���iϮ�7/���$�����B��z�ݎp��������GU�ʂz�Č$�AB��Y]Γ󚲈2m�C$�\�G���Aq��/dg�����q���7	���8��k�\+�?^���K,��K�Eu^�2��R�ᾨ�����Y����F-=*HJ��ĻIM֛)>T+b#-:�--��7W���<�X�!�'U$������RDb�0�42����U�����(gI�k�e��`;�Q"_�ǍY_��mF}xG��$-�㗴�[W�(�E�$=�b؀{gGD���I$�,*�?�Wg�j�X�|<u�%�ʞ�H�9�i�������Pꕘ�ݼVl2�n[r`��,pWC\���a[�A$&�a�N��F(4|~��`�`���\���:?Ы�0vr��Х/�Cd��rMk��{"����ݖ��X���-�+��tBH��H5ɡ�wS]���?��+d��~��ȭ�9:�)�M��D�O�m�a@%����f�/a��'�4��7c�pApf�<����	�Q�4�*����%H��;.7�l�0X� F10���n!��TNf=�0��>���FE�� ۟��}�cጾ�������"�"��r�q�w������_z�>8�`P�B{�r�j�C���U��N�Jp�yV��{�����7��щ�oh�M�¸I�n	�b���0�MzB$���=���
E�}�����Lc���J�m|=�յK3������dѤ�z4��?1���B�}����/۶��7͆�l��Dhž���:�_��DR�g�8�{�V�1���AQ����P:��K��3(��Vٌy��0�aF���t��Úv|���؋��S�|kd��6is1^���+	Uݠ�8hG&�{�.�(0�Ϊ�����[a����N|�	J�F���w7�<�]�H�tZ������d�J]R�aw�	�T"����`�1��3+�*Bv��}-����k�7�R�F���{�׌�Vc�Gn�Ǭ)~�H�Vĭv_�)���Z�{c3!�t��j�h k��+�k�?f�ƬA0 ���;����za��Y�HU�T�?�����M�g��BU���g�VY9>)bn,�]�"���{ ��N���G]�%^
� BԂ�n�Ar�E���N�K��?.	ڶj#��SI�\��Y&E(]�Ί��v��bV�ƺ¸&R��ڗ�m�}�IR\YkYĉ)�k|)(z�=�[=��g� �}���>�G!B�^�[����x���7^��K��-����/�G(��-
��n����`�HJ�E*QXY`���>��ʻ�Q�<�I�y����W���Ny�W�DU�#�y|��3�笏��[�~�\�L8���}��W<6��H7PC���͵޸C8�����k�n'����	?[�6 %�SA���BcZ�6)7��O)Oկ
��^���(#rX���=����+�4]3U��
v�W���w�,�x�?���7oe��Y�v�b�ϒ�k���S�3ei�I�@�+Vz	LUs��O��L'�EϠ��H0N�ŏ�II���K��Q,����:c��E2$2@�:�3h�OW�o�9W{`����GU��v�(��ѹ �X�GR����	b�.]˭wo���&t7�oL]�8�
r�;B��9������@��8)�z=�w���i��m�wJӮ�����up֑��c�fo�7����@�����-[���Q����vel�%Y�K�M��N����V� bw�3f-���(���¶+�L�R��t�[}�Ѳ��%����=���-���� �c�8t�q��4%=l'�5����x�D)<x�����8>8���[�xn!SH�0B<�����Ik�.T��4LǄw�O�.u����늂�A8Fm�Y�6'ܿ���B@�'f�7��$V*��׾��R	�Z!`��wh>�$X�~;@�
�9.B7��Q2�j���(cly�ó��HC�l���Ւ|f�6J�m0̵H�~s]�:j��BPC�N�����cp�{-%�� ˟+�/j}�9�a/cZ������j9�NiY����P3�=�Y����8eӚ���	`�A+��3 �á�e�{	�e�(�����Wn⾘�F�����11s�/��T�I�ͱ*"�����QBZ���ӛ�sK�MbT��ݏ��� �I�@�� �����V��[�pQTly�Ũ>٤|�w+h��@�n+�Z�#�h0p7�W��Fr�����+����o,�ĉា僎�YG�|�i#jw[����
�
G�k+`�b���)wp�0����L���M��jFpJ�i:���q�����$Q)���!���=��L��e!�Y?ު����L^�zz48ՕӇ%h���n3)x�c�t��x�Q��״��b��~π��᝜�ĉ>a"xݾ�o�m@�9{&���U>.��Ɨ�<37a
�ޮ�c������/Q��J8)��%��l��C��\'�&QDQ\�&Xj�+j>5\��+����Uā<cT�sKE�1����Ṯk�{�;�ו,�9`��΢ƦY6�v뿓��Q �0�'Z�r�Z��լ�Q3r\�X��m������1�H7�)��>J&S�����1y75:"��TZg@�|L"�������>��0�̤�s��Oz��@���H��(��=~�^��*(#VgŊ
���o��n(��w�gS"
P�@pC��
�SP�;���&Q�b������l����2غD�F�^��to/Q���>���1�s?�7���zǝ�׌�£��-}�0�U+��	��jO0;� ��{��E_?�8��[����ģAC��g_}}��:���M�Q��p�M��zv�'��x����|z����$6�zL�G"�#b<ջp����Ֆ�e���V�w7�O�f;�v� ��?�����N�+w�v������h�϶�l8�軜��'/"/E��",�P��lH���b���� k@���}^^���]�P���������$��� aC��W��J��;�(*i�����P�����P"zpYԕ+2��n �p�4���k����l�T�X,�p�t�Y�H��o���p��x	N�'=�4m�i�.7�2�J~���UD��FRЇD�����U2��'�� 6T."�Pv#+'�D 9]�O��d�a{��xJ�s� \8d��Gf&���A��в�
��E� �b|L�꿵.��
���Lt�3�2�fo+��C�iB�H@u�,�a�7d)/t��g؛��s�g�Ӛ#�TE�^��N	k4tYq�3}��,�xty#���s�SJr��߷Ldʹ7���ZD� rM�	��{�������Q�׆��U�_�H��=�Ͷ���Y��RE�����󃢭�T��C8����Gz,z��־j��"ޥ��2g��"��K�g^���~9��9�Jং����$h�H�׮��d� Vy���2�ڂ��V�v�.�xe.�}�at/dN�HxI��
k�4?�t�g���b:��S��:/}�K`������m_Dh�����M�j$^L���C������#H��4U�NҶZ��r�<�O&ݹ����%݊P=�*zL��Wݡ��T���ދ7Z[��R5Q�l�o��@���0�V����.�n�����(i���r��f�͑F�<�N�U�f�4���`����B���f�@�Z%|6�U��~�ʋ�����U^�m	���&p?PF���=H7�H_-���|Ny�/��`��pYcC��m!����<9�-7���f�`y�����q��ln�RJ�ƹ���NN��a�덀���^��U	�e���X-�Eh��w����5j��#�0�b}�)���&�;����h��J��(��!s�j�5�E��1�@��HG�IA,�"�7���6b���r�ă�kz2��p�\��BG�V�D�E�#F���\[�������ǿ���IB�$GP̩��!���ß^������%�]0���G���7x.h��˒��L�+&2ǍO�P�8z���W��K�*zV�R�	�v��6*/A�h���g������{Ψ�FH�P�
<$�X�X(��?s�آM����x�4]`o!��C~��M9/sb��VmA���"����֮?Q�^�S@�V��g�0'�F\n��/w��"���*��/S���&> �(�bqr�a������:���'ə�*�:�L��O�`z��+����R���^���dS��z`�2H����Aro׷\���:�:2��^#G���6�k+��T@\�}6��0$���Zf��J��|\ ��T���BB��L��9v	��I����g�������F��@�λ�>{?���Ƣ�W��էI���v��sqw�:��{E�$nG4y0�z�G7�C��Q���J*s���a�L-�B��M�6��>��-%`I�w3*��%$C�����5RCX�s-�c�ș�ԡ*���YH^�	�gy,g��隋������YN�/
I�YǞ��zK,�i2��8�I'��V �3}#����ؑ·�H��/c�b���t��J��
���a��Khj}�Q�H�x@T���+�g`Z���!'´�JX{��\3u�y���W��TU=�+�@H{[�3�e͈�����?}2-ߛ�ew:''�ش���fk�h�F4C�܈{+��I�~�`V���*��F�H~���#��꽸V���NH8\y(�41_^�r���_���+�1�ʫ�Dwg4��c�KF�;�7�c΁d��,ށ���z���.�~,���7'��@�g�G �S�a����9�:�×���Jڼ�{WX��Z��d'I���u�v#g �>,�kN�����61n%��9:[��\O�	��,BC'o�ql@4�P~����m&��e,����No�Y��o�^�"�|�i��1�3�������W�x���CQ�ng�5H�IKu.)�cq_���%��O�����$��!�.��%6\d�L�,�x	dto�'x�<	=IZ^lH웧��,9��4qI��L�#>s�f��]��S�%��0ܦ�*��4�b��̮��z�\
�b�2]��z�x�K>$`fdE���a��]d��Rq��s��6��$+NLE��}�6���f]GU�:��R��j#�NZ�ުW>�_RW��}.�وJufE�"�mM����PAC���I|�S"��δT ��ľ��<˲�TB�Y"U�87�u�L���Т����%�?]*`�Z:rk�˰��2k�:�2���ʰ�}��T;��|�oA&��FD��p����0�m��MM'���d�t].�HŸԗC�T��Ў�r
͍��!<���|��xJڼk�;*D�)9p�:��p���@]��6�ܧ5)��<�K6��wMy�#%՟��)�Γ��L������
?gb	��ܬ�S]=.0lQqNb���U���f�UO��Ry%����jN��Fwa��.��*��MB�b��F�������LD	���_�lʲ�ݾ�(q��b��KK%EN�}�~ ���c|M1V�i Nu"�H
%pȰ����: ��tS�ӑ�n�h������RC֠�0�.��Ռi-V(uN���>���F8�u>|p�m�h�HJ�`(�@�<}��+�O���fu��6�A9�$9�7o=����A�����&��<E1�m�J��Y���!&��[C�����(��zgb �d5�6j?U�c�_~C&uǰ�V�����P��	��W��\,\��r�M/�{f��1��`|6�eB����N@��?�����h(n�Jqz�Y��2W#Ky���~.��!����	�S�1_���}<�_�eC��	�i�7b���;�[�a�Rs1Z2�f�V���?'z��?e'rzR��k҇ˠ�h`cEd�H �ljs��Ns���ż]��.�����o�睩���Er7Heh�?�ӸaV�/�UzqB���]���|�,���(�Z�R��Jj�ù�si�Aѽ)Coi9�|]����;�k��!
�����ܓ���Cjr�K�Z�,���,N���eq�9潋���EHb+�n���>��T��q���3}��X�?���џ�+��9����@~�c!�2+��[��xn��E�:y~�~� �G�1`���a4f��n�V�>���+�6��[���h�6&'௅m"C�/C(`"����47d3�J��	�7��G,�/��0�͕����䦘��&�s0
��Kb8g�L�J �)���ơT��ߐcH��koZrd�|����@������N��Ue�#��t�VE��Ib�Z@�/�����@�gýrK�S�p]�G�"_�'e�4�a[�Y��h��F�t��'��� Ld��5F-T%V 38��Ղ��4.Yv���o!6�|��V�2r^RqC��a����`��|�hi�|F�	�>��R��_��2Z�����z��ޭ_=C&J���{�����9w�H�D9�.��W�i��q��3H�����i������K��O�X7���5�+Y{����ct?�����K�[5,,�'���+{�j�[ �}�;�Y��
�xL�n��A�U��t�At�_P��ت��`\f�rB�	ہ�B��x���%�o��u�7.�Cq��ߕO3�(j۸,f  ���.L���[i��u�{7�P�a�iU+�r�&A�������H�<��a�d��:Z�K仅ϫ����jZN�`��E�2�Z��IdO	`�U�2y�#r���eҩ k\N*?��x��ލ�����u��CYbk|�9X���qݳ��Qj���/��`���.����Y��E�/��-�[�� j�++���>�em�ӄ�@^g	����'h�9
Nr}���}SLz�2M�!��Lg�h][��`	[.eX�@����T���2����V�b�G��H�ݻ-qQsF��rX���
�V����{��T+q�dO+�� �wS��,0	J-�����<9j��7�u�X�p_ת�CY��g��,c:@��z�-W�b2Tn��P�k����:�k�3o:�������n�/��d�T�M�U���c�q�/(8�;��(�N�l�^j�:!�
@[���a���7� Ҁ�w=FTUZ"4Pi<rM��iu���CXБ>��ġ4���\O^�~X�P��!&�y�I*����Y���󶺌��w���M��R��w�)V#���6��&p/�T0o� �N�1T�0##?rU�����c"+��9H� ���$,H����w��)8���P=zY��j��:oﴟ#�"�U�)��E�f��i��T���£`W�)���U�P�w� D?�y�1A�+��_c?^��*α�Iv���<D!���c8���+U��oP�a�4ܒ.�u��j��2*V9ٸI�
׎�A����q-7_�F��_m`m�郹����h�I���j�j���p]����y��oG��8�V<I�H�YeQ�G�0��8��-v�1Xj��Fr��#����S�w`H/�6'����|��Q�wch��p�οm=ad�.L����0�ܴ��6)̌i����Û�2���h��c�u�!F�%!N����:?ۏ�С�����w�������JŬ_0�X�h퍀�{�~�<�~{?_ AJ���p��� 	� �e,�p��qQI�������^�W9�v	����t�t�`�9��^��y�ds�A�0Y�řG1^Rf��!6n�=�y��X�,�i�EI�qW߷��%r��0-R���'�W��Ek��ݻ��i �)!� -#Gl��o/Ֆ�����U�2G�R��'��V�C�xq�����0]#�o��ȖL���p�E&���Cj����֣��<���G�ܚCu�Z�+�h٤��ߞ�՚���s�7�<}���W͂Nq��9s���Fb3��n�b��qyC�I��g(��
o��h`Pt��h���Q������]Փ��62om
�:�q;/�A�/��pTG�_���&��0��T��l�@C互6��:�L�J�$�;�Q����0�էb�$~�xTi�P���n>��
��&�T��o��f1�Z��N��9���rQ�&�(c���$�m<� K�E���H�1}��s���VŠl��)f۬��rT�::{����@MN�	%~P�#5�$g��%�x�ST$S�g�5��5a�֗�NB����m0,��Kx�5E���c�V��9�e�W[t�臿��&�f#ǉ��gZrن0���(��ᄝғ&��<�(�YY\.ʷ�I�&�1o��]�%?ډP=�lS���i�n��<La�:�J���_�a�/d�h)x�qHj�^�~|�`@�ˀ\��6�I�2�dΌAE�ܭӜ~��?����5��a�5������;���#����\A;�[/�5`gm �����;��'H�X�y]���^8���]�[Bd���{�e�Q��g�m��C &�T$O�G��
��*G�E�\1ë�L�����g�|�:	LO#�q9�w��I�
�l8S�D����^1�sC�`�/on/y�ц%�ګ"����0yuJ
g�M��Pf����}�#��}�H��w�6B�����qMM�h)��e,�,*2��?%�'MkU�0�dҕ��W�Myw �n$s�m�K��V��x�`�Y9����Q/UYj."��
_��p[�j/j�g؇z2�h�~'�CC0P%�^@~�Y����:P��Z5��&?2c����Cy�W'���M9x(S*-��zv�R����)�R�#J����9�	�_���g	d�ɷN�F�@p;A�fw�H�?H����A��Hb���L"d�(���r�E
b�#m
���LJ7Ƅsߙ��N�<Fz�4B!!ɬ'�.���Ay�+��qDpr�u�3�v'O|�w) �r�#���=�{Zjϭ�)�攍�f��6�l��
xN�h	��<_�>��/헾Ǎ
��CY>��oej�0�К�"��u��Y�%-y��.��0@���җ5��jy����-�E>ԋyg�ٻ媳-V�^�ꕁ�	����ҽ��CV A�I=pk�f;c��UB���y���>�� w���}4K�YX��Ʈ�����5�w;�p�P����dr�X�,p�4�(�nښ��c~��.�&�av�=�~R�V��l_a�/��lO�va����L�Q�d��4�S˝3��KzM�4��T���5�c�鵚��J�2��:�CK�cOe������/ ���'���i��ZAv��Vں�l��{f�c���u#�Ү�	�!�r�A쿛:���Q#>��G��=�>[���ɋ�][����spٞ{�|�D<�󙴣tI��ry�/ٹ�a섾y����.�� *2tE�t��:�x�z��\�a�X�)�����C��Hܕ6�� ,n$V/s�����b�@l�����os,��K��eR�>/bV���d����0��tt���=v��@��q-%-�Gj������Rz� }b�F��`�����rɢ����ô	��3Y�m��K*��&�P�<d֝��¿�
�Ӯڞ_ȝ���9���ᵬS��H�d�y�Z5{�c�Le1uzȻ���@�3t��Ŋ�H��`�ӻ�Y;	jr��"t�+h`���.����Sף�+���'1�'ڞ]֙�-�DWad�Ny�.�}��;Ʊ^������ɦ�&�`"�&t��bC������y�D]�g���5f�������J)���:n��!=S�Q��8�7�vH7���5?,��Q�Z6����j�'��G����z�z��ً�����p�)���h*�K ���@���W�|NW��,��Q�{�-Z� l���͕����I���& �D�'MU��W�9�;���G$����y�V�s��LN}�ߪ�����4&� 6������*����'���d�[�cK���GIB70C��=�;���k�^��w�8w��ŷ|�P0չz����ba8%P%(lp5@Q]`Ŏ��i���+H�B���=w|W"�|U-b{�fP�� r�z�U/�)3��\�F~u{����\2sJͲ^���R� =g|�A���O|jy�����LۺA�:A�	�K7��������%�p�Fס@����wr��Dh��٨[$�z�O���{�������uRg���ݐ0߂KR-�u�fņE)�0-��6/��ׯxp�e72�'��M����>5|_�NM<>hlg���B�R{���G�8�,�9a�LCL�o=,e�PӁ��+�ԫx����l�7q�C��$�ͩ�g���#��m����j���͓������#bǸM�<��Q����%�{��l�5ħ�)S�]���q�>�8�NNf�)E���-���a���;�9�XE�#t[��7)Ң�u7���`�� �i7�1w���t��_,$���A���-���60W��V��Bn@�N+Z9n4/��T%�]q��cXz�� �S���r�'���_o�/�2t I�y���4#�;\
\�j�_�9��׃H��w���;�8�63y�U�N�:��� �m�jL�=|����bO���j �s�Ւ4\3���%�p�<��u�$�'�E!@?͝�u/�٩z]~D1&o��,�!��9�j�{8����綽���r�j��_ŜfP��!�v�b$+Z�[h��AT}��HĂJkx�<�^j�A��*�p.5���&��5Շ;`нM��*`C�)������V׬x6'��{�4@Q��&�bL{��9t'��λ����mOGQ~4G^pϓ�1n3Nʇ��N[�nH����I�X?	��{6x<|5'<�s�ZU�Pi����hB�ÿ^`��mn�`���uW�7mJ��{��A��Y�Jd���g�#<�n�w��*Bi��E����wlXf<��H�1��h.��.t��N������J!�so~��U����	�X��k��R.�D�Ń�?P�}"۠�&O���]���b��d����7r7n;�C����M�k�췋�4����wߤ�/&U����g�%��eJ��5�jۉ�5�����Jl̠��͍�6�ܒ`�I�ƥ7N��Λ�Ӑo��bEŶQJ�h;Gػ���H"�|�6�m3i>_��'�t���w�LD�_ ���o�k�x���h�g��%��?]i~Jt����eb������.MG���h�Ν�2��}���tv���#k�A\��W�66�fV͢6��r-�i�����v�[UsJO~���C0G���V��ܶN�mR���a��;ŭ�E��
����I� ���'��K�k���LJ�o	�f��3���kVg�Z��P]�C�wN��r�:�Nĺ	:Hߒק��@(�����yL^�S&�$��� �&���X6��;���Dz+�}�RN�7�r�R{������ �-�C�[��e���}�Far/ǩ�&��6�C"aT���_�2n?VT!0{^:��x������~Z`�T^��Jԃ9Ʉ�����^�P?��2e�>�����������fo.��F)"͝���bOs ek�"R������$RF�j\"Z;�
�݀v⥩�����.7���d�`�iw�=Ύ<(�b��
��A;[�SB%9A8c!<�5����K���/Wʱ���F%;�\�B�XY ��0�s����_3��2���n�	��А�����!�0L����_��I�9��HDf(Qϻܸ��#���O$��?��i����l�,����W�*�%�\���h�%qՒ����H��`Lws�v؆�<;83�PUS�sb�(�_5���sn*�܎]��J���<pja��)����_d��]]ؘ*[	Q�ZO������:\�f^� u3�=�`)GX�/Ȯ�Q���W��	& 8
Cz;O�TS��品�a�����]�w�I6��|q*��ѻ����� ��?<��hpK,�j��vn�Rn�e7����v���/ġ%����	f��'�Xz�e���'VJ�w�x��(�z��'�!3P��6����J2N���t��m���3�a�Y$�n��EN���E��?\�m~��"ר�:Ԏ'7�� �$Ѽ[5�9��{$�1i�����Om���)��r���m/���W@
s������d&#6Y��L�pým�IŚ��sf*ֵ@�	����)*�"�3���[�q&-��G_�Ɨ"��³M����v�]�N�;Ro���s�=�����\�%Z��V�Õ8_p8�͏_�2}�J�`4�$�q�O�g�!����5��I,]�f�,�(��8FC��>��u�7{ڀJ*@dOu´�gg;L�炐l[fM�Ӭ�w"oe���xc&b� ��u's��S�?�~�i�{v?�0�_�&��
]��ܰʗs�l�dmw�7D���0�v�[#%6
95MF������U��ʽT�FOO��&������˅,<�<�q]R�/��Mu�,/��Hs�8JF��Lg;R�����������L�� k"��v`
(M�l��5�����N}X�Q�a[` QBCcINk���Q� �5���+��I.r�;�պW,�RE�iBP���	��7(�3�E�^kzF!8�n�y����TJ�&]�@Z�Y�E�����6� ��	a�M�h;יPQ�����4�FN��i'�ʉ`X���,C�ޠq�����V�&�ɯ. ꏨWN�/KkCCK�B�wOܾ�C����� �Cд�G�e��L޵���$M�Ӆ�3�e��p<�`9�:p���N�:'N0.u/������<�$�5��u�HC���V���І*68���a�o2�!b\�zkU��n�ݡ��02p�E{����fDgbr:9@�D3��L�|il���[��A�=���PR��T��s<�b��;ӳkʈr���ⱶ���,i���ps��8�Rs��5���7?-�7k�2l�ZN��Pz+����6K��ɍw�<~M��d�� ��(CR6�=��2ik�bT���,�t���O�N�x{6E��2b��`X0���`>�Ri;���|�08������PU�7W�����}���(-m2��Tb����Y�C�(&��##�UIAV��YD����{���_0#�@�4�㎛����eн�d����WO�3ks[��Q��$��j�>i>D�Mw�8]����M��7�=4�c�\��B����:�O����dU\�2r!�G��`�A��~_�+H��Kj�`Ͷ��݋�%�C۩.�.���v<����V�b앾M���FQ6F޶rG0��!Zh^�$ �05���M�����K�:6q�"N�xԙa*fi���D��XÙ&���E7���6^��bQa��Iǯks�f�$����{CA	������Sgn�ʤf��7�0�lm�g�Vυ2�w���[��S�8D8��0�"<�$!�|X1�[���=��o�Bk����A�S���dh$�����O��?�he~K���K`�(m6����EN-���k��H�D�����rY���QA�K�%�1P�Cf	{��t��ex�N�#c�˾Sn�IJ��)���<{�ԓ�k� ��v}�?���au��OH�q��~)Ֆ	���j7�o@ʃ���� �܆�L]t ��:{��\�Ah���i����xz<|�-��k��U԰�\�8�G���&)sVnڦ$ �i�z�n�L���;Z�uE���U��@���	t�q�8�b<�)��n��?�M�z��p��N��`�"Z��8@n�����%�a��w�o����������p?�8�r@�u	�@C�F��>����U�Bd��X8I���1�\�^�>L�"X���Um.Ē�u+yEZ�����fӛ������K���L<�>#����0$?W�)31��Ϡ[�>�7�6��	1Y���Q�_�d!��sIq�_�z^�}I��{y+\E�A��R�*X�@�����nY���a"*��n$�l��!|���]�pQ��jnz�$c�f滂�&�	~3���z���IBb�&�LDk����4j�zJ�a5�� {�#{Ow����v�ߴ0��]���a�B$�����9���9�P܀��p 3M�8�T���x)ؤM��kX�������-hC�Q��������լ�@ ᯚl��-4Rz���OMȸ����|1V͑�nxۿhh�*q�OU��uLY%����}Ya.�� F|����K�%�\(R�k�4��4�ۋDծ��{wa�h��"��|�����2@x>�ݐ��7+��;Cϖ꼣a�/t(�1�1�E��1ԾC�ꀵ"�����T��/܅^|e�m��_Afq-qT`���z{
��9�-�Q��nP���"�7a<`|VR.���)+�	j�����^]�������)�D��m��H��Bv4��qoZԙ؃~�*c�����M-|%�>v$?q�]Haʜ�4u3=z#��_��k��~F��O��ӈ��%�ĳ5����
�	�3�	K�V�j��PPxzQʽ�sY�[���:X#��{j�>Y7;��beD��Q��7��*@u���<����ɕ�8�gRZ�	����*�NO�,���2Id�P�;KP�X�.m�XtN�ϲ�M�7���|+��P�$��x5�'��*�O�DX�J��u�ko��tC�oFI'��ࠍ��]f�p�~�����w�D8�)`TG�\���.���$�	�0]��3�������!�P�n?�ٌ�D�TiB�ν�A��A����$�Pr�0#����J�e���z�F�Q�	�-p_�8[91C'�ڦU�2akɧo������E[��{�!��ޡ&�H4�.�!�3��&� -�v&@I2�4�@��i4�Va�`��܈�m'����ٸ�ncŚ��n2����}�l�+�ھ�f�ZV<�&�.�����5͕�ͱ)uݽ{���T�I.�2˜�>�[ʱY��U�+��/�m�g��v(��́�����l89��W(��5*�8�p�pF��þj�z|���3�|�]8����ѿ�K�2��
͟���C�TQ�Q�����Y�@ .�r�Fz�>g%�Y۾�I-QhZ"�@���ה����;�m��KM�n�����1�<��~.��W�'l�\ٖ
@l�rh�]�G1�3W�ȧ:w��<*A�:>B�p֊�fb�S����(���3�it�KiX�k¡1�w�w�戼�´Y���	;������,�ds������O�t �ᚫ���-;�ު��;�|��LL?�f��M��iq�7S�1wS>�(/x�'��+��m[��B��M���%������Xn�Ko��Cx���|�-7�e��tx��xض�Y�K�~�B��Q����g�_�_'�GQ���$���i6�-�1m�Mc��� dYR��&-	0�2��Ow�HKb�2NMZ���`�?8A�9�W"�h��f��2_i�xY4�T��)�u
��y�=jl�A����_\kjY���ZL��E�&��p����5$5�[�v/:�'"�l鵛���Kk�_'躍>'9߸���,2����b�T>v���,�D�48�]j`�&Ч�]�g�� S����������l1�j�@��R\���Ξ6?�,�8�B�̟���|��Y���v,�(֨q5�=W`a5�ۙIEa��h#�l~&չP�� z�6����w��I�R��"�$��d�h�g��:=���W8F�5OY��2�!��#@<u@o}Ҥ���]"�m����x�s�v0�긞���K010`t)G�r�a�]}C!�#x��]�n�HF���d�pe��"j�`X�Pe;}d��b��e��,J�*��ȼ=�����s�� ��.��	�V�i�3��b2�L��g?͊*�5�o��O�C��E{�}!4c4���]~��O���|�ŝ��Ν�}z�|Edw��,+�n㚟�*�8�0#)��=�X]~��\o`}�LK�B}Q�?ܴu:����×α|�u��韕@zqV	v&��9Q�xf�o�; *��sw��(K�ٕ@5��NX+���dr]sHܛ �ְ�թ2�zd���m�4:)���+q��yu;w,�eۿ��[�ń$Z�`��G4�Y�}n���DU.K���R2&s⿜�'�-�WlT��2y4�>�c��x$��I��m���b(qn"�P1���Z<�#������g/\��k�A�27�i#6"��s����Z� zV����d�hƱ��0w������2���m%`_�g-�x3ɭ%5�=_�ޙ�Ez;��I��h:�l�"�\*(���w���W���� XNn��uB�Sb�D�_MBo)����tˋ*���	��Z�M_j�6L9������{�n#�3��t &+���ī�B��(2�L1�= ���֠���"���Qf'X�n�p�u0�y0V��f��H����S��|�)k@`S���k��֕xvK��DF�u����'�=��j4wNò�J�� �;]�i��w��s¸b�$��=��v�ZN7ClY�`؍�"�u�� ��y�LH�wH^0U� �[tl�D�I'Ǧ,^${�
#��F��ܨ�o4�����t�y�>nvGB����/�@aP_C�k�Gq�u}sb�˗I ��ΟF���AZ�ޝ%nW�"J&��8��������K�C��Ť�H��y�$��<{����yq�⪲�÷&~�n`���K�f�}�^[�3��e�%���s��ܼ ����������U!���J��#�T��Ohf�qǴU�ocL�4{��sV�L���O�V���d�W"崂'�lq�S�s��3͸R����u���
q�$I����z�d<�%��������H1{�;b���S��k���\(SRqa`���0�OYq��()��.��3�\sO��܋$8*1�z�,��%��rsF��6�x�	Fk��pvv��䰜C8�ڤu����^�
YL�D<J|8M��-A1}��;���XG&�Kj?�l;��
3�ol��9��=�_���>N3��N��A���&��-��c�J�{�Ikj�:��k��s����)e��9��v��%(�s��os��Z�!2��������� �9k����8����kܹ)�6�Z��葼�uup���Ȍ��Vd#��� >���h��ve���-���_{�bR���q!��ߑ@�״*F�͒�YY����#������)r�Q�� ��c�H�����Fm|Ut��n������<�����\Ŋ��7�)w��Q_ٵr�Z��3-���:�3��B]q���f81�L�q����E0���gY�R u����w���-������ßN�P�b��#Lz��,�*U�� �Y�xhޝ�-�P=�!M|i��`��9Y�	�����ښ�c�X,��L���Qg�2�`����W{bs��ŧ��cR�hjj#Lc0�}�{ʓt�{����.>�h�r�s�\�Դ[^+K.�>X�#�Y�,�5��h��%�6���o��ǺSl�1r@>���i�R���>m��K���ъ�H'�U7�Ar�m���C��SCe3�Dn�[��f��`,��Li��j�z��,zpT�v���j� )E����W�u��D/$�����F�p����L]�"_/*�#4�&=g�9אr��5d�NN�B���츇_�÷�u���*"��v�ۡ��z�e�oYJݛ����Ԅo'5��a�.;BS���_�nl�]�ݗ���8�3�qɏiL��*Q�I�A��n8̞�oS1>�P�Κ��H�t>�m�-CQt���@���4�C�Mr��-/����\��)5x�%9�������`u��	���ͦi������B�yJW�tU!�m{	ZzF&�2�0R���s�������v�
o�߀��ĩ��V8�;u�N"@��9a"o:���:�\n��+Bf\��>y2�t UO9r)��
��1�3~P�Py
��� ��LѬx�@h2���DQ���D48�tLn� oe;Ƴ9>+��+��Ԛ8$�SDT�h��G�H=9�d����j̬��B)����8#��*b�:*c������dn�)~(`��J�[|ڎ��*rq�W�Q��r&a^��;��j�ZT��N��l�S��0�b���Z��l�|�F��t�j����w��������T�ܵ�u�����H��M���9��ԓ@R&I�}7R>�y��0���{1�6��S>#�Y|CX\�Me���Bˤo���%��P�r|
�3t�Y{�*�G(7*I=�����=�G�w�Jd�M�a#��X����Y��@�O��h�o9���s����A��OZ���m�o�fx���)^�	UAE6U��~^���@f�L��Є���W���S���kSaw�"<:Oi��j_;e�1s���䅪ȵgQ,K�P�h���!�.'��F�֥pH	n�mA�SWu����(ѻ�5��j�k�jp9l,������K�lNdᯌ�B��#L��>si1�q=�������K~�9O���[��^��+m��A��*ޯD[cRv�nl���K��zd
_���4���H�:�=�#���'����jz���Iп7��>C����	߆��Q�Uj��i�ۑL7��"G����Fs���qlՒ��m�p�Q�T�>�O�����"`6zW��˵*�j�}�9bm�.����� -��H��p�,��%�ѥ�a$_̈�d�D�^≸C�z���gbeF���>�5TF9��������������Tx2TZ	����x��L�Ƀ`
���B��?:|N(��ܽ���K��5��#��Wry�|�	�z�
��h�yx@��0Z�]G�:x�g5D��j�!�*G�q��׫�v���=:� y����W�޼�_�W1�M����O����\B���>�/�4\�%������k>K0���hq |#w�s���l�W��w���]�A���	����^�d
F\D1���E����E���6�}�h���K��<p�|^���>h<�Ϳce�U����
	L%�fy�S515�{ԅG�Ya�A'<5�)����x�	b3�kHQ���L7ʆ$��F��麩d�����nd�aVfxV�ӷ8�	_A�]�5�r =Fg�=@����H�|�$!��+8��Sp�	l����uϣ@1��92�;(i�!qx]Ew�
�_�@SYN�z�{@
-��$8/�2*ݳQ��i�*�YL7oF���˙3�گ*�8�:f�6p�|Ny�S���.��Hc�2E��7�ѓ�F��
��tMen���@"��D]�å�O�8�rf+5��0�
1p���J�n��4z�]���>la�4:!hiʻq$y���t ��"����)��Mڦ~1�볞�Ȍ�e�F:�8�� ������� �u5� �p3ze���������X7��tl�S4��;sZ�|k�ׁ#������pT�J����?�"���T�&��*�l�i-�s�:�(�z)֞g��Z��Y
�E8�m`R6s�þ1�?�~ɛ�g�-�R�Cώ��j�n�c��W�w��{��2�
�����0е���@�}�̛f14��p�'��BH���2�ZU6�N�ψ��h|�-���_ߗ[2�]��`u��7t�oU���Q�o�10��0P;�L�ɵ�A�V�|��y=�e4j#��^�{��:��H����3�(����0��*�v�P��&U���Cn�[�аg0BC�Encj�hE�WXAĘߌ����-�ou����oO�%�k����������8ZA�<�(hsj�(�7�>�zo������{}�i�뜜��$.���c,�$�F���5���=��:2xJ�}]{��`�M��5a�㽙}�H��� 3"J=n�ɡ�+�"��ǋ���d�dz	�o�cYϋcG�U�w~�m�|V3�Cj�p�?s^�1���﷚��z>j���Z2k��zvz+���8u��g��op�f������nR�� ��ϖ§x�ƥ�?b���s ���C�J~���7�Sf%Vß�K<PPH\�3��<J�{����#��}��r�p�d19�G�b`'��ݍ$�ad�Q�3;����d�7�ۈ:��Z4�z�e�?�?YƏU�a�2�<����t>�Kf�pᙕX:��5�Ŭ�~��(e�_�5sX
���c��wROb+��0c��uV5Sh}l�d�D�e���}k"[�SE�/':�B����5��R[V1�>7�k���%�Õ�>�a�)���#�MUMu��2��`4g1^�V����������{~�`��5��dN7�ߝ� 㢦�o���/y&o��q�̬4$�퓚ĥ�8ĠȆe�)��_V�?G�J���[�:�3'f���E�)*���>*��u��,��cw�5[$�K4|�;�,�� ���->HI�}��� b�L�Е
�Z�߁[���9k"�jcP�X����B�b{�עZ7Z'����%�:�M�QR[�M��g+�\�nUECP.�P��9a>�U�g'�n��.x�\c:�Ѕ����r%FH��P��e����&�P����
_��R2z3���C/���>��ZH^p�,wC=+�w���	�56n��gy%͢<�ӥ���7����"ۍ��t����h_tPa�����рC{bw�6���z3e�5+C�+���ED�lu:��^�t���2�HJ�䯪&L�P�΂�od�9w8�o_����E/{�fRz���01��]UC��$=ࡖ�}v��"���m�����`�@�j#Sr$t8ލ;�i����>�7r�W�5Ǯ���Q�S8p�n3��-k�w))�Ȇ��5��X�rm6hY�/fy�L`+G�"�7�Z��|��fY��سk��/�O��z%w	�� �:������zh[£�ΰ�6�j�0�p��b o������'�F"����ECIy�嵸W�~p�>����]h���I��Le�O{�B��A�!�F��G���������j�(��gt���eO�1(����`�H����;�R����l	��Jy�*j��'���6���T����2��ܜ�
b��8/��߷�����+0 � 0�@�s�%m�]��P�����k@�� r�*1��N�t��$��W&l��%��ĥ�\��Pd�ލ���A���# �w�z��JK������Y���h�T��x�e�Wy`W�-F�Cd�@ks�ed O.������tM�ޕť�!Y��κGl �C���9 ��N����:���z�/�;M9Ը+�W64.�A��2�.!�We�#�zL���A���C��O�I�,�n�Mť�k���X�]��ģ�V��]�r}���YcҚ�*T�ͺn���o��$��T�V.Dp��)%����4�K��#��o����8?6j����1P��|�EH�3J5�t�cm:nGQ@���S�`N�	���V�u9{��+�E�W��I�.����cM�%{_wy��9Z�Ž����ک��>�8_��٨����yPt;Qq%vAL@������o�F��!!�C���a;�ӕ���*Ech_�b�횺X�7�0�+�R����+�����$%��rZj�����geK"�:�����/��������,��F�>�B	KDM�30t�H�1��~�w
L��Gb���f,��P�	��:)#Է��`��j>�neѯ��	䓲��&=Dj�e���[R�-�"����"��zuĮ������2|ʝ~bl�ߴ��A	3D�(�Hx_���[����>��X���N/:h�+,��O��[+͏�[zx+<8@�-g���U�a�A�C��)X��!q��u�qEsz3�.�����S����Z�
%��%�Z<����v�m�$у�����e��QX$џc����<�[ǚM�"|�yW�gj�%+��Sw��^���Ts�pT<jVWܶ�)b��}Y	����4Oe$-p��~�$?��r���%a�=�d���x��)�}��QH����8)���"m��}�+2�r@����bO�ʅ��ͱ���#��M�{:s_3 � ��fid����BȔ���^|T�ȏqj/�SE���xO��Y����[�b^���������ic�������c��u�3���Í�i�l��|��ٹ�k}�X�̢�>��7�"�n�.��7|B�e�1򀅧-,��-���������$lc�!��}��9yA��jɔ�3��i�i�i�!��2��2�Z��1Y	ݯ�?� ��<�Y`����,P���]A��q�8��aw�~����q랼�+�3p��"ZY�:��c��9� 1���7�ifҋݹ	�7?ш�W��#�l��sqW���g��:�~`��U���?e�Bhk��|���GR��_0�l������@3俖\������}�����[��:p'�/�P�;.���嚸'	B�^�A��sl���TNU�G������@�Z�-�n�*0�}k�t=���(j�$:]��<UՅ�
OB�&4ArrF*6f�>#�պN\	�C���r�'a=�~�� s�fU~�h�������^���Z�i�Y㨖Rº,c����Sc�AɅ �d�0m�7�{RyW�����㈼����"۝��Rm�+r	S�Dyn���X�	�7�=���'E˲��(?bn���1�O�c���s��S����B�Hsm
ֲ���`�~�J"�wt��,�f�p�nA!�aK$I��?!�.�581��8��E���G���jH��E�vGZ66��VKY��X�=�	��@�[�a�rHF��i�����)5����L���ݑlQ|M2����Čr�+�)z�)ݜ��~���-��|����WF{�'���i���0	�!t�2>E�
>�K��.��r��U��}c�Eɞ�K�zzJ;ts� ;����5�KB$�ǘc�1��w�#���lp�b��'�/6��>L�]�s�U�r�E���[W	�GJ&]�9�]>��7zu��iF?ubs��:K�ҋȅB��v���/�<>��md���䜁h ��t�v���F귷�Z\��D�j�K�v%~o�1Jg���	����&�f�sL0�+�Ђ�/�[D˛�v��d1ʯUVE���Mf`�j_�nnj�@�K��ѿw/���@M���PI&-n��v��V�@���5�H�T��HY��+Ϸ��L%Ly�~�|��=���$�$��2�V��c&_�q�u��g�`��
��;��4f�$mv�\/@+	�8��̎�J}2�e[ؼ%�xWk��R0���#�R�̭�ʡI�ȁ?������1+���㜄�5r�]>������h~ �ju<+K�?�����]}�װfX���-�l�^�?�姊r����K����~�x��'��s��RC����`*R��8 �!�ӗa�{O��Z��4s
>W%q�l��*q�c��H�6��[������l7G��F@�p����y�D�(Gy^|�1�s�_gӁC.'Wm�������<�5|�gp�?@7�nz����T�w�e�����ξ�!8p
F$�	���E�^�E�_���Ũ���=W7v��*��R�
�ڗˊOQ�OR��[��fT�T'ԑ'��W�>�sLm@�zdS,��)��U������XF`b��<��[t�����wW"3f�Je.���W�g�c1=d>�6��s
�o���^8�ȩr8�{C7�-�h�A<��������>��@5rE�Q_<xt�N�����~ٙ�n�CeS��PL}U�BK�Gz}��+L��q��B~�ұ�*��_���s�R��� ��k���w���ճ&ԠjNW��KLT>�x~4@ȁ�w�
!�כ��b���V�8�a�+l3V"-37��NfG�ّ	��~��)�h�'Jo\6o)�V����1�~
rİ�2 d�'��%1�^�U9����>��x�w0�4�,�(�7򻓖͋;Q�,��?��.A�/}<��J��A�h}A#⭐��%��ڃ����,9�k�4$�+�����8L���E�����J�����9�@G	��sBP���Q��jB��L�L�س���7Bi�7M�F��(�+[�,C��ڹ�81�q1]�ܸ+�1�)"�_�](����#:�О��f�д�vǖ�Vl�#9��o�O3h��I����Q���,B�8� R�������o�!h�;�\�1���0��2��w��7�].�1}������H]zR�U#�!��F��[8�@��{�&;a"��������9����ۗBe~��9L��_����㺩e�1���H]rh#jn��r S���Aک���͊��.��k�@�S-~�猯}����qՖx�8�S���$��X^��G��؃��Z��Z�u�i�P�#*����=�9��Q���̙�;�:�\P�W-�	�CPs_��v�]�{��NtK����6�K�i�:N�.���옕����c9NL��竃�Ǟ�
�E#?4vT��	�E�7��D�P��7�go+$|� ��[A~ht-�㞷���━��?u9;�D>JM�:Q�f�%��h:��Td^ʷ.����1���[��-�i5���&�mx���g�.��]�^zg���������@�v������Qq{��J���gpӗቝ�{�@*n{�T=�39w��^�˨�a���h_�[�T
[���-CD<�!��L����E�B�&���q/"8ag)��g�����H���a/S��E�v_�y��|,{5�� ���ǭR(��7M�{;OP������q�ӂ�,˓��ED�#WP���(�E����`[K�0]}��iT�u��p�w\Z��q~�����v������x��II�!��Epg����*��x��(��y�E�+��� Mcp��	b�Mn���p��@����?_"���e��)�����
���%�uW<أ�:y�E�6[d뙏�z2u��r�^�� ΍�F����-&k�D�t}�Z��og[�?ks�B����G��3D���ܻr'������}�B@��F�Ot=�55�oXs_��Ŭ��L�(Կy,$Ѣj�vdT��.�$fZ0ц�i#
�݋v�P��׋4�ھ4�)\�-C�i��g�5Ǹ��[PMdۣ��ȭ����$��L��_��>�zJ��s49�U|��WD\2j� 9y7��_���I��q;3��AR	Zy�Mfj���X��[��K�t�2����ʖ�J]��ڧ���p;�t�zK�f��ң}�J4M��DE�����9xp����N���0=�|�t���3B4��B���U�k� �̄E�%�Ńg
V��'�L;����hQ0VD׈��hN;��u�__��CeӒ^���z�Ha���F�����f��ϚX��1�6�
¤�����3J�=bG�� J�[�t���1����0��{<�q#���8�o^)m�F�Km�%��9&�/��/�2�ia �\Z�ō������&6��4P~a�.\�NA�K��i��ҩ��G(���{�g�}��)|Ѿ�(�V��k37�S��z62����|�zÈ��a�8s"�j�"�p����\Ԯڸ7�ūX�$'dDhQti�/r���lO���]��|�����[�TZVB�Rg*M������H�T&E�Ã��ُ
�]6���m�qr����Q^Lk�G�B�S�V�9
9v�>`W��f�������XM����5�-U�$��a���,�׎K� /��������6�v�3
�}�3�H��_�B[5����;옃�V�/���K·co����ڵ��]פ�I&d���)y�="AG�a	��hc� "4=з\��O��Mt���61�+])�d�a*C��e����"�>� �%{	��M�rL6QlEX�,���+��J�;B���c�V�K�x\���_%�Ga�q�p($3���)3�5���;ԁ�cj�3�|�ݜ��v��p�4#��J�P3�S��p[?��FV�ꞩ|�FM�r���\*�ul�xō,��IdE����.�����h�,$�$#k{�Nv��̻�:4�!�:Qz�?W�:�Oٔ~��d���$~,`��{��v����D�\nx�z��G$���1���B�ry��ˇYK$cEH�1m��X�Ztd���T���z��5p~]1!����d>qR�[<Z�x�����)���[�C�>��1�H���P��ҹMAuoJ� �*1��dhj�@��������GYO�7���qO�H�O�.͏ڦ4E�Uᯧo�K�#�L�xC?��N�u�<dJ��8�@	M#�A9�C��e!�ޒd�} �u��Yj{m���G~,p�����/G0�VxKW����ud��
�	c+l�u1���^������m��l�(��ټ�Z������%<�U���j�f��/
;��J�����@�wJ5ӻ�_�6��k� n�b�+^`*׫�4�m��!:����}@�_ݵ��)�X���l%��b�R����[��_� �?è)�������T#Dvq�Y��b�f}��2�{��~�
�tƿB2wxVQ�����q����.uRHa50�G�H�xo�lWL���!�l\窗0�����d�6%�tL℉���C��)�H� ��隉�a�D.�Jy=��S�����#<`g����Q�����83�D���	�*F��e�D����+��pڢ�ub���� �Cٙ��W;�(������(Ē����#���^ˇ�X׻�Ք�r5�/��bfd�8���|j&?�H�TH����\�ʸ���(ͮ�!#c���©M������IZ�xF���/��<PXX��0�"��g9H4�j�σ$AKE��8�bu[�y_��uȘZ!�� �G�~��uv�p�����D��=f���G;"L�D�C�eR�#����y�P�5�����W�H��~�=������B	I��cCx�Y������8�W��j�cI���E�*�'�"
�A�f:��.?��-|Ǌ�=R���&pj
�S��d�j1������g���J���X��:E��.<4�=��F�7{v�p�c�!�q���"sE�B�]���k|���8VY��
��NYv�����q��7����w��� !8�~�s�۴��ֹ�uxq�|)���rLO�G[/O����"P+��H����ǀ���,��<�"k���'p�b �1Y�L1l�r�{,w!�|c�V����@sW0W��gW3��4z�C�� ��:[-�0��"kF��+��.N�5j
[�K[�{>S�
����V
H���+Y�Q�<JP�"%����r@:�o��&�&���Μ��e�(�W���&} ��/!׬G�$m���t"h�����\	Q��͍*�s���V����:����ޤ����R��	;�c�W����l�9P ��p>�1�ѿ�w��pV��dU�����:mb�LE��%C�i���9�Gb� ��K��S��g8�A�N�dFG΋jhQ���,&f�R?��3mR7�� 3��R���v�!�Wq��1����sV\�~�g]<0���^w<�:m�V��P���?x�����'%��ճY����#�yJ�`��f���KW�4��æ9s��J�H�',ڴ��tS`����%�M)�RN�$��z�|�6���x��0(�U!71���y��`��`���?w|x-��˗�F���Hk��u��9��%ڦf�{����q����Ó�5\%d�.�I{[��*K��.~L�Y�S��dN�ܭ�VE�o����?��ɾ��H��x�3|����/�K#=	-��(1]��Z����z�2X�-��ϭ�x%�T�q�����# �WMU$�q�=���2~�UZ=w���<�0E�y��ز?-���!zu�N�`���Y�Bѭ9@����F~���,�CZ������Yiw�T�$Q���n���2A���>!<����������j�$�]��u�v[����/������h;Eu`��n+4(/'8�.@ZT�(�V'�o�v�n��j���P!o�Q�&��髇5���3��*W�>���9��L�X`�i��٭)	]��M�ϩ�H&�}�o�Gu��A�#����mƋ'�{��q>S`��7^�Ҕ�<�I1^oyIx�� ���S:֊2��!�y��S7f��f�B���Q@�px[���c{/��̿wO� 0sn����̟!-J��J��_���cW�	�_�^�f�ʶ�A4�9���0�v]���[�⍳>����uT�s�Z���	��4����������J}Ϥ��Os����	ɝWY4�"ۜ-����4���+i2�3��蒝_���f�SJ�?��o`��6}A{RJ�����+�=H-��=��\�>��+i�(w����^2��Q���+i$D^n��2�ƀ���(�A۳���c\�D1_�X<�['X��J��Z� nr��.,�n���K��߼�\ݨQ�+i@k���й�v��S��� .��4u�l��ݒ�ÞY�꿒P��#�+�A�\��f�����x"��<���*)$L��i�UFZ�G��,����O
fc��j��H1�!�nIH�G$���]��TN������Nu �F����>��NA�
"��@'�149_A4�ۣ�}�om��s��(V����Oѫ���ԝ�m4g~a3��u>>�|�#��4Y�>
[�P��\M�L��Z/�6|k��fcpPI}y����z�Pv�!��[�$�����ƨ�<��1��Z��p�?A����Z��TB��Ez"b?��@q
1��Į�ٟn�KY�C0jN֎��RN�����'-8����*�u����Z�b~X�q� �T�v3}���GzX]���Ԛ`Peu��P����j\7�|8p��>��<���w.�e4  �ټ�2������(T�uP���f�}p���V2�d=��#�e���OuN�G��+Bx�?�H���(wC�_({N����ڎn�jڬ>���y�]�,s� A=�^r�g��;��RL�[�G�d-%��5���l����μ�a�+�4�?Lu����Xt�_4��!Yfp�;_d���E��}D�te��H��� ����/?zX!t�C�#Wfs(��u��D�Q�WrS�\aJ�~0b�Iy�#��mא,�4�4܎MF:�pl�oÝ��֬���mu�.�6���*������iɔ̬z��nM,�*j��_�;�Hȩ���)y������b�(���(��9#���M	��0��ȩ,C���kH��,���3���n�~���G����_t��v(�05	q�5#���f��h����9�֣��0�-rm�%�8aࡽ�U��m��D4��<Z��ه�%[Q��&�|�q'5�:�~!/Я%�sŗ1iוֹ@r�ʫ5j]]�n���6{�������L��h�Y�`����"�~�{E���ʟ��m��D�c�怯���|3C����P�m�j1�����i9�Gߕ�|����:�U�-�X�7���6�h����VJ�-A9�~"L�K\�fF����z�~0c�R*9�Ӌ��x�e���_o������Lϲ���%�6ۏcMk:�U�Y�v,친Z/��|�`��y��%'�0v�]�8��v���@U�@�C��,a�]�Zcj���sc�hEц:> �Wg�&�;��CG�n�H��{[�(=����s�n>��2��?���01�U�>\6zeF�����ȑ@K�mF���$�a�[N>^�g�gH�G;��I^�Oy\}�rV�f?M�Ҩ8;�p�"��&��ԅ��߸ս�-�+��\x��͠����pI�@;�:?wM0��}v�ݩ���w7m��w*�f��Eg��|�u�U��T����Ek��4W&�qTr.jf�2N��u^���"�,�)�T�֩�2�[*_�P���lԵv�&�l�,I����z]W>��P.X�g�����Ǹ�S��b��~��
ܯ�����#�y$����;$�{Q.�GJX��v�k3Kt�#��]�9I"U�xh���_�f��F%����A�f���??l����� �y�>�r %��EF0���y {����2�"c�ɢ`@#>�B�a�(����n��R�R�.~�^�úi�=x�,�W�$�j�zwx�#�q�B�_s�d�����_�C�Y�N@�}���o�.8L�:��o_=,�G�e�|<� �X���V����^K& :[��2IΤ|&��$A�T�7_5�Wu8�Yre��W�������\;p���1�c7#�����d`i-S�N�X��P{��~�?��t����o��8Q�/Gc��i:��ɏ?��,��?u�(�<
�"{�O��J��ǩI�:�
ŏ9<3AE7�.T��ػ��Y[RǾI�N���ĉgࢹcz�拶M�	�%���\0�|��@�)x��{L"�\5>z�Y��B�_2.�0OcĔ{٨/��(�U��XF��`��A-�B��h�Ӛ�ۮu�/���i$<��$8��kj��2��H�������0#��K"�����e�W�'���Y���Xg��1��ٕ���,�t-V07묰����J'��-7��4hd�����k�Q��+�J�|���Ob�[n��/��^>	�
1yW31������S*@�$L���szF$��0�J���(4��3R%��ܸ�\�݈`P��M^ðbY��e8��h�>���'��H�����0	������S��h�m짉Q�ȼIT�H�����?!�d��i���vFQ��3���Q,�-j��Y�,�*ň_���bD2:��]�}��N�+'R�q�b��}>p��..�C��^֡%8"���joW��yQ񟻁f?�n�cBI�/K����eP�ځ��{�m��;���$q<vʇ���=�1�n?��q�gm�Z;C��D��{L��Q�*��>�T���^9�%��bҵTYc�h�\.��"�܆��1^X;/�A�D\�y��T�F��r/<��;h�)֚�}1%���J�a��@@�ʑ��b�9��H����u�떄�e�F,��5��7a��)�K�FC��w���sp*�oDx�ߺ�ׯ��X����1�mV`$��N�@p𖭿�;�W�+�Z3#�#�"�N�9t@R?��P�q�l-�
��a�	�>n(m�_�с-�����h� ���-mv�fb�F�uG<;��-64(6�y�sC���xDU��]��E���)0Blc0M6^ѳ��9_�%��Ҧ�þ���=P�?e��9����O.vF�{fˑ�0�je�c���@FO���)E���N���9(-8J�����U�cJA�A��JX$�Kev4!R*��4��ji9�E�/�&L�i}cA*�:a��F�Z> ��k�\L�~�iL ��Cgjq̠�PW�U?4����m �w��rW�ƹ�K#o�F�d�?z[B�(I�5b#�ž��2�Ca��5@I��b������/�?�92�A������Lе����))�q��=���k��**�2Ye}o�h��{�ƈ�nn���rӣ�����hOo��!A�,�Q$��i�<�؏8�g�{�������H^��o�n���^'���4�ӱ�$���#�C�֑K��U�����ٴ2�ށe��4P8�0��j�e��-$�������w은��o;��N��?i��I�mt}��:�7�|f�-y�n{9c���<]�r�[�Pm?ݎ����Ռ�t9r��.�
�u��J�{�aPuHD�K�}��O[
}:8��ޗ$9>ǣ���,���j�h�zM*Y�3\�Jk\ѱ#���*�iDf�<���\�B�9��̩�!�!���_$�,���[ 3/zܗk��] z�e8}AX�؋��7���88-� j��N��--AC�H�O����hT��d��t��?�h�-Z�7���m�����-�g�h�aO��Wc��u��ީO2M��Ԅ�2����
`�Q��G��z�%q�^���}:�[���d�R�lI��2�4n�)���ғ�������Pk2S_}	u�oTsA@I�o�\v�Gk��	K���ȕSW���*�KO�F���xN�����a��`M��8]f�$u��΋.�G�;���2ޟ�N�_,�p]��O)߻5�uV|��~�Bl���<7�s*���� W�Y�������,��^,;��;c�����y`$�P�/�6�dc�!����O�� �c�,��/��yk�%[�P�
�iZ��mM��K?���z���i�;Aw����������e�{/7șv�g�{ڡ��2T������
3j��XZ�O��t��5F��Ͷ�{g�s�%&�����R�'�����ra��P���U�rl��2�V��k���ms�3��G��b�Bz�7>�J��O�7G��mHo��^i��	4(���eM��0(��(�FE%��+�Y�x�h&h���I���E�|SI����D�Hw��>�#?*����ښ�;�j�-�pM|wg�����u�x��>^��ug���!<ۙGq��<�XO�&�~A�F�^���b���zkt�A<���!������ev�{�ƒ���?(n�Y�yrc�z���4����O9ԣ/���qڌ�<��E�f/��C�D: �ߕ��0�;c�j��"	~v��39mX�$1@�/����F�/׶�uK d����� D�.;S��S��)Q~�����0J����]�~����a"P}�m��;'C1Hl�.�]@���&x�)��U�틤�/���>h<�g��71��q{EM� �Q����㫁b��<;$%W��L8>_������%/�#ŭQ��F�-ʮho5���}�?3�3\b�)�s4<Z^���d���sǔ[hp�2�O����iY��G6 ���yVU-��� ?qV��sB����i���j�<�ג�m�vO7�Ҽ�pơU`���Ȑ�Q*	�3���I��ԉ�h#6��20��@�E��bD@-��<k@^��>��������c����F��5O#}m��!���ܢ��՘J�]���SW���LDیW�a���!a�@Rm��O����B�}�	��v'aT䕑"��|�K�f�d�c��O.o.Y�$�?FՖ�-Wm�<:v��.�&#a�\�Od��S�-����%�]�ו��>�b�����w�7�]=b�U)�Q��i�g�g�{/ƴl�R�gJ��L$�Tg�f�ץ��
�1��V;'Hv�ܸ���=�س�MJp�h��+���C�oj[mL�M(h+��E&i"KV��4!C���D�[P鶌;!��8�l��@ Đ��!����{�"�"aV�J)3Zy����!���T-q�y)�,�y��S-� Š�Ӕ ?>��K�FD���0�*�F�y�X�Au*��X��5+b=fu䬴�߽<OȘ䱿p9��Ù�r�����|�J�4��6]��Z�b�i����Epm�$I��;��:�P�u�
-T,cn���\BA����� w�� -�Q�¡~���A~ٺ�"��#�j�>z����xXj��B���J��dgR�� ��!�9�T^��g.9*LMt`4�}>�Y���
�%cq!�Jإ�*�-u�����8���ˢ$�����	 ��	MccD����5;ω~#�j�� ���rL L���޿�|\3���T��_ӡ��h�soyi�X9Ȫ�	F�Nh7��=�=��8R}�4Q��Z�a��%-��TT�~��I;�P�ĕފγv�??�jSb�=�c!c����Z��W�~���������G�쭹Yu��S�t�	��w��yO�e�X���������lS�_K�n�Se�����lw�h�]��^~���9���^4�8#^�{��Lv���WɅ_��#�Xlބ��T�y��AtU��>��ze �p�_>ղ�o��q�8]+tU�#B=O9�ۜ};p����x��V$A �:}��?K[904��j4%����_P�2��@�_���1�qI���!�%�=��ê.f�I����#�Jva�$�{-�-�-jȅ���>�=�J3�q�܈-X$��>���wF��������F|���y`/������޾t�b��!����(�A�DU�J�:0��_������r�\)D`fv)�7��Ũ�_o�)���u�{a��ziO�ϧ����z�Ola��%�_q���� �y�b�LD5�$En���zk�Tޖ~Z�w��=E�x�e��/R��I����H�&!s�q�5y�Sߵ��ۺ&{��1LU󀔆_c��k��g���Nq��M��(le���W�,W��5Q���8��L�b�������t�MT�6��
EM�W�`o>(%-�K�������}M�ny��/��ǡ�d�����	^��kF�)X76���uY>`w��䂋�H�t�?��ѯ"��#�E��(�XC�(�z���T��ǟ�f?��v��%�y��OU�=?�kH�Sb����G�0�����|�S�
(q��ڷ7����\[M$pJyҮ�WH3��al@�5R��Kn��2���KR�
���5��ź;j�`Q��ZcK`��<�2����,�f��Z)�'��+,zÊ��j�zX��-H@)��M������2\U�A���M �H:lck��F�ӓL��=�<R��ܾ��7�_��"]��U�F g�#���훂����������:}P��7�h���
X�x�`X��b�W���/�JE�̱c����#�F�N��=�L����o�� f2���J�U��:;zP	�`���r��)s��/� Z9�Y��Q�:��3�����\��O�j|b��t���HI�V]`��D�?���VY�5�y�M�{�P~֝���3�x�P�� ����Ti*g�$[(��/��$�}�/�5y �<�'d;tl8�f�I���Ld�)a��R�����E^�צ�x���5�����&��|rO�N��P@�� �|�<��r��.�Lh���b2��`��Qo��H���Z+�E1]�n��&����R&��"õ�����E�'�c����
*f�䇿��3:꓉�E,	��8v���7����c�!���6�|5��?���y�u!�ї���2b���d�f��I~����𺦢�����K�rC�\�������B��!5�� �A��La@M�zW_>��.�Ʃ�WQ}��K��tKK�͙M	|5|,�#�Z���G eĞޟ�A$��/�{/"����oP��"���+��KA����V��./���I;�c|m/�Q̤��M���<.���Q��9��C��&/ϒ�K��+;����>�Kd��1� ,D!>m���F��O�������w���Z��Qć�X*������A�Rh�<7�}��c���Z���(l�Xz�/8���f�B@c^/��Y(odJ?�=9i��@ǣ��/H����	ja,�5lA���b8���0j��Ht�B�N�r��m��r
˄ �bF
3WKE>�~�t�"mcKJjT�˗��弮FF���fv՗%��� ���s8q9�8�?�u�<)�Q���9��-�m�M�5��E�Ľy|c�NC1IwX������p���̚]��5�w�×P$f�����M~������:��h�&����3�t\zEJ;�u��v�A�֔۠ퟭ�Rk��>��k��?����?�
O�1O����
����ߴ�p���qv~uy�#��S�*@�c����F���.��%�_�/~�tr�@Ik��B���7�M�\<6
1���>!�,䘶�!H��Χyؘ���̱��I�X�(��EWS���Y,�0��߶��=t�7Y�t��d���6����^���Q�j�O��o��I6د}����%�R����[@�@௴B�P|����fM�O���WLi�����spC Ϻ'�a�p]ǚ=���*��y' r�h�7c�H����	�]/z�{"��~�~���#�����2��2k�sߡ��*F*iV�& ����k�w�&�`���o2P�Nyx�Mݎ��;����/i�q�YE����fX���5\ͺaq�x�Ėo���1fu�'�5 ز������>[Aq�|�,\!ը��H�v7$����rԣG�p�mN���*Qe.d��c�%^W�kY!$؍�"ZVO�� /�V�6�Z�QL��c��CJ�b����x��xN|�6b�r��w֮k�Cz��i�>D<��I��u�a3�)ఄ���9eP�8?9:��q������ޠ릆�4:��Q����M�5��9>j�S�#Hv �����Џ�"�}2�r���1�����A�Gw95BoA3���G��Ө0��T��1<�2H��K�3�Tڃ������!���K?�^�\��{y=?���Wm"pU��޽� u����kR�{sl�b�,4O�J�T�|T�b4¹�Ke�N���?�!(h��N6g�Se�O�(K��:_n�R���p؃nF!E;��\�6F܂�J��(�	�l��,(H!��6�Hm)�d�_�+�Vb	���g����>I��H��6M)��\es��#V����s�T(�F[e��K>����i��k䮇OX�N[��D���p�oS�1W��2�BS��c	j%�ˆ~���4�Re�z׌�JD3�^����]7�F�JX>aFg��m����#����^Y��
r���t��`2R�qVQ��
l\L�?���{�_�Gƀ�Öp2��r�zO��Q����2
d(��N���o���S+���%�?�#,�9�]�����^/ns���:�#�[QQ
�?=!M�k��FI ������&�|W[P7���}�
�v�l�G�U#���!+q31�7\�]=ЮxH���;��Q[�G$O�v>�2j�DR���%����X���Z*�e,T���u����[�q�?�N�T6N�3m�i������/��_h0�@��I���/C
s����"�{Q�8�q4!ks3��LЪc�1�7�� �y�����P��dJ�.8�dpy���k�����+��>n�Jo�|I�j��J峓�@�K~���A�y�D c! �mdҼ��pNI[2U��	��a)�ƣ�,2{�N�F�Ւ�QO��C&�g9E�Њmh�/�0E
��&��SĖ����t��6�,0�+�Æ/,��� G�$�vz=���>I�4�?�TSR+���p�f9����&�M���8�.mO�� }�����u�_J��b��Z�7���W��6i�.�#�L<F[к�x�����`q��4��ԡ�J��w�ζNh�t�	ά�C���,_��?�g}6�wdJdɯ��hK�W�_���ϊPl�,�y�����g݉�%v�M'�dk�-u!����s/��J�t 5�Y����w"�p�v��"1;�ȭ�.��M�$5��7o[����b�~��޵�xB��]���z@���u�K��T�Թ���Ǧ��}�l�[D�q��0(��w��9�EI{`���-r��nb��(�e@&�S��Q��\�%@���� &���p��g��;ۯ?J؞�}���c�J&�r�99 BUJ��I�.�E]�ॊ�S�7w ��?Oa�٬4�:2�-�)}�!GF"�s����f�B�����:(;���a�1���*��+���E'ᛕ�R<�ū��$�(F
�����m낰VE�t��C4���ě�Y��Pl�RG��W�b0ES�vW�]R߼��Mc�}	�v�h��U�>���fZNZ�H<W���j�������?ۄ�ه��|S����%��턾�sQ�V�VbB51��L�mɼ ���|!C��Ý����7x���NI�9��(t掋�W�����i�<�
�HГ 7D��ξ�>
�p��bZJ����n��Y5��Q��B�c��I�u5��o�ZP�+��$bՅ#"��J��d8�`
�M���!�u��B�2��fzu���7�s`<�5⻑v뿥�^+�ݣ��7�WqR��#�J���2W���CƮ`x�)�ڲ��ܘ�����/e;��k��x`Zv��CԧfUs57�%�,f���I�<�G�����x"t=���0�8�r�_����#��fpE�0Ţ(x1z���M�v�)�>�����ըu��5���#k��Ά�&a��Xq$�
l!#�6Ea-?�\���;Wg�	 ��P�oOiĳ��{�^��s�ɐ���L9L���Fqy�z"@̣��B�C�)_6��ǭ�'_`���F8�u6BPZ^��ac�����<��ox�Vu���QZ�TZ��g-Q�7�Y�A�fa'VZ�	R�N�h2W���'?��Z�B�K/ ���q��RTP�d6��m��GHᢈD���T��rǯ�c�����ۧ~)h�2�n��9���*��:�����3T��!z׽{N^���Q�w�}�5�����d]x�P�_)��,�p�h�4R��G�V1Ë1���N��Fp��n�+�頲��2��+�3}��X�L`$f�2�%5��9��8����n�y���jAA���50J��=Ś��X��9�?B��� 汅�'ǒ��1�V�b#����Q�F-�.��KOn�:����1w��G-�r��߆>8��*�'ޝn�������y�a4����0 u�X�_/��|$M��e��~$�4�t�AU�]U�2�Ɓd��p��kԏ���j;N�J�� �$
٧A���4.��8�y%�S�{;�x�H8#�v?>�&t��Л�`@1���X��O-o��������ĻNg>Zz�Z���;% ��_؋��
�eG/��\8�y>����m~&�[�02~�)��?묞�;����u
����R������xr�F��b9RjV��R�*%	��߿l��-z+>�����C��Oa�e9��v1풪-u�*r�9�ԥ�3:y�,�Ӧ�
������T�O<v�o���=�N����4�{G�b�I�ғ���F_����Q�)!�-���8��:�[cƤ����PtUi0F���Zҵlx��9Ī�N9���]�_�$a}�-�J@C}dU�k�Z�_E�Fv��R�e|h�L�a�Q��@��q&��G)c�P���'�n�8	�b��pbU�P@�c�$�����?k7	γM�� �'1l��l�V�Mğ�ں=NM]���`+��9�ޚH/���r1�T�_�u��J��/M�;7iI�t�˘��ug�Q��� ��e�D��U����UD�A��f��b��%!�?eARl�yp�v�!�%�BL5rej�*p�єB|��cήSe"wk6�K�z��i��r��;��8��	l%9�8N�j�{�������ʞ5���IY��)h]_1�D�Y[6�o���$��./{vu�P��&���㳱������AQ1c5y�+�jvcsĻc ��a�X8�<LәT��s"�����$�lH���=�����&�cӯ6>��?}rZ<�H�k�-��ճz����4L����!��Qo��s ��kvD���wl�c�U��<�"�yN�ъ���xv�o嘑/.��<�́�EV9~Iô�S.X����$xi� ���a͠�C\ذ�m��q9��[��R22�	4��r>w�e4���+�թj#��6�#޽5?�a��_cw���V,E�>8�ǐa���EV����:o�(�ۚ�xa���{8Јm*��?� ��d���]�|P����#��
�\�'��:p0t)�/�x���<=��<��;4v^b��B+	��I�͘utFP
�A5�-��S������Y�e�N�ǣ"�S~�2"Z�1�F��Y�-���j_���\��Hb��%,��k��V�=齞Ν@#��ϡ*���b���|_8��Ԟ-�M��_�:Ыꋁu&AG����n�#�V@��n��X�t7�Ϫ�5�5ȓ1bWv��n�ɤ�wr�Ek$��_S�p��f���ё�K��v.k�9A��rdU�MA_�z4}b��NA��nC�i#��eÝi�m5;�JGLc���@K���1��_��},u��چ~��<mW��+0�̌´�eRf��S�E���%+q�$������~@�k�W!�G��YJ�n��v�N$�8B��+���yn=aT)��Y��"��h��z�����D��$���re��d���ǏU�ͪ�0]a���賁3<���)�~/�9�g\J+��4�j��w�!������-�{铅-�^ dA�����Jո�(ۼ�d�>�ڬr�l��4�� �r[/+�|�
*j�45n� �J?�u,[k��4�����ݝ�O�RR��n��!T-r0��k=�>��T�1��c͵@�#��#������!J^^7��H!��>ء��ؐ���~���!�T�1���F��'����;���C�Heo9���C����-��h�$A���E9�-� R�SSKA8H��r��%;Co�Q%���9���3^v[Z-O_Zrz7������p�Q3֣v 0��8������w��2�^�/���Kȉ����큎���?�5
eC��}C�Q��m��ٸ�����Ԇt��)�y� �߇4��Ը�Je�w4��f
	�΁ͣq���j��K#�_I��u8��-��������Տֻ���~�-ˏ�*�ėJ����;qS/oT'�fbH�s�<zD ͥ#�!��z^�ɑ��]��m��0uE�,�>����o�y���x1S�[�bHM�0s}:O�}'	��H6<g��N"�m�[��qaY�r텎Ǥ�ɒ������f^1���QKw�>�&�04[�W�M�o��+6�l�໮�Ρ��k�̤�u����"��9kf����a���6*I?��C�dI�D��6e."�3�Z)B�i,�Zd1���������5e�x�!�¤�_9�+��D�rDz�Ovd�3͂�*<:��p�K-��r,Ϳ�!���_,|�-��KZy�?��7E	Mr,�be��+l#>k���5��hY�V`*w�z��@V.z���kM�K7�_|Њgw3����(���9�(Ͼ��ti��C#!sc�b
LR�boH�o�y,5�O��Oc�}b�w�$J�	���������#�@w\�%>u�_�*˧������xCӌw�u/P�MrK�U�����I��#�4�������YG5m�n���=��i��>���FIY`$.�c���:Z~C/�e(;����*t�ӭVq�9��ߛ���YZ/� B�H�p�T��	$�?{��c�c<ͲIj�7`_Χ/��t�����3�C��vŇ(h���	�L��(7���I������?:@7A�����X�Î�FT��m�X��^zful��(�+'�/���`z��d��L�@���C�ޔǛ	_k�s��!�-3 �J�,eY�*E=�-��Z��#n��A�a ���S�"��P������a��)�?�	7C(���:�wZ�<bś�:
�䫥��vՋ��S��(�z}[e�ře�^��D˲��o)!DYse��v�>�*�(���b�z��*H"/u�][���/N ��d��{
޾�Ö΋9�닥�S7���,�c?�ʋh���[�D8��h�O|�ӱ7�r�
09@�+0>#�7�H��G�N��ʺ�V\�]��A�H�1�G>�.�2�Gan�p�bV�t/ٌ��)6A����T�{<Ӭsdt�+]���a;h{����Q��QGҠѲM�z��@/�#��.<+W��ԃۗ���8D���G9[��c̯^xaN,G����vT^�ZCBkAӞ,��:	�Ez��dS �����TO���Q�G�]Zq��ɌE�a��r�nx�p��?kMD6��9�_ +�	��5D���D�X�	���'[>:Zm�~�aq�S����#���sX��"j	d[>��sm]a��ѧ�b�R*�'�L�5W��+��tR�g�tBF,?Q�z��#��'��]�DTMd������%�]ױ��	G�~I�t{��k��jѱ�$�J]��˾{���a(2Ĥ�iyI E������3�~6o�q���9���,�}or5G:�t��sd�iN���|�i ����[�`�~�V�Ʀ�4>�Ɓ��R��@��W���$��QZ�}���G���K��-(�wl�[�b�,nP�����<�[s��%��oe��Äi�""u�
4�{T˼M���#�}�$�����|tn1�6���7��Ix�} q"���+Y<޼;�V�S�������"������K��b��Q�F�r�Dz��U�� F$�@�uw:8��>��W��g���<�9�Rؑ��W���-�'�[?y�Z�p8��O�W%#���tfCB#�w���0�n���>���[=N.�����c�S7Q�V&,(#����PB��G��!��y�Dq~?�s���U���K�!I�!.��t�󼉋��Z2~��� ��u�١E24����K�`�!�'�i�X޽ӼeA"����g�#'�f%k��\u�[h���wSN�O�#ִ	]X:�)~����a *,����Z{��������p*A�_�)v��/��1���|o� ,�n��:W���x3S��2��������p�"�Py�\k��@�@�U�?�l�o~�/���I�3�k�$�@+ws����g�j�f![>BGo0�O��`.� O�ȳd1>������8P^��w�VK�ַ'�E��jO�H<�L0*��ɜ�J��7���Lg��]ޣ9.��z��Hi�x�A���Mv���I��}��v���m����t!KT���&a;1,RTr��+u�V����Ӵ��8���z��2!d�[>����UUƆ�[��%O���/=�B,��4�>C	�D�����_j��vh%�E�B�>�v0��M�o��f7�CD���;δJ��ks@؅�j-C�-`�t�Q�Rk����O.'Nk��F��Zi�����'cOKEs�h6�vU��4����%gb$I!Ä�3 V��q��J��� �*����l�B�S��o�� z�Ӱ?{A��vB���0Dԗ�nu5�}�O�I}�@oK��C ���fS�/Z�	n��&;\�r�4�9��(b�v�ݚ���x֬� L
/j	���B�ZJ���bס���)�TZF�ZMD�T�ص_��]b�	�UwJ���T�<�~�BG^.��{zmU/�H۽��h;�����w�J��I0I5"��Ұ~��7~ ۋ����a�ݫk�D�K�W�V���n��AW�݅����ʊ	m��	:�$yk�o���"o)�E�P�������������:���߱�I���u�-���튡�p-V��Hn�A��{�A"��F�i0��v�Ӱ��~J�Տ#�`1�l�`����;ɘa�qtĠڹx�}B ��h��w��H����kdQܸMw�n�Azy���T叨ъ�O�)
�0��>��B�-�2�����f|���,�x�s(�����WV��Y�e�cU2�F�Q^�1x�̟D�*h��˯Ԭ��P>ܼ��Yj�߉}׎TB�#���g7QD�[)�f�BMf�(���B�� �#Öjd<TxBO~��?�O��t�JZ���r	B7�B��iV����)��.�l�+x�����(��-���1���-p0�.�\Yӱ�l�
s8����ˁ崔�����y����6��-.뀃S���~��l:F<[Dў��p�	3D�һ�%=��˴��Zn7� ����&'�W���+�?ޱ�$�[�3�����h�y�8�]�gwЌ��K��s��L~t�%�.~�m�����ŷ?���Y����DK8-�����
/����s;<̉2G	�\�j�SV��27o�E!���3 \?��,�����J�m8�cim[��]3�Ag�dt�UR�SdXRc��CN:BvX��g�C�u�*χ7`O�;Y����&9��ᬌH��$��Oׯ}��:�*+K�:�C��)k{�U6�J��bf��!�):F3�W�������r�nޙǝ>�'�#�tr��?<��w%m_ڤݶ0;GNg� ��f�hK�f��a���yb���,O{��A�P]��w���L��}8�b����A�e�s<�����ӝQ�Q.x�;��"_�d�OSj�}w�ZKrN]Y�!�$�5�o1y�c����B�{X_��D��F�L[��t�0�<�JI�#AFH�P��)D�XS�F��+�d�;lm�O���t9�����2�5��yQ�w����w����|�>+�x�/d�'�,Ugu�+%#��@�����sDE��T��z��f��˷9�,yp>�	D0чҽ��f�CL�Wh����RPNM�T��L�\�/�5:sIh���?������*�`4���N��z�Ta/q���Pq�G0K
��1�������5�����n�m�� ���&n6����7�l4��"�:m��A2mT��G�N(��}�1�&�Ҏ�9w�|��%�G��D�|�^�q�-ίIN:V	�X�N#���T��`�N�r�i���׀@1
Z"��Î&�k�Bb�cx�r$�q�y�d�VKGKK�0�����=Ju���ns�m���~؉�|��K�>��|�����] 7�s
��I�/��P�%D��5
�v �)f�w�Ӗ��i�:"S��@�N�\���$��[|MUE'xj��T�C�����N�w�U9�6�!���{�t�t�A0���W��6V�H��xL��)��XX��z�	utjo�v��H��h�_A��Ȫ�G*/�O��ܾ��Ts�����|�Ar