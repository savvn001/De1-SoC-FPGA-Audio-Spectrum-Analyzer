-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
OYP/eZjl7hvx2RUFT3kbgmBdevomvgymMD9XRPXPKw0wHKlDzSvw1C/HwPHl0BkYLZZT6AH8rxN2
ks6WDMoYX+m/0QtSXpBq/6wqSpc+P4Mv23EbxkUTLjZSaqugN2gnHd6cKOhAMCrO+NWDRAlgi6Z3
h1hT1ifX9j3a81tQHClt0F9JBlC5QFlq1vAPeA3D0g3UO+Gubi/uG7uVCReHOVBa0mfCDRlVm9+e
4pxjY31cuPVxdpe1hQnfrciB454NgbxcWckjVjxf+Rpfm+kk8SEyZ8z6cE+OSz3bRLNpXmQl1Wp8
e0urGexBi9k2jQ0JzPfcjeeOLZnXMGQqVXNmcw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
4YYjO5uC8oy5NOm3ycCe9yfnuB7kdf8gi09mwqq8f7qH+EJXS8pvu17Gw5sVdqn/3YMHrRG+1AoK
gfrJcKeFTNCX6L5RRNIG4jTY2ZVUg7vUJt3EBYmf5+ltGKOCP7xy/6rkoznbyaOKbswsGDSgyBs2
pZ3WJSsmlDFGIP5aqpM6tFqZUQeKI0//AMSkP44zXw5+C1Gk7hpQ/JcgCKGAIaUE/khDtNVbZgto
/o4w03lrGwWlFUIBPUNV1Xw8fxrvHYtfEJxxs6iE5d7bWrmn1oQDkX24RY8a8bJD08iDtshcBv7N
BoguYeYQQo5LcMPi5a9jrS3L38pFt0DwSVMmSWmwGLEEh2Xfffvy/8AgJmpfZZvPOCwzpXNcedtp
ZLMnVeFSwe7vxZ7pZRr65KLYy67htw21rSanTWZO8A2gpefqw6r5eWcXjdVWiCOvdUeJMAbH4qlX
3Hvwetd1u+hbTAMN1ysyS+NKbOxY7NyjbGVW9kbnLKLucLdHABG+5be7CFwqeLIxM+9Kv/zMdJ52
Tx898Zsa7wFzESDd+sVneHNxEZNoq4pZfkNAmCJGUY3J4qrU+d/dwLJd5n765p6xK5ajMZox9+JM
qrx1X+LAMNDwoFSCS3nkfh1Y4uehzOHa7YAZ3+xxc5BFOVF7cEWdsy5nFYVDc67wqVC5xIUjFtld
0wqdlnqPuwCVuOQ7JrOiVaFEklu5lci+r5LBZj/5SxOEHvzUZELnuwrHgbpib2XGlXm8AauuSjno
ImVtEl8+afzu1p3Vi5VEOncQtb6i8ndWyVyYRBFnl/nxOSRkHTVFpxR8ed5CBxo/VvnDnZOEctr/
GiT0EFlfNM2Xm5Ip1hB2OVWtYFsuZpTtzANXCrmtgNy5htGdvjtBcxiRkAjgrX1WqofSZ3kfnW87
6RuuoR7dHVjGeMg17zs7y4V1IinRqy/IXOf1yl9gxv4t8AvCGJDdFtB8l3RYPHHC9/ocybfSUgk1
IWo51/yU3v9HtcqK+kqKfE+XcjEpASCsMGXoogZC40E7DrkUzpPN7HCrmnOyyXrM70638B7HCj81
NIScsqJ/F1PwXggVg/cfBtuiLmOG17Y8SGSXODcFEYKTlmxHNpq9CgDCxt9soODNMdcOYDmME65U
PmqqAEfbSQU6vrWArkwuUV3qB7/0LikPJY3GzuIqlw+RtGRjkwEbak8Jin6SHmeZouTAxqwkKs4d
8Rx6XHWunPNnv0RyVSayQFg8eJtmiPkyhFmfSCxQ1hEF0kEIsyChPUP8hcZYvQtACLpbv/xKbo3O
bgd9G07IZ/ZmgI/z8PNTpvz38NzHkHZba2WX3MUKv+Hfp4JCsoA5htyQJDvjixx+2/zcou+KkzZb
ZoQAboENOeLlMPOZB18TUIdjNmF3CSUcbocqStpTaF79HDtTmrCDWdTTRXYfvjBIGx+pLYMKfqoz
nyP4wAbjDJ13sGT/pEoNSeWQ10hO7BoB2OVrsG/JmQGqHKAWVupQYPcLioX7ixLww92s6Q+g1izP
1Uy1gRq7ekQsXnUvsmFvAOawMHtvJ98T/XHh1GWeV2aWMOws/aiZn9bx0EufYqkWCrX0sqWqRwUW
eT/gjkfck+XnVhiB2z8APaBW7Zio3T+s1X59kMMFs4CJz1M4sEHT3lVV+4foCt9jPalLK8n/V/ql
+jZ/l5+w7doMoZoUFq0Ds4N96muQ7tAgBe3aCk2VFnIOzuB2qeSX1yh/+8C7oDni/DSFdrZG48kQ
KY3A2yCHMujK/jv5C11gp86IAyWikjhAZAVHdCaUhLteNBsYl/klFeqdoOFQp0rDmoMy7Gw2qk6/
j440ApLw2c41P7DxRurfEvfVkA5RG5LXJfKZj7oVXh/SaqyrxkvW2QKRFD/9wzEk9X5Jal9XSIYS
4ylgD8aGsRBeOB8Jq1aNIqclfPgqYF/hlw8NtIvnMBCH2M9LPzn5p5XlUIXStFMGM2jxN4W1bixL
x+82tmQ4GhGRsUnyHlzZGLKfLenYJnIfBMd66itwAKhWuZ2bLoDw7vvd0jhxIyEo4dNAteQLu+8i
HWDKocW9tQ3xmShu94P9xkmrSOvN4I3vXc75CbOVqF4wixPPOklHfwxTHKOAhrLJxj8w8Id11wj0
xcZr/qvABLbwdqgEEOzi2DDpNPxU9Rn2VJpyeG5dzOsElf92xiTb9mlWotDlu0KX8y0rnoa9Rdnu
o7FFbE175rnANiyglUATaueFY7S8US9Iykd3g6RkK8vENIJtq9ENU+mwKKkY+ZsoWY8WMtfkuT1Q
6JjjI3VM+PAJJdx4wdhra/ALOTm28d6A+WnsdZ0t6UUo8cxzUWx6N/b9q01bjfI7fWN0FS/PKVuA
CXXxQvLp7iOrSq/cnuETeILCiX7bHeBdDuMenlg+TfhhKU4K1IditB/PaNhq1guWDiAejDlPcSNP
3ARq9lLURiMUzmRF4/Car4mJgU7aB8fAs71baNoJ9H1TSEcQT+v77u0NMkn58j/OYVrQnQBvXTgd
DBn0W4ZLdM1xvwJ4Qrzb2t38k2548YnDEjF/KI927X5mlWm77OYAnzfXAEk7GSuueLF/GqsRy2HX
GDzSnWh7uLqhmpPcmKrL/s41SXwL47M4hwlwr6Eay66KJ0XDcdabUMFXdk+MWhnKWnUD/HxJUjsH
tJvjUFyEDFZimDhESeQ7FzaN32FfESQU4AiEPoyxQ5ZneghuK0sbFkkoB1du1oXzBR+HGfvztj46
//HiJw36p1fn1Mqtyf7GeppM+igzmOk1UHs0O4ugdQ+DEbdLSm6hmBCDGBFNVUudigoxZQkk9IRW
OkUDcOxqd7p7YyKi3VU2D7xaVK3qleKe8l6b8HuXihtxOsQSRK6tsjz9pssVH+CQoaoqDJCVWUB8
1hGLxHr6T60/nPty6egfmAo/OFk8rcLBB8aCA5bQ3qyzooYNlYMASlbSAaiXy4ZzskRgFNeQprp1
M1zIDhd8KWI4qpSnj7bQahUWE3SklnxDyohEBqkLiLgcCZUeIrh21fgJJnk6CXTa0jqa09s4fvJE
Z8/G1hjIU78/sGkhtrOQkhM6DJfY8v1T16bytY2HUynniQCBVGc3Wmo4Ate/V+R0xA5HqahA1kQ3
uhdQCO5M+eTgkid6nH/d14Y04xEW6FsVxVmmLUy2Cky4hUMHfRO7/Yl0iqMuX+xA09OqBYQtALqR
DU9783QZ/c/jEFraICSdWUWaDJhB/Nh0VzpDQ0pyE3YldRX5+SknDcvs08RaKwGqYQFA+prh5I6/
nsPBOilt77oiGjFBNtEBpC/xJER1BRgqrLE1vIzgDVzQ90CVU7vKCfCvKOhXzGR7ztZBygGBjaVl
iFFF4wIBUSdWLY1WGxtXI1H0ofZuD/CC3xnIXtJi0CLqLo3+qIrYs5dpqEl0ZMB7ywn8a51+pLlD
wQIrW5T4kby9cAg0HNNDdoQIwoNeRGAFHRWx4M0Y6DMA7qVsAiZg9++wqADwavLLam5agXY6oaHz
qW6qybf57n+aFWi3nzv54fXbdGHf7BScJhCfNs0D+EqA9TnGNKhq51Sp7yYov09oMWW/rf+gHORy
zOcqW8LjHuPDYFxmbOR/tEAkkLwFyFs39O8TCt2TV7XnnZ3ZxWvp3nl66LTgaQOQ/PYDoKJp+7mN
lwBkIWMD7fvX7BrkusTwR9b8jX5uJ64p9bLcXDi00XVnSzefQm8oNikKCjlaCk0LN0BDD2eswvdr
P3b9TUfDRV8RH9Cc7r+hpS5uzBcoXCkuZuyGpoj6+qdViewZr2xmc5R5yCQGG2D0bCPR5ovy+D5I
bvaUwJBZXZlsooRQHSdKLpMWcoDNSP0/LYTg+GFVcSYWg3sMfn8rkTw8Mnr2cIcIk/k2t2N61jDE
NaOgnKw+rekIjcMWofLeCv/kQdHsZmpFr0caI+GPowQx4w8BYW2vOcPDnE72u4TRiK7C6iEJP80a
59kJLV+C5j3lSXHNY3DBUuD/pD3JEF/k0VFh+5vUsNLHOe6zS2C1ilhvIBAC4qUq86t/QXat/a1I
heACmo2gLhLPgbBtG4NgV21vDllqhVK0IYmReBZV5AknUjGQJemUhBOtQAuRziGLzrHKXmsDZSOh
BaKcydRdswIHziOF9Sxz1skyW6UgteyhSqATtFFepRJNgIIrCEQ9OghBm0XBBMzJR297iY96XqU2
nUfzvvY1TqDI5t13g2eVGrrWq78+sc3oO9zgBKsTTRGM//bOldTUqAmpnvK9nnTCUGaAQ/C7/RsK
YZzwzjxAv0O2LbME+Zq17Qxwi0F1Yr7wMVo+QkYjVZ7E8V2v3+6YW+6eDXObt8rd5Te9wVfC1MAo
vHDtaXMt76rUnprAkLdFxMM1Eq3ZvP3ojNzkkRHynx4c3lmyo1YbswgjRxGfCBaPyw/EVwI42Xjl
YiLy+Ck3nqezYiQzMsm33YK/z/aSOihz0JCgAfydCZ6lLPg8ia9yVCR+OGhM4YrzcMZVKFqQTnfc
ojURQlpY0zre/Zq+XdHKnoh2JAm4AfiZn0wbbotRoLRsYiHeFEEoMU5WDkVC9FjuDUjTThPKA6m+
XjzxYBjO6lixVlzGypsUEUbSIbxQVH/lHN8dER7pMRy1tdhlMi/PNZGxos2IY7aWJe4YJ6E+ZLOx
KoxzWVGE9S9q6rhOp6ByueFdIW1TtUElp6YSIuVWZ4seXtV9X4pCoIYRjBEMHTmznYgzRrmUc/Z8
LzA1x9/kP4WMwCCvQhyxxjWZOin7gAbLl2kHOF54eSUB4a3zJVDdHg9r1gwy9eP2M6QUNVMFsQtL
kfl3+9tatkHbSfshkZYTmFu+0H1z+seu1Xrwch1vv77ZpGJF+zkt+ZyFqX4YN3aXNkr3IHeznAPW
Kaok8Ci5gyskZB6XkjGQpEFGJeA8YsTAab/7eyuxpgqrT6yQ0t7OE7TwCkH8AtEztJcH00BpD7Yn
jboN6T0lgPT6bC1iyIT2j4hvAINtOxn6ldunMcg2qCSrivL6O8D1LEejYCXtRj9Iyjw98F9vdsve
ETeveqxQy6CTD62jTVRnB+0549i22npdbn4feIz1uCxRahVlKTgpoB4xC0pq4PYjStb1AdTRfY6U
Me71V07AzLeKknP6wgabSrn7KBt8t5I+xilKBS4n/85VpazSeoFNVhWrmmYuLLCtvef1QB+kirm9
wX1439zE/cepMwLQwJ/5kXgFawUd9giUqTowdjqofMi0hjrdzSqdmyH0U/50xLDDUZBZOV5ZtZro
CCneVPmeYci3J/G3ieU03AV3g8g3LF9+zxyQ4Qh2g/RS8P4HPrYf3x77z4rhYMNRT+lYKqrZLpuc
mJ5onqe8nsLxheg7xKNhOUBOAqyybjVlQ027zl0qvtpYSLCEJxVLBYglwmpwK7dKmiJtNmR0L6oM
johXWuPHgL56N/OMVndNkDRUhO6kxyj9NTGxVprtlMG0XI2JYnY5iCFBqO0sjfDl+pOG/rjIN+vz
u2CdSJHvpIzBOa8O+BidopWXcyxCweP2WM6STED0/7EkmgDxLOe6wvCM3lzOSM5+lTjYirfvN8c+
t6R844vs1WjSrHgRcQbqv75uf/uaSq3YNaUgBSGbvEIYHhTHPeWTES4YgG5hsFvEEDyMQhzI9ddM
q42dblxVPf6hAhrJ32m+i00j3XXod0v9Nj+gPzUY8hq9wiLsH4Ro98UYD2SK6ny25Eemdi6nsBaJ
kBujtbC4VwLH+ooVUYnA5l5q1Kt/CMJgbsyPRzy5TWsoxdTCiqM7y4LAqaOTQcIZjHQOtzz7g+0T
82DOh9HlidIrvYJP5erTnLdKcO06qPX+vx1Ub6YrD0keXccsKYacCdDQkOpPxF+9yuORRqYa6U+0
5A+61U2HP/BrbHzOGSSGh4JMGndXkir/7ofcf397lWaJIhHc0xGX/u5iCaI0xtqzynqZp90xK6PB
SM1TFCPjsyogzkhQUNYKre313WIRve02aPHc2g4GsK5GDqx0AjMmV6+e2jhjG/Gr4PMFkeudTs3i
REc3WGSiAwO8ieDvVgQqAR/SRQisSrwAxDT5F1P7SCULxnXbK1AFTg96Dj/khI9b8AGi/IHQq0ed
Q89v7Lo3oJdcHoo65ivacASp/mSizZxFpU4bStd2qXE/dSYuNt1xJnana0EBPTeEJSeO2HVAT/bR
g8EdMDvtaT/tLVLnXTERQaOtZ+eNxZnZf3FC7cyb+I8oJtIM9dH90/vLlLjTfxNnPb9mt5uyFoFW
aKl23QEeEg7NAw+8J3RUAbVc8tUTIrxACL0WdDfROLCKjq5KmfpTwHwHE7NJurIyd3Qu6cDtYxpJ
zqYWo9nc+RvyxgYXNB07NcHGLbTkawuKzj2oRugf4wjzDNPXe/qBWBmOUAXMkzpPPVNw9pLzsKOs
VBswD4W8+3O8KXsduirGOHaNopoGgCje7lohpj64IX1pTxP/4Fc8n7H2m5WVZk6X6ch02XQbv9g7
x9CqCYX8rlHehjsVSbRaAa2I+ZFDhlGlVtuFAqnNUvlct8rVnUOA0YLdltzKasSdBJmj759KT7JI
TK1gXm7khs3gA1xMi+n8yo82acVfpX2gbU2pYSJZb6CvkL4QU8tAf9d18Ffr6f1CRVsfbAzN//hv
d/r4pXRnA7AYoIpt63XDSJQT1zYguqgNORJ/5DtmdySqchZYuP6GUWS8v4ez2o3fmqTBmvhmG/jA
zYhIPXxdWhOGgR9tQhsN56au0cGmKsyub0OXB/nUZ9FsYAPvVl6mJrjCfjR8j582XrHTpE93RN4j
zrCfcTvjOijvrhauVNNyqclDZ+52kG26VeLu4tR4M7iarsgO1GLTwayK3pFJJHwO4VasvO7qdAlJ
oEiqJhSPKD7GzNAWLe0yG90QoaZUKIxr3Fq/BYw+Jfl9glnHt0lucIC4OhSsUbo8dw++rF24edvz
ookbp5VRW2WsjVlPBTpN5gFttDJgtyed/bw2kOIO+/LFjKJ3nV4/N+fvN1c6cuMCBHk37A3jmHTO
Iffjb2JpYGSNGIJvzyxL9n7IV8EMx3ab5dfYS44TbdH46xUJC7RROTjhmoHekY9sdu+rAMKqQhUO
Gu8DlffSnv8Ahi8awyOpjUT7MjZmLVnk2eD1ppUNCN2HH120jLXq/cUo0PFXgMRcNAmVjXHCqhGg
XWOASgSydsgtsfKECtRQ0X/M4WqGCVlGM0Gkv2L/wSe+kY2qAt6MzFgwEhfx71d2flQzKaChejeh
AeQ7qXufelc5GNksvZg1TePjgnyb1mXboeGQ/u1tb3jWCPf3VswzaXFQaZQLNjqmNGaWKmmNewX+
FyoES2AnB+Wz8fgyblZBfLB2SsL5Z01aQH1vbNTOFmccRz/SqGZYAzUr5aNCzm1ox/oS4vSVBRB9
uw9ee8u7cyrM1B/r33kr6UkFUmPscqWnoifhyccX63OyH9/ustAdUemsw2lWYGWshPiD+cyxuvEk
ZvgoRZHpgvv6daZ3Oui9thHoFwrp8qMXSsQeBFPO04MuMsVWjZZzAmakIY19FrPey/Gk8lByZVHw
bmFOmP7l3sL1lmPVSsyA/rkNF2vPENiHyigLaMELuaWIrbEhBUX2sQ7R3633WohOuYdRwBp46CQx
7zxly8vhY6wsHQhwiF2XsOgb+xWpKn7DB0TaAKFM6zLZWQpJrolrDQz5UupWM+5tQRNVYf2Qein3
zhaoWXwIC+KPifm3A59kMvWUfwlEuA6GM4p99qD7a1G4GI23mjUQ1XodhJThdsCH8vXHZQJJQ6Av
4BJ6Eig6hxdrNWRwq4oV52e/G0lR6SyBsgu+QK5Fy870Yb+xQVUPINPdt467Hcab2lJpweuaZZaP
kEEPTEhgbqqdhVN7Z4LKJYZTCPbK1L7KMShSz2OUWD1vBXcsQ4rD7lBr94kBYjh3fGXbl5XqD0zy
tNpaFw/vZwI/wlftwbm1Avh2o2EDKRmIjGvdiqXtal8KcPjo7NMVNdpTrS6rTr+BWU0UAn9/6ytA
217TOcCWLJpyYhEx6EzJNRO/yKFaz/AOuSd8qGIvYO1HNmfvRzOjvr2bt1SuyAsRkIwIuuj++fvx
/1amHBE9BrATyZyhybvBBE4ofrBs1BdCVgCeazTTWw1mthoIwJQWKqu142K/WgIEv1uIySYq1MAX
oYmIlCyr9JQPZuYIPg/hEuUKTEA1ehGbEJzQJGofNLjVJePrOS2l+bdempFz8rqrUwQe5VM8q2Tl
OnivbFUlRPkIbmNYxnNb/9o87FoxawtRYHDxaxuPgJC7N9v8V7Zlt97RINaH1Qz9GI9MURtWc1UL
Aw2YVemS73+6NMHlLvHF3NVtQ+8HJahxlZ8tIqiJRPOb9wKi1ei+rXdIx/iKP42eo5Osx1/k6g2h
cI8ZLG3/f3YDjuJ/Pbv7wcggCPbpFofLSHcvmI2ahtCZ3/iI0yTha4ngUwZKWFgLgFQSCOfEWOEF
qTNvgcHV31VdBOwgh91dzOiURtVag0TnVTenC4UugXKwL7eFpOxxCQQD4sOD13p6iFu34nwAxWW1
iiJU6lYGDRJcl9WmNZ0bCd/o04ircW1FO3IHLaynFb+6ao+3/PzVyr9H3euI3Fb1p6DUin4z6Los
DV3OVosJpQ3Eix1Bpd3qTVBjitOW2B8EWFcqIWI//1OtcelJM3ijuvtFLRKnTHcqjzpGLrNPDCLO
6lIt6S0UelrEdY+oiKk8gwSwSVGvnQBpHXlyefBxybaugCaT3Yyst24Qeh5qhNpFtOGNEbzE38f0
7zpduEr7PKeecMpq/XzD6YGi9vgpsXIcT+a/G3DpIKIj96iVEOCtmu1Sf+7EfbP9QG8c/TzwW87/
gE1HpEJSQyLXVsGcA/UCjGshgXrKM+su0fg+N2Ns3w66ll43dybIfaE0E1TtlNRTRZHOWjs/8oC2
bTuOfc9FKj5cyyPdFnDDWIIXMmnGvva8XS/VZxUeUD4Lyg6Upb6YaD6/uLTat6kL1pzFnUPXwkyb
BCrWPG+HCe+0HrLa3YSpafk9QrIZlu9E0KhTvo2Ps8YN5i6qpTTZV6U3QUBGJvZm9fpS1j5O5Vij
QBjLW1J3MH+wucT7utkCGe32z70s3MUptBQVzXc8ZcF7hEYCvvWPq/6A3s+co+Oj1KKCm4yl3FAs
vjxYaJS8Mloc6BMDqK8bL3GJHX/Hz7mLbOziSmbyIqRiRlJ0vz7doj8R1GMwc+E5VXrrp3pN/0F/
55pSGm7Zc/xf0DH3RhpcYp/Ow3SKK+AFSi6HZXktzaF3NyqXu6wy1n/cKRaPHLBxq3V+f4zyT2qV
UKNqcy4G4l/HpI4WNTp2idfHeU02Yq4hfAPanUoYAuuvOF7NjGPqYWjHnv5cEEUnMeQTk4TLERt8
+scZBWhF8OLS0C6JZBIE9JMBlk4mFGu3tsJtI5rRCNJuehWmvlJ+S9JiNWjrQ95sDQ4sl5Wb/6P+
ti4e9rvC+LWmMMtdNsJAxSPklNesJ2SDS5eiou8bPAX4HBNgJaEn1gHWS1d4BGLywetCcvag7v+S
qvaKNkwNpMsPQr+g2WkbYOUNHb10gmga/R6Xp7tStRyo+DW0BLgZKIquQBA1vJRfEo8pPJrkxXvU
wWFSt5GZvUnfgOKfCYOJCvVaxR0WHqSX0CURh5RJOl4AYc5EGilcfycTbdpG1SjVhpQfKXumE/AS
BWz9C04KYO0P39UE5cn9jEDQnabcB/g29XPsQaVRVTZ9fT3mac7EVZTW2I2f406uoPv/ONiDNYHA
A8xCBs/415J1sQjvpWDvxPA/YjVKptbjv9A3eh92l/jpE4rz4pHDTANOw6fNhpVANBAZCk0Fz0RG
n7RkfdEWWNnscSwKiCdS0LSpJk/VXdOXsUmUIlUnDAZNUKZBXyaeywZsun93LKEVLsLXtxx3xNvr
TDkVqOY4P0f7gzCahnQtyayh5Fh61kv/bsLbJEhNWpPU8uBsxG22lC46qJDSq3AJS0Zg5tipu/56
zQJ4N8G36UMGxdhQHTJkZmU1XIFAvRXwrRFq6z/dy0PKFh+3XX8OUDGsSPq9CHnHz10S703nQmM/
ESV1FVGo3AY48/b7CQILgY1yQEtfd41Q0ScB0iylxYRlMIv9nc2BaFmMifT6iBiMMVR89lZ7JQnG
jjwkw5HXfr3+h/Q/3FW8ehcZG0yaYS74kPLR5K3EbSTJpshoxAecLO0Xsr6G4uXQdqmCtd/0w4U5
6oCg9KV8P+jeQeKyF1oim1/AGIfz+rUmn8Mb8cxpsegapxXFuRfaNcS49Ea6PX9F+fpcAOo7Xyyu
RLYE5l3U3Ml5kOHtpTs45DeFC2RnlNeuxfO7vh427qWoVkTX5cZ7jJmIqL08QB6P+O80jW6EMlU6
iZiMJhYf/bkX+MEG+6R7x424C18Qo3t6DLeNUsi+1lgjgCwlFJFalpEgpq6O04vCr1iboOXIO5jY
D9U+en4cJrgZt29P5WQdMiOZi814SzohHXAYfdJJqKTWWjWWU8VtQ1HO4cHFyaqMfWPePDqAJBSZ
HxxX7NQs5Un2cbBaSx/EZGLjzhYa+rt0tp4W0INWG5IvWnQXWGjh2cuvqvKAfsi5Gs313HLTLPwQ
pQBQDBl+Bd/6SRmtXvCifsCHbs6XO/Nc0A/7SwOoBwkU+tz+mDL5nFRBXurv1qJ7lBVHuEzwGlCF
ImxXMTsmxP4FydKf/0J1nK+Sy5VOo9xpZ3GozSnYIv86T5PUxObQpD5uVgeK8YTNuAErJl/EqKjy
7Jif4FC+zeleAd916EZMX4dgn2f4Vw3yXvqHe8JkJ03wmBtKhkIuWMQcJB2Xu1rFWPuLGMbWJyJW
9Fkst7WMqS7GFIRy0oiu6BsHQ+f70fIuz+QIQLnugC02heM0FERNLPaNQUIWh2erJms/5UQ6u787
4D3o8JOWJ2bdjQc049k5WWMf8BHRdbHvLYFGDLOh0Tqbd57rBCphLuSt///gwV2w5k/wohD+TFbb
U5E0V7rIpiFHU81Qxd0A/eRaffPJYaC5YAEd5ru+OeWY6I7++el92sdQpfB8fEsrFGfnqQH02Z6e
uda+RIEeXmMx4XJ4C82UKwB7bkY1c2lWeSfAXHKIXwZky2m98d3wSK2uf4zCdw4InSsd7f5AoH5V
59nvvIBBLBf3vT7AJqeLULZZEWvHiZ2G9YPemPSW+UEhd3qjqgU8V4PratMJcUIpLp1lnyU3DzJJ
/Emu/7xS4H1XtSGYUd3sOOqKEQ1jGAOcPZo9yQkp+NixcXiYZHRiinmpqmzzDrxYyUZNxjABWjT1
50yZtYNDYRy8CQmtAJGgQaznGULCb3JQRnBogJcTzRX9fmcUsLsagFxQc2Xp31UHR5RdZ6byybbd
E60r7doHW1Hb3syEjkUuc8PalyBpmQBmfFNN6d1p7M5i45a5uCw1xetrmdWH5blxnWqAbS7njish
gKg/lhOSGEU6KmEJIEbXNPGUbiX3wPeHQ1P3Sj5rs77ZI4yxbp3AovXgvZtgej+GEtCY/cz7Tj1L
BkgW2BLqRhkwAixrNgCQcPJXnGRf/fHx0X1HWDajbfo7qj52BTl2m8Z88lfCZUuFO2b2P2fLA01o
hL8bNoh6mxGPUqCi7Dk8c525NqD6ZbNLoIJVnXbKNHArS5/iFtRQhd6Zg8PgFJdoDSsZJjsQcmei
x0tCq6bi6QTSNFHOeNKrv4JdTGT9ySMD+1Z9ikSLFKoHYi1Byh1FLeJit8k2rYOetOSLXrxApbYP
jS3V1KSU10Y/rmG9IPTi0dwtg/J+KyVPy4V/xPs+Oc8HWEEnSUV6t4HmGPaS6fnYv/aZeTnYC/gG
pRhNfLWoa43rJf1e2lRUzb9ZTNyMxiwmJNEau8tKwa+xWjyoFVfi99Aa6lAO7QygKEyAe1NQY34D
RR6d0hS1AmAYpQfr1YgCxGciInR3d7m69PKwOSMKYYA8JrAqPPWoCuVHvVQmoN3ed1CaqDYsR2CP
qucO34Mf13lWkWcyOTMl46yGvh+iUJI1JVkbnmmqUeAeodFM+yDNSZ/nswzzd8O7qSuHtpfpBKJU
NPP31WLkUJrkVDQNiryjHsYy1w0cqhUg25CFy3mOnj2tnmHO4MCT5jnYkDD+uKzT1+YtzSejcI37
ioHJt84Kx2/1j9OLi/+4Zo/DyUY+jAtLoSBtZxXNq/v3lrdszTl7r3QzH9tp5VIauRn5Y9TQgHz8
rEFcHJ200mFkiyxwMn0sY/1ufxurBCI41xGX63clNBd/NqzxroMWhd7MqbJCiKq00UTW2NAoACNW
cZrnJxm9cVUfxnQKlH69m5q3BN0GdkewL8HqCYMeOG7op1APV+QbzM0uYlC2x0f0ws+tP+pgj2cm
pK6M4Y/HH8qxLUJQ3LnpBdzD7Wx5e9UpMiNuKQrH3Cz9CTGXBNxlBioCi5LMIhts2Qw26JcrXigf
hGWJqzaS+/ROTYB42RXOLxjL8+/LAcEs6i+FGvmZgG6PpRWhXbk8rK2lshjn0RaM3+cbejNV5OoP
CjmFQAOt5CyMS3EdvH++wjaPrF8xgmuULpXDZ6EP22GApL4iSDhTz7sLrN5B3T9fz3zEOYjbtOSZ
vS3UtJImikz6lY9nWGZOiabjLXtrpJP8oj2DnfK5JdCUwlwDaFoBphO37VBQ9ZLWAdxUoFkL9QmR
7p+D1BwOleqmoWZ5hNcksmXmjaksF+PFSo/NEI/GUK+zk/IwC/Hef4PPuKShWKFEa+squQA0h8dL
1JQYEmDmiFtCh551HLAkJPz8FR2dmc0C10GYVPdihWIFCpka2Ge5LHPG5R53acZt25YwnWU9nNNy
5Wk7uHik8vc7Lo2k/JuoMUaGHyLwlaVP1FInGDP+VjmT1KFLQEyUvrs3NDwslTjMWxXGwI9oTk99
2g5dp/rPaEus/DlhCrnB6ApteZv0Kuefaxhojm5Hk/waWgwIfOTQZJC6eTK+KBNejs3TN8VPMQSp
pqjwuwX7oHJO7feUN3jVjfWypwHLFD6/Mqtb0NEGQHDYq10WDbFfvPlA6dUqideqWj67uXqBYCap
NXNCvcrQapKTK5HgRd66Am/7yGxZLG0ThiKVwliMrVkqGhZc0nQX5OKfhLl5zK9cmlAb4FgJle9H
zgHaytbINtX5491iemT9dL7BkfyJOW7rbm7ytJhEyo63aCOBDtzQSHLNcEQQNKcvlhAzBGKGK3/l
qO1jxdwVkwfiIMZSer0UxbHWQuNItW/Ye+GuMOr4Fgi2FZ4nHCLDRFd671yb8VJt1PjXEdtCJpkk
4MlM+ctMgBksCYTeiVphfHIyw82TdRKOg8OooRbAi+7ksTJ/tc8nA4I5aLOx3QS/jL7D1oQhfUWG
1StGKWslPwopvNZxXEC4W17zDOq1v90XtKNK9AmbX9h4IDT4txy+jQF81vg8q5XsU0z6lPDB+MeN
m8F7tnM/NGa0kC/SKaN2z46pBvCbs+rg2kFBrxE1rVEKEE0+I+3JC61pDgo4xgNSOifI6uzPWyZK
MxkeEYXbtSzils0eAzXT2oddSrVJZ1VbJC2Gfxp/sRABcFgsrxxI/VhuS4UKhh3PS78syS1jRWU5
3QWQjIGlzC7+s38RCEOgTiJ4AKMIkX3aJugt6ge3iW1HxgfzaC7MJKNg3kvf/0tlg0FC3qcPaQ0C
oN+Ngz8hljdqBLmCyJJbewnBfTWzCVaZm7ikZqmFpeQCbjk1aZoJ98zak4YRjiTkrtbs5l7+vpHD
Pd0UKQl4RqxO5bn5EGLn7VR360lyOhFoK/PMyv/BgXGQASmOAYPQzjiF3sYuhp8ZdLz/bO8jzrcB
mgF4gM7HzbXnzsQ7TU9bBiJ+8XtRnSU9WD9UnNy8mS60585TtmsVLdF5PKMQAu4o1qu4NfPA43mb
onK3Js0poqC4Y/lZoU/CrL8M4S6tgcyCx5U+DZLHR6bBhBLOlser1jmKzK2vfBSR8N+EW3hc6ehx
LRPMPZsfVMEV3R0EOv81DccCJeJlizgA/GAsgWgYfhse5232egp8xv8W9HKLwDJef3pXKgjVniGk
ZLSuywprxAGBkLQxH2z76czKWyzjdwmreox0xnZ6pgcF1G47tD4+2o+BFwFhAt7f8B82fShByDOW
3QYVrhIs9SBMp8Feajy3HCPk44H1j/ZTyDbqB6/6fkk6+LKYvaOgmDzkcALVNUj12/ULv9hL4IqE
6GhmO1l5hY1AGiEJRuGh/G74g6yopDupFGZS+Orbwg+DjdZeU521xOc/gdzsxc2bk0d8OcLGTiT6
ApGMTP4HMXbd48DSw/i8bes0UczDoeQfAAqiK8/3Xx6/dmdgLolTxGQ53wtPmhpI0ksgtpAi/S6t
9QxUs78uYAexS+mEXCtPkM33DeR86r39hzdvN5wJDK87GOa4ECNg0aLhyaTn74w/6ozK3gs9ClO9
2Jjo7HCI3Ijmh59McF5Vyo5kOKrKo1hcYTyQCooLQVv9ewb8YBSg1l9m9S9ERlROBMYukK9L3Qmv
kCKp9USpAYoQYJDayYprX8CPobA9J8vnfSc3V/9wV9b2rN2fVETYRS5NSY+xmne5EWopry2WSIUs
1k+/mVnU8uPYlsSrb240FavmDOUxBSP7m1issa1r6pNlG41kNWJnGHrnfHU42kgKDhhas0hIXjzR
MrrvcX10tiuPSZl7R65ilyIXnI29XS3RQNtVmMGIncd5RHnD8/ql3E6qsIrxuSDFaVRNwGM2A2Vg
NdYHUfaHlycu6+nIIGBZj8AECGbXvuxj9J2MvZGqwKLcwAIFb8GoBJDsGBKjvk+gAc+kCY6//vBy
e5aiDHSOu1Y1UHVrUmdAE0EVQMo5MriDu8t36DJoqV47WyIEkBL9GeoJKaOI7ADfsrvyAOplzxKJ
JyzsmYSPSwiWJTkYc/zQcr1rF9Zb092r7VZxaQMNCIZGysun/z6xSNtqoQv96SR3l8eBJVtnqsGu
lV67a6qb43BZMiU21Y35GOrQskGLZFpWlc07xrpquSPoOvpE4eYpHg5+s+MAnmmrYVGOfs2I2L/C
oapNNJy4scDDi4CQS2eS+uG1B3ZifXEKzcO/ICwM3Mud3q05WfOIbP4r95eic1EHZGHMrEU20HgJ
aScpOmdYNWn9q+M4++yVgfjQM4TgerrG/n9HmWogJ6Snm9WJmjb+PRHBJqXOlTh2Ai5IR9cMpR9Q
5UNurp3EI9RI1pFBoA9iW4NZTi5jmU9XiVHFxMkW0sIGz1qSJPl34Rsrpv7dXewAGVz/S6RB2BBu
kRcr6F623egWf24aSa9cUl0W/sgkuJDs3jPiwjLTz9ZtsCdUedycF76/XvB0HeIJKtwXTEmb8ZhZ
J4/MUDWPOshZhs6Kokd2zDYFvtVld5YMyUFUX/HHUVSlf3Qa1rxUYwzEvWiT9dsH9RoC/xxkwj1G
D5R05f8+2t0S39iMCZA1SP/yh8ke5xvsx9/aZ2w9+hFws+3lzX0ywHhpgkcrXPlu3/FUckVRex1T
UZeic1QnOUg9wwRUvlv0uXRor/bb+PVhWQ2zu9iyR56RG446E3DFy0VwRvvdsZDYvMSKD1C6ZjkW
PDheMspQfBXGGdas0M4QhX0cDg6JuhwUQb350LDr+BjelPTRK5x6umkTMeNZsB0TwaiqoHehn44b
EO+ZNkbxsOyX4roGeER6jERdhSHInhf7LjSZWGUvzkidxXvy5E4Nn681ijVKW2HKCUqQhEknULvP
lZXh1JSMPTxmiv1qMtFR6PQRN0F8nu957FrgtlvJrF/rVALFp6FGUdj3bFoX4qUn+o1oUH6YhcLf
YK7ju8ZKV2ZGMtUyC4EDWnN15WIZ/vp2f3aTcnEOLv0LXFp5n8l8t+nbIwK2NCqMLwANVw25FltX
INVFG1sONdei8jGoNZ35xiF8RKhAJiDEZ8TNqFNgJ4JKEsm025dbpdipduTseTCqfaByUr1HpcKC
2vGKx81Rm2Q6vhxf1EatecoEoDbS26L/VhuNueKSJ821JTXCyCNzJr6lHXGfKFK5RhseE8/TG1dK
np8ORdu+/pG4VUyI+SWpCHMTKj3eVDq87z/wnxuNaq4OFu92la2AibgGWtUVl7I0RfNWzFEx4inw
ELG+6Vyd4FHr6V3HWtjB+ivMhGgLll5l/qDqSPzVrROc2MWhAmyh9puH0jU5P6UjuHJ60FmJ0hTS
y5k74XgbOZFeFJiSh9u3O+21ScRbUqwgaxk9x4txP7TuJntEB7ebuRbxdS1zzeJF2PHJZTaOyvEv
jCYMGs/HaQDfj4svBXDdFKNjp9Zaq75izj9seYN8MAKfIeOr8GNXyzGALoyXnL44kNsBtMAG1dYb
tihWJ87HqG642Zjr5eO5Uj/J7z07w6ZCHZpf8DkNgxP1MZLMGh384Gt6AcNQ0vDCqmM/Qmi0iL0K
OHEnOVv60NNesHrQIpHQkiKWn5CElDhz4CJqxjXm1pg5KAwhDVrsQeNR6skyEKnaXNAoCrHfW6Vv
FRtmtwCHdXyzc+b4utcEKrvOtlf90/743m2dR/c0GMBOSWzKgra0kxfpjLpf7MhSPWjMzUrH8NbH
xjlhyFvnOM2WElOqEYlk4Pprrv1pQaR5fn/5UPiVSoRCjSJoRV10AEo7fMuSL6n05MuaLo/tz3PB
D9hD6QC61FnznV0FnaWAWMZ26lHrzY9t79KAbGVnFhCHAr49+MqgnWC93fQIGcqpja5stwwp+vwy
7yGbE9z+M230N0Qy3hJyggIlHSlWjkdQi8UvxGQOACgSPlzqsmUIXQ7RvFKVn8lPbUC6D1CH3pIi
l4A6mjlZDVWQTq2TBGP2bKbl/OSym3u7OTD+I2kUXFVvIltLzT/gZwM2BOJdv+tkwd4KkZ/IQ9Bq
VukhQXANhemm1d8lALAOOqOIqPhpwpsdADvghJVqsDKhxjMajszUhXtQwWHAtFi6DTbuPLAfCzix
RJFfgc7iYu/Ri70Kj+pOcZHyw96+tusrE0IjVNArGyySFnOLkCJT97kR/eAuO6PFobVndzPRSGXm
LmLAi8g5CELRgcAfkgpsFS0vHxglPfdRn3E68iA5HIdmCjVWl+Km6pTG5DvMWzj9XXsVl6peClSq
3xlnciGWsfiDZrG/RnFuVpozC4RO3po5ilMKioTAVAO5Q71evoNU3PfigxuNq/ENz0EjS1H26aUo
Cf+hr2+62zd/r5WkyovwBZ2tbWdIkSy36W5aK46ppsp/kADIWwv3+S9cHhyCTfCFLIZUl8yrFgT4
/HXbYv3kR52BbFh0A/rW6qyr7lR2OShD9y/pNBFHr4M3NSenzVb1VkskRdPMhG1RB95CqHGaj9P6
yFqt23+3ji9STTcAcw6PC9uaPRn3h0sag5pz13175xSdoOVcjTb24UOSSH6YxtkRyk2cVu5kQa0R
V+b06VK3b5GHZa+d63BCH/bNzhxAxlpHUIHbFVFju1LY6KrDPenVbIf4bZYTLmHmh+Xu6/tiqIvj
bPUcoQ9oc/BSyf+romG8iJhlsnxbvMG+CRZP7zo4UsdAC88hB8OdDv7/TsRIq+7UO3v3Dcu8sgjy
2h23tRD4RmLekvKzmT9EAHmCQ2eoolkYCgBzmYpSCEfc3GRa5HGl03dEgonqK+l54XBP90DKJtvy
5SpHBu0i18p+T3g6ARg9wH7OK33bC50db7VR8cRgsH8U5wusSrz7PsvSjn5MRyzhcYIlvtmNQ891
VBNI6R2rsxWe36EdStZoMVQVEFImLwXofqEfFBY6A1YpuaZ6rooWZXvRCQm3MgXLyyDMBYdUTF//
v7auPW9TnX2iO66Y+7N21UVRPVfD18HpqlmKpDHgWYXyLklqVkIFRr5Veafgi6w5VMWHKaswQT2U
zYRzBE/kvrqwMT7srC0//IzgpAj4huPx1qgqYbuSXXTzPEpilXh9eqOYLm9rWi7t1IS7buAHuA1u
QIor1hWfw9QXNuPoJLm9gkcZcji4Tfe7rkMERFEF4p/wYgItnCRTUR0ltkeCIsQzHLE1vTHgmsLi
d1bqfPA7RFGW6PZkcKF2GYgBvZpUTuKSoXz8HZZgwwKI0vdmrRn+PMjZHjB5QcFbcQlnJprfmzAd
aFw+TIfTCSE2xI3reAXkgxDRide978/zZ60v9yM6knp8NoJjAe2npcrnvvgQ7fvN5lGCUbglXkQX
PZpQhuk7Ea7kqHWVq1aWaKINiMJjqP4XLDOT3Lm/HrNpW5SnPJLv4mjE0fX5Hq2QMfqwnYzz+neb
adGp1xay5Wk6PRT0/Coo6V0vI9AEbhPiDrbo6y4Jh4/0YcfA2xQE2vt7G0kfVUZe+3wZJ+mzmsdw
hsQQGaY/5QJOM+nA94ApttcCdjYwas+Xz4JYDEH3nTQpm3cUYfIrYerZoiYlzP5/D4rrFxromrh2
+lW4/E3KpqlFKY0qcJXiLmHCeldOFLlV7F3qtCocfi0762/CPLMt5asMTzWbcMCh2N3tqoUObDFs
IPfrbOpDf0DifVBdUYq0HQs99/WHUFXNsvMx28RLA7zvS8KAGSELlV1pYMtffkr0kZh3HiEgMbrO
zGHeaGn/dhR8XtTzOS5O+zptQtIdCRjDgxasMWzpFbNI3qyYNJ6dStYHWRbT9Cd8aNBAxpdy4WHY
qzSoeWdq1ZfxqWpLqkx/JQylgAH0qGjm6tGkOmSwkjWQ80V2YyMKEmyoz0B5tH/nRymX/HrsjSKq
Lm4Yo9r87FhHq2tsrNfn2P/VB2JFa7VfkjpssdXnM3vJbrjaiHUU0S7uDHGRiOzLSb6IRSMDHIzF
Bz6QfX61yOTWtuEU9YO1GSBJBCZRts1CvojuQhCccukytY1LRIuEU1o59BdbmgseO50JOIjyKclo
R99rnK6qTPlmXYJLYWtHiNQqD2vGlQbkICFXblIItxWWXo7oqkLINWIt3/+R2udRg1ylQK0a5dSQ
8nFf90NYs4gXRPV9YPORFar6p68V7z8UeOK0eLk2PqL4Ud+coxrTYzGLlD9LHKlcBQoBE9ERdd6m
pfb/GgtKBtzzROdikzYw0f7A1vC1TX6+QtzprNR25666nUxIO9Zwu9eBbKmxBvGYAus7WXKKQIG4
cxenupj5oehgraAYPSUelvj1PC/rxlttuLHgcOYn/TXySe5MiH5Ggv7UHAQf/rQsPZ00j2hcPnnS
x71FbYIQp7RpyAk9HiKcTM6zdOakCrov/+NMxmz9doMCBHvMA4rmJx2l5BV4S+EVOzuv2AbrTocw
YgtGN13KOT7jn2ad+edYbFLDaIX5CiCdRxMfuO28VmdvukRl7IHFNjuQLSj720vcfhBgPlDjp5Hd
ariPN85ApDQhG3XM4jbsqtU0JGc0/HqXkJu0UMMOYztwL4Fw2PBEdcabPHIOOM7TaGH9xYmZ162r
TJnaopW2V9NsH4FpHSf9/opqSb3SqQNpPrIoAuuVyg2PCO4S+i4o0nmuZoqtoVg98JUlAHnshJA3
cdYehfHfPOmwxwojZxqwbjpGiIgXYe/OpxpxsAG8B6NCrMGWrIwIF/xJt1Cji8SSsk5+8fUyzFUy
GpMrCnmcll0yJTF9fjknAIpTHqWqqMa4DZ54KGnZB1RGOQDCPSYRKBkV9DiXHi3COeb4xs8L/KTi
+gEeqXUsBaubvLNKtuvBqQyZa9E+lUe+igyOIBavaEb8V5zs2ZqqN1zBP/KhRuIdQ0+sgT+x/Bt1
LmjOFXp19EoUHoJ8ZYFAdE+omBqDe+bM6Wq4Q0HdmBOfTAKrUF69uAtv5WIQfUedRSS73MWaW5rg
joHKKrT0otiJ36MmTP8PmBsX64tAXobD3oY7AcqTK44JqJfbZNcTsY/N/gxc51tixdGRPqw6zt1S
qEzH1Wv4V+PRSRxX/JWS7aArhrh+MWK8j1kMoOF3EaF6ZCPQoce4KAud8ilqHOJ6tden5ndeaewl
kPJLACkyK9MAHPv571yDTeVuL80KtXq+0xlJApcvW0grUIuSo2eo20+DT+ADOuKB70XalCKSjroR
PGI3pDhUfOC2QAzxIMEglJ30mvy4BOUoiegCdT1p/O9LFCJbak04jJ6LsFpzzo1IVwQ0YRorunIy
PwSKmvRFUvVX+q/Aiy2iSaXegkk4x6l9NWLtRNkK9z75EwqQxrrKoUlHtDhzyANhO+a5YMdur4VO
FrACZ+qmpwhxOHEGsxV1VdmFExaUFBKsAKDptXtpKgvW+9dbyiQdqP/U7g96bkvfATbUvYrktqrm
CoR7hoiGakJqXki9Tgt+nvU6HnhIUzoETj1+KRdpZR23pR9ICdw9MW82KABixtJzB2gdSl4YMz8h
QjZto8akQeli/fRV5r27pIfCKpKEI1h9j/PVn7jmzQyN8E53J4kvd5hYHFwixVEWxwhsWsDt6tWK
zSaWlEpsuv9p43W/0a38W86AAB41h0uxnnqKJwAMJ4dQJBMqgcghcszF99DHrmzOQBikn5utjXHY
oX5TMP9T7Mh9DwSEZuh972+KIRijZwBdrfG6P5U+yxc0FDCsOOyxvNF7lS9H7h9sufAzK9sZwS2T
Bs1fgWCl0kJtjxblb5UFzUMrPhTc6ZdgR7gCdQZ/1tU3Y2j7Ie27+a5RdtEVrjlVnzhOVfKZnFmt
EKKeXSFcbeYQ4D/0hkNtycQrt9RzL2qPf/P0eIYVdojnlLkz4MYUrCZ/+eMgJK3Pm/Tp6mN5jhLY
DfVaFtJ0LBD4vL2dvRBcb1TsCKzvXqbcfSFXvlUetpOrQTAQBgRA0kEY9d2GTpO1tv/+lpm6/RJ5
nk2yhyPVhCXpbfpdWSEyjodJ9Qa6Ym8GjPP7hKgIGW3r1dGmLNvLlFfhPnL85ll8BxN3YZ8iF1rU
cWijBRxDbOV+b4lhooecZI4q99f8+Fde3DexvrUzDAYWrc5zow4SwVQ9tLgZRVRVb2K7n7LqQQRe
v9bmyVCEO++kQc8PaMXo1rxdpu6Ux4tspvBItWDn/7lS5FRbR9EMfctoYEvZaG0zkNyA4BrAB0Dy
FLD4WzDWPTCR38HGvw/lSwqVcAvN7lCflW6ITjw3fkTdmcZ9i9igJrgSsiKUKOumvAFM9IKbfPh4
RSF0wWfpAdUyDtPDwfIR3p6Jze6M6cP6h+yWcXipATY064wiL207T7+GCWWnAZp85ZounbfecX84
WDJXr7rCyJzIJ0K++a7BJEOSp/eHx+7P/eunQZwz26/ktXIkm9B2E4HYE+GMdBpv623CW5rLgVnB
wtEo4GzanMDHmdnCEdd+NKx9AYjNIhGUfCRZMZSbL7OIDTnCkIILISjEAzoIRWbGDglL5AZItJFb
J35aKBDq60FtizG6hrC6eArH/ADl4QTr1J1t3wV8crIdjl24vzYIFm8+WMO1MFg0/nspuny5kNxw
xLm0frlDxPFgL6320girKGj5OXlTK6ObbqNRgyPy8xE/Ntx+0bj2V976lLFxoNoTEnbLPGma78bU
Y62YVZ1B7UASTIVEHBo1ZLkZQQlq6CjZy4W+YjQ22NCPdCbmwEl5YaAqqmLvowGljoRrfJW0Fk03
zDA2D5lQhsn6YRIKaz3bC3qIS/bkgxFFrSft4BOt22nMGnfNHqedCmusAEDsDuHm7dhJmzRJ8ZhG
nHdu5dBzhkYDqtgwE6o50UsG7GxzShTIxS0SxBAvl96b9e+xZYYALjliA9shEYAZNlblzIl8yXW5
CSjgzs9MMqN47Aq9lHEWOni8a8GkcKKYN268m6+fbo90hYShB9a8Oc+NNU5Pmj+WtZGYTpEkvqfO
i7JIteVC3i87CriqJJRnfEC0M9tA8N0W+k8L0L7UB4cigbm0Y480E0T8bqJVgRzCGO6OnDMr4+le
wzKfM6EYT32rtylUxpEBxWXp3VEjHiBsIxJEQgqS6P9TFw4VjitgjpOQVnGV6NEEIjZQ3eEZ2bdr
FzpFiGWoaCUQWgx9BHIQ52dERYjSj1iW4Ne8/SudUgCJ3NMu25ner7N8AQRECizYxlHG4N7Ebhx3
CEfn9H9z3XOiOpnblwGpjBn/Q+CcLHLor6bHmj6jWO5IGvyhCrXaSemj03lZPmOCuGZZzad5P58G
ZdzvS6G7ZzJJ4sZWUjlx9gFFaXl1tFqBuN3/8rlhJwl5nfPpwPD39PeS7vb6phJIvxEQ0+yaKvKr
AdthBowpznAM/iXjImX9wR7dBDHk+aWw7YTOVjd6Qxog3T/Otoiwusa8/nLQT+aFAJd+aiO02eRr
YPm6aBZWeWoF/4xGaqewAwwZWmnhmrMvFpSJuEemqtURA2ZP3uZMQ54iXrb+g0INOsLQ5SESc9PF
zmBRKBFZYpmhZgJH+hkzKj8hH0Q1GBnK3bhj4u0oyIa9NLZt4ttu8sWscE07i4pUNV+AnNym/UOm
5hAfj/lxb8UoIGa/UgCoGMURXEL1NV9ZyM8+NwJaGeKpe4hBN8kFypa8TRLFLVpOiH/SKMzX5gex
F2KCTo/eBeWD/U1fTKzDxcIWvTv5FCYjNQwq8bTjJlWHiXtbqQS18O4GtQTq6T2wLx+9ur7WzcWZ
5l3gEuqwf1XcL60sqOjqHPtwttDhg2VimVtoMSEI+18DXtgPHZ2bgEASrdB5XxqepHFbLekT43As
AZHEochCsIOJsjlzQfsfLEitbP4HIZkhCcsg/EqpmyquPvVup2ctW45r9lKeSHxrH0009Rtw3SNg
W0gIKnyTGlP53InjaeE22WcORQoJGPTql5reRfuK8I0i3sjFoGiwKknOAxhgqbe3de3+3rH5WbW/
qG/wrxUCaHh79z+W7tVP7rm0/kfjnhXgHEFt89MoE+B9+3gVseqysZ9YAC6kAdHXe3QZr9RGD8Jy
JayVoiaY3Rt9imVccNyCs43uVV6C8oSLegQ01Xsy7xQwPQSuAh6DjIINgCTQQBSAWIaE50KH2v/w
3Q5JPEp+fajprQ/rK7NVCjFnQVxACsCowmG3cb8U5VbWLAu+USrvWhN606p+KTlS7l7ion9YFPnd
vpXmrwu1WJYmSIyThyWBqzhT8B4Q+ViX14DREkmM7OUDSh/JIkPqiG9lXQUOZ7/wBby2Z2/oHoOx
NRkOLUMYHXdyzp9/Pn0CD3hq78z8AVPvh+R1JBlHCgwIGmatKxL1UBwyGxfs5WXTaSY8AqbIkRlT
1dlVa1p7IqDGSUI/3IQ3/9F/6Aa8ujTuMykkdf6zRo+bmEjXp0nG04efYgd/kEqiqeKSDz6j8HuJ
TLNEr4b34R2ucrfz1C+sTwKeFzh8zRPcHk3ppy/ivPL0/aqZFeer98iiT+gJbFUFeE7LjULSDCFg
By4budIO6OVnisgkTbI5rkgzNyrpHGkVIM8MVvv7SRBp3jkaSslUMZjifN1riLHFkQDQ7fbF/iIZ
v6Aa+uVBjyPDUKDfZyLKohdO4YAz7l1+PMVzTXPc33XB0o46Ty1GlcjrcR5OX2LNAd+E6Ws+aXGn
umNXA9utsXbFQDUxoDiyeBHsjb9rDMTkOmw3r6Ni3mbWZMiQg/yi3GibbAWrFh8mpFRSjp3poSZ3
tF56tdh5FwuSglsPmh3RvaCCPtEcaLb144qMiMSb4I+VFUacr205KIzM25s1d/AWkHuHyiagsu69
b+Fxs6MrN0cxYk0w3aHNkjRVvzavYNSBY+NuraIiDaIVegqu7wyP9APx2W1yCxQUjAWDBCNU4hbT
B2CjsVpVbv9AY1HQDpi2VO2Z9L4HxFDGuOuMfAKV7xFLjTCPAXciaHgNPkiw3wtM9/3KkYJIQEJs
q32VF/TlocPOA6xL/CZUMLIYeFRWU8kS7ZTZT7edSC+5sCovNnOSYOhcq5eg1eOXhvayttvgA3qX
/2AJWpsZVHdjzlWMexAuyahuWpVqC2NLsxUFuUjT3p4ekXEnICTXTsn5kIoPB1jttro4bpkvscm6
rXCmJQ/BpwHj4hd0ldiaBIePnbDuOp2PLe8Yclc0cELZlA2JPtGoepEFRIctoNFufQvPTnM5QokD
pRcWbUWD8B73diaNoHGrN4oAwUT2aAskkgeYaH87ogZLuN2BNvYexbDmMEF+vrvU+wM8Obx2txP9
xz2LcDZWnkk2X5U2u5IJdbNysx/aRuiyYLEbcGCR0bKo5DZpLqU7bjka2kWlDr1dTGU2P0DFQ5Cj
TOIEf1q8Dr0XDnFuu2o7lW6uBCrweYJpV1VbKL2twU8F6X4Nf2MGjjkJRxLDBgKqtmAd+tkt7Kv4
mreS+EbIbwz4g8UWtZUhmiUUOe5XdPjiLTVOUBiOXemDL0Y3EY2XPJPt9YPBFr+maGaoisrlawDr
3X4mHpHqFTJvBTi4N0gNAFkm4EsxiMrlr57uFEnWCYDT/8lILxeCLkBPCnqfUJaXrZiF8YZg9xy3
Uy09aRDbM++23XJAwICa0bz/sWOgnGc19A7MqFRKyaHm71Vibh1eNU7xnKYC2wUiN9/zSqatMudm
OgB9VnVgeI0q+P5lbsg49Yo1W1SOXp/StMh0PupsNcGp5IVV6e7u54yIIQS7w/DOGnz1r3x5gkxP
IBdpqO4qEmOOKTYsWFnYqDYOCRURV+LZEKDaIITaU+XuoHVWzgThj8aywCaj5u6WDBZurUz08z1q
InjZDUtFA/pVU9RrPitd3o4eXDgNcKjiemu7pe76LjLcSPvjHclL8VX2eOSAr8Qtx8Oo+naWenmw
6Mf/ULt3upgD9qIhHirKzAKMGQAolDL2p7H8cM3NrA20G6HoeZ7el9/NGszJIZGKOpBDNXgVq3B6
4CvOr9kmKRkY5YFmJBjH1PbuJLcdHwYxmCBMj/HuGexTskz4LotXP6Xn4h9mnVpPfvAZJR2L/FKf
UmpsAjBX2w0N4GeoKOQmCHV2Bf/fD0SDNCS1kNQCLkTjUIdurEZS6MQgMefdTIB5Sd2L06ZgEmWv
we/wJ7YWMPIFa7EO/NW8NxKE+TwKGMWI0AusNfN9PrNuw29fYf6IckQIS1kOqqHSol9HN+MI6h03
PB1rpEuLbR+YZo6Ok0AAkuT4iFZTcCqqu5tsuEZMJkqbK8ek5si+0Hy5M0lFfiE1HBb3uogourIJ
2Uz27r07WRv1IRiXV5B+YjwNRPxkiIKKh7NnlzLT5A74AecY084UZu+mjzZz5CCh6YK9B/wTUK+c
QTquKlK/1ILBY2C5TcEUPsw7P9u+Da6SyjGnzd1XLZFHZIAR9ompE7ODvFtJhv7NjHImL+vqdYDt
RIo1VaUAv7wa1zlMOp28okHCM1TiDh5pAHCYWK93VsL8OmEDE0ZrWf/gA4TplNq8G1eei3c5MXu0
3w3SR31IPdLH46cJ/0S4xi/xq6XkeT1vUD+ohn5tRpCfsJ50C9D7eO0xfRqFbYHYLL+srtdYRG7N
ynuwOysCx7wBoDsmx1+FyeRxhYaj1vS9/dCu7sJv8tM60qQha53KtoOsQv0FRTE9eoY/1gfapp/7
vpYyCAPgTcdba6qY56BsdRCLM/9IngXLV2eUJgYs6ZNrcPrvHvUYAvOe250Z9cCAZjN4fKA4nfcc
VLVj5OKqBywrKDgnxjPmskTdSrb7xCfuQjqP2+E4vcHoCHhsZBk9g4WjM95OHSzzE//51gYayqGB
vd9UxakLXOxycFvQ05u7kIRSYOJxdZQ995L9xRU4zSthBwOzIxEqC2yn4yi31L1zfyzFFcvzvY1V
AJCUp0SBKM717CygsiTJffvI9cIGN5wz5VZny+mHqpIpAs1CLXA4TnXYu+Wykve8pNLJ27MUgTw1
X2NGxNgYCGTPfU2ZKuPKdAyiwaKk53liUhXNuj0zHPeLSks0ObCh6Lk/OY+1s2bdWq9nkVt3vYjo
LfP06eUekaVCZ1+wJJWs3S9eSDwoR3EGcUeStc5GMRPEu+fLaB5BHvu95EBFbmgIKfQ7Sp9nq9Uw
7qLH/47KISv4v6u2PQIbYDV01QHnLpKUH5a3GPU66b+rFcX/RHkMJilwFb+KfS9+UGydqcZvGiDr
fMm07Kc31+1ib6e+TfYKJVCivvSEzWUf3Pwc/bnixe4PxZfpGnU4a8jdIXdNMLMiAJvAPU9SMDhY
DdYuHcIH64ox9UzVtPZPSd9QW7IhrNm4Ry4YyuhUZC7/huMRQB3oW4gULnaP7nSCAZk5ekiNHb2E
nAQDi7lXrBO2RNAN2pdEfNBd37CCHKytqUGYkCrpVeliJJSOJKYCtBT+tcJjobgdRhPgcSKZ0HJf
jt/Osex+kNaNHQkWikumZFDS6ItyoPhAriIEQRrrSQhF914RwZcFS2Wns9otSTx7Vkn0T5o7ae8X
LFeCPeQ3rmHLxCTlD7afU8Ox1NchY2He2xrfF4YXDpfhzysB7cs4OUVczyYt4lkpWyypKIWu783S
bTZIs20WRy6xkzfAuOSbswVz/tRakGp9cUycJxHU2RCEwkzO+z0FvsN7rULXMaYQmFJB2q+G+qPj
+1PoHwJaMcOWKoJX4LmlCzxd/ym9aJNFbfBRmO87+Wfvc0TlaSXpJ+3qvxvi+lfIo6hVxtfQHHG/
Wb7/4Nz0v8wtaG5aQV75Chgm17x3LYn6YeFxCXhkopjKffA88nEIdjU1BVwUAscf6jJydW6jorH+
jbR3DlHUWe9rJ7ouHoX35K5z0OJcUKgzX2K66gzEsbyRzLy4Fp9Vsce9w5VdEaRJpZRYkTbD4PoA
DPQbsPFN4I5XeFHTvZSlkh3f9OfEO3HGA6A7WAdgD0klgBOMq+hU54pfv2/rmgbygVGvR/gnQG2G
jvDc1pAlEJUbDoR3RLcF4DeeDwP5SwFzExB9adxktOLBzIID7liKyEs3HhhhkE3ssVkQr39ZhTLg
VSYwYd/YuDmzmoWZj2bwfZvNe1kYY1EgJId+T611RFuaK3ZIM0vimBodgSvM0VNXq6/YtSFM41+2
RMIaiZYBxf7aD01NLAxpVe5SJ0g60L0OUeDBdmtgpU4CAKVgBCk2jTMqnf/fY2Qr2/hhA2BeKPKO
RtnhejdUw9FIAmuabCcCl5uRWTUIKZUHUR5hvFkn4VXlLbpMClaHadFmPZbOhLbOP/VE60vhcw9A
ceDmdCPNWbcS5ND56s+b/7v4r0xAeCPDnWvChHmKFFLIf+SyxwI/2NxSlf8L+UFBj7bjHu5jXmYh
XK5JzCB78aeCZcRzxH+23de3TwAkbiUKXxIockId7M1GtDr1Gy9ZDGnjYwU7xNKSFXcHp9yG7yVN
DI7WqFUqe+Hilnub/noIFC2AeggwDgXa9qLQOQO/rMVynVIlATx7B7jmGHEoUKC5MnzKsVhjxoPo
Ps/EAU3o/apiclhPtlyp7FuufXE8p1BzgUXGK5V89jaaFhcO8+tuzCPK0FtOOyAfrFba1eBawtVi
rIwIwi0VNoE7Q4It2LP3wdFeUxNroeuiI9KDoOW5nPcVFytpRkRRyeNHO1iQrPF+MyBvSj5TMLML
Un/mVMDRYYk9jqUowOewxAjInu+tmffCCYRs6LklqsyFggflAM3s+U91rZa79gYJykvDRKZmF5sC
57MnrSQPyAcS00wmzkee0x+VhyvheI4ji17L0fq337GSz9guA/gZn6VZ6pPMwSB2j7CgxQqm7reJ
Vcc3EUj9Hxj/mTFs3QZFDATj+caiKxG0QoxCDW95ZuMXDfkErE1Eqy+kO9UvUSGtifNZxkmb8bSN
Q6cACPlCgkkOnjve7Ym6IsrKll/6gP0vRi+FDhQ0mVyTethYg+mF5wcjQWZXLOeGsE77TTMxH0Uu
jaD8P6DbTvdnUBt5srU/vGvHZAQ73YYcc9nZ1t4NI2jlT40TBD6QOawL49v8nn/IB1kOJSCzB4Qd
hN5+0hl8qh2kM7bLaexZk8UDyMX7MCa9C12guxkA0c2XaOwITlOJeOQzIQ+58VX5Ub1gFAerAZ3H
MOgYPqyROAlVTa7k0VyGZ91Zyj7PcLHj3Td+5s2hgwVEh4SL/LrdugRCpzrPjeYWM5bSFeqfOz6u
3ucb6oTsoc+YwxEu1I9njcDP20ekpED/139lOXR0qIasGU84wcDYbnfvm1245iPkOOuAmlt5s5fa
mXB/U5pPVfp4OhvihlqXID4dENDrtpPAjEwoIuE4tgZ8wsMQ16TlInMX6IPai1na7Z39XbwBJQTU
wEmP9/j0abf4/Qof3Zpv8rCSQ+tAWmYhGSnb7VWG+0KzUvDhqDnYTJSp5m27mNsuGm+obYIBIjos
Jo2v0hEjGdL3+/flHjoUDUiV/lH3xaixPNOisytX2ZwOeApvKW9knOlMSX7f977yq/gY9zRsgYBW
wsOuOeUwpwAYRy+Yy7htJNGByvRQTQ5g6q82Ci9wgNbL0gIB8zuQHHhcSM2WynR2Oo9jh1NN6Gyp
29WT6AuoBvtR6IMtvjB4sesgVAJMD1QUWzkeoAYAQedh8XvN+X8sUSZUCGvo6BYBeDDsmw99geRp
cG98Q32VyaTUFbZDTofFu77Gx6rI+kq9+wrkVQBk8P5row+Zg3xkVMQCh8PC6bQixQsZhx5HkW2O
KXz9VguKQcC8V8S/vXXZP7STW0DT2wolaCLSTcimkL6Daiy9FbObk3/ZG6MUQNAPnzmmPk////TJ
fdJp+h+5MZUGWExNDU63D5+qU1Xp2u/X4fAAqn0ajH66pS0KGtc4O0jmnfMEHgus2JZqRU48yNKs
VFOm95fKVknp/bDZxQJEM559M/IELZrGkB8vkQVI2im0UR1YLFApOkBeubbLZYKZM01ANzLi6mSs
k0bPcSno5UrBjQG5+8uy9SfrgDJWZs0T+OQkVNlhqmv7JM31jpNBKmEo/rcqC71FpAKd7NmoDmh7
y/Ug8O8D824xQg1t5VB+VZebVfG06/hED4lG86O9SNVUwixXJVKHOFChqSVD42EB0mu3TvsOXmKd
y/DBUMUlh1Vtsm9+mJf8/VBlDK9zdrJm6pbrAspXH9g68OdlUH7r8H0AJ+oIzAnQsbIy37s9CAoV
PbnZ2p4ZyCQW2zOTI21akyhFuzzC5457fXPTZX3W0lJIKxvHl4mv+V0+2F7Rxhj5X16j3GasQrIq
XgQEYAbi6Oy80rjJwblIF59Palc77vZkrWcOuS6OelPFpncGBEzNiAbjBgoiUE8KQvX8SFa4lCOy
wkSOf/s8HsAMp90vMgW9e380hJsXeOeB/IvC8N0qV/y/bJ0D8kdyrvX8QTRkS3BlGMVzF+317fdT
/Cf44+lQ1CvYTrgeAYN+Ypz1Vz7SivaNshzysIbdR5+tDgBGaV0QlgQip78yTbpxqnpur71Oa+rm
WrD7m5qGbdM8+FV7dszJLiVGzhKBqSiSR9/C+SI/Dlg0dyIfC5Bw+DV2QaVx2Dq9LvtEEI8K4f/y
3yH1SnPZVDfgIuNgQ2ha1iPNj8UkhQdW9MMLuLTEE7efAMUIWVNGjwSsgHjCEyyGct2qLhfsDYaU
J8uzHleMtKPE2mfZoc06HezD8FQ5WnRTjk95StVs6PKK4QofvKdpF6b9xZhErNRfok5e1IlwspOI
yDxoQFL+EIrtCketw3EFtkA2ZXOr+ZuT4R3DPNFOq47glTNEhoOeGd/lwrUWd7mSIdWNyYDNeKIC
hUL0ow3gH6Z+aInetgo5mJ/MQTJi2HPAIiwCSUCgzoF5qt7XLcya0OKydhyufIepcT0dyRoi8m4k
FB7bOKZvDtaZdBbe14ndLGD5ArEc4gH9ucVmIGQ6qe6XRR/JcdE0MBOCGgdV07CjoUy/R+sHOGBB
oVEN4k8Anr9SHjBnEpMhYwdOHomw9U00aErVWNLMB8MyVOP64tEEPW36OuuYoA3GSIXDCRlnOOSC
RCY8thVeyikiU8oav13uLZkNJOSuuM2mPShhLLTk4cfd3BNTo5KR0PK1EDFhGW7rDBAu4BxRNgBL
td1cxT6G/1xsaWN7ZDv3m4g8hn/LcH6SOG7tlUYBJAtMqTuCvihiLffsKMnXkhirgBsecScaXhwW
vEwQiOge6B9aBNYpDM3qk6ua/StCQJGcVoL+Mbg5sLkpwuz2fldumsIW2hUdOZVs+fu6YPfYNT/G
n+hA5OTjzub/yAeIJu0Kcxe4s4RV+1er0Voj2UrPamk01qBAV1eeQuTB4w6j2bHqwHFKkUv+ioSB
lAJ3tc9PQvlRgcs/HNujTI/tq/oWctj4qlfw4zNHvJoYREa5YSFt+XgOsx3jexJg9Dqlp9JgemO2
joctp/uF4na4J7XI+S+cSnxvntvxK8kYSHLbySko3LfGLva4DfcSi0kPWP6NF7NUqMeashaDGNrx
sMjTVGgfzkfuvKR2Z2N48bxq8GvQnlDuhvWgJXFE/6VVhXk5jN3Parnha6MBQyjCZ3m3TEYHZR/i
wKkk6IXkrpjtPw+ZYkIRmAxJ1oGe9XBWC1jVQfhDvt/kBxcRqEwLJqEl+75QZcL6B3u4pjmGDV6+
vMvEIf3riuC3sVWgaScz7JJcVD70FJdd4dqIGONxV30N2PN+RuXBcKtfp5v6Y7PcKTyiLsbb6jfG
yYovp+GRsFZliUzEjDQimo87eO/37TwQE0lcUpt5cr28nyslhj2iBasthx5XkXIVph9TVSEGbNE/
aDu8uN2y/xGW1Y0KjSFPqQgmp3gbDtUJkMffb4N1ViKVDJ90NGktCMz3nZkN7/6BkpARvdfdzdPZ
qfUoHAs52hYojhL7Gbe+cgCNp2xi4eUcGkfgGlKQqgFI3Jf8oulpLIQLFeJ64f35dPEy6q8NopjV
nwuODTeSBPPtgGxJaZQAAlUxQytv5JvjM/GDrnrwnIZseuEg7nFgnlQu48lNokw4BIK5nMF+y8ln
CqAHvmYM67C4BUo+C1NcqaJRFkhBG4Nr7JB2MZz7X9ZqG/v8WTQJIOTMNlLas1UgOixiGHbwDX+Q
iw/g4+cOk9FDti9OQmLJ8wBwIu0aOwIRXXGJycc/qvQNypyQOR6q8nTwp/0ds+sRx25uUjYbAxPQ
1ayOu8tIJGxn4N7Yo0exk1YV3FmHrlKLkQAAYbZAZGHEX+++NhpcaSlCksXURi/fV3qwYgf3UYLy
9seR3Tc6Bq7q0CRlFFc3T2aooIGmJ9eresuSb2ZSwiMgP0wrGgqilu/ibXFGSSXHzHvajAmRAWuN
vfY94zDA0v6LNb9h+nwEv01zWUgDmoJa9u7twiMufvTXyuqu0LIUPxUTzxyjeahv0MHpFFgrmcwD
a8i6aKMLcKtZr66ssTi0lRysSnkXCqvJWJmhkHgCGP5HuWyLSfKeyfPhWktDGitWW4YyAz4XSiUq
ncv+R9o2dDi9rBIsgoHJNUTjr10BA55taBJ5dmQgFarHXNfcrjU0N3ye/PKp64m3iyVDV2q7Vfvh
pKOVyl86IobFzXKJEzeSy+RIdLtWngKp0yuNCLAAgzxxcE3VoibKClsyRdjULOuJuNmsm0EmBCFo
u9EMpyNphg9IhwNt2WkDfwxNBsiil6c/eqz52NDgYNWQ79sSg7gsjBF30B/W5UcwIBxJNP77BGta
zWivUefZWA/c1JEvKSsgM3rcNvw0hF/b14LBhNPZ++B9fGImbR3rhNu1GTGwISExSJ8X1P0lJ3Ef
GXusDjN7/EoVxqCD5qmclj8VxoXI87pmD7O32FVFFH19QJKlAA98ultA5J3O9cOfw6numESUECUT
gk9lOhrPVhH40cMs1Hb7j6DtE4OtfHuAhfZHiPzfYV0/37vnZ+WDryB+/Zs0hvEIi/ohCRRiGK3y
IvhbMHkxKxc8ImyYRzG2CZMeMeIQztrx5N79T1ShaAP3COUi1tkUysYBI1HmgNlfdq2OD0LKTJpi
RWhlsp5+JQllPpctXHDTWB4dww77E4/lgY94xBP1he8GDsFO3rPBsZkd28OJa/iftik3iVmTa5Cj
/nRF9/hC1X0zHUJ3jbFzywcMHKBaXFW2f/p+SUceUYKJXwgvgETrVpmfj6KK5lT0HhRyVLHVBB9L
Jmik+Mi7527G2nLgiAOJFFExNeSHF7Z788u5by/ZBQ7IYpopwkB6oIg6dO/vfhGFz7Pzf3l9+0mU
qYE6ZNaNFTJHVKJ2dYosDZ09FJBy9+V7Y+phCrIGdJDnc+sN6Z3ijZRaf5rvc468EH14BRya9nCW
N9gRovUadclc3OlF1AHoXyLBSUE5I/mCNOns28DAl5nvjQhHbQKwiYh+VAgNpAGiWAo4u9vG8iHe
WpagLqLw/s82dQN40sxVy2U/UaFxyLzex0Mh2Ul7RigsjXGJ5010p7LM/YAtazfPliBoGPTThwCw
94xJog0vEim2M3Hb4wNJUBy0TjsjpALLrenpvkkdHKUw6drE8KNns2l3COeJhz6wXW/dzCxhbdED
+1YH/JzfsJhUpED4JhwRwpI/AzkjSFEJ+BjjBr5iflGyVx3O8mJzUDZTGr4OIFFy3R21l8uEfobp
do3PciPUdj+3/+tkKuHlMgAf1XrjCH1aiTsjNXyFb75Qb4FufMRjBzaIPp1KMxzdGo5kcq2LHmR4
gnAZVyJvR1xt/S04Drq1nf2n87fkEk7fsebMZW0vT1/eIcbrTDNFz5PEoUoLkRPGv0BAVzFWkJX1
M321/xsZRsRRTDzKuQAHTUhraoosunlzNIIul+kg9CKzjVRZzu6K/gKxhUj4YiqVv7igR78hVBB8
gbOyT+UA52doGR6gOn8kkdW8rt6LrY/+X9/DMHIO54xiFWoTHoSqZ5Ly6BQZYOSYHTXhRCu1fjpd
gkACUi6yG+CHltojGsX94txd3FbfYW4cCY2kxn9HMfFtNNryid5PbyKSIJ4VeGSw0010vq3UdbF6
HSe39s22/sh4NmfOOYe7N0qhmR13oHcOzxMt5N3KMqt46eupDGhgxa7aTyYbMOvJHGi1JuvskcBe
Z2Jjqh3R4flVSNfXAI6PKIw8981jNu78uoji1zFqstUwsz0ymBk0oiwy+fgIVbP3FXD41R4awRkP
D6qUpjQTFXOieEdSCmSVrywSlp7PtMcJbwxGqQcOgQAVlA+VMG+nDZouQu43rylZwlVK+zGRRVIX
Sv8Cx4ajlSR2R7QeUB8/xBmFF9d8dRWTvYN/HpgQvTw1yAydCRPqUh/kjn/tBT0M1Jls29jG7qHM
hE8gS9fdlAu1CXVCAB8YfQuINZHkD/1kAU1DaexQGEbafSEfzGv5OyNcVmAAguzbt8Iu9tJwlSK1
yPyGKIf9zLQPPdObDlKT3tjx3+WBECXFHG86SuwbDGv5Z80AAuajrPexg817dPMTOGWDkA/GQF6v
DpDAH5ZMUyodAbULkG3aBBg/FKHXj2rbJqDya1f0fp3Q/tHl3XQAzkWS6CfpCe3m11u5r+t2wOMn
ZzIDMN48obcjvPNH6TKzJbJuWo734CK7IwqeERi/YFe5RefcHYXq9vHBAfycOyqvLHfwl9wMwHzb
0oCDFLneWlzvXSmHFNBB3OxhNG8j1Bmdm7AyndMMHlXIJ7KrlpnZDPHK99zRNmJz8ZAC4nNlYOKF
6leF3eQmY6tPd2mjUD2v3n2PbNNfSjPAm/d+9zQhajGp3i3GL6fCX1CBQbOmsyU3tbcUyk5qlZao
dDaIdX1NwNRGXPFNG/jMd+jQ1PZ4G8hzZ1pADD2AyfwW07armNS1sNnCga93jSECxviMZed36Shy
ci1kFl7VEYArFP6DpDosH67Lg3X9cgXBdxglOGrGb1bmFHurpYbGI9EOlVIu3DeymEfc+l9e6ww=
`protect end_protected
