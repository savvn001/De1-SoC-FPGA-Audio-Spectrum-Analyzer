��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	��ς�M��R�s�5쾴�rTP�~%��ٮ5,�7 �Õ)54_�]�[zPE�xR���,�I���� U �/a�x�)69pS�����y�I�j׸��X[m�2O\X�r��P�3��J��0FJ�5aKו��Wq��\?�p�������Sj���6^G���|͉�>9}b��t&��ث���u������~C��qV��v�M/��@0e'��bQ �K��S��k��T�;a7���Ig��̊([�?W̭��~x���l��#��X���m9��-�maNƖQ�r'� W�Pq7����Qlwl6 B	 �9n�Al�]D�5��Ɖl��j�oR?�2qހ����e���|��V#T(�:yk[	�����ȲT���ٔ��q2X\���.��f7s�z�Z,��0�6��$ˀR�/]fәū�V�K%c�H�b��גg��2IN����Q��xn�U���|Hԉ��N��G�l�_�p��5�
;IO�NS �n`�`��㊝T�_m/a� ���vm�B��~��y��V"��UҺ�/le}��u5��%���'M�~W���̕J�Q��&VF$�ZZ.�-%�/�Z�A��JtiD�<���{j��IN�岟E��@�\��L�̻�y�^H�2�5Y�scy�Au���d�q�^��$
��{��C���D�Z�{/n 4���r)��� ��� ^([���;mc����}��y�O��~��7�&aݮ�������?��P,�<Mvu�s&$��>@�%�E\�����↹�8eL t5 ;��5rN܎�i�1�'$OTQ�*�	tٜ��.��5��E�;db������KOjE@_=���r��ɢ�!&�P%�`��Sۧ|ŉN�x[�fa�o�X�=@X_{��Q��(������z<��I�z�t���T�s��Qָ��;���$'<�蛠1U-k�}\2��X�P�b�~O3O�4����1��@���9�w�΅����h�}��<��{Ԡ;�H*q�s� .A��h9u�r��=�=�Eܬ~Y�	��a/R�n�]��Ě�"Os_�~xy���a��?���p�l�&t�\h�����D~c�#,lE�p_���(��Ɠ�l/$�r0 �~�1�;��ޥ���V	c�$���	6RB����	�
�0tj@�ɤ_�+HT��ݣ�p�3��7`�̻Tz��(��Ў_�M����e�|����?�յ����:b�6�?J��} H�����B�6d��n_�~z��~_pMd��_��Y^Kć)&����!=�y~<�l�Ϧ3[��ꈃ�����,ȯ)�k*a�������N��=�?5t(��oIv7�}�����p�ק�b��$��n�sZ{����^9�p0�U�5>�
!U�+1�;WEl����h���8VzI�	�HF�A���;��W�� �H���L��j�� �NY���Ie��B,+��gơ}�>P�����w	+��si/T�k�+����1� cC�Zu:Y���}�e����ͮ%����!d' '2��~�\K���gԔr��;��6)�:?�g'�k٣�Z���y���t=�z�
�z��V2���B�j�!���Ň��K�+7��!y�O̢]������7�>;Nĸ*n��~&�5$��~L�[�r����k8���u'�f���d���!8��Jz*v��%����A�:���ݟ*UaY�je��V��u�B�b�Tđ��Nb��`�A�0��0^{$�}M?�'��\S�[�V�Ѱ��m��_���Q[�!�m2N]��D��Vup����6�֯Y>�||k �i�k]��2��n�����Z�����r�흷SLؔ�q&�qG�=k�M���O��:R���i(��RT�a����G �㑺��)2���M��yYՍ�	6|�S��R����d��غӘ��݊%�d��@���U{���#�u<�ިM=�yg�����q��[@���+��Tc9~�uz �.��)ka���,zl����}^�"WD� �䨱��ؐ�.�&\��$��Fk�ӱ�lEe��ޭ9C�jl�Ŋ-%X�5/�"��Z�4%Ct�������-��gEҟ����,�nD�Ʒz���r[�"�i�R�����9F�R]�2�ԉU��O
�f�^K����Pbsڿ�[�k`i�>�!���Cer�%.��녴M��T0?��L���sV����xY���En	�c��nx������z�;l�&�X�?���8�4�`�#f.��}���R��wo�?����#���ޙ��У;C���T�#���uU�Hg*�&����]Z�~".I<�~>~�fz�U��b@����,��g���G6�������=Mw��@�����6�,;��@Nȇ��M��;'��}ʬ�;<
o�tU�o��Rs�g�4�ׁJ8���F���K6A���vW�F_R[�s��)�N�k�n�4D�F2y�Dmr�T�,�o6"~��D�;$
I�j�ƣ���]�O��/o�",�YD&.���Z S��@gˤsN�(���|���E�y���7�����3�����c��h�G�x����l��2��o�]���]�|�
F��X�ǜ��v�O����T�����G���`������i�4w�'z���t���Y%r0P_Ֆ�#-�Ӱq�g2�"k�3��w�$ ��ۊS�-� U	���GXhJS��Jz(�M�O���>�g�*Պ���eNg/��o2�4NV����ڦ���5����R�d�� Ee�r
�1җ'Aװ�ڋ���DÎ+�<��}��Չ h���l�O;Jja�R���Pl�N� :h��W+�u��(6�b���
�N�{T�
ܛ�6]�L�����C>��g����TO��0˫j>�'H�6��Keri��>�����B<|o�.�� m�]��iht\ǶQ*��\.�/�����@�����8iA#Ŝ�y�m�l����?�7���7I�|�}�&��=�!��6nT��D	�D�잲��D��}�E
H��RL�'��O�
��G������7�!�Z��ۛ�H;b��p��c���6�j�s@j`�=���z�m{=eP��t�t�m�`0,�*�#�����C�P#�c-
�BԠ(���%��E*�X�Ɖ��d��䏪L���?���ⴷ�o��3!��U��u��@��
��3�Q]=	"���N��h�H��3�B>�&4!ϋ��xd/El��,U>С�Xl���ţB��e>�4�׃��yR션����r����7'��t��z�A�t\�@��Z��Ȱ�nVEBF�(3D��KUx=
���7zW�J��p:vb�*&
*���Y	;fw�&M͑$/}�?q�ct�Dd��oH+���-�PU���H�9�P���.��h|��y"�褳v�Ϭ�)X����������{�|P�)��w�3 5#�j��:��{�X�*�c�u)�Wϲ�Ji�����ٕ����E�Jp�U�F��=F�$&#� �km�Y�0�
&�\�͙�	�24Ӯ��u���K�Y̭	)N�6�[�y^*������x��־���؎Q���{�0�n�w	gqW{�^ ƍrghȷ����VRt�_U5R�Mg�_'*:-Cum���)'�>��Mс!�$����0���)ajq��������[<�σ6�q������h~��(��P ~(�YT����q��kyMw�9�}ב��F|���n����}�VH�Tը� ���������<hd�>A�8�DR`x���~*���#���*G��Z}��`���m��w߿�� �Ѕ7:��kY���.Q�5��mp���1�6"�IA�i_��D���k���>�0!�S����_�n�����Գ`����c��dG���~-mP���	�v�8+�l�]����<�+A��8�M��*�����[���?�����#�.��݆�����ld�%p}��7trʥǃP�v[$����l/�E������~�<�g�����zx���h!��Vn=�ܝ�pzK/�.ul �}��1/(L@�a|����p,O2�+���y�?�Q@�h���ǰ���%���6�ԁ֛TI�,�^��#ۦ����SK:6& ^�&��}�bͺ�F�����BR�pа]���a3@�Q�Nruv��Ιgk=ˌZ�i��7������i5،ˋ�&�j`JKr�a���y��ue >c�/-�k��]� >�[欠p��"�=e
�����9�
���)p5Qu!b~�	���֟�B���:O��>#��C�rIÈF�8�<?�;�%%y�՞&0�	��;ѹ�������iY��ƫN�g<�����$�[$=Y2`	}�����j�h���.`�|�s����%v�wP̗��]��#y��tb���J��ɺ�/I�K�k�I|{m���g��Te���Բ�gcNv����
�k���k��<J�wFڱ����N��+���K�y+�-�+��;�֐��/N�9�s�9�}eOƘ�*�<{�[�%�w����b�{P��	nY�XV{�Y��K@�el�@>�@p>ph0ߙ@����3Ъ�غc�J��ρ12�[��[�rV�S@��宖I)G�ݤݖg���iv]��]3d��А(�?�����|h��ݝ�"{p@���m�jt<3G���CO(�,&�2ʦL1�;k>����/D��y��<bv�=�X��]=f%��A�o�c �7�7;��r��sO)����p/��g�}73I�n{�?_�P��7*�

�G?9�f�	�[A/6��N��v��䈫DE�L�Z4U�ه��|���Ԙ�d^��Ž�2�(�@��������a��vzR�oS�5TfA�H�[��&��*��� ɦ#���!u���T�J��>6Qc�뱘�x�?���� ��a�[²�V�u����-���;��0��s�6���T|���x�&�=*��3��dI
�����R�/�K_+W.��QBE}T�洞.���H�����$4��y��LB0�ε����z���l��ʺ8d���m~��e0\���ÓF^��Wd��˘#�a���W��ɽܟ�P��)T�8͈����D*_�M[��h����&��&RMT>1�s�����+;ž4J�KfD��Bǔ(a�������cXy�D��'�����@��>��m<YXG���@��&����&�*z ��]����b� 웉%%�2����	ԉ�&�8ӽc�a��-P/v�x������3��ч�S1��B9�oYK|$-�6���
�f�u���U��3���֓z&
B�k�'��s��s�8���B��Q�_Sd����p�.��
��X���z�t�� �/3�a̾����C�S�GI�!R%(�1�f/Sjo�\aW�.�g�cjb0�4O����aV��/�ƣT��6}6ۙAw�c5��b��c-�p���v��{���9[(�[g��ϴ��AG�K*?�P�MM��9>rb�Ǚ��M��ާ�eм�C��R��m9��i�tx5oָq��_%�D�	s�b�)��ԗ�xOnE��ٳf:�j��|�C䧂���)�L{�^�HH,���1����m����޺�P���W�������'bZ�>������i����߳���(u�B�m�V�	�/U4�� �J8�NI��"����t�Cj��
pƂq���ԄB��:z5W-^@Jq@��<k��^�5��}�D[>s?[(�ٲ��Ϻ?�5"Iiw>����tܵpic	�64� ���_T���F�mA*��)yg~b�������q�pÇ�utsq��g�q���
ߴx���Ĥh}�dEk��^�69���$uS����U�ղsܚ�U��/[�K<<�5�(������=t�I�����X�)���0���8ɠhB��*erRV;)i0 cW��	�?bl�y���Ŕ�qq��
�ђ����e]k�	2Jw*�Y�c2"tY��D��aN�ɇa�/o|��ݮL�Qv;���� \��F�4R�ZG���E����`��-^���+T���Pk�s�b�'�=U��9�ǅ|��T��cG�{�U �<���U���U��V�RPg c��H�ڸn>�>p$&��_h2��K;� �p��1��i|��kLZ�ݦ��m�D��eS��:����3��L����h���~�,E����vaO�/��S�Py������
镽i�$��h�����ZD��l90���TJ�I��T"��G����B4Us/��f+�{�p?��p��T�A/:a��ފ�i[/����y�|�Jh���AeWrr<3�x�+�	��S��L�O����j�[4�Iuj�i�8\�+H���ԍk�+�E3o!1"���YЮ�B!��H�E��+��%�X>��\�t���1UA�}z���o��E���yZ ~c���<&�'V�4��g���	��/���k@(Ϣ߇�Y�4�ݸ(D7��K?*>S���pe�2�5$H��C0U���5���.��aB!�vD/zh��|EjZ�4��lW&t �2퟾�D���Qot؈;����^��)�V����X�֎r��<�O̡;`�z��4���ρc�RM�Ua�r4M/s��3r�� �֜�x�⑜()��UX�%�xJV����o(��212���u��}ΰh��?�u�h6�����r�����W�G6�����l	�W�O�2�t"3NC�	�}��*�@v�:"�k��UpX�������*��*w/�u(]oVS�c�B�S�� ,