-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lM6HIntXSQTThgHoOiYSqvGUKSbAxq8vOhmUh887nxxHUz1W4PSlfrbBTuacQKZb5tAAoX8y0iGV
W6n/O30M77LHnTSpncidn0wBr2yTKewWmsAwUX3vLL25ljm9zd7/Pc3qMiB7anmkUIQezWf6W+Rn
4j3/I6P/2/v6CiE0s0sF3s3MVaJyjaUKXIqCjaeY5Q20E1yZYZqYyPXZOXNdFSbChiCLf45R2c7t
PJMJPv7agLXO53pzOWCpoqEK5Wf9DgxQ+yuSJGGuxUhjWQlOQWMUaKPpnBnvrWkjE58KIjXDxWif
goQLKImVo4hY6jKYnOSXvwbLgDZhKcmQbQLTrA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9472)
`protect data_block
Fx4lOktUixpP/KfpefGk+70qkqwYUGNeYDo6hOr3qJtZiReuqbNlqo3VIoho/7qbUCBEnfhJqnBV
WPv5B2tDbtHsGLEqHVzHvNxa5CWyAJqlK5y1OEijrGMt4olu/h84TOaMGquLQ9NhOrx3o+R+XSYd
QhUk9bDtPXN48D77rba65W5/BgajX9hpLE3XGKWcotevpmAyWYvlUeI7Cv+n7ZOIlA4mB5BT1lXk
staOMhmnB1Q44MqACgP8+YizK1an8R82nDjEDNia+e4LE8Wn/pljVoPbFS0v/QLI+JURHBLBZfKg
YLgxrCPLG5tqYII4xibkuBKZf9aEToWUTuNN6HuD5yHruYK/hmzBq6ftX46ucJCcE9vRihHQxXXv
+TGmyCqg/spJJ+/ltycA9gAEOR9uwfNeazNt6lzjcce2QpZGStH6zxCGDdsgopaJ5MJLhSRorb/1
xzxtooPmMo2c0ZJfQNTltbMGd0PoY2mNK1Kpaq466QJYDFGLNxsq3C80gg2MGiv5BhztIYymGoV4
HKlhtYGu5rpLN8nEWWMhwK66oCt0F5Vjl3jG0WQBS6COK1sziDvqprDT/Kf2OUoc7hksMgfNTvCy
JjehM9Eh0WoSp5EHfz2d3ClKJyu/5zLs1xAVHUOHeToM2m4nQK3GexBiV3/lj/GkJW7daeHGYhKL
rc9BBZ/70YvQS7dIxmduCDZ0qS8nOjRh+HBiSvcQHt0kptBNjkjh4qpRWnkxPMehBVmN4RG30DGc
IC5T9HHqUJgqgBwayQH3PZDxViY9Gk+Yl7e7sWEjNZlWandv4vJa8aUwVKEzu/5Jwvfwce97q3Rx
J3VcbmjJpx81HOfNxPYA3Bq4zhl/am24ij/SWXlM78dNhlMkp94ZmRrk28jPq3DSTBM7t7FyyhRc
vaZeujOPAFjgvKph/hyI1IYLL+5XUixa9nvymjjUahCvXGJzhUtanaMQn5ThCrp4iAvhGj1pdOUa
5VrKSvCysH4kCSXdvU5W+1taHNRgvF9e7IrT1i+xU3pkEgYOy5FWGOoSAmhgK1qTq74UTkz0qz5z
CMfy/xjiLlJ2Wl0i3fYxKu/CLoQTqsKXtGoCg/nFF177J/GmnRP1ERodKFYAdR9qWXqlBfE7EYMo
1US3hsMYG4tadMEqGHz+kJG0R+ju1ZLvvJJlBeczQK0maovoQmPfv+HkrvTURb1LXi7xC7IwQ278
W7jcg7bEJnFaz8yv2+B6sLdwe5bqLy1DMIxxoUj/P1ZkbIs/jPx3ZNR1rLQG6isTNiUPcV+KtJal
sCqy9T7mxUdbl9JxzQl4aJbc0r+uU7mUvLi440MOguEC4Cyci551gBeSubh7ip9Gxr6jkctnztDy
coYMZBYIH2ZQO2YX0vpBGTnDF+9klGmngNKUWKTAiF92c0UsfGtJxPWHUM6G5p3DmZjrW9Dfjq8r
qEo63agHsLRFNaO9D91Y2WvYybscP/Tv1/CSPSKebHblD3H3bdWpJ+K7bAtYImECw8e6M+9tCjgq
d0vrhZ/ar+zI875cnIqeVJG0ujEVp1Pe20yFymuvOHf09iKtMdpbhDAg/JnW+IwU+2PT0TLqES4U
KQdVQm0aSbDV2wBRNUer4lGW+gAS+fn/jQgE+pRHD/gJo8qYqtV7e5y/XpdG45bCd/PEkFPdhvpr
f0camMR3xlGDQLtBL9VNSAogX7QK9WxYEeAiKM02OYmFWfKGsifWytS5MArDr3cAUt6p+jYPhSW1
jfRf7mtwoE3cT7fwnRl6D8HF2aUGGpyNcvcSD5VdQi0YEzbx5vC92b+WlGCSPiLCoZ2/ZynIgp6m
7SJ2duYs9O+o5coPofJTaZrmzVS6ImEwC4f82K7i9q4fK1eWv8ebGv+Kq7oRUo+SrXp0vja7PjzD
8HPsvMqCnOSgzAhqmon9VvG3rCDIUV6y2hH+aisEVmP98iXVZqrjaDwwdC5auJ0qqiLphKcVGUdQ
DK/vFYdfOYHey+j19P9f6B5hwzeVV3QjelF/PaoKj2sT3y4PMrKbIgudV+2RgJ4YrFsnKO273XgZ
/hwUPuSr/z3nunkz7RN/IKtnt6HWBsD3mS4aW7wcf9qW/OacmKQes9gTIIYC/PsYK7aDm/a2fmhf
zN6aJ3II7WFTtqflS95UshOKsATGJshfsoMwAph4LNIbcqXuB6oM9WcAZ82qWCRC0mI7P3BWE6dF
m+t+ijpUBOAPkaGJIQhWJgcIMI6yc1MRB7zE9axk2h6B/uOmeaXENhCeQOrf/V93+jxggtpP4DWE
+xUFq3B7xG7xW/+X7Sxw5BhX/yS3DYf/1ya4YNr6MmVb/TtxJ/+5uq/IN1aHPZCnEMBn6DSjOQpo
BMOX4Wpz5Zw9niY1a0+5CtopRzELL6MY+0/1cQcWflh05KIdx6oge4dbp0gKjZCZ+YiYEk6DCrsi
mi0IYSc0axmyncYjw/wohCm1nqVSq+AHfyRxUoRqAeXeBmdIY9bvd6YjtdH/S7T61W2AhZk/vlC/
/vRh5ZL9uLanxuFsJMQtVMBpp1YbLEqroySw/vJpimfoG19tG3GvaJW7kq/MmWqu9BqhR4sJfcbZ
x8R8Fjj3xWJ24ULgobXsyI3HvOC4PY+T5rlSgdDv/9eAigsTyhcFZFXRGb8OL0Nzla2x/rqcaoox
r6wjppQAJbGeMdIcU4c18Js6xbXWJ2KOqW6U33olK3fpfTAWDbgjd/sMPCNnA0UTjEdEApkrqCBG
8MsGroBgNFvzahLh33GArgkkGH+xAuHG4bNfWFxwoR/e1382/xq/l+ZbOfRLDEhGfEbp9Uby3Ps/
6aRtO6zuDw3u0KgkLBGEQj+6E7Hwm9p8urAIN1uAOr38ZsQlOM17aK3mAwtgKi2CwtSMLqyywteb
OZHN2ZEw4bjqO+FAWlBGC/9D82RofDH340Gl/Yu3I8uxuHtuRAxTC+juLsNtY4RXlJs7sxyPeIOJ
WEJnvO2lXzYqGbHhC7MzOI0jE/d10fR2X+gKkGQ/3WRyWDklQ+TaF0lSKqu+e9z4hRwScuxUlnoX
Ue0E7nEiYUobBK/UEo8RGugb4mRm0ram4xvNuQzc5MaXwzGAKYIwcKWMCLcilY+HxoWe1uL0xkae
L8iHRUYLktnDaf6IPvyQm+Ch/SrBMkdEA3lfumsPNDoIviAKK9RCPlRYHsksoGPxI0Fl9swXfpwE
Sc5+pE2/P+um2NVDrfHJU7jjjipnBgiu5npKtkY/Lw8XEMRwGpu+eDdIumPibIhC/PyovwKNcwbj
vs/4YUUBVG8Gl3eHd54Ast4YrQwI6/XZTp3GNsDVMgQXqqm1lVwXTx5RJDqjav0AQpdfE406rhaM
K0CaHEJTlJPhnOlHJJYMckYGrfHa/d4icMED9/NHcDUXFLbvIoFE4SL6QIl9Sn2+dQSrinJgMaa+
3RzX3/UgOyhsi1MfCwPJqSoUKwPaLnsxkpQXn2Q6uNh5Uxp86QKwU6XV6xli7B51nj37VtKOUTAt
82qNVRmtfe5BkXmySigg8+/GZlm+lrrYf8li80eOtOLdX7uxbI2W1ANmdtjfzGEvp+bIRqtm4FGD
mBZvPGq6pptTCYHh7qt5AgjdEnZB+cu/xxqvwGEhCdHiDr/K5V+9KeaLyP73qTXfye/7ItUfkI6C
KXuv0Gr/tBuyuuvJarRHlJ9vpuWFByJt/x2Kr0n6QJEjzygruXHrFxeKKvWApMWeNP4VRL3yqnFH
026oh3quBRDHJyAIsyaO4vscy30sOl2DlAII1avol27WEnuRjMjPO2JlZwjYc8vQhCYNPJ1Uj6Gr
be7svWRN3FmlJpV/wluWA53+3HPYiFz0u+vTZ869+n0mhebG3EWpRpBg4hnMWLau+uAzf+SDmozD
nnFX2aBoxuEymo6QGeW1bOni+9LQntGF9U4GF+uVdpUXGfqBVaHbIREQP0vJ50Lg29ik63PhcmZn
y5zyvr2QBIqg4ngEFp07Z6FjWqF79Ga860l4bCNfW33d7fjtDJdZ9POjcKTHGjq/17TO5tPkTxiZ
pXQddYnPiWVjmKeohFYWliTu5xtm3jE/C5NPIptfvCC9a2sQh1uVCVJ7IYmCwygSMw72NrUOCONz
wRvoh3Nnz1o/8yiGjE1RPqt7HxgUHwWeTZ+7AR9eSZre0T28QkuHWNOE6hMv12ZwJCaNhCKVhj1u
qJYIHmcXxmuCad9oXlnaYjm9FERlOYLT4fEnXQqgqZx1SJRKNqMYaUHXqFosXLsYieq3ao4w5A9n
fvOQ0t6P9i04BzIGm4lZ79L13rZbixDn/11Va6PUjiJCGT40ArN3vZLnWh91Z04CJD+VlMfjYkX+
USYVQ0nXn/Sww8N0gLQkg3kxcT0tAHTWv/M9iw3v3Na0yJIRvQ0OmiE/+fNfoY1sBlhTuuLPS6Bf
E2gvJB6KsJcarei3jQC3QLF9EvTSDe1yFBnlSeYE2Bz8gLArgBrQ7MZO83K71igsctGbNWStVDPc
gn+Zx59BiY09p5nXu5HDdfMK1n102K44c1UcFWYoiv61k6XfeaCeQsTL9qivMK8JExArQGfS7QQT
uV7cbNUBKWJJBxNQkFlWZObq+Ugsyvkc2v7arBD+vgQL8Q/+nP9lZ9K4xirDI3X/iSv8/1pFpUu+
Xx6z84tHUQuWgnfonnMyou2efWFmcxEw1DvmpDsUjD4yTFP59qYTkXISFjqB93EwPSiLOloi4Lp0
OY1S00VcEikqagRDVOOZHK0wzlI5xpjy3+i5GhqrNZoSGgCjvK0EhPR3uwgl/tXJ+wMQyHbU66og
dG97CN8jN+3wjXyWKRTaiHw+wyVnHXGWkujHKa974bFF+/bEjphLCEPHEUyWsVVZYhoeNjrTSTl4
ve1F/Z4dzdphhyhlukl6nvmbPJnwU+Su+Dse3OhJiuHEH8SLLy2E1Az/cOg8JV7YEK0Zrt7ikxzo
/LCiJzXuNVmPw2FIvl3jmxUVPqRihogfHaUhuu8zXXjvSogVQfGB2jGNUr4QDy2Z1FkbPwt6Jx96
JPopWO+5smiEzFCFieoSVyvUY93tgFyyXRv6cXa4CmCtPd4rQnO1GnoGhTMu7xFon5j/NH9Mm+CJ
fwNE6KVw4PE01ZjZRKnHfkyTuF8GtrUK5lf8AmPMiA1LFcvdj6RzbMmcjzPyt22mrpzNPHM92SU2
UiWqACRuxEnhVWegdkZNOHBiVCjHqeHdE94uIcstWJaWalIUCkTiBjU7w5yTMMZaOm/6i00b4/5R
sGBO16ju3rmmSzC6ArV0JARwfBjY+r/L2I++GX+RJut8nhDykcuc7TDLAVZOKBMjijf6bvkyuQO8
q4BehCLnOOcxM0BjT4MkufUdMUg6EyZDQwNGacPvFQfuXRK1ofaKJ+RaXDe06jVzyb+1D7Q7Zv3S
LhoxNwcH4go+J1EuA9PjKWPEtDWlx0hr6wfCQe7j9ew8timt6GwYY8uQcm2SSU4vzAjkJcKigben
IduqilDSgj74z61wJZjxM+cNdhCCDrB1kWkztqAwJpud9nlWX/zUr4l1EHqGRv+IY3lqhhW4h57p
d811h3xvmOuOsbthpk7hfMh2qaFlfKGNCBI7p0XbEURw/E5IbtqHK9wJsM4Hgm9UtgRKOLnpA8bQ
gL8AS++xhXJmq5HSfiQjvmPoQlBJFtfcEQWOAeiIqEJop6na5w54aD33e5RNcSyDQqyLba7jYZP4
sArpbnIumvgkPic8HpCyB+/K6zFYZJ2fN4cU+ONEUYptPtz34W5sscv4/zNjsplcT2gfypEKHpnZ
RCdfPjTfiqS2XO3kRDHteOh+hwUReC07qR+0OykaxCh8LYS3ugB+pVgqD0iY1NG0b9hN95Y+Sjzu
bOaxGkXOBXKbG+1S0wRXhzqjPpdGJb8Ugcl6+Z/kfXRvTfxPYQ3iB+vzxpQixviKigFaSY96kQkM
GLbe/4EeEEtla+fAa/0CQLdLCFKiLK9P2co+z9TZYS8Bof/DTzEzzC6HjuKPC7iHU0WbV9IqRq5G
jnEHKlR9IOYxPspAiKQVfzxiTTgFarYu7ilTb6nwuXsQrj2BpFr0xNhrxWvjO4EI1ZPi5sLEUvNt
dbLvNveqO9ichLU2kj0bmxZTuc5Nw0gdGsJYWpZGM7/fToFWpOujZfAItCRDqWp/TdieTwHMkBDF
Lvc7KDl8+djxp10a6wPZmFtz0tA/en7l4sm2WFaFl3WkSPVlYzt36YRIAiJzfD8EP1EKsaCpbdvU
EjorbVdaSpR54jzuGoHz5kRCYCv6Hh9qCQ61wRz9Gx5g7ACi18Djm3yuYpCP9s0EKkymTBWj2A0f
H7q1XPpxrQly/awVko7oLTC79VtdLbm/GMOo+VfKOvdRYGEBrscMyhWLebR9SaCP6iecqCL2W1DL
vpeUvYP+z/6Xik5y7ru6rOE39Dx36XHXRBZTBpEknOeAURV9zfIogTqbOxNDUuap/DdqwurewFe2
30Pj11UcziSWlif2nJL8sb2SreMENBjT6pciHNrs4co6xIm8+V5IwyxKDFguG5Txm1dABdzcpy7z
8N+bCdQks11H5xP8wexqG1KfJPUY3J0b9eXvIDzBIabf+EsdyJLBmRt+zFPnXel2zqRBOxqOSKuX
sTLQnBlcwmAn7h3i9+Z8Q0LYTYalN6hdVgQlNw6P6EVPQdBy0v9bnt7aPMgupyxdlv2lGlAFbzgi
dB+ojhhffBUhUIiUrvR2xjZvp3gAtfS+lBo7Pe3Wz5YZuc/mZgMdFhbDhykxd2L73iPePlVbcqKo
hZhX8TjdJaQqg/kRpTaoKRaE2fCoX9CBYfy6Jss7dCsPy15BBGjSNIwGwQROxO6vKv1pWLl3UVea
TKXGqmQYxCyhkW1YnTZbcU01CMc73ZfR0EC8EP/84G+ca0JmqVa/tlNwkXaBVXVdbMVQWvcGXqp0
vxPVANIdgdENFu15GC1zQmXy4JAbWj+FLGfLsAjroXZ6oGQ68UM60DRj+WI43DdV/IS7QAISutkf
qhYTHF21IpN3q/6ZlyYqZGEevmpmKXgRt694Lr/E9evLBg3lRNpsQ0jGn6hbOMDoSqSQWLs6b2zE
vUsH/WP0G0jU8RLHN9WCpexk9MkHEvzS12iaxKqAnoQUvbHPwxCfH0WXoHKevxtcewoA3bOeUhmN
WQOMX49R9YbAuXEcFCweEjAnhJ7BQEVIxjIzEAf8WiR2wivYKlkRcD3NMf7Ky5dV8dlZw3E3fSa+
wg0c6uNv3+1SnV9nvpV2Vw0q2p37otVH5hsa4+hY2hP+FZ4TRHVhP1wRGtbXf1iP7LDW1ZsWS20V
S0+Y1+B95yBFR9X/xw9geg0NM44rxvIRkcVm2qTVfcmQ7BVNura4y4xRT14ehFQ9snjw5eKf+xtv
5s4wG47GVO9NV+P41gaUqMcj0ttdb5sxliTsJL1EuvLss3UJ0jaN4JwKVgkY/+vjWsCB/KKEsxRE
sQrr35GWLY3KDPYIr+4vCuVR62n2lFOzpseE6gQK8vElNINjnAA5tMWFgBAQBMMNOH945mvCzNkc
qw7pSY+QN8rvqaD49Q8dnsuD1nPkWs0f1//kJjg19BtnfRzQ51Kxe/sM1n8oU1ED1FPjSqAH2s/N
8IzPvdlemjACqWs1MsvkW7vlq68qS9bI6nuCbFU95UMPADj51B8Lzw60QWj+FtqHXnY3d0nxKi+w
ea2TsGPvSl17bwukFJDpV8S1e/5BO+CovtIemYbiTb07kGXi9Ea2ty4OQbt7EKghjdUfG8xDN8BD
NjNY9jAQ+awlicmzfR1r9BTY5zkm++YEIQSUP5iz05O7dUBrAMQduXvqe73Ikh/x90R1zw27um1j
5TG/ZZkVN/T8qn/W5kzQs1rDG7zMUZhynPAp07tKsTQ7AwmZfiXN5jSld645O2ivki5barw2hB1Y
Yvl09iEzUpHgtBphkpkOosuzEl6dMq2nE0kmZu0YisI/xKFUxGgSOdTRfuNmN6bGP71MCs44as61
jr5WRAwY5n3/zhUvL267bFqMhABdzV3FzgOI/HE2JPSaPw4jlxgqz/WUgYdi8rgEyFKBmth5AOQ4
pPI70KMselTYQCSL/5Yf02XL3mWTQ7MbsnUCUUMx13giCeGfeHxHFKXpxw2PZXFkLGPUv60AAhge
NO2wqQhdu2YZYvZGOFUkc0lji+QM85nIpKoNQoPymobQRarxSmDV0cRsOHj4rYNylyGc4uN/PWSk
XVG/i8Dt/HfhCPu8NCmaHsrbpS6/hbcaS83eLur4qVF7e8XMv3Q3D0M7Q56qBZcaAHTfADe9u++C
rK0tO2RuxYJo44jo2+CAmgpNLHNeTcPQjBbXjxB16pKspchvUsuWR21GFZU9g12kS0eTQmYyDJ4P
Qa5lcLc6S3RkXLIoiFamK2wUurTjubK8gTwXbwfd1XMATE3+TnNHA+V3NaodzMiME9siAyMagyFt
0P9oOsUbPV1oUFj2zk5Oqq19oqhZf+HAzudFSOp2JqWDI0mEIVkxHce9g8tvzprj4v/EFbspEeyQ
h6dqlqBwZJPCE5rY1lVykZ0MP1v0AJxsp6EwD4SBvqgg/jkE7gZJsNyLnOd3V1YzYP7gj/0AyOcG
Ci9a0FWszvOJScOuAfhYsyIZp/ttHTdAQAtosoZOEQOxnDE14kPSmd/4U0bQUY6pZw2PW7mpSgFh
4uynS2XZsCN+xzKMeZ+wNWKMR0x0lQBymw39RRoPxFDV/MRXq1DanLvwmZ3gT80OEHlmgfeuPufz
J2yrcQvQL82AIJEyUH1w6a7iDvYA6IjNVoqAEWO30y8ogo610aqifkC1WUV3KknEpa20l0hyOaSz
cM0ebK7yFikfi0Ci242SxsZ0V+woCO/4O8VYYrSWUhrY32Z2mNssl07thmSaleHFUSjhkywDvyn+
mXsijOASBsxc9TE2rjY3LFP/anb/8R0ytEHlDQ68meAt4tJQZjooGlQJz+LgzOkZABkgwjwAL45F
1c4EH65pNsBJAmP/UL5cSsO/jLNdwZtA/gj4gDVWyH1S2OaVGJAUyQfcs9KcMm62P2vdsP91xAr/
7G00A/Dl6Ka8SuXxI8CBljrLo9enBjZ+9INd8xAq2bzNsduwfT3ou4eWCotUb54/9P1SE5PVi+Ts
tqBI0LUnK9TiDC7c39Y+Czd+6bsPmeHiwcX02wMKzpbNMP8A8hXWD4NGJ0pkj3R9B+RZ4AQ8o0c9
jYnwKVzUcn1psqLnEkVX1oxZlkTsaN+wdyGmi30fVOqrdci46PieVekoAxlWRtuPq5koWYdJrUWV
+RDGtDpDhM2BOaTjoN4fT2KbJlog/OdtjtkYNhAqqpxYGSkHIsk2V0kjXBs/H7gcdMU2c71emWRC
3xpK3oBBDyqP2zokaWvYH4bPnHOxHtf80j5UaMd6lpEZaHwtRqKeqGC23qX2IIkALzhtr7F6Wq8k
GBO76J7sMfVi/WPCrCvJPj04lxCNASvrNz5WaENfmYaSjY+8KP5EgkHEeWtGl+9fbuS7BvzmLIwU
773cxM+BWRYJ5UvKcwBM2w9ag++D+nqtoa6c3reyhF4PIpW7kxLFXcefxvPbaWUYJ5PUBv90i7Ne
2WUbtcNX2nuzHFC+Dsaqo305MBnBKudZ/bZ+zfIPO0U30nXdmn/UKwr4vbVjPtirIkUa70HU1V5y
yvLtX7eBSqJ0ltB2yW/pmW6GDvZjbCpNO2mP9+321tW/J6zLi2FpYlnlykvlwa3PkhiCOLWj8mKp
YYFexX2vBTjWJYSo0ZyxjA5TZgK1S6l+qfBDpGLQFXVxVuCLGeH4g4X5fmb/dso4h6qZ/mWiPZC5
8m3LUBnLgZfsM53kbfnVtdB579VN+Im0FycuMfbMFG4BKkBebbAsLTuiEPgKACcsIORkOU+P8Dpw
wCqH6ocGbTccfuTF9uA68Iur29sZhGpMpCamU0H+qKvNXXlUZfqViumW7LwXs+0GaH1sFp2k8zOV
6g7ZGKFu/jkFC9GbbjzqlUQVln0Gxa0oiHRmawsmb7uvwEovwIWF79zfRGJTif6k5uktPfB51brN
BemwSmq+6dDnHRkXHUUIlSh5m2FQ+ekNdnBS2+AKBg3YxCmKt+ggGH/ReDPIcCN41oB2j6UgqHY/
ZyTNN9FGW6Gmqm7GT8PhtsZHcvFrkxAYRbNIQhxzBDNUd5rMQjMfRBIDqyOF+2jAKvQk/rgkZI3b
IBJR7WMqFncVoo9zk8xDO57nFjRkyMTVtO1ml4msv42Ha0Ys9Z52w78YhVrV9Z9c0fA2rnYYy3CK
+ZuPH7+HMEk/t/DV4gMO/6zuJ/fc7v2nQS4v4pgezVuNk8H6zVKkzICpE6Q/A8jdY9UPjQZZamSx
uebAd0zD9ZuSbkJMVsxNQEk3raXOTTLMQ4ClWly9R4I97p7ZVUK1bVsAAAnzjc7NoaEgA9Tpg9NB
dOkdQtKrWJcmvUsocMlQYbzfUR/TPo7u8yQYjBva2tgQkk4Y285UqICxqNujV+minYJEfwNvDv0k
nsjOYD7Qgpbw3+1ZMU+Q5P2r+o0OmNhpUEP/NHa2TDo4iFEGSzKwVtIadnOwAaG9f6sW+01NR755
YigZ+T+03Y1qiwQ03O/vMj2WtlCDmMqtThT/pWt2WjMoRJYWz9wJBMSB0KVEa/izQHJzaxseBICP
XuoKOW/0xiT5o3rv7UpWrkcYX20vLi0zNp5mY3omBYd+Fl8HvUf6XcQjHSxWKmLGgdHIa92tKyLl
2gFQCNFKpqzNVEIzwMZM11q1GI9Y0B9iIyIIDqPf+cJpu7jYaVGshlPVqfoeBTaVWysELxJFE8DM
5SmqQUzwgW8GzTfXASPa4ztdSEHU1oeCQKZh1Dq73NmaQSAwzNC1dQ7qgvtj0jKUvl0Vjx6RCmZ1
62YtnK+OqjheRzOAa2Q5Z98dbWLp8OCQkdF+EGDO29O7V58VwRnWUpraJRsuFg61529TpoygWI7s
Hw2cZd5vFoICMHQF/YE2LUrB16nl6f0LCdEjWLO4NkKNn1nB4MvWIMfDlIesWl7hbDxn6KJkQXd9
Oe7AT1JHNvquH3nPSzcw5zg/QSVkl4tOFWlrmbwXczaKmk6XQrubN4lunJG/uPzxDH3mL0wR6rbX
X6yLE40X5joXf9C9opK0TeIEWbzD+bMfAqyuwM+3fy1JSAubfQx/nVR/jSYAp3pe6j269xqiV8/T
T6IjU2yf20yc6EvpBqe0MGTaUfli7vL+phgyVgpdnkgyT78dy+4CDb72mfibGcmVqKzwvl/2oB1X
33TTkWa1SQ89Oprw9wxctKs9kqNtyLShMmDA7ooP91VojfWYkqJZl6kmHYZdNdKZ8qpdnQTKfEQq
Nc7ij21SABqAA2WD6EN5t9a8Zc01NN83nP6qsP6xcfzR4UkdiLWLFOxHHJaVKvcl4JHCCxDe68Sv
K4uKLgvRPSku6b33f6MbG4whdJtsUK5b6M7FxTkKlYO3Ms9O3kGUmqQ4UeefkTqmlQkN52A9esEJ
0OxE1ErzWFLru2SeYGpjwr+P4aL7BAhXUVxfwFvZXIXbnD3yDQ+YBmlOXknvUan4BK0egJqTNf+Q
oNTWNbBwpabHDTYUMcgXGYWSr2YjVOkHkF4gEAWmRyDbIvCw1dP0jppgvyDNIlGvlKpwiWLJICin
C/YUtAsGXLgPVpdrInHxiIVfUHzmo4PmE+M0DnUyCKJl2a8vy6Yv4ZsH94lefwOqNtNWM4x25jCI
Agf1tVIPU23XP9U5DufwheSCUQcDXZQJLHlpUH2r5fOe+D4cXHAj3s89YGHQOsaV5D+vN4QSEGCp
/rWvxS4BUyl7VoDiSf+Ot73C3kMbCibzsqZQl6Njw0iuJFTRgaJB+POCDELrkKSo/D9Qk3cI1HAa
JhE/9X3sAHq4dskCiebnnM/XRlkwmwmsTrTzDrbGWcRY3Ktc2lhQId6EvYc1ienRDAAAKxrWSoJQ
67CDoox1jY47vRZg2wumaGNNwA0LSRRpNrAVsvPpuRUht1hgNty5Sdga88yHXSGaAGyh05j6dXDU
mvVeXTK8IuNIx9pEEqEoX2noRN7M+94Wzkds/PCo8gNNM3PQbUlVsZiSXBgiCjSI1CY7pq6kt+eq
SUkek178LKnJNUIgFaIsBeXZAWorJk3cUB7LuUvRJNYpAMYbiKgWe2GPpyowIOb08Eh3McYAtW7A
jkCoc+95cJRtDv6FZpBcOhEXJ+2CbLvKtJDSyQCNU1ilpPfH9w18xi2ROOWUt5b3zexts4R9UW7k
Ep4eQ1ywkfHcYPpnrE7O3gJU/i76AxLD7SP8Cb76xYwG37HtYZtVEL8IVg1n+aJsbMi0p/1auXEM
/J7/znPmVza45L01TsFG7C7PcrYUTHUXiQO42vcj3cmRG5gBp3LP+ETmIjU+JXpdGTSt9UwdwL5e
KO0D43xgnG1dxv/6VJcR0L/YnSfzY4oaQ/p9i0w4e5jkatFjRJSBFwO9BhQcupYTGWLrKByDLpBp
Cf82R55vBCZiQ/+Gx77Bbdv8+Iv7NflakZgh1PcxDPSHKJSAE9n0ZJpQ/7DkAbP4MLpCNMzriFKr
6CjZhGwHlgBdAJxTmDl+hLk/OeTDZFFytiGJUQpliKyXExiMoXIN+z5h1np/vol4nEAo8ZY/eCk0
j5aP1f2V/cAwtA==
`protect end_protected
