-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K60kHAbwXn/aMgxOIl1KpRpztmucvWNBBiK5xDItaCIkvEKFAiyY8NxiYqaamsqF0KpoXhFG6Hvz
aUBCrZR0TgVoQVyZQfnpDJ2dNDfy4qqNYHhpnsBrWnVyjLHXoB1qPvuUyXFflOizWoS7xewM4Zcn
EWLon+aD8Vj9/zMCIqgvH35Whg5+clKiJh/BSKquxCPPi0baG55gghVcY9IbG+rQKmvfefItWFSy
4EYKRF4P2L47X4UBQF8oGbPKeXE4y9G5Tb5bYvJxxVLea3sNwBcU1CdOn6A1/q/xtIs4NXK1PkgY
5FyfrQWjlx0nDmI+Pu/X5EtcAThLmLSt+x1TUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9904)
`protect data_block
IMKCuUZZnjPNo8l4iTBy+gXTNRChjv/DwmlyVD4ojweb0+3tpJcXukkLB9E/WdwXad8bQKr/44+a
7dcXj04P+x8K04wxzcqFHWBRTei/PteyRkynT+o2MNli+Sgsttg72JdDITncDUOj0E/EhbwXJ7kF
bQ9vDAeueIpFJkQ9nVYLkiiqzvKgBGztrtJdY4TDyNxIwtVagPBdPpwCtA+QPvWaNT/GysQvXatK
NhxeHQ6YUOXgnuwylWEcfY5ODJrNd5C1DVCvnc/Ff7JRvrayrsXIFJep/8PvbXJ9tiTC0WTgLcMA
jb5J53KzoM6hDegROo5ak2cXjscocGhR4KO1AhhOkz5QMrxEJLmAUD9392fCnb2WyuSDzMo2a+fE
ZR+i4m1Wvo82YVSo87qZxgp4GNiqaczDMhB+VdMEbsbivHDVgWqvnpZcBIprq7gNuByUmgnEEsKu
guLLdfI4JnGfO5mr1gCT9fn7u+/xDiqAdJpPw2F4Zk3h7ubgG6UP9MvSfT7BtwdVqCPGAnQze+N+
IWzM7IxerP9WtwAAHBsWWOmw4r/3pkxPgXxFp21taEZKhVwX24LiEbo7D2T0/enkBG63/c2cJFIu
WFXMsWonz9oX/tWxeHqsZQKuugsQR3qY5Jk7kCaabfr1yV5E7UjJRH77dTNptQhAWqZY4S77lgo2
xaPniamciHiMMcf+pL6X9ASp/O3Ofj8XCvonHPwbMgKeAm6IK+dpYbBuKu5GNgEEk2/Lkkb70uuG
K2O67UWxorKOgfqycgfdTu0SsiZd/XTl1WwdWdZZP2PuETAxkkH7fJwWdgNWV3st9wZLVZBWgVkD
kCK+/2kD76Utl+kxbZUO8cnL75ggvYvE3hTCGv2S9O+Ci9Z9S55/Jd3AADdip2HXMIfnsmt2X566
N8vcaK3BeOrKX9baZw548VfiDq+RJcYCHgx75pKfJqwbjjD8On/rga8Pd1S2KdlcxXWTFWlAdHjf
hpxO6dFksYJtmGBK2HIAJg3jUaez4zDBEZ8xCqZfxmIX5VUHAHtVS9mIuvKXvTGn4msUeUuYqQut
UrtIGufhIZM+szFyaCchXlviCg+JcVnnhSLrUa8U0V+TOV0eKPRsZ0k3oArsu392BLcxMmTKA409
+5S97RIDVUUO357xm4tD48LeDleuaOnNBI41tZK645+GQFncPSV+Em2Wk1yqOtHuer3QwkjP4zUu
c4Hxzdfu17FH5o2WxBJqwA5gXQeXWc2gcWDlxN2EfqD3UJZrP7HdHoqgYrYdC0/OZs8J7Hd2mWjA
n29bxWBbpZ5V138Ar+rKzhW4+OnmdcDjKA8i43VNADGvda9eiIcvmzVpzewar++vwlSHM4qwXHjX
r7KSmopFdEUUciwaKGh/jxPrCekADKtQCT9sCBjKeH2KF3D5Rlr/AFo3wIdfpjHVphgsSO3I42Et
/bB3v/hjPBFdIIGfWZGUJMpb+NVhB4XAsquxPWz19liY0GZ/HiJepDl9eKa6N0x04QeTcWr+p29k
BFQ9YLIpYwB3mhpsUfS/kwL7lBlunB3RXfQLOVslqqHQNh2PFbeljqmTv+S9eKtdFxZmcIAtuSub
FL22ACD0CoGH7kuIUPzFZGiNdBQ4BELBPogX8r8cnVRapO7oaER9sCc/UO+ClB4ugl23gDnZmxwE
vMBf4R4g83OBwseMPdbiDjHfk+meH30wwaaQqYpugDZ8576koZe9EhzCOHKk9O4Zx/iHDPXtqY8U
xdvKClIyOLRid2hyngocoRKZGo5uJga02bXgchEKk7s1OMVZwnkxBHUMbESATMxEFpXJXNJu2c7Y
aHZ9kTCYFWwWBtnh2eR6n8CdXxskXJiqpXM36fTCdMA1lvXzGOLNnGRtDrT/p6s0j2/ymysx/CE8
W9p69sYtyOLxKfecVs3QGADMuXdanWk3ij+wA8sdz0J/Oeaw7xmAxjEvPa38pfuf9ThcHkvPC84k
WL/E337bITbUhES5mEup29/p8w9IWc+L0GHw6sHyoL1ZFTHKqxW1LTus7DGCg4YJCsbr9Kghk+M6
bJuutc4J1HREqjIv3lUhkbJylVl7gqFkVf/IO82MCM2gATrvJ+2AURuOry7S4PigY3f9YZIQuvL6
HGfzgtuQVF27W5lK1w6lvK3YKtlrUhsO6PR1lWmDQ8PcK0pqRBZnHbAHZBM3ghuYBpsHsU3NI7mR
Y6aWfCVGRB8qVbiNsduCEggdCWpV4Twh5bJsD8MT/ppYkf62q8+M9Pvtuypd/HePs5BBsXhQOedM
QzsFO7FYGONpW3623E+xIavIhOi22fgKF263aS8Gn0fqQB0A570mJReYZfVALpn0aAUuPMqxGNQe
PqOyqxosNumgwK6UC4eNJDjttKmBTrG1K3RS3wToA1r9SY9NfJ6iKL6ohUSOTzFWXPEwCiyUr1gl
Yk68YxwR0dk+0qTaMg8hfeCeGRYdq0eZJFa50118t4oK2hnJAz+EM1vlJiYTUTOtxpVIMJG/s+Gq
WgazaCtCj5Jw57n5IcqcXn0E+1uRT+bEsupEIMNtSydrOSse4bBaG41yhc+zhX/emKZtLKpWiiei
Ib3hCiyS5eZsCBQTUa/ldhEqVFeZDZK4kICxAKfjtj/GjbaX4V7OtwXnR+HO3ZL/ZSguQiE90IHU
Oy82Eom99ezaduSAcsCA4YZOlIeWI1FiM+offh3MwsCWOLZcdZTyHAtzwZ/KmvXnCo2wznEdOlUS
70axc2/zQsma1rs4yfvBumLC05Uwr6JYyr6WWPXwzykCkVU7tmTt1mlGWQrxZZoIS5dvm12KyunC
sf8yqaD1UOvdcKrY4nqMBnouT5kBkTyiHlCM0LFYK+wnKE4x8SJ8dQm6kNeZvp2KOE3o0MSgwJ/I
VLQCeskWtq2nhFIbzxQSwnu7O54XdKlO8G33vT3tIhJuo0lV9d+7ugdNR65ey5tW+FelEJysUY9l
g/wCG1ULI+/GEkGyhwZEfcdkQ46YGtQm+u+vblK+2P1D+nwWMSH4i+3wXkgiXh5dgJn+Mp6PNrQv
iVP+SCTBhooWGXM/3YcfYOOyvTLEceNzwD4p6HrBMIoLF8hFzwYNl0O4MYICSf2G2/LZThM/EPdR
aQUGvcnbrs0fbgfLIcdQYlmcwZSns7T7O0rG70pj7TiJQW3shNBjwPIe3sWrSR3JU1jDqdEwrtIr
bdUgjJR3j+xSjgi7LZIn4j1ThmDKyOIIT8vi7Z9ik8vP4tff6budU8O9v3ZFf3qx3/jIihcLjnsv
sgkuekO4Rjg5tlVaUBWr2tpoduniCuRx57VcIT69B/h4Nv+oGKCNqgHi6UAJ9iUgqhznH2FoREXH
kl4vlTVPIUqKtdupzJSkN68OQKuWK5+B3hc5bEU8+jw7wWrHE9bqAI4oX5Dd2CvzXLvVHRe463OT
uus9ew1v9n6Y81y0lEp2qGc1CGWE47ZXthFicCMwQfrvNNuKaNMCDcW0XdYaulYwxYsPUauDsq35
8y9iMCnu13+/bysxDD/w1c+YCy865TLUL96dY5OCuvN/lWTBvkHFjn2HIBF5MNnZre1MPhL9Fojj
PZHa2exIwHm5G+VCggq6dsPV0deqoGBsdLd82GDyCfZzmKEBRBeN43fVXoSITi0VfB33RFA3+4Oa
cHgLOPzHhIAH0oM8Bp652ahzcvFX2eB6zBg0mPnxTegry6A2riz3PYejiSZQIQ6u7PcDp0tf3qdd
ckC4o8ACJXlXjeig1AQ69rI2M1Varzg+DXVAsOYldluukMHHjL1BJFMSDn2ilyDMXEGBugnjSUVc
tmxUbztir67nCelqVCPVNmaraY6/XH3hTvhhGUrxssyibADbU/vk4Hm0H6PXNX04kbmwy4ygbO2A
55dtgZRdAyUcgapozIhuZ4ydLIgwqkA8/n1PKkDAT+1JXIz5g2okm7+qU4BguXPjZEnL6Ya88TXj
kNXQBL2mQw41hvfSi1RxvMEx+fEK8e3eFHD7Ttomd1/qcQA8IG+u78YhCgkAus1wb5Yxu5xXEa4+
LZdRycqe750EZgEEnRNvnZDSI2yG663NFxXT+y4bUnhuqMfwWlLKa/oiGXT3HHqzsRO1DUifD0AE
JVWXTXr3lePDtdH5o4AqfHHay9PntM2Ym5Z/MXdNZ/giD/MhMm8/uaIK5ilE5q1PUT4gnewtB0/l
RQ6bGfQG0eofJLgerxV0eE/m3iR5DS4aCbfWx17oJBDReUgD5PUap1i6vMoKNo4caQ9FmQ1cwyDI
Xvr5Xdo088C0MLwcVr0cYA4OUDeOhz0Eqe0qVCO72b+z0+Di9xVUGdtK9JqDXcYL4OXcTSXqen6P
Aah5RMr0m+63Rb1eMfZ5WhQ2Urpq4GPernrFbbUY4P7kd/G5klrBcw87Ljyfra3ThuRphlwqbqkt
INubYYXB0bbvOlrR7DA/o3q9I6gg6P+IQlAKHLOL99J9yXHpXx1u/mmYgKXeVjynQdzljBoo6hWi
PCvnhkkQtDnD8TZcrhqxTszmvvnkTSK1kLwYotge9y5Uk/b7ThMpxTMnzKM9bN4ClGBGb4Jb0h88
GVUGNbBbO+OeYEl0SyTkZa7E/XXyj/I146ZfJsRtNV5/LpsweybIAq3qLC39J1pQMcJeduT5c72c
6qeJCen4jCV9Yw7c9znwpqdlMOcOPQgq9o+7VVpu60N1GQwR3PF5k2l8tqrU8cP/ngWA18Kwfjjz
MffFIhDCiv50paVmPS8XnUrk6kVS+atabS5v5e0PnzZCM/jj0GYP3QxFWSmI9xuLCIn397Dz0zvA
WjnuqqagnWrbKvDRU5T3a+7vCqhCUvJn3ON/P8DTbNUQyuS8vKxreU+tl2yJcJOZH7j+tf9jcjVg
pW/dZGr5bxWnIRP3W3ttFP7XS9ks6KpBfvEzsyuMmoPC0xbyGgBrLFZeQ7mf3wXxRG+VAR2wpKeL
5B1Y6apJ8h3rY1RBczdELC5ecGLILfeF4Aoo8rVtKT3aTNXGe3yMDPnPoXMJbRn88rcvrYWklZ+e
KzR7RT5FYn+CQ1zvqZpKBbh8d3r43SmX1Z8p/v0uvUrSgKQ+Kcaz81AwoJaHKR8yy03M4v7FkAQS
TyLg3uHOaJnXye4bPKUVf9gmh771uOrYrlJzYgIE0r1KOAdO3a895BlKKGsi4/G1glxdZYjA2vf6
gGqFhU0joQn4HCbg0JcAYn/ywJ2IIaXQLn/2dUMbqBSXYtEtpvAJCsmwN5xqLNpccR6z5/tuH5XO
MjN2y0MvHdcD6mIJq06pbJ+5dHFWU8NDPH89C/6E+ATAxQ9yUuVRrMTNfQSN/yHOPr/QuZ1w3gSj
plHQllPRev5B964kwpLFm3OOugL5swwEdvMCX3iG+TcHto7xXKisq8zjBr783DfRPGR9XKwtabu1
E1RZv1DWqcGjLv+XTw0ifxfdavaE/QhAAjB6Kc9Bfm2cCK5SQXw6O/aF3jPFwnVab6vCA7N/8hWQ
JNsvqKQSWw8W/n6EZaAap96/ok8vgx11a1SmMmWvflv2U6Fsgb1vmgzrmMb1iaQHrMI/YGODyDvQ
jpNXIaTabolfrioFMNuROX2GpV6WRP2MCQorgmnizzVtYnxxnL1Gi0dGSqtDbPcglS8NevntFl+U
5oEQZHA21nxKwc8jmu3kW5/9d41xkGfR0aSzQDW7JI/quQR9kI8ggTI0wPx2TEfOOKlvTGxce1A8
NlqCGPfKPT9KdqK9r+FfifZmYCOVw4Q02tQlssmSCFwNoIzw1GBZi1cjkFhBS4cpUPnbH6KePBUP
/Pj2IS/HKzO5u4/9BL6OtDUpqbt7dWCOd7Zdud4i7GfmJgQU3C6OhWJip+gWpV+NjlhOXFqM+NZj
Jq3/foF7SG+SKEAcnE9RxLeyPpz94qm3FnGBdATZhrG5Plsqt2OD49WNSGzkhhDToVaQ8fFxNLGg
XK0xaVIMqLNARRL4e6b7WNgLMR6rajs/WOpwGKAfzhXojno/N6Rc4YDusLwvvVr4/YZabczQbn8t
E9BKw/nZ8xr2rZ8vy385Ge3Fy2+u4dfAjTZW3QrhkMvAux+VqDmBWN4rOpEydODEHwScPV7SL386
8Dn0D39zp8D5P49t97euBBZPixhZ8o8BEt/QtvAti3FucMnnpJReWdjaFWlMN09lYY83XMPv/T+c
njkjCgAEtIUjz52vz0nU3g17A+zIuukaXuh+4T6cVb38Knvhq9Xv0uDseJrguyMz3qKM9089m5YA
vMk13C2L0GoBW0DO7PY/yBqEFNXWYv832mv5QB4X9/f06Wbc7TnTcwbOJI84P2jojxtf6IM/Dgy0
T1abAnVU0UW8LPyAS7Q6juD8ETZZrZV+s+6OtMYi7USOiqloCZGMvxDJ2ZBc+DAlcaCka2x466br
vT0byWqfPRjwx4ZZx6Fx0uoPFE100JWeybo9dlV3Uuu3Tpy7PiztUnRXapI/UlvwOyG4QhXpoqDW
QMj4VJMTPBd1uQyMxHimWWnHYFyC1RgWQRqy6oqqcazX9R5sxJJhOO7BlqlHuVFQzRDW5kS4rR4M
b3bbV/5h+Yi8d1DU+rqEcQtE1PgO1TRV0Up2nKrv4xZx3rji7EW3OpziiV38HPf6aZw0l6fns18O
Ym4f+/UOIZqV3B2fixkkbHsqbEGQv/Yu6wfYQXbMyJHKXrrI7fMvxzVhEColirhXXO2ZAs7DckU7
0CvUQyxEHVc3g74h0fumJkbcHpFd7Np2PSBO6n5P7NlQ6RIswMwQRUslitcqlqeCiP1QwIuCtg6b
eHs26/klA4bWViLmspxUDxcYpxQR8SdsycMBDxLQyW1AfZIL5TOAdg5Gq5So7IZjBWT8+zgPUPX6
62R4Y6nWlzcfnBasLKxmJ+a57fcNDdAuPzydNJCryFD8hufejjUcZc6UnnphrtdnP2JnWwRcHhXy
mlhV0cc3VcZmXfsUALuv0WD4nvaPo2bxxwKnLsZQJMfav7XUzUoPXMeUagzuyxuFl0pZ89ITsZcw
NXgAxL/rZY/C5cSBHiftO1Tjo4ca37crFsJnJYVLLp98aHqMw2dDgOZrbQKfgVN9n+9sbqfjvr5Y
OdUNbrzt2Pthe/n5kjnhGgu+Owxhe1SxRe2TLjkKLae7bZBgj0uratIeGg5v5JeRFAgEKax8ygPe
CBnjBj0B/BCHxq2wwBZACVzW8329gAhW+MzouD+UhyDpXLwm/HtFSVy7YdqM/gFRORpCv43ygzII
8szmnEdgqTdgVVGVCKOMDYwyqL11xGiMvgGS8K8t5URMMw+RNo9GND4G1Hg4gYwDCAoMFBZPM9Qz
SqRc4fVuf42XS8hUBhiiqpGkTqnVslCT/NwDrNkvObZ3K1ah/Byuj3fF+3volZHWi8Thb21h75ZK
gXt9eaY+MewanrWF/T4oaJRfxlmqXYtJRLcxqGW0vqTYCg3noHG6yR1SYv3hycei0V7dEluLfP6b
fTxwqxbMegeo9ZOw+Q3s0XZ7JW9GLg1FgTvm6Oh7Mj2Xiu51OrijI6MjcTssTMPeA6nWlrlnEPJL
IfYVBCgl+Xuwum1uFsqbXGIUNAGsfWSpqag+4t/+1RfvGEqAdeRZYizmWOUsTL24wZdFZlravMo7
SfHp5oLO44rxnG0lEV9sMdnmdBcPspXmVHWrDWh1ufy63LDsqI9TkifIDKKPEFuPC2Fjmc6CcEB7
ASGkXNCkQybUo4McKPSOGgTdYUGom5ikgzUd0a7/akAX2tanvAnocUGXIFhD+HqTW3ld9Kd9SsgG
sa/4qUI+FY8CSiX7C1eHbovpVCrc2qtLfU2hcjoq4eRNNVslasX4StUWIR5+Pfitpv6WIiwkvnQn
KC60bCuZg8H3UP1jZx+AodxpYGM99Sgvkc7JVPgXeJubTeC9BLfHpPsMcfE7hRJYr2PfVQ9LN2j8
ncu4gPZBaCc2+Y/4wfwzjTwYiba1vSm+rRmwVLcHIHep/lzMs+L0rrfavrgXZ0Kyws9S/oAJnZlA
aJd0oC6OBofU7H59/Fdg9Fi583nekpKPxNY5/XOInC/73GvlGtHcPhrTVgjCM3fN8maEL5lSs+tY
NEYT1UkfsXYhJtYXeIg9d20aGDrboSDBJr6EM63yMs23lGqtkMjuDFZc/yGtOb6azxl4uRGhtda0
uOI+Lie4MfdnAyNFs5qoJfBeZCdEMQR/OEo2iDeH6y0wWoTqIgzVzAXBxI48+S9AtUZ12aTKg5Qr
tSYHLmGIh+nMka+B+TPo4gLomkZI+Q+HDJd+fgoyFGMfWcwOWD0VfNQyyVyIw5G4hftyAxnmI3LA
jTG3uVMVBAVB5nJsS8iNWbqAz/0r0lG54341RBNcdS5R5/Bsf/Bpn2iyez4vTr07JVVbAD4E2hWb
odz00XFu6yCsueTtrAQnuyMDjUv3HKzJBn1a2JyfFIcSzXU0kyrMFTd1swA5Rp/FQGgwNPhjG/Wl
5LoOuiIP7v20FoD2oPGbfMijeBsdxsZjGW1F7sIXfC59gB9td5HhfQZgcH4knOCEG0rUdSzLZeNU
Mf9fmX0691IeBNzwO+sSDW9ciXbAHaib99R8lDVF0lql8LZZPcwc6sE+hhVHZP70kD3B57TWboE4
mCWx+EBDGwI0SnJYko9m/TYxZMkTtVJQGl7eF7NOLJkQxmv1+qtl3o8ceU1JZODOUxVxqWbxA4A0
opW+fAkW43abAhG4uuUZLPKk6hbjvT9HUfDgjBIPjog34BIOMUosdM1t9Nb17dcI14tKfUo0BX8s
Bs06XKOLAEkbkPbcSr+bIPkBjmkFRg7P+MBl+QvidMkFJ+ZGbBulN9wcidwuashYmNwsPcXIFEpy
YQ43Mj2tKekpU3lqnSL4QW58vYxDflEYUw9zRCdUMyKCRYeKjM6zq9SLLiQ5/Fmf40Leyuq0Lt/f
Y/TojIWhFY+ojJDhO2DlTyessp3q99e8xNG/B9LTtVVl9BsYKvjsukznBV1f/+2wW/nd8zbve8Zj
gWS0/iGAIRjWT3apdeT8JvtNZYaZCTU2nmC2DWCYhg2JnnrkzxY6tk8s305H0nLUGKwje4sUrYPK
K98qtxE6QfaaNJBKX0g3C8t6W0FKTSayC++1P4P0ADQ55T0j7mAXuEunfxe+uGYJQY16bjyj0ept
3ss4LUZPUWwB/WGC4gjRtJKaCodq9fmQeRwHcY/PhNnemOnnjumNl//f3pDQHQ1AoIhZFLBYb3Xz
jZsb6Qo2wkKTz134lbpvVK1hK32PlE8t8OYJbgZPQc05+A+LH9feW2rc9kmwmTdXOSmhJUKbbkPm
bwPIWRVweG6WEOJIIRWtCwHbo/YUG6huGu/jYilxjVHkxPeF5A9bECfQN5yo4K79makIx4i223My
k4sW+CZmo8N+qPqctE89irKKDpOqldflDlvwha2u1GBHBlAP5ALQZCmWnbeYfct7mEjKZKvx83hW
A05+iCI6YXed53lzRbaydK67jMs0ofcCoTaCnT0aaOMwY7NKZXdfhJonju8JJELZmB7qLYuLLJaL
sApTVM9RJc0vvDZBm6m0yPHaPHTZNfZX7/BlBfo8ZNa0uFmDyx+p/SVegKqZZBi8oBDHMiySNuBZ
aMgbEztJW0Pk6Z0iJRJuQnVJ0bkXRqfKIwuqfV/4qgT7mo+kJ9SK6456UKC0gmwtDYKgUZPn69Dv
75RlhDL43EcoeILiB6gRxc38y9kOHR8qOc7OenTXmhqIJUdz+x3FEtbP66WdG+ORWWP/gjhtmzZX
ZWX5KdvrI19cd22RqjFToG2FdquxEEyCpwdOkp8Kvc6boq0QowLy3DPRgfQE4FmC4Ap/MWHXRhfP
iSFBMApDuXUxY0UKOqynEfZhlt/xCAipv5V3h6SPOvG0gp0GjJH5G6yD42+1JXP8udOcUKUmevqT
Aqr+3qxxjeivx6dzAruxyMvTPiGgZ+oCMIK277IdYM7YvXxxr2qLy1EqCdrVRxekzB1U2wI/FjCS
/vW1snxpfBjCKv63IAfrNE2kuib0EveewP8DX55I000Of9N7XrU62JbRLhtNZTKEfbuYjFanW99G
MgdG7Sis0olZEaEP7JuM4AMnnCWMKp+1+g7Vt+AzekkV+cXqVbIbPUgipB7seny6j9WA0H3uuFZy
d+W1/rjzup+hGasRqXOpLq2SuSYoWZMIir916rBzgDmm4VvCwxm5HdiaIhNf81qTCvJ+qidT+15i
EOi6xJyNIXX69buYWbI2OHgWR/aTVQ54FJ6AJM1yNt/238VOX402myxOZadRWhsiUnQvKj2S4HiB
w+c4N+afpug4ih8Bz/Tb3ciWyaAHd/i5DSZDc0FAIz3YZe3kJrqYSQ7UVQtiGbTJMOfVvjmBX5yq
Jmc+TCpd8RWJX6oZn6J11ryuWWJ1gYMaoFKWA+oSoKT0r3uJLIFc90TFK/dG0hyO0BZV55kvdTu3
W+xNUhtexVDinPR0QM3Wzhayc0KkdLgSJ63hMR5GlMIPTMbGzGACTYJfGMewH4o9Y5JGXkUM1gjq
soVaE88pbHJbI6sanhmgmySCiCF92mX6IkjfffH5atYGN0R2NNqRB/u1o/98BddmxTCXAAdCeqlj
XCSpl1/REu3sSvhZJPid1PITOn8ANAAfS3jkQIGuRd/aVrZORBkISwFmzrqMIxJygyINOPd4C4V7
y1JpVm5FuxG+8foCMOAe+wx5hRiFisUhsp9V//s1YvCfrsys7l+VyGwEo9ieAYaX7+syqxYt9cma
fzyOcLeXLOFYfWHCmzIOkMP7QVU+usA7o59S6RCOV2C8axlf0SJs2yuSCYZfpa7RFyqqFx/XIdBQ
eavxrrxd8TX+Kjd72OKG262gDV+oLucdxVGjrjqn9cxBSi/C4exuESouoaX0qLkRH0iThvIQD36g
3t/+/Nz6FjDLhx1gFPWD0I7/omUGvgl0bWei4dyJNPdL7JWmVSDhpr0oJgag2yV4h6N8gpGktyXj
0GnUuMaOthdX395jOi1U72XKE7/xq+EkswGzdWD9P+J5bmb3mCRYUozM/QhP8f6jzZX7DcgyTA/6
P4SZreIjwh8AP98azou5LKAWuH3aJBYC0rTEw2Cyo1wnZqrzmW/A1Zh8y0qQXis/A8HaNCeJY9Ml
tPQaMFmnh35/G+xOYU4hNlCmn7iL0mqmyoh03rx8jfT6aq62bVPjxtOcrUq351jb8/fGhc/3QvoW
lFXKCboXUBTKjLeGmKJDfetxHvtyWt8KniP81WxMEpi6PSecyWTxgnBkt8NPWLENDhAc6Mu0FjFA
HR9RzdwyjfLhsLBNRQdSZjAkdrzngnY1pXSyKFKfiSD5itrtptS9OutQEa+CFwml5UIV16uWIb5O
XjxcyBbKmx+kYmgoor2zxZkaTOnMKkHVvU3C+1dLfQlwKZDjGG3ESeP5/XwiIglMI4KBob6q45uD
ESo+8+KkbfwAWlP62CYupuVyGbzOxKqPLdi7P3VUlFK+ueqNelDOkP9pOCr4ZeH+/gbjFnGpoTJ1
e408p7TqOJOa/inOybVQa5wN6LR06pRvH/ju94fa7lTk3jVejonsUIdjgYg5Ja3vwHcwQMlguf6n
lVmIOA3DLEbaGuspxQ/XdlJ7HiaNvTACegKBf+Ga8MCD/iEO2w+oqwtHXrTvZeXIg9YcqoFNij3A
dzaVWOv4MW59Dx8jqwSRnRV4XovCrWvpSm+FIIOXpDtpNTqByZrfR2MLsFvXtGGjByQQVDTotnRG
L7QtNwaZ8ZdFYPwfJJ3KqcLPf8KBMNhjM+C/2uio+uCD5Qct1JWTW8/e0FwE37P1jZJ/Xv6FPW0c
6Ddyp/FsD9KMKhF4ls15CXvEduJS/HN+yTWLhgwvIb2KNe4lVvKNEe4YwYIl1IrmszaABYWKF2GP
MBA8kMuSCt+ZCubrgAPImX8ye9lRh7gH+i0yNSJbum9JcBUn3ua68qGKWXHRdtvpelIwQG7lvdwo
vgaX7htISSp8N6QY4QPshtqY7WaucQQSbsp6QzR816Ec4wCLiCSzGiYz4MhP4rB3NJfURyXE5DZ8
2fBwNx+honfuYrdoingCwgS5IYCb3IbkHVotVY0bkCT1/0xGT5wY0B6nXyaan5N0psOgUZMh+D81
va2iMeKXDo627KL3zEVrr5aXCBzoUJ/Nv5DI0CdS6hueof4ZQZWlfzFWxdflhGAurtt/UMd88+6F
AdBZLd2wTL5+49lGS1/vKt3YQP3ljhA4dhAv0wsBb59212SLMki+Ur/ZDl1aHtIId2ywHfasan2l
TqGWUOQfp/UCIn/PsYTDoR1kzLuRY9+NkiO198UJN0ZpvfeefhUuPtd64DMkzc4SDd1G4pob1N17
gpJhAVVDNvNZ6yt4lGWtFQGVPonjt50NtvxrVBDBBBwp3d0SsG1x0/ognH4p3f52g7ywEFWJXzZo
QqefsimKCMsDrmEKzprLOUOIF7zrwRNpeZIqi46BUsUaoSn1ArlDIvuw0Y+Dp4sM7xliiEj/Rze+
lB3ebFlLXTcabB2M3ddzoJypcLHj/GhfAHepCc8kvEdOO+JqiAXMFqcvuaM0QIoQk3ogCm7kVDaz
M6KhJctrtvytxqqx3Hg+Z9yU361B9ne/JYPvr51MK9fmowKUaS9O4eAcN2AuGwCioSHil4ucgFXE
LehX6PkzAHqTM73xVvJZKJlD1mo0kWmp+ppKxSQArISj/Qa0CtfBjjbM1okamJGEBxDuoL7awdM6
e8PsiXrzjKKY8XFwoEzH2Y6MSfgxuK7mSwqFTPTgwypdHTpRCsTlSSuyIAQgBis0xMVDtX28j66V
MkQes+0YvYEN1ZdbjK6UF4wF1ogObj8j8ioFgsAldmD07znFKVkTo46KCieD61lPo7xWzc2OIAzj
zrIQNgSBjRvynKAnbfhe6jG/4PC258lVNo6As2YMlXto+mpoU7uIlmsWwLMwZuhlMb3eLkla+/KJ
WF1g+pOqJ8CO/0tb15wQ1woWhLU1v29JphAADk7QeoBJs1zw5ZzIfCghVPh60JbjwMS4HbZv6eVB
q/+wEDAJYaD1jjvTubBqbgTjZ3wf2cyI6S3WtCkUGEGWs/hXAsofOsjLutm/a9L6yz1i7uTttTuO
aoGmyidsi5pIuWhDGBGfL+WFnEQfoO63uj/tjjjDZ4V9gJ339HXu+L7S2XEfcV1lVontN/bUWzXT
r7ptsv6AYZhgGyeN8qCtwhSmrkIyQyldkjBpoF6FVy8p9jRepVA2BiFEdQ==
`protect end_protected
