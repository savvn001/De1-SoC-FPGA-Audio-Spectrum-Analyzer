��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Ylr�0q(��mIB��� s]�}�I�`�/��$%��
�d����A"���7��Q�?Z�	<���V|Na,��<V�1\��Q�����:��
%����(Wu��lv%,����ڧb����z���� �ULoZ��>�IL��u3S�q��LWmL�X�Q|_����=�~���SЧ�(�)l!����;�7~,'��qC�WM�ߘ��gGg�$����+��g�9�=>S�IjJ�gR���`gq�Rq+���7"TTŲ��ŁM��-ӿ��]W�h)]�0�6MN�O�x�+�i#t(�M�%qގl.��:��s��ےM�S�c只RK��FWG�˗ ��8���g�E���u�w�n7g��%�|jܫ�7�;���eHr%|���c��d�cg�C�Hr��~���D�V@��W���Jkv���tL�sC��T"��$"�{�z�� 't�����o�q����EbRY[�x�P���ᡙ]qu��X��k�������0S�%(�b�v�5Ka'P�hA��K�K�[����c����zH��I��1��۳yQr��5�:%�o�0K���֚��)B���x�͸�=<!���n�"���m�u��t�v�ޣ<R'
��N�-�\~F�ɭ�%��x��J�|��UZN;����{�D\�!��W�y�@iU��phB��#:�
�:E��<�T䙷�+~��R�B�a��p�Iqx�a�-5��=h	#��h�)����ͥ����69q�,�{Xm���o�Pom�c���_[�C�]=@7j���+�a&a��8r���B,��#Է�hT�@k8T�rGg�z�[�X0�""6l�I���!q��m	�޵�Q��7�Vw`��'p㙯���S_M�G�"I2C�c$�<��M=띎[�: �RgF��2#iS��-�%<�h��0v��ukQ<� ��U�u��q�����Dӿ�0>m:ے��\9�[0:r�_��u�c<�,�e�d���|V̨&��ң$c6�?����|2��s�����SѲϠ�:��(�RzH7�i��� �-��BGV���MWh��y&ky�.�
0��2��ȂS݃�0�ח������Q*!�W0p�g[>�����e*�O��G��ŋކ���Wr��S��#C~�DQ�i�KC��N	[�ºk���W�Y?��W�f�׉���3:2���5ѺJ4jЭ����2$n�ʤ��ޛ�&����f�r����sݩ�d��t���ҋ]�@�F��F�,�
8�@�@�_��H���P����aݓe��V�\�>l>踯����^#�9%/����ZۀڦF��q8�F�D�����g@8�ܚ�oɏD�9L�i�1��-ץx-���p�W��O����N�ei�u	�?����9*��K&����FWH��b��( a}�Ku�wx ]����~���y�D�������t#��%�����9�:W���.c�Hқ�L�cϰU�=�w�6<�
��#�%\ i���v��I���wn}�O4�Q�$-�����b� SZ=��I5�(�b�O�>�V�}y䘑�R��݃�>ݗ��C��";"tю�LjI�͊��g�y8���V�CO�
���!E{�8*v fv����6$�hM�ZvT��#ʾ�b�*�0hvm�O�3�Zy�|p�J0���r��᛿�F� ��)���%��Tc��ia��;a&�f�H������ѱ?�ό�vE�bX֬i�|^��ոU�㍚ƪ����lV���1\캷g� 7�2'�P2���
�F�Dϴj`�U�RAe�%"����B�ٱgKL�>�����v͜Z`��!��R(W0jE��]D1�+G[��|]�}�fV�W�����&�?��|��"�N^o�1(�C����	B���nS,�ظw��ˆ��>�ú�F�:�����Q Tn�7P2E(a���W���n���"�Ix�q~Au4r޻|�k���<��C��v�:ǔt�Ą��p�{m6ۿ��ulߛ`9��E9�� !|ln�t�8b�Ǥ�T#��8�~J�iV�ݯ���4�?��%b���q$9�x� ._h�r�b2�w�oj���}����5�\��	h�r��탥��~����x�I��QcPϩ,o�G5%��������8zO�k]2�l����L��Sd]�|�4=��j*�S-��"��� �ZP������n?0��
g�,"��OUr�vo���V����ew�۾uw��̕�JY�Z�1�ɥ�9}{�?��p)�DW���`�+���љ;\	n�4@&H�	�(B������*�i��!z��h�ܦK�>��c�Y0P%�[Ǯ�!�.�B�(ϋ"^P���I��!0�hy�����&d��%�4���"���c��{�j�Z�A�P�Q%�C�<�
���9��c�MJ�	���XU�_c�Z�:��*�>&�~��8t��K�Bq:j�yTl�E<n�X^�����E�z%j��@Ef#2�P	�df��3�CwE�m�#���Oa�L������(��y.�*�/���aF{
�<��ɮ6z� �1��E팡���E ތ��a�8�FfV��!�G¥�pEO�M=�?�)�˴0e�`�x�CY��ne�BeU�ts�q8����iP����Z�*(M��p��;��=}��t%�鸬ޡ��k���:Ņ��l�9Υq�ic;Y�<v�bIC�TG*�·__�8�`�lM׹,BX�l?�6�#�IZ՝�!k���-�����V<��b�����;��V1U6�������"�\�J\�&J�0��|��p�{�ul`��_�i�>}%Y�`����N�	�Nγ��+�/�tGƓ���V��繅'yDl���-�{/B�x���N�@L�!-��mR�����>joЩ�S�$��'����K��5uֺ�ID/!.� c�]<'�v�\����V,w� /�uw,�"D�r%����@K�q���?7���iD}�4�g'�~<�͎�A��3	v�^��{ܨ��vJ�K��̝�gd/���:��:�[����=���7��˯��-ܷO�wl���8< RG;���T��r��6�/k���Рo�8i/٥���gdʆ�d�Ƥp�D4|��l��qbѰb�99�B�g<O�~ࡩ�Q{�I� D1���@����Pr�-s��ugw~E벹 YF3�D�u	��A.3z��s�Y�"lQe
�8�����~$��`�������9h���J]��S�"���	�I�Uz��G��cu�w�t���$ ����vؔ�W�5�U}��r'9/������J1��C~L)4zUO^~9�D�k� ���Hv#2�#)��j��[zP�Oe�U��@$�Z���Ķb$�r	v>:weO�3Zd����j�[k+=���c�C��]n��?D�4!��Qh�S��d	���5�E��	���@�X���Ф�e�s��������{}i.]B�
L�I���[�K��qv	>�5���F�|.�Cd�����M�`
�<�g2+{�a8����/�2�봭�����#CőF��8���
�-R�4�����D��d�"L��'���r�n߳�t����ޠ_j�9�W�Gn鉒���O�;�k�ɔ݋O���&�O,�� �{8'0B�;�ؽ�2,��q� �1������n_ÍE����?%��VO�{ǧ��NѮ�4An@0�I1t"E^L�T"!���b98M��v���%"R���P*�s"Q|I��ى��Ua~
��y4� !�N�d-U�+<�d�F$m�k�l��H0�nYJ�<�`uQZo{�l�p��3�u���3FA��qqHmZb�q \e�?�"dz?�R�H�m�F���QH+w8��F/�bI�	�.��?jߤƇ7��r�D �@�}�D,��I�T���3@rOS��{�zl��EOϵӛ8���ilN��e'�Q;�}����f�,��L��HG2Q�<m�C�F�2i����,���ךd\f)���3���/��M��m0A��sm��f����<�XK9U^�5 EX�F��4��"ʻȧ NQ]�)��?E����~�hX�н_����0��~ �ۭ̆���7�qtyhA�&�^t��o~���&dTD_�	LU%��y��W�z�w^�&8&��^�cL|#��5�q�8�'��^�4n�/W�{���Pm?հ�B����|�I�[�E��������
.f���7K|�B�Ԥ�|qƉ/K�n��ݓ�@����*r�5� |�<���Y<t�6h
��MJ��EcCw'�7:UԻT-��
d��P�W09�,]Uܬ�U�EPT�?�e��ܔ���i<	O�u��
7������#y�6�=v�R���j�*\��Qj�4"n�ţm�:iUf�H������;�:������[[��7���eu:b�tȨ�C����X�`��d���%�D��������b�*�����('��x�SO��Tï�:H������)���T��Sl��[��DǖF��}/4e3t�'&{��Tc�sNI��H�]��X��G�z$��Ip��߼[�RnH�����6�bC�B�����S�qٔ<�r��h�gҢؐ��T���x\�o �
Sm�$�+Y	p����(�{���N��p�mU�-�����^��lT���1�wm���@�6�4o�Y��e����M� ;~���U��ɻS�5K�M�VZ��g:[ ���o��r^@�,�R�ņl�Y�r)��ىHN�%k�¾B�A{ݡ�
,� [[�,n��N|��y�,���![�*���� Z3C'��X���P�8;C�/��k!����iھ�	q��3�pr$�f	:��wJ�ɕ�W帉�t(T�h)@��q�>�y�|b�>`/w��a/�)� �?Tn˺0`ՏT�as#+L��" ; �F��2�cL��;�z}|����F��"�l=��#�͓j��`W���v�_��y��t��%k�Զ8؆�I��ă�x��uZ/���#��e�W�mn��-;n`98F��z_��������
��~�A//�HZt�F������p���M%뉧��l%�]#*���.�ZW��8J��9��jq�8N��Gd���7ğcXP���D���?!��@����y���E�:�$-���c�t�[v�S>M&R,��c�,r<˺'1�����[J�f���ii��w.�f�iL��6��,)A��dF�(�
�'F
�U��I�c��jh�t���(�ߌ쥩B��МC(�?o�|5�X��F��\0��|�F�)�Y��PnG��وR������#C(��ұ��z>"��u�(���eڼ���O/p5LI����X��3_�`�)���B�W��JBAt�_�x��/JE��ʋ8X�7�%����Z>;}����9����13����@c��?G��a�����}Ӆ�̸�`D7�g>)��3{Ғ0.s9���Հ*�4=�2GQ��YO�#䣶�[z���4l�����!��8�:���e��#��?Wg���%cpWJ�fE��g����S����늵k0����#Y3�s���wd�Q�&�%��>�����yɯ$���
���ba]�앩,��i�<��#��~�,��"��o���~ŗ<�5�_� Y��G�p�g���|w¾f̓m���U�1�Jh�d׮��'	v��JWp�������[���N߻��y��F����C����J�">~�Y��8��Wm����dx������s�;T�^�Q��]͊w,��M�mU�c#YsKpA ���G��V�<B�Fj��{����QP��/���D�+���_/��'�Z�/�C��_�������`�t���-GP��l�qf̰z���Z�Fq�G�d�M��Mry��weN�?�;S��u�����K�W��uf꿿5���\[Ӹ
�s������5礯����T�lI��#H!y�P 0��fU�����9,}pՁ۸X[Jr��J��O#mR��"��l�cI�:ۣ#�!����67k:��<�~և��(��i�����%?C���ͅs0 ���W��"G��2����)��#�Ƿb_g!m�8r.�j����S���4Nˌi��	�6��Q9�<yfY��8�dk�h����H���kC;��ݿ7���<�����~���M0�x��M�o��^����u��n)��Z9��������5(n"g%.2��I\�݀�p��9���rg;^d�4�����G��^X�]��� �/�A���J]��n�u��aֳ]Y������_�5l��������Z��Jo�#0��	��y}�&̰-��cf����j���D��͒!�2��6��M��9�50Dm���c��Qص����&�N*=���z[uM�u^I
��G���e��!��9����A�^�Ԫes��%|��jF�PS��	�K�]Ɛ�jwS�BC�jh����(F��\�/*�XW�n@-Hz"���r�!B�~8&��a���^H��,mW;9���U�Y&�������^�C���/�"��(���+�q���m��M���?�
iO�4e�Ek$�gP��/uZ��7��)/�\��5�����b�N�*\�K��*t]Ӵ�?Q�	's�r�KG�V}G�X����f� �0�6���?];u���V�w�μ��B�Sշ���g�i~Cw�-�X� �UUu��6�2sPN���N��4d`3���M��C˾�ؤ+�\�Ȕ�|n�2F�f6K��3�Op�X������h��&�/Pi���2�.��n��TȐ�!@U��k�&��j%yO����r���8�� s+E������C[�tV��ƐC��/nt���Jt��o)0�
Nx ��1d��\b��uۼ�t�dJc�@Xn-��4PV�����CY�E��K��~^��_��%��D��+Ǯ:�<�:�����i�*�V�c�����&2��vӡ��QE5���M�A;+�
�{�jE���W��--��{ȓm�ɰ0�P����4Q��Όi�˶{���vI"�sM����өӭ>G��UX���vm��{�ٯ�y׫V�PfYY���6�1�v�1�?����R��:����!�^]����xE>V6P��$~������-��9;Z�&���M����v������g/$�{h��y$2S�Yb�[R�Bi�
�|��[�L=P1���gx!������!A�+��.�L/w��Ō�jPȻ��7�Y���&�t��qʝG�Q��'�~Y��u�k@ĎJ���OU���S]$A���S�����N�h�����U��8�.N.#++:_�U\�ZL �ȱ��h��yS�o_��)�^� 󛫘���E/Z��s+�y�:C����9���ǅ�u'�����sŁ��J�I�?��q��d�ճ�K�A,�焰~V/���[�T�S�5i�n���V!߳�4[_խK���-������Η{�6t3O���iB�$l�g� ���ACqWQ.��]��X"ⳳ�;���@>s��i�z.с?�ۓ�*���]Cm�5�3��y	�>����b��%Gv�hUvu���
OTƚ �cxt]>�軀=wQ�����Z��`�ד�Zu��/L����T��EDz^8�PT6�l�_��JP�zGP<�#&�K������*���DN��~S�]]� o"�[`�O��7S��9��?]�'�A����S�əagT�{?�S���0f�����j�A�sZ���(/��B{�J~�j�$Xf��	��v%�����H� �|R�{��11�2�����c�0�,Ŝ� ��2��1"������8��F"��]ejI���̑�.�� ���l!}w__��GK��+��?�ʞ섫=g(�M[�"��hmpqH�����1ټE����^=�֑��>�`��Nb� ��w��]�ޜ��vѯ� q��l�1v��-��y��
����[>��$qG�a鄠���̋�Cc@M�}u2��oL��ܯ�I
��E�V.����i���[�Y����A��~3z�W��*�����0�0�eC}A��"ߐ{h�e����� ������S ����m��\�۲M�^��X.�w�k_�;��p#٘�.�[���u*_?���ʛ��WA�D%-|�w�����u����,m�^���T��`X���
���`[)�Q�ի�n��I��>�L�c�������Z��U{,�4���]O�fe�8�����@�a�mC�A��u�i7.�k��v:M5�~�j�1�Lc[]�|ź����>Ȇn�:/(���rG�����(�E���+���GB��&�X�I� �sm&R$���%������Ռi�J�����[b-����M���l�y'CW�Ε0� C���Ti�qࣞ�z���`(g>��ô��Q X�]|�<����A�t����у ����7'Ww���#f����|�d�ъ���&�� ���,��J�''C�EE1��+}�#�Z!'�~��~L02۴�֏7��Fd�D�Qx��.V%�
:?����K���*�����\5G��2���:ܫ���g��\M��#�*i��2j�|k)M��3w�{����o�%q�6��wũ���j�-�"bL�j'��)ܣk�Hm
�]���lbp	͠�$oW�-�&�feLq>��C;H~�t���(�t���3�<�P�����+��t�L��y��d���1Z��{h<U4��!��j���N���G���v@ p!w?ĺ��4g��r���f��i~fQ�Fm./nɚ1kw�񽷈-O4_/�G7��so'�[��_Qh�?�������F�]��솛D/K�ppm#�`���-�ލ�r����Y�?=+�vK��o��>�k9��
�S��x�H��Ɲk���ɡ�R��z�%uj5�O_17���w�:G�}��R�W;=�zLN��@#X�3"�?��U)�gh�2.�:;�L\UF;����r���-Rx��f����Ujf,�q�K�
�7WFkq=q㕈���( "��|eX��aԻ�Z��s�X��� �Y7�>�;<Zͫ�|\�	��ӤdL038d���$l��]��@�G�;?*��>�v]�Q�&�Ǩ�t;"��/�O���W%�$גsh�Lߵ�z�d0t��?u������>��,7Ga	q*n룘(1�ӮG�F���5�/^ s��v���U��x2O�;����]k0�v)�$��P/��6�.d&F�já�z���v�ݫշ��s�E�?�&���j�ő�C�����_a���Ȍkf��}�'8�өt��,C���7��Ѫ��}R��~=�ؚ#��@B�۞N�7��T�7G���}bli��k����������uP~�����8~j�s$=E��{����3�&�U�̤PZU\Gɞ�-a+��Z�;T:u�7kO����e�5X鯧c���Xʳr>Ec�=B����R�� ���E%gU[����~���A��6��Q�DP�����Ni�˛�= ��j��x͚I�@���_�X����Q6�Fw��t �>���3�r3�Ji���i�q([���R�m�m�������d�b/Xy�Y�����܊�l�V���a�c$�Ϗ�;A���fb�w6y��9s�o5�
�&�o�X����J�W5�)@�JE�A����Pɮ-&H�|"�����U���O����}7vWI�?�T>iZ:k�*�I	�e8 <�����_;�o���}ƛM�8���Tl�Un����,g�$%�J
�S�dMГ�����L}���
��&6������j̼&���.7�,��ohH���+�Wc�5ǦC�[ߴL+����oM�ު�O�K|��nQ���t���ө�(��L�,�"E.X3]1A�.)��FdWL�D�,S"�p��}��.#�U9Ad_�9�t��"�"QrH�j���9?<�,��1p28N�8a�0 6�kc%�8�A�NIE���~����/��y���e���E͈II_�=�z��6�r9\)�_2S������D#�L�Q���/�NQ��+ɗ�)Q��@���C����M��&��H 5\/��IK� ��؄���!*l�,v�{����P<qT%�L$��<f�E]o���C��2��p��(�8\�0���3Ĥ��5��`�W�o+2����|1��Y�L] �n_���^��������ar%_��p1��ʖ�y�Ŕ�p���B�Aӣ^�N�3��/o��0�����D-�P@b�E���M`~�D2z9
��O��e�p����fݾNi�����P(�M���Ӎ��Y~v�r�VL�:Q1m�0�]6O���+�3d��s��seL�ga�bPᔚ���m�ݐ1���u����&�Ԯ1�T��Q��'�6^p���b�J9ll�hw�i+=�����F�I�k�e�껲/`�_�3�{��p���,Uզ��E�Q#�ŏ�<�*�-�ʥj�9�`�`"Gt�H�$�����Qom1EjPj[�� ��%��}cj�����x@�왤2���88�l�Ieu�4���/�yN��Ff�Ҁ ^�T�:�S��W�OH�3U.㽸�Ry�(���M4%���z��k��X���c+VB�����ou�f��VK�d����꾋����˝�(�]�[|m�z���䏥�% i_
ݫnd*��_�E�'b���TNd˷g�D�O2jVY��]1J�0>���HR_�M�zn�� �P]����b�p�RIgmU�z�s1�����$�\C�'�m{����]�9��l�������k\�@�<x�+h���A��k��l{GhYt5�/��F���X�=��@��QٖI8 w���6-�Ƙ��X��I	](���\�]�O'o�/�9[8/����`�t7 �: ��69	���JG�x��2������i5dl�c����r5���h����:�?�wǈ"7i�u�~�y�Uh���C_���6�D�wdjY�e�~�`�Ґ��00OP�r�sČӈ�*�o�a}[1X�L��������O��po�80�A�0����}��x9-�%(��.�+ �U����[�Z�Iw*�~j>�)�t�w6d��Dk1�����7~g��]|C��,��!�!8m�}������S-Xy=h2'.�PKR��Ql*/����V�4.Ӗ�,�&VM0�g*�����p��05Ń��?=�5	79w�Zx��W㍃~F��pj��H�ЅA����!�}� ��^�������}��4�"��
�<�a�	�a�����p�����Rp{�fx�,O�ëT.Oگ�5�g xQs�m8J/NNS��{V�Z���T�vX�~S}Y|�f=�����r��@Bq��u����?�۞�^�օC�ҁ��x�F濦JE��ݧ��t7��$� `����ޭ���\��}�mW�`Ra-��6����K�AD���h�9i��!�%mL���$\p�a�X���8��0��Q�� �^��E�T漘�X?c �]���������^��k��*0�fb7�Ҽ,K���B�CI�Oê�%����J!�GY��R�%�p8��tn��A6�-B���'�D�oEke\�O#Z�GP4b�e�����ޭ�����)C�r!��t�kmɻl�Oc�waל�=��`�q-����vDB3Mt�ir�����������G9�ti5��xv>?c� zZ��V�E���K9Ŕ��Xԉ�G�oI4G��L��Yi����������I�rsE�O���DP��S"�s��܎c7���z� ��M9��۫?{�)l�W򮁾��G�P�&����x9�FG�I)0@�'�
�I0��?��ƅ�ј\dK��n�v�gf��nҍ�`ˬ�wS^�vw����tN!������j��������6�����6Q��a_f�~���_�ە�x�죢S�"��Iƀ��7����>Oڠ��&SZ���>HC|������fq�Ϗ��g�os�p�?�ۢ-s3D�TN!���1��^݆��]'~0b;�-��4�ژ�*����%}L(�ǊpL����:Z���܂��Xd^�9;���㐝H����Q���0zS�E��z����&���&��8A?=(�I��?I�4���c#���S��Z�Ñ��Q:�8r��u�茢���}��q$� �p��4��4�a%���n�1�e���טp4;)�I�B&����y�Z>]�D4���\�m.����l���H!G>q&���K� 2k���#�Z���v�!�4�nC·Ml���"jߴt&��&��a�-י�*%��7��iV�����V����>��oC��q�܂bE�
�mU{� �֑Â�̾��{�+��S8��Ј�H@�\���*�!=�ܣH�g!7��2܈f��L����6��Z�+��Nc�v�1��B�`�������>�Z!���o�A1,�M�.�l7�A�60��b#YBh+��G�Hݡ�1���'��� \���>���B���)Ҵk)�G��$�	O�%딾"��y�Z�=
+x��;O�m�җ5�$P��;Г����M��Pǜ��[�L��ۂV�6