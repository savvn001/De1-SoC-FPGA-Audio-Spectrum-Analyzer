��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��YlO���
�'�wUّ��1K6�!%p��s8�l��������S��2-�%�OY"���Ȣ��6S�ty*`(���՛yԣZ���L�_��-+��#���p�r(�R��<z����4����R���ٞ�y�����>�
s[J�C�ɜ=F�����J��r�?�U�g���l�jl_t��Ys� ��.;E�P��b؃��V��âC�����P|�T��#��#0q�gl1�YQ���"ʓ�|�Z@����lJ��{��<��wE5|#^6�Ɲ��3���)M,aZ.�L	k�
����3o�.�1�eƱ������	���V�Ȉ^l?f4�d��#
���ZF5P���� J'.`�u���;���C�W�[��3��ʖ嫲Y�����*?L�'�V 	�/1#i����U�р�;���t��IT!tQ���M$,	�e,�׹���#��7/�AF�x%��P�=G����}khw>��g�Ѥ�3^L�����(���K�:ܾ�o�z7����6ڄ���/�k�]�[p���3��� 6�~��+�s�cv��a.ǻ�m[��t-�P!$�W�������.o��+�)���P1��M��(j�|��t� ~(_���@S�@�(��<�V��?n�C�L��0��9�łB�{���2��������:�ܵ[�(Mj�߻OG��"O{�v�ǧ�
O�Y(Zu�+��Oi6��إaO����Ճ?ÇF-���_=�6�G�"��ѭ�:�d�7o�E=�YE�� cg}��vF��п��'�0�a%{��#J�6�J�B����L*}�YT���&˰?yX���Tjxp.� ��<"�1AYp���oV�k��xO�T�|���	\��Y�֊��zC؍�}3J���;�հ<_�9	�+�ȍsV�x1�{�ԁě�T���~���^�Z��(u16x�L�+���q��WK2�$az�!a���m�.�&6W���'��X�L#͖�6R}���׾۲^6M�h9����Z#�s��b����\�d2>�)�������&:$&����s�gj�x���5,�YԈf_-okd�����p$��\�
t�{#��H���(�Q���e��w�?���ж�0���1"��kQ��[�����V�}��`�=>Jk���:Hc.`�\w+��ң�?ǁ��j4�g�Մ>p �[bh��i��ֱv����3�i��{'4��`8о&�!�tՐ�/n"�=���sq��ȥZ���R�Іʤ,�Q��v�F�L��<��<�Ro��A��.�(`,Bb%�='��t��&O�2ц@f���d��y�e��4K��夞�M;�����P�����ۣ�as��@|n.��*���B�ѓ�@ �,�sb�A�k��}߸�)��, �U�ۡ��W�l�#+���ʖ���;�D0O�΅A��k�^��*�[��<���g�ԗ��㮱�8�bB��χh�@,�y�ndx5=Y�<=uoD}�$b710VY�X���� ��(p�7��+�	-��K���ccoo ��H�B�w���n!h�G��G|�f�B[����Pp@�I���"�68g�@d ��A��X����D�^��K���ʪO��,��c3h���l�E��CP�X���!d��~�7}���F~ao���W�+������0����~Rv X覈k|�;!8AA@}ަIO�-!pQ�xV���{[A,�^쯕@`�b���w$ł�����u�h3NS~��Λ��]jk`��Ϗ�]��~ÕG�ﲕ&K�}^�;m�\k�Nn6�����nB=rl�!��'�睡 g.�M�g���F�@���&t\�9��*�sb���}o�aRT����С�Iӹ��BK$E��B"Rl�nI����+�Z1�dJ8�{�:���U8]*�nO/� U.	q)R6|3�!��[#h�Ƭ=a�	�c?����T��*}}����
e7 ��#�J δ���.�?2G�5�>@�{�� r��XA}����u��Y�~c5��{��(���!$?D�1�$�dt�RL`"2g�=��<mK���h*u�HP�]8Ģ+��߿b�E�bv� # ����d�����܁�D��[��>cNӮ���CX4)q�H�K�N�0�s8*a0V�H����!yi��nCo�����(�6ȉQA�[H����'��A�+'t�Xh���ٰv�����v�O>���9];���{�Jc��Ӣ8<��ӅO�"�Ў���Ǧ ��}%l(���U��4��AR��w9��//�Fc*��ò*�}�e76J��DJg*��[���*��S�;J{@)OIp�L�����e�?\є2�����ys::�E�<r��XQ�]�#��*�!�gc'�p���v�i5:��}^A}=�ynq����)^ڵ���Q@����F����:�kf���7�3Q��u��1�*����@���}��8cݿ�-L�����G�2������?Y��Wװn���>��+t�����xj�q���k�'}�x|*�o�<'+�R�������A��
s�k�W���o��v�m?������S�d	�=!�ןp�΂6T�_ (tR2L� ���criCf0���޻��~F��ݾ����k~��[�G���S,#�D\ft��#+�>�R�XԜ�/�7��JD�}]�mۦX�vu؀)ZY����ٛ�ܿ�i$����#w_,
���݃z\A�c��U,x�a�$�-s��1k�5����B� U%�ˬ������h���44�y/_��m�}_5�yDįtӢ�Z��x���^�@�`	A�޻b
���ښ�(G�@I	C��X���	��zݿE���0����b�MGoC�#�1�O���!�U�:�'l��j�]Ykp+l9-��%Cs��9s8��^ò���T�	��y
KZ.��*�E,���>�#G�>��;&W�Wʽ=q��R@�����^��vð�x��%x��J	=aF�S��F#s��^b��\q�+V���"h����[�^��{���F�+�w��m��T�����As�M�s@�F�<���U�.R��a;=Ta��ew�_��}��a\��>�V2����F��t&t/À>
���tmִ[WӢa���5}�S��^m���F�>��E���l��U)/�~�K�_���a_Ή��:IB�0\��e6����H~ݳA�<�^�W����_]&0�d7��7.��F���x�����Y	d�g�I�0p�G��rM����u��0�c��_]/J�=��'��ne#Oز��8�]>�iM NKm��ĥ�����@F�(*�'�?�S�vGnm�X��TMC����*�W�Uv��1��I
���Sk�6
-��� ��%�5y���?�y�F����2�r1s�kcY��"gۋt�P��\�E= ���<c�=����SUe�8!*�Uz"Б��lT⣮خ`�Ɉ�7��s��(`�,��vUƴ�B�Ӈg�d��e+WmN`�5�����y߆Z���ei��>����7T��`Lq�p- �YxI�^C�}���͠���=7��'����B�-g)�s�Aj"�QJ?�
S7?��&vcJy�x����K{{�wZ��{�ŵ��������M��d<�-���w�L!��v�6�F�2��e�یU)�0�8����_O�!���u#��ɼ��2�kb/�.ex�����	\#���M&�(-e~X�� x}+x��mc&A�L��$�.�2�t�p:�>ZW��ݯA8�� ��r�ǭ�o��m�el�Y+}�bt��<>��!P}�n���7���X��r��J^��W,ƕ@V� �%AKSA�s�Md����:�CĚ6����yh몬eņ4C�h���u5h$���,-����?ơe�Qݽo�4��V�9p�#��سxa��Q}�I��b't��LίOb��[��^�]�L�f�~��X�����h�O�q������G�x�dV�ˉ��:uhP`�\�� T�T��	���Zz��9��}�e8��Zǖ��,��2�'����v<+a����t{�	LL�:�~����ڂ��W\UT��0��œ���D���a/�fڏ���g��m��|�2����K��WX,�cQp�J�(pAIxM^���#�4��Y��KmI��{�����5�QlM��	GN�3'Y�酭V�e�,�������FwN������ܗ�e�z��ût��Z����8'�'��%��bx���1i��Δ��{ N"�ż���%*w���S���$�!GRm��x�k3'v�[�:��ue��g޷����pf�4RS�ΰV͡4��$zE[G�f�\a~����2�<�f�z�����J˻B�Z�d	j�\�3x�����Mc�S���7+5A��#��x뭻`{C0!gv�E��P�HM�k��5�{��=�)�D�����-���Y6�N�T��h#�r�F�K\�>pn&0ף�h	�Y�����,��@~�&x=8��Y�B�0 �n��^����Ed�Y�Jn��jb<���^�
e��{��s=�$�h:T�93R�L�7�!����d�N�a<����C�����|`�L�~�����>�#�/�V|�����UB�ukY|k�/�t��Wyf.���Ɯ�8��38pZǣ�R��*>�r�b�]���,g|��9����HyϏO����&ʓ��A?��!�`�x �~"�>�*����l���x '+a��'K9g6��)���G��By�U�X�.>te�%��a-�������`�,�����#�KA�J�}T�Zɦ�M��ey]0E�Q�bM�q>5P:���R�d��l�,�;��A��E"�5�[
;����)7����� �M�U��k� ��dAqR9A^�u~Ǔ�@b_�Y��B�A�I����&��z�>5�{f�Dr= U�4�aw�r|EnN�w��@2�W,܂t�~�W'�Jz�T���fbSK����?���b�D�:Z��tTC:��{�˙Z��=��}��!h!A~v�j�F���z�_���aB~��FP1�<%�Q��>Vr�qz�n�1�G��J��Q���S����Ҵ�Vg���L]�2=I�q ����^�����������	Vj�i���9c&b�[+�/��R}�0���t��@��+r؅�f9_>��t?�1q
Q
pM`i@n�w
]_0������,�A��Ե;o����`�K�4�s������ /r#]}��_A~@P*��
Ih��!��= u� �q��9�)I��@�c�=œ})�Rц��w�2}Yg�c�)��c���"8��胈S���ߑ6�M�t�~�2�1�bL���k��k0Y�����=��T���0�h��P�� B),�yo1Glp���e~��r�@}e�ω�]���m�x�*.��H�Dr��{�#�}7y����B�܅A�f���'��K�>X;�.UtxP�!ni���zV�1����2�撁<��u���_������Hc;���L��Jk�&m6�8�*���`�ưD���Q+�~'��\\*�l�mυ����x��.�\�<8�5�N��:V^5�K��r�m6�-BFg�k������ݳ��8�����
��ci8C�^��7�
7וƦ�%�PG+���]2Bچ�x���H�S�
� �LϬIf����k�2�4����R�>�;$ �f�:Q���
\
��3t'���j��B��L#C�"�r�-*a��f�y.2�"G�W3�C�xWз��z�"(�{��I������]|���xk@_��Kd��c#d70n!E惋��!4v^J�w�T���(*陜��������PŊ�fmt�'Vq�1��lv.�M��q�0ўp�G�����	� 0T]�V�7W>���@�T���\��u�Bs}�,ѣzq��p1A(U��a �UM(E���l}�Q9*brh#�u:�8e<�շ�E%�2�Ti�w��֋����X^�����-I<�������oP�.�F-�3�P�˜��[�/�^,�h���_[֬�Z�(��2|��!��jԿ��'{�W�IwP��$�-�=N^�=B��	�v�nF/{K�Zg%rU���.zWt �i(m5�P����q'1�r;2;c��S}p`�(-i��jMJy�1�&~w�L@L���ɓ#���/`�&2�?5)��|x�P�OR����ڹ;�b�S�gUyMa���x{�D�4�Ӕ�z׭����-��l� N5�@T�DR�j�/*�C���5a�j=�c�2�*_��iC�ɮD�)�ɳ�%�;^:?\����O����5:�/�J�w&�R��˻�����:Y��q���,�v�+Ds�.��X��9�(�S��m��d���@j�_۸�[x�����̭Mwvo8�2�6��(�do����tW���ש��V���lvV~طx�*L�	����� �gh_d�o!w�Y 9�O�-�~���mtP���ˢ�f�P�k�/>\鎍����pBݯ.��c�cnY�*B�>��~ԥ��[��0�p~LE�/	�·�J�x�a���2�s8	Di��Kcq��~�>��O�Dq��W@�v��t�1�����`<�f���e��.��U�f�����|ҩ��D\����S����<?�f�8�g7SB$�,�lfS~�Q��3�/�(_"�|��/¯�+���c�:�/�@����%G����+��R����,���l��޳�佇17�CX7��A�ސ��R���Mϧ���Խ����ߣ��?�Rm��#�~䨠k)*���yx����L"�ۙCbٵ��E�}W��Ū���Ħ�����W�����nB�_��'��HJ*��jea�%)�^�d�Ӂ5�g�׷ގ�z��[����"��rI�w�&�ɜ�us�@�ٹ1�8��f��}��%��ʳ�m���+ӿ�>�h�n�F��������>cy�,)�r�
Äs�,�]�7Q���t �m�C�a��
B��=!�>��IO�~R�Ġ��n}�@N�����C���=��@��@�0.�Iy`���-0מ�P�(��Z�wp6��,K="ڊ\��~~�՚���\H��ld��Jju�P�Z5sr9*k��lr�{��'ve�/{/ �z?�8R&����U�)�3}yi�mA�����:B(De<:��c��Vm��d�K5 ��Z_n��n�&P��e���8y�Juϩ@�s��*H��57 �2o�����ĉ�a�� �㢪�Lj�K"�G�(��Y{���>�r�4�k��w�薊�Ԉ��hY��hb�����b�¯�OI�C���Q���^j�Vq������}�;��q?�r^�]���?��#�xb��38,i�퉯�@@k��EIC$2{���@��n=V �׭6�������O���&�s�V��FZ^`d�6��xrYfq�6f�b�	xD�	.�w硿uFUr���e�T�K���.�ݣ�_����;J�Z~<8���,@R�:C*m���U�X�7c��5q��Ԫ�VK�d��q:�#���^�P"�(���I ?�	�84z�8���-n*{Z�g!Y!)SY�J���Nל�j��0�9񔐏��.%Vxe�
N��l��i��b��J�Gw@�3��ط��1G)め���j;����UM�K�flxViJ7�N~��D�k�B�|�xxg1��I�l��T)�Cv�I7�*k=���ȵ{�,,�����@3kF��vg�C�%�C�>X�)��ѶM6>������s�ݔR���p���H�hͰT���b���"����ַ��S��=q?tW�Y���K�-����)��Ye��zh�n��0�*�������KWo�R�� ��ĭ�$;^��ӕ#�-[��mU�RR�J�|�M�?�[����K� ).�I
F]|�E��
nv��(e�)CH�B�9�ؗz%dܩ{'6�H.&��˚�n6�ڸ�e~��0�#*lt��~�R�E���aN/P���A%���&���� �$Il�I�:jt�W��x�XA}	Jh���5��Sߌ�c�4�7�H���� iͲ��FY����BK�~^	�5�#SJ�b����������#Ys���!����mMO��E�n��Bd�^n��6�򍪓m!�3��ls�%���?����tЩ�0�Ŵ�J�ѩg���&��R�}�	^Wt�p]�6�:i��a߄�>k�8��+���c��u�i��>uQ�+���k��~�#Y/C��I���O��W厏|�E	 ͪ�Q���� j�Q#�xkc���DT�F�{���|���w��K���Q�Yi��1����@W�jI���)�疞�$-��`�Vwv��E�U�� ;T	;2,z�G-�t)�f�t]>s6��%weD��Y0���ֱ��L�t�����SH�n�T�ߓ�B�����T��zzsԟ��a?e��&��$$
Ƅ��'H�:G!_@�j���I]��Yeۆ�H��p¥�`� ��җ�>���2�EC�Kq�3�-������Desσ��/�%)��ΧP�Vei[y]L�J�&ڵ��֮I�������ǭ��������|/��:I���r=��{��o�Be3	5��O_�0���|O���>S�˞./���ğ���"����e�"U�=�/Š`�����/��$6�+Wi2���	�1L�/���nȃc�Ɖ�^Q&l�lkN� Flћ��ߟ �^չ!2A�K.�fk�~wW���T�>�fw�{@u�y]"��P���v�U�N]٨�^�$�e^�߶W,�C��7Dc���]x#��>����G�B�8ǗіPc����Wf�*I��i,�WWs�R����ńb��q�C��,w��鲣�X��VVX'�_��sJZ�@�ÑQ%���Bt��׹�ny��
=��n$�F�H[��=/�ߑ�^��A�����ԣl�W/H�	Afe�
�j:���\I��;��2pT���p�e|@0}�R�1�1��#|�U9��+6q��'����qꋤPP́2�J�&���W�xy�f͕��u#�$�'R,'��/��W^8�^������!҈H�Te�'� CB2����x������$@ԵL���C轭�@���U����?q�b]�i���?B�lݾ�
X5`\5 H��}vƪݴ|?QGI��_j�ǩwN �.ڰ��OE'gp��<��r�����[gւ����L�^�=��Vj�x֜���Z��M�����#���,ےI��"_a��_T��+�,��6�?G)֤�+��;;����z�~��A|�D�����UzqP_!�p2�)3/���!����i��ʧ��1<���is9s��aMI�vD`W����ﺄiK�Y#�����&�Խ�z8�v�O�'g���
��(��6=W��-a�sJ�
�6z��΢@��v����
�C��C��1���@lkV�"M9l �%5
����D+������g8�:��[ϲ`[���X��L��*�3��0r󏰍�@'�J6u�����ߙ���k����hP=�����ձ�bfZ�~PW��~�8\?M�Q�M��r�n��HP6'�fL��1s#��915֟��զ]<�/�4�� At�U���+���������拀��x���?_�5��
"���)�6o1B���0
�߅�Z�Z�O˚bե��ӄ��/x]��kU�
�]Q9��p�OX�=
�$�5���C����&V��܎Ǯ��k%+��[2.�Q ��J�[Չ�+<*R�ūWʥ`�"JnK�����8\���gT���������[���B^���p��]�@�5���h�=��������Q� u��a4�u�,E.oh?��z�O��*�ɻt���ޛ.#��^�X	o2ݚ�6c�q��0uU�ϯ���4��#E��i�����K-֟�O�1|�@��l�g�������U�����N������,���I�D&MI&�{��� S�|�@�ǐ~s2�3���[��!��7�D���G�t�q�+D$=�@���W�$(�͟��'���7"#P���n���ie@cր�����9��6���k�� �{���>�N�X�r�3wn��������O�KK���vE#�ϒӧ�Am�wu����	�Bd��^M��U��J8t�U1ŀ�����<�S���
NH�R^Z�3�ϭ�_��D68譋���s��Y�b>���oC
�X�2n�����[[3"2h	>��^gH����t7�c�ܧ���k	�ɐ�+����$>�����-&j�	/*051�b�$�0"O��=%��\/��w�-��Y"�M��R6"�z��ފ���My��5�ƀ�^�e����)��8N������H�K��	Fȕ���~F���'�u<ٴ� �$��6��{C�A�JhD,��%"��J|����˖��*xjڒ$��1��gQf�~��z��� e!��N����74f�Xi��S�E��-8]�����T�g�����L�Yq-D���ԑ)��1�RQ؁Q�t��:O�16��˨F�w9S�w�U�W��t	�: ߆!����14	��k���&����tvIww��\f[��W�:ݿ&]�P7L�!H������^}��{n���=ĉ.�o�4ˎX��i�����������ly	���E�D}�9�у�s��N�Q��h�7�1oi��ii�xK[9�t�h=lY����Ӆ2#V�~6�����T��1�K�xђ���]�+��WC`�w���z᪋���N����[���^��|�z`?���4D��i`��8��eѽ�
��	D�̌��H�QP$�5�x��Z�p�ɊͲ%��<e"O�L�A�������Pꊟ�c;+��*�iUL� .p7:>_�A���:�j��@�o��T��3^P�p��h�����v]'0�p��LZ���Y����o�=7�eˉJ�{�m4����&9�\���^F�i�S��{��I��!`���o����R?$֡o�%&��8-��１)�(G�̲p���)����%q/�7�c?�`���	�b��\ H�e-�zB/�0�����^��D�%dTc,�Zwn�l�3ꮻYB&�Ӗ@�}-�V`�jwm�5�2/~���Ƥ��x�l-��"-c���]����54̧2��	n��p`��t 晝���TT;�pN��3�\��4#��GPd�_HR�b	b��C[���[��;Ue����/D'�Xk<�p�c<9/9���zn��pR�0��,dٖ��c =7fTSa��0{��V��W1!_;qi'54�)�es�G��D�2��o�8�Yɓ��3����`f�����E�� ��<3c�>�C���|ē`����������C��,����	rxtf^��^��*��p�5��w".�ـ>���M��e�6a�a�?Kd����?��>�G-�)��(n�	2��]~]t���Ι`�k�2��NN�y��V� ���W�p�v�o�
�J��j^H\'����ܬ���ps#�<Z���dԨ&_�=~�poBx��$�~��ˠ(u/Z�0P��l��3�R��cG���;ښ� 6��8+���vS�j{>�[zҙ*�j�H��V=���(�ʒꃞ�xR��%GS�3����t���ơ|?!3��T�@,ե��կy���'���m�#7����pwuc�l�}D��L���}l?�~#����O�#D��0XN<Bbl
���?���l��Ft��aMv^Hi6���b98Wa��"N'��P�~ָZ{��>̆ U{6�b_l���'���t���A���o��N�DcB��	� `r�7,~�܍')���9ا^��5�w�a��Ӟ�@+�������<�MCQ_�ZL`a����(5�z0#
����J\������>���b+��Ft����׼�ӆn�D&F褙[���)d� ��>�a�n��ZlE��ᣋ�l���B�#_�-�I�}悈�%��� vhZ'�į���\�쿑|J�8ʹ���dss<�3�6_Cw���5D��K���n)|�H��De(;�G�W��>��t�aA:�f
�b�ۘ����#���T��?M�C�`_E>��Qal���_R���)��
toe�H�v���t*����xr��,�#JP�����;�W���+��z���޹��SK��<x�3�\��V�rR��` =⊟&���J���j|	hX���uT�S� W�p�|Y~~�U8���U��,���-#��8�S�໌��m�W�7�:�p�>��%����橌2vB���WN��Z��4����YV<��O_��w�É�����-ϳ�(��2��P,��A�>�<APL��i�U���\I����[�����^����̈a�j�S�i������E��~�����:�����Ws>2��Z&t�S�3M�}#��
�E�|��O���. ���	I�W0j�k��	~�lAa$?����7c�`2��5�j\u+I�V,]���S�}��u��_̥��Z��_A"�:�9(�� �K��c㵢��Մ�Еn�)�l��g�k�B��k��{�}���]�UaR�@��`�#���O���T\Q�{�߻yiG���*��	f��\�Xy�aF�ɤ�z`/�H��Qg�ϧ���|LP+�|W��К��UK�/U��S�Iq��gR�r�/ �!iOr�WQ`X�=�
u���t�[Ԏ}|�7�:KE��X��1��8��}N��5������I��9�S�):�3B�(���IT��/�C�a~���%�pnFk��a{͕Y߻�@��#{/t���{�{���4I#�BF�.��E�}3�+j�Y�Ca��_�X�P�u �d�A"����F�$#��q3��%ij��J�`5�Lf@X���A%�9��'�>0�NgI|�sɵ��=c��d�-����3P��A�w?��bd�^�O�x!|P�0*�c��F^Bѩ{��U�����هA�؞V/��:�(��|��ϐo��A:.�����@�ƕ�b#�dɤ|������D�	1�`�d�n�N��Mחɠ�<e�>�ʭq���JB[Yq)�Td� gS����蚐(ʮBo�9�W�10KdR}���#s�~�,�Ɏ5Mm�^^ިN��0�N�u��(Dz�-9k��A�N}sޮ�a��M��z��'���h�A�z�m��c���rxQ�EҺMgh�M�	�:/��"	����.���& =3�
wb�6�R�{���!^��S�N�	����3��pV\��x��%�*_qA��B��o�ȔsB
�c`uf΃�4�1d*���n�LQP3�ީqsqJ<�!D��z�Ƃ4�a����Il���n!��u�Bu���\]�߈�
��rt� �l5�p?�_X��mJ$]��.��9T�n8�K
~l����t0�3�91�VP!ƛ���`zg���VXv��^S02�WX� hp�# J��50?J U�$Āsq[=�e{(�&�k���TY���:����R�[Z&	�Rj���{���+���r\Ʉ��
Э"�G%$,�n���?:�P�l�u]J�#�v��];�DkH��l�v�lyZ��4��q�ʨhC�@�G�됭��g�U����M�si�,V>���snZ#�)Y%:����8�J3�17,s^X��Z�T{��2XM�3
���а���|���o��~�Q�+H7�Ij{����ʉXSH}w�Ѷ�f�����>=��}H&�:�r �g�d�j��g�	�sK���O?���d��x[�鼣,�H/͍�Tv�;E*�jj�h��&�5充� o>�%{�	�����3h���i��_w�/�H�'�B#�sw����nO����0�*��#�{t�J�hW��|)��U�z�E�f�Q�.��'�+&��LJ#w�~��ִ��θh2�I[�"܉����	�1(G�d�~~x��@�v��qo�IwG����}��e��=�]߁	�+���o�D��s�7������<����n1fYq(QIhg��ss��0;D�����q0u4r�ѷCM�;���Š*j����^���(�E��pW�c?5_�I�<�W�������N;Y%_�/y�ɗ����Îvߥg���C�[�t�]��%9�uS�Ǜ�銡4��*��Yc::.KZ@�9棶(]�<�(J�i=(N�Z�@�W.��7t��/��3�·�-�k��ꈣ�C�W9̔��,Qď������%�����nX��v���Y��p/��ӻ�ι4������n�cQ!��r@�d7����\�bz,y�$�Y��}����e�����YF� Sp )���8�B������H�u��R^Sx�)XTr�����M0���F��%��䀤d��@_��&;�p��^�;o�Ȱ;e<U\q�7�~܃O��E��c`3�����y��t+��*���f�5ߔ�K"\Z>D��Z����/��I ���ϲ�!7j�)�
���(m�u��Zd�L9����*e������@PO��b�
�V����ҍ6_[$IM��D��'�|�3��V����v�8��vҳ������_��Mn�S�hXy"&r�`��Y$h(*O��m"&�ܲ�7xvhѸ���x�m�ҩ"|8u��[.���7t��%t%-00��O$���0��o�V:��۪��V6J�҂���ĿW�n�(n���֕���*��<��H��	���-$�&Tu��5�+.��
 �2�&V���6�[�������@#�%�5����d�ra��8�� O��E<-�� �}�bmͿO����uF<Y��ާr����Mp�{[G�� � �N�7y�vz��voS)� S����h�L��	{O�7�3���Vd��-*�~-���϶��/�|�����wg^�h��~:y&Dq2c�#w�����_�L9�+���-s����.��Ȟ�o���0���Y�E�L�*�k���/$�;/ۖ�a�5���ۤK�3y��4e�Z���0�ש��~6aZqUh̰�	`+�CK\��j�;����\�$4���q�7�ѩ&�z���_��kT����� ڡe[a������qށ�36���0��(_\����*�{��iޕ�!�ͅ�m,������������R������V�U@��&.�����0������!�N�Q��~�>.������+�s���KOl=� ��q�ű*� �>��UO.s�/�:�"���顸��S�.���a�#�4�"�o�wk�w$�C�%��l���D~Q��󌣪H��c�t�K�3�Œ����'>�U���-�N��Z��G�d���:��]5oW#�G�>U�V�A��%;]S	3p�Zq+[)v�jY���p��˻L����D��}�	L�-Ŭ��<{��*-�t��".�gۖ��2�2Mz\�k.�u0a'Z�Rىl�p;��''r�m?-����8 ���]"�w����'zP�r@K�Y�7�Jp�Mj&T��χn�ũp���0���w.��"4KvU��2}o��F������:��3��T��9���_��$gjIl�ٟ�E2��r��v�;

��'� ���,���O[��4�D��!Q$9�'�t��V�������b�6�>�m�����oJ`RM�x
Ǎkxä�ݕ�78}s��7G�m ��jg�d5�9 ���P�[���l�R�*�r^���LV0o��yA��Wú�P,�֏Qm��� �fՃm�b� u2�/@��b�Iu!��i�N��^�2� ��h����Z�����FrB�*p�]x�_�W�o�g52���#U�X�z���1��۷,���f��V�G�z//��E[�F�C)�)�O�����}G�\��=��`�k�a�%���^�E�����Nqqv��B��r���0�ڶ��Ǖ*�M�S�${�?f�j��D2������qP��ϿxO" m�M7VF*�~���e4�3EX�����F�����[���G�SH�D�����E�G7�wx�"g ���#љAe1t��m촗"^\�:� D�v���3(T�Q3z�|��Ne�^�*��-�1l��F�:�]/$ m\�������x�w��Q{!s�βY|�CtJ�V������Hp]�] |�#�K�mW�F�V����Z�[W35qǈ!	��l�zё�b�W�B���}�@(�$J���Αu��1�^u�(㱛 k��!� ��O�uq�K3G�F��F�����&i��ˊ���G���F�G�O�q�����xm��k�����vs���7�;I���j{��bHg�5�%Q�Cy�۱�
����f�R>"!�=����|ӦHF#�h��Tz*0������N�䳄&c-�=���u�h$KM9H
�EA"G�Ԋ`�U��U���*Z4�
t��r������l-��N��
�1�	�4���?��?	U�êF"��� n�V��}{+}�ݗ�ZT_�����Q㼫��|3"���
�H쟠�[ι�W_�-��C���b�R�a�� r'�*s0�I�.��wUSL{��,L#E�(PJ�.^
�a���i懥|%\y��/>P�~�8�O�WH�4�r}���S�b���)�A(k��ü�{�$�!�L�3�ӑ���H>$=�/K{�L@�� jͶ��D��>���J�ĸ�k��q��w|��A����[Y {�Fo-:8[~ܮ7Q[z�B~�����Ul�}�Pm������;$20[���).z}	�(i��YD6�XU`T쾇�oyvʏ�[)������vb�����b�� r��9��3VKeN�\�S��ޑ�W϶���	I�ؓfA�aA�v�,����X����MT=~Y���Ԕ�7�\P�H��c@�С���N�'�����_�q�wC��bV7���x@X�o�^?��*�J�QdLn�B�0�\��^���r�P�� �<���Zl3k�Ag�x�:ou|��K@�Yֲn=$Y�G�[ʈD�1s��ܘZ��� ��UA>Ej�>9���pBc챪;���$`btv��Y�9m�(�ǑyV�A�BO�6���y���C0��c�v���2��.��{����ڜM���i�(�cf���N��|⺈��Z%����P�KG9e�x,�i��h�X`[&"��}!�)����8�Su�H���D�uܚ`�+�FRa�n|�p�o����������@�h6���z:�=˟�=S�(y��j2�{bg�0k�h�F�0d�8�v�^�9U��*J'��7��w�"��t��1@���Yd<N/��W��$�A�8!w�L�:�����S�Ml����~�B��ݻ��0��� o{�˻��(z���fht��|���$�֙����-2~��O����"Q�-~�s��PtGn�s� �4�x�n��@!����}�ĮN#"S�+�#TUJ5X�����/t\����L<m.c����\[i�(+Aƻ-�^
L��Q*�m�ṟe/qڨ��1HX���.:<K�kP�S�X�P�
������P��6��A8��d[/�8 Z_���LB6ݱ(���c�y��a��;�>q���hM�
MՃ!V�[�מM
n�;��|����d�JZ��?=ժʫ�l�]�è7��Z	��S�r#)�z�W�}�h�&�p}D1�/��uc�j�\#��p.��U.�ZV�d��0w�Nz-�	qA����O,���Hr�T2h�oZ��I����<��~���8?X)���ɚkV��f���#C��A��tmb����px�ǚGt��41p7���i��әk�,^J�?��l��MX�����c��+4ƒ����k�n?\bS��7���*�kr�p�6,ޞZ��};3�f!�[�RXk��J,�{�����T;v�>;@;6�Zj�#c�g)$����~������W�r�z�c��ּ��RUs�[�	c"�k���K'=f��5� �՗�����{z�MUa�ey�d"��Z=ш�
�[a���d��ٓ�~��(��>8bl�0;Ʉ�(�'�h��.��CS�p��'[���'����C�� 7�ĂD�m�R�AHu`� VB�s`4
�g���-Yk� "Ázֱ͓BS|$S�?e�E�\���N���N�Ľ �[��'0Y�b���A�����H��A�L��)A=��a�������Y$���k���b�ET�����ơ_��v+5j�o���Ӆ'mO�Jx?�,�ز���W�U������>Ot�0}� Ĳo׼���Q���~76ז��"5���l���\ŀL1e+4��v��9�m�	��"P����A�yw[Dϒ�*�Ʊ���/�4;�)���ٕk-k���Fʶ���ӻ}���&�I���.#��$
�f�ׇ
;�M���8�)�0	U��pȒ�R��`������Ѥ�NjD-W�W&��q����C�����ӆ�'��2QTA��0x����<Q�wؐ�@��0	�&\� � ��w CEu>���^�h�Y����d��V��������������1j|3<$����/��?k���'s�I��TV��N���峊ϨZ��������w^�䀜�������^\�<�ns�%��#b'�O��$SgƂ�c�%)�Yj�Qq8����o���n0]��J�頊,�+ۙ��$9<�Y��<F%��
M@�D��J���릙s �\��a;6N�Q�Q������]�uU�,��k�A���j����L���E"+ͧ�4���8�s�鱪�a��[�"֖��B����&��6�fX��ѥ"җ �ܺ���O�ZRL����Y�#�3�
:�b��]�-�Q�0Tb�|��@��`���mG�*�Ɔ�����������	"��ܰʟ�ǟNr]��~�&��%�dI�Z4M&#��CV��8�;[�b|�۪�q��:�,������'Ç�Mc Z�ϔ�؉�:F�{����=�f�7Z������y�Dӂ��ł��q�.�u*�)�u��K�5�Ԅk0,��E)I�o�_8}��*�o8fN�:�+��Q��U�og�����@�q0�*6����&���%F_��SLէ-a���>���ApzfE��Ϣ/[�O�X�ur�$������ G`�	���q5�YH�KNVE��?�ǚ�泝Y^T��-q��sٶ�M� Ɓ���4���?'���/!��Y�={7v��?�7�@�U��M�urN�W���m=&��C��ړ!���/B��1U��k�h�ۯ�>kwKw��zk��26[{�ɩ���n�+�E�F~$��z��𰃬��c]Nr�K!/�U$�uZ�fD�s޹��?&���;1�A��%���Ӯ0�#������Kά�vղ����Ut�i&ɡ8&;�Lծ��	@XO��/�c�!O2uU�J�lh��~�Ȍ�ù�[Q�z��W�|>J�ʰ��L����X�Z�q��E� *ami$OQH���ꄏ,Q�����7��q���#3\4	MG� �C.t (|�o4�rS�2��Up@���t�c�����-|�}H�[~!)�E�9pbpY����ϓu�5�=��y)�.|��=�}6��M�Nuhp؆�-9�.��{��~AQ�d��jB
Sl.](k��F��<�����@��|VB�Pj�E�E�����?�>ǟ8f&��W'����(��� �
}VH������௼w~,�V)K@W�#<`�s�TO�0�W,�HȐ~a�"g�0�C[�Jāj�F�"a�W�%/��!;1�Ǔ��:Q)V���z�'R�戂���_������ C,Ԏ&� q�$v������tW�ܝ��k07 ��%���։�qhd5M�7�a���C���}��P('x�U�p����(wS��xZS�0����]��L]/�߬����U���z_D[�=j�>��</��ͧq�qm:;��w�f /3Z�����I��ռc���3���9b>?�&�m�;�+�A�Dos�^�S�/�K��z�����5��䳢��x�Ȏ���R�h]����}�׍�g���~�'�J���T�����ͳ%������n%�8�.��Bʀ�	317|�xM��+��I�Dr�y���~�e��1����cSR*Q��%j4SU���N��U���	#y�l��p����(; �_����pF3A'A��,A�9seo\���<u�3L3��U��q���{��1�t���!3hx18� �ZSI�<�����z�r��J�����0�ʽ���+����m��?��]���ɔ��{�p��6�����+�B��o���!m��]d�P��\=:�4�k򱄕�]S����6���j��Hݿ�e�8�k��|����������>�H���Z�N䷖�Tvs/�[���%��Q�<b����
W<G�����U����6U[=M�+_.k�����sUKbv����6 �n�nb��kǅ�w	���$rR,��Mȶ����S�'.ĕ�!
|u$�鋩������O��$50�0DLS��j�WV0�Nz�&�:����'-�5j�#�� e~�/���a�%S�o����+�������������^7$#��J��1Yp̉�|B^
:���,g�D!e,A)'�E�^�����S�g,&��[bv��y�7��x�j���^۟ av����1��Ѡ����Y3^�e��3w4ض("�/w�\fK���)B��CI*i$���:)?J�~��Z?�CU�Q��	�4-Rd�3�=YT�4��� ��y����
IVM��8I�
<���8��N(٭�f��3[�p��l:������<{���sgM>�|MJ�h��[�x��ˌ�?�*�����5�O����5�X�%�Pd�]�zչу?���J��3G0�2�#�6�J�)e�V���jn@#;�R�4�� �$��i��G�NR����ߤ͉lմ��E'_���M�q]YG�mV��4�`�������I�e�!�m�Q����'OO��hL,��;��覟��Ǟh�v��f.��8�4�����'[�H·�E~���d�Js�v���C����u.���i���^�4�J����j��3 �ο�l�Z�M�G�Kr�K}�t�w�f��/7�?z3a�����b�(4	+`�cd
S�ۅ�(B�d7�R"�QlO�k�2�O���jMw%���?e�h=�O(�nw����������5%�zw��(����a&�W-�&<ڟ�&7���A��~��d�90��6����c ��{'\� %h$q���(@V�V�_7N�P{��׃J�W�$���v��j��p�������b�6(��,��_��'*(�(��R)0�}�2 N�6|��p�3�1-���L����$�O}z� S[!�c���C㍋�%&�@����f��X@��"����E���ǚd熐L�,O;�3�5�Y���ˍ� I�.����s�I��N6�5�c���BFg2l��;MQ�gm�oP1=��W?�\uY��+�l�+eU�_	���U�&�;g��{e*;�:z�N��
5ݼ�v8M�{k`R�ܮ�{�K�ۡB`�Ap
����P]nȫ#[Xt���,���K��^����x�{}����(*,�k�]Ӽn#�:^����V�>ܥ_-�R�+����i)���\���_N�(0p2z�����͍�2�&R܋C��~يR<vH���cN#-s�/[�4�cbG(�ҰdSMo�P����R,�.8��X���O#����p+&��ѩ[�=����p���j�|3,��#�\5��@? �gm��ԄyzA�9o�/0�go�h�c�H����Az����:4�0h(�ky�����e�!Up}�i2�:5o��k:��I��1�#|qRP���5�!�4�>��Wc��ͷ�1ΈL���4:tM�����ei-�~f�	���ٖ
G/��A�%*�7�;��=F8<��wo�l��շ����Iت���?P����_؏���BΥ�!��.8}񅲳����������#���Uǃ��+������B(b�3��s)	�,�������_��`��U9��b)2������
��G�����1�(w�c�W�T&c% f_j�|s���xG3����P!���Z03�Z�q�3,�U�O�~\"��o>/OS�P'	�	���%�s� ��{�Aig(��V#����	���*b�A�Ɇ�myw�Φ���H|3$9��c&�[��(��/�6v�!���T��h�.�K����xS�N�e�@�L��h<�f���랺W��76[8쨾�:����=��ʴ�|+����h���2��1*�Wdji�^�}���h�A���e��і�!!���7�R��H��3�3�Y�D��	===wG�K�C�z&ս�D���y4g����9�]7ꧮ��n��)�t��|��C��H�#pb}�˘�~�+5�7S>����E{`��a�h,%/�����U���:c||��/���7'�I]�'��t5�ҴI�P�%��]�B_~R���7�����[O��:��>�e~��1�B_a����*쌩֞��_�|_�;<�����)1)t�HNT��u"$w�Ŵ�ͺ<����� 9�g�2��̋��u�!���x<�K`�r=�|",��R~�=J��Ns�u8U�l��RV���)[��T�1�����":ߚ'����l78��]b6oW͢��8b�����~�;�J��L�J�99��%�����㜫w��B�Ɍ�bV�?�*���wz����b����K��Xc�*W�#q�&���p�	o����L�D��:����=M����F"+p�q�7/C��lm����c�wr�4d'�cS�M17�EmmK�l���������8O>��3Hk�67uT�%	�qՉ�U~��F���&#LD� ,:ϐ���}��X���+�l^'�mF"]1��U����Zq��E�t��_},�[p��;@?��U;;�4�mOʦ��G�c_�������uT�%�ljǗ὆K����	�fm�"�8��΢(^���l0q�s�w^�}:�:�.%�$�2��҂�O�	 +)�:)j�^5	Ĕ+SP��d·�%��� ��M�&�lLnt��aj�.LŁ�}�>ފ=\�r�o#i�5�Q�1x��n|n�1ݑ� ]F��̙-���Rј��a�e�Ct��j�%�������q�X�0EGEe���Q��?!P�2���l-����@u��޷���\�� 4��w�i��۬:b��F���rf��$�ب����ӅtxC�ۅy�	I)�Z$R!R.E���������f֘Vg�����6H%!��X
7	ΏC1S��O Ķ����r�a-���y\�m��Ce�_�qz^ɶ�ˮMA}W��tj�Zҙ����R�j�|�ُ]��l����� h�.��u"�e�(�,J��{��ĎU����k��\��8���B�[1�M�dS�V�;�<�9T��������j�ߐ|� ݯ �e�!_��I�1C]��U껣�����o�	`�E/��~P��h���=��ъ�^3艢���u�9���[�<�f?�J��7��@{�:��J�,aZȊ�p��>���s�L����.�W�����jY�\�ee�:�+�Հz���m�'Й4�������R��e���/{3MŸ����!Ҍ$?�slŌ¼ٻ�yGi���U��� ���C�L-�w��,������lr]�<q�f<��%�~�b�<�h�JU��V���E�G�x8�>�����u�����'��p��U�`��4U�%��4u|аI2���E�e����"�,B�O
����*Be0-Ϭ�!�tM�0����j���!��mQ�m������.U��X1�nEj��Qb�Jy�W=��iс�gpQN�������9���l��.*
�����Q����3(�U�y��6�K6\��H��x;�������:�÷���9��;\Eo�y̩R�yh�4bN;8\id��pU KMk)r���I��*�D۸�ǻK��#("˛�8Q`\�5sU/�+d�_ ��lV����Ub�/�_g!;h� ������=,^ed6F�SԱ�֛�n���څ�#P��1l��ޠ��C3m'p��^x�㎞E�yN��ȅa�et�F׷�`hp%�X��{�NR�e�(,�p�Τ+ X�5��y�Ý-�@>K��N6��K2���tp�
��'�С�b���z��m~_c ���}�wY�����Qfb�g�[��h���7$����Mi�ݧ��UZg���\P��i�.��>�!��nfCW�Y�3n��� �[Gx������j	��0� S���W�yV7����������H�O���ιp���G��4%Gjj�<|W���n��.�����Z«���X"�߻t���Ϯ�B6h��X�1b�)�fP������HYL&ջ�h�d%���j���U�·������pw��YVo�DN����T���MՕ��7���:�`�l��6�!6_?��Y��I�O�`�v�|�_�x�k�ψ>�}oE�ݺi����m��ٌ�9h�p�Q=���*���R�J΍�y*j*%�jadB��T��Kzj����ΒCN��8�O ��i.�(j��'�g��P]sj��(�&�-y(9�jW�{���9��2�ڥ��T~�X�l���?B���� �*�xg�0@�[]4�hZ���5��إ~�d���b+��,���H�.^=?
�ID-�O����*ڕ�~.[`�ǟ�"f�'#�Wiue�ei?a���&��b�
��ث:��c+E;P��޸��T�`:��ڷT^��B���҇]�M�H��\>�U+�J/�f����M����fc�T�f�����d������
ڍ��1��+�|>�EOM�D��
	�n!/u�
���F����<����ƃ,����0�⪉f�hJ�BL�6S�����u�Z��h;�F��!6[A�4LTؿ������av�9q]�qLU�cW+�D�L-nYS���R����������o'���*}e��`������X�;�Z`��/P4 ��f�9��Is��ϔ��Q�X�0���l�T]��Z�`ۑ�vʣ![r�'^��eh�8	i1c�T��X�Z���֜T2��6M���_c�Q�r��}���[2%�g�@f͠'�
��W>���3��Y��� ��d��h���zT*����l˃�E���L�6é�L��r{Cq+���(���j��y�H�s�(>��E�h�|�!�\Z- �(	�tm4o�&��M�xX�`��v{@b�E�eL�k�<+�tUXU���/�
X���홷�ןT8LM9a��yF�c<Ϡ �N��F��Y�V���k
}}���E�]h�/~FOU_�`�lk�\&����hG��TՐ����7i�Xˤ���a	M>�zQU,���Gop=q��l�j%��w)8U)07�0�x=NuR*"��M�\.zW�2��%��э�=p���~yKP��aY% ջ��V/�)ުS� ��,��;�~OF�i�),�����K�P-W�����nj����'��ȿ�a�@'���j{���
����A������;,Q��Q� �:�`��ڴ�k8w��IF;����ڐG���Jd2-��HП=tz��u;1ayڷM����u�);�kg��/u�2K� �S٣�ԙ��ƣ��}��p�N-p��[Y�8�������D��84r[ۯg ��*���t#\̜$24�e+L�J�v(X�a�ɋ��h>>�oX���1f��n�W�*���K����Fxpxg��p�r�N��w�Q�7��� 
��
��z��_��Kܴ�������
�pL��Jq���`���P�4p)2�8�o�`�4��!mb/�[$��X���q�]y���r�gX[��W9#u��_���Z'����:Pq���E����b�νe*�������]��,X���}�"����S�1J���0��a_��r}�ۣ����:��A�x'�Ӛ�ͩ����5���w3#B����k��`o��N���NX��~9Ҙ[5�� o�P�p
���#MK�O_V;�g�
�NO��i�y�,��p9��3!�,����ɎFd��b"�N7���5���b�,V�Ku�(ul���&F��4��[ƙ/O����a��΂Z�M��,H�|^�_��`$Z�I���o�(��`��c�o �A	�6Ӛ�eTҲ�(��#�T����K����5 �LQ�u�M����fTxE�G�Y���/_�b��Ǟ0T�i^� �ǉ6D���B���I��Kߑ��T|�����Oݚ�V�|�~�t�iL`uӭ�,��7��D}�i�d7�quܧ�}�k��A�ܽ�-��5c���%��_;�i �@��]&�Z�ye~�0�
�QDO�n��Y�z�^R���]��JӃ8��s�M�t�[�T<]}Ϲe�P�s|�1��%m�|�f�� ��X�x���eV3����=��`EJܞaM���.\|�9PV�]q�N�W��O������Y�/�P�?3|q�Z4-�j�&�"�0�.������M%��EicζZ�f�>J��9zo(i�f)U(��wlkxst�ƜLt��#.�E�����
�UD/Aئ�Q�O����oU�mR;*#f���!��>_>�F�}��K(QH���
����C��@��v�_b�q=���C�.y�bs9&{����4�Y8�R���Q99�?�~��n�Tnp���=b�NI(asxje]c;���m��٦_#�d��ܷ�|�P����S�l����BM6�M5�y@IL�w �[ߐBN�|u%;4n�.8�ܴx�'\���q�L�:a��E��{����0�����l�A̐��#��*SR��5�u�i�}+�Vf�7��<U|΍��<vs*�db+xX}�<���e����Kl�J2�M��-g@�er����d�\*��9�pv_ 5���._*E�fIj�:�C� ��R26½�-{�)~�8�84�1��&Uҧ��4/P�+>{����W>������@��/�,���gh��Z�3��|2ó��{���$P��4�eS��JT�0�#��̒if�1����I�N��TZ�-*ע����HFA��m<�Þ�	G�OO���9�KT��~��=6N�и�ֲ�~�=w�)��lD\Rd���s\h3q!զb6�J��8�r��Y)+P���8K�N�+P&,��Y���L?��<��c�R����Ŧ�@]�����$�J�������f���M�bg>K�+��ނz+u{�S�l:�W�����"l&��&���9-��E��Nu}(w����?�,U��y0
�<Q��E+a��&[�T}]x�C>A��f8=7#m��P��&!�7��=7�Y8��� ���D=���]=	#i��X�8,����i�oҪ�%C���*�G\f#�d ���rRb0}Vˌ�
,�rJf��< CiO���,2��%����t�&9['��>:��EB���7+M�[/�ѥU�(g2Q�e,��8��^Q�I({�U��m��C�/� ��t�ͷߗ�Xl�+���j1Q"�F�2r�C�J�/q�Nk7�����%��8gC��w���@�S�3w�rP��d^�)?Y�ˢj���3$�ɻ1`��K�ľ��qS7��CtI��2:��7xB�{�+,E"oeȯ�s��{�.o�˒9~a� M�7���<�/	�b�v��nN���M�6ӆ� Ehc��-����C����U�Jƹ�M ��{_���H�6�	��r��;i�^��<=�y�,q�Qc�1��c(��&,��wҒ.J���'n�g����v]FB�گ���~�Uo�����U�����J{�@��1O��ӂ�ȋ����p��X]�Y�]��i��n���+������6���y>���2�X���.e���+]�_����h	TUp��Iي�����D���z �}ő♀l�>��\�(����4d �;󥫎>]uÉl��gp98e���ϟ�
R݁4��Ϳ8]�d�8���2�?�_���ӝL�7F���]zj�%9N��{ݕ�����?�J��bw��x��5vTv].4뚝�,���:ԡ����A�����a���eq�I�������!�v�/����߱�f�S�^���Nϕ� :Q����F���<��C
0����Iw�)�ն���{B�?U1x�Y�:d4�<"�$���6�
$ؔ��y[5��i(�,���2��8��6��\c�T�`����^�i������H2���k^�����B>1�� ��1���aOup�M��Y>&�SE�-wSr�-�s��^��S��z���m컦i��Tq<A.�o)��i��%�%�~�'�<�h}KǾUe��F� ��*��M&���5��p�O�ڜ��y�@��_���,HG��<B�b�*�r�י;�%� �s�(d-$��`r�AH��~VVN��-���?�_������C)҈X65��<��]y�L>[�dܨȤ��/���inex��V��za�g�(I�@�̸=��k�>�0���4
~Y�I�!�BW�*}æ`��H��&�(��P����|����gZ�E��LE��@��h�S����S�����4�o���D��[�R!qI/�*�\��"��S�ZC�3;y�$Y�ȍ�T#D=�ޑ}i�c�e(�ΐ�Z��?/��eϪ?�g�A-5���{w�|$^tT�#�"��s���!~/��,Pg'&7��' u7��ۦ� ���'�Z�	�o\�(�I*�S	� ����e�I��BД�Bzu��I/�e��!�c��`�g'Q��@\���?����t�:i����,9w\f̋�q�KN�_�u��8a�MŚ?��	���=y�:�W��/�Џ�7�Ɵ��ܙa��5F�A�z$8�}���N��፶EX�=|�AK�o^��i�%�9]�/w-E�ΐ�*q���v�g��\���$�´߭�2-���ߦ��S��;�|;�K�$��̥aX���!�雬s���R7�߂��%�ѝ�@�;��>{6���EْW�{4�n�9��.,����8|&�U��ᴏ�L����������S�Rc�m��9�_�=6�
͟Ƥ�F��Ĉ���Q�.��/|4v+y�Fkc�`��o#����g��	,<�'(�n�8œ#��'R���@O��A���VeLL�]+����tQ�)i�ӻ�4e�5��At��{hq�%g����H[�Q���MC�/��"mι	6E�=�4���ŗ�Kh���,���C&.���k�ݶ�����;���ᮼ�=	�_� �x�ޢ+.fh-^�`�@���ePs��h9�������\��Z-����˝�=�!�(�!��j��$Cӝ&j��'Ǥ|+��}C��؟мܱ���	'qy�L�a��7!�xԂ���z3|��~6���0^'�EP�ռ�;q3�����;G3W����1�eb�q"�x��I����_��(�ȵ��/w�Ct|`�y���&l)��":�@�����G%��kw:�Z�79T�ܗ@��b׎�!��G�����nU���Ǔ��v�Ď���k���^�����a=ͅGaE��q3����� ���5y��N/-������T�]˭?��M�Ro��������c6B��UÇ�W���vE�g�$31�K�3R!���g $`?�B�⺲?zw%r5�
�K){Zn>��tq#����=� Z�bw��֠�ѹ;�8�<�8����˯_,V��{t��� y�Z���9,y���%Z����x|�xJ���G�Z�$�n�=E���@hpM��I�h�� 
ónx��D�k����#Du�w]���I;��T�Ա��V��C��{e>R �q�b�t��,lPk=�`r$-�Vw���hq�'N�(��AUNፅ+F�6��2h� ��O�m6�o�1z�M�u�tuHLC��������4;�2Lq���GɅx�D��[�}%��%�|qL���P8���adk6t�	_��঍�ʅ���s�s{��Ayk��G���e�$"o�����V��K�x'���\�Œ���P������eDȴ��eBm1�o�AM���;�4�c����/����ȼy��!���-�����͍���d?5�G��ݽ�|������i�*u
���]������(�d���8ə�>���|��a�} �0�B.]A�{j#�L@ԏ�E��յ�`�i�+tǘ��]O���N��R��U�f%��|Ugq|�^T�}��+Ds�e�`�|���>�	9���<Ч�iP�z�Ȼ�#�C�Z4A�i�a��ۃC��%8
[J���T:��@�_M��.�*�Ϳ<�S��i���@��D�w��:�%���"��)LM�e���W��a�y�$�y;#�E���&���y}I�"x�R���<ձ	CD�����;�mK�f��Ӳ���+M��U�ʫm5l�]�*��s���H�
��}��}���BC���Ա��ΏȞ��L/��H��S�+�P�x��˻�T�2�@ J�oηq.�猉�}�X��vy�jɗ{�k�Ό=�[�'�d�c4���Jv/SJg �o�4n�t�WD��p����kV)Y�rz�������݅�HQ�8@L�`�ȏ�����-��i���܇�b��r>�r��Z;kY���R{�D�F�_�!Etl,����� �L���U`�:@��P��xc�zЀ�� �W�k��L+�ҋ�k��F?a�ǔ:��H�e�>�&v#Oҥ3 鼤1��e�K:�9�m��G��U@/DKv�Hr)�/�.�i���mz�*���3r�6m�7x*rs\ҵ��+}yn饐\n��Y(���%����OT�܀R.�I"t�_�g@0/�Hi�c�+�|��'UC�ژ'�
:�M���q[��z�����D#� n>�e�c�b��6�o^��|FT�e�9�!�2X*��Ga�K0J���BV�j�	ݝm[OZ�E��Ԃ�s�ت�{s=%�����-���A�Q�,�|�����Z�s!xA����r�g^}�~�ϐ�g�)�ޛ��.y�;�ͅ7Pk����Ӏ���G��bs��/��7]�����^'��tS ��c��!�Z�P[0���[V��.����	5��|%�����pNP�7�y$æ�%����a*�����|���X`��^s`�	�f�-����m�e��N�@L�X��o��/�L�Q��?r��_g�	3�ӺX>

����3N�隴�wn0
Q<r-ۛ��|���T���CQ��3�R1��WpO�8!�y��)�D�H���Ԥ�2˫wb�Y���ܞ�ˤ�4m�0j�ޢ7��4��ZiF�%	<>�
1|K*؛�D�sY/.g�ȋ-}A��_)X{��+r�Z\�X�L��#^?���_Uw�����9Ԟ"x�
EN���z^�^�+�'�Dua*�����$�]=M���+S���;8�p0�\(�Q�N��������M^-@RC�h۝(h�s�^�Vi�{[���g�h����h�jE�+��L�#��I\������[#��1�+�7 ĕhB����E��ycPEɑy�K�hA�ݡ��'��&�h"�F.I����$P� �)�2KO����-�O9���|W�CG�q�rUh�?���s��gE7-������Wc�Q��G%6N�(���Օ%��::ES|@�4R�t�4���>j��� @^Y���n)����&itH$��}���npZpc����q��j��90o��7pnS!Av��w����LV�\�6����\	�Su�����hD�`��o۞����Uiu���Z���-[`�!S�G���ܓ}�7
�����1~`~�k5΅������~(r�*M�F�M��b�S�/����X����9�A)�+��&S.����L5�f�I�:
P�����:tf���s��,ժ���+k;� ��h��sr�f�ƍƙ󍺹{8�=V-D}�!J������:e�ô�|�{4�)�G$�y?d (
�����*N�U�nN��''�&3pWڴAl���$�4k����u>��M�%ЧDe�+'Y�}U�N3,��������ړh�����Ns~f1�*$��_%���-u�g��Yer���vƟ�Ne{�v~�wqy1����h�\
/��Ҍd1M#���-�������k/ J֠JR�[��hp�RTQQ� �����dR�� Xt,�]^qy�Q1
��v�KO���X�,�,Vi�1��}#�y !
c��B������!&�U�(��r�W�Hv������t*@N�&�R�k���87*�WT~�i�XX]4��`/fE7���y!���W�w��������K���r�P1�=����P*&��T�I#mg2:I)�����g!�h<RO�|1��4����D;d�M�=7�vO��d&�!�Ĭ2�\	a"L�mz	}H��{]�a�Y|JI�n+�YC���P[�.]��d�B�{��M�����6u[~��-����v�úU]��g����Y��*~Ҋ��Ĵ|*�#�1_� m)�DoҔ�_�S����Q˥R^�s�7���%��"\*c@������Q��S��F�_��Jm�K��7Y��xm+�v#v %���lՕ����'v5�6���}�Ԝܝ�l$=�;<�H���(M��׺���������!QpZp�	ں �c0�!��lb���Ɖ
�b����c5��Qwp�C��r��[g'&28��K�\�TF�}���hc�r��7 2�90�F����g�7���.im_�W�XB������#�@��7��z�k�T:�UAމ���_�+�K�����%��jۿ�hwt�� ���fC�[���T����$
��kv�l�������b⿁C=44�ru%��
{��%�?�4�* ��c1ph�ٴl�^Rc�	9�tI{���cs{_�y�?}k{����X�5�y����d)��ד���hi��\`��`�+�n�V�W��j$C�>�8I���G�>_^��[L��P� �Q�g)g[��w��mGB���������Tv[�>x�M�4�I$Р>�]���'+����R�t��.:��w�-,�5R~7�Dr�^˄�Q������,��?�w���?��S�����s�>^�U����u�q��'�u^�S�
ӈ�=��	^2��B(��S�O
��q����E��器�oh�ȏ�w�\�!�Y���x�<�2��Z��!E�zNm�\��}��Y�pvg� ;��%��/����sӧ��U��<#wWD�d���l=��[�dW�q������7����#_�ii��T߼ñ�� ̹�T��n��q��Nd����	��J�+e��C$BC2ʿ� ��ʧմ#s3� �E��B�RXd���K��K����:Pv�8�Q���jQZ]��xt�Iy�,�hm6��w�:,ZVE�1�(A��aы%��2(<`$����>�9\��n���gF.�r6��&z�j� �pu�I/�E7}���6����Gh�� <��(�5��]eo�Щ�Uߋ�i�����J��(a���9^�[����8����M��k� ��7Z��mELd�Q-�-�q����'�|v+�
тp�B}.� �V����-l��j�KO](�0�X<����q��L�pr�:��4�J���@���p�k�/���1Q�t�Y�F�hֵ4Ԁ��Ku5J��k�OO��G0<7��!�i��e�H)�a2���Ӏ�H#���z���C5a�Ƽ���f��'�Њ�%�����1x�)�v?��S�D*"8��˚9b9US��*�۷
ZР0/`إ��C�)R��\�.����5�`R���`@�|)��F�"�*M;KMg�}~���˩0��Bt�kJ�e3��A����
�4���a����4�D,��-4n6r�<C,#�k����Jy(�_�L�2�v#)@�A�Ɋ^jؖ�0m��7���A�,�G��z3�P�B�s�7����3l��Ԯ����@3�pH+�i��Y+�m�)ڹ2��O�S7�����`f�+F���h��M�����w�v��fz�k�8�� �����E��03[Y�3��K��1��=㇮@b��/}�D�d5-8�ş0p��f�h\�.fN>��#�|��T�Ƞ�L�N��(#�5t�����R!�7D
�*S��(1-z9Z&\Zݺ-I�Zǆ���f��WWC=݃���;}2<D&�!����Α�(��;p��_4�B���T��|>z���WU��������it��餟�[�*~I� �2�;Г�VK�
�f--ۻ����^by�Tʹ��!w�e�88�_ї�����C�z��s���������Z>�O#�(y�%��JX�|���&�jq�������4QCL��ߕǯ�s�ħE~�e��)�x8Z��ޥ�eF"29k��J��^c���w�X�9��<���#wnr[����(�Y��ƶz;��v%?�/�<�rPfh�Z�����1~G��$�
Ǎ�����:*�����^�J�%<�9�\���>�o�~�z}8���������k��|h� ��C�kx�E|7H��k�ʵ�{~l,^K0�����q�J�:�";qL�ŭaW���� �JT�[K�7#��b��C�:�0�q��f5���p�4I^�IӣzO���'�>� c=��d?�{��������=#X���U%��m�%`3O��l^�[��^Ǚ胄�}��М�y[����;?�QN��U �g����@�����9��GH@�aH�ӈ���6�������4�N����!���`̰1�g����������`9�R+3. �͎֓����]ڼsJ�t�!�O����F�|M4���?M�1�4� 3�D2|_�cn�l���uRe�d��L���ǠD�R��fƁ��Q1��?��͕�T;�%#8<�IM��hA8!��oN�]M�WH(T;m�?;��yl��T ��\(^�$�f`��~�Uk)E.�ƅ�X/j��V{c��ǋ�ÿ��	�:��	��;�K�I��f<�ѹ
���h����-¸��b)��*/�������'���ǆ�LYD���X�:�j��Lbc���,�p�����q�1����f���#��l Hk�QRja���E�xX�z����_["DmϬ���P7}R}⇍�8�������ɂ!p�U�DuTJ�����qn�@ǌY�0�$	_�!��BXF�j�z�ӿ/Њ4�� u:���6�
Y��B��MrS0��i�a�]�Y}��s��/�xk���/��/�
�9����M�A`u2�O�X��b�a��H�!N���^�sH�������[,��U~��L���S�Y��g�Y�8��<�ty����@c�2�t�<���+_����4Q����v���D��d�Wn�&Y%}�{�ᗼ�K��v/����|J߮�L�$v_j�����Ʃ��-���
U8h�X�ȳ�U��]��LA>����(lc��Z�w(�Ƶ�eq��P��TR�j�4��O1�V/v���19��rg*}��L׻M�����ԩ�n����v�
"V쯮�1�^q�q��&k�ldC����I�� 6wN�`�*�=&Q.�c�E޳�i�}��� T��yaw}�m��I��)��8�?]�g��I3F��q_^�j�28H�2t�X��1:�n(��[^>#b�D�{��Uۭ�������{�W��gV�q�#��Qv�۫0���ԗ���Ё�Vt��F��ǃCs@6>��0�s
��Č_֥�>�Fg�[��1�(m=JJ��A�k�"�L���SvZK�����/gȇ�c���j��XM�:��@�寢���ǎPW|�%�Zq�S�}c𸠜 ��⯏<)�;�y�![0���;�1鵄pw�C�����ZH|��8��\rܻ�i�`!�-��=�D0�ȋ^��kq��吼N~Tm�d��d̐4�����/=��ڳ��!��kvYT+�䄡�T�"��S�'�پk֞46?�[�G_z��>��ʀ��������e�z��E:VqI��%�^:N~U���w^*O:c鑽��5����C0�(�z��~qe�◓O��ɉ9)�v��/p�ţ1���S%ד��b�����	�� mN��e:K�E%a�v}+)S0��'�7��������|/y�Ӣ&8��#/꠵��sFr\�w��,+@>���X|�IT��x������A2ՈV�5*=�Y�o.�%p�r�Տp�6�[�!I�+��	��7��Y��mڹ$��o' ���uX�3<[����F!}�E��ۥC�QI�4��� �����3CD��\��܌�Q��2�d �<�C�v��[1Q#*f֧�@��7�r��wZ��z�1֯1ʐ���LV���\�JU�H2��O×��ҥ�}s���;F�O��I��2�0c��%��սb=e����8/۪҃�~�nk�csL�y0=<�-aM2b*��#}x�uTRU�}YO"�����1�����߂n�T�^����8��X���<g�(辊]umji�O�6�� P˕�M���n�6��m��2���[HZ��^ZN�?�	�͔]�7�ɴ&�`]}��g��d�4�����֩�a͆Vk��		?'>�z8u�0����`�����	+ �>#����x�����y���y$aɌ�`�ق_J��fOґ���1##3E���¶�����,#
�t˗{T���~Z�[ w������ ��[HW��J�+�\XIΖ���ZT���e�E���� ��2":z��416��h��Ď[��z�%0E#�_47!��"v��n��K��E�:�Z�f��_g��h�1���5d�R}�qK��0C�+ w	'���|գ�7���$��/�3�.��F)j�2R�y9K���}B�����Һ�s4��}xN"D	��:�[E���<Z���h!��:���0���	��0A���(�+#f�'doR�V���� �z8Y�^�⇹�J�v�: �yn*ֿ����bG��>!w�0�Q��t�\�Z�ǗF����#E��U 1�I�mO)b (�������q�\��ۚ��2�c+B���Ih*"�K�����'N��ɔ�>���P� 1V�-<SW��ȱ�į'1�
�hO���� ��W���^�6uI���o���!��a��9�Z��D��[�e�g��56*S\W�^kV1_��~�更�E���̑[L@	��씻��������9��Z�g�ۣ`�!%�'�����q�Cm��̈́?�z����Ό�RXp�ʉ�؀��$?��eW�`2uq�'ͮ��hN�t�U��Q��$Fw`*3�ϒb�`Bض)��+1��mVDg��& O�Z�m���T��#tc"���fY<__ZŜK�G}���z�ˉI�^�$��)�E�D���3^�Qب`��M����]�z�"F�W�Ս�_>/N4�N�5J���&ʗ
����!˜�:%��2�S9����C�G:�ni>�����e��gl�8��s,ɷ,x7���>8�6�Ȏ��7w���� ��wi`E����k$� 
տߣ;�+�oLe��������@�1-�E5����x����{E��zU�}}�%����R	��C&6��`'l_&e��ڧ��|qS�i���C�!��.2
In���:Vס�U��3E�wC���7�H��=Xdp2��ےUaFL����v�.z��������I6�\�Cz0I�kС,���ӡZTAE��GE�g��F3M���\`AX�����.u*j�������.#̶��$a�}��8�4�;�?2r6�s{�i��,��ST�H��h�,���0]�K�����;܊Kx�p�����u�Qs��^���\*X�>�y�@��J�X�p{�d�k�5��)֜�G�@��sH�u�4|hz�mf�Qi�����F�f��s}�iHB�d^P����b�x�fxDul���7q��0��k���8�͌�Obr���̤u�_)P��i|��b,����Y1"�������ǩ�"���U
T��n�#ba���x��d����ɡ����	K��!<C�������������c5�iow(�nw��gF�(ɶ؊��diy�k�_�Ѻ�i�;�t[��*���G���O����C:k7B��G޻�E9J�	'�� �i���(�Wh�r1��qÎ [�S�u����iN,��������1���7d)Dƈë�\h_�e�]���
u�T���D�t����y0�x����KW�0�m@�����Bz�Z9�}��+�`%�	y�P
��:�g�Qݎ�c�~v���L�*�o,�Ơ��c4[7�㶺�g���.z��@w�%�'��_��$X�|�*�=^�X��W��産��<�tW�5-Y������h�G�n�`�9'�B1ȍ���/�5jk�f�u�.��ȬI[L9/����b)��у�����q)�h5ؗ����'�Q���u��d�}MeX8�ƍl�?C
xgр���^�|���R<���S��A�@�p����"�ǒ{�{1���:�?��L�X�E�"����Cc�<,4��8>��(���$��j�ov��Sů����Mc����3M|4KB-.+�&_�n-B�xf�%����L^�e���!R�g��+�ۊWR�=���v=#9<\��S�
ۭC�m��c��O�MG���&���Og���2x��:��B2�M�k�x��������^���� �!R���c���'l���ދ�����o�,MVU���t{�#��
C6��7An6�W,��9P�z��d3����	�MC� W�h�Q!!�Cu���:ԯ�AY�l\���jNÁhp�2��#b]8�ׄ�P$�$~�fw|G��%M���J\��ib1�wC��T��t�iS���9��.1;jE��6&b������Zֶ+_Y�')��H��v��T�Y�b�c%���DU�1���/���If�ٹ� ���ڐ#&���ڊ����d�o@"�9�]�/���AML�+Wuq�lعPP����
Uk�HN
s7��`>�ds,g����K5��8����R����i/�m��; i��e�ŨA݌!n
�IN�ďR�kthLE�P�/���G�q�ڈ�]��HY��`�����V��$���jc���q�O�d;~nG���$k)��ģ��Mأm�g��=�݇�i

��h�`on����mi���k��o��� c�M�h�2�	{��Z�eƁv���3jG��|K;�� __iS��Ƚ��j���D4�H��uqZ����X�P�h4�jOo۽K��Y�{y �"p�C�.k��xZ��u�}�|Ŏ�������#���(����o}���3b��ϣ���O;����7cK�Uj��2�1 �g߰l�\x(𱪼��X��X}�P��?�hy3d���YU�4�v#|FF�煌����w�B΅e�:���.��w����3M�⁙�$�� �"+�2��~÷��������?���g� ���1y���BI��B�|*)ϑU%�=�7�����Nn�AC�Ƌd�֧��Ek���&���g����()S5�Vj��!qm���`@��}
1<$K��l9Q�Ռm���ɦ��-�4�OT��{���"F�FRk�������_�f�n�u�r4���v�㍇Rm�@�ML���R���Zo«��#�B�j�� 1���&�/6���U3^����c@�T+��3ǳ��NM��51ߎg
!Is�0�����e�璈(��}�v�F�իG��W��õv�"_� ���H/t��-&5�c@�<V�
S2X!�qe�>��hA"����h[�~<��h����D��Z61��������_ڦ����ѯ���X�y�(c�)�������A�򢝱&��J9�>4�R�tbǤ�]PO��H������d�B��7}ݴS�B���Cے�����v�[E��?��+������ 8�zirI:���fV
���O�e�͗55��}�,��m���'_p��E���f�T�!|�S�\]1�٘Wi��������9� �|W1��H�fi^;3�#�2	�46�H��|�:�,��0ۗ����~j`������ܰ+�P���.�����Ӂ"��֮w漠H+ya��L��=?���~�������bTsp�HƱV2�}�!.�\M6���ޓ�K�VOJIA=5�C�('K-'hi�{��?�G������A�O��o)c�$�!=h�~��},�nPV�d��dJ�a�E�@����;I�g��N�gU��f���D�A��� 2�ݾ�;����cȘ T�N����k}%'a<���CkfNM`Ԋ���L�%��m-�j��3(%\������\�E�'4�O��_�i~�7:�����2u��		>oA	eG�!�?E�dTB�sf5`����$�p�g�<�4QwׯL��yn��C5�f���RL�o� �NKXee���v�WǙ�b1�P�.8��돭����c�sFLU�z�����������88�£�W�_ӡ��t��*UI��d�:^���s����u��zY\�Z������N��&���|������
/:�
��u,M�D��v�=\���$e-��c;+'��j�ب�ʡ�퉳��!�=vۛZ -5/�8ȿoې�5�t�f�N�Ɯ��-�m�r���c4p9�nQ��K_Xk��e��w�f��/�vbݟ��N����q����>����y�T��� ���3�ܫ:�M
:�a�K�S�4B��G\d�W�o0�~ڟY=��-u�5�(�X�������!+��\hPo�Sk	���GY��8o:��v��)c��>i��&V�wJ�I��p쬵�����@%��h!��c
#�63t�V�8��w�)�O��%4�bg�f��3(腑z�#]�j�s�C�B�oyTo��Zo9�`{���W�_F�p$�.�3;�
��uCsBy҃V�'&y�.��,��Ysfܚ�Y��MN6]P�����8�CF�o2H��o�T�����Q���^h4����u�υ�m� qrHN'X����f��Oqd�[����Pպ�#�q�p�ǭ��}����D��oT�,��2Z ,�.�q�"K��%�ݣ���_P�FmK~��6����dQJ1���֩��b^~?�Dswa����`�!<� I.��t��8��b!��T��xt�I����'��?}���61�p~7[4E��B=�K4�ކ��!y����!Rsku�ڐ�X�QXٔ ��ݵ����F��C+m�U��T�w4�y�j��(h�#BM�Qw)�.��d�k�(l���axH��J������Dǵ��h匹�4n�E�,���q���k������Rl��ݍ8�#�����[�r��c����X9��ﺝ��**ok���9�E��S���W+B���z���ƕ�-�Pv���s���TG"�N�l�����~�.~�i]ڷ��D�������JhX��~Y��i����<;�A��w�1�cF�>��R��?���J�n�M �������z�$�E)U��W�v9�Rͯ\vMbq�h����P1 x�{�o@� ���/~��<e@�L�<�7��	/{�E�V�ܶ�*��a�l3*v�p�fd-g�^:�e���Q���) ����y6&H�ω���e�Ł�T���7���\��$�Z�M��~`��=��s ���&2\Kڳ��F�����:9�yy�C�ȸ��4T�2i��Z����5:�@Q����,�-�;���s9m��Q�nC����n_�%6�b���iy�qs3F�G�@*�H'-}�_��02���͓u�<
d��YǱ���#��>��T\6K�jL�byh��=^k���-�*��d��%�W�a���Ne}e)��`ң� 5b��[H�"���	��EN�{eC=2��=2V]3�����`j;~��X�/���5�	�/�%F���^ KK��Zp�%�z�&�;Ox�� {��sF������S�@	L�"Q]�Z�Ƈ�	�ܯ�4N�!Î=���i�f��נH�m>Nb	?�_R�?�/a�r�n�~UÜ�!֖�0��Ծ���?�AZ�o�����4�d�'478.h�^�;�0n�/�#r�ʽ�GS�r@r�_W�-����T���޷�CJ��G�)��.<����s�7�,�;��x>�m�t~R�[:b;��Y�.��d�H��t.b���T�Q��zcd~��$�����m�n���!�?�.'�p��R�u>���?^ք���Bf�K'���{�<��gB�<l�Տ|M{�
� h��ъ�%�Ns�>�R�2�;�ޗ�.U�����S��Z���_�m���'t�Ǿ6#�O�V��f",�ŌC&2����u/��A��0�-0M���v}��>�8�3����
ѹ&���^��Mj�=�bc�[Hn��9��L���5��<ȗ��:�#�BD�ި��)�nK���L@���	=h��F���/�^]�p�G��E�?��L��b�g!w���i���;�>�<�b³?�D�d�P��p��{�9���"�:�a�M�؊���z���6݈��apQ���P����	�������=}����eI�wO�d׉b���lEk]������7	Oq�ލ��?�ZCwD��u�0�3�~C��Xf9S���Cjƀ���S��B.F�eҺ������#Q�:o�X=���̰��\<σ�9���N��l�2����z@�1���Ül[��HIt�\w��:HS�␠���΢[N;�j鷝�=\@��\�]`���B�NE�v:(�n�"����d���^ܻ駏d|/:�[����i���[��D��-��UD?z��'����x���Ԣ,��,��[{�0����a��Q����==R��%J&�cy��ʽ)x-�o:
��U��1���㧯�
$Q��'��A���[\��{Ԑ�	b�nM�uฯ3#*	5��r`��5�B8�������2�RgC��a��i������Qh�+�M/��_`C�֗��?*�}����PKT¡V6������j���\ӯ�u�h��leo���Ie8�~���S
.T�%�&�&!�n���Q�e�HZԙ���q���Q�lhq�U�RL:E)L'�\w6�ƥ��M[��N��J��F���o�dt�Q�DP}��v� ]��RF@�*6��$���,7�$2�s_#}J�L	g�~�{��� �\�3t��@����0"ꈽ/Y�9%y%wZ�=1�]AN���	#F�Ag_��nV�X*ݐ ����m�{�Pۃ�N6�D���tY��k� ��H颖}:����Ev8�x�H�迳_5&���+l��#>Qi���df�M�,y,<&@Z�d`��ϡ���V�o�Mlh0U�qC��C~lz�n��z���&�}�+a� ��*|�Ѹ��;��7�~	tz�VZ�kN���]���=�b
�>'P^�ߺ�ˍN�p���nVF�8�`j��	�-��-��o�8An̾�f����e�~�eo���1[C/�G&�[��o2�eZ�=:a����4�F4�a� �$�F�{
�ў�U�N�pj�=�B*s?�������qM7���[e��tcU�J_�.ր�z����S8C�D�y1Qڔ�d������0y:��|i
�x��̈�ѓ�&Sv���,D�~����H�!�BHR��7F�nT\s�`_���c�ә�I0a�%cBt�N�Q5�g��O2]�:�J�����uᇝ��d��mj�e �T�����&��(s��! ��Ʀ�8��=���� Q��wOx�ƏX���x�����;ޓC&�Q(��f�c��G��>�r��gN)��*��ցW犰��ev_�]r�U�aBBa�5��N��sj��:��m<!�B����-��6�����,�}��N��F Z-��t�|�BXS�P5)'Q���#?vh��/��F�w2\0�����h�@j��N�Ƞ.,�,�Y6�Y��}�2:3�>�x�G�2G���Xз�&J@�E	��/�Fn�f�}}��=X�)1}^�6rA�|�����ܖ�h�1������{����{���v�5�TTj.�&@|Y^.��G��k�!ը�@HJX�Y'�g�tw7v���#`��J���3�����F�1�1%!��ǇvX
�0���+�z>�u*���X9�^*��s3ʮF���p�<_��ʞ0(��P��zb�?�x��|��4f��F*�(��c)�p��b�3#,�.�K��~Q�F���#�2�k/z���\��L=Rٰ���d���G�6	����lT�q���9!��n\.�� �2ʻo�g���N��J���>��iH3>��پ|d�Pg֛-��a�cA�J{�m���a>m��m�_����H7�_>�K/�e�޹�\��k�
�򕲆4;�s��i���o^�6#��O5֝+�%b�c�| 90� [���XR=i�E���Dkk����/0[wӸ_���0�HC�t��g:mN��sl3�EVX#��Z��)I�u�Mփ�D:���űB�����Cf��s��K�+�>�#"H)��Q,�jz����:��#�%-�K��A�M���7�p��,_���]e,v���8���vQ�M���p<f#p��0�>(��fg��`� �:$�!*�����N�W���7l(��xl�2t�����W�|�ؑ�f���}�B�Z(�By�(��u7mvxg�]�w�[�H���3���n�9�1
Tap�@4��f����P�z�e�3�	2�>U��b?_�d�9���W�h&	��݁T��Wܪu�k4������1�E
ص�׌�]d��#2M��m�>	��>�"�y�+E�
�hYG*�H:�/^��X���"�]�2X���Q�[��t�h�G��k-�`�cľ�
ŭ~$�q���`*�S�7)�߉�� �ع��+��\)���PK�;-G,�A�6�&;_��~���4棇�s�>�h�L��_�ic87c/vc����1�,{Ii�"�\��q���$��+��G��T�>�Q���z*׵x[�tEqO�X�a��ڣ�R˗�Ͳ�x��Q;n��
���?��7D1�V��4�y�
�)x\]HnP���5<�Zn8F?.��<��y5���XF�}>���#�S�fs�w֡Q&�(�u��%���.�vqH�<(F�7I�8�.\���O����������&~��ƫ�6���b���u�Ɨ�V1 n�@6��B(`g�TtO�u埄�}��U+���:�ka���ꇛ���H��z�<*��X}GJ߯���i�R"A�Q�����p�`��2�Ey>� c�%�4v����� k�@~�ڍ��gRh	6N�����f���K���W-ۀ}q(��z(�\S�'eD �E�{<�;�=����p�`�}%{��r�ö��tc�ȍO�#-��6�LńW�^��,��>�2��`��lm^�˰�
�j���C^
�c�~v�J��wJ���V�9��W�w��ã�/� ��f�/�Ї4�W��p��wM�b�UQyq�?�'X#)��J�)%}���ïVT[I�:���2 �~�6x_�ggE�&���IĴep�{k!t��;�	���\�`@TH�R��92�5����}�W#�g�a6�Wn���X�rV��v�0m�3`�?+5�I5x�c@�� ��Gr��,;�'@��FV�;e�ƈ  (�����oej�%��e7Xrwը@"b2���'gI���R�����S5]�
��u��Y���o'?�x���Z�Yƾ�#zGl���Y^��6��:e�roV�]�US�!�
h��mx\����:�k+Sdh��B]�+��/�v�yv>��u ���fvU|f2�e��=��4*ͧ�|�kI_��^r�x��䒞��Z��+�}L�K�q����6.�6���%�\���=�Q����p�v�Y~���%[Kov��� ͚9܉�����!����ޖ�޺ۧ�eZA}7�K, $�����} )���U�� ��B�X��#1�ٖ��Y#�HP�=�Jʻgϙu����B���d��zmu�~��H�GS��]&z�u�p?Gm^O+�/��E��լ�ڸ�n-����)'��������E3��;�5��6�wP�75�2LQ�0/�Gh#�C�_p�#Bj�1�";.����ۿe�YK8UB�ɽ�Q�em��[�� %���D��z+!%�;<�Њ���q����yhT���;t�0�>RdE��)5Ɨ�?e���5ޖK�]�q�?��$����v�h�ѿo'$�$fv�&���Z�^�{=)�u�ɰ8�C�0	6z'*���t��BH�B^�q���{��3�+�3��$QA�Q�G�0�zJ��mu���A'��l��-hӹčǴ�C��r2��!��M�P_� |�A������@Mk�n�y[��k��)�ȵ-�>Bw���9PX2�R�/F�f	��"��ʆ�ٷS�wU�=��`<��q�b �a��������d�����E�=���,�1 �]���g"E\B���l����rJO��mu���1�VwLz33�G�Q����n��:rT�A�l��s���gE#Yh��9��Ļ���B�F"g�0:P���g���4ٴٻ���&-�2��l�)zJӀU��,5$eF���'X�;j�ԍG����}=�G��MdE�x�^��TE*��)�C�6_�^%Ņ2l_J�M҃	�,y�g㚦�l�=:K�LA����*Lqǀ���Y�@������)�=�[K�*���΀����4���n*\3�y�0�d#����Q���͖hT�:�t����-�c��1�a���c�>}a��}u���S;�ך�C}������|����
 ,�H̗��[����0i�%ۢ�A��z�2z����|�Ao�K�u~�'�B;
�CK�| L�j�*���7�O�nܸ��\ E=�$Z���Po��X�����qdHB��{iȿ��il�`u�nZ-�71l��3QR�۲Η�ʱj/�^��X��CJ*0Bc�����	-%jh��5Ǣ����> �]�ˆH
O�(i��!��dM��nSN��&�M���8�@j����o�n �e��A��y�w~/�)���K\���� �V����	�rO~�ڵ�5�3.�0xO���z���e~i�O��K��6e׈
���Q�5�E�X���iU�~3�}�BY������?�z{��yD��nˠ�ؤ*��dV��F����8���] �wO��v�Yx�U��N����1h׫��
z��6i%�C?����b�y �b��