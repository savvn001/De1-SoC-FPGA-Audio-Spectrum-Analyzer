-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Kv7KdKfOSIlGiDGA0Puz/DCZuITjJXvreJO2frrdsT089wiRZKnEDaBbq6fe/W/g1sDPu6nUmEZy
xbdU5U4d9CNgHLfkqbK+66xOA8QbyierGOYs9uySS5Z1LMg6G2O5uEoTb/C8E/o6xzV3n1QHWUYM
xMytx7qXCgLnyDt2yj4A+OVPHbYqjJQ5DslSeR5OyIYhq7KphfxljTwmChZUGAGYw2ThNY4AxHat
uDZy3Jgd1RZXYUVUFc0AXwjEFqk1XypwX0B9zBMIxP2dFERrIl1pgzfDU3cRuLLEnWIAZuPalFHr
tiOopKaF7TDLSJvbJTjm6qPQTV/mDuu0Oz7Gjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
olLoZhVAa2/lO7e3CFbyqGoXA3kXQwixmjKrS7m3ZvZn18sLvUFWM34pA+rJ9A8lisxzZrkJia14
1/4ipyM9rqdGA7HdAKHJjg8Z6MLllMzqupyvMmy1YIhzNxOpO+4CABtv84/eKFZX7W9yl9Hv/H9V
izlOLU6yLq35TEN4qNA4zOJU9MpvZ+EoCocNKcHTLo1M9PHBdw7rCcdVr0X/N8u01drG3baJPGeY
A5yutwKEVgJLAajczPgs5tptwMbzC+ljz9UJqdmniC3up4sL2lqqM8GYi7/DO+F49tntRZ7NtDjd
sPzwJ5paiuqJB4j9Y72PIMHkWavFQi+yXB1OLBoHb2ctHtw8/JU5FFN+1XSOCTSpmGD5GvBVwLMi
98qVE36+tm1N0xYVu28HNTn5PApthAxHErgs9FIjagsQu8lyq6ESGrFwo5n0knbfh/P/Gwzfmq2w
o0dGKGBheZFuxTgDxkXs2F7kO5peeSJjlrkyyxHEuPRvmvbpuwyFcUvOs/dP52C+Qd668Wf0WNQI
9Koojj+Vh2UySVv7qKpcBdzL/yXr/ou3jlvRyXHBgEn5FbroQYMh/2ab8JWRCA8MsrSbOaPq/V5z
a62ie2LW2552bSfjck2AZktZjaYC0IwUi9N81BV8oMjb8/AspO8FtPD4IIgu8MY/b6kFJPwKh7yy
k3voETdqlVz9fPnu+Mp3y5HQ9XQJHT7LZUK6dIw8k9+XLCwfScSqKx23iyRuj5I6E+UrcrvzapYH
PygwmCcRzMPk014lgx+25qgckJOlNzSPp+XvNZVL2Wgdf3FDhEunn2i0Os7L/3aCQIZ8PGMOc9SH
I2zR3kriaNcwx4MTqMfjTKnLhP0gnp/og4z2DvyjP/pT2gCq3P2u5icdJKGXTE2V/mxut6Uy6lm4
lmqyKHk96hQiSrmhKS81+szzcW86SAW8VC6BeR7QvGNs0Ieso371m9siCBkS/vUxYskSSMntkblz
5OBK4XHCQrhPuTbaHMt62600B2jGI5gC3AT0jfxidJLMV7ssaLn+S7QkN31e+zyS7NsSMsWk3Ay0
DIOVfGZPZ/IqhBw1/Wtryb6E/l4USkQuFIXHdDsc9FZD/xRyWRqu2EBun0l53purh8Rj7Vv1YEya
KDIgugT7yYU54HGXQOfrTBLQhtyNdabwKrtpKRBZ/gsPFYD0kufHOv//B2uT4x5+QpWOhBJf9RsN
5LkyCt94cuCdHuA7UCH7+tpgPSCeQ0JrBZkGVzcw7dAMjM93vPP4QDd0N8F7YbNIHG1laenhvwWC
wRKrPWSfajFU/zHRivKlxOfNdCRv/mhr0HQWftvvf/qmMX8WgXbzYelsFSGXcDKWTgZ5JBgZHKTZ
WT13C6Qswh0mf3UHDMfXDabm+h1WYmUGDCXcShPITsrmCtbc7gVx0CIUZrNOyx9DXvOvfPfbiVM5
ov9I7+8CsY1OsF0XGFSkBtRit0sdeea7RgXvYdOH1E6I+2deNiSGet6Jl0KcjWXkUxzXGQ+18SFC
SdKESCnKTDBmGSA55PEF2qMe+SB0a/yXRlUHFDNObquPs+EXIQ1gEepcAsTyMqaMbxwZUvwrHGiT
i51hssf692DQMT3bNQhzOOQniVwl1czkRzgwV+BIJfWdaqqG4pzktX8WHfWeo4pKHestN3fIkE2t
1/Wp52FvFBRR7dZ63OQNtl6EYsIr4JIY0DBesh5XCAP6rulo1NfmroZcC0v3D+jRUnOFcBS8RULv
8Wn7SHYFS/fSSBNVaAyvFCoOGIMAQBg03cayzZAjYkZgjrCPFo9rY/fzXDLL2BdxFojhbmzvWIu8
j65F7az1biILHGe2W4C2dVbF98+xUjgE/Anf45oBOg+2z5GDyyD5rUJoRiBhzkoCUMzoIE4qOopu
sPts5sPDIUb6KBIPL/jDRsS3V4LUf717pPYOc5DoMkN6xRkmH2lERkVaQaNxBPFXLSSKEoBDEvWM
raVo60NxbDC++zteM8Vd/H7NCfIjs2watd+lJS0TjKSVsXZA9LDTqPXR+kPriJBo09VBxPPDCdw0
et3tHfqu+IVbawRW1kroNOT2jrn9e7ftcww/fQ1fJ1Y2Tjwf5yo1H0vHdUUbIyP2NvK0fJyGj2Dx
TzWywzhhqJd+AvQ1m8fnGetV+Czkg8AEz+zvU3ob0n13OsRiQXADtndAGDnKF4Ph2icCYZXra4EA
fmYnZeL1Nco/J+aW6sh4ZzqTm0G0TSHspzmfdaMFsTuoobYc3Ut0w4jPmgNM5YqtTo6PJyHa8/Ft
7OvHAacBq9Yezg8WgXfQ6a1T/ZJ3fT4stFbAh0hBvyb5AYZ3FuWL32n/S1QngcOYOswpIifabY48
rv0DRR+C0s/4gp5j83UV5bARZrVqEUci13p4IiiRfS846HgQY5SMC7zlVn5VwTBvS+g+D2rlTaLg
bx46yh87qyxVYgroE9sh1dp2UemR/bpjLLtv55V/QV8TXBjjl7zn7FOwT3DEyu4Tr1O+Qn3qZluR
0GyCncpZYy0yTghUUu8hnljBXGuoxu8JAApmEy2aYQ7YMtQhqX7PusGudfqmH2N+3fDcBJVVMXiP
ApqZAw+HV/U0hWwRKY1U5bJAw8STYbl+3S194ozFKjkOFC8oMPj8PWsytQEo9LD4AFk+Da5B8kL7
HbiN9oRo6F+gaIHatn+7xfAC4brc1YnOCEeRF55vQtWOTcJICyqA16FQUsVP0stO1NyuNBNPyWjO
WXR0Wl/P17HBBUXnud/gubRpAwpY4G2VwFCwYU/2mSTtSXwzw94xY8IOAveQTJ5D7fgn56gcg+Qb
YiycxO6pHvArHhfYTOaLInMn/K2gWBgofG7stu44iEISOstZZ+Us9qVwhcVLEPzEKpdWj1TPblmo
TDSvwalwHYnjQiL/gkcC8JGrSDWQvbOcVO0UtfxdHeFtqeArk3iPPynBYQdjLBOcONm7+JYlW6uQ
IROZ3JMOxqdFJacwAGRXphboq/Xfg6qVZbr2gUGIusF5Tr2GSDNQENTpJ0SJ2TtzV3Qaau37Ii3a
cnv7Lil2rXQKcOS+lU/DBW1uhT/9U8ZdlpB8NUOxyCXgrWTedOoO1a/CVlSd05dmyuENoWg9pA4G
CRa5c1SObbXyWO+9M0/6ucAqBBdAXLcOCmsayi/9/ytHM4zrAtTUmcuhlFuHnDGKA0GpLWf+X9NB
GT1Op2o/3ONx8G9w9ZU63jjWTQCITvr0h/7DP+hIjlwJ6qeODy+5wM9EiKmTCCZiIbBKlaXRHxLA
jfmlSDzIsnyRP/AQWqYNSbMjFlFdfFgakl9y3dzf4/u/AL+FICIO6UlonuD6TefbPtpKsuLPk3g5
4CgBNYSUDWL35OyRkCqxQnmyMaSeqFqqXp3NehRRPr456C2kXwbrsDWcO3matEreszAbamcX7bnC
MDkkQN4gYakF9w+AaJDEX6cuZcC3JTUHuGdU6XQXxcZ2i2NCsRGzUZ1KXmMyBAoYsYHguQhq2aWZ
YtwtgZkE4xUfYr8U/RV9fUrXJLF5PgpqVPgXvI0N5bg3eZc555m2qkq8fC4j3lHOiSYZRObxZ2Ns
tXBrr15dNinRHYOFHQVBhgolTwEMHISHGVGQdBvEZpCKN3xzDXmObsBpTtNDC8QJNiMsGqjIlZb4
U0ZVpubojD7rw5KTDRT6Ahy4gfMDGVY/xNkmf3063l1xSlEzl/YJvCMNucmzgdU4c0w8iLkfOd58
RvBWr6BnKfyhRDtjfMbwv95RiYlW7vbBZ/Qhb0LYqMpkNYNheeOYRQNHd/OJim45HNCW026d8R5x
ehxo0S6rqAkLqaACHWpbkgZZ8yax82cnTHDmdeg0BYOll07A0cJdv9FPydihsLUfcQVHusuqokXg
ED8UZJ4ZpbzZe68a/6rA0uhLkFlIWT/MKSEZ4Nf3etg6ymRv9iFoiaHJ30TTWCmZjzB/lktX46jo
nCTjqpsm2IYmXIZY+HI7xlH7scoxdh70Bpk59NAWltdpv9oY7j56f5AQINPTUkhu8gGwfEtONJpP
cKkKtaWdPx2VAyogGwaPed+k8Jjif7y868mnyYKu2covyWcuNRhQ8zsUZV3tKXlOhjV0claerNU9
pCWj+h09XFDZofkY2Tyb9KRmbmsu7hRFHiOSfGBaFvtrX76vX8JaJxXsfPkZfKnKLr8ZFHJxhIAB
W9YnVikr+nHnuDfayiP4j/PoU8cgW6DIUUcqKzVKTAhnjfZO4UFIfJ25Ex+IINElmE7jtTLyjSbw
oXPTjvZzYVB4vlXQBGelVo02Ohe4Cnu1DBwuJ2VnlTTU4Ly8jC8oGvyPsbD/tzxX7n7BdxsayMm0
qQj/lUu0bl69F+RVvGTGdEZd5jU/xv8+7AXBdeeAgkfJ8ryF1dNkjzI7G5q3T9JrZVvGnHz4IOB2
1ZfJ5oLb52dqNsd5bv7xwc4TdGt6sdlF6RHxPZxSrYQqGq03dEid+yN7q/Y3kCe3tS2AG0ZhzE9z
7O1h6Z6wOfQhZ+n05hpTkj8sYd2sS2XOO8q0di0jwwbolB110o6duPHePuOiDRLcd/o9XpI8XiRR
ewV85dzw1Yqi22zrbAXELejkWMfaYqJmUTH/KSiFFJSqotNN/ytNN65tzrrbsGWwdDxvpeiFGR/d
TS0qGJ7DtptK6NFucC+9oybzL2/sIMlrzFoYLSRKCiQYzO/uMK015GyJGslclisFgmm5DhCrsUqX
pJdiTqP9HC4WMMMD0/c2oBX8ms/TzfzpQEKomyBPdo8SsKJ11n0/EvhSNiS60WJRSI7p612cvoH9
I1L0+ZMVRYecMqo6+AgB0JD4DzOt8ULHrwVBwGzOYcKUF7YijhQejkHQ9/seHO4Rr3LaZji+zOTx
kmSN3vOpmsYPv6t0gYKS5J56sft1PDB8jvaAif2jYW3Qd+S6S0KXK4P10eIMdXNseWF+RWP6GOzw
e4hiRZIsO8OVc+CC1msD0eao2zw5Cq8UX4KGhXoQaDxYZgMiFzLKhDd9s/BagrvPXqfscU2Sb0/E
wiBLL6PL3LDd81bK2b+eImCfJmnuabKyQ/1G6r6fm2c7nG2fLrqloMIx+79dXl7+OKLGq6ELrGQ1
Pm/urMnP9DZgVXbei3M6h6fZu8EvrlZ140JEljpZcHyrvGw+K0bEJ+JTZSLKWZKwiw8v7mMBbTHC
mwKvp8M8jBl4hMrFegkLKdPjfZjmJQYbJ669Xd5PC8S0jzVutWzKUVtQhV/NBb7vtUV+CgB3QyPX
fuR0YM1hMmXTUp6daLmPhlRHhQ/jjpg0BMrW4FjsRZi8QaWpSkB3UlrbGgdCN4/711zbJWqVXzYB
Rb6IjNbjiTb5RFhyHN/kvipHyWE2WKU/8MI+PZpK1MM0ks794vei69+PEomfjYpHKmoCSHNfAZGp
oxs3EyFJ/DR0a/161Is2eErqdf+mB5Qx5caz6jPK5Mmb69XzvSuZQsdBY73IoZzCB6HiVu7AqRca
wbvzwK82pO0H8gukdrimhYuQGb6AW6GxjVOMLBDLlGXGhUSX7oTbrHySmegDOpoK6RTsrSQf7Whv
6sX9xBuIz6fbmP1wmPbm7S8tx4yHWbms0yz4CvMxcXvlOq3ABA+xXZqMwdBKxoiLPcBoqxAYlDGR
A6KTz7MaiL0qWQ8U9I+9xoEA0rK9mo+Oz8xR3PeH2168uQeCPWZY1SYJax+1nnG2mGsxq5xGkZxd
2rjpXR+dvKOYiCOLx5WOT7/1Fu1+OJqBIeJ2Q8zjoDm0FjKWPT0AIE4vDP+B2s328SE0P9fdbx48
VEuUByx94nJupVYieAcB218pGiMY+Kq20NelmtmMcrT+UaOCgdxkOUnFMqoI1qZJMG8R+Pa6mTf7
CXggtCh0v9Xf3hC6UIhyKFBny1cog/Mgmwdfys5+iPcVVnafvqi20c5Viu4ODr1JbqZehCq9I+EH
UKfxKVtBlK2z8ii3/WQU8ryfX9wLEm/dkGyBeGTJMr3TUW5Yw6C0av6lLBO3LFMgrIK8I//Pi1KW
nHgNx6rD/i1wvssnkQtnbcvPb+V6TpYrhdOVoBCLhi2lTOEKLPVGk5q0Ku8IEPv/NTLCIke3e11y
pqVRVtS0C9jpOIzVGsnAxX+dy9ciJKj8eyWtQoCY3FpsWjaNYIWLNy+0Uq36TLTFD9yTN2c7Cw+J
QRZVRiz+LudPUARW2S36k5oypRvU3a4202v7on3hB/JRh8c47AFypzmjt++1grqCPNWc2ZYA5IwT
zlvBJfKwsm9YXow1KIrAwg53eska1pfp4mwqlkBvyg2WFbd2z7WWEH34nNU+esL/WlyXc02B5N1+
naL6BsK77haiOWRUphPFMvbYDQuRHrWsiCc/6l4KeUeNVREvznRlVDFVDq7GEoZfLnkGtwEXdZ4e
up3/et587SioAhjvc2P4HKEzgZ9Lm82d0LRig4jcWaxBR83ydOAJdKFIT18zGGXyis7d7UTJeaya
4ofhKD1ZDWgW1bQvZTkViXf5CnTdWtRahm/mjz0Xyag9SB2B7hSIi7beKxHBYagQ71NRdFQby9td
TLbW8xJrJWBoTzzAxlOAktXrx2CAj+s7cXnkxUmyYXhj9yVT4XSsMh4VA4eWnh2Q80Y1IVl9u0xd
TEZqgJSYE3lYwucWTSDerBb49zGXxwZvKhIEKNYLnqDqV5rsTVLJf78da+Euse3Ew++6TzGvP2n8
T0tp6F2X9cOD0kiIgeEx2RqJX2zIXWdx817S5plwSpVwVFVr5BxIQFwf+oOcB8Ng+uXc+OVpX1v4
PZTm9kgb+jsIV8TtF/UtIMKGJ5tt9JmTAiSfr7EbJg7aGrLjtq6KQL5JjbH9aMJngh/BOKQpMXSN
2m48l0/WyYORz56E2UwvA9N8NcCkHV2SrHR9uBrB5TOjaJJxAdXiDeWnyO7fhus7TVlkVv8kWlAD
4QfYLwRx75uP4K4KArLQ6RUPCkTFU2Ethi+F5ctCZiRjriL8QUUjqLNJwv21DwslPoB8bK608xq/
8bGN+2xQQJymOg0pzfpjTrkxwrwCOaeZFKmuPA53BuNfYxIyB4wlF5RKOt7Kb5p27RXjmbhy+Q0G
Kc3bSqx0toj7H1H5vGRkeH+U0hVXkINFFOw3cZHkd4YZKEZZby7rJqjWejymOKtvigGtdmIOQu5d
wCFy2rBXNtTmc+PISO0Ep0yzUqVlGe2x3XhDF2g7bvzypgUiLnVfTskzU7M95nonaTao+e2FK0+c
JIsJKWhtsNMxQICnAaKAOVpQkj7DtpahcfZYj01yQjiuIkXLGhHodVj34rDlnPJRRBd193hQRiOn
98a3iXYC3Jzc2XuckEkNkB5yT+Q3qEAv3Wr5yh/6fwBpcGobuCAIrKn832SpWA9MWoh6DN/IHER6
oErip09aIwdQM+rVOkSMt4elm58c+j9/3pScOIRSsZiT4eR7mVW8i6FnZcB89ntNTqzt6pLQputY
I+Kn3m0ZndElCO3R/iNNVNNGSq5J0juOxZi5rVH6AP7OhJ4oYxuuIVmSk4fZs/T4MDEgTShoaUA2
Pc+R+9bmAXMqutcaBxFC1+m2IGYnnvXrkiOFweB1Q+r/lU3BwZ17m8coar6C7W1HYusCtijrRTAe
N+yqpFmwyG3H25+sFT9h2VX0yvsEWlkg8TiVKrBS6Dx7JbIsZNOznqDoIj3ndjvgxvVLEdQrK7GX
itt327ZFiLvjguHerYX1VXp069RIkFoMoEiZhFVKMnRnO6e9WFw445+8opp0eatA88DbdSGlbY/Z
5Emu45rPO9+H/sKYW2bUFW/R3ZNpbfwhBl9Q4rr2IEuowwm9zc7bdgcEN7S7LHlWB23toZ4SFjmL
qBIWwspUSn8eTOWDpKD97PF5Nf2mvwbJAVG07kM5rrlHqvHLgVofxFKBDO9v5lCQ22TOGR8A2dDt
kkNDqWEUPH2/z25su6iPFvkOECPps2b7LlW19bvmR6jZHjr0bj4A93syDeMwwtgR9xhYy05NaFnv
myY+qcu2IyJOXjgfqhgEYoTnMqbu+4zNI/EuS8WkeiLo1oEyvK0sWvSHKoOZpLRbTZIBjuTRt+mB
zCXbXRv5XlG8HhcMDaWKAPgi/eSO3brywGBDwnegPRl6vvChWqUYqPOFsOVYjtG88Yc0W1UEjkCr
As0xI7U3Wmg9DhY1Ea9PwHZxznqVdZe5qy0Z2H/y2WNUtDi2lLrp0mhm8bBBbGpATgRN9zpd3mp/
f76JSkdm0MhTuk9Z4NnOoYHYPzdipiZn76SIOhP8ksbe67N3auugme+mOFocf4Tla0y6WHOYC6hO
7w6OLpKdZC24UVb6lDrZWT/Gu8VlhihTIbsJapBI8C1v7PRqxXMrWZmLW6WRu+ipCwr2y2GYx/1d
G5pYjCUYvmQ3NBTj288FG6/pZOGSu9Lg+AysgZAULUTitz6A0Qhk0cCWsOE+WxU6LTEcnh3imdUA
U7Cq9/BXHMKQO4T7IHFMqLy7qaz4kiIn9vrIFa1J/gWR7Zzppo9qLcQlo1M/gZAs65FlI7zh0zI2
w6/e18DFJ0ErfWOj+QWvphVxC49TQzrorEkyCqF2Y6lSRYsBOl4DV4TVhj3Be04PJWPft78rQkSs
RsAIZGT0kXIliU4RxK8x7KEFAZVWEFhSelxz+pbRttOiVQc9wkiEZN9VDYoTAZD3Bq4ktmqR0J0t
1DXUPlvxfj0EPn9FnI402tWBVfiNDyOg1o0e1G1aKyRhwqGspz1C2b6w0ovDv4q9VXYucfVSU6Ya
0zhzBiavxJXIIWIprIYLZ/0XVmc6PDlEB5YgddN7HUzJkOcgfB5scLE4Qxg9WWYOBww70GMfAzvc
fjfHggI0VQ5XTa0vk86vm2/RRSYI8JPR8M/XJTOCVzknXBjR2DlAEoE1RRJz2GQD9ek+sQ+p3P3J
rscD3cqL/lxIrrGg8qe643cUUKlo7ZLi8JFE6JSCCC9k86KvcN5ME0y47GTPJnO7x7Hn6mTGb1TP
iiCp4mv1Ki3jAfzP1hQna8qgqQ36VYykq+aJEuRokORPywrxdRflD2YDWgypH8pXggykMfgrvAmL
GJUz7HxPSrNpvI9Z8GocSVBY5yzzPPbdT86dnxptm6WpyAECi92CVW2LgkTpWjT4BJoTghX9inYv
12PEaHQujHMhGARj9aH6rGB3hEqTndJNKPZUKFfccPTtovBewvR8FMDk+s+FYu1t5oc7xtvrYZjH
/0k/CTkHzzscdBMfQrqOq66DZ3eaqo/xQUftpA8HBJBKNHZshtGELLMkLJhrjMRHNggDnTkjl1Vx
G4RtmS3puP8c/C5v+sutG5hCSTyN8T8vy+UMR6IZI4+RbAcWkfPN8nhv1AAPxSZhR1gOYcsOCYHf
rpXEqeJ88czrB0FdyJ8KfG/ew4i/9dPnDSm47kkgW9W6qSCZRc6vmIXBVYc+bRjY8iU9A29Ul4ba
1av59xVBHg2AwpQZkABViAZ5YkDb3+k/DRDSlKuAWuhgJZzlZVgIM48FQyT+/JsCFqWSLEwfLO28
9QxiSFczyzUAHMDOuS6wiSpQrvabOjc4ynLJYMVNA2ME0kUAPeWoGw7c0cpLEL8cAFIGCp0fdgaE
yJJ/5vKWnGQvDs+cNpjKLEIBheRYTJfn5159Gh/98VgNItkQH+iTwPaAqfGfaOPKppq5pPbIKenP
/MeYCfj/aCBrgjcykeH5RT/sKtX2u3ichXEs5y3Aj2HiwAgAYJcmbuI29Mfn2F3D3DiL5nl/9KU1
pTi0rvdXUKQq8x3EOLyim+EInfP9KiBssWnz8rzKIlg53HkgFnxydgeCTgnenf+sUT1iKTAup5g1
5tCDBmr8g3W3O0fJBpCK9wjPGxc1tSZPGIG7YlzUggbdk9kjsFJMCbe1VrJ3s9PUJfUxiw/VGpNe
JGy55MNo9KMuid0Awk271EG2ScHQvyq9dc9eMGZryURvPCGka5B7p1ui0SCQibKxnf13dnDEcmRk
ZtSHJU1rC2QDV2xlVwyaoy8xBb+3AaFDId/FIDVmYowDWFuBJZqU/Wps50Me3r448DR9EQEtWyWY
FGAc2DWHanToP8SBOeYa27m8WnVh+1RoHXXUJqeyiJEw6MxceoNFXUeUZ2d3ym1VGrPtfGvS6h1E
mD3bsMYeL3nX/i5LBgKO9xGWzbHb8X3GJGXfurOTNdHMItG6lplOUu3ODAGC4qlCjJ4fddDIYDSN
c6pDQseIjl1uolCNUGYtw2uNho1/O/JiHSiaJmFRMmDtgrysnvJNU+ZYS9OL0404dI9Krk/RoJJx
vMsdrMemZrTnKmf22HIg1YQ0DxUiZuO9GyNk5j2ESGld3lt2iXeicLgplY3dCXWTqsrJc+TX2na8
RBlgE7JVak8zed+TOmgvevQJ1yVk5XLmywbfZMtYIrVew8v+D+mgeMQw7+gTopwAkx63gHIiL4Ti
iWULhNUCF9KKXGqLmbRzZ87XmPSTOutzrilBhyQFKAw9AmeuReMH1I4BC/ymhrFvTfjZiDL+8c+y
ou9BQ6/3NmJIMJA7w4DKAPnSrHD7G5NvOz3TOeJn2o/SoCD48wleyrki03vOfAqoIRF/goPbApbP
fe5rqd7H7mLuK46v5anvoBJpuJjIZlXbh+xrezQ467jYsjRfi7x8zW5ll6izCPXcrXEAQnQbZ7IH
pJojVR+K8/D1vnPKBT/k7nUM11N86vTaRUlCeVSrb7hqX8fQF1kxNeya0qlr3ACGxI+LBPl7bcoH
fvQnuahijI/JF2OAFjlnCkk8GZ+qs1oNbGu1Y5UmkQ1BjRrJXPIjzqxzTh/yIYixgF9JAIhJFOyj
rMru+gjAEQF2hfKy8Zeisji1dNsb5tHwu4kgDoQC3hXf71tBmde+EkSbjmuiDOkVlKVXfZxHxiLy
2oJApIUpnS0onfpLVmgwkBWw0Rgez0U44TJWLhtl07LDF7JSk3GP0JOzwJQ9558YTJg+xbpZAENJ
A5HchIU8k3diGG9R9egs+MmuHXr9rdzi9sfw983LD9O0RxnXsZtoB9UudUJFkLgRNc9YyB7aBvrP
zdA087x1yl4rToL3TZ0AIKXwHNv9nKpYs8Iaap0VXWA0r5j4u1rkIPl37SXSocMdx04tVEJAk916
+0yiAiUTtqRmc7Lmlu+XP8gGBhF3l45PSH+0zgXiw3oQJmPupJDSk6WjeOYqFWBz9w8E/8rbOZUh
4wko+RliGxRmSzK2hJmVEPdgWX2Tl64Fs0uhswr/kQlAWJEymf8T23OfQFfOsfuP0ZzEhl6Fui1v
CUisXWLFkcvptcVnGa3gsKwNgo8L9YZ91GqXPitABplZu8YNcGxevx1KchhTHXTbSxHkFQlIncD0
XZGICJ2uX7G+l6IuLqBnccwEnPzm0GiHmlWGyiYy1VKz0QC7oNno8Kb6+YVveTxJ8IiqBvPT/nus
RfFkjRvpf33OiWqFe9RWRn0ouqiZXUzppDBy0iXeGmmhtD1UTBkIG909DoVAElYvmY+GxUVdnvyB
yMUuWmogIX6Aqr4Ip0SJKp589Kq9SC/YcGcyLM0syTQVjrhwwHYFIpIBzgyRstrZNgN7ZVsmlsRJ
wofHLSvEKqDiUZVmFw8LJ9vAbgXdCBtvEIKQmxqFkcy4HbBAW/oSFD+9kzeQcl6xcgDailZs/wHn
7hsHCZctireO2pjDs/d59LWATvGNIsRN8ErzbqRJZeJrX5Lw1ey1p5n2G1PzUth737Jp61zaYKsx
iYH72/eIXLi10K4uy/dD9G+0EIDAn6CX+Y7NpUWl55ggBbRnfKIjOSwNUelqTDu/THIZE6pGNDls
mBhvhbR06dJPFQX5ZVxFMA4c8jMjo2L3VDEsZiqjAtxvjf+hdLUGVPJ/3RFsai2vlKHZ+q5a8EvV
hmdcGAWhREnxPlgPxAh9SUeICDGXKTftbiBkmgzVjVbTOW5uDdGaCOWD/7zFiDHNns16qLlsztel
gPgCZeQBMPfPmh4WVRBR7rXJPN3t94t7aCxf3i0ePawyXxTDAVfdEjFAUrHGVecAw8kFP5B5Xw9+
fLosvIxS5kyOSDQ+ZhIneU8jAZe1UEnsG605uvCRK3fsJxt6tfekmUwZVmFlP2o5peezJIaPY4Ai
1PgE4jo/qJuQz4+WAHS6m4TU/O7teR84TfwfxJgDe2PtXjWGCuOqLkblczb1lWkmKYFvNDYcw0sX
kyXNjNy5s/NZr2EmjKw/klRonlK9nU5ERPjRQqLa8wRl/wVH3i/eF5UC1Etx45yjoGyd092d25Rb
y7ae/UAyWMbzXBP7QYtcJy1iyjKwPjXuQpdSKe3UwISRxr6wPMIUZYzkssh+a3db1SBLas+s9JSS
kNWzWK64uw/2xi7WtnIGCnknMsS6C602XUK5StS382TlsoDo++VJ2J0/iz9k2KzaGZGVnvVh0NYk
zmUCBpAVAquxI9AwtsRtujSAWLPPnMYQt7ms0Zzfm19d2LBHA0Tl43B+sGU0dOAYXKe29EjQgwGR
boPKWFfwse34sw28u3wfvS8AvXpg/G18IfucTZ/tdAL/Iep0WT7d0LZPtwbDsl+/D7Rz0EF5LJuH
+eHThiA8GY6K4eNusbATHECEM5DkHlsHlYn9wyqcKw8HWdG3XV/K4T1DtvR06ibyVon9J+HxG58q
lniWHM5tBPXoRMGAlyecwEtnHm4ue15oc5E+y7btRvfSzAKMxiUmymP/EFlC03svKcAx/gHKXMuv
BFOe3HRU5iYTeRsM6G2wNLhQzOrv1W5aCzuf0+8C5S2roIGJ7hMaGKgRL1/VutXBu+5xtcyNf8gO
nC4qRQ4RXwLLrOhcn+4MBjUk4zmgl4HbcQnoLrHmmD6cd+ZC6D4QuwyXKiHvlsoNNmsAS05nJIbV
ERM6Xtt4oWMqYCOdqvXlqyH1xRVbEXOXsOm9D7jJNdcA9ZwbwNJE595jywP0CnqxzDs8AWgnG9gX
17TT3VahUOshkIBTcBedXQQmFDjYKRJZtFfjxmg/NUiYXK6sVF6VYo8iV9zxR6fq85HWtOjlLqRC
H85D7rG5ciIVFSpu5JRS1xB4M3UxpPx5evZui41gcjuiyBIpBNrj172S1itylccbhhU7MqvTBQxM
KMlsKyhlAELXDmM9gmSpnsISk9kej2NSepIfCnjJ7Z8U1Rb1uIGbF8fj10WtfSlKFky7ifOkZzzK
AcmBCCYDGDdojqlyfFpd2poiXDY/Z+bwi9HRKj50u/RC+X+fr3MdBuM7FJgXppwveKrGl2Gruo5s
+HnYn2LgUje2w7vBYTTex7WYxx2jpuF9P+qIRE4iMA0Cvm83vCIvb0D1bsBsMvKI4TEEcDPM3U84
BuCRe3kW8vSY9RWIJ7FtEo4V+OxVemNzztc0QJ9ZqSCUyVfgEgrXzus86ghWs4LhMYqLGKa8viM+
c5S5IsRsnTgtLJJ9zLZE23K67Hw9IlJ7OyXvHt30DlEikjtHE9q9GF0xLLIunTehoGD7UV/fSvQt
EcDk2fRWVBRfjeSOE8ZwZUd2xExRkdpM02CHp1BSzGxoeca2AZbmPHmF0IwCFGLBF6vJWlfecsyl
SEfQ1ozNftA19Py2VOFCpwL0czbJKLPcpLXnAAowEekJr+occnUMS6wKNlCzHx8IHV6fxOtXqBO9
5OcngpFfqpOXClOdmLgXBbLi2LPyl/cGV5LK3dEJL5jOlylZ5haGeIDHsjKTLOMvednW4/+t/OEm
JFHZD50MwRo7CA6gMFmSCj7DBgxcjzjq6bliCZ01zy8hXwBwoeO86aO16b5RhFO/MrygXOGLe5pN
i/2x6pzWzS/KStHeRMrKu4r3LZp1rIRyiQBLgZkHu5Cu3BTviGKshb0dwkhMJKUCBWK5DNPDTrhd
/hNAKlFwxFWQuYw0CfItZgl/10g5IE7vA9YIr14wHlMxqhr/5B9gjA/fhptlLzXDoArdd7P2vISO
q4De5ZR6JA7ZsaE9zpjUlsXq+9KWAj62euAOfeP1IlpnroclsMDis+zNJX4w7cFj0qX12JY9nOcK
MIgD+n8enTzo/CRPpMg8K2/hfHCq9v+f8yEKxFceYmsKXrcAzvXC1sRL1wr4Rvq56hwk5XkvgU6S
rQh+ynffpGZqHMaonegK76mO4/eEY4V1p//9TCLntTpwx3ritBryoMVSWCAFT2LSuNR65vc1eMf4
EzqVXyE/WuFeM7eeK5gVK1HXumxDlU6du8gR6H74vnL40L/A1md0SByCYXc1lSghVN2mpwsYzY4X
+YD0KhaaR5YcAScoIsSUfDYFzUJ5192GN5mts63jgIQX6DUIFHBKovNqEDFPQAvapXVsrvykw9pH
Q9vqu+ZQceBL4RvaK9a8EINyy4ezeRczbhoKiarkP/LgqyVpfh2lE687NEHpH1cDuTo26gZa+dPw
iCqypIcMQpSEgyVKtc9JLdxvoGpmeXx2AhET8GhksHBCHeKZ8frptxFVaF8ksavAUs94j6tgIDbf
DTqkTK1sHhnjlU4eTq49yULuFHm/hilWLyskvbzS6C49NuAoYTPS6uFh87XBv3QX7FIrBkQLc0ug
aPgZbnSj+PzYmOwqh0MLNM6EzwDFUDrfGf+pnP9I8vKHS7KfVLec4WoM9NvZwY3WOADZzs9bwnxS
5lDzqakaEY5nx1Awza+8af8qjsJ2GXHKDCHxoqlhOpGnksN0ZkqPUTIwyhnTeW5xy51rP43E24Bk
uCBh9jXqCoqMEtumgS9i9GPh6KJaq+M3rAL40xAgqMfFf7Od+6+zB84h4iPmn6VrMWBi6UmMURRb
rSfjlm9kCXGZOPuYPUOgi6HoqU4p7BPdwUQBYKMhO7uRVQoUANBo61+NnMJt/FW4Pxy1eNjNFh4q
5aZL2wFdl5G/OHkWSXS3vuzb5ClCqtphoQZY8WpVlLikN9KiOof6QZpPR6UD/Dbyob+FFMTi+dUw
1On8XS3+8CXRtHN6snINupX0q9KNgPOVt5sEQQFRgviKwDLbXsS8WNulEwX2fLhPuQNcSl72oPcD
wTH8NNh/iuYIh1Hdq79rf46m6eCSLL6M7qoHog1ZGl15ZvqCxuRGvudqFsM9EhcEDLUdKmcnKtR4
9uQ4NeZC7eT3W4Z4NbOHnoHa86SPNKyxU3MitFMwT2XOnO05ngWvGhFNaLiJCdDPuFvZnGTXyNMr
FpjSVy+SFUtDUFxKM8V1+3If6AKLnU7n5wYgH3Kn8y/vKhgbXgKDV5GwvzeJ152emkIi6gyxQAod
wNjWnxmr/qGDpRIw/2nb1W4MdkmkvaZTD2M9tkYJGaEFaROnPfpZeGb+SzaXE92JGXp2S4eIpCEs
wXgNgz0SitggU4d3uCpAbI7b0zFFOgREt7RLYzQiOwvmois+1w5UmDZaDQ44kt3ZoVNH3A+4oMSp
i88TfjIcwjWYPIpMJeCoI11KeDlTHijo7JGOmCWjzT4L575am0zca+NTpf73GtwNkHsgdfPUj0Nt
5o2sH7R0WopOx4IQ3hoS/JEFyLQEW7FWStppZ0MEo2vyCxaEcFVv7f8ijS1hH1aepKLjoLJs2jbj
ptdjDAM0tWQN4SHteBjrE4au26LEBsl/69jkPfWr8VsrDurQsNzwX27IfN4FpJpdXi9iJyjfCIGH
l+dQLoBinzlEWOBQU/ZzqZB5/r/iHSaeHT6xEkFmSE/QuYfFLICuE8HpWbCATe5v3IK1n6pmQny2
oGXs3l2TnXoE0gvFM3PrUxMaHl8jN/qksbqHkGFcIrnAy30odDkBzIr9FUn2l/M/4oTLiY2whYtK
KACPqDXH1ULHp96z0axUoKsaekmFgP5pS+38yilvuwZ4BtR1PfXEy4xpzxl/40V0ZitoDhd8qS1n
udEyhUUgZii/TJ2RWY129JQe3BgCBrm8b+PK8+/eb3g+wg0r/m+29SiM9t+eQxlGF0oEmyMsRXyk
lUoCqAYIjFqikqoL/rIlszZgQi9r8yWx/fQINM9JIKv2Y828j+FLMxUq20hrfDNqmPM3ozObKL3O
ej8bUf5FkLhlOY9wY9vyFFgOnzirhO1COHt2XlS2PLFCCOuM8xP4mFLtX5wxfxxF3RxSOAuWABWZ
pQVs6f6Mmqm0GAAuG6mXmFzc8OHme+NAcnRUcfKPaEj/J139QbH9k2e9zsxjcrlKEzV2I9ac7eb9
S89I8mqLvVirzUHwneTslc58Z/8EI/bLNUoDDlMteQZPc5lG+tyEIGbAxsVV2KNWDlvYxoHKXwxK
WwFbGF1P43VqSfiDJXBwnn5Q9mACdEVTGLpYFMcXTcNFxrwnfIDSlIU4/OwVTTtSdXhanQv5cKC/
5rNMKvYCIAf+lBvLK7Wv9IQWg3hsDPeB00qkXei64lp8hmgBxRn17WZQw9WuBk6rB5DEqJp3nlJV
RPtYzX5Zry4eZy8c0aF+1wfc1bQI65WX+AH+IvOumZbqDBev8kJyn2RFQ0Q1pReCEqalVIVOB/IR
HGrDll2OS6uCoXsA1E9qDLmVYNGTLgwi60uU5KFfguVgH1tLLGWhckTo/r+o3mmgzXzcJQMm1S9j
u0nmzacD6j8S/ltqbeYo9d7nat5maKF8pWIsw5N6NuTbfochkGM8naVRtHJ/bOULP3N1rqoVoLmT
Pu9pFL1DDu+jVDR24oW4NZEsHj5KshLALIalLB16VuzP1c9CUiKLKTy8aIR/RGKMiQklMLdmRxTt
sPMbZrusfglsqc+h775aEcOfwt1WJ2ZE0339ecnyCC3LJ0u88FiqOCbgi3jve3IdRbPyGTlXmzHA
baQ1I8p0sDO2KLqn7TNacLvbERt9ZEspdbytwI2TJIKCGDQlqOWZFMIBr4TtHdcRFsSuNQmIo29m
e9t+a+/eZAzWBtFLmV+/+PYVOiKiY5EHhJIivtTPSXQMLtVSKlQRFx55Rdv+MtXvczIFbsJr2jfI
ZYAoSAHiooGnCVoclM2M1T7JQr3NoYUPpYc+5R1C5DBPVUeM7m0h3HebpeQ2Kx68GJBFihgwhMFU
+aRaVgybuPuIW6R8onAt/Isa240fSkmcUSrXc6Rj72GeZau7ujZteBQPF80ogNLy9Rpb5o9mpzTf
5/zR/jHF870MmUdPIn//wkohzJw7sxS40tC9TeYI/nFFG+wJFyiDHWwwTgGBcPZsL6wKeT4ghpu0
+SQkiGFepFeJXLxtYMzuzEWzfEowIZeTvDfcfowTgW+OJFtA7M8/F9rzjXPv3Rhg8jVevuEt8idH
GsOfmcRxOMIzW10dAD+WrZkMXGQ1DdtbXegklUQk2yrjf57d4EBgI7Uqp8Lx54osv6Kbms8KjW+s
LAdgnHgksLj09Ugvdk7p54aRHtyGCbI83RMzxW9kod+s0TWXGVLOJH6bBWKdxYdzou4E33l1N5kB
HJ74TXbFPunwOw9UkINEp3Dxugp5VKHQVFh6S+4SdXAWPUwwrNCtyz48AitICqwceRykILECf8sz
YkgESF+iCVe46rGrXwm4qF5h9F6fhE/pf98ENgRc1+iwOc55m6vJgkjER01v0AZR+d6MBD+B0xAH
kveZVBQYfyHXHmSO5+eJLj9Xqs4BX2fS9O72jfBXjvU2GqNsKQ1/uORWDgTbOOAd0MyC+1OTyEjW
oC5AdLcpFM8rfeGYHk9Tp0oUL+TavR3NpC/HcAukySLBZ7Z/WRs1VDO1egwFOBFTBjO9Ck0OGkye
Si/oPe5YvlBnzBgZYoqtkGP6K1OUX6U92pb/XOixolIOXThK/VdtJWbkSZQ1zrtDSMeKmGUnE+HQ
8plAkVXEIMPTE5XU4PPxaCAB3iX+ZytY/ZHiZr+rLZDhisG1qqw0MTgTXP50g2bOa2jJ/hJKnaaw
nY2VVx/OfBfUeBuSRRa2O4JGXtvPRgVRcXBUU9jMPM1j1LRyIukZbZV+GCjthqIIIte1I5W/9mPx
A6TMBe913gafMEGt/sVbatrLgftu5V6bYlMj5bsmsk2XC9qYi/KpNkQHPTmDWG6mERprPfTz/hU/
P7wgIuEEwViistk2nzW87jnka3VdXXxD681LkwPMDGSfoZ1soAXLU31khxQFgbiNSufMN2DYU2ls
xIC4nbG3WR8tdbMjjDIbOsXXJKg5qW9sZ26CeJHOwtNb0EJYi3OP/n7255be5acgiGfcsMY9kBpN
yS200ihusZFCNJRiAqohFB5gOjmCKZXJH/2WpU3t3k7kgTafqJRG10MVfzHWYjW4uzOj5Vl/xu9c
7Y55uk/ALk1NQCMUGXZPvMvhm5LHZLjpSSXzPOL2alrknDFFEHr3Gpj3LiME3+XQ6563MasPrIPl
peuLuQ0KatybK0m0lx2SxKejmBHRWdegMHnT9FXc5ZmOO0QfiH87v8X8e61wxiNgUBdpkwkUvyb3
j+J2RsI3gUDlGjpArfxhqTz0KO925cJSIQAY4OPQdAZiO7c31UWxf1QOs0o5V2X7ZMO1rLLccE/c
YD6svOosR6j7r2QKOnebjIT1D2UxKn8cqAOOXwJm5j9DhuVoYEXwAAfa71+JPGOj+texv33vzjrf
lvP/G9wUbiqxqh31/HHp38CukN46erpbPG6tw2N84V2Udh5BGITgUk/i/YumFyINqBDjgxYNwxvB
h1sqc+nYyY+FIwoeyayJiddmsV8497jD3kj673v0SZmCKHkpYcTLhvhvAIHZjIcA44hH7sQKDJc5
KGvYJTSUlrYksM8y7AkjJ1ly8Mp3j+1tdHvDYIpRGku9f/RKwweXnnOW7OVx6OEvv+G0ruU6wg0U
8XSMdThw9iiwir8xiX3j7GFQwII5s3JaDlkmxZaOuo03JGCVFjmWNbR7XjAyLZllj+q3wEAXpgQ+
4tFFkO46a1qSzY3PVNIYbdJffhx1MZSE+UIxDzPm4peHhiERWvkMfzH6EHr1eBc8mFmIZ8W3LP1s
xtXJ0zQabIYeOmj+KSkmS0Lfx38tniABtACMlrVGK2NfDlAbYveb7Y+aMm5I2rBMpfJQgDSO20R6
5oa0MKWLpSILQvW6y/JTTO4pHXwLNgE0f/OtlGfjqhh885H9MhgLZOS5spxIsvQtYc2hm5g4HW2D
PCPGI4r8vcDB5xz8zOnqM4IQkBpuY58MvDrieRyuRpslV63A8en8v4Sq50v1I9ZR75G8OwWaUHun
/t/LcyDztwBHnSxT+N6ptiPR7sJOAXG2va7DJ7NQeubr/Mxwz5ip1p7YfJvf07Dzt8PFVqERRxef
6Iv5WDFcJI5LukzAQHlEG7xM3Yu/cdM/8lXy3NCV92D2NjbWUVDA9NvVEv20dCuogM2ZZ2dF3LVI
zTHgoc5iNDUayJI10VPZmnpCz1l2HOyjfyGTkW3YblcMkOaMzldxM/W8vSzmJw+MhdRBBQED7Q7x
Wv1r6l7uuKblJ2T6IGWCEgp16HPM52f+gxpDUO2FQtPxfcchotI6NZjHQUrvK+LhzqZd1PnpNiIQ
UR2l0rEk+fWey/e8uMpKxCtqCCSxBND8yjlGU5/tMDJkjMy+5OCuHfMP91IRJozKxOhVEY6kYGjc
oMqLRLLoHGIb+2pEFLKmeMCo0g07qUwI6pSHw7A0TJ1n1gFw6NdP2oa/tqMl6M/BVsIEazAzHADg
h3hIsyJ334fYcHGh1zNUidQHuAaC26+AmxByF5fsFSuTMTfFAAeIdmH6pKGIUq97Jp0irPIU5mrE
MjeqQtwLQp9tVg6lR1wlDMW+JNGAwlrr7Fne6qq9g4raAPCZdiXZsm+vEV91Y0EPiEYslBtZDv+a
258Vu7ZLFxVWnXK47bo24D6n+rhqsx5tnERvLst0VKDyTgB8nWEJjzIO2NhPIp1JOW0GqcGB5kSg
uQtsyKrLv4GN9bUz1axBBamxu14rTqTPik5AJYgW+reOV7LIqMLfe3+p3gvi6lhAJBumDK0R/w1P
KXuc5G/1zn4pkT4JPtae8NGaT1LoDtbnhyr/ix+68qSfTHQyLhCydVah8y7g3pu/l5AHgFk+DHoo
hUonF9j78nCto2/oSBk4jdW3slseAvyUkA1QK0dc/T0B6Ci4defrZad+4ovwtT1UXqSxLbs6dsun
kjCLLVmPJZ8+3Nc/2iHBJEainpawqWxVTVY9uyEEtYaWRCLmRKu34ZomrVXQ3lAiO5rg1CjmfKMn
KzHAff4SNWMXYGryRl8s/t98AVEK7U/hhNdYLC4oPOV79uP1wcBao3cOJUxYPR50jNJrq3yln6EX
whzmlALc5zY/wQCCkOcNkiS1SND6H7aAfZerE9yElLZOmMsebkjeiIwg/WenYDE//8Irxhg662wk
y9dyo6ypfjH2R+iajnayEYCnts+Pix6CFe1dWqj8xmcTX6ku8FPLuqx0ibfrarYDitXa/4URIWDd
F1xhYITBhYje+t8QQIsB3GbRXnPeJ/3mzBk4QM9fsSOTsHiYP0pCb8bzd/ggP/MgVy0KHD5qsaJl
Y6KcnVu6WJYB9s+cM5/P3vuHuN7qmvFQr53ysC3ibjcwf0Cqo6eaxy/XDTd41R5cy6Tqyfgh2O1C
nQhDk8aR/RufbfB1UrPGeMLenHgWJasBclmsTFic6F+tsCb2CEv4O3zM77ghGuYONPT+JE3kvwu5
K9cpXOTG4kXBebrM065nRwTsBbPiBJoJUNxiCnmVVBHUaHU08icNUVxmXqjH1cpT1x1cDBpXx9q2
eWwvs1Sw3LzaHDtftcqhpV3F9xREAJx6RgtmIbkmxt/H+Set2p1rTzclWrd8RiZPEMg9WrKUEgbV
lxOLozf8R2ILfFnf8eIiKqMfvXagW52lVcqpOXdFSKdmURZo+LG1XqFoJNwvXNw7g18Y6CoAbk2b
zm2i4b96pYBHzLeIuoNje0ULaLQGwnMOGgvOdmkd8F2O3jyHC1mjzY/cJCIC7o1tqitJka/g8b4y
0nB1/DZBMdO2ej4r2KoMbFpqX4OHYsxZD84ntZicWKSjNx4CDK21g19VWenaPq3jpvBsryAIoUYe
e9vsP38Hmy0k9R7Bho552zR84DjxqnnNyc9OkNsj16JT8VGrbUiwuT04zUDrM6UFnDvTJ2Ah0rTP
6Ya4R8Dr4RdZQpGbZr5IOJfxs1kTjKt2VtcyxTkHXl4lw4KJP4DByr3RucqBHXgtBkd0JhpmrI6R
rnhpRtKdXn4Q5Ql+Wq/2013EI/4r1qPjPJXoFhk5JtXVMJXSbmGp7hLnGAmz4F7rp6V34fDZ0LgG
0+DVgl5PHZqK5FeRPcclbcp5ptQLR+jyMBHlCR3h72278W1QAao1b6OaKz0HVdcVym2ho3iX+VNN
elDtUFrNxrKJEhVSe6PF5nESnmGW9xXgG9RjIq2Mh7rIUaYUgcuLpnzlgY0wcjdIoCBG8z+QcJSr
rGA3/gM2cWfYyNI+vnkwLlNTAxNgeRrqo7OHvnDBEeNQWIpspkjHq/cKKgwc99+MDJlRWIF1CLVN
VX0DAHJwoudaRVZQdGl3/0BjJkCqe9LA7ECQxTuOWUniCJpPRd7izT4n4OEMHMfF94zOnC33yy5p
JDepCkEa2I0uqxrbfiuevQC7vYJqSp2WUbJP4UJDrIlP0siT325WTRr6JLXq3q6zHteeFnE3R8WM
tcpFU0wfL9R/x+SaEoSqWLseh75AlKVPTv1aiXEtacvN/zcA3Owvihw+tyq96Yck0Jz74Hk+BZ2l
6ohN1PNVYTn8ILd9q7vne6aOt400DjR/7zBlVfvnAcGjyjhEWfC2mFea45YE6Ir5kK4kWmMb8PGx
IiDR4/U/Vjp/XokZpO1EgTi2wRR1nsVSSSG9d6iCgKBrfX23q0bVIRZGPf6w3oRDCQU+4rDK7IzV
fZqdCzs08g62rFshYVi7vMHLKE7XfRjQjn/RiOTwPtMNJKpswH3bsN9QJCvbvlOQ5iWjrsty9Yfb
RQt/6v8j+WwM448ZU1e5pQIzlm4k++BqQSWs0Uxbfn8xDb5z+tk4btEx/lTtm6A1OFqG9P3Jb5kB
5p2/QVgY5z1oOM0ChfTyuv1modDuunqs0Fb2MeN/di7jaePtVbxzeRF6BEl0b9hFV95Htz9OCKTs
7zwqB7zhSyGgtNqEOkXuE9d6Kxs9PaU6cFoqHY9JkfqA5t5qL6tF9laxL0ZvmJvN0ds+AA1v6vh+
YY3DnaokdYkwQnlzxa0YjC1X9ajCzu2BiN15kenbcW+UNx939ruY7u9/qcBNL+qgEA05EKSTPgFr
Qnwk7gnYEcRycWOGIVii1Y0v4gsxW5c3ZTouzWCuxzkUpV30r9A+Q3EIlst9yWNpSQtLmQQGwo61
yCJPfeNiSHsXJJPpxNKL0oihK6jTl6gY1c8ENe+xl1wE/Zke1LGfiU1Sp/6hOTbmmrBipg75X8B1
7FqKeB0XQ06iP0Vqe3a5LWjV4gMJT27w5byYVzQLh01WVzxAHpihRCp/8cjRCytSeQp9XDGaNcTI
xjvhDYZvUTtfDx5xf+NouCtUzLeuKzdwmjQ3MkvIpoAVGbp1YINyMXRDOrbvDNSGZ6G9ZF+czDJq
LqI0xd0dig7oqJPDHceh1RvsAt1KIRr/K5tpdblhVfzYlfWJfvH0C066Y2XCr3jmGU6s+ot7LXGL
ZZkF5mqPmm4XSKTndaGHDy7UMSyaUli6yyGp+oxvB0WrFsMqO41HtNyLaLDrQ77oxZYL6olrsKB5
AqphvSGmbMDqjtle9gttWJ44XpQJ2l0uxTH0lsawTMy3gM2x0SmzKLC8pEOLmEjeDTiAZI8pVj7u
mnHB4kaIv7MjfI6TQefjeYLPytMc3HqZzrHmFloAeJMnI+jhtdc46YzW7z62lj+u75G5JhYzmmdI
ddXm7saIGWRf91RxrIAWzlthjfgkap4cT/hopR/4bE+nCluLLwq8MD+ssegNlTQCpIcZWo1Eww65
fBY1Rf8uvNXD8OlCVN2cpmdlOxasJI5DaHX90v8wOcI1jEXpfLY0C0lAZrGFuzyvN9dLBVpb2kV3
+rVVxf/4mIdsd9pJSCiFI5EEbIV9KM+W3cZkOXbLeN1XPDRiUEFZ78/eYMtDnzbw9awanWOzo53+
KO1+vf/RAsPceTK9VuNzWa7Dv/vPprc78LZAThKT7lxbEgj9CjUwt6wXS1+fEMjZ1FQmGkwEaRHM
ifNek9ZvnDCCjFzG2TmutfKAlNpiGO75ujTqOkgH4qrVHiO56YO6Z15Ibj4jCIvB+nH3/4frFpXH
XNYGmcjZhkvqQnVENR+8rHQnVi1r0fmdIBk5EBjZnNbs3508vuMGPFRSmfR3h9ztseh+Q1IXqieN
kL9BLq4rvzXDQN/OLetvOhU8qLeWPUH8A4GYujldzIx3+jmJMBJKXinK7yhvNBXPEDenZJ9s8RcY
NRHlQWBdFqlBu2HfPkfAUFNSd07x0CaWdBSLRHraI8Jl9/fc5KIYhbT6Z1vu7AMN37lDQDq5Ub1p
spPCBD5EffLJYFFdrjfZImU8zFJ8mYY5qMxSSjRXs3If2YTiKg+m/zOi7hNFqArcMxcdlWtQrbxm
Cj8RHWer8E8+yiIeVw1EjgH4IEVXCL3FijZuk0EOlaVHX+5XjI9x71JDjfRWr/a8yp7bFdr5PcU+
pfSdf6WdVDBSqjDoTQHt5Y+jiJ4OiWDm846hYGFnr4WbwPXgxfU+eS62q+cX250pFLC71IL7ji37
1EwSU154E1/bWlM8eguFcAEAe/vu3v+fv1o3cNer7L4l/bMn57ACCoW0psQkj59HQ3oOQIValDLT
/KSAoZu5fHlWbgFjOrl02IlkomJnrn5JmjCz4zy911SFO1PdWYmPxphLQIP4EkRE4HduB3jxVS/R
k/zk9YKjpwb9dP0DbOKlZmxqeKnf2SHnDCK8hViR9LrHHih/C0+2fePviyLabX16TxeNYrDmGtWB
SiGtJGcsdvmOyTCrjMkW+LwTBE1XrLly8KYODu3HIZ613ZA7BZxGJ6gqmmXj6C/pO9AlqrkY7r67
OTfByk8o1PWHO+KACjn/vIx+AZYR4SnkeA+HCEDPVxWEnQPrgcjWql41xTA9iJeuenrXT9ULCFdw
c75soGwg4hARSTGf2Yop1GPpsCH3bvTmj9zgNwa5WPYvi9/yacKEVbV7sxEihwasNJfMD+UE9D34
dcf5rwvxDJghfZcS53/RMhbLeA3rJeRqjekJ7q5CVARIh8tARkwpB5BZQjQQ8DU3mjv60b3dZao5
JUSsA8GhpGiYgHwcEeSSC4gyNrH7B+MTlyaZcG7ertlX267hZmvosK111LcHNY0gkDKXvnTwhNZv
aGvsrdRAMVogCU2xa2dWb6LFKIrQ3cpgrv/+lEBemcGShd84nzxeRimTKaqJs6s2EsZ2lpsGlnFP
vSm7lw403N+d1//HkCd3eI+ioAqWlp8JHrOy60/jTmrrFcYf7IZtqywYjTUx1SAr0IT62NnMeBqT
MU9uPh/grz7n9sJAL95fiV8EnmH5AOFV3eozFCbiOe412u8RHjheuK7T3a/8BOHrIithsO87eomg
CLvKxeGmKCXVfNXzY3BWv03PWJVHGCB+qAhGEckiH01IAb5JfD6bnHCcElVCt98E4GigK2rX/7He
Xd/FbWulCr8acoTod7k3y4wPnIp7/ak1n5BNDlBoBVtKr3amTuMKkZS3tqgpoKt2XsSmpmywXuk1
12bKo+yw3TycUcSuVDM5D/eWpPIU865km8h0MOdIkpMAPvqbAc8Lvvf1upf/fWcopJqhynpBQ2gJ
IQ9aoNKlBSXZPJdugblkzRFAjL4mbG8MWMvDuFNcXfUwNStWgEzrAb5k8sDl6JYTD2slJbhlJPif
EFleb2F9j+bdmRe3pnaQmfIkzR3MtHjOy/lAc2oBnHiuS2/6YWEucVZYEdzzGixZK+5MbT37QydE
M5WW3E6p6F7P1NFM1D6i/aT4c0ndJDypTQSPtaR7IeWbheV9hct1VGnr8HzxICcmFrWRe1nh3xWK
VGJyCmbp+ORh6ocwUUhzuAxcKM9kx4mWHLby5hkMKA/UfDGUVd+nIk0RYY14y4XJc4O9P68gyZ4P
g39V577fLFhsEMl+rHEriF4GSJ4Ni2xnZEgMiYPHIQYRSoeXCSk97Z2PBqVLGzLiZYWW5Jg4CpuA
91pBlo2briNSp8vwxjvatafjTirUuMRGtIdBUjP6hipB2SE2xNnDU2vuI2RYXdMZ3iklsqJZd6z+
PU2UrXcU2xOEwLisnf3wmV2fWNF3+TemHjmRNwGVrimU3PW2lGzSovuLKidgNBoAJD8djXbKDfxV
KSHl9lqfQ5e/Fb/R/RrYq8Md7CaRYt98aRw20qKYK18gsE50H7qLYxgpkGJBmcrYWZQCyrGpfXLI
an9z79faiKI2h27mgkcl9efdcdOhrhRJRKOgNWjmLgskznToYjRylb0OyXd2y9KaqH1EqWb6+wHY
jJWa16SBhV3LE/0IUIC67O2lvSodMoyNmcO8ccYMmjylqVxVvpZ8tB3YHdh9d2hssvvTvqabNlbC
IKT6jnYo/LgrCH1BXH2LllLikes2UHCSwJrgHoAyBGY3L2Tttf07OaqY5ogUsn+nHmcgdT+XICps
rr+MNTIXFZHNApym0lwbmNwxY5kHd2UBi7CfJggwn7YE2R3W7cOBPiMc9I6XXZfqwEUrwTH9+DiY
pA8R5VoXGC0xeLV3yPgaM6QEfXMkkyZrS3oxkNP7LJM+C8y5oEVXmjKMjFBnm60BwasaJlUAA6GG
mDqg6NMWMgQ5In6LyWdAmpuYMztnQNem6CRQQYPKJIn1dlwC4R761yqus/A/+OUVCCKbuJLXRoyk
AAHJ3T/K/VvLxMxwtY5CpTYe5yTeWxmcB+Wh7g20KUJhu2cHpGD+AaZyB3OwpVP2hFq3wTKmZJbp
Oamg6INs0tFW4OXIEMzsrefboo52JRPNY+bS1xgHTjD6nUxGA6z/QmiN8qyQ8BhhjcEZMujUu/gb
gEERZDEkCD3Kf83IR8H4iTNTdffVbFZs3cCxBck5h+0oo10+mA3QhHdwa8Z7dfNm9KQGQKd7Dbeb
o7DfLYS0NwmeAyzUqulEYAqqZPmxth7xjuUuZFP5qlBCs7JvvsNHRhYENicnYE+Oif9QC7AgZRgA
ubsuo3eSaDLPayo94TsmzWlxK3SeDfXo9QcztdHfdiWfiBxZeaUCWsjX1gJ/GCfP3vm4jb0PW9FG
00POxRhbBgzBnN4GGMyyK+z7up+u/QLf9qnp3UlZFbtJo12XvxIwrzZ2PjHZQbbkAsWaapNTqWLJ
DVsodk94eyqrWWPRt4ty9U59virUwsX0Y/WZsMTBNP3F0h/yJ6A0QjDG8t9EnZY1g3y8VlOku9xz
/ImibFN5LhBpQxs0fT8gjUb8lhy3xVQ9Qqfkh9ciVsJry3D95nAXgL5AfqxIr0/VDiqXPUsvCoVJ
1j+oXekJuaXGBpBb0eqzFZ9xso7/6YR6tvqFq/HOqIZmnrEY7EXfUDjR/zOVxZiVd7OeBdKHyy+L
arznix8YJczoNiKTNyU2O5GAuNkF9+G+lrAH/QC6mCpKd7U/wJBiPrPcfVPHAFaYHHaGpbMwB4ce
iIl7RnYnhBgt1gJcQg2xpjiqvmDC5Uje18+Fw7sgEm2QV6Beta/ORqBG3I2KRCLHXxALiM5PitHA
qUfI4sPnpcDvDx4vAJ5JjUpzD35PxwHdMLpn/xSBG85HyvojdgkesoqzRFEA8LTj9JJgzf6dNAZM
UQInpI4HM//JA7sjyz4+YZWa81j3yJQbbAkyTbMTsPE+PMt19OwcgBKP7pcdM46DXGlCI9LhyLNl
hOkNLkHU1HvSPtAzqLzDTSprjTroxhmILv5SB3TkE9Gaur1iDs0HFeVFhaoBELVrP3NZKR0F85SL
H4ClkxrnfGYb3EPFl8UEz+xGynJLVKTPiBzzlfjpmOnxPKClrNltCNCDkKJVQacxDjI89s9rgS5X
HMW9ljaY2TT/8BfovMh4+PLG71BDuOB889b7TOkcsGCIjpXWrL4pCVrRwm+hh3DcdUy2sdZ+f3RB
PPW48f8XB80/skfDx1jAuZ6YsyFQrBRcIqlCcjMgRRy7OtK8NnWwxIWu+QX3KdfI17ergnRKB2VS
2YHZdy4ErPMPcq16p5M/ww8702fYKbhPNCygArq6o38uTzVDzWOzN4uG/EFFoEqsbsb2KsypLP87
DdbN8oXYgHrxWGrER5LqJOr7uylRuzoWdKT1KbpjIASFreg5gZN12EIqzabaOGylhxriO4F0NBVZ
Gtge7nwNDZK3E3CfPkyZDVY0sxpQdky/VvgWdzguwhVDImvhK4wPJ0cBzkv5G/LbbQGgHljF6Qh9
pHd+3I0Ph/NckL4L0q8PPEE2HyfGxTj5a2KBHJBDShSCXsOagKOmTc9OSyi1lVzgkkKanilz9eUN
Zl+1wUJa3MWvYJgUd0BRYGVN4tS6fXfFEkpIhGcWdbsfsJXyl864C3cfywYZq13cXiW8+CkthENG
O/1PyGZmG8iXRipk3uH1ZC3DOE0bO0cjDHaIe4ZHiJ3sU+AMVb3Nxv8UYi2k5OvfIN4xCKJcxype
XGYkFCRhtIBrGeukVXMUv9VhOWK3riWG8pHUgtq/R793spiksRRzse1lclp8w6S08iR2lDl21QKK
khgKEGuQp7QMj5nTNOG/g8Xu/wnAcEkfclMn1ip/p6lwajckR3s7uOCPGi1XlYH0iGwajTwSBbpO
yCnUniJOWvsqG97zNaJg2yUjRi5/KllZ4Am3ugRE1dO/1nbrbYu8FFvTN/EHsM0wqhU9lOWR/RuL
mDaPRmk2ZjnTuEo/AextlfTNESTu2pSzqAh+gSlGSZonIebN/QSU9ZBZB+oYxEuH3tZUA2XMXqLK
9W+/n8jMZEYD//xGcFGLSmz8wy/OXnaJIVxF5vnhevM3aCwPwZXkPqC3I03+LJOcB1aLlKvZ2U0z
7JjS4UgAy0IXsJucba7ljEC/iAoDWu+7FjRfcCdNPUfjizJBrXU2PDnmnJMw+9o129kEGa7Nd/bY
bvTEUBDg/wNfsBb+wzLT8rfBTzupopiisFLNPLA6N4rGGc/cn1jUWnPkpJkcj6bZaeWgAlT6wbJc
BPdXbDg3gl3NJGZ3kY2Qy0+6qTRgKmVnLiZLSDIIHA7NsdmvqdeGRKYChZrlKJ51DCJ4MZJUW34X
oUj3WqXnaQY2Nn/tV8Xmj4UD8jRWpVorQaCh+PvhKzE4ldPCB4njpkZgsEN/bZMN3CjRKktQKqP3
05RIO1b1Abj3U8WHqUK+ynHEYDEJQEUbbn+nB20Q5c37NktQ4KCkQss+RbSZhWm34h2r6/ik2PS1
NjPG9+X3s5tCRzxOTYiNsLw1oknz9vQQSCL50ODnez4sIXAimuduUXQZJPt523pQHMrMvt1ZUsEU
ijBJVPvhcpFV4Nz3ixf4lH+WBoSpXVgibgTTR46smRMHf1Dkc5AEOlH0dlxIkX9Y4VyD0R/L4rVd
ftDKdmbbtPmb1jrqpTV7t8JCSlRjQi4dBM+JI+DowNmx83p4Lmu2KZ8dToHyqzOKyzePY5nLsF0t
sQfXFHp+lp0b1/NkZPX6jcaQzkL73/CnmCejlLuV77ksz0VAT8C/mT8Q1uzgzdubO+qtbPshr3kK
WfXuwNw8HBUPP+sA6Yq1SKWtFVTGNC/WqT95UqEnT19vgNVTGw151AxIJsCFvSyLLuoKd5BAH4Sf
sJAKqe2W9gHCKS+8xch0dvYTm+c8Mjd7fRUFP5kP9w3DIt3QW3t9orQVtm9fM6dPOWZB1P50IG5x
gT1mnGmEaiQ2pTmpoaNZ4/qOnm9YN1rSiWmfRmTCauY9Z4LD8jdx7Y21N/ga/8mi10yIwGkXAzq8
vl/gYLqjBzwAs08mIzf7sN6qY64iatd6lvzOAlRmXAtl0eN9jY9zuX7zNZ6rMWX5R9i0CS7yFTwk
Vk2ZbaMmfxpsZKUZrdXl0Hq7iqpkDPUWqdBVk4w6aIqNWZcBNjGxv58arTY+tYBfF0iqx14wqYdR
8J7sshpWy8gh9gljmTJEuplq8wNeEAwFMv+CjPJW8qLWgm8s86lZNmqkWwsdRdrnS3FgIS6NqUhK
hDzsid4QFqnYld3wsJsHyzUzKnqiuHeZA8G3B22GVrwMfzaK5InRB4d0oxS/zSGeWcY8b+/+SLPw
hfcUWx28SN6QzBosuA0XdT+Niqg0TCPjRXltiOEw/tNqkLG9XvnFNHEUsEcBXNX37TN4g+G/xa7T
N1rH5eSM8+PWXV6hvjCh1h4ceP3xYMU9BEq0iWTToUnVb/9F9vegtp2upckYfJz5nEmsJVnMNDeu
1XQnuQ87wBhNevkWjglQnwOzgjE54z6IkAQPcLssDGE/g+1oDxduLLzpb4SVb32RWoLsl8cYEQUx
zYSUcaV7GUV46Da4YVrw/3MczjIlswFTJqGpcsQuPJXdTRoM06nBaDiSmfRcnJZBLGopbHQ2/1vR
iJsbIxDwTEKXvwydbucOHQJ+AcdxVPhRMqaAEJZ+UytIVAIHH2IAlh/W2BregpPEjgsiQKr8IkfL
3DlOQQwb0YczZs4Xb8lS9utCf7IBksxD2WK7FIv6ThliOb0AEh1vAdg67Q7k622scmu6i3nVwjUd
QmRwbQVx/mQZkcI0lJihVxfNF/EnOGSPDOZ9MUsKo3uWTwJ3xZWQJeynFrBBJPxWKdDrXzuP+rnB
wGzGxTm3QONZqrLTxJYcl9ElsY6jD1UITM8Gbx3s32zUvIFpQfVLYdird9lzW07VQPEY7Pnv0pAw
1W9Kw+RTDZCaVijwrVJUPKe6xfwYBlLHAFZ/+BMwsOQNf6SlKnt9LmFLLmRbk/Ep6ohDMuDzsboQ
9TBdd+sPG/szkT2t5Z3/6jaOz1jXNg4+eRLVsDfqz1Nxcjl3Xy21U71D4fkl/nH2Q1gZGMSRBCj4
JshJkKjN7+WRn5PPE4dzY0bZiumcDPoasT6wN3Rg1N7PY8RQj8GKB4+Zd/Nx6LiHoVXhmsdsQSXX
JgPiCmgsbVHYTA8h37s0uzjVwmD/qG7Fu6Wbz3qDTJHYTssMlDlJhhjKoQcjqYadXAhEMmnKxCPF
2SewnCuoZrBaMS6bFBrWulRscHcccJtnGAC6BrbwP/XnEHU+Roh+8s0ch7lL2hl7AKAZf5Nxc69L
SSN9Yt9MGJPilYOz1ds6o9XnYQqT6dYs22BnIUVWUsklpOkKEGt/Sp2yP7JgrzLYFtS/dU2mY/Zb
c8iif9tSrB79bGzH68oKavjMclXUrDrTZeF4suXStUSO+WikbcnzTdgC9IlMXCwdaHvtaz5PF/Ss
7hsLu48w5eIUwIXauA0HAWgnrG7LTDPz0IJm75GDlbfXBlrk3QE+hy+mAtywmPu6eAXC7ANrQVBq
YmkQpGgJMbmgsO4shSR2QFQXTJtZAakM/Pnl7OzVv8/sKzYigYsg6DRGkdaYtnUSoP8fRak7PB3G
+sB4UWJTUcL4449AfT7JB+lQtGuXN0DilRky/usPfyg0ZRJR6ECTLk5Fc/AG+m8052UsFZWE/ULE
pYsBwoc3VgKOrdwnNuSEW3nxXLZtl29QpYX/yuhXMVDze1BEC06cAUAmjKnWVjK9N3zv+69BxMEx
kqeGIXiygniMyT+K2QSWV3WoxRHoqUMWrPJt3swrdctY5/qnFznRTym2KybYI9vyJ6Iz5sEzNrq+
HbmuDoILPCi7nP8v3pySrrERABXAFA/QGzVqzv6JZhIagdh0M8H+Xs+p+RmdMZQ13oKdNrGPcs83
aQGT2GjZLrTieX0FSZ2n4+5xZZBA4G3NCJQreKKI3NvLbRvvcjqE2+CiB2XkpJLqqwnGSMmt9Gcc
1PR47jhEMsm+GZMd+y5IJpKvOIv8kw5oh1/w4baIs+Cz8sBZSO3/4EXLsPAIcGZAp5DHZvg9+GTb
zL1q4IUDJ4N0TvV6U6w6CPOESUzGEWDAs1bTVlNibt0bMthF6lwY6Bc2tkpq2ReGN33opg83TO+A
cOIgss8GjRWnDvoc/YctZCSUgTBQPbBPpKTIQ3pyoPyo7d2Mi2ySQFPBanKkUDWioxC6xkF3vsUN
W91WUA2ND1EabGWQvzasdF0pqXNs+szEKJb7cKQY2OuP0v7HEjQ/RJP24RrqnzYIsfdx9oFenDtO
sN0fZXDNSIAB8Z3NUN/qGkc/SpLiotao1nj3QdAgQgvGvEgF58J6AQ1j2C9kmNTzVIsgNzxCY9xv
KGHHYa/kG+68WTvalifrLjZwlHTCUwM2aPx8lYjDh0px7EM3uYoVgtoTwf24YpR5aD5+3nDuh6z5
WaykdfcohpHVfT5iztDzoPM3xv8cTCgnlWoi6gHoiezUDPKHpQV+jgUQZzdUMz6PAWquNhiXEy/K
/zImfolvTtfHj9n/sLzMkYE3rtpNK63E8HhWFhOz4C8YLv8tUnuHYtZ1HwRLoIVW6CKruG0EoKXT
FmKoE7hEi2ja7vbXGwHalMpMh0sR9wIeVSw1pP+boEJyKLnfwk88nyFzxMnmCp3uNWVGZJDu/WUy
TTddNCZGYwGIAPKL69sK/OKrFMtAcbHOEehMm9345kDPu3nwgcfrpUetkWUwqYtVMXagnjdsLmzJ
B3r5x3N37s0wk486pDj7cBa9Gje6WGcWhnreDKofwn0M6ifa76+AU9hMHOih8C3N3Ee3qU0uHy9o
/RgTgcsKpbiojtynuADPHGG7+Shl3RgUDdJRal9qRKSpHdowEl6mTMdGpGwy1LTB2yq4In4B7oKf
dic6NPS6rlHTIutEd9yqhPSVlnKlteXjBN0e1dFyOaaRMcGWEkCdsEfWI73bvHYimvicSrZg0Dip
EYjNhH0l3Oel8qxgSNnBRSOriZ4VdZq+xxL3E5FakEzqGrLJNOsQ2dSUaEs1D0horsgFrM9uDvzg
9PXeSIkdoMdc/8IhV+6kkTrJh/3kSrfbVHRTJZgB6qVz3Rm3O7X7WOyHzPYD70QHXWDVwDmPopvQ
b1ZfUS0Bl+Vl3F4Yj0w4wMPGT91Zu2NWKQEv18rqm88BS9JleCSZfG8HO0+6C78Cfp7bEVtkaysB
R32QDLYeZdn4LYfyfsKJCHvlVjosMb6gJsSthp/R32Z9ksnC48TGQfrt+UbAjAZybDzW/uYRSjRF
9IEVBa+BAQx1pMmc0upd2w8SqnPzPLbAVgRE3HrwyPagaYBqWeT+6wC6XesrO0VoELFbU9pPWnw6
Gq69EA+aIn/m4PPT7pFxJfK+0MASP7Io9PT7Ib4oUEuBEo7PDMYFHHir+A4AAky2GvxGvHOO4I+C
d8fOzVXNqAJo66qZ0ir9+9wYGxrWTzOumAXNZIJcCd94M9DBYwrD0Uu+j/1s8ouSruqOaIvp6Qqr
SNajOwxwAycfj1B6aLfxNgVfaeweq18JVdKQzfGxqAYg7oCH6S2ZDVFYsduBjs6GZ0pi2vC8Zhl5
ik3A2GordbE37kBaHQRHnp6WhXhafTGlvKLs3nnH9Ppd7uY0WtPo1I2s35UUYrKHinaY4n9E331I
Y5beRrIYnkKiJU/3cSzL+1JH7Es7bUFFPAD6+GB/nTIBaQZTc+ultwt9XZy4LmXCsRQGxfkMkKRN
UCk+47oYxWC19UUkw0elV2FErjwciIn3L2I3k0GEzLxCoPfRCMPBGUYVgy2wWW94lTb2pqa3n6JQ
Eizw3q05DYGqwKqNd+b/ZxC2QmSID4z0QTLtHmO8kxauvP3IjKBdmpu2rMQf0gWfszjtX3a3Xp2y
g9UgkdGK8KULjYaSHDNol2/Xb4OwKL5if5bZmFc1GqBBFIhHbspoe7HENglihndxB7ycFeNRDsCt
dfj93CuKKrdhmsvC7EpQeKIM6Yla4zMzcbTIOpneLWX/BuB+yLdvyBzqN5VHugxOqmWicCR+G5+x
4ymzmXMCI3rgP0SZ+VH5TpMMZDB70jsgJ01p8TnK8NiUPQ14Zl8ii7MCPo/+nrDxxRowHPflI5TS
g7m4N8uxnJeFdVFeC4w5LPp46MkkYjdIM9cA8756yvxsAQaO+T/2DygNlZhrsFNr5QwSB6CnHbdq
X6UAkGRO4QLjWWIL4UtaMXuKqM83ZW/7gFvsJ9rIm00hPDxR6Al7fRArynzLzAPikcpR+oVOGPzM
e0LuVdMEBunrXX8pzKg0FtfAnYNi4GrntSnfIAdwyfpjdByXa7g7gLxPYTgvWnrsOfgTNakjkyDU
8j0fcrHJGng5KR7F9MWj6W/Ug3AgisyIODFlKZ+kbtxJlhDjtCfee1lMscyf3RuXkTWPjKUCSMyK
iiBXkG0loTJHQfkjihhgZZ7opCjfwNu2I0WWBMpKU0NvENt7zn6nH5oMoTjKn9vmfrKJHjkuC0CO
XLLLHhwVX9prkYR15hDAU7PxD4OwgsrBIH46927zchUEkvwgguYhRo6XyaCbN2oIYvbStAYoSL4Y
4fl6IuRJkMxGrU+HfZG8vJWKQl9NwLXUTQu/frJ0P5XrJbU1O/vfQP9niXukUoji89YH0ZgVVxZy
TvQtni8/4qAQLNR+8VozePcltca5GIbCBEnIMXukb+uTPXqj9wG75dALT2oY2AlXyu5Pv9uvZ3+Y
lZdwPzhK9ONZPQxa4353Hn6QyK1v0zVG2hkhxIvfB3k49xD+qQMAv/SXv2vHSzmd6oBxjiMupIhg
zfXfbHWjaoAjXnx/Rm/Fh58u90ex0H9OqiNpBeNe/bKBQn+EYLo5rZr1thrjAIb+lKdXYijKveiS
1y0by3gHAXMs8oZ/Vu9zERBgapIMJdazXc1CJILBwmdK+O3rBsj6cb12exuwQQWMaIa80vBqXM72
u/ZCCuBVtAvz1i0QPLkAzgECv3R3IeW9Ir0Lh/P1P5x888RA/mVm6HwPlpij5wDJnmEptfHaKFH2
UJRvSQc4EZt+t7IHHnJ704GXPcQOWfxZsJtFHxI08tlkUT0jCGWVg4+IE15xneMJED80oF8M1DCl
GQmY5B5gILbW7QMorW/PRE7fb8Y+R4eDG0lBHJ0myIkMIfeeOpPQ1IfUupLk5N0S2Ly5H9x/B+Vk
qz9Puc5d32oOu+6hIlw8QxNLMkVFj2QEiZJb0D74Zryw4Crgp/Nxuu3W6meGlPfb5ieWPIjtmFeB
ZgG3GKcx+34OokrcijhjwsirDDamnPOCBcdQ69/1FXrvlwdc4pt7LnKbiGqXbEZcHoTHuEin7r8P
XtZaEXi7MhQkOyIj7o2Eq5RdjIOzkkCOEvjcvv9KK9oVOcJg+Qq3o0xRikvUkHOX22PX3/yFGwNC
SR7aG5t3Z8p+2ImVsOnyS1daMhJQaE139RXotPMVuYIOw+TvSLimCDcvdp+41hAJlEE28+QP/GhE
8+OdBFrxM8q4gF+uocHV9l7k+p3ctOyxcNYvOI1zCBD6kGsFIRGVmSkBejH/FtxOUEvreVhoSj34
xDlP5jMGBptisxLyC63PMjFKLyQWBe+zF9AFnrFcRLq4H6gnTYFsJT6gqsimSA0sxLZDwpW1l3wn
NI0P9kg3ekIBJLy1tR/KAGLyhCUTFnQGegTdcXt04kq76iuKUbINXz+wizkkHVWblgBcvDzZF6n3
Gh/bkJResgkEn3SV7laRHShk+ROIlJWxD6d/fZToZnseA1ECAtmyIozt3u87hnwg5fpdDFC2xXVh
71v5buhAz42R40w4Qv7Y4AgOQGJY5pMU0thQ9k8yKRmWV9X4r8W+1/K6jFDH+GlrB8X12tIcEvhk
DnF1n9GiMODi6+wUftrz7gLadlLyIH/qGDGCYiccXCTnCXkfLQLeAKqdnmdD1fGQHgZ8JvmB8Jmi
ABeR0d5IqVWKY0psPGDSdtSEnzmuRNKEUFD+rXO78i7BycqDjhwlRgpNCkXIR6QxbAAoZT4buN0+
HMJmCGhDM2wIOGlqODxcx6kBlA7nDox06JtOYhSFiSQKQL8RLWZqxp1iOyIoxW+LSpj6dlrL7BLA
2EzEyAewpKeUcEIlfYM7jqsGg5h2iJoNTuWDs25Scqhw1qU/I829L5CHwYvSIgRqPw/fcycWH71S
XHui69SOEG93hympmk0Ss2eJwgioONuD+TgLnuG1RmksBBH19+UkRQK9hiUYRyr6pki674K9Bgwx
ShxvBbDnV9Mu0HXLkU9MQG6ImqzgW9vPgRy64nifynFrWMqOj3sNsS35eKLE4yClnbLHWE3kT0AP
cRjfEffqf7pKeD+WRQy92KSp5TLehscVMHnuKRxZlws41LUv4fvEOKNDAaW3pyFlx1usdLT1YA41
38w1WrNbnQ9qlp3bA3Xi9kUFizjynfbPIJU9xOkygS8vjBVycW1AZtFMsvfqHxHh3QVNmS8+4Ih3
7SGTAVYeWw+KHsNnd8F0v8DNgn/9Hc1cc+Sn8pdsdUHP1duBESI3IGOfVeATLmmG9MP27eydAofk
APzjMDDoy2ntpmxWyTFH6TxHqO/fKB4EklQGsVA+canXxgHd67qb2wtuuQVgoLOtp0Q6YeMk7uF3
7cFNsizA3hFEo+bJ8ll8CoIDd4xy0Yys6QbaRK5ai71IOHzGN+AxL81NEMG03o2U4HlQK94NFAx1
v+Ylj1/U/1TAdL7cwsVYlQTgfx1izl02y5NUQwzwuS4OMT3B1gy+bHnikmrT/I1Vha2QiIfrZERE
lXEvSjHniZ4LOBUPMdnXh+0Kzv7TZzpizGToZ6+bdy/Vb46WLW/S80aooFA4mXB0KPl8HSYcLUCZ
32Ej1sJWq6dVxWcEn0NTbH20/i1rPUA2HttN5gJeztTvziQxVT5ZMqp1ocpGivHCLsxQG6me/T//
cu3nBIVQNpSsdJMwYChrjAowexnyWA33KtP+H/BDrwjwXDKdR0ePkTOGQMG0VncY3h9nwTZF2plP
Nm2PpDZrvig9ma0Tr237aOeNjDMdNKyAGKcDfZl0p8q7UHYSysf7y1lxGCi99P/NKKQDvKuTN6ry
fv4AGP1lU8C1ZvZ1InZxFBkKoGljDG+m59CqaEzJhG5py7y2K/niHYZYrk5YIVyM5wgYK6bJ7ufK
9cxz59sYf6dmnYltMRxXv1Z7knkAbd6DISKLpZfFemLL6qDHLvRU6oF56DYK1+cmPsI8PfYdDwzq
2Nh1hkqyTXgy0f58nbrxIiEMEFtk1sI+s9Ra16qC2NT8lBPxL9HWrrfD5ZHWaiSAnF533oEG/ji0
NEM8kWVCzjGy2YyvmLH+FXireEVX0OTFMliyVYzHO6seS2KmIWMVrEeQ4SiRt6xsT+JHUgrEjDn7
taWbV4BM6+z2LeqMfeXNJBl/IywURr1cGFSVWnA2ahaO5yBxgdwAs3W5aaeamAxAEb9KcjLqnT6b
XOF3TIZu/igI1VwbUtYBOQV7F4ZewKZrG2Vxk5vEitTPsaXlNfzZIPP3Tql1Y/lwpGcISCiyoMSU
zh78Q1dVpQO2QEHxWd0xjdU3hLfFETND8ASWQVAdtV43jUkyBzcbiZtSyXgr2w5lLkEJ+YMOb8b+
cOJ2TTBTr0nRPrh24JrrzBC2IfgOetqFmy47SYhDMmldLpkpchQ/N0kiML6R50sFA2RYIs6dvebn
d+E+LcD+PfVuTMM51MOoETwgAdXTpsBRe8yfIjGPr+/p1f65abyoMsxvYc+HkyuGC6CDz2GPV9Ig
lKSAZDBcJL2ZflSCzyT7HAhQt64bgWXYehwlT2QLtWbMsJVSI713tEdrMEXVEKXErNkuI2/XxpXH
9IfCy/iRnku+hoC/gkj5KFlBiQYQ93AMD9rvPR9UPTwnTwKSkRoky7zhv3Zuo0+va9OEOp6B7Etk
Up83F4uYW+2EHEFffjYIcFXvKdiG85cZufunsaDE/gm/UgoQtiKkbawegVknY8tZD1IZM6WhfAEh
aWABWIGutBB5JeTb1xJsF6C1fBlXLEynUT3Scjf0LcbEWlyWL/pK7sTltuBEAS4j7pUuFEiakse6
hE3l7nkT1eA/sDkQUKNhr3clF/iB325tXKfxLhrlgfbmPCDDUiSFUYrINB6yoe7Ykz34zmaM6AP9
v2cKfQxls6kxtjgn08QoK27SmZYTdAesGAffxq/ofVfvt5/P3Ipo9ZDaR9gO0tEoWB5woJT1Hwt4
yQI/MnMNW3N85+ZZEYuYN0fIKizc9sdXjHSMJ6WlLZmPZOl8V+Q1E01QOp5v9V2NTuMfYWq0Xdge
gAwGM25O+NQYB3oAEjRyxus65NI7BhIQaFSGQn3rpnwTh91D42WlwAbmzhEjwSZ17XX/HGD99O2G
lWImLSSRSfnFEDrhK9EYoJVA6yOuVxBxj48n41GHJwv3bLlU+wffqJp6GSXwEh/8Gcgr3x4GM2KT
3qYxunjrrijLxs76JRx3ThajKs79GCmTMuZ3+rDGROPQIhgPzNPm4YsmQ3wOEfPWXu6+TektND9j
Ov0rp5JoeI86cCd5gGiMqB2dZWbF4FE1okENAnj7PsBP/6Nyxo0HWb8ofrgNmAoCebEDvnrTsN8T
dndGNn9BQ5JRhEjX9grZXcYlfd3f0qQiZxSi/lQiUzgial8s7WEAm3/uoAu/E//sKGlQOyHwsuGM
+SlCISqmOVRuG2+fxiRIYprXq7dbHsXjxAXgTfPbTX4AbBdKPUxNolYaEzPi1cJuCrwf3lReFSff
Wi2GcBbp6joOM290JxaEIUSe4l2vy6sJ5LOqGb6UjAyrrKF/9/eE+KCFexZWTFZWsm8CR1076HpD
BGTY18yYVhynDkbxrhLdt8AEJTH1hHBkseH6xb5Ndt5SdmIbMppAPXuhlm2vK5DcTcLUKS5dzN/q
4R1ygNYu/ZaG8LKJXO796x5TK8ct0okXeaJoGKfOCUBKpKN/dCiRd6oG7/0KDd3tZ17k5+Eamcxs
igYW7r0R8eGbPbXnQm+ScJhU/tk//OTN05PAwIZkkNre+i6pDoderzo93ZtwdV7svXOd88MWKsUi
IYWwqhcuzCs/2iqvZXG41nwGsHZXS5ChnDaxirUVMHQGUGyHsvJ6abujQVWq9zZBhg7+7eZhZ0MT
c+3igZeZI5nhgfXi1eT5YVxUeg/IDCHr6ybSjRx7L770NMTvyOxFJ22MLG1Ok92mi6EbnAcOFdFu
PpHtcfQw46wriTVEVGcR+6kTMczv0iN1pc/GWFqWuS25eaRU1K7hERLcDFVD3creDsaF4Uhv/7xE
1YsTtwlRXTytIxjP5K3riVt5u0xj5nByRwBg1TZRJORPHVQ8zZBv1kVhHnx014CCskdJI3blhm8c
+QoYbacLHP4JzuaJbFYvm82KZeFKJkH3st6m1eGF6x1vdZl0ENoObBuDNQNp8X6vFuFSDHnVEMpg
pz/d+EULga+wPq9PPbZGPnmVWRUGnJyZYasUqXgianByJygREropXAAvGElebfytVMb4yUi43SSJ
whMEiZO7iKmn3R6potswfn+VfEndSAcIFdw9rpcc0R4wkmKjW2LKAsSUAmhuFuQsEO0dCcGD6dOd
eH6KGjhjApge14jssJxvUHDXu0ALvnFgOb6UL/QSzPttqKdIametih4EMJWiRhULi/gSH/FLtBpz
AJ+bZDtCL4N2Ie2wkPpgXGylANZyJKBNkuAAyI4r+npPZRZfUV7nYxKfyCBqjpgCRwXXDnAJx/FD
mpcIn8xKAqTNb48Mi4+mbHdkGsSKbf49TbhICYOh9PuR51qlJC/zmhvXGZypVrJJQsaQ9UD9dx8d
G68VuMrtQkFlg7RjsLAIr1LSoLuM5DukzL9Ml0Vu6HaB4zrtLZRHFepP4RJ06czLDG8Gh1pigONr
Qjn8Kv3Kuyrf8UNkKrylKiScqssIMbENq5K4LTNs4E1GZi7c1LbRkU/c5gqSql+4vt9kuwKK4a5H
q8O9ld9zkvC3ONmwj1VLlevUH2+IadOh4mldkXZkWPnsxJ63IE9WGalnW1EUHPRziBP16Gv+mHGn
eVJFeRtmnw9htwFB/ugcp4fSR1GiRW0c97OPU2rUEIveB4HqnFIB0MI32MUDNFvqwi1UANtDCA3V
sA1NZvZim1acblxhzs/ETyvf6LjHvwAQX2sofpsDKwoWVxcA3VIhBp80ICbdcX1SdvpUINRN5y59
aGN84yDU99Fhnvj57n+BjvnyjNg6NmNYTHB+eDzDgTDxjjIAOwYde1pX9JtJQm3avgGzrPHvXB2m
wPCH00K2anskptmSlivH34Gj3/QRVFD5M0zotfv/q0vDNHZ08p+S7iiMQqmJOYcHZqnLHCrBEkMJ
zC8nD78B3d26XiNlyelljEOD0hNUjZ+0X/GH2tATgoOeYvyHkfeXior84fxMDOUlrGY9aCtYG2aO
vcsb06ROHo3m5KQidOwVVtkrRaZpMFI/RgqOAIhrLdY6mL0kwB8TGLFqDQ1RoR4EQsHrlk+aZjfI
Qj6c+pT/ln7U+VVnZIVl7B7pkCsJwjMqLCOtti7leGLsiHoVjKsp7z152HHxmqy+cBiMmCQ83pda
on9+I/979bDjr3IlZSNU8Uj6xVQry3v59m0vD69xOJUJ1fpAVZM8OFIW9QEFos9iYtsu9VPNB/qr
ONxvbx3fKMLFz50Ou9P0YH2fXQtFbelghC7PMAD5PT5rKOoERIoIDPHUx3qORN6Jr8hH5YORaAJg
a7XUT+rEufa6FfHEdsaHieyLUc8Mu7Len03+VwCY71D39D9WD63dCCjdTlzUfp/l6m4EQxPI+P/g
2+BNETaqq1rZIB/IcGphpKMKaqc0XKBMOaCU5sHEvvCmdw+6olalwJl35Za0enLq0BQIfqPahpCU
Wk8TCSMrCb5wJqCveiZaD90CaiItHLM2peAsGUJHNwC/WbTdPjtHylJVbJdKXXjgOM6DsZsLZtp7
Kc0pztjQDEe3KPtz0VFNfNaro0lo7+cAdCxnRH+25Orry6Obek6xSJXT1zGO0IOYoV9iMXMnwoT9
A7kIVB6Znv37uOH4sqLD9g6wx3w1ajQKBZ7UJ78yIzK2jZ/H/20YU32BL1HiDYrM5ufKuNg8wAkV
qnO9Ki7v4ROhEYwZV54NtX5Mx2AT2DVX/bOI//NNpvsrZBhnMDfPazbHB7vK0DNdzEFouUkgCxoA
Nrs4+MhFGfLISiqndx3AeV/ImPYceMHJPUNHzmyHv3qpIVOU7vQ5nSKvHdI7/S23N6dOfnieCVdt
ae5gae9Bal/9oa0+uyGQF6GaIwAKp4DzA/7T1enkIWTUiKITBEOgyO9y0+ahyKZe+Xhz2oGj/tdu
tOvHHwdsmxcKqLReTI4nGvPaWDB8hpNe5Ewv+vQFMfAGlj6LW5xLf2qZAnAcns8W5xML+WrqxwSk
E9JfBJrxZgDTakqgHUDGXMtTLSWJ53/GkU0CvZy9MVgL5YnvvkjhDJsEf0VqhaSMDNDe/evaHhvC
E9jXoxf/oyJh2povdb4rKW3k72xaLvGx8MUgyeYw3VLaOjpqQkvQoO0W8mobnXPOo/jo2QWapxFg
32ET6j8Wkr6hkJyQ9+0FoyxheKbCp27PfLNJelFSuMv+ycfT0NWRdBfff+R3XL0DcZY2DUOtvQi6
ogKLQeywUaRsGIsdvCgtC7gHGFAxNwa9YOkhvH/lzGboj9WXX84QWWk2+XpbBqMiXTq9oWQdog0O
oYm8ikBne9cJiwb4REcuzdFlFv2fTzEYoUZ9jv5D7pukcSkL7Czvqhehut02EsAhWQTu/cu5C3bO
Lb9nUUPDIev032CTOz+EMH4pzgiOOlEagebcSWDcJ6PHiMulywKRb2LX5ArKMB1OxDL/KXUIf5Mk
nI+zgr1LcbrnyfOBvZayyp3UHtLLOYHd6TNcQDT9h45NKXNZISN9SnOEfKXRt9T/cufCMRp7KDui
AfQCAB/+BzIRerKuKEzWYCdsh3VjmM0tqGsGk7NdfF8qzJaBokbgLW22aU16Vgop8qg3vNt+Psmg
D+cEx5ZuIQQ358o8O9eeir9rjUzLedyWrTOPERCcr9BVOzUCQ9DQ7vCjMuH1EuiVd3qUto/LEKiw
ADQ+hwsh5cNlT0hxPszT3yFTWQUXMIgZOLU+vZsWJ+5S1dYj7TWgZsMcJStqvCvB14wjxMq+W/RA
8WyUSm7WHpoDzqa3xahkzQDQoGxX24edzrAE0Zo9mn1ZjOAD3XGX6HC+HNAzT9qC4+jQJH+8/gEP
MEGfzYPN3RMCze2/Rh9mav98Q927ELnSduw9UIsXMjULDeinNx2F30nN20d0c8QPJsjCWXnkDCff
ACbPIz4rHrcEJm2bOQaoXjMGYaVBqH8lheAvCU1jBdJStgarIEATyUYA6wevlWSZsUsGwbc+kN6t
zegVQzvfE43k1jz36YpWVJ8PryX8cROoNLb0usZtQrASzZdcx+v1O7tcuo6UAAOF5PTg7EqGsr0u
PztJDLP3Vata81YFacg/1tGubrCgak34a+l2rgHMAVUaqNCYTu8++O2E6QD1K2CUD3pSZDeP2u5a
Z7NwzdWfNFf1RmBvzd5yX63E4lPQvLCU0J+FRh4aZTichJuNQtdhhNC851IIkaqdS+MV7+RuhcFR
f4UnoRU2IU2pUZBS+E0vCZ6jYRhShB3IBirXF7R1E/W6tZ4Nq7yxSqBboi0gw7lZ3CWr8ZKtnb+r
TQWG3MzlLlu8e01PaU6CTisDyzmNu/FCIokQ+RdKwUE7fzf29LwoasdvRoB6J31HASlFKLWyxDBq
Q8K/2OIw/uJocM535ielmeFMzSNUSMAu4HoG7Phd1xGfgS9CffrdfRRzcU35VkEVIE4H+ojt9m5y
4KeJ1oQ3bsMOXHK8XBJ0dUsS38xesdcq3BDagTklF4jTUDre7AnfUrcntNf4FRl/pHVemTcfRFRk
xTZoDR64Eb4Oo7wfB3mrgqP1d1LBCrubhLwta2J+B3uyMucxvKYZxHu21/AC3XJ8BWjDpw06Pyxt
qSBHw04+yImY5fmq/F1P8G9jh2QLckfAuav9ZkfTBRul/FsWOe3T0oOB8s91YqJg0Q5mXyvy3u1M
lQdOcfG839N5trxzyO1yH66fgHvCWIv8agevoco86tob30C6/PARbaQ0iLJ9os3rC9Hvd4zGqc9c
wZz7TD6jjP9xgc4Et3nvPqlwCN8vW3FZm27o6YBBOyEqO8Cx6kxtMCi4ZR27RoSGaaVvV0d9KG4o
sWKnhouZnAN5rBJ2rMm84AVix9O0/1Y/+2b7ygFRFSziSysXSF6D/H+qMhSZL+Xh906SJklviixc
tLQNkh2vq4US3nQXydR8SnvYZj5o5alceJY3mw44hkJ71AFQBWPb9PN2CNYhIkhky1ObkKlUeFAv
3xBec+4SOYXGEQawy7bhct6Z+We/7dR4EyDes9CnRQGdtIXUVDBBkuY3DalSKTQSXYrMC0LYKL42
BEJS7AdgDOva9peboYlLEsBdvrkuc/e33efsf074rBzJXRF+t9uHBCiPfzhfbcP3MEwXq5+QPB7d
6jBft1WJJJSkvk+YmUV8QNOpP5+Z3sCOj3vM3RdXn1ZA3Aih7fSGVavnfi7mMbcpDHsNzG4l/RTE
ZFPDa8xep4inDW0Xw0G0JdibDLb8b+QBQi1VSgsHtWtdo9DhrFVjzcZQm56YCRIQDxv3cwjReBam
ZDDJGo9ojAoKA+MFDCV8Tce2NOMEbkQvJuG7cuA6kaW/Kme7sx5S4rwuVvVABl5SxoCRhFhww/wV
QIT2/J2cDMjYibSGR/SGYuucR87JDPNZOvmZ8QVE9A2O/WdBmvLM0ft/irQ3LAqPAnuI8POX8WFN
FaLwMFof4WZPpdXY24xHNhZeT1ruOjeSDgY7+fwgQac9yDKy86bH59tBEZL7x02DlM51GW29kC4K
VcIDV2iuirmejQB9Gy+fBGjt+pJcnAugo6VoGrXinzFmU9bq8WGHAzso6/0SApFcUYiFZgdMW2dS
cmYpz/sLjCqLTk0yRpkPo7JHSyaMlZv8L5/pvh0PzO7ZLTBnDBTMsBUaqHggMfcWIw+/s4Wi9OuB
X2dm3YfcfTYSRg632FE8wE4e9QY5WopdSa9UWy3vvBfpYBc4HmHGOsaQ4DsNNItnuDTI+ieF/oJB
9Ldb0nyXaMe5f2ng96areZlACG5f0dd7lKcXutr81nQhSzEYlIZzh6iHO3znX9u8ElJGRx++aidS
indV3uCAVG49vOkW5u7hIlD6CMGx08uX9cyV/TVr9nVIC7Fi48y6bPdqpHrAVJZ6tfmvFKRU3UV/
lC7Cszki+R5arO3+A7OGQ/NkGtbWpXdEvHNA6NRz6OSAqlINmh5YYs8VHTQnZmwXf0nRt1oFBG17
088TJxgq1wcxw4FPXlpo1HwCRoz7opx0rIBct8EnUTCF4h4vmTUyLP8ghn5tfxWY0c7Btx7hnkQM
D2O9w4HIdYvc/k+SG/GZgAX0ZLE3eVXsaqV1zkF2FdIDUjAyAirUtZUgDt3O7oRxoh/7AmtO3t7+
msSGQlCTxFI2lN/FKBv0kBme8sWRCyA3S0/J7pI4OquFpsPoc/q4ThTci1BZ4XUWH73YtYxFLlvp
bGZThEsV0WCtoKoMVDUrlxHdU1y/zMyvyF1+hakpAvxb1b5DJyHzOk7BUymCkbrUUYVCDtDSErZv
h+QcnoUL1RPYTWbF2iwYdn9bAO0Z9vW63ZKleWIHZBVi9g39BjW30My+2k3ywwZTzHSOnTF+sn6G
1mumezn4+QKWK+4NT9wftYVA6D+4+RYCOojghzXfAIkx404Qh/vMjXX16zHLw2fM/XiWMjd/nVmY
dwLWYVoX7eSzlJ5Jq9Ik0n7x9F31Fj9Gxxaj37xgEZaoxB6nm/zmt7yEV9vaiXpE7i3vdp1CqLau
VwkREpQNERjzN7ZeL7+XaxiKaatIyL2uZv5GNaGQPE9LSd0jv+BRFlEeTtOxD11PhckFgO3eCroh
ENqqMbReucvbNZH8pxCjTSxns04Lgl66aORS+hOlnTzlBbR3Tl4N6AxbK2a3YAYtxLtLAiJ+28zG
/Xf3lValPPitkuCS3bOPOxDNG1vBATElsLA7jxNKgjqAJw7svz1nv7lHVRHgHUSqA05QgPBPsI/K
4xgorONhbWM4SgvQ0WVNTAI4CrH5JM/Nwl3Rpg23y45IOLmcFxQ1bbbXHZY0H3x5gmN0pNft5bWd
hdtWVkeyt/0j+yeRCobeEqoQJ3tFMG6NoKncZgfMHQe3j1XLh/08ptLZRy4QC2V948BtkjBs9U5P
j/jZQgw+sgh2GpjN7jqkPpz4u5Wy+ElC5wnmgi1aq/N8YogF1KHmaZn+iAcdq14nyR74k98OGRtf
PPYt1oRSKvjy7UrL8WiByH3didIk+SbrQ2D7OPT/xT3fBCUEJEjT9MiMtyvFCgvCaHOWUerctx3E
Tmpnjz6UBeefYhC8twVemeOUOjENRbzKLsPIHoeo82mpKi7yMaTEjUc7tALGnagNQmXhvS0H2pcI
cDNKr/qGAOCf3q2qLxc4SDLVmdISgK4vMi8K9y71A6oqhah58tW/oBAdf0BHnSJTvq7NYNZjl9if
mrDahzLoEUrpzVJWeMScACtVkgxyRzIVv4lCJpZatQw5dkrHkWBcwZpX6HS81FRZA8VCPJTS+zaw
0i/H8NErKy/0Cn9OOU+SDQVn6W7Nf1HYPKQw3qTLx9iK9YZfwdYtvPm7WYX0PlJzQ2boHeF1vcHU
fHzGiEXe72/j6mJbBdi9MCgo2LHu7/147OVocY0dg+V3M1Iy58iPTC4GqqDAFrwwdGbhEYeKMzsw
EymqJ/QWn+ZwnG1M5bnrBOEOBFq79VNRSFwSDhDk5uQYfNa+YfHF2VDPsV18hQuMRuPaydqchtBq
+59c6TRbsMxz7A8r2n39n99XEh5WuuXcWB5poO2lmcjbO7j3/hFCyncOqkHacCevBifUn0K2boqn
h3++Xaq3kV6YBfIKnpFdR80RwUv/5KqVgGCsqqCQRkwwGDKvQqQ5P6D84p0JJZyt8OHzmR99Mugy
hC+ryDqUdrxpWWvONTs4O3OvEWnWNOtcV/3zx6ZGVVWwFykyYx5jmeVBFCeP+1mL1OS2sj6IAeJ1
l6Ao36HZo4gGB3/VWMg67SW6QQK72eRY0Qkl55f3Gc9AcAcndAYEjRn6ANAgbBYqQWOjq1Kq2UY5
+a/UxbNSchFTtGzTYRI3cEVqkV4bFQxHhXhXc1AWbKd56KVsepexXspoznO97s4YqdN/9QvV3HDL
TZ+bAHK5OmKeGR+z8rjfA/7MOQbdUTFuubG9TEoFZZQtBA66bXfgP7LM2Rp/bFo/l09jwY+RW1dY
tdqwiJZycgwED5EE9NehFJuwlKMdMfLC9TJ7UsBfVaFoGQPseaxfZoxEs0aZyBRPQHlsBtrWNAmW
ZkZZp58RgpOARMNpinVZhFcMvhXfCOIObJ3zBZlNyRkm8xARJWSViOJ6HBaWgjGvQCMPG9PJi/YI
tGckIwnrdv79B2FGWYDXLSjlRNHPiwDNu6pyHuBnGx+4kyvHN0Ax9uY6HwMnwwUNIBxZK/gKlVfr
spEYqnk3lSDEMQBempfkSCX6gTD/z2ygpacHx+o02ep37JVox3eJdwvP0ACDnXj+ZATXTNN0xZev
N/enJeifIoxJ7Hn3m23cEdgVhS5mVWhug4Jp8LMvj0GLpkrP5e5CWpPQiH+iU3W1aVQFK+04Jss4
yhD2TcMqyfsLmEggGA2dwWdWgSbZyI9Liy2MTbeQRnovC2NUEVyFl4VIrmVB9U0EhCiT5z8/k/cl
8m+viNFuT3dGeDytIsL+REIuBs0dw/p9e7IiUPlOV2qbhmNJYRCaqkO78AfQQwLQeXUKKwY1dUpQ
Bo7D2OO/vKuroDO0R0/Dqcyj4Jwzf/WC7i8araKc8hnwIzgiHZMoOb+prNvMz+2b91Tx0/nKqQGK
jS0XydlbDmV2OFeVGTlrjNszBg6ecpyv/bVKHVFrsVKoRw9BIZ+NtTZAGe2TH87NtpmU2Ig/uZqh
SYk3HR6nvThsaJ5B7DW2fFJGsnG24aU1xV3213Kdw76VzQ/vnNQ3wwv5zd2mtNhFXkC6dXjnUXeX
McqiQZElS2Gx7PMhh3HXZvi3kGIos4v3EI8idmSuSi/lvm283X1JTJMUDFddWiwK2+a0tic47z5c
M4UUuv1R4c8A/R4uLesnzJdDQdjryf0IuqJNRRIjmGrgrPBRg164JXCtjeKyoOjLeL9V9utZni1K
t4BltCY8ApZnQveCRD+H/LS+02rW0ecvQfTl/fu+CdauKUnnmmCYRE++9umhVYYrn2kPuyZx8J+W
zmET2b48BsjC+tZOaZwGWK7sRrwRRnFTyE9UBalFLLBBwE6RaiO31EUBeP+8RTgLRbLH7SEBc3Mg
M393iJQE/qWyPrhz3/amr4rd6z81F3JfNX1ecsBirP3zVdY/OBSwqxpOSH/GLyoR1LiR/Jsj2TYc
QNBwnb8i6XngKFxCOxfl6bSzoF4qsY/VkRUlwuwKKiao7FS18ErHKFi8yOCNsppsqdjogTvK2uRC
0pMXjWBWAX8GJTYMK5691o/MIp56A478e6tZgpCuWZqCTFP/pLHnhTNws2QqFr38To9pNulkCc7w
5jPnTu9lrO1epHb5x5zSg9ceBaXIAxuz3m0vnWjPe4yOHyMwbbR1D34V9bNslFmKc67U0jgJJo/0
gKkOxqcs0a4xIqP8vWCiLRGK6n9SKIJC+De0uHgYgrrZMIIIjTAWYWQ6l27lBBRicOBnEe9CgXDg
IHofLUb3YAKNAzqSVmo/TYo7c44++yx+xsmbw7dFWXPUrrWZD3Qiwpkfs5xAh1Y5BroaVfU67TKP
tR6C/Sxk6iH8Mx8Qc7Nid3JnRO+PRxkd3GUD4OMBt8GOTeyFA2zFT8yxtGl1k7oWERxTVjzu7dkO
9qhgAhGM5e3ZhkkT18eSP2N49ay/gPaR9DaMGkK+RzjYVS84v+qGBnev6yGmGhxiyOk++L/XG0xd
2tZpNg/j3f/l+1tWluy++gk11FjOMdbAqsY4DekKSk4r8nPtE+3QjKGjf0ziow9HCWMz1copbwVm
OwSioKDbc4BawNGT3+7FJWtMnc/NX/RHFkt10rNRu6kCIhKEddm7EY8xOZetosSl6Ufm8+2kPQuJ
eXIURztomjh7+9FDm6lBzM+2dDm/Aza8682yukGYao5iV28H/Odl8UQVb59I98jisLnBElRmDNHc
3nrzBgs3FxjogZOt6F2Vi6nnDgCOYewhQoC3mjmXQKRjnr0/by/oNJJeKDfONKdAupOyAxDLFXto
jRIQ/512W9c4owamDI71WtOnet0qLdnkhRqcMw9+AcNX4U3EKIofXOvnpEaZgXSil2s5vWpuJfUU
6QbmT+9Hs8HypcZY57jdv2TH6sok+q2XCPOjNL4MrM2i/UYwJJv7HxeJFf/5bjIqo96PNdJ5Nig4
VSsh6J8PlpRM7+TLXuUMB21Q5YAVMGs3O12OkkyC36kNQ6p/7ZMG3lruFWhkcRFMYcFpRuBJchKE
znVmkonj8JeJszl2Go1oMqTe7PQawap1UMK5gFsX5AaS1v8C+6Ff248eWkwLRrjFK3oHd9ycoSMi
oO9ToEnBm7P70qfKcUTfhZKrrAzX3rebis8YhE5aaMqSlRbFbZZs9jTPA/jtzQjhP5JBXwJbrT9S
R4pUMxB4GHsEvlddqUYyA6QhkdWlLSOj8NGDsGMJdsejFWYQS1N7Y0NY56iTbDFbea/g57lfRrvx
fIoUvdG2ynLAcbnbUX09evJNIM0EgPJjEljgwmLBX7CJUirt5ulPNkro2Oaz4B8Fr/Vd+2kv2Qs9
ahh0qWEifMQntBZ9krMp9fdjEMrd9zLxMvobz+o0sHG11WVGWzspWBIgLmcQwqbcAfHVKOEmm2Ac
GuhRdISGhmRL3wMBgtmYb6M0n9iqlS/dmmChgqks6GLSJNnzrT2EPQzjQMX0Lyeee/yy+pbt0/sz
qtfEBEtTPlrqVfw39Fm67lldRWqHcmVGMG1C0Ezr9BQkDuM8n2RzUdZSZaltNR+d3qzotjr9EYMe
TU/ocL9+hLY6KCvl9tWSdOOrXq7kN/2aY1Ka2gHZD7Ky6ngnLuGhIrIWWHxkizIxyi1cs7D3cwbW
toka1DBcdTe8ycAe/bQ6FAPndIFhmZRYUdaM/lE+JqnwJLoYYIINwDnpxRz7yh8NDbCFYQZvJDYU
UeG+Va1bZXgq5ddzuA3a8kwgx3X0ebl29XEkxNuGDTuwnuSXx73zRRkxppBARvMo2ENRKNSMjUSf
LwGMjIFBJSe69m167egQbO3h+ReVuMEI+95aIBwL8rZNbvthJxdPEKAWsQ/KWnTzv4HWNTnLGoE4
DtMEoEYx0y5RbqSsTf+UxEGbsSWRQu1dUmrh/ONovk+rGJdau57GiHPZd1GHaie9IT4BTWyAOD4C
tOZiWYKKp1BNp5n8QVR8GxL38vOgTWBOaKhBERmjYOUkXbS9Nh6iJ1hjmJxYmjjNWgYa98U6rQvh
pJh3RdYsrczZlbXNst3IlEJPwaXgWlTn8KEPi9iVdCCWkW2zWvhneYMQYKrp3RhBzR/1ZpYeNPQS
KOJblmipXOcx75GGzW+1QrHhMbQA/1vryu3MWDy7Hd13AGcwIVaC2S6zkhFbmls3G8Ceu9pShIU4
b9JM0S6qnvpwj2P3f4zUjHSdi2FUo6EIZ7VGWPHvDNWn3y5tq1iu43Ts8WaoGyJGnYCVqq/EPHvJ
f78YQvGCOmFmsivhPYlVUpwfz+eH177K/sfIhne1WCsYuqqOOWEFp/mnhrsL08sviBxFyCJetElu
NVxqBySi6Yg7rCYz3geSHWTXA66DugHHNfNEk3SVOp2ldomRvHFf2V/LF/sFOoPHdvMEIMpiN7zM
4HYxahE3nrjeY47zZm4BBwyPUhUL/KKsbwSNfSJM0XtDBkOdwxMKlGuTrGDMB3LI6njQIaXD49ns
dEYNsXYl/3M4kE5Dhr9N+cj61GpnTFzMWRohvEuHVu0p3QhSNVvRvjZEX88yTqlt/kmm/+9OYh3s
CaSoeYKYVj09YsK071oWF2FNG7TH7kkggXKqoLcMqky16ReDaNviCZmi9EsSAnImqXmWHow81q29
9Ow9akYb95JCu/iHzYdNm/JtqndTGJG0NXpJ3dOax2VFQVPgHBp8cmw6di2TelaPKc+em8oFOnQn
d3wRDWlMiaoYblsoyYp2dKkI87DxW/DvUa7arQE0/yV14iwssGOfpo/khw+k909QFXx9d0hrsVQz
01oHrOu7i7A1AMf3Gx/WzD+8Vxkdq7a+SaAht9zdc8IvAS5kudrSHDHqcWNA/gAcON0F3ogQZ3w8
sKEDBs0zY1hH333zYsqf0uZKrDLZyTrG6bCkjmr9zU1rxOJY2jyDCJXWyxaHeLcA5LENSpGWxj16
sRyyPRzsI5pc9qxfiX8Fw3RCjq2MOllpakaiGPDObTcqBeyasCj02aiffirq99C+4t9yCdZcBpEk
oAFPb1za19DUHk9h1xZ0DgvLQHQz/qsrup+WEYs/mnTdvvDRrdFBNTduZCyVHd/WLULVDObHnVOA
Tahfb/J0ezPA/1wMth1v+25tIMgoOpG70j9UP8vom9Xd1LTamT7R6jDwrvGodNwEyD+Gh8LrBuXh
I8igQrOQ0eo+MyKkt9R9fq0Rwm5fL+kdg/KLRVKCZTbso7vgl42RazEtvYRJNSysr+U3IovKvSxl
MqQGU3K+ATtWwtgQu/NS8n7npHed6Daj3zeRoXHmB2tomg6cX+PNldlxuRp99NIIS0sNUcj8+m0Y
MZBZgRZBpC4cY5nLlZL1mXLhH9/djfJciKOowM9B0HRLUcDm4XXVsYKepsw7YhW7WJCMoQN2ykMh
1hXfM7mX+fUJo1foBe4Z1BMB2lrFZ68PiK4Z2f8eCuVcfumMIghqZG5JD0QzD5YXwwM0A9NivYEm
4675oiLAFNL5sCQ0V1XDnS9CC2uIPXXH2U4mU0sLf6HA0miZq+9v4OzpC7SiEWzpx27y4QBiVURm
Tpc6ctB17XnJop/AwpHKIujRZcl+XrkKJgN1YjIa+hWZRX3xL2hrQZrBWKk3QV75g6DpFgVihi6A
bPFb7HUefMqMX299i9gTl8UFi7PAh0om/juz7z/vVXOF5E7Ge6W8/VwUp6aaRj0xqJ1bsfrDqEa9
XIxDwOXFdvYuWeayOdFTsdbFltLEJDKXT5Yw5BOS0ZL0HeEr9h7FCiJDzKyyMfKWqyO/2nrrhIum
FXdC0ntNH+L0se0KfzbCyOIXtPOV6DvJn4NioC4FewKoYehKOUW/48jM9RpPqS599rhP5M8Eymq0
ceKqKQrmL4XBOi9fk6jNZ3XTQIMEjkJsRt1f3TNIWzcIyK8n3x3BQKRutIy4IJLRcMriHNETFhVO
jfFyIJsq1/APP2PEwx+YPgB7D9im98ewyDxNxDlCPCaIHFR6CWlyZJ/QYJZkuewgmYnSvL64hg96
QEiEJKnvQXBnnvKUJLk39w+Vj17pItq5Neo/nLG8pGw4EBdDVKueHr7n4LI96GmbYa9GZiROWHrA
oNJDpa6EBjfWOMkHpWD1DNF5+9FBCcuEYpBXIb6vkJ4keZtRcroe+9iKLqrPRMhk2J7fEjxZykRL
JcU0nU8CJodgf9Hcy77y0KEQLimChBIF44faJMubAL9ZbvMci1BuX8fUFCxnb2lX9og73/oDN/aq
OC9vSrAMN4Zzbz8xJS0e9LvRx/88WSVvC9rnA3u3JZalCXSwR9zO+RdRtNUtC0F/1P7Tux65hLHq
1oobSxhkruQ1EQZz3k3FWfwpcAmlPBTb5jNgfdQ9T3uuAvfpuxY8xsBU9GyAEAMrlMbmAAAiuuTq
i91rkYIQstsdUOA2PbTP5svjzA+yVjVQITgvVyzqG2BkDohT3n7i+1jSH3d6OAkarwbupZrusmUm
uUjXxo1fs/v6D0ZywLUpuBn1UyagDTGCmtj7V0rDJjHPK7qoAiMl8Sm+F8aYYy+6ugYnIan1X5lw
FZVEtQFuO8QB8YCLD4o73VIJ8WCDxnhpTpzDQduXfHJx/Jot7XeHWt8YgHuL/lU15jAhQP8YRvEO
mwLAC9CsksvV0tmwF8ktX+mtIz8zXwphug5/OIsFjN8jl+arFcyKM/gzlOj3gI8f4B/YE9HGYF/e
cqPM4TKne4ugXpbQa9n36XF4UZfxJ/+W+NPl0TFtsIyhaBltP8qyJQRr4le/6J6HTKrVD9l2yiow
zu7AkefEbv93KI9yHaALSuzjPVf9hD4aJKXC/1fUpl/jnl4kJUqtqYnzM6N4ReNkOCgCBXgHjXZN
h7BZGf0RqJUmpQcJbji2KNvQAG5oC0JXxedQyZfLA7nr40JP/secWovs8m72gF1ko8CFy8kxQ0k5
kQjjvfzsASoPgb/BTZgyYt2HbCxFQB6bT0QaoMDuUC5LXy0SbTqWkt3xLV1ebdIwEzsdH+pQK46G
yFnalMnqMVjHUPcY7ZowMXMRG16CoNnGl3pLz+XNET5rWFVzwSkY+NNPS8NRX0ze3vtQR8I2nnJ3
WXqUlDsEjDyOtTckBuSSHxsbT6AqLNs+grZp6uJoYCIY/9MxrewEUxA+/sT37sulo1Tc80+DDsrD
YrYYqrP4MkgaJbyxPMml00KO6uXPkUfvTcuk4BQaL/f0ugdnikz/f599BI8CFeBdI555iHNFaetj
eAIQkgzb4qAAPyHl/f9F6XU8oMRvQEsrWmLnZ0wPrkIf1C4C50488Ee0tCPN+Zr44PxEX58x6yBB
F1vACNq754QM+hRyY4xT3+DqR3dE/rJHIgWpjlKkiAjXJNgbTO/bWqReXvZopyrVHUTKtfsgRynE
vZaI6t0vPRjlnV54oVaYbkzNmsFCitk5V7diVCSCi6F7qR+JSNjT/geyxndqzPRQqtCZcuJlLf9b
3P/+Ce1l+SG7zvaErg/ZACAIjnGaRqY4Ncl8hNOwm6bTNzz70uRgeUlA8xEdpCdIpfYOPF4lL33i
zyEYSamkp197X+d64XUNidh1YRJBm5ihr7uNne6n4GmZUwchVIjO87MxhdRQKQ/8+2NDotb+uba1
jusz/RYsG8PYZA3avKrEYY/HoCb0BUGPmGrPgveWaagk5ip78mzMUbZzLhZugJpiMjWEQ1c9wJ0W
hcMLuIkNpZl5KMer9OalIMZ5pyICwnfDynhxLm3NOaUJztEYImvPzGNZ2BgKRGAyT5+vWcrrwHzU
hC0yKZtOQnCGFRDb1rbZpaxhR+3kD1hu9cYtjYxSjwArU69eR4J6GQwFmXRpHDph8Mt1joDHihnC
/GjrV4ANtbrIgMQsB0k3/1sYDBo8GaDhm9xFZc+OOa65fBqq2kRX66CAKihRKnJ2ix4oOrdQ75u7
briqOie2xsfPTDfbmGbl3dPt+Vfffd2sS1Zl86BTvEuLeOiSshu0r4Vp8x3uC9MXc3v48MXiJsG4
d+WcEXCk4E1ukV7wjr3EdMXyONHbtXSUbZ5vcGaBkLBg/itN+2fmIjyRmqbpI4+bihcW0jrWDiWC
6lpDedJHE7ZakMnAjEDWCrdxwiYVcNoS8sJyC6NSNvOFTbk6T6zwsS+91hUwBlb4BNbHla2jQPnM
VmDJmEYOIwe04cLUG2/I0XmKpyr4PenUeDJJ9EReENbDGz/1pMvkQJJk5K4lbwYCTIe52KM1Uhza
dLAEeAelwy8CArlQ+cb4oaoJ0UcvgEaf0cRlXGH0fLHF04laf2muqMXwNaTJweHyWpepxUwR5nBX
E2qNHf9OTTdYzu8tPErPGEceoDlWqPOeuTLH6Pd0ac6qZn0IoHYVT0Yn4uRk8LC3j81I576NdpYN
2z8PdqfUF/CHyYRJu0A9Qi4PGguqMpvtTJL3A5yJ9zabbrBBUpbBimQALgyHqdyntgAWdvZHGX1K
5NB9QyuIz8RtwtLcQOAt/23zaiRaN5C/0DYg7+lRl+Zkf4y/OcVW7LZHH3Ab0H/Ok3sNIY6o82+b
OouzKyTeohvKW3YAdTBtbzW63yswG2Vnm5XwKZCxnZ7qBQdtP1CmVhZfSuTZPZnGDFBUo1p3SnFp
UtOp7UZlzcd9FOr/UIT97B1Tq67pyDOFfGQzv3XAn/bVtVNr2he7MkNxxhGp/IjRYhRu7nNCHq5G
sTWOmIq466wxr9C+Go+ohxlmNrKowc8y3gOZtJATUUx5veKsqcJZx4eb7uG/xyKOsd2+hJZ8pf5H
8DdTU7S61UzYMXrcJyojZDcARVgrNbbI0p0ncqCScZK48nhhigHRK3t9i/E/Tq4oFWT4oI6r9Yh0
78jA3veXtJtj580YVpT32bVVitNOxlBfmTVccY6irWzOsmTlgbpUErVarwVmu5uHmnJVOKEBLL0j
Padzfxg2FUaZtAPIj4z4bH7iP3CwoBxbe+V0JNUJA4LSUrpQM/G8pbjpOPph2PhB9zpYow8XswlF
75XZC1tqsWjkUipSwHxTndQXf+9vR3w9SXqBoVulOB7JXhjDZyZSRGVOq1Wg6tXiXRFaqXaB3muT
GKsrRWD5RETBQsGD/rHFN3rxrZravXNhGc/jlxQyG+/GrqYAr133hKClZBAPXSg6Atzb2P2GkVht
X0mMIVotsJV0nQhpJyxdGgVurIqHRE0kjbZPcKMDMay4RsMR6PFo+onz4NJui9LQAwN0n6wBj3pD
o+E0HziVge/Phjxs69JG/IrOGRlYs7aaaeiFcep0lfzlbRfkAcpXqC5rstlS5ZV/tIlrcVjlrssD
NULr/tNZO4wEJNvGJDdctGWbY2SGA7+GnS8/V1lo4OcNY7eUEQtMYi1XPxNkPe80z9i0hEcV4Wpf
NeqThw7KIGySNTj/SA4cMYzwHPPsfSEH27iIjq6aNePg/q8CQT1LaATN+93WzDWsoc5ElX/YaRQd
ZEqmEFGz6rBq7712d1UP5qlh6BQVVlqRSiRaxcX4LbLe9AquiloV8fqA2PadMJ1xl79Sp4ITCpM7
Oxiy1y4DjqYQwInlYZk96Y39juU5k6mbevQcRgEAq7cS57MxX1f7sVuo6LrXtnkdfD/NGlDyOWLz
5v43DkXUnYdLEAtwpBEm2ATTQkaMyhcWWQibB5D3GaDe0Eig3k4eOtvfbMODZm91nG/qCFa/Ma4g
fI4G1R9/H+bc97SXfibRXOivmQUf6dUP/CbzT3RVOYvv4NRf9DrGhw8YvZPqX18EqZKH79dBDPGs
tNCnLDuHb7zEkOaYjqfrgjnCPMOhy13MnRcA8dx9Tpb1GsjERn8Dr20+uufqBNi+yqJ9+1HUnZ2s
WB0rQS/ExWNInO4sstf/EI5p+hDtVMqU7yWCsSIzuR1vcAbIv711bZf60jK+ZajC4snvQ8ONCW0Z
G0cGIGRZbi6T3R6neQnPOo21Y7iRSW+rklrYyak3NAkXZ/C8CHL2/pZkRdHUX5xJyfS4wFMtl//k
cNw37cw2nd5JLAW7nyc67RelC/GENbfVIqK9JwcfMXa+0DNGZ2hylzXOGp4ns9t+MgMzn7r7EV5o
JPLRXPch773+V7bEqiS+AOUE3+WJUUltsLm1pIpINy+fev5Lf/O6yfnz8zWyultioKLxCVrD18Fl
2m2b235COIbrL22FubtmVV65WUDpC3ttGBFTK6jsgfnNSl5WR1lm/t37Nq7fu0HVuaRgB6PKtSaG
Ko4aUj9K8J4e2bQCgsEL26faaaYaVE06qckUZeDoGL1BL8GrBWBlGII1aYI9e4BSxZbi7BgyetJh
5xDodbC6PQ2nYybingJTUHFnaCuDpOeAw+mxni8y3LUKTP70KRCdSrvvLzjsgyieIs3E/zRIXbF5
OlYRiLnBkHSTbIiae01BQOobcXc1SddFGpkUm0u1rskcbECoZ8phtGfORxDSfGVb5vCS0drt5CBy
n1n+rHkAtQndczHMa1ypSKnq8/qXcNFWu9iTHEhBsz34+38Ob/+9DpWytV9zUwl1XgGiAJgemWST
kUlJ8JFW5t4SKvjSZGQuqPyCwes4dmuEEupkdOH9+9PxFVqYleKJGuoAaUOTeX9UkZsz9rTzWHTg
WwHeF6LvisIkzesC8qZp60tIH02nZy6Nsry+a47qLg+Meis+vIWoRglQXCv9vSJ+be7nCwnxcmsX
h4LA/PlJ+uAwq8J6gwsnkdDCut5Ok2KaN08QGJ2P6i9eQIK38HuxpNUmH1DiKHHSgWC5ZuIcXv/S
kApdjZqugzasrd0bIE1geul8UMozFuJK0553jWrrnWnzT5t5BS3+jdHSH8GMr1rXgPTtx9wxAgDz
Q6BBHJhbk0o+y5vhMUFjj531qIHQtCb29Au6XOaZ8FHnVmlTGiRogFNLJX60YmDEzNmECJi8M3Ik
7wpA/QFIW72SgQo4J7TL5Cwi/6dkTd8aGE+gOc7E15a1lHmc7hkvXF2NhsTff17XKhgVt58/oWcD
DeWCGB/B8iae2zbHUzVlVYLNPHAxz2jiIdvo0CX3nVUSkSIHtBY7d6jjdBJC7AEk31S9qIMX7Bm4
EyQAKuM8FNagkTE0TuAF8H1n1xtvdw5kutsncBfQ4QcyJbVF1pPLT1NbspUjQ0ARoiR3P9i5nXry
5InF2rt7iuW7wWNAjfDfzIo8U9hXlesETAD8EG4vYuMPAgSqXiIehmA9Vqhx/qpZeJl+h502ARGG
3TT3PA6MqLPBRBq7W9vRh2t0MEJLu5+u8tK2TQnYTKSXH42i7cmXzIleQVqs/q9SqH8XteS/dtd+
5qLqObzIdWSBPYw2sEmdjgItQpi3RjhASmwTpjurCbuMQh7edTj+2utqd9LZFdSOBT6pRq01XmqY
pK1jQ1gMqrNE4K2Z38hzRwqLgze62tg/DI/j8xVkE0ZHebgbOm76jvpWy8+Icoh+TW4dgWwKiJhh
Nm0p1EENqHHS7uuNTjWHmcQGg6b+6rhOgJNLgBTID/qH2emnSPWRLs/sOT+/EkEOw+Z/6xZMv8EK
lOyQKRTy9j+GSJFFaysQgLomOvyaS1sqvdXwRSlKyXOmBZFQZIzg7rPvLepLjWx1J0jLraec4Yro
q0xPW+QYTDTzCfk0Ak5qwEwylKYuiOMj0lM/rxBaYhpH0/5eI36QJxuo8b49IMMuxchEhsyuMJkg
i0K2cnIvT8i24aidHOfXemWmp5iqO7fkf7tAMdm1uOrt535Hb/y7jMA0pYt1ND/jYWzPuaPRkNEA
yCof37ICnri7VZcl2UepRXyylS8Dd9qcXYlvV6HDobBHAi//rFO4VxBwNpPlw19dvhw1EKheHWrT
/yBInh25VrTHK872KHSK5tBvgWCsZHp+3TaWQ//AEW0ky2HegxDsabMKU+no/UMWR0BjHMiYG0R+
R5vPqmSth2QAXJqOe3x+0rZRe5Ofr1qqguIfgbj0bGy3JiQeDGgWKwUXQWUlebkveC2edUGDaWql
ol2UAiNDnKQnIBKPAHj0Zd6TuVOEXsk3UQBPCtBW78JyOTOL88mWv4++tzN/R2cfuatLw+c6IwEm
B6YmGT1xjIu/BBG3ATloEWFhzJDCypqddlykHAaEARyg7KurjNyHSGaZ4dpW1HUc12gtbTgBo6ZR
F7dltz5NOr/AXt55IaUFmpdwNDltTekUbQuvt430OeiDPXjzKiGEFefJesdJYabiZ11HHRGJxyo1
pliG0HQ62pDY8eAKtg0tOMBnj0bfDAfKaLlnXfndLGKWSrQbndXagZL1wZn06n4RF9XLip30gLnO
/klotFQsV7dgAbuVUd5EZ/+2n9uKs3s3rjcrdcdK61REHxEDLQC+N5UJlw/anzzWovmAF0iRZGSD
OKIprxHC/tfYoy523UAWMZBPIwnkPEd8UYuQvZ3tv+dt1Jiui0FvAuw3fdl/+OhdW5FqOE7w9zrO
Pluw1KAkMqoID9B9jI8PNIgdlc7PbuugNsoy1K9t8nFIqg/HVlN5EmZ4T5KCZAgDfFpN6UbAh6y0
EH2jGu7dTMKNhhKIWxRBglktxO1ONq/Bi7K0NExa+pYhqW/U8UaR+CNOWL4fyw6IEvnlAOZkg4n4
R3YPHir2dsTQQjv5qMUEH46U6XhRcw+Mh3f2wsPAE0cLslbVS0+MY2gm2jwwh++xlXQVJGKEiROH
vkxkEWxCKzfhitYv3gyj+JYRdx4/vohVvwj+nJfgfhTwrryB6ZH6PviqFDTrbZKlwDGUgZqsiWCz
i6G8L2HjiRhHXRD4rgD+O0sjVtX1RjNCV6g+0sv0AnIEmtAN4J6FcbUp1jrHdh5i48ewibsHC8TR
qq6DpLyXPNsUxgtKPA2wlz1RPa9ENUvRPVoddIU4OTA4ZOnZQk0LZl72XFgCRTRhtfStGTzwUhYx
4BOJarwyNZaa85l5sdxfRdSLYh1VJtpokoQ5WgO2QGB7D4y8jli5kDvbMkz6n4Bs1ehGokGwnonV
cpWyx+4MoesB6/zuupfi+m/cl10ZH9YpaCYul6YXAvw9A04N22lAC79zJR9hYrnS6y6nWgztJ4Z8
PdKx3J/RYP/jMvYW3ugJH6antmLwlzVPgz7ov5hjvk1aftWxVhRHb8WADSy8XHfjLFt0LaJi5YA/
OxyoyXeqclXJmzEPlL5Z6ElQvBlB15ulW6vUcBYodNo8AgjMSTUrYcc0hyaOLObQXnhmuTulXdTX
mAvhBuQQUGqlFu8cEUHzJb4zSKoX/RTTI5PaQ6xRLu3I/H2g6XVo+erMM7i5v1EFIE+MYcTLCgTS
kqRtj5R4LZZdE3SgNgYwcs0cazxdbOx+K0VOfj6ShSf9z+yAFO+u7ISJHTjd4Ci8fJK+7fW5c8IA
9slOuJeqvy8O8XVJ/3E6vrpifmL7+SuH/NLVy+cKAZwTcHRCu+n8VHW3PJcCt0KHETsDGEUsmpMl
ZrOVgmw6Kjd4knrYW73l+NYsJhoPCeyrxXTLXrUSdGrpnvZlGwSM40a8ssnqxoWKAz7L+zPT+kHQ
p1tz/7qw5184K3yaGDx++tAbI+UiNWea6XGJ82asZ71X/9y6aIAGLNx9+Zsg20l6aCX/vdACzTIM
Tz8rcgvb7GQp/d1Sv48CLPwNmYE0pz4QwlqvNeGo0kZ+HPeOSZ8kNGU2SjA0GSBcwzqMFx3LS1FA
zzqSsSUKYlTu0/Q116RP8XjotLOr/cJqGl4nhB6IbwZGYvS+IbvKWMUP1spHX1psf4MYPEyGpIDO
euYfoEA9OHUOHdGujrBmwsr3ybI/rxy2CiwvWG9RWXw4X/FvQglBFY6ybm5SampKXthuz0KMwsxe
geBQAGepBskfscfpdfomRJzcnIx0SUaHkBgI8UBgo7mueoLb0DjAQdesppE+sq3WvByn8qIa8tYH
lSryh1N48jsejle4PT0pSQxZN+O3t3lkgfXwhMc2jpm1siU1xTryKEAcctior75YcojUcOKT7Vxx
hQGTsnfyP5rJEqCELoTuwSyYrgdx7nXLDOOup1HBV2rM9IL8V7EZR1pqfc5oybsskaFYL8D3dHPd
z6ImEcreregs8f7vDnurElPphxV/DrYf9Omhpf4rTbDnOd+S1fRxJFDbjDV3Lw7UmH9ZkW/VLQga
CnZa76qVfTCjz4Eykr4f8l+MMASjfoXqgBNSraWo8PcultrNFe2xrRNmwGxfiwTtFGY6iH5Xo2kB
7pVQJdFpL4nv4s/PCokc6PU3l25bN73d3XGdZqMQUUkhv6/8v2n3vH0hj+y8997EPTZ1yAXqroow
Tk/flsM6nzla63BmfAlOU93Q9yb7mMTu58XIBHspmqJuoT+UHBqK8Odq6ZbJ8/qqrh073cfKyfDN
wEHjxIOuuc8BjGf0MbgqNpPaPzyG8/ZMUo6u2IYIW1wpuMmiDO9MXP3ybh7plQkl2dBA1Wtf7oiB
0qa6rnU6M6B/VlQUoe3aw1N0Vk6KuKqOd+HTaOwjZAPcLhrQPwmcfNzOs1WNGZvUZw79pFO3P0vo
q5zUDwQXmdpSJ4UNGH7n5Ptsp7d6e7cKzeY1ONRwXr90ZW4Yx1mp3q3gT/ALO3c0CP5sEF9hNHGM
jdEWFlRJhblqiZoqO69swdX4u+Tw+A9V5pxOnFLCkhrkRhnuhLZ6O1AZGsi0zoJoOv1Lq5TWlJdb
Xcco8o0R6QPTqu9aLZTrRl8CnDp4+IR83qH3RG+FKUERAP/uLldaVQQoaASWqmY1vKQw7bKQMkVn
B0R/u38+DQ83FLueQR2ew63RRyxEgwD7EdmIcP0wmD5y85e9qSddhOzqw+i+U5eLv6XQR07z36QL
YUt2+XduSetRIvrevPfHFJDLDWrz6q+42pXSj3m24r/pNhI1ASMhq+szN0iwVSxA6dzuo8saCEw9
hE2ahU3eN0MRY/YUD7k/U+STo4O77kiILaDkpIAFJgPUuL/fbZEF8DJo5zIzODIZW7yXtx/7Zjgk
OZFo0R7uhQjoFPM1a/vP7+AbamexdaWc7R+Q8Ak5Nea0p7xfx07VsgJRl3Ijrd2OnhtlSA8yU/t0
2QnXA+sv0GrAxykcmJRpPtMaho+thH5HVb0Pg3bTF56BQFQ+Di2iXogkZvZDxLCx0rTvmTqfyDOQ
G3GwIATHotGrePL6ui/5ZndrMaSQcOKru5RXmxxYTKHDD9ZbhaDrRTMhxOEqftVxZTNk8HGzVN5G
P+R7Wy+ejbVR51Q6/IU5g1/vUbhoyAKo124e4GlR3dCV885kdBvj/apt9KdHzaILJSx5SnsjyeUk
qtOTViLuJT50OYH+IywPWMZQxkER30MaLNj6skznMHVK/oJQ9zY6jkdseSmxwDRYbSghVI9/5C3T
t6oYveuXMcnkkG2a4S/ndf9xAQ8xSAu8+EhwdCx235+B+2HemWDgeTUIeXqBaL/RYARv+mV8INQF
sHwVrPemfaeG6dvqIcWkgguH1Lg6P8V2XVkyuFO/ZjHb5emCV9Oy/MZVBwq5aeaypJtel/gJelfQ
3Ws0Zw0I4gjJKSemlWu/rrVTrjjWLV+wOYYrwp/PERHot43UZVvv2riuMObptDLsot1DtgolIngi
kIIjETJGJC6Ag7ge8WNKvyVMp7OgYtkZoZqftcCQ5K/RAhld5akJfUU2z0RvyKq369sCaRrGw9Hm
JfBWNt1keqPW3mIrcKCwU+kQeixySQZSSYajDk1X9Lc5kseB0N0ack4mo+8onE94bsbfdPsrSRJ/
n2oUl5LXnN9PbjJpAsB0PyVO47T9oMD67HFb/tFoIfVM/DXJ1d58XOnVCp2K0TK1u7D/sbMc1n00
WSfth7LBhQt7gLp78CJn5fZkSy9iqK/Wkv5bFrmg/NMPgOpEwSIfMRHVRG1dHc7GpgEaWmGFxE3Z
fMjExFrWX9ESxzWmvTdYbtlkPAoWFQ57yx2D3t82BVTGrhaBBGXByiqjXpP/+dvtgWeGlWnmLXX/
eOySxw8AJBkXJKHtl7hClT7KnehBKk/hUsUVJqezv9tZWhkYm1EcTLiwn8Tw75VzLcXgC+6I1mRF
FKSNf97h+mHZ+QukCtUsXpb8Raidt/vcElY0YP4ZuQamMV7l2oOOUYbmHRXLURA2rMI0b3vYC3PS
Iccji9gd60gvAxkZ89jUD9rlXosLwOif7qTe5Gq9tAMklFQuOXIVlrx1WkA4CgSmd9FFB6vmP61e
5NFvRlF0R6fbzz2bNMhmMybcfNs0NijQSMUo+FaB8WQrbpa68L4FrwrlTqMIMa4QkhWi+SQzGdBB
N6IxWbYZT9OiPWAHeuZ6DMIrue0s4+NGNgr65z8SluzKIaQNagwbcBpUbZFmVwL61UWmndPmB+m/
Tr4inmvotiYMtAl/29Pr4JHcbIHpUfLCkUIYjA1nduLsO7OfzAPzGPM8GhygWXxlwrBdTH5CajBz
iWwbSxgq91qUvgcZFl+6/KZ5QQ8LP4Hya2OyRIC4B+nBlvWm2u10ReMRSH08yIF/Htf0YMJgct2u
Xx8raTg/sdHU7e03M2Bcv/d8IWRGs0P31PRS5DsNAbSIROwlnbnayF8NCcr/6sgd60YEPK5iSIUC
pyRo2pcEqsXxopz6bLjgx4UUGW3fYgnpFrCiqajh5VZUP3pU573rKyl6wj46YVgLZ2AOfG+3oeiT
mWPNaRGW1A7HFJLeiQZsrVSKqszrUkpAvG19B7e6fgx19P5CoXVEb2EpYZXn3aTWA74gvfgLkVcs
BpkZJdO4WqZQHxfJVvIOOftRjZwHz8/V8SGDBIwgGnuvftZERS+3Pn0zeoKOwIbAr6n/qI2064BB
anAdVBJ3KIGh5n3ABn8TplTsDuxTxURL8blPIz8uHe/k7SaKgSbf/+87HkR8y988mP3ooM2RjcE2
H/9Es2NMqU4NEF9RT2eQnPav1/Zw1iG75kOTEGPCEn5+VtXSHlYofXaJJaxvhvWFXvDypX0KOucM
Jb9wB7lGK5cajLVBxy+IJlRed1gxRpCiMC/SUYgnBuE/Jk4wY9YsEUN/OlPris5nxhIOsrcUs7zF
lTxkzPi9wSZB3E0V53WKv9AOiQMOf/nbwgGnb5ugf2mn365lT2s89P3rLXzpOQYxWZ8nLAJvILKh
lX+IiAk2KhVoroErMfwrkEcH246mkP/mciN+UtFX5rWd8VX6s2SWKFxlRPpctjYBQceuTL44yEO5
jKcyV5WNX+Y4LI4wqHrItZRBNurY3XmXG6gmoaDWl1+FFMflUChU8VsqFXkmMdokFQTTd/r8bTlZ
Yg7MuaiDaVRnnRXVoj5XL0ow3OUS+QzWV9xLqt/Z7CwuJRDVkDeoZZnt3TgX7UgODkfmKTvzBZH1
kR9mk7An4d+3ORoo4VyUr6RFmEBA6V1zNhVmnSp1f5EQQr8SjgRHs8+QLJFAdBrl0K7MfvyVgqcd
plPjo71VEzwE/W3pfgO8dm8LiulYzcJ2f6nfhQTeZBnMCiKA0vwArMT+RstTBsklXWUEJhYDEXLT
esFvfg82Xy1uFMo6kZ/At3fwwAaqVlZwNkwDA5nR7cN/FK07VB2ZHA1ruvVVcuxhWJ9tM7lkDIb3
citzeoILn/+sUf6zsu5FP9vC4KKsgjJ99DfoSUxpM5g2xyqjw50B9ZwtZTPmQ6XZo4W3nqwIWFhf
S3cPP64sQNTJqhIeRIWvn4xleBQ04dxTd/SDu4t/WaWRBAP9FdU04Oxr/58k2zsh56R5FVsycQ97
vikAsYMH5tCxf+3fIXJENklOmR1Y9r2pPdJYj+HLnM9VqmCMjRfNtxO03VAUYWtoWvHkqMohMjBV
BUFM6xY5OyemSEhiII9gt/1ntGb2qUU8QuNxe/33P7TmrsfT6tGolhJ8aNa903BrOATAQenehUjv
ySJjkxpZFiuXPbT6DIAE8u800btoLFIML9TaXKiyHH2ahsNwRdwAbQvl6WiQ6QmBYV9Ha9YPrzZH
8h6qakPQaeZOSHN26RhGabLl4wCTuraNS5TH1D/+RdXTXwOINuktu6uLhQpJQoMFF1ATXXesSxF1
y29HZ2agYTyO0QIzg66e9+eG4d2LFbn1m9wk4du1zjvk+TfgGDnSY79bzyhoCui7RzwIuJRgrlu9
c0l5rQXdV03cX+QtAysegV4LUt9eHNQ5gQv7QEIe9EB97BsAGmfNbaWqLu1uTaxN86PyubnvB3tj
dbWVuzkwa8VFDhjUhDF0Hm1AK3TXpnWWg6ube1X7JmhIRS+zCWuTIcWlSX5lQtEjswFC31GjZuJp
IRAOjT/5Y0YDCrmCv8ITC8jCRqgBOVN71PGCxJKv43/7Wc8fgSNEjhwX9aMXT3DTG7bD8JewUrrF
VFlybtMoZjM77DtRHJYNWn2NikfVFJ2SOINNr32kuEwjaOYRl8NJdD5KJG9M+wTm2Tuy88oMp4PD
lbjF3bcCpLivmbpUnAZ/dzTwQhejQUixUjX2d1g/fKsCOuA6ehyqDPwRxEyhkwDeQVbEKFct/jdA
QzDrW1i5V0+cBlKlI2/YJ1WfuLOq9wYEWArFACyhpXO2Cl2kpLcWyrgXsXczJTvn46MK4umwAV33
HoM6jrdVTVTEGH2z+FA02tjFEEk+aZ4qXpeE0vAm9+q4I3KPtjdjlm8vOGY7E+N0ydD4juZfkGOk
mG9bhJ5i7kOr4yWyeSv6wvD8Kf8v/uRASd0JcH49IbFecyvZonGQQbU0sqFS4akNTJBzw6e4iH0M
gbLCZrMsN0otJeZQtInGQYFhE5raPMWTOghQwjgEpVhuIS+QyNjP7A5IHs1faTIfUPh/Y9ZGNdtC
6FRL6JKPoo46UYQU7ij73eKnu0fjrJsb4H6Tq6O/W3B3SBhuxb4ToE70qd00oR52/9d9gz9qL62W
nOHrFJIvSNox2mFGha6WIzYm7yewlkHxKfyxKwTXHquSzUIlFT8MZHQM7eAzZJEBH1YQOM1kXhtW
y0blrMtcaG9daztq7Z58Jjt/QReTl2qj9HupxczbtZuhy2e/2wmsYYJIc9KAYTlkVBX+H85AtkQE
gWAGJ8Chy1DLivFjYtlo1/dR2FdI0ujzkGFNQBHzv5sc7qutABWNFTLtBX2E3gDf/Jdi+s9B2gu9
7RzyfBIG+H82/TphLtfD6YToRRpfSQFiDIbGbQlENl048B9vmcxL7G3bzvWv0GBLmQ4Jom4LjLDA
ddMux9JB/BthXRb0e51t6c9iOZOFG+MQKyWktFZXiXnySMVqJOROPVrhwnZQg+AtTJaAXRajcdGg
hP1da25J/SNq1DQh99iyxAQB05fD8dOCM05qpCUtz84L+AroyGvkztP06I18B1cjxnJq954YOowv
97/r81Z0wLqTnusGrYi+Qs5WR9NOg65I2ag3G5hTAoUiFN0itSSSxO0XllgCmQx41uDe0vfA9sYz
8KN4NlkAj7V2cwgtmY1B33K7Dc9+bzyM/Lz0ASsR7fM4A9nipHoz0BFciBLeuUoaA5+uiLUAihO3
hzZkvZfSEmbmNXb7wOvIC6iEIQGLVzJivwCLfSodWksPTvGBEL8wwjPGrqJMSpDRiZufTnGJ4VaG
Ndjzkt5bbqhVU/E+GtdEXZ+eHWSHEI0cIFsszeQE82jPguVu4OdDj4Prmx8aU3Eg45niDRuw28t9
MNDjLKXvK/3wqgMBub+W1k5eHVy/TSGT+SWVmWE6R+CS2hmzKtK76pv801n+sW2DXiCBO9Y9ddMc
I1Y5zqgz7+lmstz+binA0bWY/WGkChs76qq4RrfGpD2szhwkEr9Mb1QYYi3CxccCC/mvTbIBBCXQ
vDBiGi+d+JJ1BPWkVl8INXuBk9eknldShc12nOTJXVWd2POnsC/AQR/4tHcWYfYg7VFHxfW6kGLD
f/UUP5qFvOgGLQXK9qTP7CAOu3XdcxsttG3yYKU7fSBmI/obQwkzyhgWOSzG8ZqVODptbZE0cfVd
UOzqX4+jRT+nTKyzL3af99wdllbHrdM4q3FRuazhGj+0ORg7PPaKeAlZcQVlBtVkchuHTS5Yg49S
ykFGBsNUOnz0YttnPtSbgtC+VEfOjg72+Zr3Wv6j6L65ilUhbodyqflYbZ9/9h8YL1jE7nWiguke
qIs2EMn4X32u4kAkslqRWSnzJLpi57aBVTwkKbAhmPYJEvshQzjOX7pwv5Bnujv1oxaO7pa4I7X+
Wo1bREK8kfrsH6vaU8bXLIJcid7VB7Cxj7kg3pCocdzT4TLPNzR5RNGVLTgqwP2khiqJWPxA4JzR
h2qGW0JDctI6i33JyqvXosjbTifV4XpC3LALk6RgTN15T2b/b7ah0mjm03MiW1aZm7l9ugoUjvBv
MPHM7e30anFtruFIH+e1Orb91NIaWPfvUZcS9LfYqFQDAMGztS14bof12rbKhc57hlKgV2sdEbQA
TnCVpJqASReNX5uFwHjPWicWjjwpOyYSxYRuK9IssRJjJyjvap1y+6cZy3VT5A9vDaWxkMv6rZHV
CorPSDwJF/IvOWipgR93SROEejKUxVWRUOHOAea2lhT+1Cicv8KXNyICUBNg978aqrktuA58cvhy
14GNRhoMEk0aXD3zd4Rb8/ljNlbOC5KchmmzveppYD2S4czshZ2pQestmlbk6bSfBbYUsYhQAVob
BSNGvxNk8PWT+a01IPNtvwjnpnIzj7dzUt6eCZ/QhJrWhlwRDS9tZuuIPHMU9mxyCQ3H8xdEgyMt
TvBzdOhYlRArC8tdG9vdv7F6FH6SUTNxWEWCXQhHGQdLiQGiOl/i5l2w4R6ixXvYSdiHovXsDG9i
n4nqZa6apujkqpO86i8aGEF/pUM+Jk3UBOA6YxMTAsZR00rVMSBlRooN026J2qL+cQ+kX1Uvys2I
pbGg5Ng48tCGZqC/242CVHMWIU+wuCZCgFx8ZmCd5rL3PG8nO5/rSqnTGwHixjtm68g8tP41kG3t
F0b0Cs+5crn3jRrSeV2iq1qShnplIHvr0YBfzUbfRK5GCRJ5g1Gv6RIH/E4n4VcP3VzukZMfPBI/
Ab3G/uONTi91Vl4Y6lqNMuycsNoKj0rxbUtMPYdQKh0TiM93TVXBF4+afeu+WSqpySqRU+vP0a6v
IFAg4wxQdLp8kkOe+uJ4uAava8c7BfWVybZLmFtjqlpeFDAvHA0NYUuX1CplxJfJtFf87SNsFDn9
ihOA4L+oSxFHAORzqUBAa8vQj42vEqKo/yn1aUEvj2ySk/HzIRQ3ueqDxwbaY7lVSsmoOkAIOkf7
a/yy+lzInXc5h0jZBDUa3bcVjS4d2AoLtayDvNEmiTpTW8aTsA+TaA3IoXbzz5n2cIUE1JlPRpu4
ecyRFU9CNpZjOXphmx1vSavCy7L10ZFu1/SJ9PR7nMXx+dABTF5Xjm2Jt3sAWBb7yfGeAM7muFym
3FC1wybi+ZXp2qKP4R2hondNDXWJbFVFnX+RjgMwk4FyKUBWdKfzXnRUSFywbz7LRJHydIwGQqE6
jkW5T4vWXhkpcd6GWWbbANrAQscNAGYJlNJrLu9Rr4w4kq9dW7/2Vd58toa0UXltz123O7FdQKqo
MfHgHVGY332Fvf5IdrYCIuq/Rj9ti8y+x1junNVQSWVBjeOYcmYu7LuuIHr9QjYbsm/f9n9NcLo2
8wRSfw+BVNl7K7Qau0QnbI8LQtHZ6gYyc6HZhyItVFHIKREbzxXflvz4zkU3TrJY1eDm2501w+Rw
4MGo9lwe1c7X73y+G6jWmzAQd99erm+yRMZxXiWF0bNRQTqptYywf/UIe4yofll40j3tG5iKuUGI
mazbVYtstZls1vBE8gZlJFlIv7ebtosD79VyNvlK70UltgESAoEse0P735HrD1d/l3vxMvYu0e+q
2WhH6wTHj/3JPHuBpOtty60jmOMW/HeEuVyMnT8gz+WW0v8PxPiU+nMg5aTjhgCPSSZWPDwkfu5P
0hMR67VqQ7qfhOJntOOZjaV5hiUcfyvcqN2/6bc1MudRJOEnlTdv3Hdz/YBmJvm7RdDAkTnf63Nu
hhprUqQPA9nHzNlAqD5Zu1dSOFL69G5yi1KFJcX96fG6lmD7v0D5KqsxupBGHEDKupZ7wHdGP5xB
73l0Hfwv2pHOPular2fCLGLRM1omIgxIJFSDcaEdBEad5urscQDt0tCjs8F2So5JTswLk0TsKcd7
xdKzdFUf/lsOemsWjtibf0SAvhLwCh17oAYfpIOUbZ8ieJWgQrentxwdEW09spWzFNuNFcqjlD3a
6IgzXuGbCQWMKQ1YoF5f7+yGSaL5RI1ejnpd3Shi5u6hOGQcnnA4ARRhJuZTeuXb672Do9pmPJtj
bY47lOVHca8ufd/9wOWq7I1qnbC9NSLBcwP2OswebkmaY6CZgvbg91MBOhBRhCH1gkx9h82uDqIN
HEuwArkMgaahrRFVOBJ7Ekbkbkg/tCclIUYXDnMbPXEB5LzGe9AMrg/5gSWc6bUZZogx1/Kc83tH
lS5dD9GFM58hBDCfZzRNDTy83iaHXZ5JdoRh/BRJ7c7aNs1qVQQtzGaqcSwWnAGv8UNE2LJM2Z/+
jZ0kmv3wE/+6j4QBQZTkhsRN9sVvOFohBrPPwFCy3gVFQ1qLVw3g4CNmbRmBwJYw+Ky9sensAxrP
/DF1q5x+Iu3xXBVrKLIKZrJBdVUjg7tyBiXUrahfv1akERpkFfpPQt6Tz0hKdk545wuJ8vbz1bsn
lPCcCzBgbxPEfpngdeziNvneU/++Kj0yevaIc4jvU2xzqiTAohgqC0YC2gTvmP81Ybm6FncIvjG8
VoIlI2x26o+K3b9cJZ06prtC4dXvu64ST1pVCvzCSSVI3wK5ZfOeApibvj2Y2cBlUKJaij4WeV2o
aaAiy0cQGOvysrUUDlky3uYu4LOjyabpUfmYl4tQNOj73UIr/oLapS6t1zLz9zCWtToUEpL1YZuv
4dPJ/qgS+2EWmi4s6eMSzuxi32StLdP0OVfc+cQ5tr/JW1cmpN1LgqkB6xTcF3/qUfvORIlzPZjO
LIEKzZDPTMEPPLA/FEoGxGWsVwnj1CJ4mhioBPBYCpfzxNjUAUzx+cb946YGLVN58+bRTWXGr4hY
k4oIb7oF7/KQi807vmgXmzKzydcR7PiKMZiCXQHpau5YBvNa+4UaaDy6vtAcipB3dmyB+Scp/rv5
61WdYEavrQ7zr5W2Id+llFC3Hu3BZsRRT9IKSCUt+TVzF4K+A79p5W/knS7XNwc8mYjpy7VxULVc
2NB6tDvqmFK0rwNtMLtRwZNvJH7R51MC5DRx33FI8fcfRAWwcbZHYwUrt14OzbygDajE5b9m1mAT
rQfzVgcfZ1WwurC9Zdk1PciUq4OG+bpCYUjz68B6R6qdx5ifWOvIMbs2G7YF6DFUDOZlqWQ8cddq
nXgfIBZaoaZE3m3OdpF0KtinIStl6VEjgcQ2URYEvgCng8ZhJ03KpflNP8Uj+kH6QRnftIouNISX
bCa8MhAazthU9/rmV6WPGrQkrRm4X/cOigst5ejM/HwDeijoauJZ3S+TF6jka8J/XdefdOHkDyZe
4/a1Dz3pgHfzcJRakWKtCyP/60frCdMVlDXHmFwiviYcXhk0xrezj4aUxHBQ8xQ9RA4jN2UCRdpW
LZQ//Bua43n8f1Cz3nTJupqKNbdSn3tY0eAGCW0uTUR29+vhfpWcuke3geboaE45j/SV341U5XK3
qd/JMqhiIoCqYFgr4iOrd7VHdwEVxdxw4/BV3xLX0Vzg3hLqtfMJ0w1ORQFeE2IcpX+M/GaU4Bv3
IIhI4aHhS1coJxIXKc9j1w0xiLEazbNzqvZwW2P0t1g6pXfsy4ZaOJTNWC3ttnHDPrtTTf2+yIxH
j/mxTP0yR5OnSYLd+U6zqkjJoahRYcfOyrKHM0qFEZhnpF6ZM3nZRdpsql/IqU6fx1a2EId39Y+j
SrKi6TxjtpJ+b313afe5Su5mytrsZY6PofthsOFqro5S+Pzt2owTeAnJNlTmVa9OCSGmwryoYWs1
ImqPICCUbDM3vQ47dfWOz0cx3hcv9QckuaNTQ/oO/lJPim2v0Y9fMGHscYVCkwHPBD97QzMc8pkO
3A0NBunUj5w/7PtJ6XT3TZezlB8lejFh9LxTrGdjToV57Q+1tnSXsb3piwvt7Ola0V8GjxEPBDGD
CQ71+3bNe8FjulDsX5RyRZm+mAcpUFs1qdDOSob//0H3ZvYu1WzSTcU9ps8vg5l68VZjohqAPiis
zS8mKJDA5bm6T/hqj/YTK3t1GIVbkfHjHE63G9AgErI67/BDG/ooBwgdV0dT4WL4IA/HBUIEYtQ5
j0tCLPPXpEnORznmLVSbeEEiMkOqXMK7S5wFNKAv9ksun0wmYfGlmge8av68SP4otNyZvFU+qoGX
B1mPiD6yhKzMNbockPDub//tP67VzJn/2KYqXerlZWwYS2U6EmH+39l7URIB6/Bx8a/hK/PeEvpu
F5FIJmFwap7qAPo7epQjxPAPOpIH9sI5ylV6AHvS3sHGBO6bYcwecoLTTILfk8+zyHt9iRyFxVtM
i+ksnZ48l0GNWn2APdYplXJRAZ8DZ9BqptIbSIEMOveroui+de8urhctr7K0xvRn3nLPVWP3ZAgq
da3079NFxF+cZ6yRvuTlH7EpIRNa9YceHoFf/Nd6E4cugiGkM+rMo97ayBsgDIQkiGwflb8cTqHx
z5T0LLMFsFX4bunhwYDHtqG7J5x+O1hpRDFYMYkckwOL30LWNRQNzog+4qRLsVzRCtqBDGA9RURd
Zhc0Dtu42JQPcJR1CZFaXHYV1LL5pCmb63UZseFnQUAdHCioLdFkU3zqm9kq8dVldJExtq+NFDBE
Xx+iFTy7FaFXhwL2L0hN98f46eooe9JRNAm+w+HgZgsXdfHEWPu/ctfHbQvOU4UuL0i3ZxXWtu2M
54HmLSSbH5Qqz55NRCz/T+ji5Y2DMDDvROCIS3Sumpr92DsfFkUhOks7SzD1Z3KaRts7bVvBGBzd
uSzZB/+B4of08+tZev/908W91QUlkr3GNwbQaFzCB1BzJ7q4YJGEzdhRERQ7anlG64Lq/gwf71SB
ETkkiArNucFkYooBtcD67zDb5DRIoeEZyfgZdhp1bx4fiCqWDe32Ju2/nzVpL7wykDrqgtPOtEHc
sMWwQg1M2+ktjImdL8OEL+UUVOCp+su0L1UQcQ9Y059NyUHKkKx1eHFMxZEETPHyRARnpahFcGGF
0x2Ky/4Jj1w73EV9NP9IDFzpsXwobCMDUdMR/VyA/Bn3WiQWUZ/RU+iKET7dbTF/zRcbVoyK+80I
PdSt4Gyvk/eiXahsD4XkXS0/KBYjgMegUXv7VHBGLanJuNmmKzUjUww56z5QCX6HqFrFjOLX/esA
/OoTXKzWPpmkYkA2+20seLeigipnjGHRsj6Y7NyPomyN6FTLPrdoK1m9lhRFknWGu7aJX23J/lpu
wtaSCOLyrD+92udVvD4X9f1xb3Dp9lScmAtVDfJ/zqZLSS24tGeADXFv+RFTvjUNxWUWj4cXVxMg
jJqeQ02nftxeVxr0I0Zr67rWwNKz9U7L7x4KxRa0QialaWgf3GrFZHqBTz2fc7zbCgW6XzqxRxZw
pPm0skcXh2E8q5ux3JGUgmf0eH6XsAgp0OZQW+h8mW5S4k6894lvYM/9K9dX4M/w1eerq808ZBXi
Fx+8K0d/JA8LOPGyQNrzO2xe9Slzint4XDFgTKA7zKoWodIU8cPJq7OEHK8pHsxcF/r9dmyWjz5e
KSc+TSwYH8D89+NRIYWo/nBn0yHclVgxV3IVXGkSemiAwPoUs0lGH62O6IxBuEVgpF0QaQU3VBoB
NPg5Mewnd0LEiOZ2rtELlj8HkWfNWrg4svC3kb47nHbqkbmn+FTKg3eJ+PCR3drFghgfjumhijEd
2eO6AmfuTVYASfQrNbTaPGCfLCCPlb058hYh7zNumwzXFboJqcwnzRiuJE4LSkbKQQBJNaUZXOfh
z9FY8zer8ep0Fpn8GL7pV+hyIbb+l3QyLJRGam0HEREAWiAd97RmSBIait9YRWzyfBFuln+Fb+vD
3Mbz4RqmSGA6/JzlQ5VEeUy7obYVW/cAjlrsXsMq7GCfGEUpzga65Y2qAKUxWKWJtWh2Sdk4ghho
pzx5p7XqlENSvtQ0iILSqLa8b5EjDZ2P+kPuxU1wbAfJm1p93Pl9/zSKgZW/NfQAlk5GTFkgE+gQ
lAS1tGn7NTDUfrktHs88HZOEnk1Ei+Pa74t7OSLNtWGdiArblYzrDIwxE66ZTFQwjOUBYQ6wF1VY
rLgnroWIley/7634KWvE335ZA4x9AsHH9st2btEWbMxQ7+mtEnlkizUiImqAdDGBz97VU0yBsxYc
D9GIRM32tieXnrHxTMA/14FPgiCF5nr3rXoGFVNf9NLILbPt/pXmpcbTHnlKVTkT5wpxN7rT/jeO
0fCy+4EuXoW3MPeiWrkJonhERM/cryk5PQZnKwt1RAiI32ujn42MmypBbrPQiNKlp9wW+v+2iN39
U3k+UrJLDlDDpQTFa9LFKn1IudlrzuzpYqCyuy9pkQD5hVKtxShwuzAd0a7bdIhGl8x++FdjQbbx
X6Y1nOHhpsQfmfgCyQ0V1uWVxOojFFr6EHYQsGJ5c1nwIOuRjf3/EfSBKAlxRWvBBsnPo8n3aUjz
R7T45RjwzOS0/CQrSOmQe5W6WhIE3AUIIEEWdMz9S3RErWcywZPJK2IzFeSKTo90qXX5VYAcWZzs
X+lJb5VyblzckMtSZ1g1AxJCE6u3K0wfffQT9zGBz/EQ+Tip+m6hWdVWGFiUDujA5AJvzOc/XAzh
hRt1MnSghZwmM+YFnvjEndFOQ6xzvS2GHnouKv7Xxx07UWwuOZmSNXgUIA4Ff7JkqomKqXIUSpT8
DiE5epxc2y4/PPWkxMbKvHRY966QMc7mPw7SLoUKKJsBLeIa6VP93DgIz54OmwZUOA0D/udePtxZ
CgUFP403xR7hGsDSLpDVX31jpmBCd0PIue7jrJ7nw0JA2yfSmGCuTZdsExV9SD6+uYh1ZG3l5RZl
Q/Og5vRajr3VL6YRo76NCgaQtU8unF5VxV5JSZsQB8YpE/RDGU6MmXsf9DCSyX3M0DkUfv9SIgwT
AaPykkPzLaXRXa/cyUtqbdPz31TFPmnsUKxI2LsEU0/1SuBKh7rVM38OQBjACogvJRfW81Cmfo5G
7snMKa6Zr1P6LyIQCU6jKyWxpNtmvQeJn/0F504+eNhp7SH/RbiEEkY+FX3Fs31LN2lNmfmfvx1U
imRDmERiIensFEv7SiFe4G6oyhJSFa5WLAXHM5mA93iXEcgU6rJq/oT6Z28ce+XS4bIvwpvYLhvY
xkvoi+00OBNWdbTOVyXjOOm4JCq1NE6EAXenk+lT+GoSRRhqKykhLzpsG70nvHUPWUacM6pkMaUT
KBNla2Tz+EWJpIxgciFI6L3+dX70tAVOVtcbsHsx7D4EqkrGIhqEsVeZdup4BYdHCghn52GcLimj
Z9/5gQCTIKjwWrfcde+r2YvflJmfK/srdjK41sqTglX+r3FzeTAbuURDPnlZ3lriY7yB8jR9gEuK
lInhMb7f0zi9K3XbfKBdtqRhDDhKwYGJGi5exMGkWyRCzd3uJxBTa1uEd9YvG15n65VoxSAUNk5O
Ql3KRlVeSWGWMs6M99g6Hp6PM5h3GLXo7NS+U2YmAcILyLeRlMyN7wegvvVIUbHhbaxvlGrXA9NI
Z1dLQTyp/GeH66c18Qr1j0uhl3Q8Ubw2AnQCrjNuNF4CKuBnR/t3PfSaeexiLeQpqEHxq5PB2Uv0
gfK6p7fHwzZhrcYoAY5ev+Wm6DtrlbQFeuIV+PofsAcC6HO+QZTUHKBwAmxbRwN8O5sbPrAcbNoK
wKkIOV4ElUlOyWq+KD+uMnLWn7ozemjCtz1nQTJnJK4FOcoB7KceMjXjeBDGaDrhAQVZvu033ut8
KOPyVtCfNy83btwYwR8oAX7xiBqX1e+WoA0eoZM93xMiEJBx+YYBMEpuK6IvWQ5W1SFZWEZr9Qh+
0/+fee8D2VMt7jVVSiY/R8F22mxkDtlqy2LMhrLGR3VnSAwwijJFc8fEj8xW81XOJajb14HKBg5X
NRqj3CYtgwerEItG1nTKtPGHtXEgb6j5f9SHxUgx1q8XzDzVw3jGOpyRrg9Xgcglsm4RFGRiJme8
Y6b5OH/IAQXKdMjzPFylHLSmVZgfho3BK98MtgBThMnQTlFJ5Oj7yW1MupPT73rryjmX9dvUqpTv
pvsrhghIg1i0gwmjcuH0eaq4TARQOer0v3PpDhxZbW9en70xDz+TJf8bHr5V41hdkxOwovYChMqg
NN4PAV0R3wzGUKORyYGMK80c3H5A4hm4PyoBoO2dWzcQsAgqX0BeIw2r+ECqUE5SiCourOAT0Fhv
+TW9mrxveum6pynn3GICEM/w3dVU3G7ZC60JgVf0Nrv4Pxb1eA68nmKuNMFwOrIUksxOwB7TGHRh
APmsVFjt6cjtzC2JVpEUil5o0RGLIifyWSGWa5ALnkx3rMgSForoW8w2oMzKnjKq0BEKWo2LO2+P
fQ8gP6ocEvAmfblo5dcNbQyhz8KIDhHMBfV0BFcgUJfqgP6Nca/+bDNycO5xpBsPQDOkliZfuSnp
DSVHBuPrLlpdMIJJR0XEUjwWZ4E7jGlU2mpWvgFKaTxzUqv44lQuo2uC9DLq/KEv9N24Q7Xn04ZW
wVE9ksR0UtHNEYfQg6hHN6+ghYzEgm6UQ4Pg1J4YmGjSNy4f5cTGgYv5K5xUNZAFzzW2/0R6j9zJ
6pMjl3zdaAiexTyd3J5hpuBRzM0Y/fvl1sgjG7j5qCjOVTl+94hB/hHht4HLCPJCXQ0RH88MHQJh
vidS3zt3fDsEyXFBVWSO9dj/2aF7riMBv29Kf2mqBMoBq1BHgWZ3lhGKulax4cQT5lEgQ8UDuxsm
5d11FqpFffNZh9ddxSqicdcSAdluzMjNfjuqTAYK8Eu6I99Ds0jijBg/Bnc31XOgVc2lVl4ym2GW
qRy4EOwZEjInrpRzyzi5vHFz6biu5F48DNY5xqo612mqOiKFVNi8nP0UpIAy0zkyPb6zqCAFf2Xn
XqJENJ+yAVUdZ98X72FOhVCC1jX37PXKrSlJPeL8yiYiZVf5+AmQG4zcYodMF+0vrDn9xyVEf/96
bzDTOvPv6bLlE3gf+TT1hO2hPZJnhW1Gb87JmZCtIYeskGfBPKNzkis7VoFbIebWsQSYtpUvSSiK
RFeBep7cXadNgt/HNm1o60VK48acSVldrVsuu5/eabYZWWccO60Dv9U2aq54P83TVZqyaaFOifbA
xAXy/kVMR3F//SeLe7sv6zv4IGkR7CQ3LmFetJuo3GXU73B3q+6klxXbEmDYGXdimSMEP4nEZ+Vk
zdEhM1I7fmNdcr2i+uf2bRvZsunbUx9PVbe2ALxowWIV3xgBAqRdRZwsjNGsSQcxXiZ0M/vxpK8u
rq1h3LfX/ntqfZG6SPfOQBVKAvPJ1lJ3H6W518XitPZQMdko07E0m+j/wAppOPi+J/kBUfnEQMb6
F2DunMbGM6HrHm4SUhgfRZIDmHp9+DXFg5InY+fLTPgP/mFu2tkDxfdijSukXrn5yK7YzRObyzdt
9dum2yMTKsTuwKXsP4aCcOvyA/IdS16MIKTFWskztyt+u2G3rfsLoiH+Lo+eNPuBxvm2pc2xlE9p
UbET8Q13pE9Zbxmt6pPF8+jGeqsuLmgSO5x5Ln3hlbyT7giFV5DmCrySZAhf7QBpJwpjZjaouNfu
OaGqkn8OCa1ygG+fesWs5vUcV6oYEjk/BpXrwZ1Gu2D3aMmWo/0fJ9VLVKy+19uOMB+6YDzj9Vwj
uDGMhdkzjJfg430Dx4BgSRCWScv5gOMiXuR3CG6fWcbRzo9l9MD5ROfyMN1zH81ycjEDQHGI7sOv
A1k89xRendO7KCXRLEuWqgu5Z5gPOBJF3JnyaMyrXiFrrWuiTI/3CIas3zFhqNP4+ZzXiepUMaiS
L40VPNUUM4FlWT1+TP13IXtyhKI5j/85Qzw3OMbnQoIJni425Womdo4uKFIL+zyAjPCdgcNyhRzB
GlFuNo15KFXiLEfe5tfpbs/NQ2OeXaksRk31+RCHjjWPV0ARatqVTqA/MjO0Tx6G0wkVIMWBsfmx
KHIjoc7ol656Xh3SutttXDT6Q8ki8RGDoUbHsuHnJ5Ti7XzT94Axc3NAfcljU2r9wZGpsOQdEF9k
WLGqgEb6xFkONDWgZTFqeIqqMzNZHne1s0JMI5EEYE4RDYZTWtn/YjxoIr7qf/qAhw+xxDWvP5nn
UbyXaPEyj+Y2D5IebH9nXbDwdcZOm3AssWDRDBNT1V5cBPe3WnetbKD6ClIi4611YhcJU+qyZmT3
qtERDvXtHyxghsoljWaPK0GiqhzrjrWDbFQ38OyUdFdLvfA5w1GHSC7z1+FAYX1F+BnqX825c1zC
85Dtc/xr+0OrRn6NIeP3+pKkBvP8tVq3jKumfaQIGFa73xv03Om8CDCqmTvCIKpyXOIxaiCYeu7n
6dwxqoYafYE41vRWiFJx80BjijbrAb26ZErXO3JYiqamObvjq82Ie5pXzJ5/J8mmnW9wJQWLBL40
IlSERQh+GZGA5Fg4AAQBOvAaCjYKGW99RZItiapUGBjcLU6DrnbvzLGRdQs6aJwO66ic6IntISrW
NKqPIPOteciou6Asib4Rb1ULaOhdZaS7UP29uc1txgudPHkwAfkAen/5+0vWj8O+zt0pY+TKbGsr
sHpuc7n8acSFjsP27dw76lHa2xMWWbbDSLqx3I9t9l/ziIE+CXjCr0zS3oOC5lqzaHhbrmEbswg0
f5vO+mmMFY+Ny+Lv91yEDyAta1JQL2PfK3rk0kAPzqU1anMUBXpmZpBKRalCRH158/vuPh3z1If/
8t0y0zSY6etfiUsRQmEdF27ZYZkM7a8dmS3nfgAHt0BzDCe6JNM2htThdiCnEr/pX+NSOKDjAVLh
gSohfAy58HDlido3kdj5SqX5MlDBvpJn2snyterIrVOEvQertUinzKbzL8GgY6OB1H80CWZBIRJG
gnMsu9EHFkruG7dIUrTEJIxi8hQbybF4eqAz8zeCQNUwfhRd0R+z46CagKuij1iLt3+Zj0OL4ijA
D2lUGNt7scLvXoG8b7A/uNekMKCrx8a9brrYhAEgGyX6A6RVdaRj0mepMpxeBJVByv/iVzVbQ2VR
+j5T7WEXxqYHQJ7Zx8JyayA48cGrxm91YbVKcCy+px1r+uEADwxfctvz1RaLM+q5k30NZRPnvev5
1P+EkZyVZ6N+exWuQtui5RaMT4J1EM84b9Nv5rPwmDF69aH2h2CjjZlZ9JcN6RlXZVNxy8LHFpW1
FnKHzMNT0IiIYCCQnVgdOmAWscqGW3XWycYQov48383mUyzS5hlIWHjo2DF9KS7gqr5UxMaLygln
iG25vx9zhxS/3Vbq4dbJhhEIXI9qsIL4hg6qvKW3wWkJQeUOt+GGH0azVUq3481yVR0V+wD+C1bV
cjTxbGHYCbMMcgAtCJ5DvZQGEDJehAes2V7TjFxlpofe58nDBjKDIhOru/xc3cNs/Eurr77nlY+K
OtDQ0XUb3LiLoX9AkGhSwdsuP4TjYt5JMnBlGHNybs9/rCOb5WWHVPnUDFTw+2hujvi7S6PG8b0A
yYVzisUJr3OWjvrwuyZ4E7TpHlKBtvfRKoJG9UMEfGa9ERnfkFwpBslT2YRrBMplkvrpX6tnXuDa
L0GjKLGEnRISes47jh1387iidHX/PAHc+1LQAE2lnAaCc/Xz2Jfc3JPUqxlfjE5gLUOzN/ETxLmi
z+0UJDomcfYKAR09skX3Lc/+4hAPaSzYJjZT+m652tX10p6gH6S3ic/SeGsKfchqAr7Hy97NxibY
siT3Sw73fBUgGKhpRdhmGrG/l0UIZoEa4LdNF1FmmafXsevLy7VAY9UpILfzqlTRKKKHqQursgxQ
/C17lQbeQErgZrflddtZTw9W5X4Vvj57oRDLXgsU34Bct7DtAFduJBWq1x1Wv5eoOOCapr2lk857
lSKI8q85SHvWRKRxBF8XGqnkovlVf4xmpFe2XrSdJw6YAdOBar7R6nXecOuSLGfp0uZ6WF7Q5xsR
K7q4OL2AZ74MyBVaij/i00XDGQfqMuk18B1w7ym5GJZ0PmTiYRfvzAYigC4sXgYPzcgL/p2/QAzM
Cbd9dMuABG9ncc4HbuMuh8Q0/VhkRipQL1mYhOoqVU69eR/as1qVf2rZaiyvtqHlkOOsh1Sef9I5
898kMgqJ4RXLGoKyIYzE1C/zAi2XgojKCCHVK7XAyZHGebPGEAZgOZJ1FRdUzuQ18535tNzVLM8g
dZS2J3yZdfiyB7aG/e7Xj90HMycJwCJbz1naDKh+OJdyRKtY6RY2vY3TTaK3DfdbVV33b0pjXP6m
v+dW70qIap1U6MebHc/keGnO7RYdxOemvPYKE8cF4pyfAUj6UdGeCOzDeWZ5nz2V0lGQ5FacfN7e
/AK44xsXFXfA0QjPgynBYkmL/p7DaWd1kef5wawsMpCIFb9i3QE/iOIu4y0wecGkFGQLilQtkeV0
3moJ8CnRj2nD2TRWgz90Xu5BiprrOFBSARlwNrBzMZRnxzu4GHHPsWhgT67esJjbDWEULEPZ2EUe
T0+FfD4oMVytp52VYv2JEXdqlGv7eZ+U6s36r1ZA3VVIH2Xw8ZiRQuz7WXUchBJLHLd6VMcJrNeo
v6SSVyXrxow9A3cevpXHb5MGImx6aMwjkRnRVimzW45WV4/bMYwshc1OWeL111sIyXg06uYFRCHU
8c93nh5mlyesVstXoyDM+V6IBoES7EUR8Ly6Mi6RfOrYKPammdO3DGuXegXOcWYIiH5uKmeyO7S7
oHuZAc/f8QWLIjdPhfljagPTo9sXJ5r3w2CceBOb5nJ8JsiRYcpscqI8hAkGWKKFGUrY+zavndHJ
Xvl4GjImv4X9cBPtIwxYMV+k8VN88htApFe8cYGlJeoo/l8JhAd4QA49MtUBZspiNGYsGaW9CJQl
4mEL0I1wj1TwthM2Flvx7uKKZmxYlHj/O7K5nDVEOgeZWSuLOBCzbwp+MNZ8YudG+W+gMhsXRXZ5
kLmXZhiKXQliiocJc9Y9ecMTZxwwXGXzm5oilIr/oZZvyVgyeK+j7V9k9vQyP0UopNxs1pMmtGqJ
7ntwTPzwDVRAJ9+ago38yXthwaVinDtxYwItmGChS5auAgHW/kkvwbuoZFYy0L/Lqjdd40B9TvvB
Sr8cvFtFGGrs38K/bGmfg+94sFXcRI8ReJ+4I81tzmwap3XosBm+UPeLFM9Ksr4d3lovoNtEdPeb
QAcO8S3GnAJCVOGJ1gAopPf7YzWXjg+RjsxMvyPRzIpm2oNHnu7tr1o74Jz3SGoTlRlBxRPaf0nM
MnAsXl8Qi6jyCb//00a7hzsy2zshcj6yrUo0s3hQe4Q+6jWNhQgzKw51fzrP+63AWZBk/J6E4VPl
xlF0qACGt0koy4yjdpjL9+1ae5DpRUJu0c5hM7wudeAvsuPAG8n16yXD8YFmZGp+rN6aOf8pKtpM
QsuTvlG37UucySY0Wy+OYAXGjn1Jls15ZN29AKxHoBgX8DZpL23WMRka1eEIcLSgeOS0mtTDHPvK
BdMAllbqlSK5lrK0At62TnNxnLWZxbRty8faGun/E7cNlG521a1w91pfoOpidv7vVMcyW6ZJvaqt
eAIfU7vF7VUNip4G7QfqQqzJIBKnh+9/nAfrN4FNGOm0bLb5A1wJY74rkXbLxPdJseumLg+GW/D+
oglxfXGTgheJ2XUdP09GNOhO2N3RcnZE/U/L33dN7xMvyOqISQhnGOY7CBMlII6V2cPlfnEix+gE
aYxXyuDN+SKpCopzBTU9Obla6yEq0zyvQolCOycK/41diW6Bx91zrQjrBdAV4kXkQx3oVELC5sv8
J4jB5pznlQN4/3+oz+qvqDELP7sO6W7jXLFbOkt2PuhkXPzbbBvp6gnUrEdDA0QCQi11E4Nok2nK
LvrXuB42wkImNtKBsLpZ/D3qVl05qLdpE5UzItnsXjdaSV1a0Fz2A1BBv2H2uCga0iVABxzJwhi9
TBWi5x3cLKq832BQ8HZUDkxJ1pcK6lTtML4/6yf2gpLTa62t8r3ae0n1LI2agoG8UwJOfjJIYhWQ
gzAvdths31+UnnCN4GmnAX1vfGB5NxWEU3xsbm/neAGLhNNeeE1VlqVobKYy3bZUJ/im7V0VzqL6
1u0KNFSCwPFhZ9zb5GpN2+lOz33bBOn6CvaWpSCoRIA5+s5wIA/3K+iu9lJfTYXsIbkgv104u2sl
G9p80E/1NHCyfo9aAyx8vE4ZHJwFzQ76iGflg3/cwQ+7FA2AM8WD5Yf17Vo2ZtSGpkq+G2e84njv
YcKGIwYzxz9uuIIV0IB2Nm2lVS7kI5llKMARt9yy0J04i5df1H48WxdXMGavzIreq9L7ZRyyfwzc
9HC5fRFHGMy26pA4E5G/0zNjCweuFcKiP/k/jd7qmWoFPwDA/wb1pTDIRfQ0v17XmoZRtbdC17Fl
DtTNCrPIJxaOY8bEyN9N22lLI8nyS30pXUunc5vX2mhEIi3pbbl3MevTT8gfbfGWwFeGZ02GF8kF
mLQ8SmA/5LhQMuAKWv1zvM6ROfNxhZtiBc+b5pfub3bUMLkqu7DkRPu3AKj/F1ZtNDXynK7r6tiA
FlAOMleMqjsLB3kA5/bVc2uKfF9i0Mv7jjx2DstwB2IJppGAlMs/3sCrMlO9KrnHXlSGqfbfHPwv
XoceOvSHjg3nEAbRzmnzrAi/vCyhmQmF/IjwRn1uiqGtrM55JBP+yytkwIP0dHOgEKxb05zK7slk
9QSxlAQG8uaauNxfCol86es9A3YHccyMghe6DRVgOSj25jpQEE6TIAG8jm5EiJZj3yikVtZ2PGJO
ZCXdgy3D937zSO4Z/YEp9cK1ya5jgagBET+bvV95tgaPWIvcMR5WLjRBG/Dr4tlaWIBR5hMEXt4I
DoQWE5jpZzQyVm9IRUbYCMu/6yDPTeOsd6RtdovLXOAGz4AzB5vENm9XAVWpY49wPT25kgqIY+l1
fNCnwVD+zdB49ULcmkjvlktJyqDacAqj71lSr9w2ijZ1oeqt9NOHAU0VTcnJ2PLSnBbGrTlvsdKR
XZYobYxVQsEB4O4d6jLWcHmJqi7nZ/vHE6+wY5vMiuGRRxmwJSvldc1TMHuaR/U4a8bUo/DACZbx
Y0D0P2+FzwSiJa2lNLB9TiNvRoMntU1M4DmOaOcQF+qor5ZxrsL4s1Yo6yju8qajH6cfb8RCFO90
i+HzhZbKw+i9n8xPvyxxcwHg+BVOKVFK4klzWFcQoT7NhWKo5nLK/tZpfExg12UZxSC3Pw56OxpX
Wxa+bAbOpCX8gZWpRUf08r5Zv2j4Hcv3V3/dt0O8p+8Ik1EbczRMk9vtqCaKR6NLsOHMNhwgGVoj
LG4Er2pZMeZDln+pV6vhOtJf2OHHzqSbrSa6CB7aqkcOypTm0i9OmamumCSki9LhzP5Rp9Kcl/DQ
H/23FefR5D/OdgSGwd9VXyarX13f4VF65qyoTqnhPJfIYwbItp3pFsRX1aVi9Jil5grSyBrvokgi
ozUH4uVSq5JYf/mrTvE9Q7S+vZDeufRNbIwCGs4FMj37MAUe1+QU/o9/arQKNJYFXZNIf3JczRmG
xhzi7YJAmmIWafY/hAAhc8tzQ8G53k0QQlk6qjLdBSxkxz/hgEST1KtA9tEeWJ8e3cM5TDem5UVl
gnfk676vSoz9lX2vr3sL2i9nH9iTWib1zujqtN6lduN9YILmwI/Wc5/1QSCUh3oZ0jaduTPhzAdd
5ZXMr8qAIV2mi7BR5ZOB+zTQGpRoE7sOpEldS1muSaxDN7R85AqSzjBISkvUN0n87YPEEsdux1yV
xCgj/NOf5zLd7DYBU0O/Fok9zYRkGqmqtxuqah7J18RHMFToTC8/KMqzKc2hzj93GpuDx2FRc1mT
gQVw0VRNnuQgiwB8wJIApPgcRgiQhYl7qE6gq6bjtHFYsdFYDuDQ1v10dn7kkAgvGgo3L7T6LMwH
bGFpo+HH2mjCbTtx2/jVkcvFFUxExxSGyeAKmx6jkHQRtot6Lxk+UmiCXJNj/rAsVpIZDzFtuOUz
kQYBWBUkgM8Cv/HNIhNXz93BsmI041m+ZbJDXqTdsONQEDxkBVVCOVsdv1K2G2MGSG5mq23AO4PD
p5rO+cNH5UYItMQyybufLhxMj1BchpXZAPcQ5MPHXxgvXd+T6eOYSUVs2y8aafH03dwN3N08RKqQ
XG1Tmgr9LAXCaG105hfsTYnMEqGORpkA3cITWEVeOMNDHxKfM3m6IoDt3/cmAGmlvfxt+VCqEYKi
rwpyhXaegAZ6cbtEPKxZA1endQFPpETTUWIM3pZuR/sbnDeZ3BprN6WBF8HBgebwWA0I0WIWqDTk
s8GWoi0IoWJ/xstN+W8jndA3itn+okdhS3+b6bMFbkHQAg2NCFK11M9EbJUc0MFdoGIHYQwacKIz
2xbIOHGh1lREq7ldsKOB8L514lAj1O7Fr4q1p8MxB2V1yd9izS5Dzd5u4WO8MOUHvgJrBEp/oLGP
fmsFLH19p108985sefQyehS111xWqdmW6tmXprNs/WXZ/b0Ck8MlNIu1jDGYWIQqmT6sUIQiP5ng
TmkoPCUVhL6P0/gPt9GXRkL7MJUCJjpXkZO4Ufa0gjlV/bZHoISJIhLV94IlwGAuPGN+GhgDuqGJ
JqBLW3fV9/OQBHhefVxgLIU9s8tIYDuKlGWr8f8ZmAxjlK5aMf0Ox5dYQD5F+/SILXTz7VXf91Np
qMP571uchhAaHTt+kr3zezASLCafEG9Ind4anol28zgw2hUccDHYXYaNN4NPEBBVUVMTislibmvl
dslldyb/6IHPBS6aSa7SHZdc76f3i+uWlnVZ8S1F/oyfxypQkhYJ/SHMcXHhR0hhzYp9pwvBtMED
+S7Bv/GE3D/kkY7C2njDD7NuvOMRi5P1wMqHookUcmWeEQo8m3Us3g+BW6r7P9SIE1kJvlZcafyz
q1yQtHyeqARRA9rp8TZ2GyhHZmEGP2X77wRYVVhjtBikvFxV+v3T6NBCzdRXBSuBAfELGMmL0DJQ
Qmzcw9xn1uaSgF83SNAWB0Nl8g4nJ5x3e7smRmIF2bCDJ6s4Iji2SM0Uu61fcrZc3vuvTkAlO282
2ATehsZ1RcyK3AVMvhpcsV+7wZ1Lkz4+8BxRYV0i2uXBMIzIytGTZHJ16O3L00Xon/R6p6HNRkTe
jyY7f6qaR0jScK+mgC5HNHEum/emwGeD+wvQz96GGtbwgN7R9pE8GURYXvhGzehpp+E2swFSquKz
V/ubDzNH/4dXOCejw4P7TS6I+SDtUkKk9A2sixQ1U+MwMmWTNY8Wz0QoQ+bcd6JlFFGZa75CdLAr
vIfsCwWqx+KpvBESbW5BfkMj1cyz1EOeDdqAg78Noz972Tp2j9qMXFm9GaPUtjU1sMJBEXEHRS2o
b0swXgtoS+vy7Geeyn0IodgnAzDcNvBZm07sBdNVHlSpFJNgTDnBYrPjJ3F82ESW49ZUfFbEmnKf
7La1fiS2gggHq8HLddJ+lDjej+a/peRcu2LQJJ/Icnt34Mfph4zHKk3z7MqTcYgODj+e90wYWNcB
RrtUVsyXA4OYVqHcTtKsGAZkyY3TAqHXw4HPDPxKkZVKEiH6HhfTkMb1MT6QLD+6AnBvBlLtispU
+q9wfTYh+lHKu9yfe19+zM6UvddtuY6SPK8n2QFciB5L6Flrm/0A9wbN7C+ga7W7vV5My7/0sg4p
7FYiamIPRBJa3Tv47TbRfE+sN2sexTygTufsPk3mNuodgqIfebo+Qk+4Lk32WMMuSVLZQS+zgYX/
29mHUDEgDW3xhkBXu/+3Wfm8dLCctIDsHMxWy38yYCmJ0JzEjh7KQ8ON1rDa3UZBmdtmMOOEKCN2
/7dvpNAAR4Xh4Lcwr/JNIcklVpffsfGsGu0iY27nEzK1KGEdJwapFlNUfXaR+y+4OxG0zz0QLcmV
+KuO8Rt+iHGKVEWNK/77z8xm/YrpNUVHjcjLjiDzEzx94uiUtXCKW3IOECAUUMktb0kiHy6HT96H
2tRsiv116+VISjceIb2nqGJUVmDnc+ppS5C8oF9UdwzhmgUBuI0zZUx+q81xMSE2bV2vgmQNO8Jw
qOPNL2mOf/Ksg5b3L6pt6Wlk7kgMaJv1ADwfZETau6DiExo90k9N9gXpiYB3S2pfyHkC7VatFX/a
DtX5xg2zsAR8PvAOOdxfyZxZJ/7hpmwWhIVdlykliDZs8u0Jiy2ZZa5UDx5SplUmcUImws2KruPt
NqT3EndYfEHuGIm329c9quDLnUnpy6sP6J20hKu26Z0PMfvHqp/GxSkzd87zV2pY+AyLL9mAgBIi
PIQny7OkZq2k5BiPPclKVIXNCNdf55+jPfphXBes16ceZ8ctzV1GdVJSKrEgJ2gKu1GuLiiIvzYa
5MVmfFv6pAS91BQ1vl31822rGzKlGLINLAt1wbxCByG4JOXGB71M+msFw8SwIrRzV2eIM3aKauSB
8xPghYpw7QVJGjT+JpdRrYmPhGwkPTH2+X1rdcM5MPeVmyIujdhnni5EIc1ITKjBN26TAQXuw1Qn
UrL8Qmkp0TXejXWidoqz9/x8mX3zSQzH6pHpF/LOOJPONUCAHMAbsoZxixFaEX8WIxy3TLvmZJBl
E/LpIn8nuSByDf7ZE2BHrUBmJAUapPIv0ONKWvNLThTytcVcnCv3S6NeiiTM/JlcTEFNf8K7dJvR
wRYyJNAx/MhF6gbHxuz+AEarZjtpBAYy8vBqEofdyYc8b0SM4y1ima2nm8YtZJboLXE7bZvgFv6K
Phk3Opj4RmhrlG20Dhx2iSgFJzSvScnrnqmDHKB77EUE+l53/cA9eAoCAobN4YiM3mri1S6g6tyF
TDmFtpJX+UFTUdU1LeU9yVHorjF0ORDMK7nlshebs6EOkP/ym1fgfO+sg9FU3Evdw4bNdkkFISoC
UttZQmEsh3DEtyDDgy2zEWqfdxdpJWxMEHBlXaqKdM52CP9S0UJ0gbGroIGUWIEG7shNFjkshDMN
MACOyi3usF4hJkA020FwCKkkcRkcJ2YsNvmNWljGIq8dsnRdKSfN8dy6zjxbrvaNpIv/td0pzYWO
GZQzRDyUqI65lcL6vHFYMHTwd0iPOUIKbgrcSlvqR1yPVTS6c/Lt+yD9t1XYaFF6N/4XJ0raU35Z
unPTMkCgtb/33xouj/qn8/JpGhxL5M7a5O4updUFh9lXoTMr+1nsga13ApNj7pNciP0a3k08ccMQ
2GLqA/GUR7ydi3TrxrjTgv/LxL4CASXLKBm4CIlEjLBbmkZhEIHanYGELmCpYtTRt7RpgITdryK8
cgXJ6iOCuwGMuHtD7PAhkUUp99XjVrwZHdOzf3ldYcBaY+ZKbd22Z3B2aQClg2k8HyNt+uZMvkwC
GqdE/lMuQbqAruw+1YDydG2uT3w+2NIm7oMqqrXPZBA6I25UItQPH3BSjiB84NDc27Lk7s9aSZnB
sbdziSS4GVzBpF2HaYo8VMmBqsRIvZ9PykFXNgGgDuFriPPP87Xk398ZvWG4IMh8Of8URniJPCqz
tLkLDqoIdRO+N84iZJt0Ki8wG1RYBdUFk9qsGeRbuIkaa5h5obxSBrOD3ehfajyBKebX+XXIGPbO
7TjnCuIhG6E/kDsl8YO0+u5dws7ujruFxWqA2Ty3tmXTxdVy4e8/KDDxxLZ7XQQVjc+EkcbGqgw0
UmRPbEgtSFAaKLNx6ro0yCsb4pBgZvR96IsrLxxaMv10ESYJ2yuJM3HuZURA1Aj/5FIxQFxp11/A
H7JfrulpP77f9L5NpLWq8W0pu9A1qD0/m1yMCUm8fZBrOtFmqKTRI/fAcGuDqZpDWvrvObUQOvMN
apVyOtyg2cdVEkLArDyw3XSNuVjykDuQzX82pXsJ0khqHIRav7Z+zqXYvknZeejrkZx+gV1cQpwe
TwxLw/cYFHp/2fp18XOPZ5B+GnHbfxRA2WGyHqqcw2180Mt+KGYUVG9lu7Lw2rgzUz+/SA4++Lw9
LhY5VV3L4frE1BLTrF1U5h+ojHyMjfEo+awCPecHpCpGXGa+Y8jcLlWQvdNF4IdIzZyoFbuc8bq3
fyJ3J20zsiIM1MgYiUHBZQQuPAOrJqATaHlSVIOw2UVaSlCs2Ep5dbOJqIIxYvfT9m/lqWqFaJ6C
1csD02osN/CBA/yEAYZitWp0KerWwBgIeHsjoOYqzu19RMqgZKGHepeyBmK/PGDWIFiZ7eft0XIJ
mONEHX/xerEUiCiAEqic6dJHGl6Of+wK88ax/nKx0RsPt9mSeLN8KsPVUIreBE/IK2RlSwEXjzZF
FGj/7MJeLCXoqO2uJoK+NMcXEbwOQ948xplnjFpYbXZCTkI49RZyKCFKnstv5+pJM5/kTk9tX8id
3YE3xFJ4UZDy7NxHrYyqvf3bTDAyBjIZzxcAtRQDP2QBkiFQUSBjxoidyzTVDnXzXFWr4Ivw9R84
hUn/Nyx9ZHrhoQ2ZGUbCFeMHx2/4y9MaoR7RdCVvz037rfJcp3+CMT8xDz5EKfuakr8BUy8gV8+Y
5MmIiuoJz6pe18bGj05p0Ed0+blBQdYb/X+F+ODT9RbX68B7qy48sBP0mNud9fR0T2d8PKhvVthH
SRi7+AXmCwR5MjnxFLv1GPK8YklZYrUsoIwisox98FDR7cE1JN39tj3yXrWRaB0sVC9kY8FtapuJ
WIvnqNI/6TrtPmBt18M6zqslzrSfmKIi61RoyRqUsPGeYpAH7f62o3DQNbZrhAB/IBs9zXxta2Y4
hI5LShubpoP9VP9cRS8s2Wboh5Hi5GcfiCd0eNGsOJcH12p3TzO5v6LngyxR++tpGQL9UDRFFf1C
CzicTZ4Lbz5sLGhrIrl9jepSlJzVRVNAmXWamIYl3Yopi2AHebnX1IJpjI6pks2KzxxgFo/hU7q7
RewQYV6BspJskyewt+VvGblA0i3omZgwmgR1EnOVaU9knDfvxcQ3pjePIrxk3DNaTfC6lqT2uI4s
iDluYjjc7M6r3OyIq8p9HMvI6rkq1Yf2jjWUOpKro2W8vSRBw4iR6QhIRJlL1EsTO6bgEXBNjetE
zPvf4NKJnewhgEgsjPuaOYku0cHfevcbvC26rCJhukrVvGGXQOAKvCygVjGdVbgRe/Lsx0Q6sXqv
i6NT5B12FzlTrZKfOdV+ocjZiWwRqmVapBw+1JQ6JfW91/bHcqJP/pLkpFrgKFnh/Hxq6afFFL53
MsIjGRhwq8P88N0pt6BlAQqXqim0ssl9q81CVQ2XlZacZ3ymJmq7y3rUb47wxF+FWiy0RWIuYD76
ZDi9LyWIWzaZVBjHMTwppm1bjkAMCmmKHpu65t3s8xmkCDX61ZiV6yyV7OMVgKCRf459Zto93RUo
7cNknUtmBf3Zszj4cfv6wgh2WwE9uncqtp+GrTH70o1MaXsqSGqfunt8lVgJeosOe41LKKt1hLOF
ha0w5qNTXrLdvJbNn352tBvnlN6xeFjpZFOE08LxxYJ0ZP/fLmM9EWw98AVLNgUOVjAbd0HbbTe7
J5Z9hYHyLVJ09dU5uB1ODVatpS7fNjIcDri39Mztm/WMLGbw1XwR+HTIvSftbDY52v0YDn+XuvJk
Y40ANdMWww7vlYxz9QA2fKK+EhnFQGNjV61cEv1TG3dwWbIlyTO63fca2LXp8AOr4ByAuZIHR5n5
vMyraoQNnct1UwzoKIJHfJH2DFwMtjHUFzLqr8WSUqX7VPZRVjZrADfe/Q2Q1l/R3JOu2AVhWHmE
JbXkuqrd4lKnKp3DHoNbcSvPgq4FrR4kPr309OlzlUiOzO1QRuD0hy6amLHQjNwa/a6jBQMEFbws
l0JIAuwIzwKJkGPCDCXfHb3pY+ih6PFGIVbTvpKAEiCYfaimA/oWt70+pmhEI1guQFs7HYFgn+qj
wi3mQmJmMQhsU/p/Re4Gxd5Me6ZWt7kziAyxblvPxiFz7G+MKX7JDVqcR3MuWH1z34TgJSl6mwHW
pU8tPFdjnqeunXox1T8SezKLv4AEfAQxNIEfempOWRARnwVcZZsnUkQtScU/cy9g9st/hD3IkyPl
NgnjAgQSud4iOXYsBV67aQbbDG8lrajr2hYMREhYX6HJzcueOD4wNxPVu1Sa0nsnZMygJHitNF8l
uy+RrxXZRbOdO3Gfrt9yXb547Nbr00kVMTH/X3zo4zEHkb+etAAmU9DoBGOVOfr+3adEsTFICL6a
6FlNXs7qoEg0EsPd3gZkfjiLVBq8+6CrvD72/MMdrJZfm6YJzUHVX1AhLjMG5DRhPal9lSzYwejw
o1BgJ1NWwtRCCu19kaRJX83NNn1vAgOIXqf0Jnw4Gwsa0N3eFVj/FN7EtzHMK8RLh1pQ8aqwHDZT
eYwlQohpopIAw4egBl3ympj6KSS/oi6fNJtQ1HyJDBXtulqATd2QypgbUUplHG9YYUAYqfkpyror
PAYgZZ3Gg5BwriM7PmvSmwa3ovmvTGdHmtxTrwwVDGuAc4wyoibPcL5dP4Tei9XoFNjYjWFYWNT6
SRrNXYv1AB9NDDxE996aTAcX4lE23+/kb3UnAEnz/LLpvrwbLPkuJ7ZX7/QMv2gqiuTgJTLngwXU
RLZf/eiTI/sQl7YZgrbzZr4U4Q0vmvCVglkYdxUvVEl/Vbdraamxf+ywaRk4mxbEB1WXcuKsjYLo
AST6Lt5tSCsHpAXxxRb6AJMU60OyBNugDZIAcFgmIFpMKkuTg9GJa4IrGxn26rbsgd+k2kIBHNxy
wI/J3z0vx+whA/dU8AZVrJ3FKvX7UauXNriBTHcuTRqoK/oCHu1NamNUWArTGHJa5zT6+TVYJEH0
cWx/UzLPBuC1HoPr2+/zVy/u3GWVKPeHm436U6VzbXugS6HEz/ZphpSLj6LZHflOcw78q88cy9hM
9+mUqJqyaPRtYIpZ6CyblGjqistEma9LjXG2BzGKsa4RzK9jtAhcYSiPos/a3iw9qxDwnJMaUXae
m+X/OEIxNqORhP/nrmKNoPfDnnJe8enTLH9oyRRITdmBMT+76NuS9jMlVKG4IjdeGjkQBz98HErS
RN1+k4tIjE92CZb2NXsLaJ5LkTQzZ5IG9BpKNBHKPffzdLu2+rFTN44C+vym3d0yXVg7hbQlexoc
rG2btyAYFNt93nFgmKMmtmNag8f10Y0sQI45OuLv3gDf0lCITNF2mLzfpLDL57o4oIVOb78iOjSW
8TlRhAVYAYjXJr1h9wCfXxNKh/BU0vhtGDWA97WgP1hSXjMk4K4KVp/jjZpcaf6eCeY3M57ulSgj
djYlXwMCo1piJnImAB4feTfRM0qjVloxgXp3VsDXIzLneYb/u7/6IBL95TJPTVwZwOaTYuHq9pno
JjP40Ebz90BYu3nG4NBpjVeFUx42RMamdiSjzEq050TeNf/tzEfMeNNguhhwrFGGB9iVKr3PToNi
GFme9Aj9XmRAhEVC4KaRbj8dz1mfZODt4ttnHH1Q79seA8rrBJnXTulL5c8DcvpaSMvZYVLV86GG
W7RA7Te+V9ob4CuczftOeo6kVCtULkP5XriqJwRD+vpbE2kXTXVzKAKjlKSxkDmu2uXolBPyvgZB
D7kC/gnqrQ5TQ7araIhYgmbQRPIWcbzYWL4z/xzbK+hT96dpL3HD3+lXcX9ZnF1ecm/T8wlNSyrg
4L2GR/4b1GxEVHuu+P8tyRVxq3UbxngyLl0i8unijKSaCoiORLJxIo55tBvIb64jXi1dITNUfy4U
ap/ymFqP2/vy33K+X8zeS8U7IIkWpzxddVRmzKaXJaN7m1iRdSqt1KBCJMkqa+Jsf9VgKEWwThTY
g0vrprVcDoDnD+jx3QQEncity4sGserf/taQDvymfUIobAzet464mFHatLqmruxBvRHcMGI2uqks
0gZTz/Cd29snAM5L+fUR+TxXF0uCq8FNcYvFh0FlCZdDgQ/rJIG5lK7sHg419n4RKy5olFGGVKRA
3iYUzsIpENgVRDHh0Q+qSYhipptHTuGrnqe44kR6xOiwFhtrAiO6FZaorNc0VqGCdsDuNDevHcE/
Udv34lEvbUj49t8tBND1O/88/gzHZmdzh4o3bScrgyBsw1NeColZSHvNqypqO3nlk9clHJxPeqAG
dbdI5N3JYKywkeaBYpAPPj64N9BfsC5noJCb9GsYZHLoRtEenTFVhgkHYzlbjyLkzXUN4yylRDMd
G5lIjssTPODvtpcfs6E0n4NQL2W1CuRX13qhgKFDRjs3o2AxCiqU2TRiDcB8HItNRbCf8JmAXlZ7
7Qemi1ToBnLx/yH4rtylhzupGxDWIgv9CR5y2mphusucXTopqtmTYLC68OveqLF1TlNqPqbm1/qD
fZm6ViIjSGGQvdyz+IHERuJoKfp3+mNhJzn3xBIrQT70X3fxd94NHeKdEW6yNs31HQSldEh0H3dw
R1hLDZNEBPlWhM7Jl4MlktqifDUEpHgT2G9cePYk3Ofj5zHQGk8ApwZGo38oButZAaU9eJeJW8HJ
O7caN0js+2pkbD8X11J4KMOm+fZO/AOTSLCbGOX6I9SqWyPeHDVcgHQ42lrbVVRepF8W2Q5JjY0R
U1De2sp81+8cji1ag0kxdsZt63a4pugILLX1zL4xQR7f6JLlSHhDy82dejl+CR3ZXMdhXqsmnr9c
eboh8n4S1903oLEimDOAiHyysfZjHP3sd1dccWSHmtgnhAVrj+q+K9ImMe6V9CABhaWbTHK1Txza
JBfjXtSlPKJaJEVe4ecwZqOIFKesSwcIQmwp3PpLY/pSaKeUQWkLRO7hIHAe7z+A/k34oF3kdOqq
zHIDH3Tr5t9muVwktShZ21Iwo2TgJ4+Fbcj9SRaB27CIUlCjixItxBNdnMIhJq5KAn5WFX1lrpIT
IiaO/Cz2eMBvwfe9JKg6QxOcC6s5LSkPc7LG4MwgpGBoIlqDZshpQjGdR/cw80oo08YVwxslPD79
6JGccNcHa81L7LSb7nXrFV7SengZUS8Ay4yObZhmNxC842VcZWo7bcPfcB1IlX/Nb1oEoYAVCatE
TsA/g0DjHPEvfn3XdKlcYInIxnRa2+idxSd8xmDvPK00VAk6XGpKjz94HBsmrxWGjr9Fia1MuI1E
WAGsDVviJij3RgrukweUTKXDdHphpH9QZJIpBnljiqxsvr6eWGHZYkgRQoqTsRaQ5mNcUO1MPAsd
7EQXpV3B36KlcoCUDNvweYs0q9dD6sJH1xfL7/Vv44NupirVbe8XTZX7IpmUz+ULS0ei8E87/rCE
LuSRbbv0vEjxMsfVpGYUbK6oAu76Cp0OgD+KdWeV+BLEwbRxIcgtA9wOcXBbnnFaZL6Ww9ZCabBW
Tf20XLfwxUXhJvfgAty1LZWszLu6LDTAiBPFR8Txg3TdOSeFdjNoMuWhNRJs7LugVhqTozpOR9xf
11SJNnbZrxO0tUsjJtGAl0kN4WcgQvhe1/O/DGBxT5Tz3gxLtBHObs7qXCEvKzZ7IgjAHggPxt8T
jx6udGkfBgMj71ixTBXxv9CS8K4WUdq5VzWvY9Q97u+pxSInBXvAFjywLPK3f3+Z5ptCA4kEvT7X
6BZazp/oY2MGh2YNzPWqAGaT5Cb6skVeTgAWh98Ck+iDWxqZFkaOcpQSTsEew6o6KnGgRtWy89ZE
9Y7mQi95zgEpiYUl3mAUj0+IWQzeT6PqTm7mgS6lyxEpvUOnx+b9KEEZxaqtewzTwhn5urY+9R3f
E6xi2J0HboXL8OH0sWfzVo8NWKMIaW9HaPviiWwHWkTmZfgg4Ql9r5/p1sq5SpFb7l6d0sD7ttgp
7tp4NncW0jcA2D9gUMtR/GcQWj56j+owyqT/8vEdcxV8TqjKaVTWL9DrECoZTHE0VCQbOH2u2bhA
2YjZSBoHM37V/87rI0I6UxUxQgY56DoUTfklioB1t3fGch+Zb90ROkUzrt9k1t1mkfbqoubavaYM
+8glebasjQyEVWLi9//lP54JU6cRGGrp9LH7M7ruZ7Qn7wepfvmqnGcjevI2NUcPKNWhqBdM5on1
IfqKBHo56mGKIEs6i+1OowqnMrIx7r+l1MTNnpYME9GR3pneKlTHZevcSZzkWIrW6ab1HpGVGTCy
GNwi2g+ElT3i4JvmHFcDlHL52LNV7FZh3SN9WLoo6kAggpiHQoGFpLBm+205PCs35gC/CHnhjU9y
57fT2Z/MwBAxDHi/BsqtrolF5d+oQ14ielKA00DG6E6+av0eKxWwFyiHIWDcvNHMnkgs9Kgji0Sg
TRSb7Ga6hNHNLGOJIzDxcj+LIhxFBdpfgVAsh5pX4IaLsuo+aiO64jYMmfZw9vOMaEFmOTEXrTZ1
RD+jqsUSqSydmuXjNp82xDN9oOOULTZKAjo9DhjFlOzzCNo7bSOlKitGoRKX/BW3TmhaMVIDrDuM
lmbYEDax26g/CocKSSl23ZKMFScWQ6MztQN1lfms8souf8vt2IFG2qDs7QBvoTqlMyjwATOp7I3n
80V1zznXDDocYz42c3LFIyOl7T8prD0Mhuh/MuuzRRBC09HM4HeZkmuZgcWmYFWSk391PHmRf82p
RrIVCLyh9RkzTqQe5ntr1ZiCbjsjyuPxSDNf9wz1u9Ph/OZFaQLsrF6N0LMPE5zPbg8SzHNuT+Fi
9X9ItlQqJKX2V2aqTi6E2FV8tOngCo4qV7ReF5W0E3UUrOJNqQLX0RAeCEleEhKoyBta3zsQJLi6
AkqaWPFW7xDglkyHBrAyzM7j5s061OwlCwgymyUUGQDUO3UBPnkXNP/0wor/cFPBLv022bVZgc2N
vWiAyNC8oVty3+AoFanW9Yx+JWzhe7yEKzSU3gfMlyOqM9ZEbmXmKKkuduUIA1kBlYfbf5bUfShP
wYDTdPyiFwXJ2MLM+EWq+e7LUTvuepfwEAB5sc2N51epI37lUFI6cwzHZzQFz+ZYMzDGhktoRfv7
gjZteYNHRMYJscXqqBUgSii6Pmydx0o+vGfZpoW9nDkw/ZAA3fSqt+885pAJtoLHsVfgIyN5olxX
8h+glmscjeWdARhkheUGQ9hJzf+UP/I/Tw97SkWg6xIUdNYSdmU6DP/PONiyUouC3xH0YVDFSXut
amt8D7zWeXoa3FCQWDXEqJqJBkMHl7E0J20JrIulFCEt1SAp7FYOKgRlTjg+tm/ktDobJ1y/OPNz
uZ94VvjB1NlL5hkESaMVdOU3ZZ5wyWdA+2Yr8AMana/uP5G1vQ5GriwdTE0raAKbctNEnaIfNin6
8bfpSZvGuQ5fVC2V6iF8tfN85YrEUt5KBgNo9nHywbqCC1UEIaCYF4DZu1GBO5E+hkSE29r7yEQN
obGKHTIvy78ZovXJ5mpsbuxl+T0onxx/MPKtZ+N14r1AnVqVLtpryZsYO8e6t0nFz2gMPVXKKE0Y
NTmo0A4+JYtbXHVXMly8P+rUlNKMh0EX1PfAnuA8oQXPJXY6mEowveQWg6NRnpp2Wa3VWScWZdGN
CRhZQzGblf6bBYvrcMmCM9gb5q6MbHBLkHr5FYi21NHst4naVCUv8DHvqPP1/19H9URevpgaJtzT
JRkWwaqGt+h1HYGoAkApy5d9UrbWXTgLRwHh6owKCpiybww+OOP+DNBx11c+JzjK+ynN19fVaAVL
ACLh1URt98fIX2+crG42uGH8dHz1ijg9Fm/F5KJm5XhO45M1T1hcPQPqvveu1I8uE4rJ5aF7mYRO
KQSvjKrN3R79CR2UbfyqsWH+5o/QBrgh4wuy//udOj6khXNtU/4kvvVrkcWNJqpC6qZAJYQpby7R
4cDV6CAdTYHxsZCz20R8X3PoXOPhcpdXiNr/usnRQ0if55z7zSdZEk7zeDHKVS6obRDeH/N5DJAe
yLk2Pdm+lNAw25n7B/H5W4K/MxtaMrCFhUrR2Z0bTvmWDNk3mZad5NHLhCBpydDIcWArpzkjZg+e
h/J8TQRIPs3VEpRz2/1isk5k8h4wW0g5mLJ8LJ1H6EjLhWEGsy8+09k2xHQ3D6s/Gu1Wq6W273/p
3q0BjYeXolWdj+AVmzpFchVFi1wh836VMYzlmWXT9LuA1FAq7Rt8sKkJRCOjpHaOl0FK/mWPOUyd
5ZPzE6w6567kJNEy0JGl97n2oc1jbNytrXOMEmALN9Kkg0wcU2bqQW6nnayesTfvcX2dXtI93c2C
mWI8mxX8foG64xczGuq8wQM48CwHJslKYkLBSgBFvyUKpvck6sBTVENnwmzUhmMFDR3gv5YvnWCb
w5CLilFcVKrGHkO38EvR0Wa5UPWEYqulDdYE048YWNTOZuY4TUK0HFXMNmuETu3vg+Y3/6SB9e5o
t2yEJt5YpPVw9TIgrPbI0ma4ZGb2lW2rX0scVyDsQ5kntbfVEE31NI9uGeYF/hY44Ng1CJBSLclm
BRzU1tgDWAEcfJtwwyUaXNWHTo4yWgyurG3ZZ4zlK7vMvmlxJEY8FPSzdnWopD7nGjP+jNhdkYeM
yiY9bSoiReVibkgAKa4NCTbmM1n3fqaaEMOlSUAQyorXsGcZKxXmlCufCGyQpDQn/TDT7TjdJHsR
kprn+Z/4Q3KuBotbVdXXfc+3qvUj2KDHIHX4epbGHhbSOvSfB8qcjmrtVvZn/fxBGTe82Qp8wt3r
9+69BK/2DkciMR5pbWP4mKob+QYZUgCKjIFdov1R/p30xCKSbCE9cgJ3YsrEPBrayOExfBYL9ByV
ktnybQjUK4nhWl3/nv8LXeFN3IuzcjtWnDYsuW3JNWPDM6IpQWFesoAo+m1NaTANymBya+k++8rd
eN9zK4nAmdxKwvmfnMbxIdSg3+8W5O6oCVuEyetGntd+5N/l+8wxIIF1UvzH7uzMjHqCISMtjL6Q
F4MvBWzHDOpiCEJMaXOEQ4LHiCiPWXbTTasOv4sotzzFca02OwaUdPgNyPy9MW8MWb6fVknavOgy
Ry0kpeqBW2Y+49CnbtBK11IlU6Y1y0dAGVPjyc1tobdnuUF715kPLSDC6qaJO6VB2gVGW1vSxtkN
sefgNtf66NLmlRdZR0lNCS764WkcnSbUoI17fY8+C9/CTw4nvFcU69iwR7pF3ETlNYaDx8yhiqj3
JpF/6HPaGkUqrlDuN4DzkUaXrfyahtgKpKNFBtyscQoa0glaJHHY4G6cPyNUuFwHwp6P099uGPzQ
m1rkg1STVxXedLurB6MJNUHtn6UfLAD0x+b+FYeCHDrpUBV/4zV93TmmuFWwWT+DnMq4qNwBjWmB
GVptswYlY92dgiZtl+1eEZPn64u1HkoDzToe6K+sTS1X9i0gUnoMCKVJMSXA4NM3LI/m/YPQno7V
r6aAS0cxzMKajaLSPTYyc8ETuMTPpUvyRh32ICLwD5d+YfD+qCWr5AUSUAZeVQLaAt0XIdduP+dK
VGTKYVi364qRWsnd/Amy1fyGPR+mAuFBPMiVjTFutnQWehdf4NmxlWE1FCixavZ4vqVUNkRVUILO
pbk7r0vNAwfojbXebReZV5mXCyN+7taFlwALupkf1mAHWngLvdHW6uruRg+o/61bGW9/GWmxISqc
1r5jyEvV5SlJQJVJzv7UH35IngohefswBjfdISmyZMypj01d/YiQ+g3baEWoDkckQ2ETQH4xBB8f
f6AwMW7orYXeRMN+DPdKeJJ5X1zaBZ+pUUgaUel4v1GBz0k6S/0asfm8RHo8lrzD1YSlSp9kJ8qc
0JNR81pbxtJcjm9cJ07MAH6uXTONuTcHjTaTXw2HdblgDN4S/2gX8lC/Bv25oMO7B7qZT2vewYX4
uueF0wEaUzukPDd9kgpSLPxY2niW2j/NmduN4HuZvAJRrHSugRTcQGJd34f668kaSXzlcUBJLXok
1X41K8pED2BUDJSrUlbmlUEi+WlqXE2T2AVehz+g8gCmaU0xsFJq/XXGf91+hW6qgWZ4EP3HEUOD
BSJZOXXey1PkCDznVsSmRRXGhaB5nAkVlrPXZr5aeqz5byeR+kWFqCnsycznLhFB7kDHz8fg+Qxr
mDlu76oJMXi84ZVoypuRV5Xlug7cLCnv3kpJbexQ8Mc3+TUE129jykDsuekGGIWhi8FQ4TyV7Wtn
+FCMmPCLYhLxV+i89G2RBWZy/LgWDw6DcXFDHpFZ+rQhNhenlrGExgiXXGButlR98MxbwtISr1qw
Db+WEKRz/R7B42Q8TR+OjzRO+7ynnGPC8oVFHhOmjrYQRd8frKl+vSOw1HvcxPLmi1WipMSAklei
+4XBoEaP9adhwRzNca7lvcazJH05DJxVxnwMMv0LOHdRlaIo+DrW+RHdNzGDjkpounNAN08y0IwH
Iu9vrRqyyKWMCpBbyK2S+93k3zGr4uvX8zcoQFazy3Pkn/Q9hOFTHdo5Pf22rx+DtNdhpig0rJ66
90FLQGDw0u0AttNf0F0VcpDHKZxcvfFjKZMzqyNI3J4dovb5+nX511Sw8CzF8JSp2cFNp5PRcy2F
rkJYeyBv/Jb42q1Y+eZLu49FLfLjfnaiQKKtCBwDNAXY3BwI/tboWwgKn2vu2SxGCJWSx2XcJZP8
KREGfjW2SFjK41Lnwl6ev1vMMl4LMgl05AUYxmXbzia+yyW8x1GB0RiwbErMvcQwd2c6yTAhkXAp
EHzi8JSKTTv1l1Nq83b65RL4N2RCpeD7nb+p+jhCV1EkqX2tnwiztWs0i2E0wf7W7fz/ZPoMwvtv
m0Sf8sPe/yRN0NkqpdFPpR+9sx/k0kf+YvXpjP4kf50s1Z2Vi5TUF4yXwA3zAbg2n2tBIWDajszK
a6tp3MUgiTUontk8HfNT7HJCkeRsuF9n9Pkd2WTJNhjAXrTKYdP6qY88n4ecLXYipMCDJQg+Rmxk
PIijAcAH/qJeWQ1T3vs/+mh0kg0pATIlc+f+JkqBKofHn+D3jgJgqN4RHCaZr5DI+scovhq/WpUw
0gpQ1/ASJLINM7vGcpXDz3AhhwlTxmIIOM5BVztupiGJmDx23yLwbFiUTTCeQTKQ03NFpYNI1vwU
ZjPmDX4dSG7v4BTRwEI4hWwr4+4SdV/vDxz3Z2O1YlYsXUMAyYYhBxi9dC2HGiWz4Wc5kTeZ/Bsv
A7058Q9wT2Fj+Ou521oyQycz+C/rX8gKju/Jtaoa09WHTMm1hKWSMwobzdopNbwHWaRoLm6ms4sw
i0tvl56Fw5I0biOtgWxUgp7YLSWfRqkUAqzkcRIdGUVVrTaKYXMJTCV8MotiSRptC/I8ajkVlgpu
XFvJwc+mH3mxaZK3mlnTjDLrfqvQvJTZ16DlNI3eoJXcYctnywFiVoJ5RVQxpwPaEKPu4nLWgsQg
ll7U304awgf4erMjblgMtCmwiHIZRf3mD4hfndUGeSMxueV4f/HTrxStSWCHTOIz+1FTfmSmZZ7b
v0KBHzq0U1EOvh1has377YpG8RVrbbWRcF7h15+B442mA0C6OWcTlfjLgeNSK9g0Wk04QDGMudSl
OjTi9emLtJmu3LQBoMC+6jLRciBEDPCgzCyRWfgZBj2jNVWuuHA1ihXMa75O7/ihbfaMhYYVg+WU
Pq0iajgzK4fEGYSAY/Yc/9NwIswiQvNdtrazfRaH023RCdG4W3qIIYVA/CLusPlgOa3M28kZH0ws
/koFy0xSRYJrPNF6Y9qLlt6kD/6/yMZ2nQ1Vmi8PSlAjGU4UDQ89ccryAvQaNqSQ9izODqhu3j3m
jP+Dwxy1pbWxz8i6sUfB/1YiKOBS1xPGoHfcOD0XhD5F9ZrbzLCOega31uDzFmSe94stvdCTCopw
a1Pw8v+D/dcDSWXih50J4NvhTf6CDFpiuXhvuVRiYI/dviMYZof+ysOWIwf6H2jWLzNWDHBGUCwD
f0nuz3q+5+8uZ1iTFDyQlMtnmWCM7US66imb3bO5wjFaRaEvvtfiJcSE7xLyjtxbXHM1+0IIoHIK
Ws38U6gVCJqHnNT/NsEB/c78+1b6pkwIwVryw2ZdRtz+smBGCqmNvrW4FkZ+DOdlJkgYkK5MlYdv
cLinpmj3IW7kmSO2uSa2qgqp47xexC0aaMx0gLbIQ39ZWeuWVbYR9w2JuLiewgTTpfjPoxaxNgZW
19JgHgD0HAAZjXoaJpnMWc/iV1gxjWZ0iKI1Rh8UBG+wxIKqD65l5wx41nJ2f+z/ux1M60QDqkad
JfIZAiJMTWCAkkUpS5OhdGlSTsg63r4cLIiayzQtf3kJUTnX5qOkar2GVDDT361a+/CDBkZu5mF1
CdcJreSfbR1qDWtqSAjc5kJm8PhnIJ9VAt31MEo65lIbfhvvfXC0wbQpHv7MQE/3+ZipUfmNvESk
IJzyNjOs04NdGc/O3qpuA+iatLuquaPYO67QwFbmHo8rCa6Vn4vFfz2Zt8tU48c9j375gjpPVJpV
uws2vCQVYkdVjQ6TsGv3wgFi1DGgAK75z84/pJ+cjBIFeyG/vVBZq3CPRPl52T64xY5eCftlWK/R
4+zaEtbs4nnB95IiVPuFHYyG6FW+f8CtI/Rexn6A7txoGc06dkdlqL7+NLKH+Mc2mCk7e9ZBX2a4
3aO/ROMLocw9T4J4/9FAZ3e+dgx2vGNTIhd7od0UsByC8Lsztfhfj5DqivRGXWwR9IXLXN5ZzNcE
vzGzlO95U6Xn9YKbJ7wtCRHwOH9hUfHdHFZ3FHtUpqRwrHnYIymE+48dnAKsRC/AC3ArDx8o8lVL
gbGWbzVzWKJqaaAV89qJZ73eLPPv8hbuAHvqvkM8EI3FW7ZnYW6Zt4HmTk1wMnRARA0YIil+9Ayb
xx242ryy71m0Ed22l7e+0hhwBqUKwgAGsj5on697S2ELYoXkHbrUoXj7M8NNNqZJGOtlivyAMScO
zwHi745OjRqujaZOadZxcBcWl0IWEMD/uAW2uR4x404GeopTa96OcWdMJbNG8meYoPoIeihdPF5O
NrNLNOnRRW9CIy0v6qzqKswEcX4pA7z6fGkbvHl/CfEbnwPe/ao42v0dsh1jSSVu/tC1aCBSP1Jv
0Kq+HihvFiLJmPrJPdfzXV2EnIvTHG27EtJ81LM9I8iuZXny9KGBV+WomhbdF9AOutjFsmN31LCf
xjPJ7lwXKlyWBEhaqBDjj04+be9S6dEn0Sr7SRwo9dQv973DablWxrh+tVXckeT8oU2FDmzWD8U3
5STrW1N6ajf+/PFXH2B0q5V5JgWxjlsFOT4S3s97SZrv+13mu+XzVSxmCeHgHJ9mNhh++PmEO5JJ
grM8V+rceWi3J6koz67hDE01upzfsGEOobmLcH5VTJhSDNgvEuyH7WEEb2Q7KHWwxQig7qXVnyA2
rC9Yy0OEaJgKpYne09BJKNl6wemmfiLcZwREb8Um2O6Cmnsw8I2Wky2KclzX2p7+fQH5Y6ZHQC8G
TFnAJts1SPtEdRLVShYa2/RBgVXwrnXblUQ5QrlxbMd5JhJxrlX1YdcX44lhAeqQTL8ppJt2geP+
q66QfNz0RgSilj9jyuOwqIJcljOlVqFdZ/I/tXkMQme/XZf9IChcbOOG+HkbrOHxwVWFDYHEjMMb
zkXXgHfNuL1Asa5VEnXu/reXJaaIkbqqK3pXFI/egqxizC3cGDzHQxiyzro4y3QMbeM2gW38fX6j
0UgWEE6w262qg5FjTx9icffpHNOaIhTpionZbBIbdEUzahmGn5XwIUtKbMf9rLdcQpVCGV7qlgrS
tgcsInf4mp+0W6Xa3H7QDyJEJd5ARS13E+DjRgMQTQ6MCpGK43CciEQYNr9bgIMGeDBJWd2qTGx5
pCsAJ1OHZnnXJkm9vJGT8MYq5cBV0xMQeIzAr4xZXwp1msjMsg0IQD4FvELIqien65vknKHr07bg
BBeKcQk/Fme5Wvn7Fv2aai75v+QKlufdFBsWlvGn0D4vZSrKfUAeiTPVsJlB8o+m/tUEYrxN1jbQ
kCLOK3ckMdTyxWP99epoRj/eo2Xy09V3k4rX8rUxyMD+uEbiuXO2rRyqPV5oatRqvHCv1fhoh053
0ZR9x3DIXRwz5yedWKiw8dS/YglGc0+4TYmUYkN6U4IQDK9C8pxtAoJc+AbGHuyV5IwwwegnZtSd
XWGShml9O13m8d/iIk9mTkVxxvmicgf2dZrwzV+dE0WkDnQDcMD5dW/WGD70YUbeQ7AyBQVzbM4H
WOO/zgg/GGpeg4pvmkDSroFItB7HRw85V+KEiGcIImuq5FyogTO6SKk1wJDMPiQJ8FsNzzFii5mV
7ENZIcnHEFMBJwtWG/KzQNXNv2dKnUXQXMhhRA2N0PPW2oTW6Bhx6PgX1AXRWPOQu/6wsBqh7xai
x3oHlmkUVVrXXajViWp6mN98ro7+sthbsycieVHOW1EqVRBMmdIFCSWxVadRrg84EHATuJtvhVcO
bRN1bHjJJD6Oe3A0IIT70Nqi/42FBGIZ1r0KlAgc+83wfGCmTDRWvWZuyvZddZRo+mGZxPXn8kA4
qptJi57xj5LXt649O0ElITAUJDJXo5uZT08b7VVrEvm2atDwOGdE1lKSGegGxDbaQeXurYkaDS/S
R3NjtaB2ZC6XkghTv9xqZIRS9vCcc4MGzyP5xbu6IfRG0/Ki2TAnYxRgPiDcK1ITF0sACzTzOJ8N
SVBX2qtxIJsr1XMqdv6USBI5iGdxlSFUQ5AFd6/pQzYCZUvUTXCedqKq1s4nTmMpvUxNpKbpevyt
veZdfYxT2iWV4UX98K3sh797K2SipKtOEANmkVI/ow6ROAgS7JlC/WWPGYlYIGGl2frQE0B/cURU
YQlRs5b2MuXNe3ExqBdn4dwdzg3Sa4V22uDyNEI1MvKWW38SsS+Gs+zwWGpdCAcq6VjIbyCOi+F3
ksegrRpp8mliHJdbkxMPqVwz3cms0urTobBJ6FhU+Ai7KR90FClp1B+jQV8R+DQLLIaq3FS7fzxS
thX5R5BzXWef/L9etGhgmXIA0s7rE92M9YVDOj878AN0pI5fNmhKSiUChBDa+Q3vBoj3byGhWjMC
A5q/U47xqo50D9bY+mkY5+rUAe7/SujLYAhx1DwmGhTxT5yqZr6K0QUbfUl7NbTn/4/Lav2zwF/i
AyPf6J4DAbFSu8Ignm3nPZf2siMqmrW26u5lN/Wii572xf8S5H9Hh9m5GlvcldqgJDFyVK86lSS7
IhRS8tmIbTsipiPuxhxRTgGybd9MSMExC9oRvwfSp1uFI+tsCR5bRNEdb96GusPj/EXTh7qpEZJZ
NHOZODQ6saDNxXKdQwSVhV3nTLDrA5iFDJsPoAICxDSkj9cTsTeBszmB/PRitEw8AVY7IQdMO1Eg
RufrR9F+bDdZyCBGxkcxplqLG2B8pPFvS1q4zVxu5p2sBM62igq249aG1yG9AD7DU+a3QubIsKOL
Bxhie/TNfsPCheJ8qLvK92+5KBB8HyluUm+N8EK8D2IPPJoYzgIo+JSUnyNMfOw+Rd5UswWb3i+F
ADSiJcKzT9JYTyL7tWg69PdlatqplZNyW+zkdG1WdvqqbBq6wls/oaV5vrIQOPNUO1dQfkJGi3fi
KK6DuCPPDhEFvJwfFxIN1jOBihtaAMNn0HzSTz6IZ4TjpfgGiFMN3+M/vAuUaaAb5dZKX+hEXLXd
VvluANVsMWQ2p9ZLlfGyKb97FZ98E2ZgDD8uEtHNG0cRj/rfOkrGv36Vcu2Gl6oqqAPDfxk0qJqZ
zykkKY3FdWOH0+xMkoYoPXhJgB1eMntTGJDdRlmR6Y//ZTbfkj+MswWPHLzizEeWAN5vxznR+n3q
FcbhDGhQXb28lFM8yonmfguFlCeqnvpLEj+EnFKRvkQ1EWabymcoUej0/9PsHsu85S2dLwoG5J4/
4+FKZOTQCdZy3vM9VbVNtaZ3z/5jZNC4z93siThmwt4+bmsVUOiyTvv61JfMzvVuaEm+TOjBZtYj
nUw/urJuUz0K93ENNulkamZUSTaY6NIb0p2B92TCWswqzo2Uc+iYz+NtRWadGkHtDzVPZZFCxR9b
3Iq1nf35j4J5P6owQ7PuIgR29OWONo/dSikBbXxi9/iZ/T60d7DatT9ldJ5Jl4q93zZ1xS70aAuh
GEMsAEFFPHCr/9k8svAgie2kLwvve06hWeZY1B9M2RhqIzlxOENemFnfC6Ot+1udL1IBr/Rrr9Ll
IaPabLCISz9oO/Hfn3DH0UUu0ZPK1k0INl56vWbIoydqgTmmWacCLwtr2WzPsAG7BGBA/m5ejhf2
X3m1eInWdZx9zeTMdQDNzSg6YnmswMVnWf7LFZ3Ir/vFAYYsWR4VukdIbWo9N0djq544ZRSIDR9+
mYnIAYBbH7tzEHLjHY7PdweylI++yYnAtGCUXbtVCM6ZQJbS5aEGLM496SQ31BmnkgqxmToUQxny
SCBxNm5N9t5VeDVgk2To7WumcKVpBvwNh3DfwGv417BEEY/3sM1eI8zoKFZavJFfpCBNcVmFnW9X
ceN3HDZrzH0+54yPM63QTaPse6sikkf+ucqTgk243VMAD1Mn+UE02SAbGy6ePlj2Wa3P+d7D+6r7
LVWH5B3Qv1MW2XkJxa7sEcHkknkZqd7ROz/06jl7Kkf00nbk6vMIMrGDMG5Oxhy2GAqjyw6AIgca
cgEjZK18DcHX0aoy+HlfDa1X9Dgkm+66LPdxdJyyZSODapTQUZzpq3g15Sl45NT92YnH51M8s30d
8/L22fC/MOkD4Xvx7IYaBLy6NxU04JUUiA/2Pe3boOPeeXULivBPS9JU/d8FDOEWS6d6jOumZBhf
swduDVRRrhnIUNMaEx/674BL5SqXqoAyo3qP2rT9SIXa1SMw7h0Q0kVYhsY/7fXIjK22VPUAXonB
lcrFrSq+/tuYwELmG99gZ6YHBy5l+n6z+1a9fL3DpDgSkJU/1ii2KVQht5NGu+LJPz/CzL496/am
s84W2NVMLHmjE6wR31F9IjrxqiEgLUKx2QTNmnYDKGA0MWIXiEDg7blnedqgzrjBs2ywsnd0n39a
TIGbZBzQy5wVdFI3slq0EG3HMnGmTPraR5U4iTBFm1hcfZl1wiwA3ZkcEckJNdzvJeDGA24zoI33
Xn/+3y6dIfdIx/wb9QA20Km++y9faKamJubbhvUpuQZBKsWcoYWvHCz+QYm9OnPB2HJ1NxCkMYX+
mSPwmxC3SBK4+nGOjvqN/gpQzwWgkBLvXi2awCZczAVfRZ+L5lB1240F9yKb2S091aH+1Wy40vin
RDwq8B77+AgCSdWd2qEac+H2CZ7BaH6OdH/nuYAC5+CFA/NYjW1Wri+QIaTThAhQnZ3b/z1e031o
uGpVBbO516PKkv6d0F3WazL1yJ2Hqh29fghlxrTdbT2tb/8i0Grq5oAA0XFn45EPkK5C6m03vf1L
ajDJwftBFwBFJTTDiklc8kibCSurebaNd7kwa+M5y2zRNZFA9eD1rErbU+qHijE4uzF282CwQspZ
2GzJlxo/HNSHQVcS+G+JtUpDVOwCKeLXuGINgdVM2jQuPscrb0iNiHGyatSvc2dAwfqCy2wN1ifj
2YzznZ7u2Wbin76dm8Z7tTKiivy0YqQx0bcIdTNBMQ+yIlWoj3bbRL8Zysfd+pYBeSXyapDeQbUN
UZCtDtD1X4BrUSQFl5SKw4mYX6BQtERQI0Q7gxUHgO0K2Dn4ZvNiFrGH2e+5HOH6l8K1/A3NDwal
ipzV6DmwBuGme5EYRJSACXNTTE595dETTqO1OvJOpL6Aju1X92kgYmZSV5UzYrLoRFFmYgDTt/sg
6kKELSoq1ygG5mh1iohBPBjI9jWY8vOYU5gUudQxnzlbSl3AKAvkxKwU8YZL6F+IgixLG6+o0vr6
8Sp9TIvHORnwTTddebP8Pj1fpEWQqQSVF9876CuQ2IOWP9QG2kw9Ws9P9ZIhDiT9HCBLSbjdUtRg
Yt3kcA+IhIj41lQgfWuBJE6FjNq3FkCad7/j+adMCV+Uyib6vgUjdv8DfkgVW8wkx6uhJQODlAu9
AoKWzHbAIGJMwXvJDQlXZ9jyJdn4vuT7beJlx3bQtDLqI/chkA5N4LeUFgaj57bRL9NX5QSY0zHD
8pI2BOm6Rp9/+TvrgTw8mWgORXkBw1Io4/BlKnr4jne+cwseQiQwj2DdJF9sHXt4EiUV5B1/9yby
n/jygWTRYkIpE373FP++5eNPpjIFdQ3T+tTN6P64gmyvHr0XY+Fd6/iEDqCEva856xbba+46vv7v
dMFyJ/6P632DSRKe/cNCvINH9ImGRYTBiY5MhAciNwJh9DDuOBMfx8QXx2F8EZctZYMk9pa4JKUo
mJLCJT5aZ+RNpBhL0MsQ+0VzxyCCfKH/2p7pbBxpCKrjh7ZmeDCOhNZmuW3/kSX0oNE9OBFoR2OS
ZerqUl6dHFmu/nReRjQFmhsLl2M3LAxIeI59Ca5IwzSxFZvhobGQuMK6lGHRhGH0GObb20XSUgW0
Pxa9zE5Qd7a4bqffFJxlZ1E63VF7SbnGuxiqZO/4p1eldh9SqiAvWEsn2ROf5kyP7NRMylyTq9tv
euvzJ5lko6bl3rjbgOF5oRUZH/BqYrcbEXlo+ybwajlAdGSnTM48g7Ltt4Hi8xWotiJvuKweUBdu
RC+HqeBA/CBFWWMZGKuMc3x83AKHI8CfYp/ZdSFBTaowXxaj5kfhf8PZlFG4I57gFkLLqdWVh8W0
MjknzhU9/wqnRupbwH5V1klZFZPTss71BCuzFSJLDVwg3ddFtEaO6NdDh28im1uJ1QR5xBApOPAL
8lDlbjV8RitYBJgm1m7GXhkGeTagr2NLuG+5BV+byNvKh1uGJk2A5ce5+uWxDf30CE56pwrtikyC
+ILJSNxyo6EeAJA+9uPWzm2StNTqoWzf8+8ScA+aBf+s7KCuwcd9j2T2xTyThWrmp93ozn2hSuqH
rHvI9t5k1HJGTHy33vUgOsryDApKStTMCMLxb9ZhAm442PclEQZ6/ans18hPnJT3lD9VjrtCPUsG
WwpjFnzVGm44zMHgRfA/fgaitJVmwYk3qc9KMQaXvwaFICKIhw7YjgZ/RYGzWBhvzCReVdfwvkLW
Hv7N1pTBK3sptKZt50pLa8fMA8doNwVSGYQWpmyJVl3Jx5T1kqvzJJDcLygbFwwl6fudIo7v/3Sl
1KQ7JmSVfuqFJT/6HgTTlcqSykWVpOdXc/1dSbBtuZsaKhd2KuRv5RLD9y2IwtG9WVPgNxmIR3Oc
bJxwm3FBLq9W8X2uk+ajJoaBL35i2XQPygu84A6VVgnG53Lh08waEmerxjHmLu+mLrJSDKUjul1i
MQlHIG2dB83/tHlm7ClbcW3bJLqSOtz2DVdL/PyMy2IrRy+GfSGYhq/bYBaIqxn2/us/N91VFUXk
ZWrjuasXtz7aQzgik7ZKDwYF+snSLGVfBtPm+k8t1qh5wL2sUAgmf4FcpBMh2tLFmSZykhuU4ZvW
Yqm6qqkY2Y+seP5ggBTCVCzZVv87gSPioeb2fOHEKXwXRmxAdYffTuh1xT4BmxKAxv1BpmnKUp8O
mjKnNxQi+mYNm5vmEO919YoaizqJedZncLnpCvtvpb8OuK1/1dSFEs9cjkauhwuMTk0i63JkocW2
xiyQA5iwGW20ztmexMSgESB1s5dytsD7OHHfqPnE8Rdx4ZvF1+ppWSTCBiQ6CubZSiu+2bXAe/cZ
jpTamCR28qrDSfgQPrbUMBLNAqD0XXBtR1a3emqglQZgtJVY+412IKXcslFJZ2CBOSV46klovlnu
mu1z84fLETzvo1r7FnPrT7Ycu4F4D+Rrv4KafVntuZl6uT1cAYy+DLnT699i/GYyWii7kxHdKI+a
RvapU54Mv/e/vbPv2ymTsMx9CnSo4zgGAlofqZ7PGq7+M/Q7swwF3K4cCeA2uqOD4AbPRE3cZ5Qq
oreD2vf+ElUGTwtSPvPz/ZwAPzM8aXgaalWO2Cc0VCGQBiC96jBxmW1eRuvTjAZCqP4iQsw7cX6e
3jJT+LUIIZkZNW3Yg+XiuYOTiVzABhCSLszlS4dsuyJqfTnhHRkMMgNCb+UHneDPzHQbd8mvk4L8
vo78E8UOG5klokpkVjAyYNpOTv7BGoMnqz3wW2gk0z7ftlNWyg411/0pw+rdMLr+gmEc5wBAmMtb
4P5sNPQvVgCkAWBdj6CiJvUxkBrixkxYlTwGCepn9mxH6URTE0hAEEEGqn9x655apLe/khLcZkKo
4FYy1hGVl9rVtTxtZUZBFuGjUotM85lxNZrDt2/67ub3bZZ+bmhMOzRnut7RpEPt2wNGwOMd1IYt
Lm6DOHbsp8XhW2QQSzKstHc3YMp5WlTw1cn6SIOU/66MkDycZYc59SlKok9NAFomFHGgRlWSOnvG
i8paXQJaqAr1IWY6N46TVrWXSIyzeVtxrWnTuEbyRwaAI3Zv3zkwRVWO09EgkVOSYsc4nJCjg/x6
Fv2EJI3QoLqmfU3sSzbH+CeIQUxsrvnE6Yn+xEHPQad7kHRO53dY3/v7kYPkEOQHOAqw0dm13jJe
tp3WfoqC+gNmGSUaPINoPoehwT7yMBvx0Z8yd5cL03pilaZ+v9YvfygkGnJzE6Ye7nTc5SlLDpBh
VEaFUlLLSZ3QtPGzaVhGeoVDQXvrvRGZ7kPW7bDx5Vl4W7Pf64Xnm+aIoBXy6nla4fA3CUcSBvyd
llnvP+8oqJAGZBq/O8IERs8q05GFieuWk1whyF3B2hX9VK9qfPvC92fCOtYx8oqruPHuHfk+CA7/
p8eUu/Ym+s0yqsvyXsdLb1B/vIP9I4LuHodj+FiaGYxuZ1RJUJrkRXMjKe1K0ogzY/v/+lLW8fbu
nFaGOehG6FEc2LGtsFsAHH5BwYnoHIn+RcJdNl3XBxEWtBZvLCghYcnyqVPalyZKZnCZy+NX71KO
3HdF7aKVtZlixD4AN6UGnRMBnRxeuFUqdmeQVmN2WMvf7/IUvu9sVdLSGKODYXm5EU6IA16QWGsH
OebBcMjHwHjN5A7eNB4M7RIzyaHCowCwAbVAW2JbEjdQT63gL8h5pxAtQJH7BhlXovi7DPzv1yhw
LGDWRkFOJggldm7l6ZMmX53VWWJnJ++DlyUsseLdmg+/ZYsHIUDCwqKzIrsrlJUWE8QaCO/tShEv
bKNku1f9/lbru/Gtkm8P78wYjRp0yIRiPleNOqYmNC3pWNVmpMXarurmKM/w3PNhuQbUOMjS57Kt
eMBt9KAU1NaoR+lvmdB8sopOs4bVpq3fPLh+dHPRVUp/aBpXwQ3ofs4EE9A1Xaxr48HpX0an9IET
4EhASqquDAcGoB2qnosnw9vpim44A0bdhnwe/Zf1VmePSSN0kawFAQG14a6BMmsEWdyfsHDKk60d
JBw7bmPmAeqxole4i6LqVu7r2VpfIhMwvAuF0w5eUzu+cSTjp4qBgntgt/IKvq27yLCHeu/jOjWB
hbqKt1nNlo4MYQ+hk6P3MVgeN19TZWQk9kh49Nrh4W8Hzt4wYsiOEOeJKDv4SMVh+GLrHVNxubv1
IrMnO5BHkNm3lEAzPMHUBafILRvdo4X/K9iEqdBbzIn0hAmgBWpG3lt3s5OZoU5y6iGjj8KEop06
1D7DvSwVrpZVvQH07um1RrCDBoKAssS63lHVqaa+226NZzr0UZvkU5pp76+iyhvY/SLgopjY/Tls
Js6c+HEdrM9w/mMiwIusztUHhaFKm7koAiICQjGpmNbB+6rKTTK0+Z0EomEXq2b6M3Y9sSv35gyb
9xjv/vCdaUKed7b6/Ig7PD2kWxaquhdRdSc1gvgJvPpstxKcWNpyt24Y7mKVc7olJ5NBFFCUmhX4
t7F/jJ5pQRmVQhmQArY9rS2YftgmrnJKDJJDubuuJ0JC6fDm6gvKpqXv6U18Tx1BlEVKcbQuSqnH
AXdubRJEbZBO/AdBmQtHoCM+ct5SnohJwrvVzz67XURqJTTRlxFVaFx+aXPrNWyMel8MMJj/cwET
WsNln/QwYdoG+f531FyP/sNWOSp8890yWMW0wJd9Ji3qdNvM66LnYncYQa2U1TjsXneLYySPmN19
VXaubuFHYvj/l2yechOZTH+vqhgvz0ffKpDA877F0SA7GKIQ35VVOFbn7BNiPqMbxnDEK0Hm2NDK
z8Lf37ZPA3W7sOWCgWAxKC8t2HepLtulTA1vQnir99oTTTTwaxcUyQzUHCBPcE2/88Fl0NCVpxv6
smbqJlINFMDqFBCWyW4ALAfh7LLljN9edu+8CKlgrhazefUpABEjGiD33ooyDQDvMaPUCVgvxtvU
0YLgjb3hRc8rBYuIHzR8E2eHxAMeqpGgofM2nKtdjs1x6Bm40YbDG51/y+i+0NXCv5kTltz/aq24
t74VnqZraKOm+bWrnXYXI/Q2cTlwc+6zvs2pOMK1lJqMxOpVX+3BAC2Tbna7NeF/3f9h4SCLj+N0
AiaUZ2tjOhdagfYmrvNjRKene6zmM7I67VmiNDZsV17I8oweZi0cz5/2EtfYuzVaud69yYNXtEhM
NBTe/q57UJ01kz4PL66qg4Qj19vW/RaV0h7xPmQDqiWkbp/9ull5jFLXHAqq6o0jMyp40011Y0XL
Qb6s1QFExoNXCD8/qqsG4NfvE9amgTUruKOMC03Sl4wHK1qjBoAP8kyuCLDs8cyZDGkS/uKteksY
Iybh9W/FQCt2ueCFSypJHAMGTBn+xeDYqC49APpB7uT+g5n3eeBDhyM74H/3i4/NJPvfmEzKGi66
KbN/MEnALPM5KeiznkjHMo7+Cfco5bKYUUwYCYZ5DDxN49bNRG6i1XZjWha4QS4Yw+2u/niHBEfr
ldHdjVMqd9Txvy9ckb7PX5J1JnvQi4aDIS8nC/n6O3SZPsmCE3Z7tJWI0tP9DyffLvljNIR2Ylzj
gb5ub/GNNef4EJZ1LW19CNiNCUCCHg+yMyLnbc0xkcIO77YQdSnIB1dHRADNt+VcAthyd6Qchh0h
1Nmlliap1e6UvPQrA8xGPjl62E80ufahBSvM2Pv1Gs6DYsptrKzKNLMGwdIgJ38aLNx7ghd16v7x
VQhH9VPt4fXeOngeR4r7/gg/lBvW97Qvyy8WTuI+BCu32LnWzWnMr0s5pK0XeV0LiNnpWIWsX2iU
dKn0WreMDaFo8E8I/3gyXVC5dZgaZYSjqoqUoUM3NpWeKlZMVvpfNO6kkIfIGamFgHOw/Pj1TuGI
x9lYGihVbZ0ykXzi5haR1I7YYTbb7559sN4SIE+VTpzIZiM47SFPNh4N4ea1eA1S150HxeEmApTU
0xTqqt+zsRML0cjpJDmADm+BToD2YGvbPibctOXUK0V+2f4SoKhsUNr7JHKUKTlXmUt7ixtKLjTd
vjWUFynt6TC9fgIRa/5onywJH3sKnmxQEZJhJHFdG/mvq4e18VHJBwc7UuU8TozQhvN+d9HMDV3U
aSJMHgWoIy4/UakkXlKLThDCGoBOuJANS0s3fKJXUdzUEyw/T7l3YaunGZiX93FcRl5qfXnybjuC
X3vtDglJ9eYwIZAdxGQzRFlvcU8EgZOxQQ92/lJI4QUvkiQ+3Hax9kwpk5uKbk5Z3k4TeDdzRmPB
FNkEdPQVv1xoKFtCdj5I32CVXmHp87pk6yEAVYHEkK6mMSmDDJSMRSXt7BV/0GVLfCqDESEk3ZDA
c6oNpUn17HdoHsfNizLlZfjbbhT1gi7XarorviCoT2U2hMQD1+e/0vRBZrPMN7mQC1gity8P19ig
8yg65AQ9i2TLOEe2FM0JL6oD6z6ami9zLX4jAbtDByMO3mMtGCxx72m334yxevar4J1YMu2ZcTsF
9tGXRkCIoC+TJatRg5a0MFhMqrRGly0RX7cHq43of9SOSdv8zV3eG+BfuRPq8HbANz20goHfWxSq
oBvSfrsrVW6wZJJpcVLrTl8CsAAWYyjU86s9TwBgT10w0pFFH/1uNvMPCiUd1cZy4VoFSwEtyYGn
XNOzz7Kl0KfpGIaNL7SbVE6IbkmtsrbzMOXisQfPhqSvaNz7nG4saTSjzsjMgwwt3W4lDjPGzWv/
Cbdo/S65c3CmylbZE1uTXvZFZp6P+Zt/U/7U4AypDA46d3e4qbFpF9lS09ef6m5QTAlqlWMRiNWF
Hpbf+E9CgSOQ3DRjOq6G2sWyvjoskdLvyTwm5J7Qw15RtjmzbLlG2/NsLj3gQ/z1CvZsdDhciTad
kUHlvlqcJTgcHj5GXYd9eBRi9BI6OgRUo4ASez2WDuRcnAMOcybQfbxM0sATsdGd0pJrfph6k4RR
0ke8YDJMRNUqiQij2BTmUXX/xH8APjYrxYtodxqfW7GW6GCcy99uGo8RVBiKe8stVsKhnRfO8iTS
ldINU1OUAo5dXK0Hzda7CRcUJ48osqTEbSO3A26vxmEpe+hembledgJImIEz/6IOH3eUTVvYzbMB
xjkHEOk/LwnJIqm6e3Lh0TWHNlK+XdC+olnoVAfUCrpH6fMpU0sVHGDIn3ilPvOQXoh+Nxyvrk7Y
IiHS9P9JcxOE9/6GOeBvo6M1KGmpHZZxhO781uZd7VEOaMEZq3aUp5XFOHD5vAyJ62kmtMrITHcA
j2DiaA69NzvR2lpswq1kz+hsmSgwIrEpZTqptLsQcZ4nfDilsqUNGEJNMQJhoJxdh98v51gozFFH
LPfIy0WJk0Esrs+FLkjapCvyad1dGKKVJZRWN7ObZvJ8NMN68vLnhe3idTi0kd1tPNRp5vu11oN/
VcsG1XheL3lmOdvsk6d8m3tGM96vlXwTyRUwHo93PPXUTEXun5zC886ECfzYLV+/BacjYA+VN3V2
bHutnfItW/94QBQC4qsZZDahpY6rW1aDw+bjt5Kn0Ku+Z81rOkA/bDliPjkc61WWt6Gwy8KxSzMN
VCYR97VSmN9bAmkoIIYm0LPqjyYOYpPifLF+NTtz11GOisLCq8ak7/4v/HCM1aeSN9//FJTPFgVa
MqaL2w6Tvt+O8b/bTpaPqnseZiSf0vrO7fPLSDty3OuDeyEpdyaRVt9wbr+UbTZ+mK3x+weM2Cez
jV0lRWXM7yTSn0nbwhdIweaQoJEjlXSwpZnqCVtX03dD0uG7skesxsB9pD4n2bdzaaSIPO2HsWcG
EkElioGIhuR8/klpoepCohCJEnaprI49FVSLpiUqt3GBr4Mqjg7aiQc8z0mkX5RCf4DTTW9xCnrm
UMwGggY0plEYAAXLH5nf/JZyRfZ6PkwlSFTEwfLBB3g69tGiy66YnTBxQNbIvbnLjaGNc+Xs7PMX
SyMtvQUFwuLg4fSuCy4JO3rVJR2rNARElRgWzXrxyaZSwiBrUMr+dc7wIIsOTSUNeH8ngXTRHWB4
Y07CQs3DTP/pwlae+oAjaqgO9Ze75ZPZANKYxaL4vmWEDNWb5OCMMVqbPisWfWxgKMXvsT+jLP3I
w1CMb/mdvem/d+mlhAHJKO4CXjJyJdK6uUFmdcu0X7SNM8lhXatLYS0Qw34mfwKJtrUU5P7ISe8P
4eD+4ceJTaoD2zmKksxVXt+u8VgpPovk8V4C69DPMXH5UahHKk/p94k59SqxVeMCcTlanPVaapiE
RHGtgY2Zq6YLHwZgl1a7MvvFmiC57v+RVQ/1rtQ+AtOvvGMh+TdJmeEiRYTLBIB55LA1edHaZbIX
OYDG1WS9mWCPJDa0B2F8jY2tx+l9gcCDO5Z1koGWIK0N46fR1Dhmqft47r3UXzb5JDwGLSgEFJm2
fvmPKDZiUSTbPOvVNU+i1ujZ9/6Yz1HWUgkrDc8jMZKL1l5yu20v+aTNsEwRUq/A0GRR3k4NxIyi
X9LJobkt6vNCpfiqboLGtAJUKGWJ9Mii1WOcKwZ5PwH2WzE+/2s4yl87Pbcxcx+r6inTOzaRyhte
zljzeRTrwmL2HZ2/c+w4jpFWi1GN7KbCOpbiuOhXTUIFG0dX0NxU/OFXcKFZg9kEhQk4vQT2b6O6
Jo+XoWuzBrVk0wt3v7zxr656XSaqitJi4GhL5ooGLbm2EZcAcam9gtxj6TxjtHnAptAib4bf8PrQ
2uYi/vo/BWX9L04UzOfYaw8jJTeexZ0pzs2ysbCQ0gC8BqmdzuTqu2mhaqMDL3QN9/K+oZI+9fXn
ua4wVHfKcQpzBo/p39FD0L1MCRqKFT15oInnrOfCacikwqyhjgePSnw590M67Sxjf6Cr80RLYkm1
oNyDd+s73GSkMfFant0M5UYEb5NC5PUg7siM3AGW8tpuz4U71Ij7a0QWuKzSXawrrckzIjvjkZIH
/W//nbukAA79lGDmAyznVsXZppj7hTyZAmkE1yc9U8f/hY2Iy6vCCK6BjuU3ooJuhkyGFyl7b8xn
W8fs5Fhwv9E2WbKmGNYFZ2Gk10hYLUY6t5NwL+w43TjSniXvN1pDV3kykOz+OmqEu1rB3rT2Vn7/
NK13zW5zYSIBdBBpgmUHbn33AS4a6j40Xc6GX9gM2/DgKreT3sjvqIH+bzVoSMSaY36cV7DgrWhx
mq8ei3FP5Q/Dv5msnvsbFYuZALSCqXGdI3xNM4r1VVR5cXlP+tKdqMh6f5hg9KVc0CfMAg3UgMcF
du/AxM4O/rvA+25+Ofapqb0prs41oS7P2MtQh2a0U8i2OkOzmkMfkeZKb6gOGA5oX0SKgxuo9RGs
MLVmxSRKqu7M+fAkSJCiN+DcTHAAFW3mhO0Ygm3SbIUjGtlKUNXsiSbiU9YPvl13KJivrNhNXmGa
bHZ9qZNQ+grntuHYpxxMXOz16I4F6ABCNWvDz9AG1gEjpeSPy//6jpJxM6zp1AMrUjYzNDuoNlfV
Pkt8R5/OBwtPeziUjM6dt2947xXslAHSUv+/eCBmj4ywb98Zt5Vw1E8M9P8SD7j15bJ4LkZrJ9vD
XGw0PrCBLxIZFNYCbRCMw62wJUVcIrz8ibyt8YhUY/2p+ksStOsVbq3EDQLIJR39rPbrKHl4B527
lB/9AnWoDJqWZqUvHOF4l46Jmwo1SMAoK51Dr9uorzWe8nbjxgmjaULrLL7jO+VCNS2k1RmT56sh
a8ZaMhqbMFkHfW5xJ2Mh6XgdZ3LLixm+XpJ8SedKBhR+WhC4PfnAq72vShqgnvKfaSwQo4Rnv8qu
FCIGjuuepxzdbYVNP5ZqL6dWJOrRTw1vg1u2f+wpcYXyG66QHOW/cf6ghzcto80V8Kvvpxd2mVGl
EQmVRm1sFKyuf8TrFBm9lgB9Z5tEkZ3BMrMy6SjdzCczhkge5DgEs7LpsyGGI/QXZg1jD7bKTIK9
S7i+quT3a5EvHhoiITHePLQRuhRAbIe+f86JGBb2DwZRM9Vbyjf8RVAk/KyG169WGHgJqgH1v5Cm
ZTkhIUxuSJijxUlS+JzDabn68Y/Fgs/B9oeHj6TB0q05Qcxrytwl41cvI4ldH36gKJ+YvKUs0LTj
ARHrkur9jjA0MdRlg5YpNzCXsL5ErvUzme0QE+16Eg3vYB7cAsIIfMEVO242vxdxpc2dy+ergRfe
DDdPANkRWKNnV4sKewA45hsARzWlGirOaad+d2ImJQSOWuZVZyRaUeZp/h1psKlmVscblqXTu5wN
3LAoTbBbxtfWQGmTcoUVy/BGWg22sZbg/aMqb7ThK1y1saBGbM8y08vF3mGCoy04Ni9gQrpAVrtu
SlYlAiKgCkaJnyFalfKyozLZg6JCxXzF7hlFbtCmPRFdot4UaeQHV8ufq/dalD5x+R14hkLyfsz2
jakV77ZcnP209IWTY3svhZNkNNUl2WLYI6FomShVCq37Gx5HtLPbzZUxUMboYNjETwzEJxKJRuWR
6cVyhfVW+ja692t8wFQEMFmGVXhFUTVFqlucWyyLQjipgSpP4wR1Q8G/dlu1yFg3QHyzf2vydXzf
w3dMlL/mJlJEvwfMt39K4LQy+He9za1WhYro7ke9/OpfsBvlBVDkGZNqhPKj+wAxR8jlFBWR3xUT
oSXOPOmkspH6luy8pSskLaRESPX/ukxk2dUEv6REFNMfHe6WHr7sKKYjgBrJs3xp3TyJRZd0S3sm
dPwYTRdz2YvY9FaEmiKir64o66/kfieFTb+j4/ImcBYUFyf2E4QP1hNn+2ZKw3U/CDGUl1gUjM37
pJn5ihkrdo9Jw3zvA6FKFr3WF5C9PW94fT8fNvtnbekTgejPPfsTMtqvlh4xR8HLAYbxXYhXhC5i
8aczYD/D5pWM3UWLM+LqkKJruudfkLrAYtGc7OQ2yCG0V5Jd5Y5y3nVozbY0MUtJLivs7L2twn0B
7GHbr8iTvNpM55EHW1IG/xLWHWVetSNfhfmYBMRdi9LQ3Em333x8d7gvaO8cCRzsjoN3+3HzQAey
x33Mqmu5RfFIrYLqENwyR0/cxyeCI7eYMQZ4eWdPULLof/60b6H7wGxw0fTg/cWabW6BIPfV6KJ4
ihSUCIzQUm1GMJ5XLEr3rx+jO+muVYiiaaf3ixE6wp3v0DpmROPo3T5hvxo7Z66E5t1A7Emfqn2h
QzkDybd8gz/wKamyfx4mkXtP0chl7rLK2KZ8Z4fUiDYmXN9QiAka4KDEAsYYO41D1mHGP6XNTOr+
2R12ObtvOwYD7tiO/Waxsr2cXw2PJ5RQddeWdv0P+Yu9qIjuarhAm4bvK0M5RQmaiq275jG6fAYP
pbYT/f1O4h/UsK0MRoqFBVe0k4nVCk7BrmTkJr0J0VEJ65u3vFUNucQJk9ivPlCbjkYVLZ1pGvvw
r3f7h7/rq4uj5VE81aHOonyduNHUoS/Q/McX/M+k+/nXruHG5PHPPiPGNzG+K0FZYr6vGHESldj0
Q/xwYD7ESFDD6y/hCOhwNJx/I0YVQpFygbk4A1C6V0SqBMhI0QyBrvxQojNqMyRtMmibsJ8tUpR0
duQ2TxayxyGaa3s5ZzsngC7eH3SFIzjlE4qxuZgGpSOLiQ6qaGkkr/GRhsztoa+Kfui8TPeZi2ut
0E8Z7EKiT04yP7Q631EuvLq9MurCxB/YGvZ6B7rhdDXwKQZpT1cpya0/bzNecLq4r+Emw9dpMZNV
Cjb+J8CtPpkqlLVj9iUdK/AHceYjYi5zHp3rPJDb/dq0ew0I2APUzwXZyxOvDqFByZdzAlPr5SRQ
kKmTMblJql6Fn3TDyBUa0rRKWB4qIEXl7fv1v2R0qIFqfbhlaDZZadpDf/YloLNVUxsq34ZkcXh1
R8I+tfddXgvLvdND/pjrIe32iy8ClrVMVHBtTi8tutZ/sWcesuRTp0LlET8VDBjkpB8L02RKH+W7
WCi3CZWANUWYZc3G9JIzkQRsyZXLA3v34LyDzAHyup2uBQNi7M8325g6ebkLyGoCABA5jGDJLJ/s
RdthuPD0H/95SrSgrgFqgqFSXCimwCzxr0FD3UuQglKV3oFABHCK4lltB7W3kniH/ARn7AE5NHyZ
IdOolLJogGyqCNm3U+oCb3/jsA0Hscjx9bi1MTrBiEkxD7Z0MHMEmyyNL1XFlQjkssrBy/+R4cze
20uMulAaRRunQMsmmMMZLY/9CuQBxWLsIxJSzNL/v04uiFkXpWgAa7YQtFHoHRrY/zXAJO/Yfo97
PAM2sHOU+YXAjRD5jNPJMefyfMSslpXByYcEKSUcjmfxMEiNJ8gqLG/vzVQBWfPIVA8X9hEm27bE
ZIJEzu42XiorLcRFT4Vj7XiFknQLIdJeYnVsdElOU9NPf4rckC/66F5yzlCp5tPn4UXcrzOgdov7
pzDmFoYcvDEjFYJ2Q2cP4rn7l+tmZ/18ewuNxPGJXxMartJU8BfoDRtIBbBZPYPmCHdHiZ4xTROu
Zd9LBVM5n5EEjqET9WpN4WytYuOipIzNgNMZfBZASPNEyEttolHwuXupR9fqYVNkir1/jM2aK+nL
OMqNSeIWZvkgQOfMYXszhrFXzNaoGCOXXWwI7whbENdbXHJezbNrws+3U7pyLMqv6qRBOMit0o7E
dVwEMYvgQsWCpRwEGMNA0jE3eBEV7uxFLm7bdGVmTG5hiIe44hVAVxhIYhsFYNdTWLA4lVzU6eOZ
U3XHc71WqMEyTTbxKIMqeO1QMqRj70FyKGPt+pZiVNBYKEVdPFG3UapUuPb6+lBBEFw2LzkEYnR9
xQHYRItMQRqjeNLiy80HXyAeaicLmqjzv9c2NLFQ1ixN1egQPn30QQ+r0MUojZpVqnLYMdNs5/F/
ehb7kDab2/DegfeuHlDGyhhBOR38EW4KWV7V3SuGEHnOj04801IcApvvbtHN+8ohV+Rb8QRBib+T
dXz0y69JuTpzEC8Q6nvXmW5DI6gFaDiD4eBXjHgdG0RrQxevql/rqWbADevam3a5m7AxUwGxARqk
ja63v6FSAKfOuHhsGuLlNVIPmvDPKEHlnXBlnNdq/TxlF6JRJhcq9MVp3kRmN7BGsiuZi9Wh2ybE
NELPUnmusLhtKx6RwBeV3T1aI+OKhP3OMj30Ec2Fp2aCEiGMl4i3nbpNCH3L5QjqAFnzCtendGZ2
2CIeFXYVgi0genJt9tr0G3vQWEkHFHqvu0FKauN+KsnHV0PoE1lepkmovHUu6Y6PspyyxIJ8POOi
dHScYhRi0WFo/OmpIj97B/FZGIMBJZiXMvMIosY/bdCajHL9b/GCpL3kCo4FeegBnUf2EhkDFTpC
JnBCIrFdMzyleWdTRaxrqXr2tN/lCL2mz9GwI7DFwCdauvFJF/hVftG2/jfHhIXv4V0VfDnQj/PB
9Bp0zaVG2uxicaKEOz5KNocCNEAKc2X/X2+eorW3TVJ5l0MvBW3PD6KMAQLgNCwlEmqm9JtwYi1w
nU+gwlYXEP1dFO+eUSJM767C+TEtD4HPkDAfUmg2TtLRKA4OOSHBf8Nkdmil3ovOcKbNJ0qTEMzF
ryOwVdWkTth0tj1Z+d5KdLKuglLz8W6FbJZSutTgVq8EWgVy7ZRnWxYsgzvAKzrMKOu5hIngLpD6
I4qW4UfJM3T/qBo46KC/FGa8Mpuh0iGvODTVxvSVh9UfN/7U0pVZTy2J0NSRxp6kHecf8x0LTH+x
sKvSAe28kvfWcgCVFmvFDUWjYufRta4FXnpKOQXt7UL9lsl+sSi6JF0p5yjQRdOstl9l+TfgwRHX
RMT/7o6WfXOJbmMx1QXaOnPVz4OG7uiG+Sz3oJbbWjC6BIH+FX6/ICDtQsKpDrQ0wBN9MxY3XRSM
I6vip+XglSpv/FndbnRt06Gu6aYlYPTeWIzWns3t/bYKoTELvWtqlTvurL3l/zlf99vTdpkOLjsQ
s6MnmfugeSQ/rsW9TUpFoBEif0y1oE7Cs7G+kC7s2JL7Bz41t1tbIOhJBlBKpFJ2XQWTzDBxGri0
QwAQYEcGP0NS8TiLze+k9DEph07Oi7vZwGU0SRtM9ql+HMpk7r6qOpxFFZJXWy4n8JU7AKQPnYlD
osKPu0WlGVuP9xmd6hI6mWi9b/KwIc05j0QmUfBGTOBySF9P/gxdx1UtzXbu8uWhdmumz8SHZRwy
CRtk6o/+J17Nww909MQ6wpTlJ9BwgN6gFtW0CuvDgrHIbWhZ5jV3gYO1b+nS/KyGEU/vjf0a81Dz
eOdoRUdFTdA35iRJhFwLRqbqfLShQJetB6UUR7uEJv+JSvNU797vUKEP9EUKdI/+gkICOhbcGp/O
ggQ49P7844uF5IN+49blwCwhJiS/bSmpRR4sF8OqYBSLuU2Ha/eH9Kf57/2i3XVhNNOzCWdx+63Q
x6Z4TnZ+7BI7eW5hnRMNT7MEOTj+I1tO/x2KPXze0pS3IKUYyI1OFQXAfZwdW1skhNGNJFp22L8F
0eYOG+xkkyD37MzPo5ZREGwtQz64lPZE9Og2hB4BA6YZAregyuESzZMf3sZCtzyzkiWMPlA8ifOo
nDyNRwvd6nFrPRhdn9BuOwbBPgzeV1lvRuUzspaW0zXWmFBxllY9TqSLP/tVTyy17rkdyy9Pz31t
1OKHxMvOII5cnbJvYB3YiftBy8/b7Upg+iWV+C7sV0B+1T1yffHU46J4Tw3OHQqKA4CbzzmDaMX9
INX7PBjPWcdof0+81fUyRSLzT9Y/Oe4Bhup6WgBm/GaidmPOB+oQjZQBsD/7JjCVHxliEd26oH85
bouTZO869SrbN9bG578uBjhlE+oaIUib28PzRIEn/71iHrY8KV1DiA49PYCZAj2wpwXKgfvHYy+U
aM4ppgHMH4FDWdVgDgaWRkl/lF5+MqBLfuWmojchTIsAd+6NWLuCf5vDxmIAXrQAnjFAoSrt/qcU
dj7LGUBW3Jdx+6wc3nFOijWZABVae+QFuJtHMJBzLloNsf9v6/guRerYRJ3sFhlRrZxpPmhR19lM
TxzbvfIyo+wugWmEj9tgNWlvrtAeqoySTEPPStRy7hN+ApvXOguWEmuOye7Sm2v65z0BKGlLxYFs
ohf+9No6RsR7gMrKOozqp41a314uBvlTinQAAY8uVRS1WAVVU71icdBdYQYjhNXiDhdJnSAyzbat
kRZAPgUJo8W+vmL1SNAHsTsBRQ+5j7ziqk6libHE4NPpMUfKU/cA8w2SncP/38pcm4Ne2Fic32xV
Nxvr5RbbXMnpKrwOsGdTYfw/2LjvCyIbE82GfNCsiXQHnC0OAXBhq2exbrOzxOVs31gwFsVN5x0h
cO/eXOEKktlo2eBOBiaLDWtnF+YqGW2nWN3UgONAITRc73b52uv1RZOwVl7qSNeI0NNf+KScozUK
ZzX08fpNzXJvD7faCrb3lkaZcCrL1B9jl5hOeQ65fF4R0W1MOUtMWzFTa+joIvp5/OSa/4tt3Imq
A3DVqoX5CKyMhZ+nyG1DV7k6vYLM4AH9PkZUs0fiooO+dUlpUf9cr2urUSemE1seShY4WFJ4aqQl
R2fL7uE6ErKC1zEyREkWLGlbAzP/FtTW44iqCh18yHVl6R2aZJy6JqJRzEWX3ZAhy7h7BMuCfufk
YSBqbmcAw6EeZlmwXrBBEcPc8sae5oy/CNgQzYsqAEbaU1Yv+6OQBWtLs7ncvv8ycvA8Afrr1P+A
0jQINB1VW7zcEZyMvjACcUyYyXN5zEswo0j1KKQHAtVTRx+I6e+hp8MVrtB2AvM/r+pVhLbumyY5
USEgasF4esmZ3HLGVzpoTQk37+EuaGsqog5mEfxtJKLaGYBVU5vxuJdaTjUx6Zu60udc+sod2Ux3
blvfJ1COeGPCa77E6EphR1aROHwNHlNt46W2fnta5qQdrzeOMudgiTbp9U33Xk/jd8nqaxcx1/1B
fKZnguu1eateY5Mvnnrh0Tvppfvq7WOfJ2DwAUNskuD6R25fDT/TvdeEA/gyzivfxfhLdsWddjC2
ojCyOTHEepyeZ0DYuXDVLVaYsozSGh/2dobEyQ5wwfFAQKAmh8PDcrFu/DKdD8XoI6CbQguiFxuW
ggGfQfRdyO7q/6WeVghlB8GWe3cLjvsEFnzXE5E3mhgkL32cqw4ad3xdAr4LT5e7/me9Wgj4zAfz
CQNvuuruyx9rNZu6nk9uIwlKre7mdH67eiHUzaokXveo6ToINV85cxTgk+o2meaSiTCstAgpLzRx
6jxS5ESCctc+yLYaJMfBN+2FsI3t5RjEaO7FUshKZZsv4SLM/+6l1vqAo1X9pytZR5rT0NYGtgQS
M2bT/LIz7+XAsQKdXSu+5eW33hI+pq8+Qxfs8HmaFi5pN1vmmeREBhGMDT3ybVldTfhy0BRVhAw2
1oeL1MvGzVwTV7n1iDS3Txvd1Rh6VHLiWy7pFW61kSUjJxkeabWyGpulobxS7dyebxsuosDgwjCv
O78+0mOZ/Hcg+htWefWKBVtGFkMTg0OXq46a2Ib8mJAiIsRNShHF5N+on9vkBcNd0OXc8mHeBxo2
dzdpOfiVDJS1+psm5SeNWcoB6yodRZ2gT32hPkE+XJcIX9PDM7hp+stqsdwCHRlH2ZtdVLdpS+/K
ppAcIAh89bmkdcY8gkbQiBWEYl2lQ7Zbk3nXMUli5QtSOEY2EWY6u5UqHiC0v9eimi4FEtNdiN3n
AdRhXFtMujj8wAFJ/eUDKSFrQZWJHvMtU5myYyqxtGwhCW6+o3ZTCZFMZXHk3KeMrNBVNBOYQaN9
CL5iHzf5dVGWJ7qCq7Qg7ARHDimNoIG2aY4elJbn9P8HWGh+jOGJ1NMT/MKYhXN8y663rcmxeJTw
WilgWVjJXCZtoSY1RLoX6UV7h4hPa8cctCvQD/+/c/yS1leyQA5zZ1SEj1dfeh8PVjVrWFaCjz86
dJxgS2e+ztsBKG3npVKihQZaTbz9hSs/rNLXwiEDY/SPEDyz+/wbFeQ4GWXopK35Phida81qKZfn
xPx+1Zd+egohCcpy8PsTyOvPAnK8oSHmkI5+LJmbVNPoOkGr+b5ZVfto9os2/lFO8Edl8hQXwCTM
da4nOradsSM4W/NNsR84MU55EiMRfKAXXHBYRoJSCrTMQWDbsWIY4lDNR8wdinB/nYeD4PWExAKT
zh90wWuOgeWFZ9C1y8qNe6zs7j3X+xdAk7CtLbfKl9agIGw6p/xv5U2oQ/QC6CWui+1gx+cwuzbp
TR8HyXleAB6U5Gax5coAKR+KpNHFN4uvnMKJShtYTUC4djy4Oz52ODC4N2TryiX2rBZ1GHn5VN5j
6LTMaaY766ykcXdp5f/QE3wdfoAy6sGvquzX/Cy1B83uozCzD5u0C8vY7mK8LReXfaIaxTk9QMyK
uFG2Kjwb6Sw73cQXyu4Pc375uH/C0rTcw9S3ChVrEzhVB1zWfQkEU0+9mFaQy+WrxTe3ai91rjaH
p8BYJfpthZfpszgnyc9tz5Yx8CqRJKvCQPjKSYJn0b0cFapPpt2neu/QfN7/D+YmStSHpKYcaknY
8nkFJ6mhrSVOg3M0MBnOVS873M4EjJgZR9liX18pH2KOJ4xasCdcKvVW+HMPDlbeT88MDG8oxvqB
O6adOU2/yJHGmR3g1R3gcxceTymTgzvqtfxeirLN1FZQiqIgJOTQBOy4a/ySyFF82PvMs20Ph4Z1
4zskn/P7hRg5W9+NlMMH/3O1e9JLXuhAPpzd4Mn93URMabak1MFrsmKPxpflp3rSmimHM/koikIX
DawnYKR/MaqhQ+lEptFCmmGWBKUDJB79XbdJ6n6wZwr20RGDt9NE0Y/t5AjPv5kaIiT2HDfT2tny
4ytd0kMXhE/6MwSKlluIS9ZjEPS33W6zVGdf0iHVVqR5jJKyKRpTjeZaydiONOwSa7IXrLSaAFoH
C5xjFhleTFDYOyxztHFcAKgAVwQuFp1hIRg0aUZzQNR/F0HZaat6WlSs8/1zQovE4+MMc2UdzHuG
T+ocUWFuuOwThf5HUA+MmKuY/NdxbDaHjQZOCjJtG3NizolurI/LMEAekkNieVVOK0zSPaY7DX8H
g06SnJAvJ8Kem12yLY+34DLxFwHaer3PmQeVqr2bnOh2W7Fy0m+P07cpI7YsBKhieiovbRKfKI+d
GP0oBgZ+sbDDiZxekK4QdFpNNiUbd0a30oE6rxkB5e5IXcUrPGAffvqHw1Y5XmMGNjc5AtKG1Wvq
tev5tkHqjNUpIqvNZN95nGQzxg86X72k6HhUMuYSPDrpMqmVB+NRi4lSiolzXsCV8fmOd10I5gqr
WR+4dflVp/pu9mMHBqnWNNUdqwJqjNheG8yCsdTSaZrb3312af73J0idVX7GXEjoMPnn+i41ccFD
YAVeRguXk+xtstlwbWbQ5wbcGJREBsHVSjSOyWjFPUwV3VQTJIa3ONM9H7ccl4lLueg7Tfu/Oii7
z4LJzlh5jeYQF7Ajg8OIvR6fgCi00pxNpfj4UGLKpGtJUL5fickY0CIDPjZRYMjgQ2J3QDOXu4Ky
vIGYA39a+iZaKNkAMwQ7ZG+KZX9NkV4S1qb764KpQ5bNUoAxpyyB1S9M1mLJcVMCFGO8caHk6o2x
4OfsaH3iOI4BPWCxsePjqTSMQk+QaV22c3hUeH5NJBDltMOaEzdtvBhsBLfeJrbLkUbnJtL1S2Op
PS+3FA9Qppqqkh9yp0z6eszfjtnaH8m96REQfy1ah6K8gX6+jJekIixzpv8NrFBhnP+Rdy+9CVKx
e0BojO9aeFWBB0ohHVHm4PHbZ4QErXIodeMPkMguYWax293PDS/k9vVU3MLYJqLcgMpRe0hDm1eY
NPq+4yzhiDGhkxYPCd6KlSY2OWJQkjE6plZigWBzvdc+bfFbnI1Q/oHseb4jlGUgGz5ATTA2miyB
jrMlikv93b5MThCnv4llG91pNR2xoIl0Tw69gFrrv9ysl7DFXlWUcwj9/THEfTx+tsJRl+VA0/JC
1+kKXZsukixwxJp9ZfntL+04usVKyKADoEMil/XrzEI60xIMesjuSA5e6WG/r1JY3rnLG/rzWuH2
UaPYTLwUBwTgV83Dzr3KLVfn1KrLQcL04D3yPQe2vhp1wigpfX7ZSoP+dftMPXwips1NzBFLJJx2
azcNZAA2ts5Qomy5zXwKGClThMbXRZO1R6Nne2O+G/upZnyfVV11WDU0JWpNc1g8Kfocbqtqg1pv
xFtDG1Se/13Z07WGto4LonkFYDD5j2z6pc50wHWHS2G6GcEO/LNqCX56UcJQLff06ev3apZZqoD8
g0tgkDt/ZdWgiDy1OdXf4B3EToXQZ+pTa8ObSCQwNdZsDSNAuTa8ylw08p+QHMMBM5h4aKIaph3m
iql0/qSZTZA9RJGuH+npViFQPxH88iiuW+h+VC1aSrHSfzF/Q4+gw7KbyftOEKxuCTxed+2xZSL0
nvGrx/ak5QUhx5yT+ul+7dTvExcVgUjUa5iyH5pK8eKcGbap55mYGvXgfPfrxIMcdsHR9678KS4U
zE2QXiprsLSbbFqUw7h6tyV1yqXTSxoFaQx34L+wMvxMcYbA5a7dz4YlNKS0p6vSUfwi/iRTpPok
sp0KRA0CxI5ysbJrgLdaCkFW7UnnMbBNnWTPX1wjF/dH6ScmqALtf8e4mkv/gJdoezyAHtSSWR68
ieffMCwTSx8HBuTQD1oIvV9Nm2rELQQQLrA51iYTXz3nvv83S/wBdTEi7lSgDvfCmTJyhP178zcS
OjPRvaCoRP2ALeyn3bXZl43ESwNZViTHPAQoPcjLKeSwjUUHFMPFr0JJidCBBueAQsG099MnViSh
UuEfFZqsbJzeDsAPtRMi8CtbzWOse+tniiUeaY/CBuxD+UhZyjo0o+fH1isfzvtkEukciQtOY711
x3f6Vdkqabefkx9vVvAduxeNhi2vuVDil+58V8LtSQRRaMf2N5uQv6ll3AmYUZoDRHmUJisprgr9
wlKfZtc9K0UoJb53/hqSh0uq9NGt+EImg5/mxK+s9hBiDYIkGio9wqS3CaNTFQ7aPFk5N82yHS70
I8VEKWG1VcN0fR/T2KoWcrcqu478j4lcZKbwgrR4dEXCfKG9a0vUtxIHj4NlXgU+zV2iiUBL9Y+k
0MNeXC49OqpwrfVUTt42MIiXtVAZx5q36V/KksqXGOPRiC9PW/4Usl+/JQm0KNHBwNvz0p5powiI
0JKyNTbn7/909U52WMfT9GmlK+jcqTcP8ChlWgXcKaLNO/emoge04W8K9sW2RWMCI900BVayrwqX
VbAt0DW9tWCdgiKxD7o+r8oyV8KEKVzhxfdO/SmlSxtoSRokdrkBjwvIp9pNYOHBh8rRDum/8Jz0
Dw4ApyPy3tjJr0sYlEmAGWMp6a6IeG3kSHYx2gO7+EVMiHV68rGtuCSAuS+l0U8WbiD7AYgZ6EBj
bBoDuQw4J8SWT3S68RSc+9XNHoGpDsk7KPOnZf9i3LRG/WUpIvbo6UuvMqU1jJMPWi1XBbb+xIeg
+cM64e7/VaGQ/xslxhdioeiJdM0Vyd9rikGRU6Bui6W9ujeBOpgE4esJbGSvQV3fMyzecaBuN5Lx
5+tIiFQo7hx6+BwlxlFd7XA4K8NKuHfzLdKqu/E4HdAWQHAmMWdpW7m2jGlkUI36qqKc3mz/cBut
3J8hkmcihGB1wj1dkyb4we0SWQlIm3TKIbvxo4bIXd61pMFXlsBBDubuS+z08pKBD4mtb2SyY7/Y
RRuwCGbcA/vjNSv/Cu5Yv6AwO1FOrjRFR6An2HZGULzMhRrUmRbY5ft+XvR+OqJM2sXFFf81Zs16
9uW1t/yF6hxG5fwmgwzpBUGJKtKJkT0rjgPop73FndZL2aG5R3J+zrjkVSR6VVdMGKplTYNzik3m
Fy83tIIsqKRk8/ntSBm4p5zbsUdm1OR3DfI4t2vTrmiYcQ3r/0aV0Wn8FSDrDWK99Ow2qhKaSIyw
X4FsA4PChe3OHOJEV6Yo5Py6pBLp+t2oHUkXZjRUu02fTRbbhQWCZsi5E0gs5E69Ea6YFMekSTRy
Vz3PwG0DYsoPlc/0Q10w/wU/eK1nsI4rQwqLqkLx4oQtofgDuDZy6Z6/wwISp+A+hurU4qq5XtX3
ed5zmcETakbmKkwYzFZOAvBwOsPipXczTkQCqbnRw0CvNF53+noJA48e+0wQX9h5xX1P6nAhASyn
jotHE4UPlwcQ5CkFHn5saA9I5msLT9heo9vMNP0IJTh85/CiHVyaCt6b05NYnM77ZFGuoxeIZF79
niep9TRCk9YFa+KJ3sI0WzkV6U6em5Y/oeiYxs+8Q4ZiJEtFOfIVyfT0RINFM4wfAwQlQ+JWeTgh
TUjxmNkQgojZFHGr5xTG0ut2urnpFSv3OiWfuQEprQTbp+d/Hdd0anBLC/FnK003oheMlQLkM5+O
06zBsuvtkLJxEdrSHBBNhQLYomauPuk/FmRsdLMbQ9uKqTmnQqzCX8O5Gi842hKra6wwXa3yRpGB
w8nrrOpQMoh1Xo2efgf3XLMLgeBHH2rYfbAyJintuT+6C7nDfWv6bk9Pfgg0XYhgrvkoxXJn4tcT
vC6bO9vaQ4r+DqztOh2bOl8t+NQo1rUzsKn2HKpj/KsQHwaSqP9cBueYUj+yC70fArTgVN949fSa
pOttL4rTBPIZ62RQhQiRnNjThDylDrywzzVjFMwnDVnwMVm5mExFunPaj6haawP5u9C7TLFoAkB3
kPFzxTNp7s/W0TcRbfaA0Bk2iKjjjPEllGr68+afjL+UUdr232xAA0MzeTGDZTARMQzubE5SYBwt
/oH/ltNA7asKXpVyGO+wHYna2JJYW8KRKMkwBhDlqYtcgt88zrZkq0QqbbvkeThSQFzWtG5k/Hx7
bszGuEnlrqd/jSrk3Fg6TT1ykAVyx9+knYdGfB7i1IKkTE0KLYf0dHOI5C2SQknBQ80BV2uOwZQD
Xz8QVSlCBoTG0iH64hSssLwCb/kpHioFAWZMu9npwy2gnLkgtm7VUv1M1RLustRJ28KnyAuL8HAZ
4RGdXLKF1lrfv1PGdz1MSSN+Xg0CYNEbDFFbcT6H/DRryhsJ47zVtziuQjRa9LAAg7o6sl3ATISK
HGM3J0tbyjrX6DHFGziqI+gyC+QnG8aZM/rUTHMt6EvvtxveQD11pRkHzeCn+yi5hbd4OZs7h/5y
2T1IUZBwUXyCBs79OhMmwBSVLyAWKOQIGQV2kcFIf9AKqX8pNyDYR2ZwqhN1euu3SyFZCxZoopPq
nx+F9BbrU5xLoTxJE09ZtBnsT/r/uGqE6meSC7GMmI9Sj8f4dSEBY5dIyOOoE8N3FDG8tHFy6OhS
NE5TpP9LGzrvqH5E1nii2m4UmvHA8t33d4228lRCUamOZlY+HJPVpmyq4/yILxAwUePV7x0Vb4CX
OktuyaBTGLg8QIqt+VU+ZsOaxOqQLV75UMQJweD2PsfoUipvIepGcy84etTNP30Lyf2cJ8CetFY9
wblb3F0V9nVtpJnQrwFLL1JI6HPPSVSGDG7HUTkxrVW8VUt4myklmWK1EL0QRwn0gvCEBDjAb7X3
ivmrxU8pRm1JQGu/Y/cCoOaT+YfA2KJMt88RDm/3O/snoGNZjyQQ78e/BgAA12VzK2bVcpC64S0F
xYp0YrEYLmrnPsfRpBYTi3dzGDdM4jFri5PW9C+xa2jKPtpUxjFFbLrlVQsLhqzXG3ycnAHR1BDh
qTVIs3T3fMF+lcQTL0US1zFpreJ2TWNYj3fbVLUgdHwZHSY9iJVJRK6j+MGKpCSU0Om1VAb3/s3o
pvJ4RSrWwojXrvnn4Me7imxaTNFRAggxbr8lTFl+t0uITyFRTI4En7U9/PPbjSWLRUYLAKKSPgxs
7XHwckyawUhYksVFhGpsm94EUZ9OuEyk26eKK21l6CO7N0xMLwVLl0lFLd1IxKn+YbkG0mJF0TyC
JJrfSYA3/Y2xHATtnV9DlmKHKcnATivxXmlkh2zO8JZD7i2PPBumujuFrSs7qnVwqPP2Em+ufMT4
LAmw2Gn/qmBcNVoDdwyK58pGkI7qNtuP26Rh4bXXpuHA27EEyWtxKjNfo7S5owoUrlNXvKxkOZot
LifsMismn46+0/yr34yYRQtWY4t4YEnmikZo56p7BFU4Tk4ANiuiZQPhm3nzn8wBP14DJy0W/qKP
MvOKb6wQWmYs1JS7BUfMA4iEDARi2iroVPusPV5tvnb5zZLFKfgBAlDdEzrgUruwHolTqTnAIk7s
pQ3WQ5gKw0OFbBYgcEMEzqpMM9LhQY+nTd56ylZoHUQbF0S3UlL0nI6XaWVTT+ey6JyEViNl4aCk
C5ZCPIv3SuN1EHs/MFtgnmL0xcjUvBzWy6zc4uzUPNirXJGUyC3NtaQWbBv+s3WFGmwub5cN/1aI
XN33JS1o9NnQTP17gzxFclOfXRBf96Hz2xtCMNaG0hHrR8c4RxmlCtZ/39HJMnFRGPfMuLhFyj/F
AjQfCgbXs02o8kd5NxN0Zxxy1/2MWCZx7CCwQHncmdD7FTn7fMRaAx5l3gVnhO68qyBOhXKWoM2f
losAUIJs86iOL/1t1wQrTcHhC2FxGGBW11ZKF2PN+ZqTvT+p53q08vHTnDtY0bOw+jOi0fNt5rk1
/duobND7TFSoixryt338IBA0zBoaVbIfgmGmM4emuw9hRJLL3XBjjFN/1h9ZGe+iF7fwWKIGAvPz
GY5utim032Yhg0OSbL0myd4MQD9i+Fn3Eo07pw/kDWz8XShNOYuOD1NPg0E23hlTMJuGexLcWSZn
Z5rndGPB5lWPAjIQ0JG6SJPqlWk9MlrF6CncoSye6Tki4DXSdsaGNMyt3sLE0orU4a3p1avrUQje
dWcKWByf01MC3N1HZEKaRDD419Ar7zoG/r6Yy22J9Hu/lQ3atQ+qtw27yq+m9Siifz+7V7jw/Cvt
KyQ7sjIcBzW0Knk/VTDBL0t4zVqGQKFInr+4WuyxF2kcwW8bftM1yiTUHevzMpkXvzth2T0bN0G8
fGeYmZn3B/O4IeTdt6JxRELNzpVzxCVAHm/u4yE9radYvIO1CcM3pwC/V+PO71mbumGM9/PLmA7h
fRA6X0oqdNDO27Ly//b9JS6J97X0ERCNqa2q5Zc8vlN+CPH5l2oCbElwlCzOjEpLI3xk7f//Tnde
b+tYnIf/zpUrxSHqwZIXhGTxh/oPAafWQJiRi+SJfy3Gmt0U9JbM7IvbZuJgCT9NTIWip/hnvfnG
NUS8wpLSp654NZrCDkNI76lmPeOzmn7BNWeUZweRm+utV68jtfaYZe6jKMHszY/VR6jiLhPoD3RX
OMoRNybK0UQ4BweFqL3RQKsJgA4x6dypuxBuciQaigI5gYtUizGf6AdSFlWYVLnUVkmg/3UOu0+q
X8198ntsfgNwcehz9ebNAGBKa3ZWGUbPR21v4vVIAdN00D90NxFGfv1doo0kfEgHOjFVj07N+56E
GsPLcMYxjcLp6ZJnyQulCjXEPJjf1z6dmnky0nTD6mRbowJ2FEtq7+Ggj0zGdMwQv8UUjN5NWndk
yvMZ69j9/3bs76UMalWdPPK4swaTk72TrQG26NnoW/mjjuz+9oWI/cZpYoYjRvTUTjOIVUqws18t
omUwB7kkiWVJsLZH4fXwpq3GafZA242l+e+3rBee1zx4j9KiLWUIRK5ZQN9+ZwpQPx5vuS0Fpf6Z
wtxx2FaZB+hbbxzIIScylpW2fDCigRUUDroGetVisqEHJeh/3TGwNsyMcx8cgeYkL1fqGWnXQ90L
R0JxXb1VKZr8IO/L3jDO3Dq+6FRVQay3AjzxZIPCoEY5yzweapJqnN5qC4p5oCUBYHzqRqD03Gkp
uTs37xJcePcz5bcM4440UXYzhoOjFf29voPhyJ1EHayhRYIddLqpfX+1/GlNZge+f8nA66NXmKxD
TtXj1T3LcTq6Ne/ts6kG0sJ6OK1+CHXjKoAjRdrBUZN6WEdW/AxnU7axRcqGmlX5gfglIbO4epze
YSwLZPHMQqfunZ2C4XtcoDB6NFj6Dwp0MNU/kXQ9YRBm7mSaQWZu+I/nL0e2WQVJ3Lc85Lonzo21
cxRdFXLDpAEgYkrp4M3M34Bf0BCb+IiPKmoXQ9mF6nYC2jutpishltpenqIleZmp3fQR4ajL2kxE
p6M2CT/1440/O0QQsf0ouahJF8HRWT+zWCrawKxZ7aNrSBZjiaX3855iPl237Elnfk96RADypJi0
9c68WR1M9mc7nVoY12aGslJwAf0021bn6Ykv+StNs/HBHe2yN+Cb8JmTm90nEwGK233PzU5j1NOV
Pi3epX8JAp/AsrVMzaMXd4sjBqf4QFCdJVE3OWqZ9sNmH9Sdzb4jX+Ebpt013X8K/0Wyaz0eZcvD
tvDkpNwLG6C/ABNrf0EjiBWAYu5+ZiErYoNgyw5azxbufep9N3Bfa2h38gevpdor7yBqxLhyneH6
fOoRFw+FWMKAbJI+mU1/eTiEQG5BTMPtDj3FwhTzuEV70TXjgdwilHrvMZfWEv0ZIYDZi2GWO2To
lcmBwy7WtPwwcA6n5Uj4bvKCINSbBgqZiBPrRsUOIj97hkyZS301oa6Jq7e9GHwoP6978tpiiSwJ
tOWLn/bi1hN2/4zhsjodg0PdP5wXFwK3l4N2PcOKQVH0buZiQAlCx+zWy9HiFL9CnbwYJXYx9rIG
6KHx1aTEIVfYThA7mFiZ/kw+9DyhrKjN8rs3CkbvlCLR5eVdJ3uM1+Q2TGDpT085hDmARFlHgx1w
dA0G+P6z1hKOvSZEn52TdH9vK0nczzzTPbm4KEXz10Ia6v7VdltuUDtEEGlPoaVcRJsuOOmEeSwp
QJ/2SmiNW8BWjNumEARISJIm5tNgM9Y5pJkK0y/1L52K6TeSr7im0Rag3aJ5Nn0hPQIrFNgIiD86
DNK/j0X0Z+AriQ67G4VE9RzjcjDo83r4O9rV5sPU4lom5/erzIlj/J7nB5ifTLIk7llk4FXtjqIc
RCAZFbrbYYJsfX76p4BBao85qXU9j2Tzq+NNXNn6tNOSswk1RO6CRZANLwDs6qEA4IS7gieQv28c
F/5B+I5SX4eu7YeFCD/A9cEIvdMZuYnDv/yTsvBGDVlAn8BCtSCDp2qop0ljPbRcUrH82e2tlWz3
xWrlNXklVfMqh9sKDMUAUwvGF5gxf0doMS49QwSGI+JyxAxMpAoK8zwGXvT4elMXrpSnnNmJx0LP
ninszRmmoRk3euPPXA+vJTCQpoihBxFxHYKd0hr50qhqffrOxwlxLChGpPQPrQ2Ex0YsK0dJA+s8
jd8rxUbotfw/8kaBVHsXmrnGt6mAOA6KAliOudesb2fb40hveWW9mkUUhP9omCH4iCQzqNrWoX6L
JiwavjeGnq6H/v5FtzFJXJUyZQvTRy5zIYPTze14zpU8NLL9LYpX96X2UQusUm2FeDfNmFRBQWnE
cqyT+K3OIxAop3lJqiRkfqdaEaMYZY/mqI1KWAu6gz+8sA8ZNPi+zEbzxTrPqCct/KmWUzjzNBZv
HwteuYZY5iiVIFrO7ugQHC0luKPsJrEjvJvfUsDYdQn9+80jGz7MNy2H6IjUaexB8MwpSJEyF7aV
UEzXk9lvZilZ0dHqJYZckZ1Zq9LB+4P1BnxgFkucBusYehG5xr4PlFXjWZJsMF1NfooslqUN8KZE
haZfUEbg5keNufpKYfdjKEtjhVvuxEyrsCiyV1p2yq5EBeoYlDmtuzLJSSPIunYIjZArNMXynp/Y
vimLWiBQl7H/F858u0eVc2iS0lVwDJN8qLI9FLTQpgzuih0pwWvCcRpscmpQuDuKN/TVLfQqkI4/
3Y0UbCckHzLy2xEBpT3RT0DprJhcmiN7tQFXugdZH6mV+mdRHwSVyVhObVZykSrNKTzvcJVzgMzd
ZA0RR4oNojdbX9Xb8wvwyWEw5yZQgL8zBx9OOnPRXLX35JeuXJHGFtYanZZEb0NtueZTgV4xXeCa
OFVHAJUwCz1cLjVw5CkCv8AHMsFeLtpG7CFKxIZxf1uGBg+FnFOo8oWETOu7yehRzu2CPaIE542T
SwkKpak9ulHXceBxZRiIVnUBHLTRjV2TUWvIsBpECIc8EcomLF5StnJN1vQwaURqnsUwSw2otdX5
Ck6uDVKvSn1ieTS053ZwQefhPc+aJ9kZeVabGKTi2DStKAR8/L+ral/pHWToVAnQj24SGx8ex1Yy
zVx5ZSdcf5i+1Sqqy5XNk+hjTzjzaeoOGKmCxvUg0+gJHy3XO33F5oJjoJLtXm2VA+f5p2zO6Cb9
YL0i6XJzTvRtP/GuNnu5nTJBNYauFIcby1ifW1ZkOqWFCUswC/BpiiJNrYw4zAQ/7zo1OE+SiZ9x
vUgKbaMGTLtky5ETEigWWHfsOGM9TxFlSbFmtvINtRtyjymQk+YFC2aCbuuqnak18sDChhFwnmKX
TjQPPrMex5V8fQSfN//NI7RrabS0OT9N34/1gutUtLlKuA0okow6s2A8Op+oWoSdCfA1pUG3efzM
UTiimnoBMd4O6NHcNs5aWr4rSv/ASUP+3KFaNFlLRt6045lzzshqeQAAPy9qDoAmrXtKPRlYY4JY
0niYwxqIFf3kAxa2B/bJbHufXjWfJ5YIR4VecWi93ZHs6f79mUNLcV/SKR+Ib/yd2hOW81BVt10G
G6VvvpiMnwsRjv/oW46rP6wF4bFAutZdyIe73jbfM6/t+8/y7HlA7F6Dq0gpznLZUlkNXxMu9igi
fUQiSSNB0o+iPI/RsLlwL9py7ray7Xidh3/daX0GiJqW88WfB0yTH2HDaAIxeuFMuf/jeIhphOuW
R6sS8pbshNe5N6BZZfi2VQuwij0N6UjeFiN64VT1Y1fUnRTAaVlHK7LiuQqSd8J27MZjUEDI3CeZ
4w3ly//dm3P5sKhBJs5Pe7jDWfHG1YVVCcre4Uje9eo6TkAUE/WRLUk90B/8AnxNbKQz6W7Cp2ee
akrTBuJfGhob4M8QN90ruZp/rp05UijulogljMpdIbDRV0jjey6nT3lh/IFSffjQ8tsqB3NhEu+2
SxjdYtJuJ3fz/WjBQyym1rt5FE1x0idJpso88ceqaee3dXAhDG0mStGW/tqTQvuwK+P0DtvkI5be
/lBhTRjH7lDVD5yqQ0QIhKFNpq7TJwb+0Ocrnz356HotJsbIzncZAevdlID2K1qSnZSBtEtE1yCP
S1Y4VRwKWf1GhUmKZO668RtHmnytFDbjv1TEq7YrDkvDIDONjnPmV5bzw5EE91nRzSudRjLth8Wg
eIxJkcmUnpwb6urm6f3R+5HEG8WEKYDKryExAEASjzYicRgwNCpqGvkXlRw19ojVdxbDyDgQc+Q5
yeX07uOGSUHN5WFvH0jv0LaB5KDjkEmArt53nUCZM2MHLebcRP74FwUUvR0Uht0FsX5x+e2yM7LS
RtLgTbCfeBRWhnEAyt2mOH4iQSxZcnacoZtcUgYbVCYlIEjlJFECyIS6yvDp8YPRWMxdycg6iHjE
sJI56tIiNo8hQUpw/5dOgkykcHuXXgshxWhgjMwvH8u7zCHsZE7nALBYuP0Q//niDuj3Ni0GHNc3
EMaiBcCIYeLjE2kzLq3fRh3y0Tvw4H53gKihmScNKl1GygtApnXrGRkkZLVhtNFoYhDH+AwclJvH
3tZDW9MLrgPXh7cZ1k0JNCHMsR2CNvWJ/fYrsA4X/LbpsgFVlXDFyj+P1reZI4eEATOuacVvo6n0
6ErVbx+mXcCEx16TaSVJLxN3k1PdIlD3+P/XPnYBDHKxDqg3uqkfswO3CNlMOrZ1d+/fxpa10G8y
WFgjc53xwsZs0PDPXxJqikug2OxvCPYjhIFFD+W9UOfJbZfA1H7LjbYnW4Q6WqTfjInyBSlSHwoy
hepjV7kpGBz92dOxj0p9aZCjuGVRJbr/5c/+LUD18sNOcMaHsH0zkH8W/Ffnc8LATZBUHShi23jp
z9j0uqa9hINLzLx4Dpx78mG5zGqwVZi2d+W+X1w+YC0lGfoB8tWisS4hIphrvtQfdiO/+vR58Sh4
xyQtHyNKXPVPeK3xYfnXuDX+E5/LFqoRoxywX1pZoH1WlTCJ7PUAvTytcG2CGJAbzrHoq0rFpGOT
gVZTQE5AvP7OPW38BJueXOktpd/2pIqZsjLqXmQxKD3g9B00h1RT5y7z5Oa2fuVLxbLD55HGpIqH
q6tUIko3nw9slFKsLJN/GImVHer4CdSPvpPKXaSPRDiCrpnl0YRdvRPjqBl6LqVRAjavePJ/fhC6
r4+0OF7StWiHIj1mBKaJf1VnuanslBp0rSrOyMhPWuZKR4YfeMmZVVGWK6ssoP+yEF6Vd971I93d
19/8rYmolD0AMZoV+Vykjt883Uz/32BPTmQwsQu7Y3XJdXQ8/ppWXK/AvHF/G16lNBTV/ujywXAD
7eXea358l4zIYRTYikHETkaZyvgZTQHxwBW0yo//20dyZIQApKXKREUINcaN2TzoYsA/vo0CU6iy
URbap3g6c4rXOEk9XxxO92f+hlaFo06syrDa0iydRrNRgBqkELzmz84PMKb9EGjy0oYu2Rh7TMFR
w1ul+Jx8P9v6K2X/DATicAameHk3fuV3UG66jwZuqvJGwwiK/7ZUyGtvO93/Coib9LxQu441WzXX
TPr1vaQO65u+wlePCq82nDVL0pkCGDiwV1w4p++gtOMw5m1vj6Kb/Bc5zcrY+3Hz3rfbs59ekKnE
9GByFYUToUxEF1kGN7sB/iRFoL1p5EJSe91GR/PUkTeEq375914P3+G5mrZ2Q40NHFkDnBSt+sh6
iheAYxHqI05gJHRoRrosmq6cV8aoWFkzuElnZmHIN/VCka0gLZVKZHZWDPB7iOyVKG06HATGPUEY
PRH7+Db3M0o6fwMkGEhzi9xYAUFMWCET8lzGJWpX8ayoMD7YItjBLSyj6rjCMyAOuzI1yuRBaHqE
KUbdGd7iBE18VrCluIhcx9qcfKqf0d7IdmSvoSVmLh0CNj6knWq2oYEyDlABL6nrrg0zppzl7R62
GSd/zZNYK+KXogOFAkoZxc4+dlSufZAq3BipkSW+xsrLjJcRKkuvRzAhDCvmISv2vedMZrFA8pFR
HcCPFOcZl4d8AaEvpqpZO01s/19hGAU6ZfEaWj0cFokNGxohbEZL2b757BMzpgK3LrPlOlx66VvJ
cuBx5uAKQiZmCtm1uJR6TCPqf5C2MIaG1A5GWD3m26P68JZkDzu6QyEnPd/qWS9HibtxRGVG0m/6
F+Cn7kNRf0lVohptL3K8dH5hG+2/GRuoYz8ZjdfeEyJ4sARaKjDDdgSvraGltF8onfFVtSK9G4Ci
mPX+BKM5U4b0SpHKdl5GQRmIf/iE18CDmEjBwuJsd+tzsWNUz+m+egQ71/Q2azQY/DdmDZ9ZgHSc
g+176KPnvBC8fomFbSiYrOKycARrTQS4uQcN64v+5Y+sx9CqoEh1tWTRecYSkmNL3NFEqxp9Zt5s
qaL4nrdmqZmwSCTRF1BNgoNXY7/WDqeH2XolpflWaOsd0pJMJpKuNCnxCC3H3XQuEcY6P7nqkb4m
RPaqmj03gVOCSElMLyg+libi/sgcYWVRBj+pRPuNBf7jH1i82a7JT7gLAN1Lq1A0nwUW8KXJoLl/
0Sm+/AVahmUzRWEEhPf/sAp1t3qoo5momwcZqixoTBbCivri52ZKuC2344qukiLYbZNXpZGBaoqC
6Vb9NnRCPql4WzfzJNcEzL8652GsJYr7dykn8O9h8TSQrppcyQnVy+oO8vUWX/Sb3TX8rpZDcIAs
+2oI0yKgpmY3vU2nePPR2Wl2QHRJhkXjq1mqetOljtuV5k49TMyy/sjUEWoe+Ol95xysts7itBVC
yMopHXqfo07yc3X3n/KzQF1qIIKfT3h+XfRvhonBf0cv4a7+E/bJmK0YqFwS0792xmAqYRrCE3jB
w3dbUzGYfwTDB6mrEhP46tiTC5sAHKsOKdXkYi3s5iuEzZucF1PYNy8iaFgIdo2ajxBhAd9ynV2p
5dmm5i9Vweli6mce/TjJlqTdxIzpBgWpnwHleHHwTeqUzbE+YqcV5VZCvgRfdSlNCvPVFKPpXzUP
jjg1QSh7nzcSDFEg41YWj0jP55pFbyXVkawNbY7z+8c6TPlwwA3AQuDIj8haNEGcATeV17mW+8rl
eLLoLhaNZ5G0s/tlof/JZMkhaZc0G71mtvzt4LwCEPkCkXyIDqJWuJqQvuHS3yG5mXSHprLx+fXO
4pyRVPYseCt1zrWtJ2uvtn05tpRU4r7BpL+cvntv9V8IndinNeSF/S2n56bListUmf6DSh6NMaS7
J+uNBn0yS7K8EK7XVO87s6x5PMB3/x5J/r57f8HwIH1Tt7zhn+IXjT1buu16EUGqTQQvTrI3YZkR
u1e3P4uJRVg3Sg/HOp6Q1vgXV48t+8MCZZy+1YPn/vsc4Ehgrg39yzxwCD++2iN/WU89uPUCEA01
YGfYa+KXjJ+eKG/cc2kuWgP1jq70QfEIqyb7B3MzPaFLxQ4ouOxi9mz/4bFYXzokI96v3DKJ0lu4
E2kny77Qpb1YfC79wWy/fu2tL8AGWY3ba2kRmkdJcYf2H+JbaCpJfzX2Fy3cDfFrkCHmTgg9FFzY
HTZ3Wmr2vskCtMpAWlEjZMXlE2KSzdkRRki/VlL5ZoeU5MOo+fz9dNWdrIxqu00tUS9P0NFHPtva
xdSA7uuj1eW21wWCAGANfDJhZFC2XzVV1KzCUixncrLZhMf6Qj3gs9hQ+Jm1D3hydv4vop05IoUi
ZZmNS642QBf/yxJloCQfoukn2WBrUfwmc4o5J+RVRowylIu78Nuaz4L8RI/aljxo0kvApSLrK96U
zk8yB/UPWIpJKHDxvz5x7utizlz6jWU7ZHZbAsNG4JejEWtBkIAukIYk8ARQAydx6SIBSKTz5uid
F49azPHvHItP7C9VMY2ed0hQpZkkiTyaDs2LL9CK64BRdTeNbOLkOe3veR0KI55sbOUnlIWPSU4V
KoCBvl35OBABf+aFvSrF1K4yAmnIB2tYOosVlf7QWRUkLTN9CtcucVIOqKGdK79xypS4ybB5sfIZ
v9Sl75HEOAa0KmVYOKHyNFWeSfp5vFZtR9kOpWglu0mbbmNIn52TtOxHpINuFftz39qFChPNFy/H
HI50G3GmrR7MkNxxJJ7gYqAInzUKl38vcIHYmtmrGlDJ6iXt7GHevUrhvbE84Uzbk1Bj0qH3Fqcp
vW+py3BUV3pgGcQjs241b8vdHUnBw+GRMdIqIBdojLZUnFu7zAojgd4GGF7T2lKGxBg75YCr0jFy
xffG/2vI9D5I9OCBYHhoBwz+uoWORsiADl8PcM7ulPuJZy1mow8aVxejnVtubaOGUZryUI/cO9PH
Rj4uW+nzYbbadM44o7uelwUEdJsoYTcmd9p5DmNE9qYhXsPxUnkWkDtGFNfdgLyVFmWcqkV4bbEE
8lxRwhPfHGasD1SgSMGAjZaYwZ5hwoFwyir8ACW5ImvpDbbvC4KInnP17VvZq1W5099CBaofXYf9
FBHmbQjM537/Xq3YhBRKG5Hk8bkT0xRMGY9toFxcydYUG4i/nRHHjUDrzVFU5Rmf1nb2CfWr7+yw
HPziwvb7eZv63b7rUPn7lYBq9yVTRaNS2ihDe/wijQlJPt6dKAgAng+GNPrsfs0+r2gOWcSLLC9I
XHL8ZnkhFDMvrnRr1IMsTQKvnp0Z01MPpM6+4sLyKI3pKT1EwH4WWxh6GGYOTiANvdAh1KIC3jF0
7P7qOQtHkvNmb8M9TniajQ5fLy4XEDFWaehbIL17ZayOGNMkltMovLbrmoqJ0VQ3TNFYe9QUUNfL
O/pZQfPfodThYWXMwpdd5vElH+donJ/UMCCbt2NiW5Ga31N98kCR1XMO03I1d63xSM/XyQx6Ei9/
jdrcPZ3JJSyIbE2gn5vGBX7R0vilUkm/Tp9IdWHqMPX9vXwvrgwI4DRpntUyCnk2Mnn16NKAZkZ6
OTUmAz5ttV4RNNmxanPDRcXkFVL+af/PcH4RAtJs9X/Fl+nuoJNA4cnsWFiWIdQKVfqhTJeBWnRy
1NQHOTHQYt2aiSvRy+l10JgpHxLBkaH6tI+NIsiw+95FYmJfzugD43R274vQKvZzaVSn1AujG1Ud
nz9kRWXu3hp9tBOL+OGupuFnBAOPdcKQIBUhA+VinPDfTcJufQdO9UrgZSfjyeEvwAoyODSFB3Ea
SAauN7ySSDtw9XUubaRxoJQqSm5TzZ0F3Bjan9YDWpBPsejlaNNCsumWBONIopd5ygkN4EA6jmSH
ZX3N0a7F
`protect end_protected
