��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�	��g���cN܄w�t+�!/� 9F�B��X�ī�_	O�p�S�/��Vfπ���&WX���_��*^�MA9�����s��\����:� o�9Wz_J�������q'fҁ6��,v�ԃ7CVs��֨D �!i��9ŦU����jz�Ye7.����g_H�0��y��?��[�`�1����i9 7a�Q �8WY���5�D�nȬf���PZ��_Bn����IW�����
��y��O��3vF���K��wdKȮ��f{(�	xp��\B|۔#3g"Q�z?Yc9��~���:D_�{B��k�x�� �����"k$�f�rԾ`�R��C��p��A���02p,��B�����_�f#<�+WA��s�eI4�G�����溣�I�{}�v;�;�u��S�=�U�1���`۾�`���I̊������s[�G���S��e�I�*�v�KK��ro�48N�냄u�N���)��$��� x��Ju��0��;���uC��J�^�̲C���6�1Z~֓���3��L�ۤD?-��_JqEH��?�[��-ʰ����V"x���N��{iv���u��]ܮ�J�����Sf���Ů�1=�p�Νk{��	�am��<b�%]��Pk�9�#��e�� R�)=P��Ⲙ٦�Ģ��7n[&�Qa-��O������*Z�2�Y.+�=��	1y	Lâ����끦+<�Q�7�d����Rm"�����oi0�t���ޓ��8j���Yz��Ap��m�j��y��u<�)%9s�M�ܙH(�Gr�"=�����wGO;B�= ��b��]�z�މ#�Xy��?*�	X�����$�m��6nė܌d��0�,B������:��d�U�h+�6E�4��Y��ϊ�7�<6q�f~dܒ�u�X�G�p�j���+����K�������\�WAl6��g���k��\���
��"��){J��8ب-� �X/yO�Cޔ�����G�DC��L��	�l�K�#�q���h�D�����/RaD��j���t���W���wq�����1���g�qP
f&��ژ�-p��~O䭮��N��B_�փ�BX�¨P���&lP?����B.��p0Q�����v�׵���c�۽<Y:5���Q����� ���{0�|�f"��D�p��9��$���J@�}�.�����P*z�;�|��~=�`t���u{�����(ݞ��d�r�tG�1��#0c�]ܻ.I����*�)OГ(��m����[��kAL��{8�L���i���Xc�3s�����p++�m@O�B,�_H<��9�2�'y#sz��IW�S��z��jZ����̻yZ�^���3��y����;4�7ipb��o�L���w�g�.��ז`����?b�L?�XH��n�`3X= ��x�p�誆��SjƷ��y��:��s����5�M����e^�%i&�_{3�d�Q\S�׫)7�����\�g��a�Bu'���:ESUQ�Î�	��J��.z���H����b̓nee� ���z��8�#�q�4��qi�O5�dB<�Y�޹v�����g��c/��4&�xL�ut~A��`<e��y{o�ݳ���,P�,�OY���Qڄ�eǈC��T�:,F4Xd�Pvc�I�a��a��M��ג�Xp(��χ�r����	a{��������.���Z����*5��O{B<���2�!��._j|;��r�b;|
�Fc�'�1g�렴��jUu_`�����R�6��lk��K3���#:εׂ�,��r�*y��	���i�,'$�B�F��V���s�A���>��#�AՈ����8��6�qmmf�g��B�4�9j�{�Y��a_wHZ���l'|�e���r!����4�jʖ�ae>+���Р5��|=5R�����CӼ�=L���Ms���2\���O
e�6�k�?F��bl����}bE���G�����d5�BD�梛�,�E���1��q_���|�k�����#��Du5v0�,o*p�d�F1I�n�o��O>l�t�bo	�xX-�4/�zm���m0�uq/u�2��<�0���v+�Ձ���f�,]8uf�x��U�a�\-B�"C�a
��0;�,�n=�P�t����<��_��?n�u�����N���f��~XC�����j��Ӵ��5c��.��i���% \��Բ�-�ă�������S1���7 ���&+���9E�e���#�.�V��8[��m�#/&+;��[1g�K�����U��9��)��FN�Eۻl��Wa�%�������Ȝ��U�Us��U�ˬ|Gm��4$Q-8dJ��ι�S���9��,L�,�\e����T���pX����%�}����
�K�C�5,�����ө#V+k�Ǚ�	LO�C[H��������8j�4�o��P�1�|��B$�^|ׄ�ꎙ^����K��ĝl,�,s��O��q�pլX�7r��C����b�x��<9�O���@�
�??Ϡ'i:դ7����B�<�;I3s-l��)�>�Aō��q����(ϳc_C�;IoÍ������m��N��[�D�%�Q�DѼ��	�;��t8o�͘�É�����&� ﳉn��ѳ@\�T���"<se����b��.�g���C�^Ŭ(fB�ȥ�
������7��g���";�{B���{��p���P}�e��tYV�Z��y4�9"	���!�@�&�a�H��!n�6=���ǚ㘚����I�8qE�΁�/���Y��4��gW�J��&&vnR�7�L;AӏZ���ݑ�6V�D۫� ��}�F�Wp�}�O.�8k�\m ���trJ���k�������Zc�~8�= *+�URC߄���ټY��No������T�;�ԙ���0i� E���:�?�~�p����#�µ��X�˒���|�S!�� G��@�Q�Y�'�^T�j?R�:�o��&���z�����im>�#z|��� B��� e�pi�.�Y蕜�����Ƨ�YΡ����}4�K�U�Z5�g��+T5��v��*
>2�f���f�),�ʡ�0_i������xf�R��
ղV�؝E�S�F�����k��� �OvI�l�(P�Kjýå	�I�/��5���z��EG�)?,�˿h�<{#�݃��@�?)�[=�Y {�����Z��ėS%�ˍ��v��-��@p��J��Z [���D������t+JĢs,�u������:|�؞��+)�F+�,v���XS�I�-�s4��&�
�8@Rb��!]���lG,��w �`�q^�y���Տ��:	�gd�6���ZB���n>�;�ñ�<G�r�N^���YEn��h�vjD`�
�3����g2�e���֘�ں�4p��?)ܨz]2|Ȝ1#d�U�/i!�#˅fVp/H�v#�|.��lD�1D-����b�|)}�KU�on�6�`����������J)�5����V���&�iD>k��ӑq��EȻ������c������xW�s�4g �;G�2�� 2O�M���C�4/�����Y�/I�B�Ds�5߾���#��`8�5�b�M�Kl&��xoLt���Yy��<4Q`[�M����.,;%"�d�A?��J�Cb���!�Q\u�V&'�FVq���Fd:�!_�1��<�[�r!��o%*�L���ҳu?�����0�6"O���٧vjMf������s�k�4�]K���4�;8�lb��e54�N k`؇ʟ�X�I��-[�Ȩ/O�IB�p��W����b큾���O�^.���[��zIo��]\���c%�/e�����d7.]<L	����{��w�L�(lA�`��p2�b}t��`A`rWy������|I��GT�!�gTe�7Z�!�u/��s� ΐ��sa�Kʊ������:�X
����		�|��`6�%f�'d�Y9��q0����@��8��0�T͞�k��r�
5�@m56�����]��9��5�r��(]�����6�Y�JrE
z�9��_
�｣[V��1J������I�;�!j8��J������zκ�'�_/_���#�;����׹��-�����������C
8�"#��0���	���������-\��tL4�s�.}�VJ����=+i �qG��=�J����xӘ�j޲���æ%�u���0�ϓ{'__w�?*�n��!+&&�5��#7�Y��ǵx�?��>C��'J�U�WX�"���aQ�PI)�<�Ɂ��D0��V�^I�R����`M^��L1�s"�Sm��U�[��3��(�[��9,�bֹ�"�Ÿ�c��{�߶9�D �_Y�E�~�Ŗ��-O� �vd��]����=�kxu'��n�YI���ӗ�Y��]��T����X�}��̪k d����_<+y8=fC�2�y�ֶ���bb��|��.�4L�����|�!�S�&��
�n5?ʶ1^��TJr�X����&��%Ya����ʧo�8i���E��D�i���mOgJf�*r��X�o.�ʡV��{�+_3��*��薑�ǁt���4�,o���q���3	p�-�<�c��K(�zF�5OA�A��ɦڲ�_��+�f@��Ԟ���_���8ܣ�'���W�F(܏��v�)���9�ť����l7�S�����Hi������ �?��bgm.<[��0^�Fb7�^�sM�aw�5Y��jlİE����ʮp%��*D0:� �D�j����m�'��Y��G��/���NN�`z\���t�*�򥡍Y!�"���꺇;�h�yB�LoZW$�9��&Riz�oΣ1]P.[�@��_�k��j�������AjY
��pg���b�ڡ/\)Cn�*{=g[O���C�w��U�`�}�.s�0L� �ײ"5)��Ї|O�Y��5-#�����3��b�)��/k}|m��H���v䝜�A���=k�	�-��4�E�b�t+���WY�_�]�k�I��_~z��5�p���&>�IF#�e�D� �؆�x�&͂��+�a����� �p���e7�Mi�|�I)���r�z=Si��9d��s�c!�i�a�U��~չ��a��oH�T��D=#(L�<�3���1}gޓ�����B���'{�KH�E����x�I�(Vy]ح�h���NT�6���y�σe�M�^K�vk{i÷�����9�2qLr�sg̴7��j�2�|X21�xi�-�}�Ղr����(FB�@��i�u���>��#��a�B��+x�������� kZ l̪�:Qey<e�p����%�l9�4M.b�sy���Q �K��+��Yۍ�Ĺ���_k�C�}C&��a#lw��ϝF��Im'����R�dT1�<��ϗ���<���o���������,m�W1�ڠ��bQ��yM��~�s6��g��9-aH\�,�z[�Q�8��:Z˲��sֲ:{��ӱI��N�f�a��Pr��P��݋~}`�%?ߚ>���crŪk�7ν�*�ڵ��H n��L�����+�h�g�D3R/��؊��Q�ȸ{��B<d�Ʋ]`ow�1ܧ����b�h�~�L�Ǖ<�:�F�1X�5C���9ci}�����F�%]Sr�h�;é�K@UDg�����z���?�e�/��8!c�h����p*:k�U.c�w�ؒ@鶥�2���9)������A�q����R����J����
vv����c���֟6��D�3C���<�3��C�T^�Ff<�����\�n�y�X s�̷o:�֚N���u1Ƭ�!�s�·�"�l@w6�@��X�)߷�ɫӦ+ÈS�&"lS])��A	�I���L�~��� h�K���׭��B �����u����{�l�4����y'�Q�s)��~�jq�_���TJ� �t�����H;�%$}us�TUEF�� ���Hb�^�]�6b�b]؋z=�k�Y����X���Қ�K%{��k�'���jM�SOM���˥9b;��1&W.c��9�Q��pn�*�g<n@��&C���^�öP��I7���h��W}��a�f�F�ϋ~?��y9�PUW>>Uq��nA�Yj�#K���m0°�JL��i��뵲RVju|[�d�.⋷ۈ!��3AI��F�$���}�s�B��U8=ڗ!z^��N��M����k��T\Came݆�ub��?�KS>tg1�=����;/�l�:��&Ŝ����&IPzi�FLrd�L%���	ry�viZ�m��y���>V��,,7�3�z����|�p��bt-ȴ�X˭[�i:�{4٩��(�![�Uŧp��s�"HHUѽ���\�IX����QW(���Q� LC�@���^��5�k�{���-���eoq�����u�LG�cg��Xǹ4R �W������i�.�BWPj� ��VI��$u.���T5�Ox/=I�9��rA7�^�v}	����|�X
����^\�!L�3/������v�bz9C�Xu�'L�L*XT��hQi��\��O7C4���SN��N[$�/�qz���*-�\Ȃ�w�@��"J{��:�A.C5�d�-�ZN4��Y�m�tWX�-T��\B�'�l��t0�=����vE�%*�)��f�+��G������I`�z���؝Lb���M�(P�+������ť��?��a�9����=y2�N~r=Y�?)�v/�� �Ԗ���hM�6Z�V ��H��|����{��{#�=K@X��v��Ll"	P���6�*�%�wo5�NYuo��	s"�װ6�x��l�T�-�OG��L�ȯ��~n��Qs���j
���������\�]��e�1����۠�s(��>��n%�:D8�v�~ٽ1��.�/XH���a��4���B��:T� ��ܓ��y�[,��G+��=9�=&��)j1������f�F��_вΥ�_��)���{�[@��EJ�K/F��ߛ5B���k>_��5kƨ�.h%P,�m+�k��V�4��r3��a�%$�t�JD����|���o8/
F-^둦x���R�����͌��^-M��-Sň���K'vp�Ro�H�����a�^(�£����qm{;�O�$8��}�pI��K��4}f_��$Yx����Qs�	��+���O�]�p���9�b������bW�ߕ,	�+��3��t|�>R�����`�W���e���1�RV��>p���[tx��Zț���>h>qiN�;����oc,�mw�&���l.��ݻ=Q���qo��°4/�2��3!(�L���T���d��V��`���%GX	����J�^е�^��m]�KOVe�P��3F
q"-V�2E���KT9]	=�ol���oʋ�N��A��́�߱g�@7����e���)�o����dl���ڢ7X���_�v���2d�֞`vx�쁲訂��j���q���"%q��o'��&e�D!�YRʯ�X�`g�ߢꑩ���+U��:�U�:Gz���׈��Q^���[�Ҋ���P����߳EܕZ�@U՛���"%N��'�, �tf�z1��2~��Z "�6��е���:��-��,�e�Y�y����lM��U�iP����&�����w�G�	@k}ƍ��+kk��e���C!!���P�G{�w�Y�`V�k��(�zjJq3��yՐ���I����}�U���|,n�D'� �Kʞ���*��?H��O�0n����ᡐ	�	m X��`����)˷-G�^�MH�)7�l��[�����FI�Z�Z�6#t(YӣVM���7�	���4���ѷ��)�f��!ߘ`�()̎�Y�8��`5��S�-W��t�����O�+�45(���ɨ��s�M!�醹Ubze�/���9�xpn���2�|m�U#n��q�%�q�P#�{U]��ȒA��ޞ��J1y���v�}���78�h�AB ė���\Py�����Ϗ{���UYZJ�X��0)Lqc�H��uS��Aa��ӧ�T�$�čz��F?SJ������c�zy%'�X]�c��CQ�3��Q~�gI CQ(r��k�-z�ۯi�$�,l���\�͇�"���L���\ ���k��S�b�C��H���O{;�����Tkq���|�0E�,^�}�m7FڈA���/�~��+v��|�߲1.�+���B�c�7�kx���Ĺ��5�L��B@s���6ae��q����
od�)���\��6�0���y�=��9TG�$��Q=���:G�"L!MS���!1掯dv�2כPÄ�Z�3X���Xfk���ҫ���"҅����\��M�-�k�� "����Oķ	Un�b���9(]�>z����ٿ�n��:W�W�r�+I[U,�;�o�.��ƗW�.$�[|>	
��Wzg�]���Vm�?�/%�:�C��K�托ȵ�	T�p�v��^Wk3#��UNo`�u��?�!���f�8
q�����k��6��=(A�k�7;�5\#"��JG*�^�O���c�9����:���(�b©������{n�՚�z8V�Z=����?|���83��N��&��dכy͙�Ȃ�N1͐��}K5~M�lt���t������¸�X��t��tle�� ���e�B�*�\MM��n|�x��Ԛ_-
׆%t�[
�3FF�Wt)N��6(�[����%���-5E�i5�ںe��Q��M9����?��y:r��n]�U��_�"��м.�t�DX�~pW�E��J��`K�z��#��h��Q_�:����X��Gɮi��J�ð�`+����Nd�( 2��>���z�/��:��޾���d��Nid�;s{�vQJm�r��-3�wNV�eָ��ڂ�ZNL>74S�nmK+G3Z��j˶V�(�
K?����A���q2�-<9�����a�F���8�/��lx��K����'l�j��<j�\NȾ��k���10�#i�Ӓ��t�Z�L˚*���8�Y�,���o�A��!E��#�iC�
�}�[��9
��q]�I�]����$rE��)��JL�D�\hh,�.*��	��p_���F�cMR������Ƽ���0�]okV��残�x���}sӴ� ��'A��#�0j7�5�pX�g�JI���_���s`�������ص��_�%�T����l�?}9�W���B����G��J/���1��Δ�1�(���'���Ⱕ�Eyu1?<Ǩ��G��d�3���P�e,�-���ی�ñP^rl��BYp���&2G�� ?�5�N���DhńQ�Z��)�qž(���+�6���tٚ���$��!��N��K ��r����?����4�B�َ���_gꢦ����1���1WI�0	�W�6ڏ�6f;�/P+�.9�\�eht�݁nԇ텵��W�%��D������aΈ0�`�)<!��h5�S����g�����e���U�ל<;�L��b$QI1V�#��]�!�T�K�sGuNUT����)Ι×͗[T!���+��qh�u�.g(�-�T�c�WE^��f�eCa��;T0R=��"����t�Bv,]kÙ�iYO�49HA9DC2ρ�y^�WR���Z��>�5wď�p(
�s��JIirN<�f6U�t�m�S� "i��b�垅�=E1JϠ"mJR0Wd+m�s�
`&�kR�`�j����R���3�eT�
zش'�%)�fk�R�h��ˤ���k���GBR��:*�S>���k{��PIS8�LmD�i- |�)�k���9��XN���+T�}�1ܭ�WW����|q�I�@urBb�&9�#��!�(�w�?�y�(��H�g�{���$KD�q�����$)���!]�����.v.`Ķ�������Խl��n�O�/��v����;q�����L���)��s�+��-�+t��x<�����Q�D�@S8��~F_��N�6��j�ÚR�U$a�d� 3<o���!�S	㆚���T�RcEf|�]���O�����?����%�>E�4�4=I�?	նZ����p 
 O-����?�������ҟ��V���)�H�Ǵ�w��I�&����#�g,i�c�M�C�i����E>��kJ�ո�72�=h��Kĸ D�Ҡ�v���' �B��ư��
��P2��a�P;[�^��-g`Yu���n�����7�)<Ƅ��r<&<�2ߥU6����53�n�f� ��;��e!˓-K"���@��%e�H�g��^��ݒ��Ϟ���ݯ�z@$np'JJZ؀/�n�j+�����w�MR�S���إj�y��M�[ 証p�?j+�?�KH@��SJA6]�y�!ู;S���c 6 n#�Ծ�Sj��w졪pʌg��*��s�/�e���Wi�P�ߓ)E���g{�u�H����JӤ�P@�Q�oS��>��uۄjPZ� zk����kJz�F�_[��c����FF�ӽ,�r^hI�*���d(�'�&�X�D��rG�[4r��y�n��NujS�Ɲ�~�����Nw!���Y0�[K�5'��n7�������`w"0B�wͦ1��]�|31}������Z��E���^(b�o�X��Rky��S^p��=�A��7�p��2���°ѪU	/��O��(� ���'�.�:��U���������\���{]00
�M�BM:QZ�Pp��W�����t��>O�~=�31�Y|Y�b�DK�L�L�_�hS���*�b��uL�X_�{H<�i��6�]� �։h���x����4ڶ(B�hE��!g�����4��oPwS?��b�TB���X��*<�S�t��i��9�$���k�J}G7Y�~���"�?�v���9�=�e��.�V>!�2��Qt�V�ܐgJ�K1a�v���rFd�`�>��	�U~���j����S�[�X"���b(�^[*����D�"P�|j��7�u���D�~�U�in���Z�A�@H���G�\} ����{��Kb��9�,2< �;#E�]�δ#���=(noUVr�b�΃Ŝ	���ARjҡ�Y{ݧ_�KOf͋���!��J&�OzJa��	l"�Z��i���6x��@;��s���9���z��7�f�`���]=e}��X)	��|m��w��iZ2R�֦��K��Kɴ��Ai���(B�/f��	jvZ�
/:�M�n���9d6}�YyK\j�_�s�ק�	V���>�l`(bYyXm�d������yj�\�b+M��b�(�8�:C��I�]�Y�H��2vabq�GX/[�P�ES���ڮu��9�-v�ц��Q�i��M��$$&�K�ზڼy��@�J+hB����B���5�Y	�������`���%F
EF/6��b�+�Kv�mn-�ٛ4"�@�R��r:������Q�*B��4�f�!���`]#{:�m�Y�u�z,[}�tj�.�����c�HN	"�l�~di��Q�X�ͫ��TW�Sl[���6[R���S[b�ג�n�5x�$"��R��J� �.�	C�)��_p���}�-�U8cJ�܄GW��.ݗ�=T���걤�m%w��|V�k����X];_����q�)Uӹ��D�뚀v��<�.��>+�����+
�|@�����f�U��TS'�����:���ω���c��\pE�v`UK��^��&�n���>t�4�J��x�{~\"k���y<TaQ�b8�e(N��)��G�i��Qꆆ�	\�`��K�����،-ҖWi"#%�?����� ��7�jp��c�s9#/XS�8�܌�Sw��yT����p��?���ڡ�R��L[�֡��~j!��FLͦ~�
�Y���,�EaE!i�7���T���7��0^���4?<��Ǐ~� ��\Z�3r;��G��hL��GL��Ŗ-�>q���c̱/�-�yc8���,�J���ck��q�\{�-���g���&[�����: (g	$lR�!1�����i��&�'vHT�����h�4Ů�c���8.2���� L�d��vpd=��a�;�'���Ъo�L��n�-_�3����ʺ��� D,����ԍB����c��A?�C��.Hq�7fg�4��8�n�j�1����Z��d�L���z��h�n�{!
��Z�6�s�5�Ro��v�m�'����ǻGn��CB��6M�9 RSg��4e�1��$�k�v�4A���ݤ������Ӌ	"��\N�:�*O�Ąb%�cQ�3�6�
=���Fм*tI:��-5��ַE�@Y��V����"u\Ŝ��a��K}��Z��`\���W��I�Pa$e5�j?;���ჄW�>�M�y{~T%����0E���l%o��ܖ﫩�ԏR�*
ߨ��6D�Z�`=�y f��B����zuԒ�g���泾`�	c0лEH�5Ը1D��G;=�q<�RL��I�L��`g�;���-<Y(��6�������"@�h��r���M���:r��4��$*1�p; N��f��tQg8<�6�j�/(�P㰺�֒�T ��`z�<��Z���,�7�y���i
F��>P�f>�P����=�NQ����	�l��'ax[��& L�Є�Gֈ��V�V'���r�en )���/2|t���%�*s��΅oY�Z�ԳV��7���T�(0���0�.R/	B~/����cl���ס*�B�mp��Vv�2�_��ٴ�pC�=E��d��~�M��5b*x����@{� ��J,r0�Q�Wv&;�Nc+M��;"���Dźgx�pU�2�aG��u[�rmG��/�f���}�dCR:���5^�НU�=�C�5x���$�R�}i�Q�w�S��֦����_D�.�\�\�Z���Ҁf2���6P͌�"(2��?�;7R�����<������NN�VpJߥ�b��G��K�<�~�)H�� �LN��s���XpJ��V�� )��Gf��6O�x�����5x�<x����Z6eΨZ����i��:�9��U�N��T��H�W� Opւ	ۮ#�MÉ{�� �7�kq���^��%!{��st|O8�^ �8Bf���7�M��_��q����g��3�����]�)��.dQs����nu���G���"�
q��}�C�m8��T��j�.i;w�����W��iEߘw�)�I�@b��Ek�݂H��0��۟���c?>X���	0��lj)b��"ܐ�/=�K<�u��f<�K�CuBKG�[^mN�R�p��,�*N��'�P5��lF�����������
���r!s��ig6cS���eP��V�=�[5�0�� b��
����qJu�dȌ�a�8z�l,m� �?\�
b����g�R��"�j���2ƾ�d�"܅�O�&`��Ǥ�D���%-�������'�#ԥ��n�/פj�~A�0Y]�D��\.�d��u����in@��_<��X�}l=�5���c���� Mm�P~(�#��q
Z��c��"�%��2�q�����eTN���̱���xĻ��A��v@\��7Q���{���$܈���"9?S�A	��[�xĳ�ʬ�����Tz�L�KK5�t-�P�{������|Wm���Gz�u:��E�회KP�6H��;;ؼ;���+��Z�M`��*���s��ղ5���C�T�fo�����4���Ta¾hfܬ*Cq
ͬ9jk3�[���&8��w腀|�'i�O'�mx���EJfV��Ș���G��ܲM2��r�X�?��!	�v��������J8�������\x��,�:�?���џ3 )GF}t���H �hB�k�4r`��q ���,�Ǡ����l�Ќ�%p�d�_����mW,ii5�T�	����R��e`�CyKSU�)��.�m��D� K<�~c��D�:��"�!�T���h�x[� �a��ȼ���L �[9���[���X曮}���)���y��K�l�Q�����0��n.���xp�Ux��oBDTn�UN)؝w��B�k�/(�ȹwk�-"��Ϙ���x�.NfD��H`�P��_�h� ��G�D��KK�X*��T���ޗ��z��鷼}}rSit�����[�MqH�<��!�y#u:,E�=���T�ړ�e��La�5�q֞cDz2oVk�w�-�m��ۇ&aOt�Zh�k��
� �9EO1�b@�j
*�~>�KM1NBˆ�P��]#�����T�7;s�%� v9oO��銸U{`wd���2q��&+��8�5�F��5LDN�ᕭ�L�co54$TŹU�})T�J��c�`7�l?T�{�9xD���U܇�7�j����;W��M2ݤH�Қ���RL�6�@�M�����`n�~?� :z9�>��y�3N>a`���4�?�9��c�C?9Ѩ�?\|�Ɏ��+�p���ř�`6��r�^������η����@�0'I��5~N�߱��׉���O-�#��~QNW7�q�s�r����������k�90P���$F	�m��m7��v�^� �z
{]!�\v$YH�D�;$��>%ž�����R!VR���ߏ�R�	�Z�s��s7���9�Q�a+���c��@��P��dVM�a毈��i��bsϭ��Cܺ��nwyN���zw�9 r��(���Q*�T����T�/��!�'&6�to^��	l�+Y�y����hM�v���&�wP)��>��S_s�@2�<�>�E�pP1�m�p�a��K]�s�u�ìZGK쒃�{�J�D�~7�~�R�j�������'��U ����H�ےu��H�Ǩ=6����t,	��˹�%�%7�.5S�a�k�\�.u�d��#�(fKd��;�$rt%���\,���(E��*�1��G���
ܭ�?W�WMp5�p}�0�e�"`4s��&b6��д����؅�u6�Dr�K�Z�7UGԳ�^
v�h��]ֺLvl���H�8FWaS.A:������k�"���g_,�W<����)��̉9�p�qFc��A�JX�Y���<��ؑ��n���2 zh�[u۠B��<��^'ঢ�{b�O���K5.�)o�.}���v��������T5]�xt����M�J�9,=3����S�٫s�)tS���'2��	���GeyKc��q|U�xѳ܋ߩv����ꈃd1�J$.�4?�]b��Ap�j�O�Q�돞��e�,����ޤ�.yBS�~(���a���������d��i��\�>?����}�2٣jo}�>���b蟚岉����~T	�����(�����
����,�����N9�*q�>[:p�+w�0�!ۨx�%��k�%h��{L������8���-(�+��D��r��=zN ^p�~MG-���h�L��<ɻ'ǨK�`{CɄ^�^?/
��;�C"ǫ;�`F��]��swSIo
��^</r��.�GmYx[�Ċ3Px��Ʒ��z~tD ��#m8��1�Um��I��N�Qt��FVm�}�VgL�<.�W4v�?Ul�6�F�I�3���Yq�dڣ���n���)����&	N]��N:�܃&�v���M�z�>�����[w"}�#�lMWR��G_k�ܝ��x+�=�g+V��4,6��q�	��~��,�$�Z�֭�g=p.権C�-F�V�m���vV��\B�?3;�d������@y?srb�
�I��Y1���zYa��-�n�<�<[U�o�������ʆh���>�r5v��8}��\rIF�F�Qda��^=op�)X�=�9a�M��k���� n<���޻)��J-Dn얾7k:���pH��o*sh��0ٵ��xIQ(����%�\�Cj�Vg��L籹�b+V�H6LywfTz�QA���F���8�k)/!�PM�����8z2���UT��"�_��f9���Ʃ�;�[�&���@8��;�P�R�t�:� n�cA�~:/B7��+mZ
����#h�I�k=4��A-�az'v����Y?�A����ĺk�q���͐Xe$��9�:��}��e2�7�Q��>�����wa�c����w�2�I������nq�@z�.�(R��c��Oc�ڻ��~����|4��>Я�7�i���^O�b���!W�Qf���6��s�1Թ�/(s@zz�ֳ# ��$_$��嶐�aJSLd�ڛ���)*d�Z�u�C*�!�k��2�yuP��P)�K㡼p�*5���\��Ө�%���˜�ݪ�1�!�9
v�-EG ��X�{��ﾧ��}��/	������u+>��ބ����S���q�7�-@G1�3��aX1�$5y��^�27F�|�ݶs�1�2��A�.�6�#�����;��	Ɛ����Yd*����O�i�c�l�&���k��^��Pk��`ђd׹�+����K}�V5��cuO5G�-�|���90�]�֨,g����(�[��)ql�~�ޗ�U �W��㔺�4��'Q�OG饊�L��0�7�z��� �ZI���3z�A�2s����lm+ȕ :6ԉ"�
�����(||.���x7Tz�����J�Q�e�ԃ����Zh�ɭL�B9}rzNr� M|��)���j�yZ���&o��9$;�em���K�|�a�E.�B�g�a����D�`~u�QYq֨�gn�He��A��;��?xЧ��~�Ty!+��j��R���	��8|�Q�`�M�ض�k.����[��j��\|:˳~�x�bW��qƋ��*a]�K�Oѯ���N&s�����':S�i���V�`���/'��8j���4Fe4�~����h*���ڴ�����gG1 �[a�C�a!��S�T�=a���G�:���b"z(��K�i<�U�!��+�q��P6�p�]ou:�C2��{	���C�z�ߗ2M�3oFOw!&�������~k��λL�>�C#�!�q��u84'y��7 P=�~j�6������5Pj
���S��=��G;��T�-��Le*0�Ҧ;	)A�6Q���l��\SX��8�C���Vb�¼��R�F۔�[�����Kq�KN9T���l�r."��,�HuUc������e�&����뫩�󍿁�[�JE�U�q����
����0 @�1{�{�~M��4��+�4_��y���;�xZA�)��0�A�d������D��A�ȅ'.s#A���B�Y�����sl�!�[sJ�p쉈h�MC����aK�{�KO�L�5�hĹh�N��߅ uQ�&1jH.y�P�cL��>��ֻǻ�0���{vWit�%N��*b:�F�.�P��AQʍ���ɋʲڳ*��1�W;���4d���b<z�#��Q�&K^��ɴ�t��#$/֋�A�tG�f��y��3p�Gq��(U�!���bM*����/���ɍ�sg�upK�M����Z$ϙ���e�ȽìeL�4h��sK��
s��L6󚆑�$�YS�3��m}a�);�^˂�c��mmbe�����K�K}�Ƶ�#��ejQ*����=��#�*)�i;�M�;��BJQ���BXf�	t+�[�) �c��i��]��؃T����
�4с\ �7y�A�!F>�ȏ�/���RP'������0�`Kj��/�%�)?��(�0�~J%1K�G��;�y^��u��V>��^i��^�4i���6�aHȸ�Q�G �󜶰Bl4��e�n��ޒ$+	t���b�W.�ώ��E`���u:�1N5�U��[7Öj�)o�DQy��O����i�����'΍�Z���/��;�OS.�C��W$N��ro+S@W�jM�{��h��g�3V���`�c�M���r���[�	��\���$u/���\?t���N�h#�����x��a~�h��@y�⃿��p��к��Gu�RD��rDF/u^�E�ŝ2��
�oآ@�[3���+l�S2q����''Q(����u(s���#�:Z�4d
*���k���1'��.] ?l��D�]����Qi�%�o�)�bM�b�3U���W[&�+-Oh.J���=�s"H�����I���f��$��v}��;o-]�C��ƶ�R�{he�` {�(��[ڦ��׼VV�\�f�g4��i%ϐ�߷:#��ɨ�>ƹ�9tLŝ�À87	I�
���k���!e�	�Y]��_~Һt�1�H �Z��?�X�%X}�b҂|R�%����^���S�;*_�>�����J�y�j� V>ؤJ�vn�M�m�Z+�^M��U��	� 4�tDs5z,�{#�I	&W�����F���X�9�r�%6�"�*����Xy@��ں�CTYP��֭� �zU)�y�����p�U�%��(�1����Q�/#ʭ�.����*/�M<�zHDv�6+�K1�b,���*�Z/J�e=[mv���i��@�Q6l	K���I�!遯&�%�֓o<����h�LWȿ\&5�s���v#8��#C)�OX�ד*��^_z�cL�#=A�G ��M����a:�1
&��'�.9rL����}��!_���&��0���_"G=4�J�>����$[Jp��\�Na����W��SZ�����E�W=����D(i+(q���h�&���@�02���K`8��yb��k�]�B�v'>���!<�;�ci���p����z/v3��2Y�-�'Q;N\h�z���6�X7��&����d�Uf��4Y=3��kمu%� ������>���eK%N�۟HF���4V�7���Ͷ��eCxB���/-.�X��?�R���'8Zoa�O�n!U�ߺu1�\F<����������i�0��N&����迿= C��d���=ݡ��i$X�i� %��h�3]��9��%<�������_ΦX��lUL��n���g�*��6`,?����׺�XL�BK�Y%����HۑX���@6{�NU�^=�Ah�y�5�_I��E���0�]&4]|,�E�'��q���4�z�����֎�5�<���Gw#,�:V����9��(���-��(�Ct%�����5��1��>a0�l�Q���G0��d�J�aۉ͞jQb�!L�����!ۧ������N �ZBtOG�������VQ*�N���������+H��]��.��"��"��33LP���Y��,��ަ:�i�EF�}4�У�hG�k��E��M)��z�n��ˊM�E�­�[�mXC�����d�>;�.�q��S�W���랲�RB��%%uWH����-0OF�>2k�p��ʉ�:�^��YI?���	ڥu�*�{:�׭d|Pq��1����S�b��`��9��3�X�6�ܔp�܀�K
�U�lEk�r�� (˻���^�#��B�APgψ=�t����+`�Ir#�6��J8���3?7}��RGcLO��#�Q܌��Ƿ�yxIʠ��MS���]P]���g*R�/QIvעv�-I&�D���|$)Y}��BY���N�K��ΣYPɊ%��r��Y�����V,��%}ָC)�D"��
��&�{�ɇD��>.`"N��ڙ��1�R-D[���\����lq�VF) �>���~�3��H�N�F>�>���w�1ٙ�E���NM�-��<���zX���[h��k9?ݸ쓓5�����EF�k��r�c��v��R�|��i��Zi`
E�Y��I+��o��;��#�xW��IB�!�_�/e�s��^P���I�Q1i�ܦ��g�zZ]AX�|Q z#���uȱ�߼��K^Ж�!=�	],��e�gB��k��H8���a�aM
Dv̑y����L�ԥ*a���Տ��<.|�$�~h�Ѵ�J�`�mCB�ԕ��'Q��&/�ö�L~�]�z����	je�a��O R�|TD���ρ���l�U�ە�g���E�#mP���Z�H:�G޳',=�eO���N�aI)p�I9D{�R'���%GF��r���1��u%�K{1 �
z��R
	������ i�7F���3�s�_��^gW������`�#W8�� ���R�e�?���H�t����aV��`����=Zٵv0{"�� �mB�>n��}��o7d����HK`�h<>�Fꮱ�+�]O�����Zj�,�[�z3_�9޼;�����Z6U���Q#�]#6�z5s���R)�P�(����e슏�� �j��*�z�P��*A��Y��7V�̿����m�XHw&�k���y��%Uu�P���y&(V�N�`ؼ�&��j#���۲�f�O�v�RZ��!�s�Y/�>*�����l��匤�!GbƳ�cD�x��������M��L�!�}:�������OI��e��x~��s8κ�Ȗ��垊��e�,":��H�6�+-\�d6�k�J*�r���;�q}ȇj��J
e���c��sy��A�Z9$]$6꫶<�=B���Q�*ͶN�	�ۏá��Xk,RU�-Uك�6��{-*J}�O�᪻�K���o�8T��p�&��ea�*Aci�c{�L����ة�{r�nľ+�o#\�3a����<ȅj	�A�be�����8C�X�z�|ցD_��><:"��!�̹}�4��xo�G,�Y!����84��?G*t����NAp��8{
��J��#���bY=6H��nD~FD��5F�ɓ'}����	�}�B �O9K�S!�~��Ϧ�ۢ��|,I�lr��0v�;��4Ԡ'�� ��$ځ�� ���BN =�FI��R��ѕ�?$,�~��ǒ����HP ۔c�L�T�� �U�ǆB���P��uA���x^��N�
�"��g���Ǘ:In���^��x���c?m�/�ܝ`(x#�Z�F��:ۃ�:�/a���9|���)K�����I8zJ��P�B"��5��w��+�Xw��O�&����#�P����L!�S�2�̜c���^bi��N9����P�]GE��jh�Z�{u@�B�1+Z��C�;���M���>K�꿆��*ѹ��'~-é%GM;;ϋ�	h�H�N#X.�.'tcUR��Qm�naoX��g|ip�Q&�^�{]���VNS�T�[��%B;"8r$6D�FԭI�Hj�*�s�d� 9`���yqu೐����\��}����<��-G6�n{��I��b)valLA�,�����:�������0�ll �}���qJ-��/[��� mG�&T�?cVK;_|o�����]��	��Aa����Jr. ZV�&��7F�x�r�X����ǫq><�`���9�r�Utp�n�K�$��؏@$a�/	c�	D�a�ܜL����IO�v�l.3 Bi|�B��, (�� �Wغ01x�Ĕ2%p)�fP�r�>��)n��i$Cm},)s^?���@�K�yI^�x�Z�<�sӉo+���B��BM����Mfy��Ǯ�jٸ�Dg-��Gӓ<�@5��ެ����DAh,�t������ґ�U�w�6&���֞~���Z-�\�����Ć�7_.�a��MK��Լ���FG�����cWjd�y�S�g�*�%�+@ J4S�az��>���{� v��}��ǳ;xr&��(�(�XN7O>j���]@Y!��׵W�,z���̚�8N3�E��Z��4�e�G����܉�t����\�ʖ?%�.kLa�\�P+f7�eY���w�	͛�R ������x4Ӓ�S!tC5��RÕ�@e�i|�K��9�b/����0y]�o�V<z���k�5b{=0HA�;�yփPt�vI�g��6<�g^�\\h�Vh}:�aj3z^�>f6��!�w]��/���H�u�|j�jչ]/�?��KxD*����
Y2g������+K_4��r�?��c?Ts� S�Z���Z�$8�Lj���J��>�eS�k?#���
�8c\�2U� U�L`	{�<:���֨�D�*p�(�\�%�c��vz
�il���2/�t�c>�$��*��]�g����E'Нމ[C��tT��X���~*�xW�o<F@7Am��q�~b�E���N.���Z��t�[�r�֖�SM^ޒl�L�3'��w���:�,W�q��Z�#Q{�"q�h\�.�f��*|W��.��kp����_�C��+X��v�m��x��/���;�1���p��Y�TBad���@9�vIf?I�M=�E����pȝz!ґ�A0���:��l<{ӧ�Μ!)��}�_���䪙&4?#.{��(�5ab<�<�	_P��dO��ރ�ڀ-G=��4w�f�a���*&�kS���*^=m�(d�`��p�I����o�����,6�h	:Ps��'.�����X�cʝ�e,�/�@q��Mc8��\���U�����p���kM*��vg�;���tj�@黴o��������d�)����}��뿤�<Si����E=Ӑʉ���&` �f�n�禎^,,��',IF�y��\gO�l���B�(u��w��㿋�N��� ��*��/�v1��x���Y�Q);� ˃�yl	'����L��S�y��ߜQ��'d0!h���Q+�	`�U������oZ{��q%0'�����5��4�oT�^�K?��t����p�+�u��V�}�!�2*F�gCI*΄CŚ��l(d`�+�
���{��O�_2}��U�b�KD�j�*�� =��$c�~�7��x�Y��P�M�z��>{�rv����䉀��D�oFZ�_�a㮢L6�m�f��ZW���ŏ(;�Xe̿�0�#H�����)�$-���(Hn����4�H�04�^:J=���^����3:/4Qc���?�Ip]'��\�E���.D�z)�{C�`\E�N�y5��]z�����L�&��8H�@�U �?!]��F�|9^��0���>7��9�O��^������Tj�p<g��-'��r-�N�o���	�)����G�ۃ^:Y��sj��E͎��<L��!�#i�zG�0��������؍�8��#@�$aR#V��S{ٝT�-�̖2��۽[4ς��$���'��N�k��ȗ��`�������K���}a��d#�`��R��[�͔��������h�Y�8��iT�j)�f|�}����E���tR�t-$WV7���yҜ�?F��ӗ/�/qJ,�RT'���yz���C�]4m�m @P.��ϖ*�F{���ئ�p���~e��p���-'�
��\�}�Ao9��9��&Ox�&ˢm+K�mI%�\��BZ-�`?�Ϸ;S�	|i%<ʣ-�"�P��5BC�Q2�cŶ�H�� t�;zÃu�oQ2gk�ؘRF������S(~:��w;1�VE���
AB��+0R!�[�6�bT�B����|�	�� �>�c���,��5~��x���c~ٓdhҫ+�e�o����-1y�6/�n���8��qG��ޤ7/�ʀ�R�n�ݾ��� |8G������˕���F8=w���qQ�'m���3�L�z�,�@�A��}�P���i
y(b����b	��w3�ܘ�T﷗����z��8��b$"ɀ<I��5m� b^�"�F2\x���3W��:L��O��ǝ�@���X��@�U�r�F}>K�h�NN1$�����0�ƆG����0Ç�eEٹ��"� �Z&i9(-�Ux�;����ϕ{pb�#�=J@Z<ɬ��f��z+���̑���1�>�8w�U����}��y-H͍g;�W#�&H����.M��䪣��M4�����E&F�;�`Wk��Ԁ��2�C��Y����G��X*��b�QZ\��+7�.��_�Z��c�%����=>+bBa��b�����ޫ檂��ᙹ�|�B;?����q�R���jm�岶^�^Ͳ�wG�81�}�%/Be��᪽8%^�)]b_F��:��|v���O=�B���^\��A�"L��_���Oƪ��a�͕u��5m�<{�������'�p����5ŕ/]j�p��X,�E�����۔G{U���%߰�
^�Q]�lZI#l��X<h	�xp�cgDz�~�S�-����R'fLC?_�WS�v�$�����
/,�A���k0 �$��0�\_)���m�j%9C�P��ȡ1�nG�H��?gj�y�REщ+L�O$���xa�$�O��� ��{)��!�c������ )��smeI��c��A�
��8�r}I�_y=��vy����Ms�e?'�B�(R���6���:voɟ��璃,�l㟖�H5G���<��2�Q��$��&MC��"�{�$��8�S�@X�.ר��w9���__@Aҙi��0rp�U��9޽�z���T8=&��;�֌~���B74����u��ÛŲϛ�ʃN0�rBiأ4h�������~|3�6��w�ئ;�_��*$%||�����7���B�t�4;z�b�����X�|�I2��'����TM�!���a
�W�K�������ũ����a�X?�@�b�wY�R[ܣ��*�}��/ ��!�]n���\�~�FŴ@��s��~��)I՟�5X��8sQ�t�1�<���������&�d��k�o$j��^!G�E�1q�T,�dD8w�5f\����1��%�G�w��R��A�d��n?�Ձ�𦴅���B�^��벥P9sJC�<A&�ﰍa{MUw�ud���ɿ�|�{��Y+�i� `�As�}�s ��q݂O�R����єm�]i�d,dEjǠ*S-��� ]���fƎ���$Z#q1Ҭ��5�e��S�H9��a�'d���p&���?6��Գ�6�C���ފ[��������
[��yc��Q� _�,�Hp"�dn��`�x�10���c�s��Ti$T���y��B&���Z�^9�@�t��Α�{͇�>I�/G�P�4bC`r�J;�y�z�9A�����̙fs��rQq�.����(��
K	~�q���c!����JM*���c�:1^^�G ��f78�b/J����Z�i�j%�,��Y�C*C囶~S��Pf-� d5,�<y�uv9��=0�l�j��u���C;F�+.���3�ݦn3��SD�\}$	sͲ�V8�ƅV	RW�5���:���/J|��\���=�FE!��MHál���*l�O��D�sD�O��*_�_��\�O� �l{[*�Mk4����K�<�A���'r�H��d遻�	V����F�x�]��?�T湋2��k�7VO��g���|w�)��M��@�`�x��u]��<�Ņ7n1�[�����⪫�-a!>�E���rF����w^���g_ɲ Ǿ'�w�ʪ��hŜ���H�Ž�eq�����b�J�!���3�Voͫ��+E��<�V:����Х}<�N�����@����0�����Z�[ao��p��Y�S�*)h���;�^R���5x8����J%���7cS��9{�~�H"$W��;�C�2�}��������ŦY�;u�9���*`p��]��u,\�n@\3�p�)�:s�K0dr�L7'#�/���>��+�(��S���vRF� �ŁhI�Eڄ�#���!�V��IĂ�*nb�ԡ�*�X$��te�>q^��$���b�>�4�A'�5����f�#�N���r�&��l(�w�����ibO��[�*�4A��#��/A�%K���(u���Pv�:P��P/35�����h�څ�D�­{�ǦAd{��I~v�t�l^RX5;p@L�ӿ?"m���<��BgX���!R�3W���e���RLaK�1/l��.;�%k&U$�I�?�v�:3˳��T_�w<��������������JJ��p��{�$_��(�
[~�r1���i/m܉ԺB.�S��f
��z�-#�q/�f< �ױ�Z��zJ��p	��!�d>�,�"�K׈ľ�NX�e�=�V�������Zn@��jt���W�A�K�F\B#�>I��� 1^��ٽ�I�Fg*!F,���ū��d�<!�� ���}��;r°P�(#�	viMB�Cg��8�wɽ�S��)��;i��W���Ð#�XO:-���)�U�A��\W�}�o��ˇ������zFD��0��kX���{҈ŕP�4���?y�X����P�|_�"CҊ���}/�{������� �����=rϬFg�i-`�|�8�	vHQ��Obl��>�JN��$��>{���k��g7��)��{feBy|�TlPH��:mϟ�h��ᖈ���Y�^��I�-��x�;O��1`��odm���1|���`��s���CH���a�� ��֕��z� � �ȗB�0]�-.�G���8�&�oi	"͐�.�I�N���{����a��MH���t�D��-0_��_F���:����*�,J���K������J��g�����oFNfk�b�Q�4xM4��Ǳ��B�,//8?�{�V���VJ^��Q�ˌe�E�N��K.[�����Ar�.d�%�f8$����༆���?G�	m!�N��3k@�{�_R!��,~X��H}��7r3|lq�\�K��&���ó�(j`���8!��`2�ݠ�&���f�}�Ώ1i[a�bǨy������G�p���q�8�st�2[�CJț2�{-�U)U����I���U _�?�u:!9�g_�J	�U	��y�4�E�˰��ғ�ϖ��LMz0S��u}E�M
��h�/���G����C��*�y����G��M�;j9�͐ɿ�[VB����ފ	���f��WS9�y��1���Tg��Ͷ��Tl�����z#�,珹�K֢����G>��q�x�
׀}':tbC��U2b5�O�����?��������S�C�}��_�A8�Y���Y��x��`����s3]�§&�4%+b���#���9HkBZ;�'?��U��$�X��4��q��<]cN����O�^��iE0�&L�T���Zn�s����c�e����V�v�/R����||�5g�'�5N�9/ċ��xwq	�j�P�##���\/��QP���gb�zd %ms�M����eP�aE&H�fJ��h�@&�i�bA>)�&��M��/;|��O�7��8�)²2W���
R-��}�[�ȩ�ij���u���cJ�g/w�'V�=�W�kc��\��d$��/����%��ߌ��GD��-b�Zb䌄,�`��3V���2%�$iه~{U�W@/$Wp�ifK>.0��4�{��èXP�����Upg_k+�R1��[Ν�ٵ!��2_LC����f����D��z-�x�E2��d�V�2Ҥ/11��5�f�!
 i7��ˋM��jO
�Z��4�����JƁ'Fa$3n	������Z��"�v+F(�I4'�Q� ��8!�F�	�$%t��IQ_
w��.��?�r�e��"�cN�t:��ɖ *��j�l�,��gqJV�;�7h�]���*Q��D�O�Y���y��KJ�!�