��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	��4�/�U�~
a�z�K��6KeW,��
����}]�?���۩��o��Q�H�L�	�9�LA�'�Y�)ˑ�D��
+�X5�?_����@|ϵM5�f+.1l�7��0�Fbd��eU��P\�!�nK�!L:Yg��iT��fj��e;�'5�ʩ� S�⻴+��[U؍�)�\��^#w"u��"9M9�$�W��Ǚȣ�:#���v�	- ]��vc��R�߷2��͢�@e�����r�A�c�}X�p$4�Gft��g�8Vc���}��BQ��^�a����c�L�Q�����Q���ѧF��
d�R\�%� ����QYC�T?�m�i�잴�E��.��=3ذ��x��Md�x�INu;.<�H^׉N܎D�4��������UR���?�̱�p�/b"~����<|����ICX�V�@S��6�o^jB�4X��[��Ҩt�o?��A�	�B��)Ag���ܲ냨�f�a��gy����/R|d�J�v�:)�@��wk���Ğx�n�v
�]��X�旵pW`.�q�����T�X7_m8��2��Xn�C�����G�Q%�{t�ig;(�l�_F�k=�uA|K���9<p'-���Z��<6
wq{��H$����Ye*PYI`fg."!����m=���3�n<��q�G��=�蟾��[{VҮ=QF9nH�G�/�-y��;@�Y�f�}F�(�ْ����]-�-j$�Μ��83�����}����m�뺫w��7O�&�o{��[o9dg�I���B������6�~z������!3��]�嵗��;<0I�G_�U<�G��(��5:V�O���G�Z���(�G ʺ|�ʭ�r�1VjN��5��{��kr��DH�x#$��� ����Zh��gz�|��n�up��θ̥��U4Wa�d��Dp�Sc�	a��!���@���Mi1���4�feɟ����߅�3���Cud{��7c���E��p\ۢ	��m����:�&QI����X��_����r0�x`��a *XpSln����
`z�h��	����50d�ܩ����k����miC���V�߀�����`�.T#|��j�X�ف#�:#J�\��d�5�C������58H�Z�����#ysw��E�KM�ҕP�3ζ�p����5���v�-�"P �A`�����+�`UH�RP���>�W��U:��vI�)���.<==�|X�{�_��iA."1��j���d�� �xG��]�B	x(���ă�_O���+ʟ���>�f��\y�aJ|t� վ�)�mq)h0�̶�g��@K���4;����_�� �3���!��X<��<Q��#�	:ԩ1������E}�s򃝴����T�b�������5ǌ,�-�:�_ʎ�}��:�H/殌��(�)͔��݇?6	Y��z�L[�#���;�,�Λ�������z�7桍R8�aH�0��2���Y��ݓ�2�����*���Z<����4� ����֟�~�{~0U샺~`d��e_�
{А�kh�B�_+��������.��_�	��c
i�8c�0M�m�?[��m%��nDֹ��9@�!�=?%X���c�e���7?�=L�@R�	�_5�{�|~;��Zx�� ����~v���d����,����R;b�oڱ;��.}�0x*㷳����L�g~�tʩ�����$�+�a[P[.@��*\��k�i��v#��z��aC�������F�����Y�2�:�fq��!�DJ�������(�Q�[	}��j�]*E������8�e�M�Ρd��$gcq��č���x;���a#.�>AoS��Q������.��j>-S^�Z��^2�rY�>�L��m�Ep��d�O�pw����M�*��� �\x��
���`�?	̀�*�4����|�+�
�����'��懇�xC�!倖�q�������Y��D�7�,s��?�fڍ��ĺfXҰ����'��8�2�,F4,��B�_�O�U�mx5�ӆB����@Uq��.!+v=̒?�V�k��H�K(*��F��-@\�9*�¯�u"Y���E��)����j���9_VRN��<���&|~<��v�e.���w��e�&����oH<��~U9���
8�LX�S��MU��=m�f1�;���H7�ok��Y�K3�7��ٙT���kd��ϭM��;>?҆�K���P���,5༖ӻ�訂�S$��#�N_�C����S5k=Qak
L�?4���}��<���H=�Q�?�'���ZB]����m�bSw�u��m3�a\��ݠ�06R�kE��)�4bK�ڋ����x�/&�8��-����F�W<�i�/�Ciˮ*ݱ�_?J������r��D�t���oHm��3��d��K� B���]t���x�t_��f��L�_���|��<��3a.!.E(/@�d���tUh�P�qn-�4NZ��R�]샃Xa���J�}/C4xhb�}�˹�6I��sc(((�n��%�;�F��(mpW�Uz��� ���ȃ�Cv1|�/zm���%Ba.b;�@5�J�/�h7�yt<�7,=zo�V#��Ȣ�>�b[��6^�@ha}����N��R' `��o�6�����T�,�U��c��8�8ԪDj+빱ʋ�;I_P�+3���35<*��$?���c��\�
R:����]چ�/)BC���@���&<�"܂:p U��������4��.�op��G��O6_rl��ч_���������%}E�N�P�({�xI.�,⨉�;2Gf�
�N\K�k:q�[�ڀ��� 3�s4�����#�	�*;�{]L4G6/���������r�z=�1������a
��1?#��;��?��D <K�@,�`�ĂM�B/�sY���32J�T���� �+m�i��U�^ �ǘ��a�2�.�B:�Hׄkm�)�K��`r�]�'ot4�91��z���o@|���v6.�L�%sZzjuD�8��f�F��� �L�m��Y�}��L�.|kl1�a�pÂ ��j���KXL���(�I�Ǡ����v�ᤏ$�lY������5��Q�_�Գ����B�@�*�m��ia:�Q%��F��o��G�~�@Ev�u;����_�g�=�y��J�E��Q'f{�����"����1�����e��@V��r|�ǰ�hT���$�N	�n�`Y\����G���u� VK��.F2�_7��eD�'Hר.��ɖ�86M^�n��eR�WӰD�B%w!ʟ�p/w��2�׎�aGmO���g���;��d�ͺ�~Ȟ�q�bwؠhZ���iA�Y�V	/�!�s1#ҐN[}���	�_�	4���ޡ:�=l�(��������Sk��1x�U�����(�ԉ��XHC|:HLdE, ʪ8�_m��V��`o�@��XE˴)h�*21�&泆���Mb� ����fX'\s_��c�:�<��+K���Z$R�|��<?~����N���"�+(L���҈�o\�01v�uiKG�t�2Χ"y�F-�~J�/Y�,�m��)�bG��]��e���F�E�Ѫ�(��ޕ�� J���Ḙ�3�|�o_?j��ҝ4=qL1U�j=��p�Չ(� ,
�h�T�13x�-
��#�𱺡��{�z��zv���.u���9q�n�J/5.�[?��sS�j���iH�G'����|!IJ�f��hM��J�A��%<A��T��Md�	�� �h@\�$�No�?۵���l���B������\K�vJ�JR�˿Պ�U�w�j�	ct�:�%G��.l�ޢmϨ����D�>�7�9�	��a/�����9�\0�OI�W��wC!h -u�[�=�¤�K��ïe)֧Kc"�98�a�V�KuO�	� �y��	zdc�%4i�$�ͼ�U�H���뽅�J����6�3���8f�4#�T���/r4�o�}��D+Zu��p:�����v��(�nuJJ�]�W��b��Wu�X�HV#Ó�^�V�G��`�-�{��._*H��u�+�9!��#
���D*0S�,��f�D�$bp�ݡ/����0��HEso�f@7ϟ�0����?ż�߷������<�rP/�P0�;R