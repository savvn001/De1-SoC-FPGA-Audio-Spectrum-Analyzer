-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
smaLaAWHEZoywA524Dckw5Db7Q1yPMAiM5vC0LkVUDJHjz2uYsJ9ptQz7X/w3reg8PMPGix7U6eH
hIBaGAWAMxb6gRz2nEmXpc/u1CWFLgQ9J6tYv3RE6jtpscylQtWBQcuER68MFQtudaR47Rgfe+RZ
YDgw+SokIYcPOgXOPdAwUOgfle6smvsmD1qjtQzJJKDEB6MWvCI/HZ5ltCqjha3M9CpdgtIP1IMK
UebYuVYTd9t7U7L52ZlZHXkQmcC0q0oDezMwd11n8RcuAONzQmoev250YHgZb0k0AKURGd5xA6hL
GnYQ7DlKcrXpSmHMHZ4p/szF7aCsDTDHwS6k4g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
MpCpRuNK7o5ZXFrQzdY+L2d9d72Tpa/cUITpGRmUdnldhMyATLrIH7vHqrHCOn/Yo8u7nYv5lHwj
rXl7cV4Vo7H8jmfhFr74v1CEAe9QtFAR/eFNPfLp/32rqpWzfk7yJrc9SnaWNfzlQJJz5D94NajW
acKD7Xm/H+edGdxbGKbu+oCfLLs4HBuacIji4SWmCkAgVXlkHjiCDVG96M5usxWNnVdFtIW4zRWn
B48vdxlHrO8vShAMljGaYKm6sZLsrsHT/J7OL9zK/qcqwZ++BmwuqFBfP7xgnOj74/nPqhyxAWBQ
t3mGIj//99po50dNXSa/Z+HMrOvnCilAYQwNyWNvQimt52JQzSiTuuwE1IAB/Vh4NMQFvHiNc97s
uapTGOPC/mrkTHNJ3w7ltWyQJ7/OeTAmm3ZDEkIgNdrioGcIbeB2SJ3YbCgeCG8bpo07zoEtLrQr
4AGZgOZ9GlTs3lKg9gK1qwBTUkvhlvtqPhrqnWVy196GkZwVxyOBL4CbgssQFfs33TO5WspwZkkJ
KNTLtyESpiiO0RHFKGfcMbKm31J4WZ+4XV9+nd+H5hWR5jUXu4eRzk1xc46Z8/Gwv8fCQ3+EPYxS
jdWJptlzqbsp4LiVGC94dWQCK8i4m4cC4MEY1z3H/O+qvFnumzBetaAtQE4OYWevS4/6pPb2vDW1
js4SBe/yEmh9Z6b5fQg6zW7yEBUmh20qlL0mHJtgqvESimJjo+P2ihCqeTP84eqkYVrzSWUuacwl
duo3DRrKwpPwbF/Td2MdhHEjUbqUiW/Cid3tvldoloMCgdnBnJdMRZTg+WrYCnXpTo7ddJeMTsf8
3Yn60Kg8EEMFBiWLnG7W77JXMfeV2jkMOKZe31XnPsreQldJrPR2932vq53QMS0MT+WRUopawI9t
WEdGLgCSyQxtYbaIl6HtBMKFBa/so3IZ3/RoumTkf8xyKf1Y+DmoqW41iGsZs4no1cUk0lIsTRH0
1bpqkCCl4BtRx7FK8ssqjb0wB8t7xJmjvy0tsCbFmTA9EZXJiMP6E7n+9MQGyCypE/jifgKp3Z6l
AoVHMqPHcELSbmHSlLjtSjW3qt1t++m50xt0d668yW8ygEPu9WV7uEY67wTJfnTnCwHi/77Y2rDi
oRuhuSNHkqeWmkGZrCUCOaVYmFBZr03dQVLxB4saybB0+h/QO3RYEDPBYvhdis71+sswvXGu7Sfm
wHKMkmBENuds/ue4EmEz5UrNZuo6ixBmmz76jJnuBMz1oiSqQBrpWbAsH1NSF4dqJXmcaxWrELlt
m1Cyc+BFC3UxMGbnE8x/XoffpkAK28yHWM6wf+y8dREmlLki5wH75VsRukn6e/nbjJmAMvSjmViw
ANDBHqV0GLd4u6jD3LyIk8JkoXjtzO8q+u12ZGhhSahJ7kL1/u+WbbPVIH7AJC3ljLfwcU2OcWMS
tMVw5Eb1O7/6Vh64IDtFpz10wduiSCgqFMAtfRYbFIgMKHrJ41maSDwjnfgUJ9GZpEknKEcgMpU9
unyuUn3cUmc6GFC84+avSg1M6fMJOR8aSL4ZSIfNylhCMzczUVylSUBl/fa8R+Zvih9Ny9wox55v
A4s+4fIDb452XOia0T1VH5oQmu2QyXqfcp0EJAjuPAa5MKcV3pGhhe1vIi+vX97vnXHeh4NuNXgx
85oYDIuGgZBuXGTnUXYK0hZ16gv7WRcqpTUtMrHTFH/5LHpb4iESwKQFwpH+JBlNiK+3Z80LhFay
34GxFtuntadlFiLAevUuyXLFM6LNhQzlP6Gi6hyq5lQ4pFRfBPUoUwS42RuypdqTOTPpwMT8FZqN
N5XtAKH+8fAuG62v+DTYp4aonAAkXzav/0FWHq8rocsFeN1pZSFYR9tqg0aYLu4rm7V4yhBc9toE
mOMReTpDsWQLV6Xid9ltsu4M1Ef2gC5+InjcCbp9Y0WqeFSdubg2ymk0nFId+zjA2e3Ur0b4MHru
ktdaSNOuC1agOMH5nKPoAQg7EKZR9eV+Z5TgXa//Jp2ZLinQs/08SjwTXGGKxW2fU0pc9sTEcKIX
0ATTdCuzLcqeo68TsOYJNwO3TY8FT3tA6jPLYVSwz6O7GbebsHdLWCqmoI2BbpBzgHtgCoiS2pkC
kMYRUtNvXJM+F/cM8Y6aZY3RM4RtD6EKg0hbb1NLPz1Nd6+dtpTdQN4W4duprW31DoFcJ9BYHmuP
RK3YfN3EDmyYSrZs/wMP+Gyio9qzR0yA7GG56ADy/JAGjp42CIX+HrLtHSQZ3fDUlIWDifOCwVFj
b7ZjMlR7+jKNDS2bbsDP+KYqBgzXvZayghWschUtMlnjZySZkTL1nJTF/E/lOIHvct97AklIB6mG
U8Ax1Pv9dCAupzoxhIRv8RTbMbxknOdUuPTdj34whvh9Fdusb+LQIgvxy6ugvBbUNm4iP+tD8u4G
a4wBxz0QxMyd91zeCUPiz4cDTsZAzNn5V9rt/rnGgb1upd+pr1HmZSqZp2GEuag0PDNP0O9GpFs1
qjig1moN6oj6gK33REpDBPWULYIs6XX4IGi8LTTu+IXmk2nmQC/hKiaP/FNKxJsSa73n5esEfEHI
jkggMu1EFC4o5j2RJegxMo8DTuQj+/eao3fA5hh3SmmcINEaTOGKzy3fGwUegcrh48XFV7iE+Thw
XmgwC278igxj89eYP/X9pjlTRxCIpPsza8bVlTXpKm3BBr55vpEv2ka3txRWdUSsPglsqGVZhGcc
GKmKWo+BlsHeiKsFKNCPJWz8oxjFohWhRs9Nbpb2qOgNaI6ETPCl6g/SH9y8y19FypoDxB7bvj+e
wFCkrZp6Dg4CpWbGf4UQS0GFCpBxQTnEY0UJNI9GF+vjz80lPUbgVCWj+pX+0/oINd3MuWRhuWrr
+PvudgP7qo4tRrldvx1HMQXkZyNqMKPYeefyFCUZ1Udw/+25fFIlgzZtwzWfYZJkAx14bCO94rss
pFgY3opb5DGs0xPL38JnRobJsiOXE0Ow4JnB1uoY40jXlAdg1hGtM61GgtdVvOuJEMyne56QJNGW
dj17xO+FpybwWafcuboASiCXo4rTxMdjPNP1n2vppnVV043bh9T4SXjj3tKcReQD0Fgli2/MrhqP
4DsOSO6/Su8ucoFLCMjyV6sPa0iR9F4P3E/xcH9gE0RY/exSLZHPH9qL3A7S8ST2M+3bd3s0cMpU
CNbxXVteFDE3EGQZzKVeif01wtEMbC4N359OxXGohL/B2zfhLH0RU0G5Ju4StXQn3shHW/+H0Yra
hWGXIXyJ1lZgr+cCA+OHWBHMw0DCZ/AoZy1h1Mo2psq+N7RanVgEgUO+kH1lVF8T7aSxJyZ6+0gS
OX34T2Kcfk8LQuI6VVYVP1xPc8eBNC2QpaXCZH/f4WPPM4PdBNEyXCcwCaFqMVcQi17PFUyQVPNe
3UxckFZnEZ0aW6jJEHmDbjqk8JrxHvAnzgXXcuivC1A1lQnVJc+pU2GquIv7bJcIfvmShqNe/7Mu
Q+2RNAyUeQoofC9gdGpx0TH+pUj/B8TP+NnajE5G/H/R1czm568xgBgE6BnvivaLHvqT83Eyvmk3
jhAvXWbvLxVM/A3DluwdJz/ZMBHxrz4A+oCdq2k39Tq5eqsDl3T5U+AaB86Qg0hj7GS9wPvGBIQg
n30mPCnsSzzEpgCN339HKg7XyOq3Aec7kReh/xT9Iymkz/+tM1wAGaf0M/hsqU1dJceSbHJhNnC7
VkoCHXJVzAP1UWK6ipbM9U1LEtcUo5jkvcxLqpnzyWTE32F1bWratGwyFGR7qkkElF4L0zO7UAF4
VSpysTsbkUynJIw0wCpOUXuX9D59ibaB4FpyaO1lZdYHXe1BWPwkobCc2QOaIbuSBSZYSS76pkHo
2ExEZaKcY2LJ+Yevk11x3D7100HjYc8KBb/ocCHEkS5gQ2bpELOGhvAqFay9m3YmCEgydjR8lGpl
V3RBnNGSzbQg3ysxK4tJUr+1M/Lffu7tYZyUes5WDNgDLzBDjd4Itjks1+g9Guc38UWS2MJns9ge
IHPDoyKRU1nuLGwonlz8Tz9ZY3UTA5uzRzxxvFyA2ZCQnexofYqISeW0hDHHNWhbjnWI7XZMR0/M
de7Vtgz/ANNM17S/HxK1T8r5Ge9N5VH8BsOgRy6IGn0tAYadHiYyQjYT/nplswzHG7I4u38cLw39
UAGChl3Tv6tzcMpC3buW1ykU8j5pu8+tWLi9lqIs390NfgsSiKJXXg3TSvP1fBVQoEYlkJ5/IdxW
kS5wz3Nlb70PdBbsmQwqsjeq7HNingBzY+bE/cffeNYwcNMXyGgqQwtP9nSiPOFardvs83l59lce
Su6m7xy0YeBP8dGyg0hr9avgn8JQ0qb8hGem1ZPED3lUhiuy/uZeBx5JPPz/YVYBoli3sHaZ3HZ/
CDxtz8xVcAKqjx8PRzYi53yMTo4TCyxHBMkRp4PrcCbRqc99Q9w+9sVFH+NMuf7LKRVIMwF4QM1z
lBOnOZIZy271ai4JAHAyOd1GHPMc0IJuMiyYZQnKEhq81UUSo5PbeDBRmi79cQXb8rJDu29eE2CU
t4AZSY+7pXXc9fJZt7jp1eWCvX2UAOV+kWLBj4TDvCJ7uT2FYGcDCSewBiTMXNEDGqDod0lBm6AR
WD7KiArl2LD3yupEZK2FFxppY1YEbx+5Y9pK39qWMEYxzLfz121ehmNJpCnueAbeYbRzW5YgxL0O
k9NRL10oXcFDa8jfkSvticFRiu/R3HZA4vlNdmhXqqo0YMF1+WRIYajNkH5f2E1VHQEoKP1Xq/8E
5Y7grm09obhmlSnDZcI8LvU4p+kXtB+1FJv10kLa1psrj4mLtkULDEFKXN1NM4C7lyRmkD358pp0
1XICTfKsC3kLHtZO5bscG6msRGD3GrGELnt9bya+EVMalgk5qaQ9toqYulqJKq7EPRthO5Ig+/g3
/HXEBnEI3ZUOJfENsIWxRNmyLvUcmrrotTfcGk6kumhPl1B9xnzbHPCyrp++qk5w8m3SL3tZym9v
3YzeRG8aREbHsfxZXmW9TZiHqxOsajIroMTeVArTTQTgpEP326U0YtH6xds2689FSko6xrpMjC2A
OxXKpNFmQQHvHoVC4/bJL1L6GMgvkuhjdcYniejQoxJG84RHixTjkj4ltmOxIwbuWkefAjwoJXw7
EWUseg7nJes7OdWnUFlcB4Np2twyllZr4He4CJXkAoq1cGcYO2S2fMJ+OL+cE1SwWJCgRwbr4A1z
jQFkJ4W+aBdSwol/vQTRiL8aRyDykykDh/N2S1qtsYHwR5TUZCFRt+1B16Ud4YSYv7fH1MDQIBds
2Vro5kING0HOzpB4ivtfwTz78cyo4LV/RDvVNJ5eiZlhv0vRNCFsvdBVapz9wNeQlA6dzVbSbIAd
GWPtZcpp/bIFb5ekqHWmUwj2sk3fUtFtLVaxq/XkJb4JcCD1MqHYgpTLiziq/M72PCh9wL6gNTOm
sci9oRUXD3PZ+xlEHxSQYZvnmvIaVcfe8DnuIL0Ifw62nB2lWv0IabAq2vyi6Fm17x6cqZBNJy9T
wbt+oAhwN173zdWUxjPMdD5ts/rk75BXeMXjx6zMgFYqCbUdcwLtxjZCGGDnKnrMCeDEZjC7R4R1
cJoXXrMdGXK0v3X2XPxFJ7BylvmcyLncm+uJCaiLKMkTwh4usPGWiBImqKMzF6K0wKDYFk1a/zF8
wx5o4HZ7Yj7OH7Fmidh0TFrrw7ZCcy780OWOZ4GDLppnPSOmUE5x15I2Q7ZOrKLuk0xQFYScBJam
XZZFut3QpeN+Rmz9IRwwzEjXcXYCI0uccH6jkLWT0yk/8E7y5v9XptdIPbD45bEyi2safrWL1b3m
Wiv77waMovzPIyPTiASHqQl4e1UIouzA643lbiL1oRjpF9RBrygLrb1P2A8PbDDrlgpXK2ES2b2K
NzivnUTh/Ljiw2GqINPapKu7x/DPMmrFrajPmzbjtAFH5UN4+QgHwHnS0XYsplBUA8XVPOSV6xLB
JmXszHEOxHP0ldXDVicSBY/W9RJ2TC5Dkm1Su3uIQ5R9Ss6SfsWpS7ZiTT7b4QaI5i+r66DIXDec
e2X6vRyIWSQyA+J68MB8GtLshTSa9wnM3r2EYuMNlsb5z4vnmcFPfTqF7b+vAm5qDcEbY44N3c5Q
A2PJRgFarW5oUqIGGn9lJkLblx3WdNB16Ycm5Gj22EaGXF7+nxK/RpqlkRzbFMIOuMIyPzeCNGPg
ZVtEVtRtOG1Q4PQGxAdcUTQXS8ocVYz7kbZXXckncRNijeph/UqFcXy1Iw8DOkf3V1XwKDGdlO36
62avCfrEoAneHI/j5jhNBtpnZnXzLeME1tkdKHmMi+b8H8+F/RFKmwvyz/TeFBqz4kiFzxgFsjhC
4wwKcGOWHwt+VBcQwPrLfOvWlGFLk7hihJoWxSixIQL89Y3Dz7SecupwHFzbAO4tDD1bW4m57xcH
OAO85xzT5b1PfKz7cMcAIHL6nOIMgkvCX+FcTk+I75Y6I6NurCd+BZhJzQWI5ROtGLeaYlg8gyyY
KY8CVqCEohmANUf+XohqLTo4JDIeVoEPy90eEA83sbqZ67i0khVIxqsfe5FV4mJjybb2eCw42cSe
saP8VYFh0SWJLL+Y+NoIHpDwMB2AO0AyGWVW19t5z/Yb09XSXjqUaU+4dJ/hKe8RUB98j4Ug2KKI
iK2ZIFuS5EFgwU9YfCTHxucCZabyIFRWbm4e51W6Q1Xcis/K3Gfmv00LG7ZpvUlBlIeIxIplA7rA
EwmKhez2JtiFo6qwi59haUkLUpr6/4BSwaDPEof92mt7yl9V8g7W3l0oawlDKtHwhGvFdc5ruvk/
Brdoft/nIrbPDpgZLQUTverxsGV26JUyce8Cq/lV3yhBVDKoRa8DecooH4AloFLypqQtGeZX25Gt
Cq/Tn3o4cdVSj5NJfUAt1AvSeZtVGdtV7Igsp7mcuT3nC5MyZwDlYBeqvmjur90H4+4u5+mk9/kr
rarq8FVyM6q8AZXqz/RbGtWUEIeLIDYEcLniWvBJg++FfROW0MTvfMkQbvFQgLWrfXR70NLgyALm
wXfFoPmCSPv0yVOsc701hP18htHEoJPxejI4cYkJMGXH/epD3pc4w+4rTYh5cu1KL3uOeLu1c+G5
M97EzkyUYp8G4Z+Bp7kU4Aa7mRPhvTycORXC46pW82QV+OW/MwNzQXKKVY13v4GQqkdpurbdhS2G
La+YyzaRh4gjIH5+y0nQP7pL1pJtukL8eoiPcqLiuYfAqk0pF05UsDk6FPUbbd6icVB5OC2BoCwS
p4cw+adQMXD5ZpZ45AP1Hc7uDgxcb6MVK3bO1yFRh1HdvtS7yRiKWI0gYFax1YvazvXxgG7UzaHx
mnkhLgYu6o5K7H6/TYIiFzMqDHhTNYkq7GI9qN2OxbLGeicihtJgHmspjgL3lHRx+rVQFk4y5x2R
PiDUgFfQoLxPqyTLv+mjJWC7Ut6wpH6rhOGpncRFrNUrUnz2dWjkis85uhJ+iV80n71BTHD7PyQx
kCbxRCWINYz/VNBEUvDATw4rY8JWPdlXFhucCghOQhrN1GfR5AwhwN8P4+80VYuYQXm/iVZG8f6y
aZRAceyquQRyZhSCQ4he4STaJhR8b6ydxt011ZD3l8EdHCrZi1O7UdfFA6EB8befGQZby/zDepF3
6DrLPQQ1QvZJk3KEJoWw/ZXQadDEDxQl43n41YOw1BJlKA3ZweAFTkb1HnqWPenpcG1vJFBhAeyA
2XeHNcAMxqKYhV45D1tsbyQSk9EMYdQgHx43P5wGJlVRxPnei9s/rP9rivYKBU3ny5QMIJbTn6us
83ir7fQ+wsEZ617ZS/6ZAYnSQXXz0qoLj0ayI39TaYUyXo1AICKEax5Pslc0jR5t0wQhkCMkFUXy
HjfZdKy3OQAoj/7opf+1RoIGSJPfLm7KM5+PYC1reEaCg77gydCDANKmUROZcgpVsJkbm5QRanBq
JVH4NUqF94TdYMSIx8G200yMZVthGCg0ZOB/jZ7bIosEhWxiJgQOxjFZq/IWzZ/8mCdoC9qOr11B
5B7RjPLCPaS3LIN9La/t/614YEuOuB0KY8TIk6GPsYNUPz2/NAvURk93g9qRYOLVQ+RAA634CLlT
rm7rDQ8OqrvSc/nURwWDqG8GJCI116fqygp3/h4+8hh3S/EQTsid1jQtewZCEEynR3GyuUfHcMU1
qzz1TpqK/9c7bswSpr4pa0BCHcNDt6Zrh5S/jh2ANneOJo3/xPSn2MNuHXgq0KNjuddax1UWvp33
Liw1jEKodunk1iwpFUJQibEE3crVjcktcLAW4/+hT+nb5HX9SJoayD2lrIGx5pvKM7E9VaX8A75t
qoPxXc5F8Hm7iBpnuImNFUXxpkAEzeyxcvNev9sjsR1SeolkhoI81+IfhNONX4bfJe9Wpf+4bXT3
AerU4cUTEzRZCI7AHKGFcJ7HTAPqUPOMxIxGjgBAW2m3Wqb9yBVPq+f6gRGdw9LDhC3wcxkXb5hk
v6ftflCNIObAlECv8i6Ap28WqjgD3ARW1YRQa9iGRTooV1SH6qyzb6RM/eWxf76zElSVxVUz7HOW
KwjFHQZ+bvyXvrnId6aURFwvxjImSjwjR/XGThSm2XKjJ17KDaRHCpkJ/qAj0jPtpa2/vPxqxour
fUHIXylPUP8qTrY3a3700TohyHFTrUNSPX71RFGSv5daGG+G6XQJ5ISWRpjSgpZLuGprda/QLrb3
fdAHuLPY8qfaDl+4ametoUvwwp0wzl6FJVvkZTgAhCRnl1k/8VwBqmb2iPUtV7jCCuW2jj0hEN1m
a0yKgqxtoFGfi17TY+bSNXcyZv1cDheBHtJsrU2lvnZDg3AkmspF4ff9R6coutlrET/Sv7PNOrEQ
L6tVla+WdeMsQZD4M5Vl2QGsPrnPtCQOZmyX6qwXDh1ox4u5U8loEl7pc/T98TCuWcBP38YNeS/V
pysFLAV/KKMG19S8N7Nqr+POrEy9V3NBrRAJDTC4Fl+no00A2fr0O6FN9SmaoYbBqFNDc3/gRnO3
1c7mX3jYW1pGoXjtTtfRz54C3RRRPF4snZKZ0taqZ3e4Ht9+G6NgCpOiayo80H2I10Vu0n3KkYg9
yezfvbrRfgWfmRdpgZl+v9fi3pMjVVRVwNSLPvOJ21oiVOhE3JVqxUDibk4PZJ8hKYR9Kc7K/EeL
lfdm1RCdLSvP8Zl6dymsd0LJHqtVG4WOTYbH1C68n4nGyfIrrJ5i3DF/bRaqh0k+Biy2UVGEdO3W
LRMA6OxMHiKw8BHJ9KsaVJUlx+DVWXxqj3TBLIxM/etia5C6CgJSOjod0CVxi7Fwf00XMrX7vm4L
bwXwWnTz1cuS/+lhw5tUoOXkxj1mSZaKdUvJ4YuTRotThOMZD49hLAg/9NfAOIjHX3syQoU8XJtn
AudQ3sZcQELqSPO+V51wF52ZRhN3hy/m28nzARQcJBhUhP8kMr1dt3bTqZAUsx5UNZVx7Aw+hZjU
nOaBNb8d8kYjBfC7C2YownMBAmWeJbmE4+gcvZFCJnK8OUgpmjM5Gep0UfBS+cCRhFeqhZZfox+T
XpAGn84N6AXtDLQ8UF7jv/2JZkGB6PitH1Pkia1JKb7ugTEIhPC5BGf4aDKcBadgGtctugEQxR9G
2AIuu5Nad5ZlBKEC7NY2t9XCP9/p5rbroeNefmmUiqntjw6nG8my074K5onwlWxZGuB59baktfUg
fB2ZYiZJZqoWc0l45R50aiiS/DWsVRNVVuoDT9OLp8sAnqj5rjcpkXLcmgDdq3RSjm/uWUsBhQuT
MrKwIXu6e/kJQJbMot5nUuTbKADBsP3lnoXmJ4sNUEtZPUFLV2klrfjAdN1VOOF66kCOy/5B5Vcn
E+zlAGrryLfVwucFZswo4X5TqEQjkHo0+vbF5LYMOV7MohBTtN6k4k3TOVcu5jjpMT2NoukNtqut
OwKKF3365pcr/2lLo8NPrStFTCa3+YtkrFuve2x502csi+JABy0SKXX4rnhI1dNk7McaM4KGvkaL
c44H3u9esuYnvgZQKtRT3QXY3GtZpqIufCLKpwIr6iUsKn3nMbwmSNxziQn4FIvmVI3MUBCxIS/x
DwYve/XfeNz3bwUXUui8MWP9dKA/vezNNvGaRyLnupJsJrKI7HMUElPuF9igoWpyJpAp8Nv93exV
HjLNwwmRJPSCr7WzTw89sXAsYivr3rbtKzmLM/MLcDbWsSHsotqCGzvZfApKzNimCWww/nFSrds8
RyY20yODugDRo8QtLSu4sEnuogtcaeQE5ILg52N3bsjZvDvsDDc+KsPq5RcuYn17hkQhF7lgmYbJ
l/4RZ8m8KVCjJ4G5hdFRV9fEHrjayv250V5LXPJQvnkuvwZG+R842DDTQgWl9Avq6iqga2y66bUC
utX/zexDtR+6y/yXGdU4M2Lxcijvx43Z70x2qHzsRrz9uyDFJI8yZ2BRRioFaPDJ6tHsTVE3FQ9S
pHi1MKiMdqSc4aXx5+n6B4DNSFgWGYIR00+TrECIe6Z3IRN8ZXkVquFBYiHL5nqbEj7+tkgdIiXQ
iCWmy5N530p+aFy/+CY12ekPlPIGYES6KEFkFnaad1b2OpjPaf4q5ClYDEnGJNfLYNKuGkriZngQ
7/UZY5fObeLcHulJeP40U5k1t0u8WPwJwLKxZ8l8rL0Td/DRMq1WBcC8kGIamPIJQT4/+y5lwl93
1VcLPksUFnlUCwXKcBYBqrDOjgcbAXGSC4I3v8BbpdjddVZkfwLlyb9zl1TBxFW1G2iqR6Jma1Jy
dzCsa1rB06UFIzL3Ha0ZNxragikDdM8aQUxcyvlB0MMciY8BAStPIv9ktkam7SoMC0PooFg1vmFm
W9iTcyn3OophWE/Jxd1nntaozto9qVfwh0prhmtkTpomrae+4O6/nsIBs9qQkIauZ5jUGcl2ewJV
K+QKTF5H7CdxAIvk1+ZjWi8mq3nuI6DT8Geb0hdQWTx8R+dG8UTHGOWrQaWb6CfZJO/Q5W3Qmf8z
EvbFXpeLkyonRql1bmQDiOZ6oJ6/IYTdCpYoyI2X5wTe6BrDa8bozDlksRcAuEZI+MDLs23iLI68
NK/4RyYBXFPcudV7dz9T59X97Shn2KKTYMRWyX6HHGnH92h9M+Qn5GZCk566unT4vZUbr9U9OQaY
1ZxdKYJwTBWP7L22Ajbi3mRn3ZoQa/U2eszFy+1VFXoHh0XerW5JMDI/IrktxCgIDjNrUBVBQt4e
GO0YgHtVTzujg8JnwYg2b2B/pNFGXK2GBwtX+/FkKe6/UbY/B9B/Js1zY1/Bf07Lh4eOvZMXlrX6
WKUwSsqPm1DZnsDH4Ta8dJn65KAhEy+dDyoTCwz0t8JJXUvtWciNmMCJ2223nxvf2MG38YruWDrr
hhR0XcBg64vknFvGJgdGWzW/a2l3WMilCHTCceNvMWsPESVU4dCb40Lt1HO6hlN1PlXt9Ip+jZeX
4FJSuPsKFktEVMqGvclQrasSaMPLHugvcMp9ny5SUfZWH4ZavEuMSpipRFzgCewtrHWEeTFYNkt8
8BLoshFjyPCPd+vvjk+XIsWA+yoVf35ZXuKHyZ9rHMRQH57VGe3dfsv0eIGvb5LjgPt/pPJGtU9f
vjvaMnoLcEkDa/4s7blD5zlLylCaNL1ZN8sIrHyCsF1s2YMnmhmBl5aZ3kc506yKkG9BhqO2Rl0r
wbnc7VXRekngj8ZJItMR2gY3ebwZaac5/egwwDPMdrSNcgUZ9aeuFKx9LleUUl4aVfLYywgbtWy+
QOAd/99lFKBsHusr8zkT6zTs1edoQcTUQ1EAOvX0tjTDHoLsKRuGsc9DRj8qmvyyYCtf8ac1rO3I
YrDSTFFiz0tXb7H2St51xd6jY9z4/oDkTTyQGytxv4E4qirdVshbsVSJCxK2w+PSyuyFkA1JH5LE
tT4RPIlEQD1dyNt3jsfz+c62v9y+HbfdlLMm6Dz8nD5plYwLzqZPXEkW8M3L0nGvtjK9fGpupJt7
QDvEAlt8qyWvfyPEv18qEwp007gsuTC93kZ5onsEi9/M5DFUAgYjhkTSLfUsigNHsWnIuTK8kT6l
95tggghzyXYjOUNVANnGnsX/zIlcwUu0fWH6lXC+n0Q0EnXyAMvcdyhiCSZA5P4/NFCacxpF2p+q
5zNxc09lCkCcQZGriTXfmGJj/IqStsHOhEGCbfSihOsRbhZkMCzr7qzBh1dhhDLOKS7WHI7//GOD
MhfX9/YXR7QKVnS3rMsfXsQRVU9cgqEPrhqP7bXTPsTXF/NtxKwlWQAEioYSL65syoCImsw++7yb
GSddRHLU1To0eaEGuqTk4htJ3iduHvIEzoaALii8L/2FD91VMXV9QshtC3NPT7wxEzlWFUMF28jR
Fke6E4lPO73bI9Zo5jSejvdLvKAIoH+07gU2B4yfNn6SWF5fL28TMBmzokyjqGXNDREQagJDBA1U
T9v9DFO8B8hoKVWc1KTe1Z1zyNprnEFL1XflwPrjWxQ0QZcbRhXc1Lp938RT4bSPvF9oznRpuu75
oT6i5bnK+kPhsiIYoR57Zo8LtDGd9dJ3wFTCYrmM7rQgDDQ8laWm4UlHlMGnQFBOS8crevp0wefo
FwvD3IKGUl9KeMF4xO3hYs8bDwfgpSWi3uJe8yrz7B5bo9YEjh/JPSGomjYd5aRJteNG5iHfmuOx
prCtDGeU+cutJNLjEVlHc1MDSuhJMeM0muhUWdjPx3Xj8Sk7u1YLcP0owc0EcMkZLsmPWAxf20A1
Acg6mKg+kFutuwGmGjSkIZpyJLvsvOerUBDmCiix+SkOLmOtMUplmFvTM+ZTXNAyJbxZnFAkcZnu
fBaCspo/q54bYfuwvrz0sNEqHatjD/b7DPCJuDmS9tDSJQI/Ox0AT6zz3ErFqSHM1wA9YMxiCoCc
/NxXyvP690+iQtdKBw8naz+I2CaV1YCP9uM32ipiauDoY11HjVr11azOE++EafJggx9aUTpgi0wM
3/w5vLeD508K0Tdx9iUAVoVbLflViMXfIfSoVNadvzggqw+9RE+7g7Z5qil3V17hQdcj3WmSgWRl
CPrGZIY6QgkGHVudunmK5X493LZAdMnXvuuMjagdWkqSxtoWknfxigj2LqZAjrjTmHRFMOYjdhub
cIG/+mAuVJKpKYHGYWyheXzjbyV1+mT8CYyvGYRVubhNx6dxx2MTJ1MoUuf9KwudONtDpk6QXYBr
lA6q8IsKZXHE7/OeEoioe+Df+alIzrz0t89/pvrIKZ6HZug8RSDIeWen1reW0Dx/p5pRajcBcYYe
nIqJzkQJ17wVXXrbF4MhytWZ0tUdTCd2B6C0+RWXqWPyDs8xxrd/T4nHAMkFlXjYb1S4o06ANSpE
TnYqmqKEfVd63VV1hmfwIWq0BZa8joip0P+JFiTVM1m4bqxeBCdJn5mzOMcrxaZPiny958CusC2Y
+wKIp0ReJZUOlKQXA2WgaL8SivjsBV1qQjebLVyXdU9D/5fmL2B3qrdIB62jO437lNzBNNKaJeyd
8WxPeSe3r7AAZcKQKpdXmqyf2djA+HldTryMJ0bNREP6SfoDhHQBCAbCG3GNzTTavT3Vg5Vd71AW
vMHaiOwGR9gnn8O+bJH/tOFCDs/jajvQye7pfGdhyk6vdwDW53lS4PlTIg8dDsm9pGDSGBKGn5X2
E87wlREmKHznzNn2i92fLp+DmAcrNtSkAV+vXTzoTwpVr4ThxIYnyePN0wvo9Mpd5Fah9ZVajL5G
v3pDD4g20ez8cnri9E4mdB5UryX5Tm2YFBB6bdVL1MTDcB0652xm6bfCXgAu+epH3fDYF9YqhqW6
D+VJAc6va+ycIsUhY3KYhZ59eBd+ghEgo8oGs7Beza8B/Yk9SNR7XBLSbvglSuPJU0pIR6Gf7pA1
7BS+HMOd/3gkIMhbnoye4Mq7v31Qp1xXOtMyCluArIDxc1IazWnnZFnmcTUOUuIRgb3esXd91rw9
HFvYvQfebm6i8gFqwRL3loknI1jO+zyXDUC9bFJ9jthf8ltfw8H3Q9Z+E1SPE0ZZhW9INbsj7EkP
plWBM1Iw0ov9SAgrdGO+HAl/wFwebLPSAHYVWuCQtEZ5ni5n2RFXL1RjdadJI2JufD6OOcbcAL6K
1NxILyPxqLQSLWuVFokkuQU/jHGB6HpCXE7o/10/rQnMUri/nNf4kP1FSfTU7376LNOwCftdbVdW
rLrph4RjlUj/6y3Fm48IXF4+I2BEuHXHEy5Uc+TJfyz1OlP3KnBLYluSbrwNsKZDL6P52KYEzZqO
Ip2WsocvqXQxUlum6FNatBjQ5pLI0qLCQrxr8ErI6DbKvfmI/a5DhQ9xu5jCuKs8rv8gkqbOvI7m
x2HyDIzI4zAncTs/jqtz78r3STfEcIIDmyvHGgTWPwKEQCsIfwyKuCfWmv9A9KRJEf8feDSoFgrK
2Brn6mrCIgAJS7tYR0Z6+wVX4c0ICTNzwq25pxtHR+p09SDzZkWxrofYu9kYDs5M9BIAlO5y9BCB
26b2/gMk6Sl1z+dVxunoMuc7Vd8oNOWOf5VQcY3mGY51keF3p6CVKTsG3TR1QhaMn/FtU32W7M9F
1FdCdDCcKws2I8iAafbf547t5vBHeURGfhaz4FRxpeLcHTwleh2CIPM7PY30xnY5qtHsJFtmMA+5
h/NJHgwSimcU5a3v1pH1WNYp8FLzkz3LxZwP+6KWNV4sw+67cL1Ex230bJRhHCE9N7wVzVp+8bFs
OmAcf83q6jsCxvVSgDMkHqO5ZG/xUG2M1Ljc6C2vrtvOUu3XKO+vU2whX6bhedAO9dhm9ZeL4/85
x7VTMzk0M06Rtyc5R1ud1TshDrhNzO38wl8dw+5og/0oOT6EM/Ay+ZerEJ4O0AciBS24dnNHWMEa
CZd6vI7U4jmmPQt6Is5raKT48ZKUJlIn0AAsPkVUuYIt5FGQ54UbVE6+SxLm8Wo17vWeI3YGh4yx
rPhTFIlZHNMCwBEhcCWA/LmFxRTwA8TxLk4pZIPmkXz0n4lbW926W0g9hAvgjljVmjwmxKYDUsQv
Ro2gOuK41CUom3dCai6ftMTAgVRyNjPiHSjsI/YktmamqM34rNBPW3mLCAewQ0UVY1+RkPc2Gw8B
xA334rBTsLGxsaW2ZNBjzY5QM120raT1/Y2jiZsBo26G0v6H/dtz31RgSANqE9hroBYQeqQLiNFD
4JCtrKqQJZvcuZFpbpTS980aXS9q3abpnqJcFjWDpDE8kNhDjDWFFVXharJpFwZLqhUtXHA2Zibx
zNu99JX42Cnq5rJPl71PMdQjEQObBb/cUYVONTWVrBC69i0HgN0zjoRYdmuoH3idGnl9BT1YEKZq
dV4M2LubftHT6w75cjsuyhyb3zU3QvqF8rOhT5fV4D9DSzZwytAiQTIvIJOr/RFB7HH7iU6DDVGA
1ydWD6SStWV17GTuP9DbF8azvjllYF97v1Yw6JDbWfr8pHGuWrEbaYsLSYpUFIwp71OI2l5EFpc3
WGSbMcTgH9AA/jAm910s3uFAPY27ZK0Bn8pTgcGZQNnJNA84KwX1ix1xcMqB1XociTMv8lPVtqDB
2SrZJ6o04K++gJAhoJ4ma9tsmGOCzNWuzdwd+5/SmEeB2ZI9nXy9iN1HP025BVHm3lMaF5SrhVVl
FjiMM8fRCO0gnRK+dix/mJgrYgFu5ArRLT88q3FP5ReGBjyUPNMRk72rmZxtVnzYC91n+Ex1l7TX
kqwTSZQ7rEqwPi1LoZkXrMG4xKCAOHTdnHoV2zdbgLF6pkw/nwgWzIRhPeFn1TqLcvaw1LN7OqwY
IwMK/zsf4e2tQc46oHfi5myWsQKyEc1Zx95MdyhkiGGQJiZpOVnhTedHaamoJyvIC/lyMYmAfDZz
Tmkq+h2Y1q1tEs7TBTX0hKx5kuVlZdyA/cNY/dcx+fCanYsCkzSFzOO+LEeA8cFQPupmh93FrvTq
I+uNwM96MDwTjyFC8fajhLS3SoP9PIPRkspqqw/gHvMsIgu9JhLm1o0qLPVkYvXzPopaUIyjuHI2
bRGf1p1Q6WEbaCr+GrJcdOaqvo5zYFLVaHYNh8dUCKHD4Vh9/GXa7Bxdj0ilFLx77WDqcKV9yE81
4LVJIMOuyGRI5svOwiH7ebmo5NOIoSx5wQKDRVTNJy6oIoAIGCb4BN61FQlnGB8uAk7k0RT+GK61
j4VgfnKga3H+drs2GgulihsloC9bSdQup7kDw7jGqnWXiMN/Ojf3veULzmjzaiYAWATFpcp1Qhkz
6JIUtGvmipN9U61FavzJiseKciLpvSnv4DViQwuUTzeMxUDeyLlxcC7jC5B+5331nCT6PSY9UX6y
rEc6h4MZJv/GkJkKTWqrrbNNCnpRuk8ongbTXtWTyWYZtF+1VN6kEi29pHCMciosCMW4N8UyePpQ
fjE6iknWxBheTAfZ3zs4IbiqEEi4Wt0vevlAlXgJIXc7bkP85VwnKCpTghIznME1brm9ANzb0Cq9
H5LG2OBdzF0Srite/TC4uocvXDZ3Ydc+zLuvx8NnWXSgIKnhFiaAE5Ak/ZdGEp+PMSZBplvYjVx7
1wdn0HMXTJdcC0Id5DA/mVo76pjKoYjf76f//cnaY1aAuu5dxFLx7zVcTx5YjFuCgryMybqyqOS0
ODvKix6WWZZ1eNcXzU4h36oXWztlnvrQZMhTQL95YU0XTxuHTdfFSM4Mx/gDkSKv2klYhm76NhHl
5yYs0P17CDYH8XixA4c5udl17KiogPAWoPqFBopxa213rj3jXwTLIRg1lBykHo7h3HbOoLQSpoXi
d8vGqhmHaGmCQp3VOfCkWsIa318EZnH4iTxK3aQ2UAEjz1+lSD6/KmwsMP6afYJYWM56j0vlQlR0
edDW6qjcPp8Ca7TFZOXTuWyfEgxnHyqwIWBZOFKB9OJhTfSY0fPFZ6lQSmxoy7oUMVDZwCymGa5h
D22nBmcDaVJEVtFAPMyc9c9G7Rq+YBKh4ontg80ley45Mn1wpN31C4LBbBUPCEyRu2A5gyy+nz/R
MOsCC0W24naIfXvgVkKpu83AZNBxXvHePWyyMPLmlY/fVwi33J+nijAhpIH1+0maZXAZIgFxku9z
w3PuWLP6+lFO6bOLB8fA1gfAoP6YMdv2hyjyxlX0SGpOqdRRcADV2z5y3zQBMujWhNcvxAaT7O4t
QnDzRbXJLwtub8sJF+AcrZKLELbgoFot2S88sEGPOeVgxHPaWyJnVHS0foWz9QOaUDecQZc4CSEH
j9+3/s3MqPR6u3iB/sbJmFtnijfv06Jg7+mq01MYEYguuo0YQXxNu65CnA7R2UPgpQlFZUQBBYFM
QY4zt/BtcP42X+O1VRbx1B+TPchBooHr0O2yKQi7JXRv+xbMgAeJ6LoNi84nxzKktFA9kW+K43Hl
MIH3tXGI3F+3anFAhB1IFW3nj+KtlGLEcbtzsJTyn3feObDjc8Q9g+QxQdQkZwCGSweZQyGbzT58
9dFolSJtHCR+uln+II+XeVK8poUW6BIvzv7ZCVxhk1gv3jkzHNMMr86jL28T2tefHi6aNkskcY3R
KyBvdsUWrxl+oPDxFpIaE6bjBtAbTioltkYOSyfHzC0RByRuXIn13rE/Jy+f1D+2d2U1sQ1bMaLS
UHid1YVkRgiHX9o5+bbDHJHWnxUYm0tnjeDLy4GJR1eFvo/TetcMJI+U1CwE83xYvLNSkRYEBRq7
LIY6dhvQFuptAhhx5KHiaOX77v8pAOo3z1xihH2OoWnFofBzu4Attga5lzvb+ipaINeLJSgr3jGO
ZdGwgnuhFXwV5kohNRhQVIAKuvEW9Tkz0/oO3PGwscaca3ZcwW60dOPw3DKkDzne8+brsP8cf/kd
V36V75XRlsvSdYl+aPwYsgozcPzRdSNUEPqVPM1WLXwteTzf2KJfT4/bWMO/9FMsKD5NoZCPXIg1
j6b6iQ+TG+kzGXvSAIQjtMuBHnDSBYaafXTiwtqsE91ZQPDYo05SpcHokBTQNmHrakwVxyDW2h22
/BIgIBLe/8piq+UA0eMX+3gAZSFbkrMpo43Y9L+yCFWp6VyGmCFK3CRdCcI9oe7SpsbudN0x5jKx
Q5P/03/6aWrFkmhG4y+iSA5jH2cA83Dp0DLHuS7Db/nBskh95RRUNvRn8f7NCXH7TBkuXykeHFkt
FjBeCiwrDPNsSQdBhRRfdCF0E9EkXoJf9JYZEdmdpPxuW4ogPGSjjsHsPYMhkEIuaEx3VHZdTpax
rPwPBe42rJ2AhAI/WdVBYL9DGev4AiNJGNr8VhoUQYgKWr1yD+Z+oHj+anfhOUkW2KR3Ldh8GcB+
QOgDknELOhH9H6fT4aOyKxITwHMUH4tEXokU7YDRc16bGGHIce1q9l0cJ/ISDaZTW4hk8Idh+jBs
OEjlyhuocaDpmrEARnjVUwfeIT6VKOnN0BFKlEGCKRxODeIWpZjClY3kDGATdBJj9J7Ur/7VZoHf
cyr3dtpSnn1afhQhW4jJIhnWenXgG5QHEJQpY//rGqz9AEmuvC6OOSchR2bt6eCDDZYSw7YlciQw
jPENyl41bkZwm7NVuOyFM/Cjz7WyTSs+0yUVSF+JUFntbwfuTqVdDBYFy33BUqFeQsVm7ZNxtpSQ
mNPIMzDsFzntYBrlCa+XG+HgZZsd+GhFk7CEWOGBxeN6iopjX6h7lC4LAyaSioEBwRfSA0uW9wbS
HZsp9frAh1CnMgh/kx8/GBo43bL3x6f++EjfuThYzYPXyCQq1FvWlHcsSIELlGWwoPnILO9+Gk72
01jhYr7Ojb0Y34Ev7FfC6oDlKL0fNdN96s9OrEl2XAzxRP0mkFxk5r6vp1RaOvVTaM7Gj9QLOyr/
gAM2jcFEsAKyIXCIn2RKkwtlG+ipxdgyCsafDgYQ+6ml7EGVshghgexaN9ahpTmpZ8EY2c3+U4W6
lBMBTzpRgBq5It3k4inMsME3Q180HaADSrHTATNvATEmI4aYyxvZuR/eV3rQ/7JR/M1c4GPMmV7h
En2ZQWqGOWIAxZ5j5BBPrf6IZM6KD9fZINdbcJqMUC6CqmPMzTo8JKCEGIk4Eg4yeDIyci7V6Ysr
a8xUmfH/kUsAYAthznivWL/Ty6tC5HGFYkOKfiRKvW2HiVoTU+G4jSH8iAluq4Q06lNelfUC6eLP
QxB2GrCF07Zjvh72rQrAct022SMvCLwV77R+5p2Nb//qnGiVlGoNAXZ22aliGRFsI7/yQmTwug/W
vvLpJDMWifXQ2yMRQwfV22xgFuil4usnWDTxE57RlWKvlw0VNyrNoYVqpI4shkKpypAmW4nudHoI
LkrS9L7kKTnj1jeWk6oQMiSDnTVDoW98537736ursDMvLY8lavuuBhdAo3vMYy9CAOVPFAYRwvnb
N57YHbL5rwBFUVsXOg4ZsQ7zMAH88WI4/F/ypStbqpfYnak0+pI21zeQcbhrkVhNtauZoNqadffL
kI1Kv9lmArA+YkoX2wefUFcmtB12R8DAWH40JGMcJBxxLgKKiss9RUIKH4q05VjV8laVGiS028Gy
1z3u9FBdLPgnNkhlo1Z4g2JS//GK3xKqBFq9GVi1q8PzC72NrmucjGwLN2t7gY/bYuMo42iSUsb1
NJVvOKJn/ZNko+EXfJuEeFQo0IiUXK9PfL2QBJ6hTT9Vph1HNBbW6rU/78VfvWcFWa3+UZNT1FsQ
/minQz83WJs6vMRDXrgUDY0Or0mpI8vM81O2661bNaxWpG0Q2OOltQ3dRfE22HmjvsOEUhJjZbug
vUKQQLcZ9wFEQKaZf7c0wkmEhufAWBaViNH/ilzkeTJENNXjRgZ/XYfQdNtlE7kqJlMUMZZ+1sEv
TToAfqNLgczARM7ZsZXjBjiHMEeQ0Z6c5fo2Sou0vqhNw++nmH7JYhxeGDjFLXO6yga6B7TmUygc
LNaaU7ZJv3X9+E2CyXGWcmNNgBVs8pj4oLp+h2p9KkNzMa7i2hG+EEGITt52agmGIvurpCK9kYeY
1A1TId8dkBmKiRU1ZL33kinmh8ShSYN6uYyCwKMzipQHSmfWk9tOMpsq/elmgS0PQBkQs5vF1RhU
1qkcoZv1v1XPFi7VWaApIGfMy0xFEcWAwyOhYAeXQTpWIo4Hc+/uMa3YUoZJUpj2i/a9jWtR61Hc
rQq7XJ9xshfUwoUjUvEmYYw9y4sDDdyqOtSvIlyXJBOTIdiZ4sJkTGT/9P868mMtZ2DyDLuyRucm
emzygMYWVra4ai/+nsIvUR2yxNbgUV3sBSShJevSrSnmw8Yu3B4FV047B/F23ipbmEQJ9ZssXkk3
H94oftvl8OgA4ekxs467niqHToOk6Y8j0U0D8XfMnrHzFLEuggm4d2fMZP4tG6n9odflboD+yKiS
AsNV/zsgVvQCPQgX9muD5DqDBxrhObal1bRC80cCWAZzFPiXeprJ8tkwvzs6TccLwqWTavIxx7ii
w+VRTZvnyoXLtKr+xzzmPg3yX4wVZcuKQMQhHB/qnS/Rk+OVNdomly57v2me2HvMGsbf+PjqedNI
rUPj1gTpZmhEPXuFK+Tl8MLpKHdw95KOASmBRBi9tYfnvRgxAmPgbgSpbbzKDLm1pI/ozh0NLaJR
0ofiu62zPOkSLDiXD2t7O+VNcwIs1ZqWRSMKptc9UQIR2pIsDJVI/KMr70PLGqMNfsFUEXFL9fGd
hxDVBFRu+QO8wpXJB0rNZmkE3T5/RqRNolaqy3iP3m1X45MKzViHkXTZo9NMzqEL0/M8FgDXPzwG
WwniHjBNLvDzTfAsZpW2Ag3KHwO0tRqj7PwtoCMZGY4swv3gKBObgnRaVUVZcPfG1ifvMB6GdUvN
7zJlF/H6oWSVXu1h2eWSpUn1S4Sh7Av+r5kNohfgDa78zD/BHw1gjylFGHRF3DhFCvGkH1gxKt0t
zY+r8NP13yQzzynTApJcSxvp/bLD8y363obPS7nNk6EnigbzaBBxExJPjU/OlrKNyaf+tLRlPIvC
a5obYxtw1GsWCfNWUTE3aabcw59tpqaRErypwHMBjC0Dl2dFbUiGdjfbsdtzSq1Y2vZPdHSlqOj5
jCWDaRbnmC+XRqSHijcnJpzfPGeg9VDbSA+nVqihR4n6JBYS0pxL15CCPhD6UgjTfR1V/B984io5
TSU/4F8faVdBjBUKp4rCZj6QypWi5pmDNxFIpDHmEKEviFMpvUScZirGF1j7ND3G2dMRUvK7vg+p
yR2AXgbe/+tDSiDOwvGhDub51qfem07ZkQLiuZA7zKtg34ak0PhZTllp9XgVr4nFh0cwu3OeM/CH
tTbH99Jufv5/S+XkTkntJ+OPU3uNMLXvSGhvTVioLs1tX2V38p6Rzj8n6tTnlC6kZA9gfz+kAkEi
OWNP7wccptA7ZgaRGqUlQmdG09RGF9XnT2rjF5DxWe1IvJppSKr0luD5TTtsMvRGBzlM6wmCwetH
H3aqLZXogExUHqbVvxSzrrEW5NwKMXaciQWO/s0El4GjfxXQ+mGByFXJ/Co++V3/bqlumyYNYCyq
9Bwp/vDlfpxGn8T+G0EJyPPVwsS6MyCJGh9sTj8zbJiuKBHHAouZt7BZQv9nOY8VdgH28zlrJNwM
8hdjFqQZCnOA8w2R2idlsUxNQrbxS3yujiMroGCH6lEQYRSjygCQgtlGLlSL0HfzYBuAM7AYD46k
aYT0FdwYxpGipZWMf6/V5Mp/3d9y2Bq1AkhO3Lwc2djFsWBNP0zO/KxSiET1XTQwlYvhCKWcO6cb
iXmd86m8Dh6ACzxRYlivwg6Xbyt9ydc/PDnz2IEJvmuDFxZV4t67Du/0EE9D2vvHYpfVrrabqMfL
tdmgzK35sNKKh/2SxRkE5Bf5AuveuT+cqm48h2wAs3aeF4FXk+BD8AXI+beJLOM7fonYoTYRuV+J
OznYU4Ma15oQUSvh9VMBcBtDhT1uyLb0+9xKJum95T3nYRsGJSbnl+6vSgjXMnWGcJ3uhfdXkkb0
y/KNIEMbJwLS+euLhsZf4KKOeOf+AkJFsrPh+vVBSS2Yx7AqEWndg0Wv6td6zrJYqAWdtZX3SSG0
qD/bM2XyYx7ANFGIWSNxf6ZjKH524R+i+92WrxHICtRj2pJcKf4yo4sb5/gz5JmchRAr4Nh8ClSm
90dEmaTgX1Yy7FjSloz+0dJ11PybmvXpFGfl8LUYiHw9u0NXTuOgMS+9xTxxSXVVdrSryNa4I46t
DLiL5B3GFZPEL882MXZ8At36CkZ7P6qUE8BcRt7UHzwZBSoTIvLWaDNq4hRWu491EskjMn2YEvI5
8nx3RuqLfZisRg87JTyTwl6nNlYtWq4su6g0A43HnEmCcFp+54jHqXooDk7FJkhrcoLXE/QtpDnQ
Xai0yqR3qyj9Ibr0EC2UaK1HE4XWzf3grPy0fA/F2ZRaJ1taOiRmBGg8gGnZfbbqXkSuWsZCESOR
rokFxtFC7FlhkYmQUsLtUzlx7uZ0ZE51LphdbFIi66x9ib4iQ1b31rQIKvWdZ/qvGqEvLWkTvbgB
2gUi2wMqqA/TDSwa7OasGSqu0fbhx7MRxAM/kJwyQ2bLSyVteIECUs65JRciBE447wGFgesLbBv5
118f6VeYBtJITZjfTtxraJb9dL5CpQF448PeAuo2sSGAJVtxjg3lEFRibXcKD/kzLkkbzRvI8twI
cq88mIH7qKVyNiWKHBLVsOlxp6GOqZczNM3Z1B0ljMKJf3Jh157E2DQYDbHcH/uockw32/JcIiYO
KKeROExWLYqh4A4Cg2DR5V3ZxrhYPq/ekKdY5aMZnkV0+KnIyNDIvQJBmY4qvKtp77wTbDSE9XVq
Fuxy0lUJ9n72Da15f1DNmmbkt1YooEUOyHOubBvy99CGQeezoOJCRnRuwK79aNCb5ti6IDJvmqwF
kE/a22TqLM0e619W1qnxMFiXbff3BI6KaEpSlc6PefY4XkKPlLiCVKvXV3eQMMslptI0Rsd6cTwT
YR8YyqzG40+AUp6xoPSXaFrKCubT2HhKQ+taTyaI40qvmzqOPg2bmKo3kaH5kjVM+jgtHEOh4mEQ
7Yv0y5PPjkATgLjY/lrVwbrAs5yVoRWhKrptCJD5MAviRLcWDFSRib6Pjn4UXrhsGdIAAn+s6J0G
Wa9Js4COHGX2hE/VBhQ4Gb2W2JTKSeCSiYecLres4blrIJ4v/49UHCPLSKX2gkV/qG9utLKGaNHr
drCpopyHhtarHoPKOMoPn+kY6jxMujj7bR5N66BhEvrJisbCUz+EqyTOvYngANpaIorWxOzxZMfI
4W0+fdH4hcXaQf+aIypcU33Gj89tOvp0Awl2q4yCK6K/kyO6WXGuPZqpk4YUagh1GDEseb31/QZM
pZM3lpMfQjcb1jqGyPGgEGKn+KlWFv378qaPyJyIzpHtEQclqL/iSk+4OHMG0cmoP9lmKQpileZA
BqlzZATKINC9sYp9bbQywMZ9Kv0af2/dyHfAyxhRTiwFRzPxWYWRsyqWLLH6F08WLFQcLsOI5/29
ARpGZL8/ZC22AAH4IIoA9zV8PuHYUM4T1WFBqpOOvVChbm7zyOVlB9GEhfUbgDERdo0K9+NRTu8W
aKVXFhET+hG9h6WK9X+3zGjKuuDxdpIm0XyQqTpUrLE7e2ffptFSVJfmRu0OlKMKsBPMHzj4MZpS
DIKPIfnhyffmm4dKoFhwU95sYUOtHpu6m4xMABwgLCyLjIvO4Iifbi/kiJYGAOTEZT3RT5qJIW4V
YwRobN4v2Vl52TFAEMPmJzjdBoV/tmV3vQHhfYliuHiQetiWh5ucdzkx0dAyoOKtpD7IyJAFluU+
RS3lsVZcnK9OfNOVrmQKNjesn+0rtD1hcoxZ/5j+YGRhTPpxfrsBfugHh+KHwoylwOXnAxqS/ny2
VDhjdTNs4JKawXApIRl8f+c+h79/2mUo/wmMMFnUqaHMztAxi7D4KVlZgRfaa4Oi4GAS5HGScrw2
emzB0WrQevd/kp1uMdHnAQSgKXVPQ5Xo8nIWfbQMt1AdD+KXFJC+4O/RT8/A4G47mIOIF8yzJhDK
/hAKOMG9bLQFV8vIxNMSP7O78wcZWcPfsg3d4DT7cS7MPwGmSYHgYCvqBgXcJOrUtoBjU13WE6DF
gJodUbPB2ZJnRymPM9nFkoqmmURRt1ce+wIga9PyAF9IPqwlJmi5T6qHjAXfQZCIrnE4r/IDho7s
NSBplnaQ3PiAKZqrsACPa8sPwuZTbzk98vWZqru+Iqv6AA==
`protect end_protected
