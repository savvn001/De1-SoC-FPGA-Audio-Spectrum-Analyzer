��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	R8��&`XA����f"�T�H�"�N�i
`��)ztb���Q��gG��E,l݉ �6f5t�0I'͡s�uX�� �i�ď��MH��R��Z������\��ă��!a�V[/Y��v`�K����Q?&J�5<��L�k��.�Jn�x���x�I�����Y��n�7���ՙ#���БD��L8߹ᓞ�lC|6'
J�3�P�A�\-���&��݈�_�E���j�P�8�_�7J��L˖a�o��y���[�]�FD�N�f�)e��ǅ#�D���c��]�����l�Ԥ`נ_%�Si���K�Sy����,�X�<L?w���:M̠;�,�Lއ�"NeA&��ΐa� pQ�	����(FT����ڨu��dR��|���Y���wHsy��$ts�GD�c���秙!
��x��O��9����'���A���Y��[������&ǰ�/<B�M�ol9(�'' ƅ &c�ܷ�c{�F�ƴ�`�������s��:z/�L��!��~��@
���7���ȗ8�IŻ���ҕ�����4�U������R)����CɆ�%� �����D�ǔk�S\鰴c�~'�N�k:/����;�ET}&QΐS�Q��H8	a�k쏊�)*�d�¤�)a�V������×|f�)�=�"b���xEy*@c1am��EnL��ZV3̴@�L���hD���[�կcC�bF��"���v^�����>�� ���-#`��f	�,��˩��I��Z���[>��^�I�.'3������D)9�+�F!�%�#x���	_�gJ���bq�Z�
V6c{�I�m|� ��T����G��!�n�0$oxB/�Y�LB7���!~ 0}�-�2l��� ��L����op�t����Ce�^�:�:Ԧ�}����o�c�=<Ϯ:��h�[����H8��
����Eʱ^$=���C�g��w{�l�:1�<V�QP&kK<�I��Ԡ���_��GsoEb��	�zt6ހ(�y?�y�R]�+WT�A�;���s�C)ƻ5ϛ���g�I���Us�!"';��̉|5�ۏ�H�)V���t���U8���ke)��}Įٹd�W�y(1�;C�4���ǨG�EY�xӸ�ClϏV��f	YԂ �KP:�0&���@�8m�>�E�*V���;_�~�n�t:Ǧ�n���k��X�H�I�5@n���tD�*d~���$�=�e��1�P`R��\0��4