-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RLuh0mNovHv3vOnQclKC/l+OAE6EfSK1S6u+yYZH3K8Y72UATMEE2U03o1pR76A9fu+DJ1bWDcSa
gCudB0O/yvRP77KnZri6ap6DxHu3umgsGTK5QbgeP2NBkctwcWGTVdDlTy1DVOgn4VgCPCHYpV6e
IILOAIFVQ2nWXZF8ahb9+zv/W7uSXAe6KlikRDdZUxIXxvMke0O1EYx2cxmvJdJpP9wOpHE0fdpC
2h6Zf9gihhcN80tSXpharaBVIOMCxxu9W7l+VmXp+GPcutiz/rwigE82Bh963cKJkxyotNhJgR6f
jNnKbrjw0D1sjDYCZ3zIUcrRnkNt6rjzoT/WUw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
jIfYt0VqK+IthpYYR+21YD+jdFSQAQ7WDpGEQ8VfOFcYj85DMZglAmgauw83fkMB/a8M1y0qlayh
tB4/BIwJB6csNWOsMYtKosQg+SQm0L1swEAF+9tUwIPWNqZ/NFv83VtY8x4d3JG9quG1lIuM60Ac
6dKeADEOeh2M4IcLTafvIomC/+r5fmTWGwNpXEoO6UWtt0zuJlqPs6DxPjuTAGAFTE1cpa/m7lox
rfRD/N+AD/GEChOm2Lp8UUf9neBXDTNpJIx77zrGE0F8aORgYqYptb4KqPJ6ke+JF2X3DrXpBjNE
IYrSh9EXcUdjf305iTjUxilvpi8CiMyPP9zwwuz465sihJJXByGfMpsYRaa4+RX8RFsYkNIHpOVd
7rZGoGUzi5BPKxT4MeuRCJql2uSRFjUK/Q0zAIXvQZKK3ad1K9FIHzkJIpWG8xoZ7TPBJdBHsv+M
3hCr6IJnKadv4a7otgEIuerm0iiLtDGE8J1Qg2r7cK4HI+AD06OEFQpnvaIIKHI5g/fIm/R3K5QV
Coj38SIJK82cGtjqznI3T1H73KeXGJF/qbL++lB2cxtDrhj7CRWYA2kNJAVt757e8voDMk1e6Fuw
hLyobT2gRbVsuNZcDIzcu1K3xSZ7XH+w0a8nv1PvK8VPOE00trmRwHlfHZ5cIJWpsXwXT0N1a9iR
KVFRWuOBfVhuMnOlezICthekfAshqZP2MmCcdmubqcN1iZFr1Jnp7lbx+IIuJX1Na15mhrjUYa9q
thK92mXENzNOO8EAq+rxV7Z2uOXW+LbSi+elvoaCaSKYRKOjEkRtMrESWYTjLL+gKZTcNDv/48J0
ac2M4R99DlaywaziDEKTIfeLH/tFY6XYrkp+XqdZYfe+zFUxazt7b0w8L57iqKUrSM/kVbXTHqjT
5pUb8SS4pD0K7XX5ZKU5gD6sjv+oj+O3fWp0OHpvK4hVySVAilHyvhq81X6MddfWqUHBinSyigQQ
3z8N7gHQ0bQdOEvfw/GkK22vp6X001/Yl71EnsGsSWQHMVc0zHDJn2DSF9rBGKmovKxVN6E3PoUp
PM3gZo3cvGGEmHOVlF37lnEJ4Zhb8GUE/q+squys4q9cmtA6s6gVoWHIvFYVwjPS255iRaMZfG3K
7Fj6hNLaYLsq4v9OvRsEM8yXnAU4rpZorSEFYn0g4U7xnX2DIocdjbVnsM0w+L8No4SJAizJn1Ly
yjkUh315zrrL8z2dQfSqfnJ+xgocGz2uosdePYw3d5/2Mh4D0foyfKv0GMhYm8sfPa2w1xkEWotq
Ax8u3otE6S2SsIT2fOellb3CUMAv33slevEJawLAEx+x1Jq1g5U7KOS3VJtwgqUzuOB6iIJ6nezI
ffnSWytIB8brnnVniirno4u0xZY6sfpT14JZOzRJveQOOIgo3WZbsYontUuJz19EMS8BwJ8cTUcW
w0c4dfXTwNaHOfQsRoQaZtX9uYxx8uhihVTeFIrVr9cOjlG5Cv1RtygQ/tGqQ4F0fNqPiXWYtrXD
0Uh1E4ks1Bs9HNiRoXKURnf2VMeViq8KGMOAfwLOZJ4q5odGVolnhWhgsjbCLihLmb4qD1rZOCPH
4Mqn9EcDK7ZSazhm1HgWiX5eFYojSM1EvUmMlCthXQIG0fusO+cyqzxZzrMst/h66WPNXO3NnM+s
UT6qO5uYWsg7bzchVkcR8ABFzP1MDOs5PKfHt2Ld+h5CCbf80XBo3EIvWRK3wlEkXr+e+ZMTLPrB
tZaCZRVETtHj8TI4rDcknGw3arkrxPFlDqu6BtzirB269TSR4Xcf3NykZwHb7kSHARRN7UOp7DDC
cx8ANTAKrHbupNohoHaTzSD1Kd37LXLOAeFIae2kb2htDDo/G+4j+PTZb7zG1oa2n0tJ02LrJtkN
x3/DWDwV2GDZckpcFRDp65jXupWFKbVOpOpDh19rhtBNt+RItciYVYk6VGkh50BhZzSEhkiHuK7R
OPd836THwfBmQH7jzH1B4bovV0UhwNlRnoCkbUdfH72zMNuWKcEpmxNDVFwlvd6bqNG/6PdenyMW
BEvo83RMRHQoW9stvgtm+54WzlFtjdyQRuckApPjg7uU1zMfckb8AwV4lpWH179xRGFNVD1tpW2V
yZu7qSjsaC9zHSt3pCXv5pYSPDWY6KeTp0wefs2+0nPM23SVYeRlUrq8rPhQOS7RvNkmjZXBiqYJ
khvPHQbrxgmzZIjXfkIdbYeamk+oOB9sISmh4vFeXiUVknpwkQc/YTrPb3SqvIG7y9dyYFgky6fL
G44Q743CtJwHdL5eKWOfD0FKIJtqpRaafHCtGyRxdqSIQV1J6KdPODPBoHfQONiQoWA+z3FR5WXN
6gutVPi3cjmvLkHBX9RfeqS9mbBrJLxp2egsmxImH7EBr+PaBiHp6pK+2I2pinmxMyqj9k4JVDP3
GA2HRzV+qte27yRc69hvvA6yJKP0XaT7poV3vP9GRTeNgxm2tFg70qR/BMCuk+L9Bgc5wQwK1/U3
UFfepyUoMFpJFjADJyBavhFBrSukfH+A0Tst+Q4CkpBsaxUwQQMYNz2HCywI2qGIaVhO9L1IwUEh
AWQZ5JXuS3oU1x26BWqoAeqZnf+WCLom4+uVGkSJ6u+FYE+TrCHK1IE5UwRYufn0oxDzzjblr/tQ
cN6FAx3SwItj+rt0omObG+PMRKNzpEqH2ROOM80BpQiAc19vZz1dnT7YK3HC4wIGSOBRqipEJ5fI
ewdqgLev5vbz1NkajTrTGF2LvkVNP5Q2tJhb4ZfO2WflCs4ZX+ofjK76LFCazYkNYrZQH41dgD80
pMQMUGJQoaqyD4gmMa/Hh3fxHp4+XS3K6DCV8uNf5c/cAsvHxftAjasjQhglKKZx3r/3mSc7oO9r
C14WZ32ReVixJOWnwWphHkWcRsLb4P7PPjZx8zSgS2sZcA6GHYuMthE0nWGnZkP54nMcNK5j2vXE
GHGTUry8kJoplhcDbePnPYOovXtIQClJA0U9TIWG1lsDERtVbLHsuB+JUUz9uY4mdzAXwCgj7t5F
lPINH3WC5udyfsOQFQ0gbmfT/Wc/P4r1RsYOlzIElsWJD6yXsJ5rOtUiCnce1dZw2JRPvRcX6gX6
ik1TRh1xiyBKsAi6jyS3QCGteab7pJqIViVWXEn7z155q7OEfu0PkYPz/yK4If/NjlYfPyltjhXJ
BxW3rxDwAjC1BLr759UDyY78/7Bk16y7mt5bWqjzKX0N1liOYzCHkjaODtLVFEubPp3jgk/BlDWg
3XT2TzYXyp5fkcB7vD+HgekA/ibLU1hm7WZxkhoDXNIB3DA51yUFTcVmfjHmWaHLM2WC26PqNI9K
M7540i0V8l5RNZumMPS8vtNofeHaptiWL0ohPrUArbSHVsqf2mOATuUqjq70vtxG5DZq8dxp+ZnM
5/sfLNk7lNtwKapOufICmNWlEK9YgsRhK8oDlPXC+i+r7nymD3Rx5r2MD4VXZ2OmIWRufusCJfkl
JTB7cys2Wx3PfZRLyr+4gBd/6vNLR12FBTFNfVv/evpRwKG2IUaxVLddgMa9wI6anbZadu67DjIT
ErIbEeI3anuX54ZgAChfwFldW2x2mVspGwa/eB1KnlY07dF8s9pE7iuE0esXSFSGWoITxGcEyjy/
JTmlqcw/eJRwDPhx58k8qNQAswfcyWtqyMH1apjY0TR2B4KXXpY+OGrN/3niFqycjVFa3RtQ9ZVV
oxPsd81brGiOdm730XNeVTkRm5tg3Y2CLmHYF4CVyiJgxwaJqcglCtVaooFrVcooXiaN29CNplYv
P8IT7abF1kM8iGCg/OX+Rjbc2QHCLStLKLfdHmOHd+Nc5FVLIY8Mc0gkzWiL6cq49Tu1dmfn+Q/o
JZe/ts1Fuh3Ts+cQHJuwuhnDi9IcJoJDv611d7LRIqQpWrvGwy7XrOr3HxB5Aaz4NjfN6OL/jSvC
TYNdsSVbMkJIJ7B5B/BLP4ecBC5hKq4z0FTM8UbcUR3YnQ4mVDTbyEmLOFt2l4Q+vid/YtiKT04S
Tl3A+yrcOAvyjPhbvIfFN2IRnm9ykEwvqfvHii1MgQN0xfCirx5wC+bMF3kqoLv1ZrZSQInpOpL8
MjLmiUKQnKpdYPtDNdXCACSmkP2CQFYV8Wu11ooNCE7Xst8nmdcIJVBvm8BqgWzmAEc6iMuegeul
W+bwacF9NwZD8KD5Wiaw4ocElPoaS0puRvkmJCba/uaAjYc+sWnnrQG/FMJLehmnK1xllW3PFRXH
Sxvch4c0zKIY9zh09zh+t3K4jRmAyNggCFK302/RsyPoOGPXUzs2G1rzof5hML2fSTsa+hHpxjjx
G5Tt7nGU2w4cedSUH+X4S5dWN8RoXAIThZbWth8f0OSVD/i3qv9GUUm7YuiNR8x2w+4m36EbvKim
vDWPKgEPGurviZA9a7Q36wBcMJ6gwtsLbdjhLfC9Rm5nF+ZIvIt3wVoP41gYIqs1bB8KQqM42yY+
W7GouZvZhAvLCYJAIWp26r4tPWHQ8gG49FFdkqHeQBD6HouifLUgyoyUTKzWKPKD/zUh6V+pufuh
zZwBjmfOEZViYzpLHBXsMuiok0A+evncTAT+cy/s5K7VZCCPsf3GVyXCGnrtVCODNf2X0gE3qpu0
kgrYVv/BnujDqUdZS/TKxr8eND92/+qpGu0tfomln4v6YX+GK3rT4uWD8oEjxTw7/7sg8+nuLs4E
Y/QdDmGyJ9yjRUqe2POrtupP/f0uhOD/CSqe8y7Ad9Q5pYMkXYAgv0c6t3Yv/G4pQ3Xf7kcA+oen
ZjKnksfOrOUmcSU6vxsf5J1vydQeuHa0ntDVqSkar/sSIr15KdeyUdppa0HgbyrCYWnQJtuL6vaD
Ill+kX4xuBZgRwT3msLfqRumK7l0lhYiP59wtpBDp6GUmqTmdBZp6nan4u3ZTaToR2tbAL7DyliA
vOcvQ1mZ7shdTFoXJPCG1KHTc6eNbPEkrYQe3BHOURGAvR3bYjRwzJL0tZKbLI7sDdxJHAlQIajY
tHi/zZdRznrWNSbDWtVZuqcDxXuOc8vir6RbgALu+iiuojcDTulidMvbO0IombGBfFQcGHeCuBhd
CzvIfDdiRFiP3u4zssRgLEZSEsm7gDoVq+AaLfjdwICcoXPs8vuI/ou+2EbRFQ5dUApkr8xDHTL3
6QIRZ2DJ2FUcBOKTBQFXkTFvpEScnUwQrtr+cgtkffvYPD3b033QozQD/ipLxQ6noyeW11S/kTKp
yD05UUu6YlOsowZHnleYNiKJ5GDVHtxCgNzQ9IrNsTFGaWpdFGSHIvC9j2sWId2zMfAJDzLnuABn
VCHSKslUlhLSLcRYGZd7nK01124YoDkbgoWgmh63rySPz3uE9lHptRRkWChod9TiUowNkNeSpYkI
bX0CWL4nDDRkZ2FK7kOBEdP4OsyCBagmldm44GPrXdiFAb5od+vgGcGxbAgufyAY0eyF4zR1hUik
+PM0Db839Fp/P5EjosSEIaJw2MyLQjXLX/uBmyAxJnvclZDp9nJlFTde50yY7bZhYo3p4iiYCKfZ
l+6QoeQCVp2LWrDN7Hf7cN8g87rr53sXrskMccIGBbSATtY7cpADJ06JdMdf420UaPBejuA1iPeI
Le4IiOJVgo3BUleI5YpmD+giX7kLdgwUgC9/szKyIu1Y/EPnpIgSMqPOhsW4It0WhE4Wwvwkbqst
vAodTDjNV1HM5XUU5sPZMEzhbrXyGKum8AGSF8ZKiKKRBYymP3q//R5cMPWx5m2Sldy05i+upGGO
KuRW8mMx7yPirHrQyUj9yvx42oqQvSho0CtZR2k6EiDIL+2GugKTLpySNYb5gEcAdwtQgmZ2V/TM
RRZL+id9LjL85n12ZXOhCDslbzsUHLnO6T2A00rc+8AHvPji1/UZXxLxf49zVsxU7XCkLOLNnZPg
0GdA0zfjygzM09tpa9vTlZKXsotNc21nYs1Yb0obJ5QFJcJ9tD1MWeDLC/4ZqNhk8Mu6mJfYoRjb
bWr+j6MKwKbUTBj0tKQLNdySpYkU63ddEIFwmtpAI/od6TZRBVu8WjAyJx+WoL7vCW0BeR3tx7/x
w9oKJAiVPu6yifZHtiLlQnV8ers2OyTP0QoUXUUEZzdHXNOZjOp2wIkFFQXkvoHvQk42vpdt7/uE
yepssjzCzQPvnBJqLXy+lGTsdjHFrKZz3GjZ945atEXwIOq/bLLZKCaLEduxFI0gjvc12d5yOu97
d/DVqn18YHHs6q4lE5VYcyq+wXp6vtmzdjFrsdvz+/lM8dybd0DcpWAOxr5dQi+6dE9yogk4PhnH
d34NFK5A8/2AkmKWd4OYvnblYBAl14bDs5qxr0Fe4FxX5jD3gbam5fDFApRI4dawkWQXn7fIgNyY
FT4jV9IjackK4HgW2tdMBYCuQqqn3zs5Kq+cx4QbUNKpe6aNjYBmrtyrYDXi0iyhGmFieIMeAn0g
hm9Mi5EL9xwnD2huN8L2vDlCWYdwMg8H7Z82cIJj6l2GdL9MrFZrNU7l6EWQ4Q+dEVr7uAUp+dgc
mn4d+CVMonxTBvfuN/p8UlMuCVnI2A9Q8ccRquMPBS1l/bghatLo3ok2RFbeOzHjo+2LUOpsYQi/
YlL865GNLuRpr2CNvsyoplFHFd59EH03/tOYDPjYi5mpYzP6ajsLBVACALfWgn6pvmkRZjJg1M5/
RSb5MoP2ugTHWsv7yLdyeboRGt92Jk5rWrsMX3S1lLPwJGNaTCJeLkUHuMWcctCco/STgro0NqqI
BhmkzVmtXw00xoxSO5k9Q+KSL+WMvE2Qu+CrOlE4MICwLLsPSyxyBLFIPZzIVLgPTltpltXy7dkV
gjFiUw7OWkBc9H9AYw+dzjM18X4AH7VvIaqYcGRivwVfv45Lf1XZQrxX62Vol2H4e531AiIP5E78
oB6wMwf6iWUh2CjhquitmxQm3Lfq7i+z92ZOxdTO+VBreASZHxJsvqUDSmVZAEU/06k5e5D4B5ii
ImwqolLOcT0sPafoTe2oRJqJTqVWMZYQ/pDM2Odk/JvAIpm+2IZICqZcWhuiixeNNl0LU5A/JPeK
tFGa3yYw4FPcBbCnLdfNl9F8dAyAhNRPpwWD1qOp3SVG6jxaKE9DGxvaWY2vCU4qglatlH0LCIeq
hq9F9/5sq4+9NuA9IkiQkLK3KmRvlMqL3Hyk32gIFDZw9p0FivWXuUFD8pmnseUgS88QOQu37Dur
mitze1XNsAilptqwQl+jDl4khItVPccG/yAIGRXEngACmit+U/2knOmaNu3rKSEuUuYX0NoiAlTh
vjWdRmUO+EFbdEimEturXiXer0HNzRhiYa/+yZp6uLJMi4anJS6HjjwVFuVX1X20YpPzUUbW8+23
BI5xgCLbFoZoAPJrnDDYyy/1SQOel9nItNtoM5XHIpvRBBnWDvxp9g5CdRUkoDiKJhwaNv0akjOC
NwWFe9PD+Th+AGoGMe7+mPiSAVZYgBIve9qc4AhAL6ZfQ3ZzBIe26+xWCw0Q7C2xL1EuFiCdn4aI
aBwtalDOf0EPPPVD0fClmzkhI/1+HzBeFfOHt4Ygl1ueImMdA+li7ayD1KG7XxhXPUHeUGyD0FHw
/EOPgDusgp1DbRbDkR1POANAGyzWH2DcAk0APhS/4A0gN+9eogiYu4+8BnHNEaxKXTjEs7FPxrZ6
974IT+oSjGUljJgxGQeGkHNPjnmohn1xQxSXIZPOJRo8/x1CI/SUtkFsvMVxt+G2qer9NVzt+cnF
N8YsMG8aIdCH0An3x4PjOVrZ1107gMGJQHooVojcoi0KndJOQP06cAhaoXjTfskC0v3cOEBUvSmr
1WsJzIjVV3G0OSOjSkdkc0UfFix+Phq8OzrmrRpdJtUM5icz4yDehN5INEjHUr19roGDWdNMB+D9
n8hrC1sdehAE4BARm1oImgf4vbyaZRo65IIsZy+WS9o6NxT4ImYrVPTriikqXbHXn9cf3Fg5wy9D
B5Dp3r4I1iAIg0z1/vSgj7p9Nj+0JlPEv8VjQTVWeUJCy0dHoHXSMD6IR8jJkIU2wFr8/32B/K72
gFR/EtsNH5O1pVVvwZ1kYMuaq1WLoIFVCi12lb5QZban3gQTOsWsLMRPIo0XGIA7/seb+GyFEzhF
pzhc84WANHZpZgRsmoWiuaD1hGiseWF7TkkmDYmjllSv9NQQBuikHXpErKfH7EuoBzyOaecYPE5a
SsFQqsPzmaw1xqugwuaamac+mhwUeW3GFMfb5zQIVD+t05yRwktf7tfb8ulGbUYWvxzKmdw7r3Ag
8XgDxns9fsbYCGNKcnIr53D8lHI4z5Ly0e+V9AcWWHc1/BVYpgz+N/LZHQt7h9ZnXw8MSYpaTMPW
DggJn3flQvrAyJ8ww/Xrn4uaVzLG7rVbrSUFGJCyxvMBQKpsTy4WfXNzf4SDuc8gw3fnLnPzy77X
gnwasoJbxYhWZuEQPFCZP81RTq8SryUKiFfUriutXGkRA+DyOHWhP89H4mlWtvRWReztVfKlMlTM
diPlIr61xRaJcPxMCFu8jj47QEMrB7beA/mGawKIv2O9uhBH5mOO7Gut5LMmLrngusX8X5GgpCHB
L6HT2W08tl/mykq5EQsTJhJ0luHS5tutIFEtirh14Hvnm1bTum52V/iZ5H0DIxsuN3o2AIe/ea6c
+AecXS6bBSsx78xijyVwLMTr8NTAmjX/4rQsG1rI6aeA1BDKHcQpE3v9LptdGXDBB5hhGBVrQjt9
krYfcCaTvs6IqR0JGczeyhkzKesnX0Ukf4//POEXdiaHi2i5PtpiphOclsDMvw6n9CZaZGxHiHg0
ovgFR29LRn0VEM5E7vpjHAWhIJO2n40WEJSOYMjK4XwBoXvag1og0MkwQkw0SyDY83uFNib+QBa6
EjD5hjcv1qjPTolJjFTHVVpRBr5zCo9gCBEcUWupQvyI3ExrxFWU+8zdiD9vF5RVMWshy07KlmDx
bTVAuWHNzyh9KGvDSKiAydraiBJFARlfBXSuausoEXzEFcLwnqaY6/0iTFf6/FQfRx1uik9DetcQ
pJJysIMWOHbJ2QEdPxd2F7xspcuIHT2up5dV77x351hGKTZ2E1TbOs2du8nSBqr0RJeI2BaBCQTN
O3JvKlSsLLmhOlNWwPBnFWy0c25bAe2ystaNGv2ue4wDH9IGxN3tn2mD04XmWYyn3lpJ5lRkCSs7
R9aWt4q8vX4NPz/R7w5iRo3Vn+qJJe85pXdTA3PGPy3UYAELEWWD374k5v1mNiZBqIoFSvtku1ay
r/QW0FaqDLovQj4FwwMqAwv/67cRrLSgGQXT1R070YRwRtmgi6MQizll/yT/cWwUnYyCffykDJPd
GuIez8Ky8EmTj0zPPN3hw2vNBaMWOztGySuZoFvatvC7Tuaxno32dZ/HPLNeC4KV1+UqVUzs12t4
taBkQZRm5lI6G9OAv5sn2mWi2NSHOwSu1UHaf8jrSDvOb1+ASxWDq9ZC9R5lkchTdBXnF4Xlo5vU
qC4svCXlRTMW6KoFWwBKwzHwaIn3nfc8XhqAhUkuOTJ9iUGBg/ue1vge053kJCkpEwLsQ6Wk2jSZ
xFVQ525qf8hXDTjaGodhjXlcXlRgn6lquPlbIbpYgm5v5bGeX04RMtDq9WcT5HxrVWd0oUcqjiJM
LbbuDA8wzjcut/yM5mHC0EfICofCRYg9kWMnExY9zOWY6D/8trnuzUtc0Qj5FERxwupmJ65TnRq1
fdE4HvZYbTcje0+78eMTg7jsQpCaxloDn/ByBQPtvnZWj/VtUb527s3xMPMgTWz8UB4IFacBKPS/
59vKFMn7mnmkJBCSDl+iZHn6Ra718tFrAYMuXg3Xk/YWGZUfOLY3v7E2b9IANmODa9PIKbk8ADLP
D1HkrRCVKo9obq8Z2R27Vv9TL4MClNJitSmnlCDiyk8hluBxY7jakPI06cXCojCTmHZlppToJk5R
i4I97yVAutlv0xdUGginR9skwevM3o1+uxhfAcAJao2YCEuRsu0yAUYnoRoaXgv1NkPMHwjk73Fd
qGow2O69cg5IZ5975pX7Q5yy2Z+nI0Yr0ur5x6wxlWFeJDdQsMVZFUyzO6K92FQfWjvPb8qVUdAD
Z9NjUYktCF8xG4JgFrZr/aQ5FA3XtXsujB+xfLan3LcWQsyGJEi5XSNd5MfyfJaR8WnaD2gZYcf5
hxcdZnlksaJ7EgC6+1T9z3qb2FmE4XzIpVppdca77v2PGe+7yQ5kL1AZztYUkDbrfmnFTy5Ag87W
6xvuIJEUqJplGTvr14I9X0YBML56ahSzwoybXNyMhAfSTxUnkHiHkyM17O7QBdEeiu+f0K8cyxhO
TADgIQGcC3Vhx+y3xcsndaE9MvSfIzndD4jYJf6IBIU6GgwbQpfPySmEiTa7eNqUddF2SCu9UipV
c89F4IblWEkq3I5hw4MGPR/5HdZn/3/Rm9BnIniZQUL21cKIwLDCgy4WTxno2McxX5T4noj5H6Fd
bUSwawApaH34DiCTXdevfMI6ydNqU+G/NqOpm4KyfM15q6hkEXZO1BphGdcZcW6pJzo1A84cwnLH
cyVb4RnkPM5jzY60M78BnOgMp4wsvSHqG4vS675kGb1FG6lwAgfD/LXaEkDSaWbIM6ZzbIUQPuB7
LPOzUpjNnc5x290T/Skiw1Obz/UBC5fKoSKcAaIB4mt6Z5+Kl/jHqCyVgK30vl32DvdxqpIrjpuD
MmUzmQ5lo9n4NhB5l2oiSl+muNsmgTLFI0Q7o2IFtO7PlydCHwR6OV4Aa45umCwursXdqET/I1It
WBS2vyD+AaQ/VW6J3yUQZcmHnPr1zBPi3eeHlQXv2XlgIihc5hF5RaSEC9hMryBPlwGCJqlTrxay
PLPDpIJqFOySBlKqS5j3N/yFfdBlApeUOW1goDXUT+jGXDCRXGp0b08y9GPVoFg1w9kxLRdhUkWH
XFR+5TOOGdc1ZGXEY+5/nGA0hIQdhdFFcvLkzDRLBiL9WBc7k2VSOM81epVqpY5YJwbU6xPxTKfl
f0Si5iPXAlhIL77BWaJrOiVYSyz9nRvtc5jMG3+gjFoYahiUo+e432kt3/6ixfqcOq7fxlfGRCr4
ddr3ukIKFZbd5Lm6ZlNEDDWaQizVsyOy/joq4tJNYsOSWynoGH3d/VGx2p7CEoSSC9mGTWxyb9jG
hO6s2TkyKDRLkF4u/96oiHdbRnUs01HB+UgkhpeanBZUfQUpjU01Hwgf9xtqKuWW7mf63E8JPuy1
VUMWDs+ToymkWc05eNKUZl0nhUUfDGJFR3acSNrbdqwLGcCHFr7lO2E7Lu3f3zOwHdlaxt7Xf1mh
k/6Z2qxwg5Vnn4hnMiTTcYxHWOeuzFxoijyGWAphpBSw9iqYshAtcZJ2bHC6iiW/tKhE2uz0cO2s
/z7G+hhkRvOCaJgBsAF+Bt7d0PjWKCJy1qTThrP9s5sFveHQXJ7mKI5jTee7oqJ5teaffiY8NHNE
E+Tju8ot7cgaeiuMwYuRpJy2i3pYqiIQdokjgi08llwAduBBUIGPIzJqMjx5nbQwreIBz6ijDVT8
kP5PCywhFuY+95Gatr13d+41xCO0H5yaGNtvVyaRKrveIuZjimX/aL+IQKeNlhcS2Iy5DPc49/aM
PAA9ryQD55W2sW6HCUPGWbaJdS4XPMGJrzYdfkUERZnsBMrJYRPGnMPI8nwe2YKU7JOU4B22Robl
gs8eCovQtuSDB72+7UopmLPhyGG6c5mT9D7xEG/q4hvftogeyWzBKS5WWi6H803teZDazfVPxowc
8KaGeD6mz8Vv6WBfmUta2XfKTPaL8bNg5E/uFSCEuIn7al0AeRw2y7dC2CLbJet4/GnOqwo/SE6G
BLUdg1ldqEYcbi3Z1DKLJFHmfH0JgJb2LyRdbmiyKaJKXwG9ieAr2En/afgw+fhkaSXyhPV7Vbjx
ZLZd2JcjgmZfMbRpE6E3PUpP69WX5L9kZ+se5qjoq7puPtHZIsJ5bD2tkbh13HWNohtBvr1TNTDk
ikYZK186XLUswMs8GSp6hcbak835mUE9e9S1x9PYAUHFgQ/7U91rGv4Pn6jbYr9XnR5Rw9c1JnMP
DQywq8xKTlJqdgXhaglCgr2TSei+GKtxmvNfnMy5kuR525V4qrNltgO5vDzO/Kv75MJLS7O8YLvZ
pkx2ZOG2Tzotkp8kqEhrcF9pTUBcmV9S4n3OqB/38MbVf2farUASKmBqIn4ZuM1x2slkD7iM+rF3
YavrODY2FOQuwE2BaYNU6CJFHB2gaKsS0x/WMvvVU2KJekSZ03dgtcMsP8E1QeeKD8ZQ7cGO6i8C
mIBNilqzTJrMNuDOcjmNmwYbVfrUO+0kiv2pqwGwlubAiet9XTkK0xY2+72NjVo2XHQCoJVRTsbq
k0FjuKzwh13ZxvLYwaA93RcVBZ/ji0HU8QD7Kl8p5rYyNF5WbR13KiWDQcgAZiX+McH2F1kG+VB+
WX7pzGQjuFtSHfJgBLFiXu8rhSlOc/ztjoqEUX+PtXwfoLIwtkGbtnhak0p8eytCmgdz/Sc8guok
ErmVic1BBMWz5dqIkVYyLqfwm1uslyYIQmy7XRc2HnwV3uKk0Z+LJjCiEVvgRjBs4Fn4/Pdif6kd
USKWnOHE3wGsEPRxOKLlMU/tJEXVIROe9xMJgyi00Bda5L/2oYYswKEipAhmSKlPqid9yPmb/evX
OpN5Jr4J9DbNbWIGWgLlOCPKlNBifi+jyk6rNTt5hLEwzDOSFwYH7Hnv/qif0slD9O9fKLJ44m87
eQ26m4T61eZnsbNtoYOyLuOIMjPVbJ6d5L6JLB5hhrqMQqB8ZeX/HMfIbhz7FB6dfta6bw/GZLyU
fnAQlNsLvFltroiHQOX4BFzexz/jGaV+YTm9jCWU3dxysXVVoaZx1vab2nKxAtwIL+h9WgBSsGdB
OC2mkxyKaPUfgikPNizkvTN4HwyWG9wpvBAYTb4U5ovW80BmMj995aOmG/Mt05cm7SWyhOMnt8cQ
Id+b009rQ12rQr/vVp4w3QcOzbzHMEOz9lZf7D43n+4/211HSig8xUg10vNnRLeowXbs1KtZOQ+O
RAMiWUQdyBvNwROe/5mxvwi2XscXMxLfWfg1X55oukxlLqkyg5rWBQDfiINw6KAmy6417/rwLP8E
5XUxTf0Q5j3TGLa3tLANwXTbllZA0FfmDojZTsYd6EEM2MnWlMFHmCDLff4+k9+R/NPzT4qvEP24
8qYKbaSyLW/HBlr4aD5C9/FDxEq7clSrJ+lr/rvQajnQ1QgeJtMrWxFYx8fCXbDVnBK1J89yYC0g
CYMOS5MKdiVs6ZBsfRl2LHLSDC1hnPYakHkIiH1XuZYHhiDpKD+XGJ1Z3z9tBxIoSxhCEHXM1olZ
ImWSVNUlg81lXuBIfIS2Sc9k5mfACp5xUb5lWXNCG6uVq9sFyOQJFciU6xvCqmf7wQpim5SZHXCs
vjP7ipQi/ZtLZGCLuhOZfbNA3aTSU3Wv+GaJ4ej0d+W7ObTZrXOkhmTBAh8xC3+oKna7fOlY9Jo6
lvuNhm/areYN8ZpPeZ2/kG8fnqjC1DRvZriwcpuNsKg/uaJIdza+EFRCt0D5NhgSDi6QZ4BMWMxP
fseky60WYVIbnpGmb3l9jLLzEPG3Dulq3oOQ2AFRRIPJyTo2MgoccDJCT95GcM8pwnBqXaiYcsuf
Hp6E1wdo8CpnOz/3ofAnCd3cRXbbvSATyWGgIBjByo+n84ZNboWtXO/63RkKLohtAme6aoPfNCyt
Pf3vGszg95gIf2lr1f7KrUEbZHA920IDdJO2xEk7rRE2HR6o6CUM4GfOWQG/1DM2TcOyrouhh+TT
Ooz3AY3sLj7Za827J5rJqPbheMgjp7VwsZlIbAUEyTI3zIjroEJfSd3gJBxChNaooMLofzeyWF4q
6GJetk2l3DcNhFRL7OeFnWqrC4vbJ2OF4FlMRfmr8G2wPDpJeAZqiPIiEDkPYygzheSAJ89nH+2j
svE/U9jZIpTjRdfjKHgriZnjeBXH8eku0pL7Blgy6fZBg4k/OdAcQ0r0m5Y2h+VtJUWo4Vib9Dh9
HkXRBFGSh/kJs8i4mc+yqoX1hMSBJRuOaFdl8M0m1gWstifaD0MmYTDsNsB3JcCr/6JgWj0UkVDE
dWNwmmbSl/mmbymwvHSzrjMQ8JQ0eZrZemvEMtwjrC/q2AqPXcLEs1LMSrgw2ztQCmByEgL7t8o9
cUG+c+K3lyn9MuHK5rz5AuPSqOpwetSn+AMmvLZe23D4R5lEUrbJBJToF3m2L8RgKdugMGCuyNZG
7VakRMTUE6ZMLydbqn/yKrIm0H/VC/WxV4Gdan2KTmfZwIrKAPzOQlArMN77OvO2pRw/0b0fXh+a
3f8LYWMTxz0USZ05Rz4Ou7asEWRDeeadZZLiEHr2JR/EEeCbjq9fs3GWEJFfG1i4Fyg6VjWRqPS1
euU4/gBRN0T8i7kk6T/VkNhP879nCz06fHWIJ2vq3y52vDAyJCM75g/+wwkQ5lEjclHpnvPlpO56
YmXVu51DPpNnGo4Z13iRggN76BZos1t0KLFlCKcgAHkyefpdclGxkYccaPWQUxPDSM8sjnGBf7y4
0GN/WJBMhb8R/ivlG1cGDkbUNE/S9v6Qh3chJjdaagabX9V/Az32KkUq0ntZ6CMkmNPxORJbh1b+
rqg2C4zJXf43ZRRu/HRrtn4KRNkEDYdsZaMYNxxieybirHxosrh2tS6fkusjrPUAjsrRwhdQPZ+P
qTvBLEaPfQu3fuyvkE5XU629QHcA6Am6dT6uecJh1J6wcf+F42QRyP4iHDL7+wG6MQnGYiVSWh5A
S6A/r7TKSau2m3dvgefhCTETjj61kdfZftAHkDr0hQRxE8I3WGybkuisEbixmPOUKUxMEuo0+4AX
xvcCOXlOmjYui/E8wRzCiR3RBXu9wDPQRwwW6rAjfAygLiJ+ydOCCli/KEz8whIw+H46YTG0Ey1T
enKgtuzzMK60VxrLoVLFxDLLFFbyyO/4sbQ9Nfq3XzVGDFqtRPnWX6PSZVSJaH4POyQd3c3X/mRE
okuFAARIvIeyWYBw2txRQcw/o/5NqDsg2yDWktpeth6/6moXLgPw353m7Bhc40t+MFteW8FMUarJ
slNfuN+mebn/Xw5ZHHlzFS4iQ+AFSLsahTHCsJLn+iGsk42BQ1WY7kf/SYC2EiWTm17dwQhE2SSv
87GFjbA1v4T8HhnAGm5g8MWIBnC17w7Rmh4HtGwDRgRapA57/UtSptd4qQOdO4LMeWCpNFJoXByu
TMivdCuyn8XLOgkZQbt5mfwte5lKtIVOzmtYFoa92MRXRPWl5FinHDaxSysDRLVrjLeY5p3hQKlm
lUuhH6OIBM1GVJy6Z6/GUTlNryjZeGhoDsuZIMmcH9Vv4PKQjWT8JhunPqvxo/hdhIA82cmNIRcH
uwumNdUqSaAWPE6fQPN2bJ5bC1wUMMlJNOEeC+DXRA7dJRVUGp/ycdcyOO1VFSdtCEaCJGQ+im8w
S/xSUpA/AsjLfMkB+hPcYZqHR6vInnmEspHdVVAFfBRICl+wuayQZZOYRZJ1dryF1sT3kW6F+V+E
xy5m6GnCuVNhJE+rQ9/Pht/WXDiWgRMW9BbAgq8Z/JLLmU0wq9XzvtWklx41+HbG2MlOIrl50k/6
lDImiBEU48l/X3JmYJ5mG8xir+EEpe5F7kM6ReIfYYphm9p1P6fl5rszvglfl9t+EhkarOANwGXl
GQk2WX+qCBBx709tAgPzZ5qH/pfK/fhVIcqpf2e6GtVzniDZrqYQwGAz7s7qdBbugoewAecWQEC/
zWYEFy0clzULJIqupTb6WWj+O3vZYJ87u6BilBSxT01EM2A6FJ5yzN9IoPCwaoZPVCHyaZ/LtzS+
DkOCrX+2RHLK6TTTK3DuFP9fBZu1e9gtSUSgKelQ22oolaWFXsco76yDQnNmDvsi4DI1m65uEpOD
aSyml4qBc+GN5TKgkygRriMLnGmPj91+YiDzSSYvBJ8jrxAxnKtci9NAI/zuaauJl1VlvyrXVXvv
sLjfw4Zr2FLbFFR2msVbRTU0k2Nyu1nxN+p+g1l9VJ3QFEGjBjqCaLFD+eTP0hyN3Eqg0sjIZyUF
yNtYsCao01bslcNW324xFdF0P18JuLrZYU4YDDdLH+zmHoR4tTXsBra6gUoDU8TqWDxcZAlqASVI
r86hIGQY53SBYcT34EG/uhY+urw/5hSp3tU+nN6/yMKiImvcoMHduPzuOotpCYk4nIrTt9SJEDcU
h4s7+xe4D8u1A8KzZj7imO8QHO12M+7M4BLZKs0Zx5zlg3DzKusUM3PdQul9MZXargw1Zp01wiWI
siCqWD64xJBnXy7t16PohoLbxOZWucosket94eAi9F8Jz2uP8ERGtjuHFPjwhosjzJPIbm3vmozn
UwrSEhtmM8ogs7rDzDBA77pXylxzbMd7IjPHP3AG7pGdlZvQXbBzG7EIDNrPaiM8Tl22fVx/DYGO
HMcTmfNhORq3XvmO7AshGskd7g91Ebf0i75pKJs9Uyzigvnyt4luv0k9JqhhqWIDqekPwmBRjaPl
A+TfES8H0r9aRzllWIWHXce0pEHqCbm7gt+O5fKWq5W5LsgoytatLmRHB0GZwItqCmDx9sBtZ8a5
WFFvN3LcwWiGGZNNyiH3KFcxH4RZs01S8zUAmdCG4q+3kW4bClpKbUxlmSWS5q8aN2FYYH361Qrw
dYj1uT0y5P/bqjrzj7o1G3nMzpwkXp7f3FfCA+fGErA/kLFBxLWE5sVBNUv+yBjpwjEe4X+qW/0Z
f/1ibWcTjV1a7O4TtubZu0TjqQrRxxV/uWu3xhzJOyPtM4uJMNaR/VYujY3qqreByOXW/gg05pZy
a52nLWuI5MG5nr8SqHcgbsqcjxnnEvGzZ1YhZURSc+l/xZNSmX4vP9uD4lzuCxgjfXpUyaJCu8n8
luH1SWq280gSPDyQObzBA+oAdR6Swuf2pJYj5Rh1yKZ8TFE0uZK3uz9l72ZgA0zcmbi49LnzHEi7
huIJNlJZNksH8LwJclDa+NcdIzynvkCUoy9vzYL5+6dZwu1jy6+wo+6oG+F+KBOAvmAydzMYOkTk
6CUbSc9Q/jlxNh8nFURFxvCuBSvLDDxUpyeKnLn1037NkWIlzhz3gzaNsukz0kPERHlN4tSMhvVB
YdvUy7mKORCe8/NUI3wzzqk05XLPb29awIMRNWuMWlUiDKLjS93DNN5gDRltW6bjbpHU+sLO5bgx
VmlKjt+9j8KrFK32mxojhppJxB8xmdgkGIRj/LlzaDKnNag/AZMGSNzjdhr0HRUYFVL0d9Slw0hw
fPsMY7jvBrp3bvgvq8S6NM7XF2w8qAhx/QX9PR6lkp2cWtas/AIYCPRPz+1o0GC11OA0NM0oGM5K
t+N0XUkJCWdzYF5tXfWfLEaTmoXDNDEtsaXLWzgQRWSC0Pg8b5bRhiErWnC0jJNwzCM7lBbOK5xu
/rmpwws0bFtBC8JAkbHgMezMUNNETw1RXbP3Iq6foFcF1MoBbwsxtq/6e6TyKciu0698+ueXrVpF
cycKg+jgZ3/elvSINm+i1F4n3O6BH8yxQS2GF4eot6eLD9TIc+1D84gKE+RxcE9opJOZiZn0WevW
Y+V7WAXyaApbF4zYoT6OHJeTqJDx9uviNHd9brn6e+qyITPhoVuF3quZ2zHhZs2xWwSs4CTZKLzv
/qEyXaTF0s5Uz1SZCi6H0/IYNqDOcXEyb3BtOenVoKy799QYzZ+0viZq/1yNYQlfr/vvf2w2KLyg
2CFCo3sWcbCJLTLbEZN9o5L+D+9yuQOKshhVl4mMDpsZpFLg2y070L+KYNtMWdwEl89XUa/6fA4O
MGLBPY4ei2u1RjMd4rVC0izfXuYFB9m2SaQg4kimOvQsilQpNIWzyPxgdQLvxxXtSNKcx4SsyYL2
eBnS8Ny/fSHkzshMRp3OBHkH4EBzTzGHco1IO4nnM58dO2CsWCawzWbF3LROKYkO9QTux44apiOf
PaAhnxiQhiUFHHtj/ygwlm3j9JHrmS6JLRBIahviyo9m2PJkmzQWk0d9oPuwJG2moED/9FO/kOQU
zEIV/yZsfIVmGm+ibADC7YenmJcXmnu43ql56AQJJL8aA3/o8/IK1Tg+9l8RH2s9NnjXKmtrM7C+
HHfC5oXDxqAv5OLX3CrBlvinFHqPrOhkgcJtElBjPr0fI6OPMdfBQcr1vrrXU04spsOkho2BsSlB
1f1NSsgH+qOUHPEpByhpcol1Ol7cE4FL8jab/CeRloKw8AAgD9Y78EU2axHBncdpQ2mbbF2LjkI4
10Im1O+2w+ay+2CNPRIWeyOJOajdtshpNI5dPrb9YM2qFPY6wdeCwcoHBTZqumlEK9EFXw+tKehv
dFEAngYGczD+cy1ExZWYLAPOXZF0bsbV3Md+D7ThsT1QJjez/gCOKSOunkdkjOQ7P+FqShF5IWP/
HE/N84glkcj2KYPmrM7r4x++F7QDw/ae7kUoxv7IWzJp7R+y9X44ik3WPGXxeMq4PAlNrPTEFsfe
8Q1xOPetBxMxECHfVmRm2g/F8mMBtBJCJK4zvlZLZa6k1WL8TlaSxg1EbWsitVaJTahB0c1R+sYS
ZAvgLV8TqXv3bvimlVSPUl1oxwgEShuKVn3iv0M7EzeG9f8+TJYjQQr7HumvBfrJTov+0hnsE3dD
I+F1Xdo8hJm8sHE5AqDvODamy9LGMfWR9ZHiec8MovjQr2CEJ23b998/+ny3Pn8f25qzMHnkU7rf
ffIVQFKEX9VNbZr90rb7TwW5mep3m437rDq6c7hiliCBv+HMnaOG9LV0lrliISbfXw1haNYfDUK8
KK/UfqJuh9n3OGAlEy2s4FSTnQ2t34bfeaz9zWnlboqYGc3pFQqs0oUKC/o3xIqPlRca9z5TjQT9
ZtpWMZ+QIfW6vLmZAw40DMGWw57BkNiHhdnn3DD4YIvF2M6Ldwk8gWTPfRR+27msrDznYVAfa1KJ
yBfnqXGfFW5S3reu8RdLTSjSHx6ujQEXVnlqsWyF6g7y7enPjPmAnb/4zwk0GvgvDrhzxhyvrgs2
KWxx+z0uWw7p3ir+GiI9LcUL+ntzC3i6kGC38BAQrEThCbjtTE7j8WY9ns6gCGKMfrRVdEIefdOg
fua79813z8oUOed52gcq94oUDzDWZxzSzbqoL5nj2AOFNyan9Kxffs84wWwFRoniGLi7bIh0vznj
KSI9U2bLY9DMvxew8uq/ff/nDPY/pTp2KmMhVLUP1o9sZfsrF4qhfDZRlDtUG82bg8vOX+BIIGaY
2MlvnpIT2ozFLCQexPpRYaVvuGzjJVfNWUJv/eQXJBG7nmOi61tvUMjJ5GkwKG4wd4jvxL8M7C6I
Ki7SLmUZbbibouBD0KnXESdW+Uq6TPi4hTGWwYKtSsqNN4R6lrne8ieTJbuyxHk+VY8YE+8Agk4N
VSyu4TI1yUOAW7gpfKeMhyQdIZCCY6/f23HMNGL3R7m7R2lCJzjXpCrMJZS6H0hgJJhQoCKVcjL7
pm+t2/OqgGAEcjioFkmVSVTLLkWrMsWaZOmE29J2YqZ4X0KvDlea8Zs2X/Zs/oNnzt4sXkNiJzmu
JdahofQKoIT748a1ASMg7Yt4JEklx2UezbongQVh+VWhXzudtypS9UARj52whaWXs9zN9bazXyLE
eTINTyTgfkPTV3DZNiIjdrKePI/XHOCyb5EugkirggWCsvcbtOOPQyDXKZ6W9eZI0XKS53Z2N4uZ
JCyWtEKL/uAE8a2pUtRwIiRoOwMsYz0dlEZX/RJQHo9QZFZ9dmrVDEjLqbn/gf+sbkQOUTCSizYw
IhlvYKPOgTFRbiABiRVv/tjCJChNHKfG1gRsE7IyFqSZEhRV7djVZLZVOkOq/VgdqP8FeDKnICiR
wyjIuFauoASV0TN4MMfSct4jg3cv5j2UWDKQB1+VE/u11E6rQSVclKacmsCRQHF/bVMXi8Bi/zpN
ZQY9XylfcMWB1VylS8KS6sLvyTw51UwH0XNDbnEK8pSwJ3PFivOa9xRhtHdXUnnL8MKrcPb97Wm1
Xpzq7RHiFfVKUb3f3gauBCHBitR42x+emCDr6FwvCy91n6VWnFzM7iF+OVWcEtpWigWFHT5j3AOk
+vkg6CNhUtE3eU174pvbQpvMMc5sLunj6YhnMCBR8bFiHpKU1TDFAJJ/OjwJAehQnHvSwSl9Xry+
r16dVaHiDkAHwN6br5dQPUr5H+OXVdYN1ggOc+TgPN4FNUJqsr4qtEstL6WosQks2tnbgN9/urB9
N6lsx/OtRO2C6YGygmK7s1VbnnrMu5i/rDONTVQO0mtYB1oq9fw+h/wD5GsBkMXCPu6iNwW96foa
qjT2fyUQtC+N806ZLFhADE56kpEPprltdcAeASqJGf1N6F9mydqYXZQtO0ID4nAhO7mCrO3iI5qO
ZAAsTbKGzmHGjVy3n5hLusXv6i+LDVJbt81E7O26M7zuYB/S+MXJt4y6iLJStRPg/dkwd/uZrV9U
0F5Yd1URJq6bbs8074etcDB09ZlXkxYsPNs9eavAKiyFiIbV7d2acsHCli4ydrFcYoSwGi3I0bVJ
O+x4vu96X0PJdZH2BOf4d9wUytd/M38VxJpwu0X67uP6NiTbzFNUkHjw8VUPlTBMXZ/LbofA8xTU
j+1QXV0YsDYgG4IVLby5mHTG8qA20R0TGuEWu8OfHcPJBBif7FJgh2tOgUAzpOheTWqZw9J2yWMJ
xLWjZuiOwRn5rFK6IDAIaTC3LV5ZcuHYKy+52zKYtz2npMbQ8h2mYApKm0EGL933piTvu8+foPdT
wt+4rUoSVfwFY582yidt/Ns91ByJWhpkMjfNHKsuNeCnbShXE2lsBHuaROiom84JxM11j9M2EUki
i1ybmqzdu90U9PRDLiP/wotH90xnqSN87ktVY/HGBCFotR0AtL1VtEWqKSt3F9QK0uwh6VkTv9w9
h347i2ShIXALfcWM7XTgkL56ZI7DSuqxEUl7Vc6zlQ5LVGm4FVa8yjPLEtBAhcnP26R3Gw6AUEL2
uai5L6qznPax9hIi2DObVBzTfDMIjeuO2Tqg2cbVr15sYbW8NAKki8I+lMXJyAwY9h7pGwMA9Jmu
Xjq7RR9YrMceaOVtTF9oK5NwM5gQctjUD0L8RLaRPM5MUmby3FDKpWx21LFsUntf80QgX4/OJr3r
lUV+7ia41/HrduJzcFHKT0NF9a6gCJv77Zr7acqmpzcPr26yRHI7dotAxSbDtaKGXQJ3u2nNo0Ua
05UYHePRCH4/Gf/4cnmrWEQPl2cUAIsVxcHw0e+sITujmRpnb9oqlIJ/BRcRglTsBtsaHpBGeMAm
1VKGIGEjqnazv9Mwav/KBukIvjK/ItjE7uickaANPPgn9hUO0XqqjC4TOr+WKL5GbzKrv9MA7RBl
xNpP7LFQcmLf2Q9O6927A22at5MtrguH7r0+9f1YMdHtdpEtDkSN10RLSDIkRzJyWWpLIskt4drO
57qCsh7s9ptug1pyVn5KqiaJNAUkAVfvi0ORHlBoS+AUxh6us9PLENtOTXjp8H6MCSCP288DBL7u
PlMU/Vi6cHHBYzz1peC7onSjtLRyIfY41gOcfN3b2yKJkBUgXh2MnXPgLhayEHcCB3VO/y1cVoG8
/ULdAP8kSG5+s4U3VuQZwLT6RZVZeAXgdpMQC7QDmIduwvlere5V3EnO0NqOohxXB+Yzg1wk36Cg
VOk0R/+vvlIvNhruArv/eTdb5P55FYRd69NtzVA/WA7Zx8vtivK6Eu2wF0U1KZPZdcCGpLjlNpmf
FyyEl/SyT1SUQXcBovPCE0fivlVqcViVLOeHyA1tbTGdlkq9Ieuua86K0JQ6nGv/K9rfT0MJ6mK/
brKju/Hrxr6AagLLqqKZtI/t/z9ozgt7aYYRnMtjMDuP7KRSpA6o55HCE/V0JGGRhfEszRNCXtbf
ubpwhx9JUV6/4v/aCZ3zV8E+tKS9NPddJcF5BEO95qiV/LJaReiWajLPsGiz4z+TaiHuCamYWajd
cHoAgTJDjjOrjfXVyAV+KBPyN6JPWw5y7z7So49q+NR2/DPl91PtITpWJP08bA/BAUp7TrLEpzct
gKerAMVfHQGF6leEmqBpHGo/q6tOqOrIGIIHhh14w0A9mhq9xTvhdK54jOj/xEYjRBYZtbKXuVV5
FF7ArUo73fq/syCGJVRJWy/34m8B0bkDdFGAYx32Yg3kxEwiTtHABVAlPOScRoLkloiQKyUtyDS9
KlxTkiINYiv8cAiezIBMvBRyGMD3oEAnQ1aNKVYxzrZYgOL4eBa8Aq7xTwnHZCHyQEmd3n/+vvrU
AxSqYj4gQlQxUdt/hnG901S21bjPxKjNqqtNZqcFZbsEef3u8bHa/l1vWczv3bqJFtQhAikvNylE
AgdQAQfHx/T+zb5Lk1MmXkKM66BiURM2PPa/O7BlSTzgRQKX/S5uW7aawoL36S7UwnHCDRgpd6sw
rzhw0MhFh70goz4+j4sHNatz5xOgamBGgYe7V8w77FHiKCaM8wiAbIiV4WGEDMCRvZaztD4kKBgx
INbvyPpvqSgS+qZ/nY4zVba39uvk9QdBaAN1OwNGpmz8oT8opQR5+9wDmM+C9L9jkc8wn1c1SUxd
lepK7IqrKtBMgO1d3PixDFAYzZdTJPNZEIGYd7G+mqnvopuIdPy4Ett0DC0BXI0G7mc4frWjinMM
kWEuwZBzhqrN+rE+XrH6GTRdxPyVQfVFMnLo1p+l+Yp40HKVj+zzsTwV3eZxf4khwGKbNyaZ/mzu
q9FEGvnp+fK914SJ9uHG5vFnde1nvdEHL+6PteACyP1/9y3rsH7BGuBZMzVtycI50p6LB6r8mHWE
HLVSW0evM0D3ldD+8PjoBuDIZhOBdepZLC7/HDdPvUiMRgTcM6tYUXztNPFfwdPiqA1QyjJG8nuv
utJGLrB7hUMoJ/hEUWNKKZI1Wp10Vw9XirU67UwM/0Y9Ty0rtoG9aFJVmUA6lFdJ+NWKV2ek5Geb
D/Y1ON8XaEfCBbamAvDHKAlxhbtCBJAi8edR+vuYrxZVxiLHbOZfMQb1p+QuDG49u694TqpVj20Q
T3Wkr+p1G+kH5EANGuwOc1WWTa6JsVKEqMxWkCArElKefzlcc1eDGMgDliKNmbxXRN9utaVFQQe5
q+DbmyMEWkP/6UrVsLrd/gjJywuGN3SMI4CY7uus5wRAiRjFWKqm3IENGhvDSRvLJe5+Xgn2zJxF
OdSNOxN11zbf8zzfgIL1xLnaNaWVxvdBq3OdRJcRMhNkw39kkbjdBZCUClThS0Mz3CEbr9iNElwq
4zPyVQwvAcCOWFx84+CXZS+imSD6wETCI9+wi9L8R27dXwaH6qua1TxA3ufmMmiEk64Wyns/DIN1
9CDG+7D4rIqq+vGgTifXKkp2jXNaYq3Iiu67EbxoQkdUZ9SD577oPK2AmZ2UL6XRX06Tisy4COPF
CibcruzomKQsJYTH8C6NkTmKvBNFatnzRftOuiYNbQHIyDiCbYE1KMyfH/dK/tIItyBZ9yjGEPy/
+S1lKG8uf2oJDcv/2r5pEdKiXCqLB/lb+nEc/SDyjkG2GenzZ+kd8fKXy1ikMq1vVvfJT9tY4NBA
Im5srUwT1FvuTzrcF39NaL+krkntG0cUqCciGG5L4PjSF/I3HXEU4NgLLmbRFWTbM4iAdrMof0N4
JFNJTQXCwAwtmU74K5ltsqKGhZ79eDhcEz3We611ks+dZMscIXQVrqv9DlQ89qPfzqY0OSlR1+C/
ILAKvtEyJE5J59JlLt9x3T7ZgVw4bv/AMC+YKMHtjB0iFYqGFt+cMk5GOeGXjvHBNUEuOQqEOxhP
Io71dEijpZ5kcaNzqbqaVu7MwP5Ug3eZWt6mT/EB8TgyAPe+qF2dRCMNw91eRWZlLecMxg2wt0f0
xCGrxMJb6MZyrU8yUkRTMNSHSacnx5DaMxtbsvV8VQ5RoSvP3hQ5JGhFq6krx8/90gWJ/kVO4vlP
++ELFTiOLtne4wq39zEcrndMoqbt9SBm+TRgIEKH8FhqoMown4YLOqBehAMVYqlQ8jHBA/7p3AAx
XoQsbdHJGMkdRF6pEOs0eU7lihVyLhU8m09WRRVUy1tRkWKUkbkqOdrzYsBvj2sKrVFKgSFYf8nR
GRl3sVucWGqDzkfk8wVlh1Y4yMpq0QMweynMSra3jwQyZgLSDrwOKHgApfKuRb014zABozerCsxj
8vLoKXIzDrQphy3Kz1UbwCtvX4Vp0RdsNFcMqiD3oPspMWvwHm1P02PWsN1BtPlSwIWSNcMIfArA
hTTCLI2rxPYIIyqnuK8+pijviUmlD65FRarCX7q5pi8dzjimpAcMNvnzYn7mo+imzGfJnu6v4bCK
Br97xvBSlohMG+RwMkW79uQukQ3I6y7A9y9TYGlK1MjEOdIrANQN1B1slubhzsWEAD/svL6foJiy
w/TNILw5YrtBOSeUeR/bHw6qlK0Ng9iizW80K6csluaYNTnU9PSPwnx+peDjV+WLmthmzajMQ7I0
MWKTUyW+Mm+Tu2WII1wKqf4pQ0/Jl7tkuAL3fwknyhSxX/UaXLnBxiuswkWRwXFMSifWAEC1I0bG
VkF6WsOYnF7PZDMHrda+0N8ui/o8QTzSFg9NbP8zH8X8gcbMyGoBCyDoJKKvc2O/Y8VELz9I4xHf
WrhLDV9XReJlp9uoCTmGaCy6eK0i2LRNj61B3DLDSYygyJ7tih5PMBbUnxOmEvlsrrjhGEBpXH/p
r825j2D6Kp5U/EWoWu2xax2SfA6hBKsrXmr+fxYSP5fjW5yeyUtkmmQFjD3OMd/pT3b7e36K3feA
ynHJx40lrXGe9eepgsc5N7CcUqZ2PdeQoAjT+FcCd4MCyWntcI627y39BPK7GbONMcNyibKfCplC
vxbgCUTZ42uq6dbkYiimik1fheNQudrTrFShlVk+piihbeSijCq1VD7NsA38VFTcAw1LNMlyZw32
9lwtiIyEWZp+ip18A7LXyexAokOqmabcJu2VmWQMRmCFTYu5KYgUFEyBserH2y3aA0ADoWiZB8Rd
bjb2leDb4j4fac3H22sQRtAzD0Tx3FeWOKtWQ/juEVjSHYhkdwJLYj9qYUcC6irSuFFVFxV0PyZO
ZVLo4MjcQnm9n6y4z0CnStl9894hJLvIMd+wgyjOch2FcsM991aOSckNJzJvqgWl7feqQMpIAYmy
ODw6ebbhr6BScYO9Qrbem7nH2PXfibWjWdarigz4zPxcknZHQ3Ic8wAoXHp0PlwWIhgU9+s2FxqQ
2KYG36pXLGAMwc5w4/pIK1Bl0LCqTLFuvPfaroEv8Sh2WRcwuyNNOzpq3xR7rJXyvfgNvoK8eFtT
gcQlOUZRJ2gkwQn7U0RNRCz9DmJZCas7OECxlAoxjpL5lMZ+R2o1+OjxEX0UIUZoPxXzq7QrMatu
ctTyHHjHikwu492zC0l9WYEuDnFa2sZv/kRf5BCqXyBDR3cqOHR8KcGcfVpUcxKo6rEoqkluBg3b
9sg1XBfpjrcA7xcDqXS9KlsrXrO08EsPUhevbuSP+YPZH6NGeV3s4mhacLdIIQ2udkv699Bd5DAN
CRsu9Kkm7f1TemZaH12C4PBZ559ibTpxTEslf9nCK5k2yYLbuu2KGpDDGQrhkxoF/NZJPJeKMCD1
5zfRkBJ37H5EUOGGwJDl6FhyRnqkyxPuzgmou6hSh1EesbbkIhdNE9x1+96oCpJ8UBcTVDGWfNpA
mDy/Cw6hUJDGCr44YcsF7HTBRX7gQmxq86lK8vgX1wMS9RrzhmpERAhlp0HBEKH1xOxFG8tCc84Y
85A33PG1lp8VmYtVQpLXI8HkKyg29diBOtxNegg3zoz6cSnmFReqJnpPvkMT1rfTB815oj8/86Kd
V1mKKGrI6IUAUKG4XCMYMaxw3zCTL8mh2lY6s/KqCLvskVK9yNHGuvkTFA0yXZZhi/za2idtGUDd
hZTT13S8zHafdvo4W4EJF8me/7Ga4NPaaLRHxC3UawlawaCD0luuOb2v/wvwZyCKC8jQCmZYA8d7
lrUZ4HD1CDtYJt28KKBS7uq73aEJqjqKrG0FvUJSCxxkHZ4Fo/znc91HivD0/jcWmu2S/3saISeb
1wmInrqbwDwv+66y39BhwlRdGtVX5lEVq60qihBx4freRw81B0Ul6/xhEC1E113tnPxHEWhz3Q+S
wFWjKM2VTOKsxVwzcyitsxO8CxPMgKGjORgY3/r6aVaGOAZuY2Y7t97DvM4X1j+ipwPHF75vcMX+
hBqxMmpN72piMTKDHvwMGz6tJkJ6BoMDTJJxi+DYSDoQiUBmbNNIac6/M+5SrAOOQxtUNHeuALdF
IJmjOpzvVhTGz2lN/bI+HCgRhQ9XEqZzSab2HNB1Aer/jWckSDVYN0eBA+wwI2+WV2xNFdgWSdNx
a1uqDnJ8z38ZZt7/2ECOwIlF3HCmPExTWuMVZd3I966rTJG7/u5GLgwxFyhP/POlCcLvonLG+Tcw
+WF0Du+RkANv3RFE1v/LhWZCEPAgDwMjmC0CRtZoYbw8qJP6sOMzG/FBfdS7l0tYKHhnsZ/SHATx
+fPnS80KjFCwQF9dntGRMYuyEW+hky3Coq91qiMNTr38gomW1qv1ArHa7R7cDB6Uy3W61HWrwe/R
nVggFiuzZrbZj7JE701ftuqql29spSjsM56ZYT8vpRlFS1+SM1YK3ULcNklYV8i4VZa+Wq+SX6St
LtDFqs104TUP8tGJNjCNS0zSZiO2eyuZ724dZjOL96uFym7W1RPU+PJR69wuvf979Wutzacx69+N
CfvWJ4Gnh+tPAFYHfdMZNdSesHwMmTCxActqrNThQFY0GQ/w0rnK0ElO/AjvCwamXMZ5HdYCBXaK
gpdZ6iV7tKbMNf29sbm8PcMO7jbnCfs7f1CKZbjXT4nLGqQ6Eg0EB63WaOVI3pzJ2XbCdKUImvAG
S4tkY0sxCzKrceyBLD9d3pF3m8KjNAO+BB8l8+sskW+rY76Pvgk5ue7v0pQkTWK9GoEGs0mIhyVY
XE44LJ/UyinayWgdWIebIyEAT95JIOdSwhNhokJ5Zn0E31W+bj6K7EsBSpiQLgv4Yk32o1AGF290
Wo0bfb3hENr8bMKhPMG7BoyaZuEbM8HHmCKUn3VCYONBs58dJ3D0oo236jbh4ND0ql9aiuPq4Fa2
Qqy0R6begzKCzZGtBY0qw1p4ljh5rY1Epj2531o45kBM6oxC8exsxL9CzORZCMaRoiICRNrtbIRR
hxYJjP3aRjgUKg9RywgvRvMNV9oNeug3e4X6wZWCx8RVy0qtdJ9S1K/7V90gOqId+59Mwx9oqiX2
VGWGGDD/LENgWXI+rv6ES9pIHGXbsRQbhDRSlsLMyaNGlPZyO/n3delkcahJZ8p0rdgGPbYaZtsg
QtEim100bDCQu3dHfEBRmqvvE4k9UBSqj9WpLAUlCOyeT6TYyUF8eosagIAahK64b7Mi8s3z3/2d
k0bHatwCN3KGiR3HU1QiRHhLwsdrAUZQDBy5aQsel4HPXgXCVEoV/L3kZqGgdbGw8MJoluzC+TH8
Fu7sMky8QhZrRKQpLYtaJ079R54CQUJ5mYqlw1sd+cKKbfsmCrE8EIfI70wK/HTN3KZkAbkAF3k0
gw1aVIovR4JxA2N/exc36YhXofTUBuBjwg/IjdXz3XcQJvNVNZKUWerpswE0J0KZM6mzLkXi2JvO
N9kygBw3CVtpVZNBqSlVJd7+Z45PWBmtRPanA/o5Yik7GTkr8BBVqJsWkxqK+IipxjU3P7eSSrD3
42LT7ZoPpLHifeVQ/uVjZMsWiBUICMFjV8OqLr/gFV/P0DK/zaUjtH5cO1aeIi83RWJVvPdelw5D
0kI7m6WzR78qDh7YROSwAwyBcp/aen9jjh47xNw2AfBZyMbmmljtOrYMledHzGXSRwZNFxR6zFms
CI/3PTOmie4RZiE+VxcxsF4ljsQvkwT89gi5qHjBWKRWzh4yu9KaYxL58b5w/CfBVN3uRrMbw/W8
7DuBG+a3N1Ir490B5KyNilfluPiTrs8Sy21WXfAIK63zdTuMA69m2xOWCE1V1LoZVTJplPJbY5V3
uvbJW9h1QvzelCZ6FOG5KvMSK+9ShWrK24G/Pw74Cc0/XQuuIHLXGaC/IYUnXNmqVyg9nk+X1f+B
S9t6nv4VGCd+wwNlWOcFa6+4Am+laWq/RI3QVhXULW0H94l9yt7g23l8qqDQd6Ap/3VaTMN0pVRI
jEz3cIui6ft9pUJKJVSDXIJY6tp8gmKN2gCJwYyNEzqha8GWo5QRkY/USFDUuV+v+aOw94Fs3GZV
stJdQGZw8z5SF1fj1b65XVutMc571rQmkhRO86/9PLuNdtMiYn4ErNHa5RqbPyTI+64Fpob7tlky
945xkcBNBUsH4ffJnM0GZNxkoMy3bkY5aBWHMH6X2AFz6IrETxdmDE355rnc0ZO/+uhH/vcUvi0Z
pJB6abFlGL+Hy+5dO6eMOC9fd0IycJDsCjTjqvhnlB//EpOxE9zOMEj0MWdrQpMWD0c4UyP2oeR1
5BsMECrUMArJNhdTTmaFNy/b6AWsjTFcg4JjhteR6lIyLed6c0ga8U+LlCRDVmf3oNowLEdLaNAV
AuvJ2fvuddx4dXAOpnFsHvyZrmqtfZ1gMbUhSQvGhkvGPDTS6zOHmFa2mYf7ZbUCm10XDs4xidsK
Rpy44MUw5w8VESAWg6t4+G2VIt5rOUpHvXvol4dy+ssjSL4F1EqN5h3fljhUtNcWYW5EIfsBGZ6H
LsYJE30jS11rXnZ32oVO4jYII+dXCqo8S2o30qJZ2BVjCqQkdAwAIIlqQeHbi/2SQbCqs4C7hZQq
7Oo3Iat5JF3YPg0U62b8DRXvbvq5UEzO3k4iutwnqU02jGe1UVOUY1NOq6f0UoCMvsZ8vvLrOCr/
iofThwtar+QaJ1JrIZQRgZtZ9iNfnXTsvR4hRLe8DtU5nM47twvdxrzubZtgyXn56utU/E0MdY5N
G4/RWzWNT2hITUASdezVkbkgFQ+g1O2j5Z8UtwtDiLKvb6OPaOLK4Q1nduv8SSEwCJBLdyEAgrVj
dzcV9eKiv/T+P10TLsH+zqNw832yt5555PifuEEuPkzBCF5huUygPRyuL2oIXSI5E8E+dWo6u3jZ
pGoJ/VIIIU2F2A6Sy/1q0IkhunrnNqXi+JydFw6jNmkNWnO6bcQtg2oGpZS1PpW5FC3/php6WKXn
AVqM0NI/cn5HBfIaveB9SE0JsseLEJFnVhYJQxp1gAaHRwn2IL8odYZjdoJK79znlnKpUemjcHdD
feVi+nyZKA24bFy8zLvC0fN+M+zR6hM4SWpQlYXptIwZ2M/FY490rxZDLrL9j7o261icCyJjeK21
i39R69SktdWrw88y281pcStISZX5D6YJTnLNxeapRQecga7FNZMlUv3BAzYUNgQybBUt37qLO4A4
Xqh86oA1eeHFg3L45WCzWdxzv78+rLjzxIwjrdYG1HnSLl8IX59PN2Gd7e3mMMe6ijRdiuZDLORA
IAUtz85n00uEV1D5ill6BIzM0RI5eN34ZfDwGSTPoyHltIwGN7peG50BllTOtatdOA4j9ObIHAFG
55ijlTWYWzQ6HEBvXe/TJPFhQpQemFJ0dVPDOqJD/rr90m9yPHOWoyDqu+wXIqKr5tRDCz+Ljn5q
dNKC9Mx3V/puymN113v+d0EgFqyIGUTReHOpIpHRjAKUTVuAlmmWYQIki9gr0oMVOfUQ7IxIL4K7
wnY+MZQIxvLpS2Wext4ptZpBXZWyGv5HRCKQLPZEXCr2iwjVFXBmHQMado+gXqIw9o3zSRm6r+V3
VcAUUpbBBFpGAypwHoqdvijnLPeowET+x7lDIFrhonvbnHSYXcky2dYYUeKhxrejg2utJTM6uR/N
aPpqvogpUdVeOcySkQbCcczyWl3RvGDtncxYOjVCfL81tmpHH3bfNh9AXoHTdSQLUdAxnek6VqxF
RNcaddrvmodrb+F5ngYSIRMsWaB3+GWDCfMTTYRG9zksRpOlywwBqcuMiOseHbvp0KdOIDe1fJzy
+EtzStt4Amn1HKnBJFI5K3ksB/ktZO2OQs2XArUK0q/DvXb+wia+xRSjC1wpWuLYUMo8y8ovTmr6
CZH6G5CMJWDvUQJx4RWBPDIokEw8oPhkyEvVd84BBWjNOoYGqzYBEVy0ebyWoiepk2vQMl+wdF/U
La3w0NR8EPiugcvu9jbigN57zgO4/N8k+Y1excwNpnLIPwnnyzN863gKqNTIec8BrF73otAdoSLS
ViAqb6V7KKAdJ+ywq0xRO+HUqJDjDAUA6udIbHlHpXMxhtOPJ48YHocupln1qNcDNqb1meYBt4Vq
O4aOgNiCoHHzJkmMi+u5VJxhBgP6SkjlaFrDN0OLY/mSk6hAqnAj6phhhvkL5R2mbOSfK5y+smWA
zN91cEwhABw6f1brIbR9KD2oeE37+kpRXLVo7GbJwDGokjg4ipneHNwXDnv+6uDw/7enNadVXRf3
tH9lfUS84WlFO1HCCUZoQMBCCtBpkCVksuoVvq31wNTFDR2CSsf479WtXLjMmB0dSscbWyifBhYZ
iKz3THmQm2/A0mJvL2Gi8IDUpY4jybTZCeoP5ir1sbGiMWQDUqpxlT6B4gfCwalPmBy4k/E3ewrT
aetlUUK/T22KS5LmrnDrnU5T/cus1UYH8P/lYjHe8mAdvSKlgWFMvbQHzUdvaUNhYWA2WFtvhZvU
9sfAX789A6B9Lyu/u2e+ynout8Qlm37a3r/TR0UzHOKNESUqDJxDUnCUHFsfjcRvia9nMvk73wNr
1+i/tqwoakeMjg6VF4q96lVH+0Mzzaqk1PJ7dLnSlrWiH/vu4sx6PG15gDs6zeLT3IwiXx2pzWTs
6x+LoA+HaZPMEbG6xEyXcXvdb0WNrOnywZAo+uqZHjATgh1WycojQBu6Dap71l/dVEhGIn17p5yS
AJ9cpk9Ks4I5NM2tNG/OQ6+JygycxX3UpyVGTdKjKjqeHJ61VrD2TOPQbbMD5iPb/MzPXV+T1JWn
6ejRMJOeEPzbYvmunaMd2PQkS1JBQceVjoNIzBOd/M/Txpp93ouxA+24tQr8BZdxxMwnxAADbPFk
4w95P9DEIYoQmmMqqB1iM2Jn3cKEp4xkXc5ACymEviUgRhbfMQa4OgvD535Tk6wj93/1lCAOhNLx
G9NrzI+44gig0P7WtFw7+rdNSwrMWqa38UaKN45f/DN2aStIVkQrrTIT7/rYMAIZyCqLqk6fTT+T
Mo/eXSVSisX+WLBR7FQD9R+dJXJ7b/jBCjkvvWFM3DPEsdQyZwyUVDb7AO+FLme3DkickwGgbULq
3QaWtlMASyO0nZfsIVwM5MjaJ8R/8W3cdMqkPMpEJVs2j43pS9rTeXgjSVout3qcfjnBHNh9H5JU
yuXCvVx0iLBJFh0HBmXmWPHkR8PO5o4pA8Lvizl2ZQ8IeLyn5ZyjyKJQDDtNdM4Qe4RRcaVJPxbj
Xo/FovndHYG3WmF+mlrZaxJvjcF/vG+Aamppht1U0V0WvRUcoYQUkI7s5IbGYfk4pgMJcDrIiBkn
sj2pGamrQ1QRuHAI0rJuzCAkiyuzavdEfD7kgkreVHU1wNWzy/pErQRFWSa0+qyyGWivXexAzeFW
EuLwTQ+lhsWesomg/RiHH4g/9eyPRdSqz+xani0+nvdUXuN24qiECGV17rZfpHXYpWgUPrayiRJ6
OwSGZMEOZZ15fEcVaWzQOcV951BAhd5iJso0e62ZCHQA/sCHiRgOJ+zXewFuDlG4dS/B0PeK3Mr9
a1gY00iDTacMcVQMsM/iN4EJJBWQ7QHfcC6MGd4GaLrSydo7lOMqIGdsCCAV8cQZmq7oOyMsc12J
NQ3DCpClp/awuiOkgoTh62ZxeLriC1BR/5Vl1mzSDwhH+mh6wNRFQi+rwFmNu/koATpVaR88PZSM
ee0oFqUBomSo+ybBWw3GaHZdetVvv4/zbk9Vr2DS2xxXe9XSLc1sby2xvgHnz56WiqV+5hFyz6kW
no63m8sqStbFhGc4Ff7PMqfMVuJMQTHyqCOrVziVVO7DxYEnOhFHl41clO4oqmguT7BZ6RDg8bfa
rt7Z+aAOg6ga/7d7QNPHTVV0n3J2mrYPPI4SIfHR0TTbC3lwEo2bimHgMZbB71nq28yTeSB6ZSp6
s9HHjTeEW7v2JymITcvkWW7UjOHzyFr0mqTxcxs5Hc8u6FCj2ztzK/EjVDNB9NmVV+AsVbjae/MG
ry/BHgbWyDqXw+U+jJcxoPTFNQVsi3ebdnbjoEH6ANmyj08zxWwrKlWum9kzBo7sESX4FCcToy5o
syR/NVO0Xi1eOWcHfivxJ82lwc/OYSCkU0LoRYW3ykvpstLsRXU3oiGByapGHB3Y3XhQwaaNUBz3
CvlUpvqOw2YlzURXYduJJFMYiHYt1o7dEDkTen9xXd1hp3Rnnn4EJXran6LOyGG4zlPB7dOhLWX0
7Y9V05UWooOGWsJbYLqEdaORzT+4OG0K+q/qBNnXmnRinezIeNMwuFleFnPkkDrjR9LMO+csAXbj
fmy7yy1gJIShwCpiXWCKDvc/+4v5JAQ133XfluWoIebziWjkTYdjhCZFl3I7u0kwBYUJSiP40jua
kyofgeiIoC3uXXNZMw3OAy8R4VL67BYRWZilv0FGyfSA4CjnZiUp9maN0+0bIk716wmlP+5egtSZ
2bvZ480yCABM+RjAsLQv0io7SWV/Kk4vfm4atk5L0nrgKOcsiLnY7f0EdAF4mU5l/xVwT+IaMLVj
DyKA21Eg2X+mwLLL9xGsOwoqZuDCA8E3ahrQ0AL+O0QZsQfuahlgWDynB48hOyHGIHvI7q1aavO1
b1ed+hJ33Bgc0/b29RZluO3EOBrKg2FE+kvAjoJF9ZMpfitDvP6l+NvZIPsvX0R5Kta3BSUssYL1
5z/QcQH1sbZJ+sIw35wo7zufU9VrvfysIoavqy4c/S5mZagGUP56EdXTFgmP6Y9Vu4X+JtjNz6Fv
WAJsBvKPMKkgb1exK6See3JXe94gLgUz1EYIg/G60Y8i/ogWSvXW0EvDIIivUJsaoeG1jlhMzokV
nvhiNkRoLv0sTy6kis3pPKZrSe7FO004kor+OoHruCgIY2/s12tF5pbsXiG8YMj/OTT5SYFfG/Ef
rtBxTVviuSHxOlGx6UUsABIdLEoyeUlo8BoEuKhT+zjvx+aojX639yIsHcEmMWb4ztAtJpTddWUI
jw6xuz/deZGzqb6+2CiNzQcfVHBuDJesmQtB3UlAWI9xz+kaUsLjz1kJDh8Zn2ZRbQdveQ/dz2G3
QsbV5UNQg/yVsDPXwaEJgcTM7eQ/UGIU0EAdwVvLtTFQ7kzjvAN/dM6OwzZyEJo5v7rvmBZNnSo7
5OfrvyZ0g+xTMUTeiIcls7Fk8uf6nkvoqC061SGNtRhkb6AJWmrtG1jQ4vO2qrkbU17B78dHqeRO
b4z8tQOLwtotEOdLsP/w5NfGltLbbSpnbQ6gmY4YaAnBocUTK9+BOgyQ3O4ghrbzRppgKQnk9j7u
hXLGevBaJflR0O/DEPEyhyAftEZK//GYFTRX+795a/cy0ZuT+6ulR+Y8WoxnNKnaXYb6Co5jAG/T
JtNt8Qfm5tcbknbtKn0q+RRQhTQeNfhR5f4j6334l9I4NkDL9kSTu+kcEGzjrDFTUNnDA4nut8dW
uMBYAtYLkmKyJPwCLmcFbQp8uzmIYvXJZo2nOWFpUyjsM+e9CXixu4uH0B+hDsxJoWdXna2r979M
6xG7RyUfh0ZbIBRUzk7LP37xkkjFA6TpeVwr7P1lmEa7vGNe4n8YI+3pdmgQCiMkIPC7y/BiDmEQ
y8DRWaaju85Pcf4ToB4B1GCvhTeFsiTaErsEFuc+Sfuf9A5VA73gFsT0FGQpTs99XVXjRARe8Jk4
6jJAy+66PP6ubvO0fS5sjJOr5kKASVC08hsp6Zp4KXl7d0RuoYc4V6I8WKdIysooR836BzLXeGaE
tK+jD6QMGHTYEuKy7HZf6F096AaElheUn77ciFEnKdfxReEcY92xai0wW9kyJkNnNnSoRTkAOK4O
5Qx0W1ErCSNI913CFE3MIJCiNfNGbR8q6g6mEEYfgywZjfr709luiKPLehjcGNnayf79BtNd//jj
UhcSMWbWAHAIgQb7RieQTPB3wjnz+IJDvKuHC62xoo4Ey5WoJhBvn70odjybQhY/Pcwhvf1xvw1J
zgnIna0npM4cfgz6hN9mTbX4OVSGUiHRO33dc1voJpo2rhBr1AY9NdMhaitnn6RPqM4vLYcI7v/f
GJpcRdtb4G5+W8Btoj1uVUGLJXt2BK33wQpyzzd/1WAzTmcyz2oYzpE5gWjZFBbksfONOetxDjwK
q7zKO7d1VG+nit13RIFPJQoz+d2y46h19X5DnXFqrZDmVgpm7XA/c6na3mEzptBTDLnynkUzi/Nn
98KRhzwa+vNiWdSz01H+KKyVTexr1Sxewd1S1M/01BwpaDIg0xFPrKuoTq22qe9yNZcetGANCTc8
8k5K3OTpFueDq5bG15sXGkMY5yMqY56EJZB9DVoMLiPVaZSVF27AsYipsGEGxmyk5EA9mAJTjeFS
Djwbv1T6CfCJQ7psBvWLk6+UBELbiC84Y5o+51J2sqTlWva1UJ4JNyUZLuZkxnjRau9J0K5Bm5aj
MHEFKLeAQboTqc4BdQpwcy51IW5gfs4aEbII0hotnqfGn6KvftrA/adhLGzEI/q3N75C9gohmOzY
u8Z/XXc4wgEFP4NEYAjudmD8C6sKsQuksXf8UQtQoU4tbTFpSKYEyBfiUCel59CmmAadTScNuEQK
uj4TINVsfNhLFWa7hA5OnYareJe6McrfiSMZJoF4XLru1sZKUGDtMjc+MsWChEMU3lO2f4P8kGGY
Hq0IdFa2BLiABFYftaPX7+zrX1lAqe6vzwZUQIxfHcPChYupqp+qyX2QZrD2pvp1aovkRHC8KJec
OXxvv+yrDFsopqG5zvqsGWA+89p6ORApdBE6eYP2K83csfmjvd4cVWdxMw5IhPGujSNuuJq5ClcM
D7/DUBFVEIufkaQVbeKWfDvHrFbOZt6asNryqp1FWhNVofCL1qjb8dLlBB+wyB4WQUxiDzS8oJYz
t1r5fhNbmxBHO8VN3L5ItSao2PfhNyIq1vnckmzJoqKEgczg4U0Ks/sVkQQOGMARKonfqOcC36Zp
JwhIxZuOb5vCPuTZzz3U5aalSInhrE2oglNBygcyLTl6TgVWabzI5Mj4MIjTWI6/gyHtKU+xluLQ
S9h74c9Wz/Ka50GOs4ZmGFNNm804lWk4QAUkXetZjoeLzM5KgFj9tMY3w+ZWIRLFWMJTVfSZ9cxv
84wyAFQOiKiHe2dQA+obUsPIPpUzCrJxu+ThC3PdEpWXnU70yFKWp5tprIVmTz5EzrIKnlhV9lng
5hypk1FCbzxxRXKcJbojLVA2Q5WJNCuQYJH29vroX02AepE0SFGP4XjPL/k3s8DMScOTUzthAuYa
i04aDsriBcSWOEz+N8q4UTpx3wYaIcuI2c43Y8m5AhREHDE0KBrq5Iw483NoJ8YGsRGz8CveaGhu
FiyDUTVgiwH5a90aVt0FERnwDHxgsAYTh9abledTX2q1Uo7PbBoglFAIbIx3j7xocG8me5DiJAdF
6XI3W0kC8rZczOrUXeVJbztvE7JXWtyzZMXP0JurB0inUYXfV4Djo4m34/Hm3LCrNFhqNjtJgEhs
4mQFeWU/YPeQJhJ21H9gVQdMi+MCFG2f4La2HiHa6fvDcBsB+3qnFLYZB05xfg7j4M0vJBIk80LR
pzpHddiOEhDfX3fTIjoJUZ4dsoMdhbyUJUIMezr9xQMdusEJbx4aR7dwRYwOpMg5wC0N0OTBlFhk
LmkJt/CBJknNFAm04D3Il+C4ODiB6EiXf6ItDgJx4m4SMZQysY6fijT6eDnLNLOd37FAlNJovYU3
VVj+5X6xW/SlEccB9I+WkvrGPvhDIxgstdc+fiqVuzux9G1ctDL0BwcCEdqENbvwbLqv36VkWqn3
EUUdALOHRlzbtrqlTcyVcC3P4tX8mWCynKzWBvIvf5d50ChrG94PN9JsxJyegvgIVPV5p7SobIwg
Qsa3O43Q7yCUhBN82CIXA/ip2KRnJYWcK/9bCFLQP7JY4ZN/Bg2qUJMMoO2OuOoJetUHdBpb6VPJ
gt86kXCtZUAo1GQ/VkWpBKiyJ7VVBbNLqh6F1q8OiEs6UAwSHOi6CeIa5qovsRS0l8Kf7NVn1FAS
ilBNxrrfKtMgI6jdulIdmrGpYPDQLJGs3B74aulDV1ykYgChqHrA2R5W4LkkWcJGSdtrdmdQrSuM
vi4+n9zzBM2mg4b/Fdwic3YR13OI9rkis2Z+qxpSx3/jn8Ru++PQD6fIEt8lIOYRNuiyQrGvquyV
b7E6xYCfwmY6W3uozi/MKVSNhidqUNfXlAjSIM7KqhN9ZQyB8MD+N3S8KgEJuehmuyHqykEymoqz
mdWweYXG3and7MNtnyGb/UD863boJgpOYgCfoTC+/LJWD0TpKRKAJfg6qDgBxWE+ohCIH3z5Eh8c
jFX1spdOMo722gjuzwq8k2s9XBY72XH1se7Go29BnQOUrO/8MiGN5Y4h76RmQC3pTa+megWKwQDH
nLBFuziDge3Ev4Va98YAg0k9Scxq1k5E1aGdogUrhy5oXyQegG2u5XIWVWRagTepDF6nM6KnlmkY
PbAsbNOSeXWiIA7AjdJXdYsIBQ3o+a54rKZjuxM7elsomRRFghc1AnQpqseHoBeE0hI0SNBTuZDy
FDUnpr1UKB2hCDx2a0Zx2Kkn8KCzC6P8WfVlzj86X7VhQfoTs9PQDuICbHtFJiWhj4iKHi1RRFOp
CECpW7d1uiU3hyrxg41GXr5HgaiyaXGj/ZUVm9+c0RT8W9/Pl4onRe07vVTKHDVVfQlHHNYJJouD
dEpTYTEshE8sIDBBtf3SXhIL/ygvmOHofYMNddaZ/ymGVi9u4ZHLzR0fUak6LaKpYwO0WH1s4fAK
27WsSacZhhxy3Y10iJ3OnBnoerBDo8b2KJeD8Iu0gEfjAGg8MwzF28N7N+lcWb39alTnli65arLK
cYQZrH4C3vg69xwwUXad0Vs/bP4FyBEsrgSszdtbI1y2Tjiy9zocAvfO9gaX2T98/2mFgCjY+KsH
rupokDOXWy8QzDDydCYHw9t4Rz5GeOSh4jw03l0M2uO/MDvakE8HPm9C/bX0i5GIxrdoxlVQD1f9
zHLgP+5ZZLUvMlLLdiY+k5buoBeBs+GCjLSPQL0YDJKgUmF/Y8jEUb1Cwi5Hi6QIPbksuIsUf02R
fkKzsOdWocpqWWjTF8hVF6mPWhWbi4BDTxdFeowVjOhVX/L3IU2V6jsJiZxHMGumSug/tAXDrB2R
OqvvqnY3jbaenERQFDR/clo8MMq3i2OGdgkCkWmiGH1zOncDSsjwVp94c1YMfikVVkDay6Sfu6EW
mUKjeoisL+g81kHKtTiAEEkTX75sgzrkuhU9MSTJqt2I0x9P6B6TaTRmg5dsFK+ucFsUcf4q0wBW
Dfq2bs/AVCG6zH6LW/jYTLjKgS3MC74+mgpOALZ/nPN0M+YQM96WYn2MD1Qz6V9n5V4goOh/niY+
9qQvouglessK4keC1vzZo1TuzL7Hnsd+Hyg0oTzKefiPW60dbAA34wE5+k0m/Ct/cyviga4o7jYZ
IkNGbe4i0LAFCerA86cnxwH7183QlqK0/Gw4JWAe3d5IfEvANaK5DsSthYVHyVNQxqnfdPigjCMc
hFuh2IRGOE1VUjCEt9SMpoH8/GkdbKpczbmktO4viknnBHLfWkMheOF575lX7LX4v8nLXimHRgsr
1meHfGX/bSEMZctzjzNtnWBTO9sM0/FOdOS5mCW59F4cK2bRHdbd1Gz6XZduGLBA3ywkkP2i0x1+
OKBdeMCB7KUH4GGBJH3KHzhNR9bCMKrofGcE8jJRp0f9cZd8QVX5Qz/eiVzx31++3zBfi39a2APv
571rBkriYIn2e3NlCaRdNyo38cv1wygqCEAdNLMs1TFhBzEqWOu7oc7eaHcqjg5VeQpkYpnSS/X0
FXO1jD/VQQ049fWYiqPaKec8AEBmzeg20loaetEjvGf+cZJkM6gX0e4kwygaWcGXVNt7wunsTjZl
k5GVT1zAW00bC3JvFOkPmh4AAOuPWUb5yFJzVPI6O9XstSBlsf8V1RdOv/Fwi9eH1L77/5/To04d
flakW4IdpJd7EFXrruTOjkwSJdE7y+yu7QqiLeI1dQkDDTGEWU926YMpPdHujU74jLT/ItmoVZbE
aQbSf80kFMyZEvB3QbiPOVdU5AcuTMMkHqQ40n48J5XaBJrjYwvfnXEroP9crvEylc8dS1bxP+XX
TvIiIVwRfaH6YEMVHokddsWTBs2J6aPu1Albt4wNe+iV7lwlQavxKO0/UX79nrwS5KstP6Wvt03L
t/+fYmh55OqB+6IK53neUxmCWI09R5PrA7IjzQO+FzVizAjk9h0+hJf0fzKrs/V1s2FU0OzSmvgR
vfMQXuhzVQS7YEhzXB/FV6lBsBfKfy77LDY158Z/3hU+tKy3zn50AKwadtmkptfSzyWjelQiVAKl
mAZpxsVG40zLawfLc0nEitudgLtR7kUy07E/CrG1ibIUaB27i9WiufgrZS0MoNItcZ+10VuJAB6t
/W0VaEjVXPFkbO3yXLYZOak+598CzKfgG/qom+5mh4HsCBq8OA3HWuXaZVBcGbF0yUKG2nyTXv41
kE5gOkGDrLZw0T3eEmbXe+S+9aLM1QlGYZSoupZRNtzkcwwonMWOWlnD/Ytv/1K+bJ4kN7+CFmy7
zJmih0SKEs/zx5eOnOxobQl+4oRiDJLqgJraenfaAXp6v1BRo6gyueRhcARcie+Qz2NVgvAdwJYR
4Vpi1nXkIMsSVCrfUGsVfTtL964SaZGCcg5U2u7dguj9iyvjVXt17P6jFRk9RI0bOhlzp3WEqn1T
oGruEmD8yOTUKf27mogesYqa14yjVFg/GZLU8Gjg3Nkw+2tvgVH7Md1hjOR1OeN7XR+Vcw4VADRr
HXKCRQanjogq3juGwxlyb78IJpo2KjsaB82I7VH6ma8y0RP8P0HZbCI4c6rTyxOwOHdptO4ntQFc
sedPBBdLc7ncSKEnvh6yy8IH9KiVynGSdtkihv4T5uUpSXBGyOGDN+ezK26yBLYof73SIeTr/XYI
phy8RvLeCSiB7AHzRmn/Hi6nIE+S5J/tjp2hCwUpq8Ab5CDi61aROy0x1P/cc4adHTFP8xEEE62m
/UJ2E3qi3QgPw/ANgLL/w8RdbYw7IDAV5GrLkeDEFQ8pzJP/4U6Jcq9wNPYwamoPDMAWHHmj1uWv
mhxYjjDmPggxB+5Y018u1BXBxtfcItY38K0Y8uvsRzuamKuMW5Up24x/gpu1jQSs5Nd3H2Uq94Rj
C7LNu3J6qNycJ4CivPva6VlJ1/GuAyGdiwrsA053JPIK+mCqE1GbIPmGQbA9m9ib9CiOd9w1SNQq
FjCQ/OZeg47ZTlTRBzc8287DgeA4fajUJX0lunVUXnb1ModE4zee/hGrpIQ1uQppNCxtKLAfnJR5
yGgkc+Qprp+myXgIAWt6d4NuiwhLSsnqvy7HQ2np9SvGrDx3HZ1zDtiGjO34sDMq3z69fNNDG9Sa
+UsBCjG58GbbNB8g928nOgpOFHs5nExaO4zj6tL5AEGuD+36CoNvAFcGGJqYGvHTVDPJClcN3YC/
UzgevuvAGgYJX3l//QB9uNJvelrzEi/EvNBioTEJ81PIijCigW7X53yy3B+PsUUtVgisAL+yEeit
9/tb3D2IxXNviZ1kYNCS5gwQ+dDjyRIl/JP7aBFMVajpDlAXxRl17ggI5UmGJUtcpItD13VktaaC
z22C2let+j+WWmzOVmw1k1t71mUE+9FnmUBTOg7tGZkpJZSuNHDwN0gZZeBkWKRJAhTljnaDQe7G
2qhOdSOrIh8eOIEhS3KOHlf/BhwKxp8Vr0Z7Uon8JnBJsxLkfr4yKgptrHSbZVyQomTrH2JQitTs
iujFNu0qyn+lfBg22HUZkyiEij2Kk2HlBlxc0Gr+GhbD0EiBLQLKK9Ub6gjnoIIUKwcMsBtckgVN
Q5hDpvA48HM3mhG8k9BDczHLOlH8mtfR97I6roTUIvBq2JIREMGFnWS70YZQtG4ACRPtSVSuxsX3
UkLMfhuZkfkR8PL9dhCzjQZP7O4ULAdupSzX7WzVIPDiH/Ojv2l9eJqCrtoPDYbGBt6OJWEqrTLd
dEOW6b5xrzvk33JjEZECI+kfm1QqOIRoCmG1x278rJlBG0oCKiaEozxKyFhVoA0QUOPfzCFAXo6t
2X1wcQq1+dUkpkVcripfgkrWLCEtYOibBREmiiKxzWtXvKOPVBiQKroozs55l/MrjewnoPP4KqTt
S9ty/bNFBOpfPQKh3DCh23z2IvEGckK5pWUi3KSBnGGxFgEL659EIZuKg2tftfjmkHM+LPnDLtyu
uDV57+nTqGKkN7kzfctB59R1dDxxNoTVhMGOcMuefmOl1VixHlyIzysy5o9NU/muLPI/8NO+Vdfk
8tx7gNIxuXtEjkaSd3HVwzV0QAjZZMUaHHbNBVDuXYAWwlBiIsOSYbqBqrk2m/ZR/fDvmRJWyh1h
0XBsPCOluWYAL3unhwUWxUe5iyTci63XPHghYATS8/baf231VIW+X/SoMlyghcRYTKsQ9pKcun+r
iTjy0i453IkENIyS5axowzDZxQ+mxHCj4omYZQ8cBrk4DMQcAp+aj2KNQ6uuZNpbjb1w0qbB/Xod
tD24ZlM4XOGcCJEt6U84rWkmlzZqG7MmjAb74uQU/th4lzevnkCK8Pqj7IeAnXqxyJBy8ubTRMth
fOSRVRmYsqJ2GAE2HkGibuKIL7qJZRSC9fQvKkgQOFIIkQWrh6pzlHsuXHIsYGlifdY6JoUogzPa
8iY5LJSgrutvsVr2yFNpojqvFWmO6B1qlwSlYciukYLuaApkqybkmHPeXaHhiMnKvieTnPtcmImw
u0D6ylJGrWUFlQNFxtuD5fd9/EKj8AUcZEaM3cdte/7XqGqMb/VwUPJGoewpVb9D2t5t7CVCOi4V
8Tp9Lrgo7bFftu8jdjLULv21qclIy4WZfn7egUKghh3DUnlw8Vk/ymmSQcSQ667m+A/L7pYf7gh7
oMvijklkLPuOdXlxiBirGbpAdhcV/XfnNT70u/3xaioEwmjlaVMoP3qxcOJafuzLweoe4Fo98dZE
E3VK9xJl+Hoc+9opS/92njJ/yxSmMhOAMed4g0AgsdlrgLLWJAlC3xhNgJr/lWeyi8OWMQLUNnUa
49hqhoq388lhh+4NHCU2mGcNR5EEnylUYJWBjaLv/BwjeixJKz74qAB+86J7/fOkTHqce/Bn62k1
w/p6CvlN3amG4ymM0faQvEMT1S7i/GbSfPk6GPaW3V90UdkiT6jjg9o4U8nMtzx+HuF8TS/mCqtP
GSZD5Dp3AmOVrBK+o7gGOt5XVwBAcsOBSejKKkR0FQoblEhR+O6jyE7fECDN6HoA9fRWTw5FeuIZ
RwG4EirPxAHOiWGI2Wm0mS4yCwSox06lk4gdJcdbhpVpYkVVWOoJ6LwvGxJBUyGhkygN8XL1AQRc
x7uoy3ylpZi6jph7SK/umdTeZ6du7A5UMXJVnPOLmmwg5ATQpovwHrJBxpWFwPH851d8btam3okT
EMhspPg5ruKvyosmzED2GaE/Gz0hpFTDhRQ3zNid4trthJ3uRO1WDyhO94IFELIi8ElR/gDbGTXn
hQXKca8tmY9W62xCMUAyoBtpwTubNDwFQOJe8+l3SV9MiTs07M0j3E1I9ATbEbz/hmRjqEw2BULU
k55SpW1gJzCnwB1vmwK8YdD0hhk9k31nyZjwkhfSBqYyjM3gYN1fj7KQjtaefVigyccq/SlKAiVy
OeneDW/EL0/0yZWlZ0AqaU0Ta9Dgb1vuILSQDTgqe3tLhoagy32OmIiCE0zK2okrJ2HlSyrH7+9e
atIZfnpf7euJ+Of3l0rZcopoo4ZTMya5pzCmr+iZatHy8a1GJJDEerAunJAdpxwtEKRG+QRR2obk
7Eseqs5oeyLLpjpsp+9mmd2M7DUVujmij1/5wNJIFiFp5y/VyhydQzrFpcPv6slrNxlbtWEpnzW7
aQl87EU+ZSp/PH8ZAPUx3bdeBntoUXAd+69nddRvSJZYf6GaUUpwkZ3s7jvqBuoaWBIFVI+PncR4
foA4KILcz8tVhy/4VhVz8TDoK7GRnamJ/iNoS4SnRihFKbjB2M7LXzxsHcFioX/xehY0CDhx3DcX
MDfx5tF5A3mMH/LZcwb2JDiaK3oeqZV4IjPdN1eCNWZvLTVHe+n+hM8VPyIb2MV0Lq8W7kh4bsuH
Udw8asaD25M4dWqjS49k725hV/gZcOgeFLW1Gep/z4IP8Zw4tpiVk61fv3q+KexCKMgWL5fn2JHm
+nx31C4mnOIERK/9Oc146C2G3Ct79mWmqJr1xo7a9/ouHY8V+9NEH/AEtPUGOw8Yjx1ETxkffNr5
pN6cspEpI9PCMHR1QDuNI0hlu6t/sDeUQ25u7jw1mi7D4m+fMuJQtAspfZ6K2AgMQYVoKpE08q8T
4wvNjQypxg+icg8GocIx4HMsu5kd3se9nF34m2WRXYKQLrIkHlsYg7b6By+l9v57dj8X3DnSg/on
XX02l7lbQ3Mp9dViEjxpIXoXzTxMvWd3QsD8LBm38K2Vx2Rscju8q1wbI0ezGhI/yeolp2UUyoSL
4xiRjcwHuldsJSM+HHbswOyP85s3+83kwcaQijQRc/dNkNC7FKk6vj660Mg3uQFm1mAGmClX25dW
trutubs2aZHpsZEsPut1hQRXjKgoYugspgLVWP4wU4uswo2H12ThO+ertDcmSvzsaiymb+PdJrq4
hQZmYC66P5agLqXUGnWUjSP5C2EwyBn9AG7B3v/lBnglkADtyUdArAj/Z6hYyB6FNu9FpHS4OafS
Kx5TdalXTq0o5FQJ/kZgLkvscpVAu4fULV88Gsuy6WciEA0bhdfANMEYKlwJWSHk2lDuZ6fKMY5v
0OrhwKFX9+4DOGJDIjNE4tO1hdokPwaI1a7gY5nKL4TScORdP+A2VoTgI1CeJAm0d2eG5LLNw1Ii
bI1hCycYY2O/7h2VqyVL+689dqbJr27BL592CuFkFNUM5gMMvjkZAl4je+JX7HLjLQUf9fMpinyt
1Asv7JjN4gkOyPyw0AzOyPGcsnVW/uG2Dxe3zlHUbbiFK6kRHY2zzP/T46xuEcvD5Ak+j4VxzK7B
bdEJSrntqoKGLdUSvOjYLIWdaIPBCzhydFYkdWN35R2n4r2oFpkp+zjwwUYqNMFaVvB2JkAx5SOn
6X7un7J0wHYDGU3IVfoFNIvGiyi0SQrvQ3qWqz2aJSKYLGF+tIzWHGtqpfLN0QUw8fjIaXy/GW1V
OiTiBH9fBW4MdVal2NwKupvqj5fJCkU+aCPczgcqV+sy64YIfKxjaH9xHK33htoy64u6xkyxNyu4
vqju4fxVI3J+QQC98j59oR+fKx5eYILKvN+pm2+dExFE8PBWVYYiTj9mOTsdRKhkpnw0I4UYNr+8
PvZJs2VqZKJqkB5cxu2RFNG5DHJ8knswXxcpoLdLDG81eDJhsz8eWZa7wVLXe+PZsWbs2LEL9W89
I/JYs18D5+JliD4l9Ux3Ri+4k3c9ToEtTzDNXdhR9XT94dii255pb1K4WJMi8qCxIq5f8v2kBJES
o+4LVN3mjaaT+o6yW7LAr0e3YmA8Rfj0SITtRaQUYoxF+U4pDL0xsePsWKfsfVouYWGGqihNzukw
FBHbJA29Li5/3B8bQnqu6TuDE1vAd4qhTeN8HNF23wTZDdHVgTMn9Yv4asq5UQWDB8G/bW1vm9Tu
nT14gE41+dgbZ8w3KdoKS75Sv/scj35PB1bXy6U8dfQED/kI5EY5c5BzCmWLEGhWAvMkXuH/Exv2
FJWiBIRiGRQRfRy82EpYVnXoQvemuwxJkb4t7DkAhcvASDWjzUWbvGitIN9DJTBFhvFUvgAZRuLX
W7laA0vOIoOrmoNV9oYLCO27ylL4vW3jVgorPUoB9egzif5SnDpad+Pf6g3J2GRmwYLD7A6DjsY/
uNxg9sAURJ+7emfsa6ioJ29tCtUfaRQZGLAa7M1ymRf6GAK+9+ZrB+rh2fkKA9ya6ZGgkTzYvuxH
vuMhl3ZQhsQJQu9rAM6ZcUoBaY+S/T+kjp+fSsxmXmxPBWu9S0eDwKDKIGLlSClBg3iaDo+KN2yD
z0wQYaYq7QUIP0N8lETt237FFshR4IQSFJ0/vb4jxhjaLdWl2XgkLX2v93hD0T2ovDi0pJ+VSkG4
MC+ZRy1oj/w5CRF3MXTup8UT4HZFoofjskYCQhbQGc8buOm+3aD6V9sUnYv6FUu3x7q0oljdd68s
GjY93iCUx8ruSBq047AOov5q2/d7GNXmbr7NQSdmv630KyPCkwH4TX3F3JFpKlMoqWOCP890qyLQ
XVCwSwFZ1/D1m6RNuu6huvwiTemFKNwmySSH61Ys7kqrZ8YDZuEhqXNS9vRHdbyAPhvkBo6IiaCI
jNu8TfBz/dV1NMNPdLIqW23+bT+D6ERN50/R1cjnigcyI2WqkalCBhIOW65f9jm/zf4pP/RAjbUc
fh7Zwge6IECUXxlmAxR/DnhOKnACQbEsORL4c2PfHLwYYuq5o7y99exKZOABtIHBaXGVmqSrUaZc
gNUdmacX6f5NLUbS6abjY3AcWLPGm0ZUWbPfBciFwrtC12OT8xi/qkG6Bt9h2yDyZO9bxYe6KmbF
UfftDy9MnCM3oyzS0WT4yhz+HGiGiHvdDGI0b4JCHQcmg5gtRgkjIiJ01sIzFUzBWXvMpQV/k5sx
OVLJmG/Hx0dG8LG8OHwCHfFjhSmiovmMVzQFcDH6Yh1io1PGMoUzdg/n6MZnFe8FvT+uqv9sJ2ky
W4LNeHCk/vk/l2es7aZVhOuCm7mE80WfVgJNYUsknGD/7oJ8Hjp3AGTqXetH3nfU6pV/2tBRqQi0
lezWB5ODGpSwVEcKycxMn0x5gAVCr/Px484PHL5H89AB78v7PLbHF7/jq89Zo19Np0S05nOl+xxD
yNPc4HFE5Frsbti28p/VEaLKa8ApkzicmIPONp0pLx5yNy8M6EmSQ3kTFMB0NBsgN8nsDC3Ma8+F
6zB6ZuwF1sH+UCu7tg31Zt9DztfJ0u6KoDeLFUHra8hX5hP/LhXKnIr0yj9+fYyZawO8FYEjTrLa
WOYAMQm3eXoPVHKFFAspD6eB4jvtmUra8ZVVb+SHH0G0HcI/yNh93xWJUPNEbswjp08eDduHaEXy
4lTyAx62jPte9dxA6vvzKQVHi8s5NvV3HJcHsofHTEpHw0LUU5uAcDfS5VjNbl1poYW3plms4Gc2
2zv/wkqiNqoaC7b2w4Y31MxXKRugleIcsKVye6u1l33l2r9tH21ueGnYjetABEaT4Swe7B3CcEWj
jHpew01SYbWAjFQ3zngp28DF/djhd2pfsP33x/DFzLYOpo/36wx6yq9KlUTf2JOsLaJilHzRYF/f
tzRnjrSAuTQYk+QRmWv4CRV9xz9Bqc8tA9bK+Yvxr82Jdj5qg22UHyNrFQFe6ERJwNvcxadakrx2
XzT47EJQaaJb2vBP/RZeHMZrzDG8GFWBb5q0W661EfGMPvv8cIOd4vqfD2X6u/TMp6hpMxXypg2G
e5TodLbtOoZ5CC1E5BrHrsHRRpeDJ5cbrmgqEWZKqn2EM5X1qDz34tWTBY6u0Mva3uWRNBce8dUD
FEVNbRq+dLGgb3cFfO8fucdVd2EmfN7/HwjJtNyCxWnp5zjyTsgmSFb/2+CntTrouH6j7jkUcJXW
8rzinjkrvWLMu41Mfb+gOsc4Wy0lhEJIods/LycTU7Hp3DxUwiG3QBEHSGp6cnO+wb3LHP0qOIyM
iCzygtunBo2+nwypPz1Xydpx79ka66zwoBvvfcK0WiqAiK8OLqf4kCZSBbBG9KhTEB/9oBll4e9N
EW8bRAUrsEl56BR1v1m2leMvYv+LzZkXhLCweSxyYtbAR88yr7V5REObPHrr4yDGdvDtBTZDsG/V
IkF1Lykk3pEkRBOqccIFj8RYJRlA214WC599J/j2KmOsFUbU7fBEHazYB1ecowrZ0vsFbvRoYsay
b3BjwX+HKdMifPCDeFrYCUF6Dx3EgZZFGKRFROV2mYOVT0ZzMLDDknOJq2tcTAGWCHxBhAKDs7xo
pBuCag3gzUMLabOarwWefPig1R0WuD+VyLF1AmxKR793IOjPQImbHCmGl+gMlzfsr2C6AGIkkl8H
Qhi5GMYbhTdViMQGGQIyEB7obzZt2DJyt9r8RDVApA2eH0f4HyWCb42/5pTJUbSkYNv7P97hzBly
4Lyyqtk59iiXciFROJMyug86b7rU8jQiSfKtlbOW/G/vn6Fge7dxPaDFKwJG11GF9Lfm03dA0nJF
FyxJ/oyV3mHltWjMN2e4qj1zXIXqjXBTQDrwkzz/2FidZX2BT+cn3CGuGAQX9Gs1ZiJviWWHAWs5
N5rb4PkOuhhTFdKVyZcK/jMVgjDI89jIdGR3QJOjlhq/UH4OfwKYd3sYiJ8HSmeqiRSzuz7TnwmP
dKqHCO6X3W3VFyIQ1Rguinv+GfXpTzF/mU8I1McIWiRCebB8/+S50lHpiYBIug9HpeWinzexzn01
tYyoL6moP43vwIigpiAtGFcy6D3KZbd3MFyLAjoMAyRpmJYpnbLVNsjDjI6oFlzeaq56p/PegRrm
KYXjE9v0LPci4188Ql5RJSGmj0eYPWbC9oXqnE1j20i0U36Wz5nyBb1p32lUkbDfzleJO/ppQm1p
elUplv8if28vO0VsHa7nWr7kyCCAlfor/Df2Xxis3YiqnowpV8Y6HHF3HpexDqITH+u7ZmDPg0cm
pVnYPrwCcv5K7HH/GWn5eniIa2rRzqqIjvHu6SMJpmxdCmbkcpzRt3/kyupdeoZyl9MOGZWaXRFm
m8zjbSIXy7IxSakP8o2zM7CwcjR9PySXHA9sILTbtxaG3etwBv7XZFXAqr77ouatoSRi18vkRxDV
3vyh5Ma5It1sNf11kyPelb1+cUxQo7k3XPw8w9J5qOD1K85GEXtjkkRwfiURaEzXhXB0M4gsPk0Z
cB2iG4WKiIqJexsnSeg7Hg/1kJZJFIDLj0+jeD5euuraE7HSkFsG6JdB0vijrH5TTKuPH/KDLJCA
Z85ptSfC+RIbiL3SFh35x+jl0mp58DK5yivINeRQjCAu20Fcb5plnVyzQuzSzNKViTbm4g7+xsGv
OrTCiHxwYcJ2pkA7U+xxJoDmPkXSNRY8ecw2N6UvBTCg1CbQoiah2BVmUQXqONhLVQhRb1I5aYqm
2+SnWvJ/NcU/JDHpo3V8eLDGj3ttqaZPpWLCBqSfzMpjan5y6bSJYS97ibZShylMgASoU9BmW8cZ
oCcjhf/kzD551HbDtZnry20titESq1Lv+xOQoubOWA1TS9mYKWVR+0zPa8aOrHZnz3AqJpFHxbP6
/NJ1oM82gBEKe7W7w0iEm+AZE6nOapka+V8MUFrREHyKna7xdY+TdTRbrsd1CSAXUYzdbLRmq7F+
Bho8U92ZKBka55Fjrcl43BLshBYFZhfYdGnXqKJYvJjGdDxErLsvMtalFuMqREF1zIdk4kh4C1wJ
pNz383IlzfHwLR1LaM5HLBLJK2eMT3ip3IeyBXUo9DUBgFoNrM6K/wlHiNpjSRqMVdB9rMEuP06w
YENNniD8VYaww5/WvVcONq5gLaQ9o9Tx47/aWuZYHjUeBRbZOPKSIF928jWp7f1hr0d8MqvxnMHx
jssJ+Ey+YA5rlUP+jp8BqxpBi6upxRUI4FYA5ziULVAK/1EXr5pV48ZKX/pG91SZ8YN6Fd5UEzAq
1AYrsucHzyWoiZ1OaRnxQ5J2Gw9cDVUEAKzxarrVb5Dd7teWLii+OB4uJXnhRHLncv8fVWHse9rS
WFfV2mrKNXFuhR8AYAUyo7GeOLFcO1YJSucE5nY8ZWJUFaFbF+k6b/XYUkR9unDj86PEvOAAI8OB
wJD3w2mBCMYIDJCToGQnBb0lDBdkuQmIPIlVRSd+BhlofoxC06zFqBtbN5GSvFeT6g98cGjiE3Fb
jcUH2s5O0dl8koCPEMi5UyFxaTxTygsCpZ2kI0tjFPJ/7mCxvtfBLDSfPbU5BjRBKAo4T/AZ1jKE
16K92cGdtgXk/VGiEU+gEAv/Z5voHeRX5Fq6NuGoQjvA5CGe+7n6Y36FKeex+bOhKcXW6iGdUz8A
7w4Y8DRzyFHQ5umeufJdVF77waXGplzFwdNMTeu1RELaYai2MyDThSdYVN7GW/2CB9ZtTewm1z6q
8+WYx6hMMAmSMZ4NqrmBtJeCjT7U79UQYNHd2FJQID1BIQGmitZ8xOPpU7pJZPevuK5om4hZxIdL
9qNaWWVeXrNtXdnRl/9AiLzJzhSaH4WYFf/wnGvHFPw6mqK5lU3YSShSh/Xyz3bUEERaix0ThGAv
CvlLASKXS2k+2ajgcB3lSuotF+CMgJnFlPQcL3NEhHG2TEplbMh3PF1pasnYfFPp8Fo84XjiMCFj
scS+2l2n9WmXry9hKL2/b69vvUabTmXRhMhXoA5s+62Qfd0CpYFAIpFzADiwBB34y9UQMpBFGzWl
ZeOCgxtIex5wihFFtH3F3OYiz6rTfqDk1WkO7K6G0ZZ2ikDhJ5/EG13okzttv/1jwQI4Xffmdr8/
6vK6VzqDGX7pB+6nXFFtQN9KR6Q4vDJsqsMwXWPzoDt3+ugZmOxs1xe2F474Y8CZ04QVf1PHiSYJ
0woTyGi5K1wiCv2J31xXZCqhu0oOdaUFaW7/5OlZ+KGNJ/yy7/3dHH3c32lREJoFC8NiECNtkTSh
EcRwcwdP241EnLtetW2EDOjut7dWCXQiVo2qK6BN4b6nGo0bdepj4FAkN4Va/FCjy0HOq0EoLrMk
2cAyGPUh45MVcmYAxiISmPYfcHSfy710FkEtbt2Js0YuzN7o/lVUY4Nr1kOTlIf/bpf4GShWA0yC
OIDBULtmwmxDbOIjWGW/4isv2PZ87Q2lIn5WYimaG9BQvUlZ2S3kyAVTHK9Ukc8J9CY1LbfYNaBT
rr00uL0WZzVMNDKUPCYTq2SM54fYxGbWysFZUv+E4xiVSNEqogQdydDk/iVqVOGbuC7ueK0DEZnd
5XJyg16Gj5pqTICBfwwk1DKXtSg6trvylmjxXLQ/rjU4QvC0azE5Z5CyLb+/UElPRTlC998xPa47
EqGXtxPZlws1w0OLSbFJ2wU06wNIXtvmP8Tm8h1db60Ih7tof7XElhI1BcKvUkGBYDZkT7XcnYRg
zaZJoTODnhT3bMn3RWTgfn2/GijNnutwAo6VK9wM6OLpWGF5Ah4xFwyBy9i6wnu09QreXz4d0exd
CRe354nOChfhpQzzB5TwoOQ4aue3XpH7pnkpUWZ7yM1aUe2BKXRs6cRv0/5iPP3bSUlBbtea0nYh
SrbWhk3i6qjbSdaWwRCNLxipVNciHwokjgMxj3BgWiNZo0SoEQsjRCkJAptKtNRviwrUrkyqq/SD
M3E6fwUCiNtVbkx/rzZ7WOA5HnS/t5lJLExKszKaFGzCVjad2AWNOnV3A2fyO2Fy7F44iDTUXJt1
U0PTh7zgHNfwyq0lsEf/F7A18DNaes3p/0Hlv8AeAbA40ByQL2v4Auc34+xGW69ti2bxC/zHO89l
gTC7GZvHlK68VQDq6WfQGZarhsiFI5OvCykggRYNVUTscqFplupMWGlKB5odqs0nW1lK59BBs7we
96edj3XEmQNoXNFj+mK3jeeyuegS+Hn4YPbqZYLKLKTXgDHuZaCVnrpF7PGA81M4XGVruGXNe7sv
h3CoXjWuFkxpHdZgfSWeuZV4bDwOjNTivOykiVB1HFzySdpa5hGEE6qqOBR8vgN823YcE+zTxDp3
v8SmgLbvNg29bTKkIVN4kzN4nUgeOlo2DfSGa45Qg1/y4W2hFY/+1VH1UMo1MekGq5/QZ0JeQ8wq
mFuxOtDXIsU0kdQmDiBwH7J5wm76mwfmT8D9aC0+zu45IUyW8zuFYxoIaonDgdu0jKi6mzFnYfdt
yCdnUiyy5p/hbJdXhvXe3t/5dua2d3hBJvIUTCanM51TZhpdgq1r/tCyEef/mqkDLpt/Yj69HE8b
eVOxz/SlDQm0Pje21s8D8sBUgpbskiKH7czLL+7oARX1QfG109o04UP7r0MFw8m35T/mdG1A2QXF
eigMzoSyt+CDh9Gf6Xek5zDEBqfIAbfaniEt2Y8SJyOnIRxYBChcJticiLCCj3sv3bcELDEgntps
GZ3OqIEYp02J4zMDCkE+WymWTneACOS/VlPchQr9CDBZdKfw3togCoU3OdgLx7KVdfJ/MDdud2o9
WFSG8yZy8fgjRiKObcv1+5VJhQxoUDsvz40UzL+8AzCiAwY7rza2ZA/EtLU6KO1cxBKbbcKoyTIu
u8UY1JCSqEcL78nGjgTCzrrJlSvR9NTYWhjzeGATmlkRGGpnHePXNR/Zqv3S4tFshHP4FJNc7Ss5
BjPQwQLxup9DCRk0WG7Oce/vP1SH+B7dVbRtpOXONNgd3awaiaMlLJyATi9N6P0YbaoByYFRf4le
JMSe5asQtflR/t6R0i+0XoFIWTJT+oWWBFuggoo2Fw0rb3vozekU+szNPKxbvdGjF2vWgCkmLJNg
jQMB6YNyE5uuymrNVJuhKWS2Iy8Fzxyp6MXhv8YNd05C6BjaA7/yva2bhRoqE/GwWoDlbbZdfR6Q
wuOGoOYpjmDba76TBq6THPZYl/S1H5q9AKbi+wTTbyPk4MgGbeXUCG0W8hLOhIpEVQ7MRL9J2TBJ
gFtRDduAO+m+9FkmXV6S2Zt0jg5SOCxNffqUuW61slH/Cd6YHIlM72RBqe5JUO4wPztITKdGr9Sh
fAdUSYRAuLkwdH4gIdPCzP/nk5x0NFoWk5RA3R74LT7tGVHKH1ukFU4DENMxDjDr2vi+W/M9iLCu
4OqRF5v/Uhp++OenqhaZrpXaK/qCGTGaVIzRQ/s7ScrKJ0lKcdz2kZGS1QESBepY/GSwfDt3ZRtY
ucVKgaZ3YkkNVmntoY1/gfEN3DAMYYxWjTdicyhs3jBtVO0ymLAoOVrjpW/h6a6p32Lhh3Ug29sE
6Lx1DzQ36nyNzy5n/aKwJ4ATEZlpck4m28rqTONZoelcnWp35TQMCnUOex+ZfkyCmfcWayPJRyop
snKd95fsdDtY2XLiSi1ORoiheJegkGOicxft31BsjdEZmdSaMQ+iDdKwxO7ikcdpSfIeLhO5eW2Z
EKMOuc2kQUhe2e9pXvC4ZL5/j++pAOvU/+1ZMkw/gNvnkECANrj59jfOeHw+NaiBO7WIUAoBZdON
z7vp1yXNGkOS+UsCf0k74JGlhUbCa5xtQ6DU94k8gwFfBczVy9P9LRL9WwkBJPbGM/Miz1CqTPNT
+4LJ6SlvYZm0aOiB9ZAgKDHuja1BGFtktnudNBMu5ie+f45hojGfzoCG8ZQMFpZYiy0HKQK8Y9Mt
tWJLryOwMrST8GRdkYOPVyNrgh+pUavoXQE8/KzvT1Ircg6+bCWeMQF2Sagxbpqk6Wa/wDD41TvG
zJCxRWeJxZKQzV0FrBKfai3dMeCRo0fHmzfTzNsiQxZhYp0u4kls7uLzNT26KTJU+r0Hgqh2nX7r
9Ocjj3T1CT8Xht6BW7axMyLARNVqyUJvffCvOC7QhjxHJOOTWOeLLLLLhCVtWCnzCEKf7lfsbZV+
jdYcSoCRRsX2nciBblqiWcXx8fmYHryI8z0XEV//FCYRFcUQmtNa22a0bJDRH/dx7nTqLRttt3NP
t9ouy5ldpxEw3VoD2mYpByZqJG2hZxDOiuTnBWdxk0pZc1z8thEpGYbK1nVj4XghdCpmCDOHzNXW
O1iw99Uzqx4M7odSYrF+SMgYLst5CHeN+TJ9vrXyqFgs/rYguPmznSam6OZ6MNXVlImgVJ4mQDJ4
KGuXh7FpLf39GbJXXQVJyALG2dxL9GjlsKtSMj3l/d2tq6kSqcKhejiCgWPtyDXI41lwGfF8pLKl
33cPoAZoeHgjordYMvgPMq1zHeYscBZipMv/k6TebUS+/kEmoyYcc0bvWO5PPzK56YwPxTozCT+U
i46dGKOX3vXju8+cD+9dDqO59tzkhlhvKas2YC9FvSsk2IwpcNWpcesaymftf4+JGlMRf7on4xhs
TV/sXH6EVazyASJikgQVUVoddM/1LDYG9XmF+aBPesndO6APCHfZe87N96fOcuo7JcHkPN4JnlRl
aa1ySU+JhRlvM1nwYIYFtDu3u7Bx/jqUVhcp4Y+16ZqwwJnzD86noKFWqaKzBaT0DoZSMbnv4Wso
JVlgqFGi6q98+IW5djVFuWDFI9bFNTfZ4zYG1BxzHAJrkX2o9gsOaw7MjPggj/hfrUvlq9K4oodA
m33vswHDWLFcqGzq2WyZl2c+OpPqc6D+YaQdCXU0OweXwFwEwUdPSjd5IRlROxkPbelbUHr1xiY/
BHp3+Hs3TpRaDVBmhERzhlVozjnJJS2GCSjT5VicM2zdZclWXLcFGgB4qSVDM1yMSlarrDTo6oSb
0mbax00ScPxWxlH29nVE8nb7otCpPgikA8f7YzZiLNA4im1H2MVA3RGrA0CESvoD9tlPN5iRRLeo
ygy6nqF/mvgRTGAJIdljjY22NgBS1AVdl+LTxgeHiNUhldU9CALWnv/7AAh4b6j/k3eV1F5N9NcB
AgYw8rOb7gMvBJu3+aI0kjLuFEKke68VR9aqEtjQBcpIf1vqg8+f0mRafA7JYmhzzgb+PmHKW+7U
HRFfhckp8V07CqGOgv/n7g60E7CRmaRf9Accnls+sfw5NlMDD1v78/ZJ7uY1dtjo4Gg5XxwanE/P
SoYekR8K1fdWZikQuLbcLyHchJ0hxgc4RaVXmPTjescmQVKdQcklLSCF81ugMpFuRPLGxGXZ5UIw
K8zljO3tWYwfYYDcLRoHZgiIv4UQlFeC/CfP41FZkosKTjc9oNoD7dA1m7ZsCgRz7QCvOjx+5lOj
OobwNi2FU1QGHz64wTNm69tujU5tjKxYvlwWojno6WqnI5j6en8MqB8UDygFOmLlGqNp0jryyFht
r+P3Biq6SpLdjFbtetKutSZYu3au9tDgki5Z5PUzihDjJw6l5mUxtcG1UISSIF3tj2RmJKhvl/er
YNBSbRcbIbTrWmLM0g9Yfh9iyZT+17zcgdyl7oRGB/55z89NVbiTYhtyaIWxY7CHjhU5ykT7b33p
vURrC4A5YH4S2Xm2wsaWPKyNcapBjjs5HfXpUCQ8hr1ul5or4UnQaBU1zxZDDBf0b1OGofl+ZK5s
tk6FpZk3idI5hmMksd1JiDeP7qwskFzS/KSsW9BUvFcKy0KUwU8VBT0wRQL3XJ+6goQYdpmyA/JH
GHSco9SdZSttLhHWoOrBG6hfR04lyHbsF3sX0j72y2kSbZ4EwIXKQ/HFHwRmJQel2NfliGatt7sB
0UjS3IUAVTPkDFYpdzOL8hKB3tkvPtO7RkcBpNXlD9GkqPr6rUAYB0fjx/yIQ2VVfgtjcn95qYXS
f7IY0y/NrcyJUyZYilVK8hRKgxPC1xtPguLKU/XVAfJKc+iSt7lJYF82xpsqKx8LnyUwOftlOe+7
8rOr6z3wnRR4OKE6Dcl4RkQeog0NM9jiNabUpxId3XzOfSqYjn0y553SWjxfYl5+B3T6qkHdsYrf
Fcrgwncg2S89SI4MToXhd671Lg3EDoYg6kczvyBGLb8adT9F31lYcOMFvAHaKd3ntJbnSGtJ3zVL
rnVPn3pNh/CwG6r4kO4sXqjkviYxuPzPZuOGePi4zNfJUkEJVsfl7xWSejq31CsPrNPi0CpeDAgC
9ZLnpbWZQFub6wE+/IA531cDey8wF1oYJ/4vCBNg/gz8SLesKT5q4e9tJo8Pf+24HoJ4BxnYNHW7
Tq8i2+0z7k+JQ4N3W1cbvkWpkOomIymYxWwHQyCpCTPHD6TxW9h5GijCc75+odfhqNViaacAE55l
55YACLtM1KBVC1IjeGBSK0QwVHdTv1nZiKfO6hDfC2UMb9i6To+Hb+bd4q0uAU4zCEIJ54Ub7HM2
dzOEHNXCtRXWNB0Y2aO8vWIwrYIqqKAji3X0rDp/TK6SSkgYWQYMrnsDRgZa1sYp6BkAI5ycPI+1
ugLdlRL0h/3EcmxSB14PoCN/IFT6cn61sNrD5jck5AAxC4fmn41ty5W2SgUBPHT1MngB5tpC51PV
6TIrWKVyVgm1sP9sZWt+963GRDWbiB+OMGYYNZfe0Mqz6zKGhNC+Cgx7QRiX4qUPLA5556yk528d
fJw0kdMIQ+O9g7u5ISCiBhBcBXjQSGw1YdALtOTvZxp0mWEDhXXjx4nBgo2sY7C7foGYVwizOe3R
19S0+A9NWCAUsVeb0OZ5cuWh8wzRrqCXrS/aYVVYu0X1h5fHeVo2CJ/hkv3rBmP+vGxvKfTJIL4b
F3dWRCRXFXOOOG4O85FhgcfAk6kQBkDawXYwIpz1Da+GwA2lqo6qa0Sx/99Di6yQsLO2TrSIuSw4
8yzox7wKw7Vt/lyV5wo5+LJ0JbkZSdsgij2FGeqVHSHQjdVnfDpx7bMnT7dVXtiYZe71V4vKWUNl
8KQPqaLWdr3ARH89EYzJj1kMTs8rQZJi2DUhSRHjLx6nOlV6JAEaMxVnapS9XlfQvrKRRPAWxtPD
icCpu1MKv+JkgEtopVbfLZ3boe6iYyCevggkU92rJdguf1t+Ps6xrLWTzz3q3JYChWoA8cY+Fo9A
6M0miwzJXugY2jrRtQTKO6Bc58qx9Z4/kz8iDGbgVu8nlHNGwktOXjzipdQkqk6iayvStt1FwCw4
vYuMvyekDUQfsaA6M9sDDwP8s16rRMZU2cIzgfLyyI1eykA4wcyBrIpqLq3OpDYQmyovkyxdEyLx
CAvJEHQ8EjA56IsC83kHdY1x7M7TmJt4onkSkg9oMeqHwT5N+CMwgK7ukmJPYfMyZ/fT4SbGG4Ec
D2xPV5JseaqVrmu8YxSkh026u3QXuss3v7c73yaM90BzNOsg7AyHC2wBOLIJwR169oQw6lPlmSeS
/5nSE9xnDMdqmpoUZ0pSh7WiNmGNSsbLFAZE2Fw2DM0sdyD+5o0RMvOeZIpMTlszshKnY+LThbEy
KcUKty/rje1ZStYEfY4G0afXS3rKTZklPF/MuCAWw0tT5ZHJ1BBWqfYevRf0B6OdyBRc2rA1Tnp8
/Gj0rVHykHT2DYGJBHYFLmX9p9/uBSaLEMldekioIdVN1UECAurheXzhKwGIwb3XfGXyj2JbKcUN
0Hf3AjEY7zC2RAe4XDhGAMLDyrRjqHVgDIP3iZZxSKmXdZMxsyaPeJFU9iF+hv/wgzpuVGj1+hrB
WJ3gg3Xmq7siYg4hnwsFK6u/3JBxA63lCi/Gg8eTNnAG3tnNpArIHXc4GS/yyurpXCXEGLCxnRuK
8yKFC4DqTShIdR4j3H/iM5DzZ6IH326JKyhPAGuXTYvr4c/ezRfHZP54N1jqFwA04io7zvXfMhmU
lOwqyGOsJnCSCICopbsyiMvHCP/4gazqM+EVMhRl5oxZottWucmzzTdRmepEalM8ZvCtm7S0g8di
FvYlF/t626ALj6VsMG6eR9k3Rp2WmPpMjabaM/yob+T3hLovad6begtZuUxXcKfh2oRt8oXKO3ql
xmDl+jq+5YDkzD1fMN/oGRqt2+5eLtyPE7SPa5XmTOmVlwyAYDHEgAKFEFXmN9+DNtBTs5xCjWc5
ru3e56qhpOITNvvN1qGHkaESK95r1LQTeRF5dloweN+B/zaGZkL1lAjsMfxVImH3CnBId9y9tfYN
zvomqNfGbthAYnaqk9wpK2oVfQ6R7c6xsrtKaqUlDXCvethsC5O8USrgC6xoZ4Sn4jN2QVhsEYdc
nkbghHzK9/rPthUJglWAiqpCVrLVORaVRBnGxv8AzHR6tPOh+avQkGY2FeXIFr0gsqSquZ1uWOQN
3/TlG0s5OtvGrWWgCjxuN5YaQiYM9gQ9ym9Oq43cE4Mya9tEBeh9O6lv/rx09cH/KldMBw+tA1Mx
wOu2tZUpiHbfWcizeSUAFcmLwup0WPkXicqW8rV30nQ8wYZluNwQ0Q+nEE1t+3WF2SUuybF5ytra
7KSWqb8hzrXjfCIyAoguegc9wkn8oOnJAkLRnJc5EimWFJzIB4gRKoinb7dSzwi2aiwIiLQPRXoz
3+JPrqUR0ofAyvvXeMAdvSVXanG1LESZNc4mcdCDfEW+hIbucqR22Y7byiWEiKhnJOhIWT/bJdOl
ukrmMbIxjaxGehdcYe9cvjDQbXnUj5ypOWR6QkwwAm/axTK9igpd3dPI1nb2lvvGJmwSSijzzI7b
miBlfQ2kdbkkxMQu7wpTpjhpN1Api234oC3m3SAfeZNWuWrs6cucnZ+KK/5+WRkw3gOMNnurqh05
A7NAuvM9ziNH03VePJeJx3k31qF8NIJc2RzvxV1cu5+9Sij7/2UdDLHUnASYyrrZWy6AyP8t/juN
Zd0BcQ2wZdTXBZ9eGIlE0kSkVOP/KDELWlyZi41Zg1Ia7QGBhW1yH4hcZ2edxM9Pcdo/ZYasqRWA
1d6ciIb5WE42CMcc3L36eHVuApWKUFl0IPea7ovxuxzx5hwqyKg8egF9ZMt3fBLE7vZgEzk+4CQ3
h2S32gZuhnMg2d2AKlCBcTK7AYKhYyfeKslELd/xGwrs8u/W6P47SnXbWT8ilaW5sdzs44k81QDK
PvsyCRiQXqxcP1rpgAAlVyd8xKrWZU/psePWjpFRc2rYraGSCyFLtB3Ijqf+T1gXmqFERMZPSC4D
VTIvS+M1HuZ4dgfnTETbPsuiYVBdp257s1+eaY9HkwWwkAwwHhySKSqU5lwDYjAcrJaDQbBvpL1N
eVOpTEOozqHE2KZlRpj6Zi46VEif6+g4DpL6h9mypMWzorjwDWMvNqPXsyEmQDcqCOveTVAjsNc8
gTdVU/HdWlsELAQtFOcOuMt+niT0UOXoJpfPSa90Lr8+ZzFR4Yv1IJZE0QpXEEqwaUwwol0SL8nZ
wdGdeqqN1dmzaO+fgaIMLwX06jYXw02zRmuqrCzuXDv8gkyYGTBZTGKSKla+fWQItuqOLjcyG/3r
r33+J3PLZrYBdKH+edWL06Ue1To1qaZkMzUuNS1KDe//dmX62nSwr/YxQ/UtTsKyJK+3IB12L5uX
fUN2qPotrCndNhC5x+NcvD5aE5FCEHbnzkI4OoJ2b2uUptKjIAbXJRaY0QM2WDbc9Rp4yYyox5Mo
H0sjJIuf797UogY2V6ZvdpCbswQ7nfVUh7m0q6G6P+phkytHAUSAT2GfxqypNTL+px1p8pEtT7CQ
DDhIeymavlCwUDFEGNz1PTA7BJ4OtSJSAmmuDpOvT9mDs3nlAoMU6c0xk1vcVt3RIUh2sdP5LR/l
LdzK2+/PJMbgoDwHBZbEGSv1CfVFu/9UAO1m7uNRtKVu7mP2U9nbZgbv8Rc5dx3vEOqldh4wqv0W
UVMT9AX8l77gDCmz9acVubNcp/fePmIkcTsRoccuRz0KL38c6UVwR1CdC5PjT2ip6WX0efsAuCjU
wsDOFq+6qQ37qvrE2M0IreMnu7MM9oPZKF5zrU5PFa39laf1PXVDSy1T2Cb0UU1GuDZtMJBQejW2
LC8rq+ie/PHPIpW2mO7jXWVWmtVdrQuwiP/qgQbzHdQIrnj/glOUkTpgOz4oeQmEsINCXUCP5Mg1
Vifa2oLiA9CH9ljrP3ap2Qz6QRXuiTzyO1rb0w7IwAg0OaJoRxp2ZB0lpf9fVZ106BGRttpffDXA
hYyrjaIeZsYk0uDd1LKwgn0rT4MSqSs+PK/cmtYvt6uIc78Sgs278ydwmtOiXmoU6+HOnh2fG9lt
ZHHlon75Ux4VdncC3QNzI4SHHDuOP8vS6DGyhkPAiLgKVzjsIepGsMr5LaoqgsUpJqtjjQgv6R5f
DsUM72oP21A0hNXRp6T+AqpcA65akzL328mTwNvgGRW03hN8sdEBsM1hmDpU8YzrfIGW2QHSmCfk
5d2nB9Tpn+Y/0dCuB3Pc3edPLDBKqiU77i0WjDHZp/t1B1p2KgGYAEm538Xw+D+HXaYdOXNhyy5c
lNJpaqWAXulcxYvBwx8D09yZgL9jagfVop6xER4GLyW4sE5l1UGpRm6wcsa2UMi1w5OtOgV968yi
3+87l6Nq0Hkv+7zwsATJdo/Tx4BbOfodaNoxPnWwcGylDQwBMMy10NdET+aajeP9c+cKyzj3xlQ8
5jjp/rvHbcP12aDQG9HU+o7GFjO5FQpmcqyS1oEzMB7/Hi9b1tFG6sggXIJxKydvyvVqBTpziPHA
/VUg7BptPDkxUg3u9JUZudcVVDPk6TQY3oEj6hY++S4sciHlWTDQlK+EQqkRealvAe5zEhsi8b3k
MHYm+jswuijl+5Gol1xMQ8AkBdJAdt0aNW4m7OX3qhtlMP94kpgFHCDva73Ar6V8k0YjTgZxfrNg
0kuqUgTKgd/yW0p6kdaeUhEHhgJhBqRy57HeZSJ6f7urOtqO81aHMl68yNY9JEnhmAGoPnaCdCKK
qBO+E9aubRhhdtvEOpj3waNfzYYzUYB1HwmW/Mnim+xrAeSZA3IDkMgX76fLxJjz+vfzEzDLl/vC
F4g24cNVUnMGRQ+CsIywNTpAMIGv+hg4rDw7ZvwYU3NaQOIb2Ahs1rxyr6qxldFlm52eiVuiqwj7
BNqP7Je7uKTDyMa9pf5Zsns7BFRl1T2A2Zc/G28nAf9JqLvuCJ0I12KpiTcbLo1WN0n59FMb0rwV
6rBFSWuOE0d8IaA9YSZ8uO5hH1OFRyhUZolp7wiw9qTSjXRBTcfrwKc/6VYUt1a0N/DF4bywCWSu
2NWYa+CI5kRfJBNdzTbB0dyW5ZMWqrAO5GYd4c67zsb6qJwnL7oBaSjnqPN7DUPH2m/a5u6jhi30
aGDkcntzyoz/FhkkYTu63DqZh2b9QbC1fsBMOQyvVlmL/ElEtf5yMjYHipTnULF5DscDa0mqAfbA
6XyYrMgG+ni0LzJUz/2d1ZrkT2r7Mw3ojxxR8VPkKdTwXXSi8ZRZszham6KfEGOBEHtcBK2jzwF1
tL0gNiaDH8ETA6X2LktBZAZ/Bm9Mk9J3gW5gkfsTD1CFhkDBANNf6TV5wXTUyT+IVSTOYjXg14yJ
ETGsBgh6qaXAzcq16OXrVxYykgPlU7GXYU6FoYGKRmxccUy1iozX4p1yNes5rgGNrjY+8wF3bxsH
Z8ShJ83q8XQoMxY9V7gjw+YU8PkW+Iv/CwxjR8wH8x/NUIzepRgepuLNZagxAHsvHDZuh3es/2Zc
SJ4Ob6MRqitLZXMOVVsLgd64hGZ9/ZkjuW5oGSuFGXmPRsTwAL6X69tLimEdIla8nTNsAg6OrwEi
LDwsw21I79k/UkrZs9tWyACfXyTCf6Uk0y0Q00zhcicX1BAYBrHU+CyZjmqLi0bQZMzpV7+EZJno
tHlZnVHFWXGTtU/WQ4WmrsFsqJo8hMf13JtCV2hyNxg7xIR7FtMmcaW6tki9nlXF74R8XT0lXOpu
o5eSL6sGsDq1DnCXeMYCNVVj/1Ud1VROYT+Fmym/twrg5JGjmvvjggp9sAEpTgpmhwtPMjWuKoxg
D/QueHa/qNJojn1JnlYISxwBP2iOqqBArXQdLIEPNUaNlB8s2iErbN0eFOSAYwKeplakNnn69smp
A0jRFPceH/pZiaA/Ufrv+cYrfuGRo1pH8vw4SRvRl+ur2ndqUCrhy4/nQyvvUevynXJYgb+28z9C
mnoN5JTrVi0GH06FUDBLtDFj71nXuJDHwnArPKOBYGbyGsxPPEzhJT4SQH0nyXWXfhVKf6I+ILZS
94HlPb/GTsZkvRLSaa/MqfYA/5UZZZW2brH/Q60psv4jq5K5JA3a7RE9Mhx44DhDVEuMqe99goId
6FX9MRaG7NAIgAG/KRxowJG4ma50F+s1rSgcmcJlTtTKX3LfAoQGN3hpQY+w3w+XU6SwPh4e+g9K
50B+/QmhmiCexxXI4I1yhc0VXb9t6fIMcxsldhOChG7PqlM9inBfo+i5RTj6wfbunbGTdYpTRyz1
c9z0GYpK309r8p7ovP0dGkGEDzOoaaqugLY7gpqduSeIuWoeg0zO+XEAxdA/+wSxmvILdDdA6WYW
cFfmuve1VPuJ6D94jpnxprpBVXEUa3lHvCT8tpx7m0OCvq4bycLZfUGm0y5H4DJoEXVWCYjYV18Z
U1tWJxuaXo7tsqzhvfL6ELaz8+8fE3KlBzK1/SpS/32lGPzhMK+wFUiK87CvSN9xeCfIH7gaFuEK
cUlURsMdUV7RQSyPt1TYcn/2iQA4g7M98+kQLjDX8Uh+8qHoC8xcIudMJqD0Y42eu5XvT29iQ2pD
pyEmOcNQEUzKe0n6oO3TlH76DTret6CmT3y3koEAnQUb91QYxSYCAB1y2MRpYvAzF42auYqs6C8m
7AF8oRKrFoJ7Q3+QBN9YneZCk67OI4TB7gj3IV8BGoNb4p88gOLSbTBB+EozkECwn5q+mvGtouEr
04dvpmKHCFgMmYB+nDqh4QYvPaVssXSJpCzDLj7/0RXcUAgi4s55+2mL4YZ3pMPKR6ZjeHMc6qsR
PdhLRBBH1B5YKxlfuDvOJ8CITycLo69prmjGaMyih+X40BAgQupAwm+WjsWG27jqWyDcvHhfmuyP
8EzAOz8OUlIFzb1ZMRcgobI382fguDW9u7XVBNtno9atpubmQOLyHM54FHky0a6ZcjFQ1hk58V5W
oFGsYUsk30Q9Kmt5A+U0auSuL+JafzjdoApf6Ez5qRviAHua9UW+uJSZnBrPB9DnFxzMV37by4Bl
X9TrbmEBUI9+iXeqrpHkPhxN4BM5j3+VaEaddNNhTkHnb+qBUAcFmTe3GA32/WshO9kpIl0GQ05x
sfhms1zbF9G4ZdWxG3GTadsm+PCwyVVxoFDM5vWV8BZqO+tgkKNg9/XOEM2H6VUvFm2ucG+5tMr6
LcyZv+gF2bAOgsjmhXD68q+LKQ4z3C3vWXal0AnXThRBC2r9mTk07YnERAzpOQWS8lIWyHoS5mz0
VZQQmLXLaRWYzX/wfxVQPaZiR+5l1/BNPwg3qsbRmXhvlPK1E+BpuwGgYW+zxLmFDq4qwudiPLdV
LXEbJ0loXXQT2J7woyuOo0XwPj2Ep5sPM/+mCkuYcDhUNtMhBf+vaizEUJuiDsRFQ6q6MSAyMOGX
uMNptgT99PwmTnMLGC+IfLWVgsOpM+DbkbJfjsvv2qyDxsJivpWskCq2aYWf+etd3Q+mnYTYAl0O
jlKM3bZIWFy0GjzFTsrXRqOtZ9RGZizs7OQXCD+hOpBScVAoXQ2rwxOuncdXUafJ7mt0aS7VNKQA
pUzQGWDSDdZj1taIhIwPB17tdcn8Dt/3hsLSsKY0EWLRqvxqUkreVbW51HNfLoV56CcWWwpSEQjC
HCFzvIz2QUWazbfFPUQbcB01zEWB3GxyBszzdDsrIwp4JHI9wfZRWhzBOthNMlkLounsbrJOz4+y
5i+rDulO1HCDFjtfxG2ccDgsuss+9DfB6v3iEqT6y0fp0dzVg1ctPV6uIgdEqgWfKV171ECPxcrs
jwEJu8msrRqYxcOSkNdQrnOpgR7/i9nRDu8KKAAAPencJ1H5OZdqPTyNU2E1cLhBGS2WjHYvZ7qQ
AuTMHUFqM2hqlULwtr5q8UdbMEKctIdbpoESjFh2wfdu9MZxL1KJehdQYw7pMQ1eleva1ZHq5fSn
SroaTi7nRGhQHMRlEuocURe2FaYsDr42Nc8iZDLGK6HXP44A8pzz+kUnsqVC+d+QvauhczP0EYZd
g7J0mkK/3LetAsqR/OE7U6aAWHFh4y0zmwFhHtEzvDPSyd3bXi6jdmWtbzdBLd8uxyMuvi64Bxet
kZX67Wk+tUXiQq0G14fWx10CEHsVxxeY95TZsJiKzAZET9HsazvrOeo7lHpsd3KCqZjL3UvQsuSM
4jfVO3Gj2qwfAOimWp/4vFCYHxNCPDX3H7q4IOnNkIpL+/NCODpXk6hKhv2Rr1/d7YxdPCelwYbP
huhNQmm8Gk88eVa+uh24J2F2ObCHizvnb7NRWl4hRUJgCNf3bXvtkDWijv+tfjA/rXvziFYgrCl5
/Ypm0IiPoCV2HnoX2ZRaGDIeqWuE8S4MF1GLOE6STLYb1wPJEG4Q+ePI6AnmrDV9SiwARsH9KryG
LLJq1QbVXlj95bo+2CyuDhZcDBy1hFE2/q3ethkeXjBJPPZIVY1xE3XGBsyvEZA56pShhLoADWvx
bnbj4suvUhfkBCqQKIDZ3fwg7MjBt+gy+gxw3gOWM5TuL1fGfXBYM7eJkf8VuEgxWaKU8hDoBNs8
hWs3n9CKo93X4zht81nH8VGVRJ/nUJKn6qD8wGkZuDMOLKQM1Elhcm9m653tpeVjT+IO9bCMxomO
HqZ+QqhbEB3MoooBo5NHTwfQ2fXqsUjk2JSFPMAP2oAmGN9pfT9VIG81DUh+sFog3NNbSQCiawqe
zKT/+NM7b85Tbb7kHKzuX/ZIbEfAlG64bk6CwY05xwM6vnepzbHYvyDy6eS3xpYWAfeiWooWAIhn
en1pUdUieO47mUwYMtaACmqmYrCuSisy7GUm80vlNbs4SkqxDPlvRoX9HOVUcad3ShAEVzpNNTwZ
2C/TqpBPDd23yqEJQMuF/wcgjhIbchXFNaeNTHaAawq2uWAiNTlAPP9ApgftDpYWIU/J7PhGANSJ
1mqZh5rP5CZaZePL2NfEXy1uHxAKMEwiP+GWqppRc9HILqTjnb7sQlDN96yO3QeHwe4/eWb9ROkb
3J+RKMCExzl2hmVcpifMtmvEf7UGisu5T3UCemXEtZAgVKLyE0zTIL1uZ02uEhE8YQwkQG6Ie9q4
deAMsckLDWkMlaFFXnfzMbYSlWb+/PhS79mos7byRw2O/pZLNgA0eqEb7kKHCRnSXjcZcK7pZIIH
SHZgxW7/0daSvIFDNBZq3GY9Mt+ye7kYKSieEJes1lOdg+BoA+TpkH1FsL7/m6nPjKDASN0223as
MkgexM2O4R+M6+g3mGUyng8suCxrzDE5FQ4eJ2GQDvCxZHrK6EZM1Ux7Fa/i0nC/wMcQ0zYwGfdL
YUpof4VCv/bHfxfCuUyzZbLS07OHGkDekk0A/oumqv0+lzgay9qgcx+vnEsi9hd89hI4npjUYi3P
7HkRfxPxPJK4el8Fp3ooMSMhJ7mYx9jvlnmorFXqfHRMpi8uN9VbXzXWnM7os43MFKmQezXU+LS3
fYrNpMBJNe6JFifAIYNiP7R3mTUhc49CY4ZCz3PrtSc7WfLtESsXFgyP6ltaP4axuqfXDZoy9ITs
NHSQpHB7Fba8toC/u63jT54pt3l7cv8lV2ZWcCXLQ7qwo4dSiJ043dYc89Ohzry93m1ihNOB6m0c
X1wJMXvyO0ZmiMStKZpInYZx9H4tH/S25+YNWUmey+6aOf7rOXVtj6o6FHED14Im6n7BodZhkSh5
+07gaLB4yBWvAIci+6lT0HX0DW54tpfYlx06FjtKZ+0zmjz8nbZ5Fs52L743L8fsjkH1U7Z1DX0c
ahUMUAgkG41ITKEXKOeQP5SYCv4QcqeroNJN84q6QlES8pxFWj7px2Is0FTt4TnsGTA0KGTWfgQm
z+XwpDrohBvnPHw/xWrUErIbtclqSOiB9xg/p1CYBB4lh3AfpyQ15DScCngTqattbMK2rNvYdx6z
CMR6HlGh/nl6RrA5/f3cDctzhfGJ1IUpGnBwN/285q97xsZH80EEdqLWRMwWehkrb3nKLR9S4TXy
EYo6p6B9mDczfy6DQeQPA1y2ElcDILeG7VgGsgz+uxWKfOnHWfs0Czr2B4wkLYDw7Om7DmQs3VYj
tlY4DflUbqK6UliJ3mPTPPIgbyJJcJe9U8LGVQnh7V5rPYbCaj8X11W7e2p+QBtcSHJrfrSPmBGw
rQAW3NcSp7RunteY94TAA8RFlz7TfUWfnGtPjiSAFALtgcB0kkHN50crnFwhK79CAnsyLb8io+Ft
IMlJ7YpWzgG+/5fTG7/Ggum4MLNlW6ndRsHqxLSfAuAF84EQAAgwoAvSgxn5hiYNA3vHAT3JGW+i
fXY9hXnR35xiji2rave8/tfsdpNjO3qCtJhNv3DkFHxHxNgwjzUEj2fenW8dtZVTVKl+gKyd5oQq
OhJ0N+APXQM0ZBO107IXCHXcweWhBl1dhxFj/ZLKhC8jwjCjiq0+j68M5p+W7HtVYbf2tyu0uytq
Gt2t91NWXLuI3rrceY6A5Bpx+MDPN9UWzaOs9tacOletYOYwWZ+N6US253/0aC4oEUgYutDQPS4V
k4xL9cQDmqEY82vftfaD7Kftv0h9RJ5WMedFTkS9sUMeLJSeokp5K8ouIIiobZHIouWjHEB6PiD4
hk8azYAPXBhn2/UQE4UFbrvlaENBXXXjYciiyd5U9CzxmPPe51qgiezjE/dW/aVN2jUq88DKtxFY
WdETLu5AibcKpNi6ns3i6MhB9TEkNMe3b2mT41tPdDHcS9BXK7edvdIp1MKdyNdnMemIlNgDDJXG
fQmvxd7arXrzjA4vznOXgMRpupf6IW0nXg8UfPj09krH0Jb9ryqvNpRo6mUGBkCfM4odAWRQ8TMQ
pSSqoTP5zYfeYbBqVTLamhs9J2vYJv1Vh/WS01CkrXF9wPgy/fGAGIuqteu1pLpk4e+FZztGxrh2
Asl1Iom3IVAOhpBwSEHsV18U+FeeoE+DVZi9yHZ4iFOI94Gr5gZkrs8xATKqSlbnnwL8VedfkDU/
E5xndvsdZjE9rXCjs0guLCFqwRgMKlY8gXaVP5AVxLZQgzJ9rRDyHu/i+8qCqgAeX52SDrUdBWd7
6OEnFQcB/aqpkwKVjUQn3Xu8amDknqgEffTYn4Wz0NoX9JO12rxacQrMw6aTOK+N1/AhHJmBOS0c
ONBspZ/wWxiyJfyeDbCe0NYhhDyiiP9JY44TuqshZ5qNFTRafWjbs6LXjbwwjZUe5EzVqtuFa/u+
y1gtQ4XF34uthSfBR2RWhtW4/UHpvjmrtudsRZ/YkTcHFjfWTqToekEiQiJOxB6vCH44gtkDjMGU
3GRTOBj4LWCLE8qjMWArw2+yGFRsK6HF+j7JJC9AQygV7zSonuKcWcOcwCgcUhi2RDeu2gREOCJ6
tDV7rBRE5dNmqwn0eB8Fa84I6crXIOToJGNVtNxKeHaNyfri4YkbDdnb+Roqqp1dzd3l8FRmYenr
IqPnuzhFrbvQ1So3MEU1Js9IJTVoK+h0QXcRXPHAh/b3eH+Sr8SMfRsDKABgAztoqZZvNuwKQH4o
GmRzMlrILO2/1lMqKfWMl7UybstaEXzn9+kWV7Mx8GJKne5RM7z5sQCGXZ1IBuZOgLcayTR3Luu2
VSwZALCL3PbDdT4iiBhm5g6UOfB5pDWr3CPqWP0FY2uxFvY9LMlKgVQbFABt/oknoL1dmRE3ioRk
sFil94RS46awf2qnTR/yYkIjeEYl4l/+/U4vCzp9q5l7KtafylXP+S/C+a5qU2eIcza7LnjJ0nh2
dJTrUykPmATw1Nqd7YRBRpvyAy97080ZqSlC6eTuLVKFvHurizwcPZTgQKBWQL5bEt0APXjxceBU
DODP/9NRsBPbAqonDQAV3SXOEudR6bWowO8ZVmNNtlgzJqU+TfT9LpGElwvcc75NU26gL/dWVZOH
WdVnQIl2Nsfm9jl91HuxOaD5efe3b70s2EIlrTU32VevAZJe21UxRvcb4svo+5RGilukde4GFFuk
myc8yojqGXrCubw9vuG15KXIfaKQpxxkVBKLZvX1IPaRj3tjZq0ezTrIZCnmewi+VkR80kklL5ln
NHy49kGsNnEc1GEGn9fY4XnQTbuNVsauwXIm3zYIQs6igQCyq/N4SjBm8ngVX0uhBttgX5R3DL7P
X67uIVyoamT4DVB+L5WbPff5wIklq28DHj7XQe+/3twIccprEQdgljuD47ytOnQkCNJ9wWsIdIKV
gItbVlNRoiImVeLfzxw/6QOGBoVTeIi3/ibXOmjQ/8AWTdlZTmrk0efGeSJx897Fyybr2ct+dhjw
is1RjJmqVjll7VY7o4SyEB0ZgjkthYPTMnD5PKp0jDhUKrqiaWi9UMX1F7oJ785M5Xi6gKIa9nx0
YZ0SMN1DJsbtTedDuUCIriEw2eP2qr/EnKMolToAkoZWS1XoJA3gwAb5sCLwclwMocok8nxarMXw
cUTwqgkdqBQdV73Mi8lR8ZBbb4Q9u+JiWtvWwF35Y/wTo/3isfAMP54yWC1iav37iEW26l8HOMem
Lc3cj3PRFtq1XG+QZnVUOJ12xilGIBnRSpX/hWsp4dum5YT3p0yiccOR8ZGdXvppnJszYYp3J8Pa
fX0IMM6dzPcorfsdEx3BlfzTGFp3iBaFvpxMDDs/LStCmeG9sAsL+Mf7FZEY0HK3+pYQ7vEnDq0l
YRLL3WYo2B0mgY0FDIabJTsBYh1K1YIfsEQC1DeH2/LOOPo5sPzROdS1qKYMwOPOL6os9c7p9Asx
WR7OiO2N634u48gogLvRkCPua1zNbNMeeyy/BAG7I1vuOBz5YH/PcebQZWZmeNOPuvx0G3piyD27
iAgoCQZK0guXYP/VIabmNdbHhW7piEqk1y68TcdggpRHO3JlVbiTKD+fGFFR5bH7vJZUFl0uKYm7
WVzcVhsCUUISUvnw4LL4w9QIDYUvjK4NxxT5YuEDiNgvdeCB4mAIwTN0sAVkeguz1S/5Ive9m2Lp
W/6+hGP3X127dU8reLm4Cw4lox/TcYOlHxcprYj/ZyYMvxaYRfoFm1QNNPUopSwgPh8O2PM9xrps
5jiVWxpkBNHkB3QFOiZchq3WmTCmPxVaC8Q9WeQGX2jA4mfd8PFlZCqRYwYpDiFjEiblw4Wg9g/P
C1aTnBINs4UEVm39N2130tm8l0ehKBTRWEYPTFjAcfHX/uFjg0lv7a/JLyOXC2MJ08Fc3sIbl0fL
6eOkSGnxmEEQTcGHbZUIX1JVh7uGFxH/MVpHATtiRlTkpw7+368bFtxl7aVsn4R6SPDFwEgBnw+a
PyBpGC/uETbWIfwZDpqj49OwPEdqBeitMcoXzZ1/kZa7JT9+F+GIzF5XbRx1luzteuUdAZ47DXpH
FhI7rRESkwzVDWikqQ6c0AEgL+rQpCvzk5gHoLflTnrX4RuaC6NGlcjVEG/852aYItLoiLoYmGmV
L3zMNXIwzWQYJpAXsOixkHa3qqpuL14jM0Jk32D/oQ2dCfraASbWzquuZFqt7smdfeXEqktAhdZX
k8KiBilHWRdLc/Pd3xYpqXpWOKdTKu3SVWYxw47ulQTF2eMECG3nuSklxSa/FtEOmxxEdCMofHEK
b39LrOjZbr+AGo2g9WkDdW89eyQLiybH1KVNi3+aRFxybhzKb7i+0+dbGLeSMVzr2mtIaO3hD9Qp
idj/bRO6m+KkXg0gWxszhYFSywbwgr5kFZ8tblM26l/DfOtc0/bmGjIWBFaQ6JuQuFgshnw9agUQ
YCwJIUecnEqgQBo8tjhrBDHMjY7finhws9rkezaKTFBopY3CeQW5ZS60oUHK3KBl80xkZZ1enErH
z4gjJxCgFkaoaAoM1recBAGERboCWQvobLZofbbsHe46ACOH3rj8//Rhe7+u9nCiSUUErZ0Vklvg
KfUlAybY7hTQdASnIw505fu0e+BrcMgGNDCZtSDfDLs4aULReinlP1uU+/JIOsymEz3xdVAstnro
MWYmG3xDkybYVPnd8p/zyrUJnBCiGTjNsuu8bcMJCvUDN+/JNwgtJ9TxVHvigYDLBLuqGCFyo7ck
tbBRStCNkPethgLqr5sDQwDUsFCYr6zpF+mS08RBjPwfdH+PdbgkmRlwdzWxA6tI4yEngzL6lrPK
lDIbl/8nrjVjhq1y50q1EyUHgXfYW4k0ffMfwMGRlnnP6eVHuqrs1+0Ge9eoCKWjGN7QLPHZrZAI
GrHK9Enj8KmOgez/ei0vVn1SuypLBPxWxdAKFzlTnKc0nEldDbUZ38qn8Y9r0yGyXyZOqs24OO9f
g86KiWWH+5fkXL9WqdHso++PwgApRTiuV0C4alKSfcyA7VE3wpBqyQFZbBFsv+cwBijXuii14ZFg
KlFcE96Z7f2/vflYJZ3phOus7ANuaTKIT1LVvVOSXyEnKd8q1aWOTGXbO+pZjsue6M2GrqEQAkiu
QeZ0pfDQc7E429b15xi+gbYx8nrHgzGBKtI31kS5LGzSjQ83UDTuQwuHquCsJ6pQlw7Ir3BWYzx3
/ugsZ45vmlu/sCMqRk+TZrZMLXChEewDLLakBX++7FP5KLad8L5SumPTOxsY6nhE/HIAFDJqJQ1u
limT+dIfVXwH9i+OS2+0plq2ovXLEfSSAnE3vC8kSQB22GQh1HLIoQD3J1xP4F2n335W8biHopw1
MhCkRRJASaxFn7ODkLCtgbS3JycSO+j1+XN246xTVSGgc+0eCSA9jKIjb4OcAHXZ7QWFeBFOfhFL
0T+bgUBAn1nNyPJIba5Dmr9eeOlFnTTfLB7K4HwNwoE0gAJQ4qLRszzgigt4N6YDWAZjxuVwVmm0
FrGC2jkUcJE11Twx31PmQ1FLlL5/TRJphY4YmrIZ/2OW+sBwEqm+70QXOazTOsmW8hNoGVx4WRwK
1lJgxkMGaQGc4kKDx5s/DzXDPB637tbws3tptXTqw7Qczug/S+aZmLDrId4joFVieDj/XGy3z98/
/FIe2xTYVRnJtb5HhRxWYzZgCaYTiXb2fQAJZz+s8nHTBQvVohD4tVg5EdTeeVC8pI9VzjyHur7b
Bar3aXkSqYCdqLW2hoCBQ40UpJpI1MkYBvlfExOmxxN9RF+n3JlmxKzpkUmfMEQikTWyJ8PFZGA0
rStkVM9ESH2Dj9LeOBTOkSnWlY6bCTxkBnPX5owYNBq9ixJNGX22Gbm3Dl0LmBVO0as4WEJANnE3
lFesdy0zNk1r2rBgiOn8qxV9jmNN8jmY2u4ywniMaAFcebOe1+w0sZrEaZLeCBK4/cHUFKxqGvTJ
lULGSL9a56rssRB6Qx32KBKD8OxPTVbB6+wRsrIst1CfBBSVqDa9PAnliHAJWYdIbHgmLKdqEXUK
gIuU+7D1OdUG5qouum636PGDVRt0RIp4LjJwr0FUCymZywOed6I5YDPkKM6yvtmW2lPty1Lu/6GN
ieKT9/GoxzNZxdmJ2VsNJvLStOQx8k5kDN4OjG5njHB2b0/9lmpTOuABw7K2iDrXkXgc50iyhlNI
2o3xmbUp5qSJsTDzrQqH07rfPHwa5ZPXFofNLFbss2SX2V6FQg5qIxTZ0WWMBPcnIG2mXyuCCo6w
42ta5bCPr1G5VYyF+VQJ9aUptOr1jnzm4EVH1/47FCu5rLy+GogpOG4OZFkJI7uPyU1qESIn/skU
GhHyS4JEm82awaMshZ1tiv72Ww+G1/8lky1Uex/OwMRJit5cgR60KLxBL9sSuGyjC3M/Bop/ijIj
Dpc2v2Vx/JRvDQv3NfRxt6cm6t+eQ63X5jXRNU1vvUiZdHquhQXkvzfqw9XDMPJ+NHj2VMUgn7Gg
7Cjj5As6xkzSFGTymRPNbl0HXeg1GdkRlGqKfB3jE2imIhXrjM6SHC+Q4QBMtt98rXjrNwrDy4mx
XA9c2jRN9AZpVcL5k0khPfhRvI7fgxv/cK0N0aKQx9AouVFAqxvopc6JGXuHy8jd7+FX0OD96kp6
PsVXb/vP7qa6Xa6JtuWoUTsauye8BRsyOnlfX9QqhycAEB3aTgIMwlwxjWX+RXeiKKVUPsK+J0eQ
TS1bDq+eKZLzmtI7UuKSnCWOEslTwdTL2e1Psu3abcqc7IfO+t8VUUIHU1AfxFeuMkdj2Ggs6J6k
llJmoYvkNJqlsW+SjivX98P8saAaSDs0C5+P04uUQFwLhp6bbOMMQnZLAlfrKXQqzSK1T+lJciqE
S0Lxbu7cU5la1jxQuodzIn1NHx3DrsttJ7bpmbIYe48xkj22v2c3ZUGU/8bfs5T2uPu0eauG7yxi
upXd0YJmj1EdkDWhhSOT+8c/iAGk8a3bC5p6WcvVLLm//OMp/y3T6Plj+wy8h+ZYvLIGqKAiUmUC
RZTvxjXyDuA4tETjAnzL/FgkSLMQQag3gYVOk/eAZcYA+4ygv4p8irJy+9/E2UNkmwKDkgjuuflR
pPusm1YVjBHzSCzUCtEgD3zVL0oi1+ZFdNicOqF1DxSX1DU42SbBap1G6Vw+2s1RdptcOui44jML
Ihf5x1jPDJuE+9Bhtvcp3R/hEDgxYIM8APDFWOon8FLvlGoeDAEv0H/qah62fdnlf4Q58g03puo0
b5WI38f/Hhc9ly1jYn+YdNQ8rKVi2RjnfgNmVNKIotnr7brN83rID98YmacaKChl93QN3aNG3mFx
CIoZQJk5H1V3QQvHqr+2Bn9jb0kRjJc5RpXeZk+jlNUT7xMdqw+vSBKD4r6uysgl7qBSHdFtCG94
iQoJD61pw6yfjjJtLkEA3tkR95NLfBSlA3vo0UdErnJPuctfJSr+rUlvg5/AbtlBck4h5vwEeVw4
rceayhLuaj0JeF0vVfd95/7VhB+9Z8xNOWCxswQAyy8ZgOYPNoiCsdO3IdzQwCakSrdV9rdipbQW
WWB2XUOcq/ukZhGhCZM1gCu73/zKF0C4KfF0lJVpU+RVN380VR+eaLvfnyuKmy4z37NcpurqITuL
ib7RM6AbhMyLlYp/nMisOEHN6eUSjuZfeif3fICgRH6g0Izhzyc4qEKNRKW8JwYm3dV0VTBRXtr2
H8M77K8bxAVHOxx3R09AdWYOidu3ounR50SC0wmDsJtI9/ZEaBt/foBZi1FeUK4Hgy5Cw502uQ4d
dzFzLzSWHv/JEieea1O67V7bOwnB54GGdG3jHhGG67AFsQtFthvOUv/2FXevyOgW4X7gQCffbKZj
B6rt0cVVccApFkcH35YPK3zkUI4Fz+LSR3h7OWFLbTquHc28O7aOoOeCjNBfckq8PuzHV80LSNzL
DdwURFa6hyOqkIVhxhQCvqVWWRAJ9gJp5aBZb+7Y5CFytC93Zh8vvlVqwBSDLQ3tP7E8vhRjB2cr
intX0GiKpArIRj5Sh56YjflxpKQ/w5/5l2gfITSCoshZD7nelpMHELo5GlFQYrNFq4kW9JVo/gZT
IlOc9useAGMFJQkpl0Rv4sw0+yf+O8IIK8WmBDkiU3oEhWX6eoVzFWknGcpasU4HMEI46W69NvTn
IfiQEfb7fM3+IeU/1HQum0hqzXFthUCwcPQGol1viZGrxTwLQNkYi1CB6xc8qX2Q+r67wO9jFGA7
uh8F51fC445X1iCBAEuyGLLGWPnmmqSIsbcYaSoeSosfV/QEblputDWQbGjGWYYSJ34Z8PrFaGYk
KN9Z3Abxp9E0+pL6Ywuk+JibEVHrcuSTA7rE5q80KDyaYCJOhZZbW2FkhIVM5+iBE1fT3An0rvZ+
NEFJaXJ/7rpUJmcuGxtx3RFbcT0YFn0j43IWmMkb9AOSFIzZrDd+httC0POMhRS/jQGPEveFXMIP
XiCIxWPehTNqIz3T2Kre1WUxyLxsuF1Y6SVT8yD5AzEFHq+uue8bp4zpbifVt3xuhnEwvHQqxgPk
dAlQP17An+DKxc+SCCTmLWc62o0MkWSm4ay4WcvLHf4VtAF/z++KuDCvjSKBUBvzQWoXmcrlvfb1
076uoOHDmu6m1/HXeVGykCgWR2PH/tGTHM14JLXF9v3jSyilzgsJ8PfPYBtdGtnNgBCEWdIb1w5P
uGsvMpMynKfFAVe0/6w/oUO867ZT8OHk9916tE6AX7+T97m6/ELU2lnGhQ3KkJgG6lND1/WZWh0O
Ps9iZe61cbFFCDLq8Y72wo0ZEd6YMvkVoiwRXzL79mKvknQ4b1vPgsyVfbS1TOFC0gXxR9mcPHXG
VEtaeyMLDFetvdIaY0XOlJtWzCsAo3hSp78zHixztkD/iuTg4cUkWQJpTzwgonX+B6143912Vn2c
1h3I67L21DYUNbtKYnSq+V1A0UyoZG0ThmFpMgIHBgttAtZfff1S0DyM5bJx6Nv0ySnGf49UJcNN
pj8OHjadnd6mlimvGrORuqeyQDTP1dclC0FxhUCQijK9gfHZbFdzQGxxdqR5b2aj1cjdnEO0ObvR
EYZxvhUM0Xyab/7f6cUu9O0btF8BUAQ6idRHzXaVp9BGVSxNNNAsF+kyXAJxVnK5ucZ572bHNqfY
h4ZILjH9SDPTIYD5PzIJj146MXEHMU/WhFXXnCBTFAZTEJzrxmc8cscveH4eBCufdimTyNoqSAYb
rqhGmT8fWVzFixe7+wmAkUtgPBd9H8Yieb1j05W40BGgRsedhVSicaGgIR6Xjlsg7WeJ4u2kVlxH
62knrm9p/+AHrfKvttu6EFoDabFJ92HFOvPhu/kc3dNVecGH4g3gaKUmaAu++uzJMl+qC1bzWJrj
jxjWdprS6h9AiRsnjRnMOqpU3kJd8sjia7Ba3VMnqw4tk7yCMSRusCrG3csTCcH4nTAqIl2AsgFp
QnaXTPHRBnX2XaL09j8okQEuiAbH3Ty+WkXh9sf7pbikP9J0VK0IyQx770Oc3UtDqVmNRTY3Ul2F
LiScpL1yjGfU7cNy8EUSZ3VQ410SEhpo/iaKoOrDTIRlQI05Tk+fiE/UbpGV0WcoXj2J/I9PUQyt
lgRdXX/UuY0c535XIqOmQ6SBfgXYxcsM3KQYRlpXpm+Z6vW8XTWSvvNY6eeJC/hCPKrbO90TzsnH
zXzkAHCy1BVjpqb37UihD7ipTTAkzakCpU+6dL/sNO/Qmj+Z6LcZ3FUFrjV7zP8BFSXPWCbjOtMi
lB/U8fx1iVZqngjhWkDTXlLqYg0mumohfF+y6IGPBGbGHc/VAHpwOsCNFgQQS88us8wsLfHgxgdY
/vd9Drbt49bHdv38S+9VaS0u0y8pwkz5ra6zV/sPqhHZ4Vid8lapnWd6w2hefJ+qPqAWknsiVf6s
iqixm9EpGVIz4PvXi/MkijVtVlFVDLSyG+Wu9n3ZnV34W/JH9J5ke8SS1OKma1j4p0/b9seBtbaQ
t7/aEPlZ8oi3AVU8x7f51TKMrEdrhuUoC68V4Aw2ex6c4HwOIbCQzUceuKSqq7EXVpAi2GuONeBt
/JM+szKoWYxr3/kWGJZJ4W5WK/fTJxzR3uRCm8i62+rHcSk8gN6mFdIYUjYHcNz7gC51BAIOEu4o
izi4RYekbGkQ2hp02o7wSiJdu35wMAsO7k4BSAvTxsQ4he2k9X2DyBns1ZadHQ0uDhf30+krLgYF
kT7qGhNRQh2/s4RrSLyRj90sTE4mRIqBM5SDMzYXJkYHQ8TBkYASQ5R4ffks+4dSj9V27qmb8xG+
ZtCK7XPhG9og0h5zWri80PRDn6H1kkWBrhX75MGwxdnNWqorU6RejWeBrjVAzQtYzLtR/tdfvh5C
7XjSu3oiohYLOT5nRiURb0SjsvR4JXIgrrYNwN8xBrC7bP4YKUYoF8vRDQsuT48KYWo+MkTba6Sl
iPxSWSryZO+HRq30tB/isXrxgh45N15o3IGGeOqbqzxfsKoVC5no7iw0ZTCXps5RTBcvl5J5LUDS
5rKKQz2N+oNrh94q7/tj9G1j2BqZpqS7EsVI6BzDNgA6RdYhNdjvz2qQi1NhMbuG+LKath09Z2jI
koo85YsDJrT00FIi+qfg5YlFA0oQaz56/mGrF3DAs+2dAy43xS4sYTAL4/ZxVanZRsSV42no3XL5
8SZvEoiH3zn4o8FzkHrYq6Un6ZxToxo8Lwryj9m2TXHC1NnpTp/I33rJHIH3FW3MyROtgtXae08W
9k+9onfNlTl/Pn9ZG7pC/ZFH/EExf5Lb+gm+/RVYDkjbiX967qj/hp/lF4UOWzP+2wNxQx9Q3cSH
3T0ykosckjN9l/2ElpCUmGTbuJIz+fFDNJsSJkvGgDPyq+ldppztyqBDlRKdhozQkutKmoYZ/zug
YaYbyjErdBVrANXtGZ+AgvSkNuBG8I/eQRY77LqsPPHHp9QSw8g8HuJH4PbS5rXc9DJme60S50OP
MKmTCU8Lf5JzCOa3fT02UGcKrsa+GxWapi3JxIJsmKpC8oWRgymUdoEzyRoGYGA0O6oErb3+VOhu
V4rceBH7PbxgllTyKf8ilYhid9fBIFTU6WL2h5b4ds7XzqxOci1KxWgpx3N1eieY9/hHONooZsb0
+atgwxdG+F43HDH6DfkfdldQkIAW8Y80/ls8GDdFuls5klBWS6beVtR80T/RxufwH3C13Q/1xIvR
3KyNN/7L0IDpO79WXRtdHo17IBiMvSE2Jc4qDyCH7rwvIjz/5/MqtYiLJ7dWEDOW74+txqfBPBxS
m/aUoo4QBAhXkMqM0E8EwSbGO3HgabyYb99IKtnKlaHMYfrnClSPlzCTlHH2f8fb8nkfKNTGlyVN
Iq17WfNFXna3QfYyE8DvoacxzvC42IraxUfozdKg8I4wGXt5AScv0m9jI0WWjFPSnO6P54loJeil
FbBAK/vm6CKlo4OV5m7HqVcYeijYrMtwv/v4ZtRrnj5e6SWl3RShmsW6q6Lzh4UvPckDqewSXjmm
afZt1PHxk4pGVOlUdI4D62bypAP28guvddMtb09oWcuth4pJ1OkEdEnep4LWmmIRUgngGLuEYeJB
hxW1oNJgAQI9brPgHp5WoV6vUWt0rImXukU3KVKlEtRdbidsTbdqn6uFkxwS4evkmVMWugiOhc2Q
ZtFNboaP7EfXIyznl4WSSqTChi/REh7dFTuwEl5GUwGJSpBppdkKf2tksDgy9M2X7zJrOJfAugeh
HL1hTiKw5ZAB9y0DRI0DfGWcjmaKSHUIDlcioiSlPADepNLGltPw1PrEx0rX+gyj4SddrOhe5K37
rb3cgYdJuQAoWJs2ZO7xgYlKLPChPMomRR0e1OX5xJit7gaxwjaxEf7DRNtQFLcO+3g1rz+2kIlb
NWLEtjucO9oIsPaVAoaeltA+H/RzyMPTXJ3FrjZU430TlnuN/TnFEIaPbxo+i43odDZDFG7WJNoP
EUaJrFe/PkY9n5s7o3Nd+b1s4NepN2Ow6lcjE9lEzSLV7fCtzdAPT6uud+YCYzX44LmUO3uITnX5
1bM3KqpfoUUDNWj5IPU1FJfBVch3ipI7KCc7+jIw8ceXlcunmrythnGiEp2j5OWMtAHa3D9nthF9
89OY2CiRDpuJEZVnPHhLbDgouyjecZ78dAxzq5sawS5zUILTigTvKWjyqkD8IXO0GqMviR4APERl
UeGtajkVk3hjMQcf3q/ch8ejvoxs7CAc2HlMsiyoKOZje7jPR9vPDjIiL4H0zjHFT3wt73ULZre2
buia6LdYhxVaAI/CdogYYXmR//1Vpg6QYSF9qA16acehzLSyr4ylb9JkAlPKKEdciLkQMqQ5Pb++
4xttgGjDE/vfOr4lO5o8ILbA+nU2FB6DEr/PE2t5RLGJQT3asukTVfydKldj/tuw+GqaDccLtaT1
CEXj2YEiwQfvwKlm9tjvn5hF5gr1fzEED8B3rqJyMJ5NEoLIRPbBZiY6TawcvnrqVGw6iPUCaoqe
tH5g8g8gIe9+L3n34WNYPMA5YLjxpCmeA8a16Pm4JGHTbv/mxWiDg04yFny/lJaM5oFRQlXCufxN
hpA9w7Gaf6//0Mniwu1do2VmbNa6SenBErgfUVz/itvhCPf/HqCDY83E1xRWVwIgGpLtKLgy3JCp
x2TjV3n1ZtlW6K1ZFttNNgDRW6M7lvLB440qOoTlMUNcfb6cK3pknyGC0+ob1wqbr/NFMt65Yd/U
PgUGHc6cd4IfMgqwTYKIcf1/OB5F/ZuaamDrv7y5p3uFUvchd4JjUFleDVwoqPbPgB1zCst1QKzT
mojTDY+teWSgrdqeAWIoVzjhgbVxmbHrmLk3mUrqQ/R98qi3iHQ2LCJvk4CgiAKu2SND1QIyL1at
KFGnPI8IPYDQq0nlMcJqfYf2K9VWLIm0QnkkrwJKvPF8EENDdYN+op76I1+opIe9USNdQ5WonumS
g0LVV8Y4jMbzIw46OMAsBPajzVrnTSEIQLXl/KygBY2Gn+SnmOLqAuMWmSQW0Re4r9LAizlVmzse
HWHJzfo2UVd9YzqkH8AFEBX7HRF5oIBlNXDKlw+W6UFt4KM84ligmHY+uDttnXOVR3sOf5G+5naF
0IX4qPCF9auH6PxUUioLZhQY5aW8cChEUyvcEOS6fl7kW4pjuktRgX8bBuisdVvpjcV3cg+jgILC
RHX1Okid8tD+B7yRPNsJe9LoywvdmXwchI5F53g2eLwQ8BexM+1ulgb86YqjXL1BVBPIPLfxZvL/
JEJgqSTaoGsc5hw2i0ZTaJ3FC4z10uwuC9te8FcVi72aE8MTyy2Vi/BexMGHqGTnKUtV+KSrB/f5
ODutbWjoVPA3QbkMslL8dGFfjnc43hMM2ETEYFAJTeL4d7lKGi8v9wk5Xa412c56g5WR9aaoS+Wb
ZtIJsnZwZQxmA0q2Tsdd+dO0GsBJM4OkFFtc0/daweP0ViwpAfftXrdyQYTAkLQ5KwvpYRQb8/sP
HZSlgYd4Px/A8PEfNXQ+q03DOAiHEEX8PBBIV8nSa98zrzsuA0ivbQi0aCDP+BoSWgMPsWjedkAB
LKuYJ2kBxlZ7ymlPC72kIDa7SnPn392VBXNCSKp7X8i8LhPHjABP0/AyVn5NJxFyXlIdnU1dwkfR
kWt2AFUeNOzBIYdYV/+/kB9bra9zbZnYC2G8n15U3oYV74G55Atbq8+nxqwxVmO2QjUnb1TrWsXi
uFAx4fvZxgTzZn+MxrKWw+Wc4BlFCn/F1qzKi67nxGDIidwKWtjpR1dVa/Gs7FLps2HrqCr77r8r
kAK6vnkgghb8YKZQ19jT6yKWQHk2us3DxYBqR+SbIeKG3JK0wkntcq+MRsX/4+Jt+w4zcy+V/1o0
AzX+qpHyHzpSvqWWoXzsrhtnrmGL3q6aG81s8GBnOVRKRt+OzKJY77DCrK9LYl1ylTtgldvk+XdZ
Lzu4AszICe0Vm3ZrKbmhtMLWj+23EI/DXkuZYG7oya65KhBpZD26teHWeJfE9a+Sw4Fw7L4U3MQy
PGafqAj193/OMcJz+s3tZl04nGbhO8Ln6Iilqi2iwqAaxa7vKPGf02Bkf3uytPZXXgghrhrc6i8Y
tyGEnzzs1y2eosYzT5wnOCahFPuTU96YpM+G4c9wxv9rSm77WrR5fn6kcGaHyZXWRdh0pPnGIJef
xWO9ZwKXfEgOioEjp8fCsmiCBWW7gWu/kTuGw9xDjXKY+oUiqajeTZGB140jx6x/pOG6bQFF2tJl
dbzk/4JAFQGQ/lhgu7zhnANxddNIA19zA4t4k9nvvjb7CmoKoyQ5yWTvKKQQ2Nrof28DpShc8bDS
9IDARH0AQUrOd5YWShs68zza1repg6+Y124dv0OmQ7in9fKBZW0YPSl9tyaysVw4HMrz4mx3cqrd
NCzVVIV2SSVOSyUshtxxKQ2XtTP13+2sb3FA247iguJ3Kp89Hlal4/U2oBWB2cplW7hHJtqi3W8T
ss52GI5e/gt4ZBNP6B2qha0CBixdlJ7+r2uKAAmEWk9OdFTB+5ZdZhrKC9u8H9zngQX+7rsuPlfl
RXZ05PxI0qZr6LHpwLripzG4dAogXZDPuf75vjDN/sCeUNt4V5uIykTtiEdZiLmLqgyDrm4eOdN7
DCXzkz0TNwsLNwFxxI5gfslxaRV08cXu2b9MX1q93bhrEyQK9QYt91g4/3zNJbvLMxzI1v7C8Wu5
I9jg3W5gJbzEhNJYebcvZbkMYEeWsyBz6CKbbm+Aw9U9dCcnqH+IKb8LNcZ9zsiswC7KTvDT44um
RUuqNbPRPPBaxXdQ/83PIQb8uR0mnXuYNICRM2VJqtaqknJpL8TmBH0ANVCodsIEHultfJfdnxSh
Lg0RYuN6+wqc0BkqCpZkvqGwWyrX35q31G0sa13cN4x767VFzMEHBrboICfNhFnqaxNhvI+VVT2A
Homy3nkhtyif1NAPiKFvmMtfKTLWwOzRY3h1RvrI5gEWw6MK96X4IPYApvgYD1WIkfbDjQs7Fb2P
ZvcRHjQRIrV+F3o+t6TsRWxkjS/jZsFvziSn2MQ9Gmq3DyhG1fjzAT5yI/pPyd3cEDwFIdyVbkPV
s78TbLTZ+wTqK6PxKmyGlpuo7jGX3WyxSEQ5yDUDKzTy+gu7TQ3LOwHkZGPpiF49P6u2zE0pyVy2
T3/QiL+4kwtpuc3aCh9oCBuE3nTs9UNmoafhnZwjpTnwZEH273Uzw2ADNk86C16it7AKXg9GSUtj
BSo4//DzxrnE+57GYM9oRI4KR+plk4ipKmpKAmJ8nGsk7fMVTk2XzoDCxvVycXA4UIAwtLXGgkqX
S5iXUUkU4lsj78beKkJOrAm/wIPYFw+WdiwZv/glwyGsB4mJfXcQp7RllabYaRKlHNQsplRys4Ky
Jtp87v/sEP4CB/+FpBM18A5XQUNip4OTu6TANftgVdNrioSzmjtxOeGtdiYFNfspHke+bQzKXRPs
Cr47i3AupXbiI6oA83DG0qEBkD8fqgHfnTL4ghDdrAxLAzOivqe+CGBAlDkT/+1RAcOOExpScPGa
FYhcyxZ7VUC/gr2l9cNo63p/rKxwPobwPoREfe+TJeMq98XhOeCu7lLcsh69sILAX7xyfCfbTJsn
QmW7mHfXnHQB9ln98scA+Tv2LsTdux5tJmDy4iJf86kNhXl8aBt9B7RdfY7GMmQpDT4iKkyqk01N
Qq1nr3+tPOhB5qZlO1Zsnz4VD80zTTOK4yzBXdFlaEtQ1Ol1ma26w4Li+fYmyDXU37F6v5bgzhsB
Avv2Ecb0+y/SpFDB7q7HjG9LVNvrnu8FMxQcrMiVVy242uOl5Fh1UPEFRShO4CghPaLhMt8DC74K
TNt9e7d48PPXgXve6S5rP06GNNAZQyoy9uhh1pSVAHGT0IVwrmcVBp42NkN20elBLxBc+L5HWItR
6pFsbOztPOeS6xpWLlrunxBAJKFWZhTrXenNIY58glMGnzpN+hMb/pp2fkq/5Iz+Ad+uEdx6rMGI
WrtTTTSnBVT2xZn/oPYAyq0l1dXmuJIof2MwlTh4DF00y1CqI3zRHszSURAzlOD0h09q0wAUgElc
jWYS+j2Cgsuf4HrkmKpaGj7Hoc9WtmlI0oVFPrVuwPB4eHFZZS9gd8pf6Svv+yyDeUk9gEuZX0g+
bLGxGEjbKBWp4zYKRydZvBegm5CwHkTUkRruR2KyZUj3mmP2Xm4DCtiig3H2yXDUHy6rY+cKxi1n
R6UxkjCbI02lnKFnYeaLAdhkK6RELnzOCxyzryXAkRUa3BgtmcYJ8e6WsCetiaEnhflFktrHh5b9
gJB+PsxgJt+LRosqoCA890YiHFVA0ORwY29hRSYe0aymIZvDkFSssOJjgkun4facZRwlbNhWUdoE
NZvMueByPftW6lEOww01BmhxpdUaIekBCTxMAVRa4bJTmxG3p1hn5cXRqWFVmDRN9lJFAar6C28A
SCWZz00h8L2m21t5WAgBvxlu/6vPNNHV8LG9ApWjHGjOOzME+J4+wz1vJCLgv8JoWf05uUctZVrM
Ra3tjS4JGEd/+wbFb3kyUvTwnDgvgHaVpmn2HrHVdMkQ/G26ygglrnupQpR6wglGnmx7TraCld0U
Kwr16CQbtESCqzKndNYRm7f6plkEjeXi+f1JBbTo7gnLcqQdjEodE7vKfwZV/+T1tA+NuVripU+i
M3hGTGMN2wrtfV9g7wNHGt8BFh5a3YuCqhyxIsvwaHP2ux8s6WEiTDAwE400ZaVuTDiiPGUgcWRh
gMpq8IqjfuhvhrypEOsLT+ajFcJmZ3UPSrZJ42Wudo9hULDXlafff4cMOt+ZXwMo6sVClWYqH4Hl
N8hamDsy2WlsrVAqBWZUQNXZJL+uSisAzXGRFHQ35SJRgqBI7dUd72Q05OtAyAI+d5NdPjH6iVF5
fKr2Ke081SZk3op3qYmtysEP0RVtkVfvtDKx014R8gP5752fr6ZsE8q6fFqVoVEtZStARR0kDPEM
IL7X84RLPOLwGg8SOLU3TB69Ff2sEkD4ieaYS4Q3ucWrRYtKJuLgX2qxQs50erdlQLgRRkRZKbPp
PvycbITBThxFtXhdNIrJmW9aTg02NC043tnr5CQoaB8lSEEXN3eH2AC3ZOiKtoMtyutId9oPj1Ev
JTZ1JhCnj00dXZM83hnCCWTe2A/IdNMQ8RJ27KaxLwmV1rjP3jhSeRzuFqV2LPne+VmmihWlgtWg
ZJdbFLzEACbc5/iL/aVw+/5DT0po/OSl4+XkGy+0NPuvFx2M0rRkJOHWgjcTcJ4YZ8/2E5eXkMr6
LQ0Q7JcvZu+Apvv/w6kpQ0M+4yQm1CX0nMeBxO4qgaanzqHfm9viffsqx6vI77JLo/GWcpbRpFp6
aUZPrJYcq25GOrusl7mU7mZrHnq6AQP/ss/G1QhzMdxvoHfaI3elRrfz94pKd7vjG/gChobKTZN0
VoPqDTod8JhwFXgY44n7GdArp09e4QBOViR3nkITdQQgO+GRGxIplctyLFnRkIS0ZXiDEjecQ0oG
crVyUoCP/zt1AflVBidh4mN1gpjPPj6uwErTVryIF6HnV65txsOJQsNE0i76A5m3VIAMdJp3Kf83
msI6dSUwkZXiO/pQC+R8CUG45G+pqED97l1+qbi0bLMunRfjAyr0Xol34Z/h/t2yzzYMD8r1QdlH
GSuvIwtpGybExIfGjUpr7iFVxlMeMTyeMl3mzNdqtyN4REnG4pIOo3MeAlODuy3zNRNThNKHyPGm
8TDkN3TTnyGQ9TIgkuEEycpEdGlgQxQ/QgOd6pEKGysC6fDUaU/X7B1p7/8WSf+RG38xekWS6kGu
mOdIhyfZk2Dsesbz8iBuRbjyUR2uf5VfMRKUkDI2ErDJ1xuHSCD5JPXWulbYua/MswiulojlxK63
PhhyxNDIyoMAdYFF27RybIb+HGCt+YT+/aI+ojc6Q90kRUrsotpHwr7QOB3XAvEZ9ib/oVdY2lXj
jJQfLJIgKNvvUmnJhsJBJOR4sziALCIfOZMAMwdyVQ9TP7PFe7VUPJ1V+l9s287c71r6WpZXDqG6
hzxaoSsHhXndRfQaB7mcF6AL61Q6Bk0Lg9l6ZImXeUQZfDW68vJyhyZgG24fNzMoNLHzthYRLJuM
Pi6EGeuuuOfPNrPvAhEGbiDD0vV3M/vtjUftLnxEUGFVBKUbDlOXn8pakbpT6MzLV4bsmtLodLyj
sVkVcV+8Ek+Hjw6UNnLl2G4EjbyVAVEk+wfXBaGFhIaS223QltgTEkv1qbfCuh2vYQ0NgYahDS5/
HBNPwy4WZhPRsNr4Iky1qhHUA8DMDh+yDKy14dMIpXnaDT0JyltetWEQR3AuV9pO58KfZeD1kZ86
zz/CA/DnLGDYlDJwRpStP6nVLj6mi78ejDkLdvtzGF708pZZSgGdftHmklLj6ZWDBEyJa7riEva2
VW1W0Ycw2epI9bRF3EgBTJ3mHRIZp05z2IgkarjHF6U/f7SpzUg+LQCsBYyb13A+xJQ9YafsWuN5
dmZ2FjxzsvlG604FJQFJ1DKnJVCoEjnfU0tZ0oCz2LiKkey0sr5z8o3dYhKzAS7jeT6fHsNEJcaZ
PrJG7UmIzX0ooKcid4IYdWPSmTIBFfr1EVSBzqHjB9IK4XnFTfB+GUw/7sV9n1yL22tybluPKK5f
QnJftmMig7WnDkdPSGwZVZzmIgbNvciGUk+/hgS90eAHprfFR38As0kfAjQ26blc4VMn5Z9pjyYE
dp/YL0pjOQyP+DYE78o8Mg3mRh0kRBp0QQ+5RywC5oU9h3Fv3VaMHtTdLRPqgq7yyeL4C/kcFw39
NSnh+o1YQ9el2cPap3++95EDnLxy0nnfxMKXU+Je2B3U7y7TdP0xRLHxRfBnGGFDA+wEyy3lkplO
/5AUg4MOtc/8qGnjiPyUTmdJR+eN7ow+2jB1/KNt3bL6UZKujNAPfze3EE5QbZS82gpltf3xoDzg
M5iRyWNSxG8GgULe4k2oV6z3lIKOvp/iXSAcGNn8QvrRLrMADC1NMyckhJ/3X7EG8KiQqKdJ9+10
ciuk9P7PVTCDOp7775mibcW3DuwwFOd2xMPXHj/J5pMem6HkNjvHbYbS/ALrM81VdZJeVGLsn3UW
Tj0anUdjxITbaDZQzV8GBKwIfOiiAxFVCZLZMRl/ut/nJAyrjjZJmfEFbqwUM0W0IyCGGsNhv6SJ
NafRv++eizPpi2+amElHqs384B1X1PBONP+t+Pzpp7Y2MAIJJ+7ra99B6UHRw7HmJr0N81drXEd9
2fP7OQ6cgUo5EPAYV22L8Qs28Nu9UB4zaLzybQ4Q8v0fPX/2jSuIj/AonhcnV2+ofeTBjX7Tut+L
dRxkqYEqSDsZwPa8TDwQtqyQ5nbBkbiJJidxE/mABqC/jY9eQU7qERAPgQgsN7+JV06vcJSwIm/l
UlpoMV1cq6ql4deGsDnpd1SQrVLX32F4FuMXyZiENUqGNkAPeMN4QW72RgWBZp4qp6rwib5q+ali
LgGPdGcP08MAp3vSEbzdl5XkrJHP9emKonnVF/wcGDcfKaB7lA6dQfEBlGYBABwMqQuekO1sgwfJ
ASkEGZWsAL3f7TKLDOycCk1Q8TLQ1nDrR7xeEIBw078SuH8qSc1aYHW5KW9XhM2dE+lrJZNQjO53
WoMi7j4kVlDBskWJqKPWmCV3AEXU/SMut+vh/EU0QJ+ZcAvU60YVgp5ZG/ncPnDzc5up1J6688kx
9/RvHxtwcTKBUIUT2NG83/dE0K8OLRRuwZB5NBn+p8T4qgDMny9gus60xvCDTloY5yN0qTc3vTiO
RQoakINYziET0Etu/hBoranJaTW/BxvQ7p1yT2VL9+JILin5pt0YuOTzCGoBqNCNUDwciOa75bZ7
yugnYyBeA/bT/2A0a7/Illfwn2xT6FvVosVW4K2b+9Dg2RAdybAjs33vNAh87d/WBEDG5dW84+iC
2nAViQ+q+6J5NChtFudPbbhWDU4fpPB9V1RQU+L/o6kJ9U2WikUzdoTggcQMJpRHgwYXdJKighFW
od0JGxpkyNqTtn4v3By4ug6LRxmGNRlZijCxqDm2LKABkexW5mfFkVNyNgENcjbsoc2kgQ44bKKH
W3wR9Pct/vQ88o3zaIyqSHob3ENiEO9wo6XkTREA8U1bc7tKXY5EL95PnMewZ5ORVt0yCtnklkyD
ZrfpZGmmj2EWJz9vnLxVZj2vUk1XW2rYYUptksnfPrlB+7ivx+5JRZfVpDCyex+OzhQrgS2Ni/VS
cDl/MgPvBSm9ABtI2KyzD7Iof6kYPWLK6yq+WRZbjukm1cf26KBvrOu06ZGT2WAtYMc6sCUngJfa
h9G1q+AwyllhKiAyEFCnGlMIOpkzlnNlD1VhC66x9XbHn3CsAK5J9+bCBhmehRqbU2UKW0U9PhbS
vMoMq2GBhxznQXYkw8CNRFrnj+KHTbnQOAfmkI/gbc7ZebScags1/J9IJ+hnQjRHLLIkhwtvg0MM
rltdtLD6cHlKvDp9Wybx0Swv66AKWoQZjbn1oQ6nrvge4TDo2ZmeGOuivthwJJwCc/pdaYJbN8ok
Dk7/qotlR2JTCq1LIlbkARChrafvbFOXXVruDuE16SYGO5CqyR9rooC2Xlue7B4vktvupquIESYA
c1lhIj5bz9BRhFqyidKUBQ5cxfQ4b05IMsg8CtNp4OxW8aP8nbbfmxFzBvWoFpz91tnboYslI1ON
fwctNxXII49bGGnOORjAgh1dfSP0U5/2kEa/eHReAEXSsqn/Zt17xdU/Hs4opVYhxD0BDsoPyn5v
wXx998cxHY1MjWjtyKhA3Ox8H16KK8AHcUR15OokpDob2WjXE4CDWCp5pNebFb1jFgoGHBRBsll3
MjHKA4FM6IWefF6q6G7zcNcln+kUykTsbgKlT7NhJGpBL9HydcoU6heEpy01JgIiqjOBceZQ9Wo1
HApj7npPKaAt3PWIgTm70TbLMIIWLorozEQEI04Hz1QmbZTQkX9Ismm+P5+5AsS521Cz0gLS/Qp7
mpJ48jxQzZcAMSMAvgPu0HLx7m+gwfsQ9baLTjUD563ChV+XPGgcwexpiwlH6h8Xkopy/ixnEjeg
S5NCR5S2z5nzVx2qoC+FgZvr3NAvyesSBjW8rAVXoVIuA8buWuBtcngemqBsHSzub1qqySyd8Crj
cufafTTinMmZcwsMc3wSq703bC2NN/1pXPeBFuoXlgx0Sgd1/q/7wxIXxdPwKicRqXNJFB/KiywL
b4B/7jLHTp+v7X71PgkqDeiuv7gdzfXhk5sFPY2jty9VcIALIGgG5JHIS6cuPRtc10QR0ugWv+bv
YWU+ArV+tBBN7Jz6ZbJCN8uc4C6PLqGQPbg1prjx5COwcEajCFxEW04pw7FC7J2rByQdr4j9T6/h
7UB4QmaF5BN6/VlSUW4TD51GUrf2aim283gnytfdlIfiNs8HWL32UADG0y/eJqjTP6gYpHpHlRdt
3kRzyi43cYBqWkjhvA/mJW46Mm/2OhkOVrtJOteIXRc6GKQgvRazfTtc+BsJ9W48hmenimB0oyHG
3Xd1Gx9/7twZySEXghAtQkqgzb8k6Rwg0ZJ8Lb85cXP5O/L9afS76X3CofQ1rqC+pEFOQraAFzXB
TdKM0AoDpZQePJWjmuWlxrG9GPvkqd2e5M7Jj6V722QpJJog6T/AAjTwae68wEZH6S450T1qJMAa
M2cLbXeAydqBrv7518FV5tfZ6EbquNPfzZx3ZCK5RO3gAyO8y8up8hxq8wU2ZprZ3OfzIhZNa1xr
W+CScPt3Tj0OWxZvDCFV0/i+WFOr7+mEoJeg9ajqh0ABSw5dnh9p2xbRELHgAs8E/sI9+PtWt5o3
CO+3Woy+5vDoamrpmIMaUbyLb90VEGYaaneMFHQ5Oren8Oz1cFLHRV0Gu0khH6k18mhYdLIMneTt
asUx7eLaB5ir3OZbw14FR83+jMcGguOCtYOtk/YsyaR7Saq1MuBYdjCJ8YhM1zh7xWUTb0f2q4ws
4J4bwUHDilu1RjbTtOClN7dAwQxI/WleNFf25FCusm0bFyTJL1k6gXqEg301nYKE3f318W+Uv+zt
rO27T45fo5JSp4K2XXiG+a3qRR7+lmkLAq+t8R4u3aXkjULsvUYghTNfMFsy5E4HIFL+rKWXMlHp
Z2UlhezOucmXxj+4IWedL/njSyMML1eHQsT/QaqJJDWSNnnajgsUyR5C5YfbwL4gU88QYUaTxzCg
aCCmn4WAgY8/OzZXvadR6zh/Lp5cjxPnAK166WD0tdXPHrf2cJlCJpAccDFqdzwUPViYzUKpCQwX
Qj/srRtzmoQ77N1Ytl6gTZrHruw2ty53QBC6kZNvkru6Z8BJ+GGUzErXS3fszM7k15LeWSRraOPZ
Uo5SbqH6CE3afFfumJKw+NzYu8dk3fHOCARQ7KPvU7552qNKpuuQUHrvIgXumc4DllKli/ZSZ2QK
DnQo56Y38TxgVkjt7udprJIWKgeNPNN3a4derTJF3jCMbkCToeyOeE9NHevBk4ScmKCMOtAkASrR
yYr9aLQh6EhOpNcgEIqE1aIj8QfFtHDOKIQf+NMWSTMXSAFkBfysqCUhJS3rl7EPIBLoGpHYJSki
eDa/8mFh2528Oxm1+wyWp7rkyeYxYHjeqn0VgnqQjJf+1+ccBD7LTztYZyI0rcsI5zXI2jnLVgq6
RVQoMm1Qt8oYAtfbKaEosG8b1H7cgBHG1nh/nOU1SpRMepqiw/2tkbEwRA17ewExJtOkKFGzuMln
HG/CYPK0jpZzh285Y9bXuIMbY7Hs6T8zwZD3oB0WlS3uXEYrbbAFQ49Yy1QsKWxJaKoA+bMqZs4q
Q6Fz19Cpjoxwi20m+/7aKCBDGOWvOBYcMo3m4pb4ltc672XBu2XNXY5nC3D5OX1oksRQeLYdTSF3
/qd7Y/EiWLRj76q2+lTfnwN+fD0/KVc/7viUUT9kAVZl1bRqqGB9m3aeAZHVbKdmA+wndR+8c1v3
C5PQsDzUXnYU1ATAkJXnOzRMu6v/HA6b8kCH6wfr0FsqUHetmdoEquT5v18kNgNZtwb3sGJlZ/BZ
xZVp1R7HuTZB6RCQIkLXrcFFW8UIkqpOY9BQRdf953oOc8C6IloUwGanC5KcMhnWID7Z2cM7luOI
YN9pM4aXsJpTmKUNByb/FshN6xAFBMmbi9jCuI1s3Mx0P0hrwKO9O+AD2ofaClegsBe/04nKMzZ/
pKWzKSpACNeudURAO24BFuWKGs1NarV5GYAbQnK6xa0ZVtsnF74bW+ZfXGk9aa+0P3r/JGmMqoVl
H12ASNwo0+RDcJrPVD5S42YOAjcVo8lgLUEuonsBGr5rEQAN1efMLeV2j+v7kZaCS12BPSOubDlk
sG3zPCA01myCxXvYVKbQ9XVv4Refx9Mwtg02Vf1GyBTrm8Cno23jFIYt/qdhESV4tZExcdGTVY+c
oKhTe4pGtO1YLFzfz4fCG/lpOWh3rUIKqm9H+ZK6qZpVFgQzmu5Otk4jjWyJ+ClrtD1uNVQ9UUoP
W5/2iOa6JqEx0bkAT+ioetdIVO5XZcF0ZR2sMtas8xm9cnnPQkNE/PngjjNMKNpZxk6prBeIiT8v
FdpJ4SLxjqF4HR0zJzr60yklwEoZ/B7nOHztY4IEQsJoITV3AJy1Q/BWlnPqy+pVBOpGG0Epin+/
JuhYpkrZSQsSR6qkCXYR4dN4lpHfY+gWr3G2yIu6OviUK+xzBMI8dnRQ09anBNzuOPDLNmSa7V5v
RBX9us0sgmvRslmisB/HgQTSruXY8iIo1JCTeWrBLK9fqIYUWs26rOf5mcQ8F1PUHDtsrVM5DR2W
/Xgw6Xtf92Qil6EhYYRTzKMeTumv7wiUEBaJ12J/MHnHwHJgvA8ANYxROiUZyQt0YRexQlsoJCL4
x/yNnCnNoj68F0QrQs46JmtK5VYBtZmZQXcSIRLcJ7138ujfqQ1GbWb5Yq+1Dh8QF60gSB1R4XPd
++UX/AkElL8th4BbfiEwukoKs6cEcSJrdkQWtvkXoYW78dtQff0I46Dnu31GPRCWIsE/4kQ4OgBc
c1rrpaxhIxBETNU5kk91lpypcmGBdexzYh154u4kXSYhR+h21OkREhiQ6Cqc2MfBlAkO/9bRexfD
9Tb56AZTBdsa0BAxasfVmFsN/fKECmZPLXIdqqCG7mHEitVwvwL+tyosuLZ6y/6ah9xBrgGLaopm
FXqW/plJISavouQ/bupa1fnDJjTGKh7ursj0EUCYBTLeV+j1YwGYryjKm2tMWY8piV0G1hdj8+As
xVSjL7uEUrY9a6I3gk9Xkgq12vYmZrW77oFZCZa3cuZjZM40S+G3wulx+Z6a+4pnPqPk6cIYNmDh
VQRH3EnX+euszqWpoTuekbJpjA2I7i/qCjeAeLf+9pBog5hMKfWAdciIdXBQd8OtHZqJ9577kxmO
/cFscbCLqWvHkuH3DP6kl/s95QUZpWOHaD1O6e2oU6biWaguiW2q49go04O96OpalBMj1/TMvkDA
9Z0nkHQOdUefg+SC3lMTvubnqDtMyk0YwJxZ/2hYTsFfujB0SnrdHHJYD7IX8rHj5iqyxZPQbCtZ
qrx05uNjAc9375JG6OrT7ZZOErQTH+3sIuNZf79G/bB5iMA/oT3utwizDEjslUlX4ODpi0ez+5Di
wGtWhh4YpruI7qpHqSHuaHmpu+bhnOEWjdIgns/ROjYi8oljxeTcH27XZS5GBYZ1/mcrNaftXfCi
XV6DR6iYmItUYGg7afFovXQzGLfqtlbXReA9qjKHFddtTPVw4AXdiSw6/lZBDkEhljpwX7/jwgdU
xp0bfkBtB9hzxxXrme8KHLn1WAM6n1yDmJRSdf3Z5Y8pM6IrPlDteD6e/72wf2Zm3vrGeAc/q1oh
YbxWVxtNESLShVUlnKRZOIw0xBLt8Tmbsg1wXpIrBMDt8DDDKJuv4LfFw6ETKCHQ9aiO6tG5auLR
mumE4Dz3CX25rUIFXnkfIzFEOiwllxcJQ+pXnrLd5UqRTLZDzwNYmvXWF2RJlsHuoqxVev5CHhLD
FVJG1HEPrFv+72oFjcozD0DGMxiFfGhtnIzlGeRUj0FVaBwzdCFEuC6EBjGnyXX59Kfin6EVSQKD
xaWxXRDIszTl6HiLEyb60OrK/RDfe8710VQkC/mIOhYOEGgqBaz0RzTM5dHmDtga1QrtYe+8lDnw
EAXA4IF7OHMu+532zTXgsIvrgtiOgQUORPIP5amxMJhgddsx8MH3Ethi/Vj+oM9bJa9pUGBViEDp
ddiGJeVGf0I1XdiV9iNBX9RBQq1alsbD+ZTpxjydYjkVimwRNAq0fjuQ5tjj5Hwlc7ygMNsb3bgH
3O0j38Udl1SaPQFQKpXq5iBN6bTXVJyDteElwfRBl3F5mvIkPiMifCDiMYtz+82ZqNqYMg86jrE2
XwELeumNi7vW4TRXh3uIHmSVMW3sAD3R98MI2R4ketnvirlkL5X5ODUaQdS3FWFtsdJ9AMQTWyxY
cKB/pHj2MGVaXDbtd8VIncEhwZtsAlPqFhQ7NHkAOEX2noTtyr8E3fzGK811CdgJgvOYd7Fdmy6t
V1IghLCXruNgAPljiDYsPRA6FR29V65ApxitkxDFu7LW4CtbdRsB8Uwf4J5uEyWVK0uc2JJKQk3N
obUZmaszLCpj4eWmg+L380pYeSKl3S4q5R9qc7TGfg+wB0xXYdmOe+D+WHAX1X3wWVCqSiREJHnq
yXLzcq4UMCuo0JIDEAYJZxQqe3qQR2P4yxnk9RDFcg4+DwShddOiwf7vLsMZGH0C4gk5EEspYXdy
qzyG7rAWsAV0BDcPgjr1+Ee4LtbYUOE1TkB/sKaOTl5jdLKTtreGvu2+YK2HR/7MDmAaxPeSlymw
V/pZg3JyNc8gLq6RII+Od7k2FMm+RBA0gmj9WyimY9+fgpmUW6DV1cw1thTaHW9f9tAN1Yk5FwnF
W1oHDv5lRaDZ6ttwU8ehd7rKMwoBBGwlt2q6DROjlpheAbSXhjqt4q2rVFvHvDMr9kzn9PXpTynu
F/nkDZijfQRosZsVJo96KeeX6wZ6+GgSFSGQyaS8Mq03UkOVG7rULLPy1oeFCqSrn/5o5rcAiSQs
RnCI5o8NEyhSCvUzCalPl1MuMWX2TQMl489/ol9UQ41P98D82eV1YF2viwt26XUPVhNn2HKYspCC
u2kFOoIeN9g0pFPseahcSqpQp0ynqsbIQ+dxcVgWFeuxYXQpzz9aGhYEYi2YwVuAPmNjYqwZ/wwH
iY+j4/gpIywg6jIbfNegJDJoVh33qdpEXWZ2cukFr1j2pD4wZnwpeAHpKOSzZf+rbnt3+AbPq2vT
V17tYeZhC0gK3IbxZNGLG2Z9kpU9urWFM31xuB94F82k6iCW7Tt+k1pH7NeTN26VMHhXFiljYNQg
3Z808po5+L707xCCLLkgCXmWdUK/w90HCtU4bDAJhaEKP6pTZKO4DWnxR0eSjDBtuzb7/u+NI2xB
vFdi9oc6c5mPDF23I4pYMkmcJdaWkGKvrS1gkJIrL49QPn8tQIe5Qb8Hchl/s1cZ9adnqLhG7k0b
Jr9ULnSOM9M5HKbr4Ys1Ho2WLfuUTUSt/v2R4KnF6YjGxlRHq5Bw8nOFzSpggeSL1QqUt4705wR9
I/506qNohF4+6XurUA+fivEeJZYyrEpMc1jAhWaCYr3ThorXxwqZJ/Ju6WVTuz4onyVatCE0g8ul
OtEDrfjjn4uOLt6fj0qm1o6i2sXaAG5Sy1CEy/EhNvyMmNAkIVKX1QC6zBox7sTtb+Yv3fQcXHNl
d3/6TC407EQdKG/xRq+U/9IpQLgbo10fs8nZnBZeZuVuj4tCF8fefd3e/VzshOzG5wSg1WYwAf0Q
1h424nCWC4RHg4azU55DcABYmu+WbhMw+3ea1ovzP/4O39AbWfejUYPHIg/Qilw6hGGaVN1Wn3Cx
TehXe/Xx8+QGUvwa0qhdY5EJv4rCN4uDJa3Jzt/M21o1o1Nwvya6oVO7vPbXEEGi0tqdKxB9tJAG
5xU32bmkOrcu2KBy3Jh5IlIkNNvlWxqiuYNvKi/33H1tY27QOyBCNzaj6YLy72tu2VC9EW0/1Pye
zlNrcvptACkTQ9cu6F2ycQoOCmv3SDSZIjmJcSQIOUihOzVNbAZP0v6pDkFXnvB39kEEkjyyaMvV
X0eSdGBQRi1WeymMj8KZ3CBy2K/yDC4FTSBN+NuHA8q5lwjQMFOHcQ2+YfC9bfGOAb8vaJ/T/S8O
PjLRj6VPG9XlMCXukzXuqG48xEtahkQMHzVog8AGAd9ALfsyahZHZ0og1qJLj5c6dLEthBxqNL/Q
yAbQE7io3Ud3rUXBOl1+Fo64y29QLESCbNxG5K+BlqFpLMmIITn9Km7+z3NrB65tpZg8OskUp9ZA
qSbH9HKWKase0OqGIVCC78zuZl6quTRGRKxpqyQLW4d/qfUC7YW0CmHb3cC79/J/XF3zML694IZX
6Yppf+4g0jM7Sa6LJMQJamicOje3LG4GS/Pz4Qsi76NFIn6kdMaIiQBDqTIKNIvCVF28Ei7pxhYn
xuHflRx13Hf1UcnVT4YdIc7JjVnftTcndlCuyOeRMPCu0xQNM5+Fnj4WW2QQHXcXhi6S171pzytu
sf4zO6F8hFHf8D07LA4uwjIKy18epv/AbBXL2soFFeZYkRK+9X83k3y9R/fYEcn0+iAu5LbpK9z1
V6EghwWZ4CLMXj4PzaZBQbtMyampaP5Zthx1YNsM8o1bPLcbNpIyHvmhu1rqjLlgeQR9M85gZqzM
o+J5zT+lq0cYCk76Hh9xi+rZQTqMS7f4LbG6imbfpK2HQ+IcsV2VC8SDnJ3cT15ZxKqpqpXJRFFb
1HgRufhsiEKIiodtgSh/Ix9mIG5PKtoUHJtFY62VOCb60umAnjeKrOK9SpVtjn6DXdd6a/uUW38d
Hplf5HH/iZsyxowdrNiI/TgDxmilm7Sj50ytHLPyA0XUc/MStxe69LG5dYo+YlNB4rEDZlS7J6Je
SJ+/SfyBkz3iVXkpD7iDXniSRLshRodGmk4FN+ncbC9HaFu5zgujiPHiYrMb/uCIo1srsXOzh6qP
g4+5Nm8KlUHYARm1QpniW4+4xYGdmLVEd3Iymzsr7skNFIYn/xDCutXPOq65qwPmLVdvPf053yrq
nrY2res1nxB28aJ1ATp895D3EuVfYic9uBToFEFj1Ao6OXsmjXMyD3vry6Ph0AMoAyzjVRJFzHZQ
IAbFY09SaofU1j5V+gEEYt8aPhvVEPesIGOajtY91Q0zqzdqSKYti8B+qz6SG6d++O39UJJex6yN
80wkHDLnksF9wcbBAcQzF+EqafDU1PgkGQHD9XV1/yYbEoKs1Vg9dvHCjeLdbA3GhzBtWeBP5grD
qe6ZDajnXA/E+1m+Z41QFk9h/1egULZBTzSaghotkV/97PNtgPIU4GucfB1ndIILFgN0v61lt31v
N5EyklacJ3VKpWy4DnzMmY6gtWX80JmbcnYAfF9HW5YKIQRHo43RRh+D7QRblSAf2Po3zZsHfkl7
ofj0NOu2BW+LDb6k+VtSdiIsF+qtr/yRYzddqY/Z3MAXVjOWv2SOjuzkTZ1qZfm2K7fpSRM6F6QN
IvusVjzz/n/GglFapClxEc3dJGoLrL0DPDa8ymY3G2vL4uyfULZ47xCQQgkm5UV8fMrlCgv7OeU0
48QlA5hwoL2M2PFOiCdKri2bLWGQqRMg2fuGwOVF/gOSXTXGt5aUdCewIv6qC1G/0lSJrxtqJmnT
EwMnFTkeJ32c8PNNVUnnwfqLq3cDTBf6VL8chzuJjsuHbyZ/vxOskHoJyvbWFNwcsaPZavnvCKXN
uET5jUG0oJ2kc+yc2cO45WfdbN7teETmcJq5Mj+fgza6TVQF7gW7C7K5+8COD6ZHx6q9k57DkOlw
UXJhdyrn5M9BSGAEY1Ikr/d1u+BzDMlbATtdBrKAiHf9MCMjRD1MhPSeFucExprCEfXueeTzcd3F
RZzEEK1eRgllCjZ9ymBDwFocTFsh9n2Paf8UqGr1oh0yhxAi9rcrICAsb0FiYNzPURbHwzHg2lKm
mX7zU5XGOLvup/mJaSWqZHkK0pQfLFOgQNR5KXMk6yc7ka9KwwGZsLVpE2BEDKpGpJCGXxFnaqmR
UBllsBrcyh7ejjqF2L5Y57O4rYpgwtd3WDMde+EMH/0PFRYmWVPgxLWJJBBQvLL3+W4ss4QRIq/F
/L2oMDi7gM9pgMJntxYPD/m5mS7EColsP0v2swvW9qsV6n1RcbEg62Ta/2CRJLjYeM3l8AOFP1Rd
c5lMIStNgN1FdclpB+lh7EUEY6dLGUCnS+lX02N11GJAWJuhu7Z1u/6FElP7jghr08texwHLQnRV
Pal0g+Y0S3ftCCgAUjUQ+Zbq2lyJuxllDZ+7H68vju8qnPnmD7ZkjMasZ4cHP2qxT3aApyEvSqmG
5l2b2C8Z4xo04Db/N29kMH+YOs8J5hmdnqlhjWJLMdEpumYH0zRXCdhbkgWtR0O+T5npjptwoNlT
vvIZdJybxcpHtMtour1Hjp9NNfDtQcInOEUEUI0HeVsa0O+aU5cKijvs5slI8SsliRTMTcckQ8k3
DGHdpUmNAaYzdk7GIA/GXhIFfW4s55n0o3XR860EeEt0ndkM8UPRYEFUUQ/C7iLX412CdxFVfdfw
LnCqiXymBj3oPUkbwDtqrqMn192AvRgB7johyD4jRLu1ZTiZvAeRHzZqk2Mf2Bl72ScEH3ntnbEF
AMEj33piVGjgcqrRdVZ6Wnyk7r5TSZ7qIMe3kPJKVnyN0iO+d+g6XAloHBrBt0uxBbGUCn3lZu5Q
XJYfQ3FwaazufZ6P0AnkUyn703KJY5FZRPpllU6dMRnMeaoXnKVArerkjypIhDTCFNlc37CTyueY
JuKgmNQDPLncIc0U1T0erLUWqjvm5fyVud6F+h9+OLfPhnfBmZ+q8C5Ilg5WHJehISMo4+dPPpOX
FL4R4Gb7CQNdxbjY4LJ9fiimGgrIDcwBcD8D2Du83xbE3zk1qjKXH0kJAH/FMY4+J/He+Z87i03Z
KYSNMPPyL1QemBFOM50dLOSP7L5jEyDQ3t3kPWBlIgWZQUCD+MTbzfQPND4HUM+G5iZxUZAugghz
f/2ccGIPUozCpRozT0iq/s/tbFqvVywu3K//7/kmy51CXEkPmL+DX05ryCTdb+Mm3CQ/l0fE4KKU
YNwMPAC9VIaY5pXp2GDMQOslc5bVufmFh8c58+UXzH9gj73wAELZubJJHygwSvg6Lb5PDGamdRS3
A9fiGOttUUf0aC/XWQ/vVIc8qpsyh+pxC05puaUPpOLYEi1ggc2Zg6TvSdDm2cFvQ4HuPVl4l3BN
+iR+H4C1luskGtIt1U1BFw0qoSqgMDvJ/fKYiK/xS7iaPEmWMJvSVul2UeGmwMfm48nWbfXHpGIK
XMThmA4Rmq8fXRdrtNgyJm+XAQtBgnxgPTgSEmp2sJy8EAX2ISAJX4YnJouqFOcDpcIr2wEROCMC
HHadc6xdL8jbWoNjT8/PHTK8o6NWpi1IlPjm5cRRBLgLZ4ovwH3yN+S1TIp+NpbgKJBjQJSAttGt
5uPPPORHhRAwgWnasBLAJZAMGip8JhIpmj6Y85J6SXP+MnYg5cBE2Sf0bYZ+H3JOTYm+UYlUivta
T4aGlrZdRZCfGS0hX0xk6qQCCQq4W38iEGIO61qMIoQm2PSTbjzuhaLShl9sKuPCVAgvlWy1iTX5
fvPjF7B67j0VWmALL1uYKTuuzg6BIu0GnUcBQip2dQg2fSWq+g17nwK0jCi4Xwfsrnor+OfzhCIQ
YOxOWIvU1WTD0ntw/593j2HzI0EcTWuB9VVvo+3TDizf/AYFtYksU0HMMWOVTcbjW9llA6IttbwP
/efxGv1cxxEdKKHz6J9/8ylU6/YWLWq7yip1hUMLas+wFZeTHLzgznung0mvxUnIZ1mc9eM+iejS
Ea0RqeVsijEzNte4rnlha+hS08sG+tB5l0TMBrhEEcdaTEgHviNfZGnMkqegRcYDuAiB4+eqKeYD
3cCInmeIAYwkRMEUZuxyedPERygMYtDBUncuNqWoGm2CwzUypwYIP3RJPbrNg87HmIzBBTOfJtF+
6gG2draY1n3iL2cpiP//LGGAjFr8DZoRnRoHPfTCqBwS0tj7kLolkv3vM7xPAAlNTIcnu6ldKUEK
gt5TNLd43V8JmrLKb5MKbOxNwsFxXyaO4u1i3l7H4hYDY3FMWGJcRiiJ5qETHYg2jT6U5J9sxOMK
tJWbxluoqHoo3qss4+pjunosq0KjtBLfzj2YWiHvSlbFk/DXiUgdcGVvh+bNn2kNFunylKpI02EV
tbemwgG98874Ynx2KUbRueHq/nGLMZYKk2ZMMTxdU6V+UX4XqMCrN77Rrge7YRocKkpbxiHMMdza
kS2BS1lNMWLcvVXa/ZsL51qKEE4C5QJPgIAb3AjbVmLVhBPwO3iPGFsRPOlD302W59K0mjpob55W
UPLCAOA/i0zFR7mCiFBS18phTNvtzh0px3VQ31Sn1eoiQad5OIx9NV8SAjFjgraUNmM7oSdDz5g2
SpBn3kXipMn0BQQaoY3oBO6Q59FKPdr392DrF2c/IZB7uzGFg1wyGMdPQBCbXXWY+8irtsJ0kZcv
eGoWqmcaPJvuW6YLbSnTbxMJ9W9VYFoLgbxAQ6a2cExB0CWMB1Y35ElqeFOx3bUCy9uOnkSXlMrk
X4C4pY2k7T6yd929/ZbNFWkxZpRbSRn1ZNc7p00sNkpQ4hu6kAqxYwp+7+UP2iDOENkE2aMdIIlf
4UGaOAC7xYc0CXiCw47UwiekWvuO
`protect end_protected
