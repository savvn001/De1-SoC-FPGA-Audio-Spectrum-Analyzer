��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl3y�3�P���Ħ�i�X���\u[vW�ư&�	���E-u����b#������v�]4�L�����5H��[�������O`�=�զ���)�uJ�VB8�ݢt��&� Ϲ��>m3�ZXN3�Ӹ�f��]�N�-�	�U��n.O<��.�ue�Rܧc���~�X���/g�!іb�����������:��#��]"7�{������&���S}k�f1�,�:�'�!�Ps����z(��;ʆw��i�d�M���y�VD��.������Z�KkΜ��{`r��}j��.�?�d�p�J*υ�|Q�a�����h��N����d|&�V�+�5ih�A�W�g���V��B�4�S�4d�vH�
��l�,�ճ����l�=uP�E]y��c�&þ�PЧ�=Z�yWj\��(�Q(/}�MW��z�����IМ�8��d{���t�� ���J1���z��O�K����}����p�n4�3����>�[���Q$j;R�T��ٴ��& ,l� �ˑ%wl�i�/#�~� �vf�S`fqۙ|ɦ:��b@�%�&�C���1d�w����P\�*�:Ʌ� � O�c�尥a>��8%3y��o�0��Λ�׋�(֓|�X#Sx<����\*6|r9�/败���=�>��[�rURoP�;���?U��Awl�n�W�;�XCn��"\Ѵn�KG�]��k���MI!T�)��S�&VPk����>J�����ޏe�J�}��52�#@����[DM�۴�̀�����}������}��E���*CT���$U�i{��Ek+�G��a�Sg�����ǝ`(�uD\� sk�ϠW���*�n�#���K��k61ei+lw��ZW��rʸë� �ݙ����&ȼ�m���Ѻ$�k��^��B��P����+�1��؍|;#��m4_�����ǋ�Y}M�3\��f>��bp��@�o*>�*%Q�Tl��lų=f�۔IC#���T����^�W٭-�^w���#s	������D�bq�2��
�H9t-Y?n�IE������x&�w�?�ܮ37�mt��p��9<��.�Sc#�]:�5a�]:��*r���8�rY�DQިLljZ��:H-H0�*�,O����L�V>� 0�{�����8�B1�TY�{K&N߷&|ܺ-�^����\I!5����li���wB"����"�Ɍ4�k7a�dh���	h���}��"�@`�q�X��ou8���ؠi�y4������/����Z�� ;ӟ_��14v�D`4Q��9�D:Ω�%�!�9��&x�bM���"I�|�8o�fҿ�>���d�:Mv��6U�V�{�����������B��k�H�m���(��~,k��:W�����%�1Z������{��6F3�>��Y�E��&��Tx4^5�P���M�Y�t���^̓�����1&ȡ�MM�f��,7�ݱc���Y����3]s�s.ߞ̋�'��d����!����i�A~ieҐX�A�x�8Rne>z�����2���X����FE��N�\.ߪ�K?~��k.и���@[=3�vS ��ܩ��t�����"�����J�k(a�/rA a��Z�ve{�z]�CH|��Q�e`*���Gsý�N7iٟ��ؒ��~�8pv���GN������'pz�����̛��R>2��+d�f�$���i�6/��D���BI-��5�X����K��Y>gEM���k��oX֥&ؔ
���u�cSTБ�Iu#�tXX�@�#V̷�ŀ�O?
�,��SF��y�=cM �l����VC�^�N�u}Q��鶈�WX�F��������'ޣ��ʪ�֠t�I�:��r�2�U�}��-E&ș2{5��T��ʕ`o��������'���L6 u�O�?��r���eS�Xb����Q��x��P�.^�/�k1U�6�B(�8��L��2��3��(lP�}%Ƣ�vFI�m�+Wf� �˻e�@ �r�D&f38\8��+����s�x׊ vD34���r�~�[��"�Q��"�F��p���%��Ϥ�j �}��0�$ҥZ��D�~4])���\�ae��/��2���ȏXYsS�mZ�&L!��mq������A�a�}� M#.�uՕ��+z'+ᅥ�fL�T�+�{_
_��]�b�G	�'����0�]�V�s����ڄ7Q䁲�7K�ZU�K� �h3JӍ��8��>"*�7��T��J�G���r���Z/���!�h�O����U�����<{Kt�&�<d�?���:�60��zћ������g#�򹐶L�ns=�� V̬͒�:t ��h�t4�1"�i�X;9-	+��R��
��[~�S:nϦ(	6�Y�k�PF�.Sd[����#+IrzV�)��6#O	�x��E;�[a���D/oW����@�"^/%�p�dY:���y����V@����\d��1�z&l���m�Ð2p&у����t�}�U�5��b�*UAn|K�����"��l'�k�!o!�_�v��ht~�Wo��e`�Ƃ�:��ߦɨ�����d��V����B�n����l����2-�)���%?(oWn
ţ�e}o�M$�^���SQKiCv�rԬ��K�s�f6�(�/���L�?��Ƚ� �׫��T8";`4�nB����3ڙD����^\�D����4��֛/����[�>VS�8��u��yL���*�A��nӬ� ��"��Yb{*�E��7�y[���υ��&��4�7A&�B������]랢8}
pI��䆗OH�?]qyw��=Gy\Eu�cd�v�Cd�3�Z�>�rV����[����5�UF�<�J<��=�U]=H�NH��a���y��-u�~aR�j�V�����W5Lx��[0���8����g#�Y�Fg�x���H
$�d)_�~ؒ�Υ�O�����'�O��8n��
�ynr�e�� �r���r�C��H��^�� ��(�����tn����/h�z�{h�g�ه��h �
������ZicU��C��~��NSW���\Z�ͷ�:��|d�]���V����?����f��]@ f�Y�w$�-d���/�c�����ۏP����P�yi��(������7�k�ѥ�k�=�E!����lt
���	\I՞��,s	����Cn�d��j��SA>b0A̞~{�֍�G6��a��h�{��nx^\g2�xf�����r��A�	«`<X3�D��Kˋ�Cړ�_' L���ڞ��'\��=g="�M�MF��1��σ_<)�)��V!������b�$�!Qid�i*��SC/L��Æ9h�E��f�V��;QZ��#s�U�+5�6�M�"��<�.<��t�Ѥ��!+U�z�ٯ����yy��,��z��4<O�2���~���1�Z�֍�Ȯ���I=���N�B���ɍ|+W%�eU-U��0#c��J�ٵ"?��X���E� �Q�u"��>��|�p�Q�s�D�ǲ4)@%CZ����D	�Vsb�ŀ+�[�_hLuC!�Z�{�T8�{�c�e��H�u~�N#t�.K�J5P �|"Itb�]��Ed����������o�A���9��S���1�3���o�luEs�~�&�,V�
�1�Cܥ>ї���ظ[��p.q'`���},�%����[�{�i� ��=&s�ݣ� �TRY�~u1B�P�m^��k(�����HM(��)���p4i`e&8��jB&&�B�b�/u3�ƌ�o'm1��>��̽
R�@9j�Q�8��#'i��4�s���]�ZS;`�H�Q���Dӝ�&(�Բj)��s����S���җΪ�e��K.$]��}�'�����>���K�Q����/�-��8z�v�N� �D���hA�l&�� w�ADx~�7�5iО�f�D�~�����91Z�\���2���?÷��4E �ԋ@ds{6K�c���[s�>
$�����{2~�Q
|��.��[�M2�i�%��P��0u���w7O�=.O0/UU�]t/�� N&)�؛G�2t�agC�1��ts�����{%��i��6�|�12|�QK@���_	�/G�L���,�=QK�U!/������.R~[Я�V;�$-��d��h�N���q�.�0o�B;9��|���7��Cy��OO��0��N}f4�����w�\��830�vn&�T�>A��pL�d���xiW���7�3w��0q/My0N�U�9I���G*�%X"�Nf��m�-�%{�`����oŮF�*(2�¸�;\�]oe"��c]B6�p��E{�����*�/w;�Ox	F�vާS��@��]-!q�d�&0�YU��e�H-u̻�<�p>W3F�'t�C���mZb1�޸�w�q�{$�`�YS�aYO9�9޽3���}�VȭnGƓgz!�j4[.�7-���J�%��I��GU���q�j���ڽ�N���Q��ʧ>񖖿R�Ê)�����7����0`�U6�_��&!il��m��ӎhC;�e�O�P���߳��/M'A��?}�})�	�5��E��=�\� �d�|a�au��l�;R�E.�8�g4�-��"�a�]�pF��5�h
�G"4K��-�b,D�ܱˎړґ��%�� ^�T�c�Gؼ)�T�  ����N�W���*�y#���ws7\���,����*���(~���-��g�/Gt���&>~�P5
`v5� �2�~��7��'
y�ф�,׌�U>��*�X<�f<�#�_]�^���6c�}/���fu4��}�I��z"Bg����ؖ���[+9�����IwUlxHĺ�#��ݸR�wn�O{�1�J$�~0�*�2�t_�LR�c �"�.�@����&%�icj{ �ש$��3گ�����ˎ��I3��~�z��J������F�IT��~xk�}�38ݟ��UM%u�_ܩ�ʤx�|XU��{B&�ۛp�ţE�)¤+�T�w���*�+�	����6�;�
	���q�+��@�@T��<� -��h���#m�ӔS&�S�]��n��è8z�}a��C�N��
��E��sԟr.��+�eA����ԍ�G  	����Ԓ �˔�oѲ�G5�+�$�&a�Y���V��J�.X	yې0U�Q��V�`��2�X-vk��D�*;e��5޺H���08��\�t7e�W�����fկ�f>F(�����lkq�3*�V�v��j��Ƒo��"΍��P%%�y����£a-�O�	)�+�:B��(�Dw���4^���5�ܚ�D��(}�I�0P��s
[�d�oo-��)D�;ӥ=R��f�M�^ܥ�8��Ӄ�Z�D��h�,��&��J�ֈ��|7��Z@ep�t77h�~Q�͜\�GG��?G�i�ߒ�?U��5Y8z��R����7�/�E\�C"�_�;)�W���G�5�	�Y�n�m9� ~��ˇ����̫��d�1<k�	/����`�^ܼ�Ԇ���|4�I6Y"�	�� �L[+�y����!a3/L��C��	�Δ�ޓ���F~2�H����k;
ȸ[=Q!qo���C��n/D`-�:�-���cq���V	�D��AJ̥��_&!�S��8h$��n1�7���L-������ʦ���6�͉01C�Z^J`F��K%i�ڧ=B�}`��w��]��{f8����$�	M��$#E���0R��E�ۜ�n���s^)sc4�Īk��>B�{hգ�b�`�3$9]� E`�n36�x���K�z�*4�
�:.v>B�%�~��42�'��o3߶��+����O'���'��(���)C1A9�1
%�؍�n^�;.: �Q21���1q���E�4��8�{x=��ݖ�W�*�}s�3L��"q�ccW�5���Q]5��g@)Y9�ׁi�5 J��>��Pt	}/TsL�ڇ&�v��O��5�`�+�G�;��_�������wBVqo������g����`����c�ַ�Q�?I�d�x� J���AF6u�N�h4�����ɧ�3��n���Afb�V����?Z{�^�	�P���r�n^�1��x�p���T���9���)g*D���	=��|�����b���F4gT���#Q����>���tWpj"����q+���$�>ӲS��厭�5K��	��pn�_55KO�9:���׮�غMJ�>�#�R,d\pJ3�	ٕTO(w�ҿ������h�8 ~�[�ճ)��d��g~"V�`!k���s�
��~�}��6�r1
7W�f��-/����Rh�ΆǴUO����4�����C�f/�X�t��gx�Z�F��@��:��ʄx60���	�\�v��}��\PL����W��OgjN�th����N�%_ih�Fj����(��� �w]�ON���D��5;$�$��W����8X�Ɲ����X��q
��z���z$��A������Ǐ$Y%���Gf���4�ts�1���L?$���$i��G��/�C�MR��z�ƞ8A���sr�)p{�x���ֻ}��%�aa���G���= �NY���r��Y��Ǖ8G��<���ǎ�Q%�bN:�I^�00Q��	�X:�s��!�#��X3✿A�]����\���)�+/�O-p�:e�o���#n^�޻�'��~���@��+����7����5�P,<7�pM4}G�_׺}">@�x��D��=6�-��~��.�'+�?�$�Q��r���}�Ф�t) �aW=a^̽�
Mҿ>��s;�c���XF�RFLK�F��5��˲�/�{O=��n=/�����m���{�sx�-j"V4aҌ�PC��EWu�|��#����n��4��Y�TM��}S�Pt��Г3���}���ۺu��@�i{wj�p�#n�-3����T������h��Z0]���&�]Kn���pA���a7n����o5��Uy�2�ô��`?�����K����F:{����@4��At�N?�-����4��\��>#�hѹ ]��P;Z �`��l/a�D#DP���=����l8�㽱n�98%.Ƴ�.��$XT���p���*��+�X�?��N ΁�� �_�H�$ �&�ҽ"�H���Rb��h>�p��J.���amY_�H�X�E�
��4��*{zr E?�����^ť��2T��x6(-=!��o����7hs��rڜ�Р�2\��H��:�Ë\�*g��	0�r35>q1'
$	k~�F(���9e���̐�P|�co��)��
7��ۓ�'��_��5z���������c	��]���w��Ոd���ձ@��(`�ߨ]�>��
QvC<����G8�>й @D��T�سj�6��X��ܟL׏0tȺ3��5��'u�\�a�� F����B.������a�t������5'��]�Q�]�it�58�͊M�D�q�ጃ\v���5��__,ÒĔ5��'�Q�΅�+l��Pl����H
�[c[/H�i×h�M��'�p\"H7�[[a�&�y���������ɠ�sآsc�M��Oy����i:���½�r���S�Ꮽ�𧉤���H��#t�yX���?/8<�k����߉�t<��a��p7� r쟶��������{�`�	���:Uk��x7�0��Y��+!k56�� �wp͈�xd���5���;=n��Oe�Z�v�]y�����-%f*���GvC������5kKP�;�g{��B���	b�Բ����e��3�6&�[r(�Ћ�=k�ώ�X>(��q;#�RR}�����ئ��Z����'^��?��6.�5�S'�"�2Z� �9�SΡ�-�&8e��O*�4�v)���C�ǰ"�!"Z'�И�W7.��/@!�ڕ&��bit���=#Ť��#a!ێr8��j&g\�����$�D�D�G�ˮ��%$2�X��ę�&�pK=�Uw,<�[<Ƥ/���X$\+�1���_�,|�������R!�Dx�pb�c�{hH���_,��Cu�|���e��g�A1�ބ�D���+ ;��72�jq�a�n�]�*�i?�B�#m]
�6�`8���ߏ&m|X�u����Sת��H+i�|��I�y
I��+{/��얊#}�!RA���O71D� ]���Ș� @��d�RLlU���e��-��w�UK<�TYGt:AM��]C	�z&F��i��>R_L2������j!ܶ�z���������U��~Ц�i����K;����K�\3P�ܡ��P��d	��qٗ��u���)�F��3ն� ���r�_���-L��lT���R���y߰9�cT��H�{PV�)�L�Sd�R�~ԃ��M�>��fj��/��Xg��n#��q��_~;��i�����5�3à�T;B����?���7�N�>yP����"U#�02�H3�6���si)�{tr�!�1���p�Ky�����̴��X��ִ��U�K��:=���a/�r��O�}�u�>���&�}s�[x�#Z��bB��8s}7�$`��[:��($��e����g��R�ߢ4����BT�ϋgz��k���4be9�F��ή�������C4B\���_�`��"�)z�*�p�����>�ǥ]ܲ�{f��y�o&�C C���	��G:�K^?P�>��3?�q�T6'ϧ)��p�����Vp�,f&&�GF��#���C���7%�L�t�R�-O�A�ۨ�$w:��L8H��@�|p@#cVd��B�j�!�5�J�=|��[���>�`���O�:@�[�d3�u�R�H�ȍ*��2�V���6z� l ��ز\NqS6a��ο3��e r8ʆ�ktT��w(��=�镈��ZCAߠ)�	}S�
_�t�	����3����P�*�/���6��,5��~Oz(¡[�����u
l#���������|;.R�����H�&I��&�|聅	���zQ�?y�[�B;3�bL�~ƳE��Q�&gB �&��?��
e~�6���m ����Z����g���N���m�3`M��J��Lu`��������ل�����������!�E��E�h�����q$Z,R#R?����v=�����P!L�*��\��荼�;&Bzk��_���oJT��ܯP�X�zpx��>�+2��5��Z����7�J�f��A#nJ���O���ݱ����]@6F��"�"3U��s�ӥ;J��3L����`!JxR2�x$�ĵ��vL�<���!3�/�L�������m&9�s���mñ'��:z:��6�&�dC�����m�d��m���3ʼtE�S�Qe[`��%�&��Oy�$�?�;��uM��Rϡ��$��E�Oe����`��i����`��qEݫ���ș�T��ȶ�l WQ�]�`�[�~tVtW��4F$�
�p	4�Fs�K[�S�Έ���nO�����B�W�Y�Ly�qƮ6�O�ZaV՝Qv���$�ȅ�*auhd�J����ҷ#|���5�������%o/����94##�+�G��F'��$^�����:��]g�����\B�w����da��|�3������3�YF��Z��U7RJ�q��Az�h���
�8X�,��`HǞRYV^�롊�h'R @cx�CE��i=�[�١���?t���W�����q�W�B{�|h�Ej�ȥ�/�ς=�Q��+0�^MҢ��zJ����t���RD��Sƃu{�/��*Y�u�V8���XQI<�<'a����?��. L7�V�������3Kdy��!v�>�=?Z�ؒ�EӞ.u������">ŉ\�{��ӈi�S/^�����u�]=��C��Ӗ9%�+��Sm���d_���^.KԲ����^��=m�1�8�BE�.���/��UyC�(�d]-m8�KY���i�ՕLC��u�!��D�D�����&�rl�q҇�)���6��2��a�������`�k�oL
������75c��;~xy_N���!:ձ�u�I�
ί����yE�������$�|�p
�t���%��Z�ʕ�c>�t�k9��'� ^%��W��:dF>���Ds�&�z��0��c�z�Z�K �AK��u�[6�r�$3&@ 73Oipx���a#����q�#���F�Ԏ�*��H�T��v;;�$����Cds<4emp�*���u�q��I����]�x�{��&^�Pjx�6�6��Mw�)6�������a�����V��q��R!.�� �,H��@K�s�a��s`gх�93^^jsm����I���&ՈU�f:��4�M�|g�5؊��䢯�wK�ࣵ��2k9OA��IdZc+�zb~}��nyl5O]W��C��oī��ɿ�w�;�S�<:��7G��Wh֫f�1K��� ��F(	��;,��۪��O���Tg^�NL#=Aԗ��=�+���橤	�!l_�>͙���� �T�hZD��P*�nܚ�t��݄+|5t,�w��|O~!�w����JS��du�UV)�����L����[������Sr*�s&�vp�λA�)#�y���2�:�O)D�t�$��b|q������&���L,�uݿ�P��	�&"J�E��7��5$�
�COЖ�J5�U��%��������&Y�+$�����6��G����8��^�9T�f�*�
,��g�d���C �'�������j�=�	�}9/�]�l*�0���My=��@�i����w�_�&B81"��	'�}i�X�v��c�l��"ӂ�-4JY�)��Ʉ�MoR���`�I��}B����~�!��H%�Ӝ�Lu�����J�=�H�Z)c�6��I6��:ضF6Y�,��q�I���^�qs4��{b����$0�I�Ԁ�wB숎��q��: Z� ��\~���/���>L���k���5��x���,%�{�Q_n0/�EJ����nF�#�<�p��H�nb��+G���� 'Ӕ�?ǲ��}851'Os�E6G.��3��n��F$����C/��q�N�ͦR��D]w� ���<EXv��!m��_��?�� \zw2���a����e��ف�35��D..���o�K�/�e�xh�-�9+蛓'^�)�3~�j��Q�gu=�uK}���.�q�2n0��j�����B�o��>'j�˧u1�u�	4}��)�#��&�=1g��C��揋A��z��8m�x;\U=u�c�G/�<;q�(T?���>�19���\��� ��8��oj8�!,ց,�>�I�z���B�W�s,��(�)v|�ğ�o�yp�2�RY�#�5J��
���e��kCa@Fpe�� y��=�O�mRt�2y�xpt�A��ǲ�ߝp��8��D2�TY˖�5-���jw�UNk��Vw?�*u��[��^�o�:G�R'h!�4}]��~d_�%��;�O�3.C��!����2D148N�5#�(]�c�������ڟGD��o!­��J��ˌ!���c��f�$H����N�
d����'�"����Ka�<�ǵw־~�_��-�q��	$�3ʙ���ݷ��i��e�l�O�,O��a��EuC��@*�ԩ]ŎA�!F��z�Lڰ%�ցL�6	���J�u{��[1IB8��C��g��0K��Orܙ"�I��9�MM.��;�:�}�&��|!p�&j;�1�/��� x�7�|H�P�m~L
���x�s*(�x A��Ɔ ��#���z<�����:����5�8�e��a��^�C��| �vx�l֗�����M�y;~ޕyu`m�s����W![�`�w;�7ndn�J�b��E��Q|سk�P<.C� ����W{��-ž5��*.:&�HXv�\�
e�-��+F���	����q�hɟ���he Qr�zۻY����(1���`B-K�諙��UЇ�1�K��H�w�(Bf���}<�R�18&���_�h�ŋ�*DF}�'�֞ۻZ�%t�l1[]� "9#-׺�G|�J��n���].'��w��3^�,HCg�[�|i��Z,%Gס���3&s��^d��k��� e�}.[�v��Q^[:P���S�Phn�f�$����O6
k��F�r�i�<��\F�(��8�o9S�9$��;+��d��=bd���<d!-X��ϗ3"
�v�m�4g'rq�8+W��k1ƨv+���6���R��+��&���Aҥ�Q%E��}|���z�Q�>�T���O�` ^Ar�g�	�lc_G�
��g��}ч	�
{h�X	�ry��Ҍ&s�∴ x"3�:�0�G�Ք6�v����� ��uv�������L���-%IsBv�!�_"Vn�$v6���.�iO[Ѣʝ��>7h�\
��A%��_�:�ݔV�c�q
���pf�,D���-�ɯsZz�&�)Ұ.�?��H�ԙM*0Pp�h�\ȣ��'ɨO8M׃s��$��&�D��Z�݃(ܴ��Ck�����6Y�,�$i���|#8�jL2�7� �ؒ���{5z�i-���>dW��فLdw��zK�`�8�،�>c����&���Iy��;Í�r��\��(A.���1�5U��������6\q��|����8��Y,���=�G0��h�s^���6�(l-	?�']BZ�?]���^�y����w/8ϓG;���9��A嗷`=F��[�>�#<�*#S�E��s�2'DT�$Hl�ʟ��JYɿӃzKC�}�����%��	-Joy-{�Oֻ6;.������&"���S0H�]��-����n�VmrcVK,G D6��ݢH�����s^����&+��(�s6�^�5H<N��~r�˴u��m~)�����[ik��ˈ�18�҇f�k��h��l��3�������뼬!�I�H�s`�y���� ����drH?��4Ō	6�;�X�`��C%NΑr�A����%:;P���]���{F-��fj��\)j�����X4ˌ�-�J�T��ݥ��p�`+:�����vL6#��#6��[!\9l�v/3&��ۻ��i��c�:l���F��#�=Ӂ�0��A�ou�9�W�,J����":PX���蕰[�}!��m�~�M^�����D�[�Cq{Ƚ@�0�_$�G�Q���}��$��.��qc�ٴͳ��ʲP�p�]�"σ�D����;��f+�����ڨ��V���㧺�=w���h��R�� �2Tg<绉���x���=��cy���2�mOC�M�KW��c�.~��GXm��7IH2=CĀ��E<K(�zM�j�ts��o��]\��H�8�>��)�d1M�cn�����X��xo*ΞV�6��x�������75���?�Sea}=F�3�`y��͜;%H����j$(}��}�;���2�}���,⊗�d�)�����OL�|R�Q:!�U\t�����9��L�dK^����p~�e�����~��KXB��� ����H��Z�v�3J tc;!�<�(��q&��3�|v2u�)X99�j�5�i�H�w�K�E3�A]I��:�Z=�ٸw���e	�v��ֹ����ܰ�ۦ?��Yo�v*ZlwT�7X[��Gx =r`I�I�X��j��b�+F?�3,��౺}�{o�@Pm;s9X����!��N�*Q��&~ʿ�W�5"������xx~&�R�Cw���z�9� �`�-���Ǘ_�X!���ٖ֋A�Y���~��M�R쾯���C{-|gS��_NO�x?�&���vf�`Ɣ5�M�[-����{��if�h<d��R��.�	8��5l@?=)�0~%��"�L�)� d�/69��΄L9���~��-8z'x�!ڵ8;�9�yMq���_�����gdq���!L��;������\�� ���3��d9������)�J@!
H�S��]~�y��܉[y8z9�wf�|dI�`�fX0��t�P���u���/���QX��E�Vz�qB�n=h�hS��*���SO�^h��c�B�t^�)����0�������#z�0���c�zz)g�C�%��{���"�i�∄�@c`���H{<+�َz�[v[֪e� �	�)��G�ɨ\nue������77�)(�&'���Ε���}��o�k����r�	���Opl=	�;-C��q[)�*;�*�p?w=��%�}a���Q�m�XbO���K���!C�6>}�g��^��h�#���k�v^�=�P|��7  �6���Šq���l�BSRNV9�)=o,�TM
9�Wy���l�U��6)�-�MM�t�cs`��Ⱥ�f��S5a*�b����bN�~;�\��1��հ[m7�w5ֵdl$���
5g)�RBGL T|�˶�C<)���.�:'}[Ƴ��.Q���ȟ�A��Io��!��g��A{W�0��F}e�1Z}���U+Ni��G�p�`gaEB,�!sT��L�RJAX#'��_t �7�z�C$0V�b������6�W��\�Nf���D��)�.|�1s�I�Zveʶ1��q�7WC�x�� �9p���J���
�E�Md���v��,`i�M霫��{���@"������Ygz׉at���1���B{P����!���;���ҿ���X��_����9�k����i,|wxl���h/�$Z
z��	~?'(j%�F��ʞ���̼��|��9*�8���
���O�aO���J��A$<)�.�Ǯ �N�pYp��X�>����ÛH�~X��jZ�0oU.��\����J���jH�-3=th	N�0����W���i�AM�賬���Z���:Ԥbp��B�fS�������=��l�~W8,l���,͕�W��"T��9I������2��~�i8v�2�m���l�^]�Y�4�,�N|�ToE5�'�Ì�NgM�G�$��{x?G`��7�4���$qFE#'������HO�+�R�4�;A��G^�M�VK|#�����6�l�g�쇙��n����8��ggT�H�����!�7��+`5�Q���T���$��qw���DK�����&�@��GĝgM|Ӯa#�%d��y���_�wo�]?,��{��Kߚe/<c�Sd��`�%���-V���#�:����^p�2�W�$�qf1�ʻ�uP0I�p$���Nv����D��.�d��;=��9���7\�Wu�*g�����<�^��c�:9�����k�a�|�>"ڞ�j�u�>N�"榵1w�N����TL��tx;Vk[�{���[ϼ}+��]Ј�ۥdHc��B�L��+t
���Ha�9�~}(�2��Z,L�o[��i�;��� &艘AYڹ3�ף�:�i]��+<��Hg1ߌ�r�1��A�S�-۫���g�X�|�K;�weљ�!����K&�H�6.ˀ�D�A�. ̹İ# ü���Dɱ
��21�;�e���W�KD1����b��	�@ޚ�t�̉/���'Q�g�_����O�C�.��4��$t�`ެ���&�|�d��!7���Û\WM�0U2�?x���2j�V|g^'z�����
e݇X*�FJcuê�c9��l���j~�Qe�	�,P������t����G�Aq�]�fm���.����0�7C�~����a 9��;+�j�V�?�  �>��h�;LKMt=����<vo�}��h
��:oRBG�|O��1H?w�KkQ�u�l�s�����}������#�S\���--��s���U�r�Hɹ��a��5.��a��0LK�C��debQuw`hL��tJ��~����x��_��@���_�n�N���WVq�3?
�ܱ�����W���s(��p̍r;ǜ붠��#:���ºx�4�����{��×��FLg��6��{;��c�4���2|?ǪOR;m-%8E�׳��YM\��MC��y22�֡�/�W�W 1|k��a}.Q�ng���F~�7�y����)f#9w|c�C���d�;>/&/rp�]���M��
�_�n�?{T>�=1=I� ��\t���W����nY>2%���6����;�����#Ǘ%����	���s���U)p4;
�#t��o�y�bBv�&��kG�;H�/��$wz��(��A�|�6�B� W���l�ڥ���#e��6i�z���1b<�IjW�������q��n ����4��ϸ�*'�T>}�֯�q�h��פh>U]�2��
�<>�^��b�g�������Bk_<g�mvvi�"�>l�� �������'IL�7�C��9��@.��Fd˲ͧ�e
$%b\�[����h,���p�&|�\1MNm����:��擷+y����|G�m��y��İ�F�T���� E��X{�_I�%�>6������޿(��VW���s����:ɉ�����Di~cH�{T!�<P/��m��LX?2��Y��4�M��~�♲x�oY�T�ز$�-�s\T(��o�0�Y��H�E۶�m.�ik�b#�&dqx��{gl6Jh��������>s�\�6��ՙ��,%F�n��s��r�����+{n�T�4��Ś�P�9�C}A���NHb����%����T�A���_��U=�S�'�h���z[i�d�;���^��S� �1�?���z�w�ԁ��K�,4��h�̃����W�"�r�/�BF1 0��h"��:B�	���#X%W��b�S���1�����;8�/��ȭ2�R������RJa�j��BHS��[�_e������ث��΅GT��ç6���E��B.?�D�)�I��ђ0n2���@Q�Fj�B|���Gm_|���G�}Z�/�k*��Nz����U��˂���}ys��j�5L���҃�y+_�Љ��h�)a�	1�r��5J�H_� �P٢�XNܞa��
�U�ސ��l�3�TYUA1h��!o#L6�	�j+>EC�����[):�� ��sN�>Vjp,o,؟�ҷB��7�BqR����kE�6�PQޭ��~+cy4�y��8ښ��&���0��.�����j�ƅV�+�,�� �!�w��8A谫Z-���)~�#�Z�� _���ݝ�m�#����sN��G[����+��l�v�AE~>�O�լpJ�@L`��}�-5�R�XB���A����z�#?q!��(��5���{�F��"�#T[(�4������u�8{��Q}]�`�8��>i�!%�.h�y;�㯟������bX��.�5���	OP�yKi�+��G�p��c�-�x�F�4d܇��W�ޭ�z�Ϭu��Pt'G牵�;�A��+̅�yfm�,�q�r+�O��.m�Q�ǧ�\�{\O����@3��@�9�
������CUHf�i
EY"�j 桀W5���}PQ���v��t�qo�W��XPm�}}O�7�d��t�C��-7��´TE��*w���%rJ��)����@�-&S[�ԇǕ��b���Mg�S��2 ����������������o��{ӱt+���<c����a9���+c����sKWEo�����d�-��ol �]��X'4��fE��=���]����r9�Y�h���3N�����8�~C�8��a*�J	���"���sO6VuY?��^���PԧI�'08��&��}�L!cu�s����.�O���#A����Z��
����dl��z��J�҄�6�Ee�`[�O-�~ ��5�󂭺��.ȱ:��!p���g�.擾�7l��e8�ыh����:d�\�:G�Th'��w&׼`�䊄�u6!�K����
y��|�'��
ww &���n#	�)y���:f����D���u�e���"�R>��̼��,P�JD7ER*k�a�ǈ̋���] ,�%B���o����X�kZ~(=sDD�Bn�b�+�&����ȱ�-��}k�p���8���S�i�s���@Т-���:���"�ǯO�x�
��pnH�������E��i�4폈6�{Eq�}�4a�2�X�VMTE�e�����NS+���z�%Up�J��H��|(�0NĠ��;��!��봻3\�-ܴ]J�Q�w�$�����]{�o8�PKq�����}�L�M�U��*~�C����4a}���S�pP��h[1�N��nM�i�c6��1˂(h�8w��%��ҒC�G}Ѫ���WU�� y)o��PP�r�_�J�i�ځ+����DV�V�g�6��A{�L�VR�â�q�>p���Ѕ���7$
=�ƛ����j��FD����>޹K���Ml�E�+�Lyd~q<�*�=Vn�$��]m2$� �+z� L�����t�z���`�BD���tN{)�y5���'8���
�����/M���d9��آ������s|�i��K|W�6o��4��R��Rǧ��{'�/��k4��p.��l8Hk"Vd��>#�������D��%�g�&@6\�3a��:!s�,���&ЫQں��X�l!z��)�o�C���??�B�S�*\Vo���Vb�I]ݹk��ilLKQ���Q�t�,�}�7O;�����W?�Kt���I�%�}�K�v5Xj���ٞf]-H�� y�R?;�Սk���|z�f�{$>Z-�K:����<��YL��1����}������-�|cyp����,G��@M
�]J�02��(,;��3�ɑ�)�.X����*a�Eq���-	/��垥�i@Aeg5�5���H91���UX�A2z��E͖�?H�������q��Xr���u�o�a�S`Z�X��]�B�4)�4�j�{��O��I�l�\>�����?_UY!s��Eb��k�?+��D$��R�k�j��<Rhz���-.HiWّ��q��"��p.'�:}�ިpYdd�b��妺�(�oS��0f<��r�[k�{��>����)�@���-����BA���8��K��K�^Ul_gÐjC��z�98=0�Tk� �l�1$������7��*�3aȉ�|v�̓�ø)��X/�/.���(wi��	~��8(�-�0y��)G������4����nd�36��
�ӑ�@������ԟ,�Q��@])��F�㈏ü�y�@��$��ﯾ*��s]������/J���2�hlgU"�c��i�g���ˍ�`�1�lXq7k�?�I��PK���S��~��R��-A��ՒK	$�#h�sZ��b��}p���Àܤ��;1�4�X#�!Ӟ:B�9��g�zXzi	��ǯ��Y�ʴ<2���0��Ɗ�T0�.�y��vjt�V��D�����m/j���%��k���=[��ڠs�2H�q|Ҹ(��9��u�`�ic~R���^O��):�h�$��iu���0}9��~v�ǻ�f"�^��w���-c&���Ȱ?�P���h�mi:8\:U���n�B��`��Qlqb�������႑��M����rXT�(�NɁ{͖H2�q��q>���?	V��X�Y���q�Z˃i� 9�����h^O���Q�]����E�0 ;O�ϛE�����# 0Cy����x܌,Γ-P�`�c��C%I��2dT��t>�≑DHid�D��݇��R^����MX��\�� p�{��e�	���و������P��V� ���	�hb�΃��Īi%O���m�b�,�1��	�� �B���qk ;HdSc��2����1��&�W��8�f�8��X��0o���1�Ux2�D�H�}���i,��\"���7��&�[$a+^s��$��tP�?7�i6h�*2��]� �S7t��r�ȹo4s�ò��pn�*t����g�?����Ai7�FI��bD ��,d��*�S�ݹ�J��e��*�s���MI��*�_I�r�z҄un��f�
\a���8��xJ���(���v6�R:)~fv%��gJ��PK!��~�#����|u�����]��Բ˒���Ɖ
qLʉoh��N�1�H��� �i�6������L��%it\/�F�ٔ���v�ˠ�e^Jh�����u��[/pT��y�S���}Ҷ:Љ�:l�F*��/	sZ�r�PD�Q^e�d �ςvÎ��\w�G�^���S5 ����C�� �KUN/�x,�S�$��
��B<R�*Fֽ��~�I�%���.`����30b�e���5�D���#\��epf�J�2d�E?p�vd�HzV_B���(/�r����o�˛���l �ن����
�﷽cW���q}'=]�7�G$ab�(=��A�s��x�p�۴�:��C�!{ߒ���Q������q�[��Ηs�� ɥ��nkN�#��[������!�<n"N>6!�>Y�gB�'��O��5�˳��T#?�һ�)t�����+���k����B���'&e��	Y�K�+�e�	��}#���	@��!�}k�����&��R��g����Z�	��@��(���"_/��J�{)O����qd�6~�����:3�*� GIY������'I���O�^�y��*�d���|�SNQ��{���~�L׸�I�2�p1;����������M����_��C�zpF���tKS><���/mm$r�tMho��L��X��1�g�U|��t����'��>�ҙh���U�CaE��ʴ�yɻ�,���I�leߝ�e�i��:Tso�>v��g�xe ��$�0�Н>Gdi����V�KH�R ��������=��������Iq��9����vH���W�n�IfG��?�4�'��mX��T�|J�whX�a��Gaf�h�Q!=�����h��(�^�s6N��x�̻����@�zH��W�&���LD"�M���T'��g����ڤÚ(����h)1��$=�����	-H���[ggr���7�t�&x��{}�����:|p��uB�W�@e:�K�Y-��;����6&��J��9�j�7�������l4k%���)Px8���a^�;%���y+��{��k{��0:Τ�$���c�Z� u��P�(�HN[!��TNP
dߌ�.����7����)��H�;M���k��^a6GQo)H��(�؄���p3)j�����u/�4���
Ʃ�
w�r/-��o	�U�|P��g�(���^	%�dg���$mc�كPZ-Q����=/����m
lɝ��yI�J�c��[��'/����Z�w��=���;��"���.5-}.7��
�"ݨ�����%�p����2r��u'���s���\�腙���H5�0$%)� �A*"�qtf�EfGj�>Γ��MK�MW٭*���� 5��3��C�pj��1���!7?���)<����V&L�^��
��ISc�:�3{�*\���sEr�V/yz�u2���26` O�+=N��Ӆc`�Y�}���T�	z'�^J�ۤ���i�!��ϷR����y��酲��p�R��lv�켛����^�\�S�H]���{���(K6������Z�I��B��D�Et�`;)R��S���	<�;�<��L:
��æ?�n̔��a���S`j���:���4�!�;���x�����6[1�O��%�D�| ��Ќf;�����u�����O�S4��)ۿ(���G�-쑎U5�(��Cd�=p{�t��J#W|�"Tl_�����t
Ut>��+oc�o�/�q�sY��i7�6P��yzW�:ڌ6�e�lOvy�|ZǬ���n��k����$b����'�Ce��N�_ӳ�"Q9� 'X�I�WQރ��Sh��Q��>�~S3�sپ��vC)8�c��%Q6]l���"��{.���4�t�-����v�*o�W?oO�%����X�IP�uU7�:��?��J<��^\.`�Lo����5�-���Hw��o���|2��^���#iA�,����A��.�Ĝ/P9�ܶ�M[o9D�ﮞ��@�'�#��%�+D0�+�U��?����+���
Y��-�Z�Ja}�=
�x�ǆ�KO�XV�L�	���!.�xw|v1n��S��*4s����N������Ro�Y����eHºX�V�t���<��b�Nz_�JG�7������L�q��lf_�Ϩٗ�(V�!��%�3��>�P!�=@���{��}Hۈ�)$=G�|f3ܖG��$�Ƭ�7Ӄ;�~_�����\,��� ���"r�'�@�6A�e!��>��O?>W���n��fU5�� ���d�f�5��
#��׃5��ˬ�s}+*��C�)�=���|x�\l�j9��3�^@ J׿���|\#�t��x=/�7@io�M��1���9��7���}nU����m�����b�-kӿ���� �j�w2����/�Mÿ��*����W�o]l:X��8�/l<�@J=аQF��|�7.�(J$�]w!7�.w/���N��x镨.-�0����.L�S�\Ң9����F�u�{�Ye�}��3���!���1���{6�FI���42^~n:���%�/�Y�����E<���;���(������N�"��g���G6��6m��Č�n薅Ȱ�V�K��|=xu����[�� p����q����bu���S巿پL�GEXR�����r��VAEu�2�����Vt��<B��~��h���R�������ڶ�\��1�C�s`���jG��Xe��y���D��<�,p�Ե>^��H��B�I@fFұ9���˛t�v[�mp;V}Э�a�V�\��9�84K �1��~���5
Y�!�^���=�h����0�H.�/f	Ujw伖���Zt��(�]b{�
��=/�8�N�΍=� ��ϟw7n�X�/nN��e�������B R��r�V?� �Ͻ�V\�1i�
3����a�y`TqU-W��>+�F�_��uq�$lƸ���|���9�����y('8�]�^��>M������v�I�u[��~{#��U�M"��ph�V�\#R� ���:����[�I���M�#����Q~#�XS�R~Z<�����R���1	G� �I0ظg�����M��x�ZVp���D�U����s���N�|�I��� ��=���R;�M����
!�Q�$v�)VP�����K56��!�e[�fA��ؾwt��b�j��=����[�����lM�6���k�yʼE�֢�;��g״a�2���0�\|<u��%_[:9�GB��;��F4�&~��U"%�5����eZ�5�2�%G����:�;��.�b:v���i}�%�i���$�{��wP��(��7+�,j������	���M�u}	��\���C�QA|n�"�+�0(}�	{،�N\u	��eh�R'R�<HB("nN��HMYQ����"��S>��~sj��b�K��b�Nl���}��:�a��b��LL1��g�����)�9�쓬��2(����"�VP���)i�&UU�J2'��N�T��ri�D nE�s�m�4eis礅aPũ��M�
�3��?��ZDe��N������9<��>��ʥc�c��Hq(|pd+.��fU,b`�@���̙S�ﻁ��SP�f� ~Ҿyo�<Who��Xwz�v��4���0P�����Wʡt�֓��$�8X��q3Dj��tu��>Ik���d���Sq���v��?zA�$�#ި�>��[M�Ap~�y �%g��[/��)���ѧ����fJR@�[7F�8/�y����X��&-�Y�����9��27�u�I�������`�tH���*O�� 5/*���V��穾�	Y�����;?����#S��KG�V�8���>��\���_�(8+"�槖�,;?$G^��V��~�tj�R�0�.<e�{��J/�9�&��A����/Ȃ5a�L;�*�{��D�_�뛑�N���F���X���\�����;K��b5'�}��t��|P�.��3f�� ���bL櫼��#B�y(n��_�^�(����I�n����۵��2��[�6M
T
jϒ���TI��H��<
]�d�kk�N0���0�S}Í[���p~gW���E����q�¶��E��|Y\,SL�j�ySgYr��jDcv��v>�l�8;�f����-�u�V�������%<=#B�6�/|=����a$���Mu�x�Y��*���r8����	#<��z���2��O�����k���|O��o֧�/�%T׉�y@E|�k\�K/�SP
e:����ez�wi�ŝ.'�+k�J���qOOB�@̝�t`v�*�B���#��5�᝙G�Ę�����l��4���QY�ܦ?0�˺�B���@���_}������4nb0Ώ�x�C_H�a�c;k'�a���*E����]S>�~��"�,U��%9MU𩒅�I޶"��c�V��� J�q=ֵ�5!�'�����j�|=ɬV,��K����+�~Ӈ�˄"}ˊj�w)��yR��ۋ��{���uy�Ad���o[Sm��-<ħ	��1ܝ��A9�����d��ih�G�YH)g�u��6hu6ƍ2��$k�q{�Aa,�j��I��d)����)K�!������j?�>/Z̽=StN��o ��fy��dz8��QEO<�)�c���']�VcLԏ�{�0�l�P�$�O>�x)��:��F �!N�}���ο�W*�M԰��`��8Z�T8���e���}k���e��ܛ�n��!*.�<Y�B,At@z�@(o��D���������ŀ2����+F�	�Uc�J������F�J�z�}��#����D��I4�	}��@�5*���X�TQ*�RX��mgV<���#��@Elňpm��_�P�a-f�"�Gi��yuS8�y9���#;�|���P�/���7.�*cV�ve�
���R$s$2��Az���*�}ˈ�h��Vb�*���L<����_�re��� �R��t����o�%��8za>;�Eg��fߑ��{L^���C�� �P�� n�@vn[���C	�զ�[���Ѱ�B�0�#�*d;���b���u�:���F�p;�0���м��V4T���f5�T_P[�nM��#�|+��1�]a�Y�t�QX�����W�f�A	�g���{R�|�#/h^�,�������/�"�Dk������;�F92j����o�YÛe5�A��/t��L6���Z`&d��?�y���aH�կ~y��BD���'���oǥ�'����E� ��wƛ��CZ����c��#Y9@�! �����)�;�M5gO]�B�h/�6���SjSm�e��C�;UϨ��OE4��a�~^M
	�u�>b�M๘t��	b���f1���J8=I��e���{-5�i�+Y��Ћ(�l�wI�u��VI�ےԃL��4h r���~
�8��_U�E��*�!t�j"m��Mp֜����;?R`b���'�W��l�?A%ȞWC��;e`?��W,�1?׊�Ֆ�~ڸ۟�
�|B
�8�ot�|���J��5�j�mY� zEjVR��,����r�L�&J�OL��-tu��S$/�D���97�R����ɴ�Yb�_��P�W�_��\)B� ƖŌJ���W�A��e�k�G,��y��] _D�ϙ�-� w�
�^K�����L�K��X��#��²���_V ���.�:O�����"����%��^4�O�T�_/a�ey��C�N[W���`�7Qq��C$fs.���z\���f؃�A�.]q�N�Qg8�5�3�o��B�?8'|{/��07�+�}4�x�<�p���`7&ˀB��	~�v���D���#�\l���0��o�pjz@�DtD���)5���u�dݴ��$�O4��\&�I�����]��y̬����f@��]�<��F@���=K�q�F��X��Qw���y���h���Vtv ����bD���?,=�*3Bv
��VX�0�lG�=�����dJ�y�K^ �n�z�X�a�ax؏7��}<_ؒe"?����Œ_��r	V��#�[�S<b͇�z�(�S��1m|V�5*��F+؃	�ʃ6��5���3 �K??
L�睢�%o҅_���6�����>ÑswfB�E�\�W~@�K�	:��g��܇���&��-gM'�b(�'$�\ae�4% �0�A!��p��S�Θ8?�nW�胨�3��y���Ħ�y}�.A�#U;V�s=c���s�b���D��h}3���3�O�Q��.����eQ��[0�ઠŲ�
P�&\@@�mS��_�A ���j=�Zӥޕ������_���o��f��J���U�&`ق���/����*����c5�>�-
8,�7z�g��I��z1�	 ���o��*�cֹ�Y��������-
݀0����M��+q�^�zA�fS=dh�ծF�z>5��^�f�����L-kDh�r� :���66Q�|g��Y���\��3��I��f<7$��b�U��b?�C���\Z��C���� NI�;���{�'ٻ���,/�3L1N9��Ak�ՠl�$�.p������">�+�h�2��-�m�b��	�;�����粧�6\z�3路��]���p��$�4������0f =��,�4G ���^��hZ���%��!�M���9=W�6lST����T��S����bݕ~���Abn��G����=��*Q�������Z$� F`��)���GO۷JM��Z��waS�����Y��(�51(6��}s�V�)��p���
_��K��F��'��|S�ҋ�@3
����������Q��H�{�xzq�C�
�A�g�F!�C���i���l��z-�.�b8:��}���Ф\�JС*M���,{g�tDwѵ
:�rm��3�/�;>f����5�Oa~g����}}��DoV��<.4��	�����o�����E��C���2�JUki�6�ݚ�X$هq�}���v�jT����v)�5��䭭P�L<�&��rF�B�iz�:$rkX4�������Ã)���v��:���̱����+ �?]J���Ԓ�1�����K�J��<F�ڃ�]�'�z�M�Q�K)Te��F�怆Jw���w`'M}����ط\y��+�	��s��O�@���ɜ��;x���`��>��=Z�)U�`���ܾ��W�[���L���̝5���
���c�l�M+��t��܈M1�*����V-�1K7�Gb�^m�F������PZ�w��h�4�a񐒰Y�_�h)�A3;�<��a�G}�r��竸qT���+A"f�x�����TF�|x^l�,GbO���Nҷ����*w�L�fr.��p��Q)+��K+a��u��ޖ9dqG�+��$g�#L�'��(��P��!u�%l<�B����ޓV���A?ƥ��s?�5��oUPG-��a�M��I�c9;,˧hMY^�Hc]qr��2"�-QJW�/Ҋϓp2}����_N:����4��q�o��C��������q�F�zfi$�g�S����R3��2;��9����^ 5�rD<B�c�,��'��3��$����=>(ŵ����l\k��O�
ӑ�g���;�#��%@N�:j^]_�R�y��d,3�$���'i�)�5Q=�lo������M�h&�>b	F�U��E�g�S��|˙�;g�V
�t�t�Y�/`�'�O�����3֝F��M]�h��Ί�@��jK|�
�lRcV=VcQ�dj4�Ӌ������[�JN�Z�tpC�Fx��Ӹ9j�F>�w�B�+D+x�@��jG��&ݎ���`$�;G�.7�ꑥ��_n8��1&	�@��ӑ<��4V� �c��0c���%�4 9��L��%��t���	��c{h�0zj�be�ӑ�ҽ��"�1�%	�ܵ4���P�z��������2���ʡ�*�Ѽظ����¢^j�2X��~��AI��)TϨ� KKT���0�Hic6���@���'�:�����v
i����A��8`92ȉE� w������F��i��T��o�<T��(~]�k�!AQ��������c쬔�PWW�n��"������?�!��B��r�r����C�j������uʂ�1i�e�/��ܵ��(E��Y����sq�ڔ�H�3�x]M���0�GwU�|��;�%#ԘB�6x�W����W+.�&�'�$��T��)$vVy��0��_K���A���QJO�S)����ؘ�L�67Q���TX�)Z�!mxR��o�*�^�<�](^r����7gZ�4�L41 ,�W>���X?� �|�� {����L����ؤ�
�>D�E L�_����_�!�tZ�k���0���kܝ�X:��P����1���ij��+Jh������������0��)�o�-������brW�bY���(x:�J��-q�p�# �.�=���;Ӯ��f�@����ڔ�����~3U�*@&�� ���杨D�����/�d�H[�N��$٧eq=�%e�|CDW$�kE��w�LBR�����E%��oۦ�Ch����3��`�;	u�UOʹ�Q��hm>k_�d������J��A*=Cf�|�t�/�Å�}ܼ�w�ͣb��ڙ6��vk��������!=�ݩ?i��a�� ��e�`�%�!��@XJ���T�,A����*���Ɣ�f��\�*�!��� Z3�")n/��m���HNjy|����))S��t�w^��8�Ls�Q��Ec �Q�$��-��~\h�D�9$�0S�f��N�x����Q��XU�����Y��&z��+�
HBNc
[~�`$���B��C��!f�A�-i8�>�y�
����5�6��dS�B�!)��A��$sqև�1��	��Z�8�a�OPz��q�,"�vہ�Hs;�
u��q�S]O���
Y�2���̀�tZ���W�F���D�N$��T���$B��?_��`b����`hZ	0�?����_���Ib�m�/Nkf;j�H��KS�x),-KxM P�Ѓ��Jͥ�\)�e˰�����a��ft�;�k����4��K�8˓���*V �����M9wdf��``���i�K۵H������sȤ�b�~��y6N1<��w!;�g惑�"/}��n2F���V�~˲�i�=����xRĝ�G�6�hU����P�v�>���[�7U&�U)$���7���	mKq���Oڇ�(1���Vm?,��g��~���1���<����⇛��EP[w�� �,���d�k@T�gV?����ӝ���l;Ny����ud�� �,H*�^�˦XKQ붅��R8�)�H����H�������fMo�V��������͂.�e�������.��~���[����*���&���oG �~�t&U��-@�t�ka'�&�#k���+Ow���q�k?0d�d��v�Ȋi�� '�]��/��.'r�p/c��Z�������0F��:ĵ���؆����dc�,��;l�P��Ɍ�v��"�X�+EC�'Vs' Ϗ]�;ª!`pC�ܗ
&$� \m,<3�
6��qo��GU|�d���;L�A-!\f�m?���be��|�D��1)"�V��W%A�W��o��BJ�2�>�'Y����?l�Q��X��ah��d6f�Fv�#C�	́�H�*��I��hTA����I�m�0H������(��V������_��Ծ��`�<p��ZeS#�{/�=���.��(7'��ĭ���ɕ��vs�)�^��d���Lt��++��	�jq�#��r�ޛ'��>u�x羬�v�/�3���YDNO`�"���۽n�J��vIZ.���a�:ئHQЋ~J��O �4�~�	ޞ�c�*�$�T�i�d>J���J��GU�@+s��Y��h<`��h�.�b�(ȰJ\��@��1�m�{dc2����UO?����B;�x�E���N�����XK4����D1�i�Z���W��H��T@%,7��*�p6�:�3S�>E�
o��k�ph�R����x̡<��~B�w��=�����e��c�kT��lah�+1+�ؾ��p<��$1Tj;��c��W�A%�ք
P7�����qm���"��: � �{���{(���a`�G^>Y�;�Y�`���}�1����`��7���� �����!�Y����Z{�s+�ԓ"��vY�1���F)��
�<�x%mMӤIO�Q���DL���c�����q4ڕ���F�6a�*�����b��7��R���� �≹?��n@�VW�N���8�˼��V�D�wC�$ɽ�ą$��\�VH�5�C�%�B�_����0cV�o� QO8n��; *��T�=_0��?���x����Z<'�S��G{ԞΘ�qq{��� dα�6e��~2M�!s/�:�����$�՜h:�)^�8��ʇ}jR���%[e6m��Y�����Ɉ�,��\�k�VV��c����h1Ԏ�0���JD��S;ہt����4+��i.���瞙��xX�[� B[����=?I�8o��'W�ΟZ��LM�~Ic�g��~/M��d�g.�jv㻐��}�c�%V��Q�������Q(�$�S��ZqO9�c�"�<Q%���rQ{��$\bږ�8�����x�$?a���ؚM�K�^WFEJ�ݪ�7#?$����j�5Z	�@��p�H� -a�z���m�=Z�$!����y<�pZ�'mGC��x{���Ӵy��L+���(�ᕹ���ǳ�SU*w�r�u��HR�;�A��`�+�͍�.�$��&��w��v���D��E�L��˶4B���c;�aQ���" ����'᫄&uțO�5��"f���WZ7"������8E�&��੦��LS仁6�!��!:��cMf&���4��.w��X1~ze���kq����T�o����E���xF,3I��Bm<^�"A'}b�%LCڿV2�~�;����M�n6onh�8��8e�����'y�ͥ�#�P����́���+��h&l����AX�&�F��-��ߧ�D���}⟓�p����č��υ�^�Y��yˁ��]�^?��Jv~����01D��pwS��Gɜ��@�t���W2TH�3�ffz���As�)�-I1��$A� �������WiV�r�����e9�(C�W'c [lイ�J����|DOF���g���U�/�6($V�=V���'�����l�/[g��I�x!ܕ�֗��}�&Q��*��>�ϱ]�<j6,��!7��$�A!]��JF�f"ٝ��0s��ฃ@�Vz��|+�]�]���$��B0���c�}%q�x��g�EA{��G�*\zi�����t0IV�����!��_Ӱ���\� h����Tgb���w��F��^��ux��\��"�N�gY�&���O���G���F*���j@C�$�ml�j#�FmOi����ɹ��Z���k��~m*�{�?K����T+(1�/���G*��^�ϭ%��o (ߙM��F�����^��ў���,P~��߁F�y�WW8��Ō��!@ԩ�0�ʱ�#�܃��Jq�A^:��V��WTߌ�;��粧�̭�eJ9I��k���눉?:��H�k����m�UH�pPG�����?r{\r�p�ȸ8��L�~��Nf/�7�K��Io5#ɱ�����qܩAh����� &.ݵ���i�B-�t�(}�W��קQ��O@��o_<��V\e����~��=�W��d�g��폟�n��ȵM����52m����\.�V��2���=�����/n�3*�lIg����ŵ]������/T���+��,�/�	5C���B��lS��غ����@�g݂p�o�`n������X�h�؀�k���V1l7b ?\[m����R��b���H́K]��$��6ph�vno�$�A���-6�{�Q��A
1�}���|>�[����e�>J^y�i�QU�B�m;�ꊺ�"��X���4���g�,="{Os�/+�jG�딵�b�x�$��n��rw��B0��#�*������qz��A�O޶*�t�n�J�:9�ݹ%�Z)��U/�á�!F�՘���`��gX�Zt��AC�5A��G��,.�}��Zm�P����'ޠ���;J4;z�&�ƤY`���h��ݓ����6��gu x�	���Z�@D�؀F�N�~�xj�=�Q3�]s�K��u��.��
?�Dc5���M.Z�N���d���2$!��Q�. �wP',Yh�b�Nd+1�hj���ڡw��x��_��R��.k���F�uL΍��ZE���)F���' ��q��4��X��~Ly�ܑ086���w�8�u���OB1C��uoC�6T�k$l�<����y��jzD��؂��O�ڳ�[?��ec��?�NL��,����dlW~���Y6��ˆP���?��=pSE�
[B��D��^���4�k��Iv*���}���؜�#$�o�]�>նqV����<J���?� �����H����8����-��~G1�� 50N<�� ��=7�)���f��(�( z���A��
��Ҿ��zw/Rz�LI↘I�.7�U�6?�S��q���u�G��2�T��>��X��, c�ЂX�� O,%E�I&�fJ-_8�$ ��U��=Dk��F�����������-n�&X`��׾c��i�?��Z7��/��x"��H��l�7�A��M럆SI�-2�� � q�B1�-C>��8����ZQ)��EEO!��I�9��+��_���ٓ�e�
*Gx#�${��h�B�q����#\�I�d�hT��t�v%�u��hJ0�j�O^�����k��h�ّ�|}�8�KO(�ӵNC��._��y�#�'�����r���3�Mg�Kb Ð��I�	Ń�C_�q�/g��c�g�_А95)��4j�}+��.����w��D79��~���?0p�'�ޯ�����{L�<����Q3 C+�w9� ���m;P�^�F�֦�.c�ߍ�d�0�V�� �(���'��{đ��i0�{q��m�)��J�Ϝ)IpZ��&Γ���e���M�VX6�X���1�HX�"
�Gr��]�\�I��@���_ċ��j����C"W����S�26}8s\�-~lckp��ZtR��P_�н���;��Eef=�5��e�b�H=f�h�*+�q1�C��!6�6GrT$L�NM�<���Hi��|�B&&0��%���D���~�@�iB����:��l0֡3�����C���VI �G���<y���k3�?�1%�K��mnRs[`�M������k9���C;�J3� �+{�:���`k-��|��ЧJ�q�'��\{B�p�y�i�9m\h��|i�;��j�Xn��F0���q%��sy�3(��o_�,ȡw7܅���¾�t���<����L�0R�z�'�ZL~����yP�*>�ø;��ڀwW��	�hlɼ��J ��~�����Ũ
YUL�Ed��A@G[*�3�2��!ς�2�&�������4$>�|oJ`GR?�+�dcw����B�x�H乨�
L�A'H7��Cm�S9��40�>N�׃��7c�ʥ�ȏ�̔���.�x��rd�a��	͔�$�)�*�e���ON�Nul�������������@�it5Uov�y��)��W(�{�����䪥 
�,0�q�Ew3}N�?	<��g�gk�q|�ٰ}�??#q��Hc�&[��1
R��u�� F�y0���^
���~Ȼ�����)Oj��HU��p���M��/w��uY�� ����Vd(̅�|ԝHV˰����{b���9��@���N)G0�,��k\*�t�{7?f/F&�YC&6�_<9� n遉�no7�:"e�OK�v�Ȅ�֎HY(k���dN�� >ĂYҸ�nq�k�'�0H�Ϲ|���F1���ίDWM�Fl;(A�,�{�;�Cr͌G��L�,�RL��'�0��l?�;!�6vix�/�n�m��s<Lz�Y>8�\�p�S���( KBa��ƅ!d
�Cs���>
N?��SgV�]��+�������P��]�(w�mh	6�K̩D�<z��ҧ)�je�MD@��ڟ��U�u����o,^a���W�1�F/�NU��S�2G�n�R�=���D%�ƆHH�^n��;�ڂ�#pc�T�{���5	�]j�8���\8�7��]eE�ɠ�X D�%ml߮�}F�|�Ͽћ��pތ|So7(� "KG�a���%#C���'���ϩ�0�ɭx0�X{[����=|e,eө�
�,�BqC^Y��S�O�vg��f�����a
"�{h���-ѽ�GP�oN��Ĭ�Bͻ`����:%5�Yj�Eʗ[ݳwq>k򻶴�9���ƒ~�^����о^;4����xh�_�F��[�p ���6lW;�olh/!K#�b�	�<ԩ��K�*��H�mx��
xA|��#�p�aq�\��Y��>����`��� m�.�v�"��[v�d�.� ���@c��_j�ŘE �x���#r��v@�>�Pc%�G��Y���Y I=>೚�Y'���6N��h
��^ܰC�F(�Bq��OZƺ
.��=;������S�A��!cR�L�e�J~(C�E��1I�-?��0<|w����"�$Cr��M~����a�Ѭ/>웉O���ZaWC�p^�ٹ��A��D�_�:�ܣ������O
���F'�#C�����o��g.&�0aϟ����
� �>@|��XIk�їW��'P�tH8O�$q&!FB� \��0�@L�0ן�t�4$�(��덉�RV�/�e-.����P�!���q>�ɓq�v�"kv�07Qy��ZS�0�R~ja�։�.�H �t�����&L�I��r����A5��慦8ѽ�,n��0#���u��Ԛ}r/������[3�i���cʫS����&'�4<ei��aM�>�e�k(�Ҳ�-b���z;GF����"
N�:J�kO��pO��K���7��Yl2+Yލ�	�"7��@n;UN�.��nm,/tp~����j^<!yx����6�Xn}#�i��Մo�<�K=�UWc���4�]��i��䜐9BěmZ��%��S����ǚ�AxӐ��z�O��x���<7�:�
�$��8oj�*MW�S����������t$!��}�^�rP��`����h$�����  Ң)�]����(�Q�]�V5��F7������p�/	c���TĞ�~���z\�u�qH1�Z�V`�[	{�6��+5�9��p�sv��[���0�'�ґd�B�$� #̍ҩG%l�5� x���]��N�Lj"�!��ZQK d�Z1!��qN{�dg����tR2}��"J�P͐�%������5��Ŭ��?)��q��}f-�0��n�ʀ�N(����f�>��E�j��i�:7�D�.�O�oE��(ք�u=�\��ߝ�D�?�ߕ=�?�Z̶@�5ɞ�"�W�����*󏝨j�O�%���P��(^���+�d�F�9f�{Vy��B���ں��c��hD,.L��C�ݹҧ0�#2�^2�vо�j���JŕT�џf�ݿ=/(:ɐ5�Op��`��Ϸ���v��#p�Dav��a٥�P�X1��B��c.������dah �w���Oc����na7�j[�Ą�]���TB��9J��*6w<$���͓��nS�/������dU�â���S؞�� ����0/��%t���}��wS3��)�aYr=O�TD�|Y9�8{�a�nW���!��8���pShN��z���D���h����:�K� ���?�V�j��*e��x9mi�Y��%L�^ЙI��W�@�KJ�,�/i��o%�ia�e@��|�%e"�+���`�
j���K��	��q�~����������
{"
�(!v�ȪI���^5A���y���LY.�*������+�Qobi����D�&s���h?0��a�-p�텧#�(���L�Q��]�38�9�gŗ6��K���a͡�~���C~�]�Gu�2��?@c�*	�r�Ϳ��mUq=/Ď�D>��3Z\@���G�|���r�'ïhߛC�n���@�A]8�/����-].�D���h(W������,�<���}M�%0��yj���K)Q �.�
?N��p���aZs��2����訄�܈F-X��\n1��Oq;p��!S��/�����=��,ji������+�4�#�of"Ó5�:����S��p{�b��ʚ���x�ڤ����P �߿�i���8[X��`�Ռ�2�?������B���c�Ew�ШZ��vsO���a�n#ę$����JvZh���1p@J�R�,Ꜧ�%6#`��F��y��4�!�`�o��[���2�Xe�Y���	DqW>W����l��A���`���l(�6K��?12�W�Ô�PJ���<��N�ՔQ���;Em
Tk�����w�Tz-�v��<+$���Cm��@�dC��h*^o��#�?�~���k�F��Kۣ�l>�[���	�J�}��i����v��XsQ�c���W����EPL�?ٓ��|)
\����k�c�wA}s��nR�nWQKI��3�%�K��Q
�`pe�s�؜5��y����LN 9YQBDj)��V��OďZ�|����W�V�����BR�_��D֕�D?0Կ׶(����ac|ԃ�[�V�_a��1�ip�"�]`d��]�gG%�t�!g:��hN��J9ǁn̹40w���DS��:��ka%Z��/�o�R6&e0Tl�A�;�)>�Cx�Kt��*g�#Fx�s#�8ؗg_��2���R��B��#�s��iؿ�n�z�u��������>x����dn̌�3����D�oa"�>f�<��-r~���Y(���*�/�d{1��Oa�����N�C��l=a{b���J}�nr@��J��>6�� ��HАԁ���Z��YQK]x�
Ak��k�o{
H���o44n���6���I�(AT��m�&3{&��ڤԹ���n�W�X�"u���u���ƺ�]����X�w|VŢUH�X��;B�,���of�x*�cy��AR�ڕy7�x��b�%�;E��~HpUx��ՉF�lp��_p!�jӢ�d;���Ƴ�0��~F��rXnp�?����am����ӊ� ��i�,�V:���R���V�	�7�ٱ7���.ʺ!���*�"t��������W�������Y9��"Y�}�Pw���gw��TR�v�Q�;ka�4�ݼMeՐe�� �9�,+��W)`x� -�\��KC蚙���U�@S��n��5����}�F�O�M
��6�PR��������"u]<�C�Ե$��2U��U����݄�����/O��e�����\�B�G��=�����* ܰ��Γ���m��#B�U�x�lD��j�8��7��g	��M�k���Ֆj�^���ǃ��c�oP�#�n'�6`�0�9��(d�_���;���67�״�g�!b&�*kp1 �;���"!�p�\�U!�C4�<Eu�:���c��:���B�+��:��.���؉��C:7(�,���31yx��;)�Wg�7.$��Q������O�H;َG��q���b���3�1�F푇܌�b��}��O]T~T�!,�<`n��� ���OYz�U���3>%u���V$�Γ��ƉJC2����GoâX�@�ƃߕ�~]?�AA���,-?��1�=�[�J[uQ��G�+�¾�����,�Z?^J�%'���WE[�܇��v�+!qΪLD�.�-�wi�xQ�"�\i�(뀗��d���-���`���yy<y���6�_�Wf��\r�e���ل�)��b��uIY��ܽ)�;x�
�|���أd���rpM�l{v�\���ռ�2�b��=>)T��b��
f�C"�utf�Ο��'qg�z_ָ#[R�IZ	�0F)�X�P����N��O�-|ww0�83��L+zb�+���$�9B��'L&y�}?���^5�c�,�o/;���FzY`jb�u��5y��`R���T���]��a�*�2�����޽��^��� Ė�wOp�*�٩��\�9�S�������h����V�B�1��5&"f�z��;���v_��J��H�ԗ[(s�o��MV�h9�]� N#_�-/$q���j�i����7�v�]�2K��9���j	�Ł&�Җ�Է�G��ix@!�-=�y
T`���;<5�.�}����6�T�1�����̅4�_^"!#�}4���b�_I���L��ǵ�S����%[ rܥ�}F�i�F��OJ���Dɹ��.���"���O}zY]���kI�3�vY�9t��o3��^7Z&_JQ��-h�Pg),,�Ȅ�s�m.*
)[;~dAy8��w6�� ûZ�2�`��p"�t2J�n������qS���;^�76jQy"����^�TXu��㒩�T��>�ie�2Y��b�A�O�����QZ랓�덋c���O���(��8���n�.	���'?Wf��tRF��G��t�����B*�Ɋ�f�Πe�2�ϳ\q���ң��Ք:��e���O>&���污W�ꥂ�O�W�v���
�<]�E� l�1�+���SJՉ�\+�cx����or��n���� I�.�*��o�i�MjU���"��~�i^�@�H_gGNb4�{�+��g�����o�c�r��[�&3{p���!��t��TIs�� ��i�M4�/�����&m�Y׿U)�ܖ�a�~z���?�I�n%
b�~.IO�Y$��uW����rM��+`$�����;��m�׉>
����]��#q��,*e�������}�C�"��հu6 ��8OC�nf�Y��Êb,������W����Z'(��=	����0���R�8[J�|P�l���^�U`3CU��"oo�k�. � :��2��ࢃ� *џ�&�s� ����J���K�o�c�M�r�ZV�#Dڶ����$�7��!?Q�Q�P�K6���n����Jq\�u	�P��TȺQes�>a��%�@h��ڙ����
t��6m���9�6ej�l0���ss�X$?Y�h�an��Ϊ�A�e�c�	���h1���������dr��>�f/Nɐ��Go��U�?H����<����RW��`��+c������׳�Z�"�6B����u����{��@F�;�V1hs~:*���h�����D�;�
�0t���p�D._�B�F0���S�"�m�{��1��M �ְ��\�j�nK��׼���cp�ۜ��:���n�V�{�9�vű�XL",��V�l��Ǖ���v�h��)��T�Ч'�����Y���껁oB��p���*׼�k�1>��^�I�h��^kї�sA�Y�`���萂5����X*�g�!7���s�0�(��*��Z~��� ���h'�	���g�wG@��W>��G�WQc��DI35=�C�y�ٵ7�����,�ހZe6���l�?�h͞�B��l)�k��*�84�#ðwWˈ'�rEjQ�G����z:�0��I�0��)���t|iq���黠7�<7�2?ֿs��rq�����8-Xe��F�S���Տ+;V�q��7!��`��/`�v�d�<��/:-��w%��x�|�e�5���(�Mc��帎>$l�Fdy!�lJ�(��v�Ӏo��N"�9i��Q�[s�rضC�P�����z�wyƕ,e������᷸�'ip���	�E���k����,��D��ڧ'%���Z<�
�����������	�ZM<D�=߻5�D�e�9ޡ�έ�&�pr�?;KS�!�D!��~8H�1qS�"��7�)l��e�����CB�-QC4�T���n�����H�?;�=�`x��3����A�y�Ĺ���e
 o5'�7#߻S�f�)	�&�l]|�aB�]���H<�Q	�<�!��,�/��YH�
+����X�ݡ>1��/�P�9�>���^~�̡[F�t|����wx��pO�FjR���1B��m^�1�oρY��K���8>^^��)�Nq_<��L�4��?�'1�|�ɂ5p�W�)'@e�+�|��uT)/DCz"QiC��\pEl��Rn��	�w�WF#,�g�H'o�*�V��'��HL�����p�[5�O�mH[�UF��~�@��.{k�N7¾��8q�O�W~ۃ$�H����6��k�901'J�< ������ٍ�C�/gz����#{���OqNn����$���<1�f�`�cv7<$����L
�)R����sӴ6�95I��1��0��i�!��;lq42�z��r{D�<C,#u�1\0�J Q���?��G.�,P�@&=���o���iC�b�)�qn�?.�h�zrb���C��|�UH0������;���yll��Z�s�"�F �a~f��j�Xk���ta��Vk�Y�)���A}
[JEz��E�i�39�ն ��CCD8H����Bx��|0'�`Xg��Yj&U�yND���&t'���.�`����	ӠL�ô��kޏ�̐�\�@�;o���J�;f��=f����j[.���e�bOÂ�j#м�=��D4�5?�ڳ�U�Z��ܮi��t*S>�rݬ��`��1�ˊ3�rm��:^���9a� w��$�3�% _ȕ��U%�� �W,8#���Y�FCi�-D\�+d�v�f��f䂬��P�F�yY�aԄ�FYM���_^���]��Y����3��FA�XS'���B��ĹM�K�ڏ:��W��6�܀W��r�0�Ai�&M�z�?��R�)ƹ��Y�Ⴊ��C��(�:�q��5]
Sثc|� ]�p�4�6���m��b�Q������ט�jr��\\@�$�\���.IL��I!�nY�uM��%���9js���Y���@
�^?¢ �0B��B��Ѐ	SD�L��GӮ,�f�U�������Z������w������D�T�?��l�>�nΐZ��d�zW�H
C�l���ZW/�1���!��ȶS�JML(G��`���� �=�o�ͼho����:q��%���L��~,�������O1ū2���d?A��}rNM�f<�|����_��/7O��z�:�0E<:�e�	�Hf����o��
K)�z���L��-q�
"����C]N�I/�+�<���C�_�<8[!��?��'��՜�����c��H�o7NwdC,Ҿ�9ж���� ����E������꾧7�R������YuiY�;�K 4a���6��?��*x3)|���}�bt�ܶ�9Z����U����sVJD�mawn��q�WE{��c�9�(�m?�{2��};�'�/d|�e�c�e��:QB".�,��8��[D�.J�D���o��6:�#��e�����x���0c'����U0{�Ʈ��*�#��nѻё�a�WZ	D=0���C�6�7�j�q|�ߙK�u��Q���Y�51����x$Ec�_R���){��ġr�[���5�nޥ����v1�1���|_JL�+t�Dv/���Оhs��|�a��,)�h�7��F5�X���m�͊_����
Q	�:�9w�5Is���jJ�x���FO>��K�2�cWd���	Z@��甑zSEt���|ԗ���|���@������5f���JW�ḑ��o�<�������UrY*�񌮑 ����ܤ$���S�ѥzUo��V� ��N�~?V��/Q9uG���ˠ%����z�Ϙ��C�{����d��5XS���4�uf�ռ8�e.���iK~�a���!��+u�߲Ȓ,#���O!;��[�A`7APa?�`1�W0CՎ;�#��~8�&���+��Qv�6��^_�Im�����g�Q�?2b��2�3�#�
��K��z�������(�jǨ�ms�#��{����id��وқ�<R�^�tԞ�1��E��ҧW���	"B��R���qjo) {9�:��T�r��W^WkZ<F2u<TjR����I�4#��Y5���ʍ�ۤ�(����ݾRkP#Y!������V�My�>��F��7sSm0�AgC����1'"���G�y/��ԴTuU�|��P.��;58����+�{Xp�\��%4N�Bi�㚔�_;�KefM#h��3@�٧�C����� �s����֓ ��]~�TG��n'Fr�b�q��4��:��aC:�%�Ay�~4t�W����m�ֹ���P�������0��|cRd%zV��)j/�Ȏ2��ߏʞ>Ӷ����'G�x�3�!-�`��* E= ̒8�>l�ﭼ;bA4�6���ʹ�-=R&�W3OF���H<fgFFx�
J��7=�N9����R۔� m�����([ [F�m�ԏ�2��qI���X��aegͅYo�
��"h��[5�d��,7o�s73���[G�H��ȧ�,�S��_s�D�"F�s5�Q[Q����B�.�ٮ|���e�IUSu�+\� &��8cNw_/d�_� ����~�~�W�:�0p���D�uc���	�j�2*�0�is�n<�,�S},ÿ�n+��+N$ZE�E[�5w�f1�R��<����F1�c�{�����JS�!�j_ȏ��NS.d`�V0D3��oBu%�Ui�(�-��h��ԇ DJ�W���V��F��e��Һ��8�B��&0��s���n��XUY2� �ףýnm�6˯�z��f���7���VR��� p����������P?�����&>�o�D6�.$6�
*\wh3�ĺ�TU�z�w�a��0�Y�"h�i��Ŕ-�/.H�ž7Ұ�Q������(��*^�$�]�0��a��1g2�'�������?�e@���P����l���R�	0S� �ھf����"U-�s���d���)$ʌ��3Z�Ш��?k��v��
�U�Jt���VNR3��/�9�QIׂ����fӟ����Ȗ�Ô-5���c}W�2�Bhl�7����Ӝ��=>AC�$eA���E]}]I���i�۸�U
j�I!�����������M�7�!�xZ^Ψ��%b��n����ER�U\�ؑ�$���n�)95�9�()����9{>��V��X����#h_W�n�g]Ǫe<��o&�Qă�'��ӟ�4�ba��%�f������g.\��0=T;R%�(�0�Z�?��s3��t!Ck�j��<Ͳ+m�$��,S<��d\���g��M��^��}A�=>?��yۓ�N&�#�����c�@1Cg�����%�`��y4@.m�-`���׌�D�R4���@��Ox�7J���'��}an���/�)�� ��`~L�L�H t�\��e�՟�:>k?{g��AP�>�8�TF�A�L���4M�/�%z�P�bĄЩy`�wY����O�o�f�F=�bбV\��¤��Q���4kCT(�?�>⼴���0�SM��O&�p4�F��^�
��jJ�U	�3Z��
m
'���ۚf��l�:�/�^+�a�ه�{�cc�Q�������}}���=�m
�W=��D�&�Z�b]� jZ�K�k�"<E*���J�'�㖊�J��� -��>��z�׈;[��o�3}��+��։��0)aa��T�;�qގ_��J���+�|Z��I�\�~�?@M2+����Uj�>�;t`"��LG }L��l��T��6w֨?k��X���ힾ6'@��]��7�o�"nm�����К��o9�pv$r�yŶ
�c�Y@h�:a��s�e��,m[p-��5����{K����\ع��O?!Ɓ�>VX�.�d�W�������f��]&q`�a2���R:���H@�*�<�;���*�50����`��tIy^(�oz-?��N���?�Ol���M#�F�"���")�¶�NT���ʓɊ2cQc.^��O�Y���>A�VD��K~�MV_�8��B�U1�kuO�s��ʣ��r�X��q&�:{,Ѯ\~Y���w�:1��j��*jX�^D���VW>�Y~�T�۶�r.G�h%� W�la��X�fl^��lG�d�<c�a���r"�8�������d�����0&����ۦUk*�n�:�h&��8��6a�3�M��OT�{Pː*���( B!{����`�|:���æ&	��L0��H����.�����u����>c�ed���Y��y0���sM���Ρ��x�A١h�zԬþ�F\�l�N�,�^�@O�;:��1���}D��'�d����18�N-0��j\8<��i�|��v��"�$P�j�BX	Ĭ+T�I:�3��6��\-���м��Np�ͅi>xO�l!���Qo]m��TwKB��JJiK�a����in> |�׶sQ�V�!S2b�s"��a\�+�u�O�D����B�1���460x��4%��g�TѺ������J�4�WD��I�e���~�G9q���CE��`+a���MH𠱞3"�-g���-��`���g��H��3ǽ�] ����l����<��o���KHax(�@�x2���ӯ4?h�p��$�4H���Y��=|�f{e;��<\���om}�Vf����U����1�+v-�0��芤�"��A�����V�s��{�j��*�;~b�j��w�:a����X��;�n��5���<��tg-�rkzR1�-�g���5�Ev'����	�".��A[%��d�F�.b�	����sA��C�BIt�>l��6�Y���O�Т����x��Ћl��p�1߇R��Ieϧ�h8%�a����y�v�g��l��O�5��S���a�;�6���Ӗ�-�r�/�
i?�\����vp�9����}ڐ�1m:�� @d苢 �ߌOg���Y�z�������XL7]���88���K�_^E�s�R�)!�H=�-�ϑ>�x���#@�7.�L�i�gK��ݕ���g,z�ƌ��QU�n;��.`��Y?�B�����t��M?�� ��ײ_��=�A��h�u���T���9�KW�Z@����?6��<��_X��԰�c�P^���c�Q^�%u��_m׆n�2�
{Un�A���S8����h�1|vx�{GV���C�
���ZbDiS�1򥞞d�/%��oA�QZ��Ș!�G�i��`�M|���r�Y(\1��U�(��8)�ȭ$�ƛ5d�TD�lZ=�&�zĞ� O�����'e�ؙBB��v��%�#ۘ�:c�C����%W0��x������B�P69�m����(�%q�u�V�2N�f�Z����	�o�'�eO�Uh�x}�
çe�/~���Ot�G�؛���E9w�I/�ߴ�7�f7?+W]���/Ĝ���A_��jnU1E/��X^���tNF���	�ټV�o����p	<�ɝL���H���ww (�;`���ڧ��}�x��[��n����ܨ��!����R@9W�pA��q/�%[34�0�u@�$��WP�}�A!����_a뱔��
Ah`'QC��i}�lU��D�!5�c�ȘO��?����UX�p�%֜9Y��&��j����+�k@a�6����������1�Fţ���c��O��0*��V�܂�:�A�T���'.�	n|"�.Y=P9�*��^��Z�2<��v���+kō���4C�!�
�V:�ك����_I��F�9�ve�kn;*��&��7���=2�=`[�4>�����ЪZA����ʽ�M�'c�1�j��_NBaQ��y��`1� &�8���f^7�S�;�>
��Y�J�	]
�Dp��;�S�,#�����Jbp��K�t�\������yV��@+c�Ə` �Z���ͭdUb/���C�S����T<��s��z;k�U�rzC4r%�X��T#FF�W�{�d�p��Kh,��R?�~�fK�w�cGDl3��h&ϙuz�pFZ8�dJ.}�z(�)
D���-BC�dV'u&��}���aY���`�ʪڟ[��("��XRK^+����	��pv�p-�+�ې���){|4�$���QGT�U��o�-/����sv��J] 9��v$>� �?�J��Au������i����'��R�T���m� c���n8��"ҳ�`8����*s��e����'����F�^�N���AB`��Ð����𕉴���S�� n8ik��8�X��s.RQ�����_�U��pBM߷�]��j�!
����/B ���
���r���7��r����Aks׾D���#[�����Y� �o1(�����A�h��0]��N��t"��zj���:	R�M�m��i����U�1�� K�r��.V��Dc����<�R�V?)�2�^)���1!D3�%}
 �:~���eq�@E�wΤ��s)��Vy4���rv�b%��������������b��Io~}Z3��D��/�7�^�ދ�MHG`�7�~�V��h@`ߧB՚��(��M��}Ui��6nl��]����mݴ�J�Sd�|a#�x�������OD�pA�T�F�o�����A��^2�C����9����^�M`����Gr�$=���x9�$}��D��Ƚ�� 톲����l�c�W�6�`�7�BЋ��V����hm��7V|������^ܒ \��\���ru&�8�K��a�)kq��2����Ʋ��vj���������,��mb����?Y��s-ұ��{"�z�p�9/*9��g�4�d&(����)�@��]�#�(h_���(V�s���_�kfn~%��~4�����r�d���гT��J�I���n4��q��:��N���B>���#�+�9
<c8�s)��B��F[6J�*n���i+ ���m�j��Q�O�*�~�be�$hs��"4��#NلR��B��#j��g\75�<�|Q�վ�+.�R�&�+���ip��l��ļ/�u�q�r���0���A�]5o �C�~�䁞;�5W����%�ݯ3�����?�i�ȀkD�dDc������X�T��ZVZ,B�1n^�woG;��)'J
��o�m����\s�ތ ��9EЧ��O�?�cZ�GI�X.��Ҡ�" �P�˾��g�ܑ�x޴�}[&,�$Y-]�R�Ȭx�q9:���r�M ��y��7�Qڎ�t�K��T��i?��iU���X!��`�t���alw�3N���*춭;&5)���A�F^*��Zc�a4ݑ�5;�[�KK8�ϩ��ZP���a��ݫ��`�q��ӭIY*��2�j�<�0W���v�</������$&q���H?i_'�+�z\`?�|��S���U��w@��AT(��6�V8\�|���9�Ǯ�c������J��o	��80����u%�0�6�&�B;[�ld.�`t����$�"�R}���.B�@UH�����N'��&����D�-��Jlm:�wS���~���qn��Bbkـ$`���x�}��'��w?�}�����p���'�����+�(v4�6��A���~��|� �%�|7GM��\
Ǡv����_͹���?j� |��ɖڒs;kv0jh��S���k=�
5d�Y&��L������N�e+�*)M�0���1����|�2�3>3���q	��6��2�d��-Cغ�g�K�)�CV3�P��}b������:�"�7z�KD����I&]�2�|W�W6�XKߎ\�\���dZ�Ɣ�J���??��~f�R}q�&��˔��nq�;Z�_K��0C��G���[=n��q,�Ӝ�AX)�+Z=��f�4���2q[1��
�o(�3��Bٓ��(��yCC�>���LC!��
�����*ǹ:�6K��`G�_�t�=�����R3�Ձ��K�������
*�� c�|"k���)���|K�;ܙ��t����5#�֡���'G(O~����(Rģ���&�t���X��q��p��r3���C�:�Lfp�[�6ص�.Pl�OʐW��#�B��7շ(��@h���S#�V][PWo����N�D����F�?;�#L��_��f�����E6w�t�FA�S�rp�R>G��Ƹ\h-��(���3�&��ek�h�"(&���ߎ>W�H�0����M>�}ݞ3'%_]�t8�iǪ`�h�������������]̙|m�ן�5�t�{���Cl21�)�[¸U���a`������G���IK��϶�q���Ψ"��v7���`+�E�TZ�"�6�Ӯ\��v��"+���\�4D�:�
�{�'�5���D�oߐ� N�`�h��c$&�ո�_K3�4���A����G����E�:���_� "RH2.�_~M��;�U��� {��;��$�GU�d���<�X�עR�R��i�%W�����.��g�4��f,�%���m�-���&v�]u=N^N��X�]̽Ҫ��#g)È���-�ǳb�Դ�X��=E>��1����6$[��� ��TT�t�`S�.��u ^���O.@Z��a�8H�G\7�v|��2��!�����`/Tv��m�m��P�9@O����򠻸�&��Pe����ى/�����2z-|u[9�Y)>@�q8��C�-Z���[*��Gyi�XB߬�:���Ob�I�������������1W���t�����|r���b����Un|��6��+.C�*��h��]���4 �D�?Ʉ�H���(�p����c���DA b�+�8�c.��XfOZ �pL����Y%p��w9������a�B��<U�S4"���*�S� *a�C�K�^����`����G[}����jK��r��ܘMnv[�x�������S��N�/.K�1l��eM��x��憁�� S�Ipݏ�^��V��T�+g|�[X�W��+���WB��x�04��]Y��&!��=�w�x�6���	$4��O��Z�dCOE/�̞o����� ���1����i��^��
�.&�#����.㍛��K�>>$�a�ٍ��^�<F��3���֗ƥ^C'��b��~�ӟkc\�T����^��m ��b������^�*6_�˨D{��9��R޻�EW7Ot7���p�����Ɣ���D�r(�#/b`�66dJaez��r�� M�,��w�6�gY?�'��ߚ�w/����Z�k�ΐ�BM��Cc�- ����S�Ϙً����B�N����z
HXx��ͺ(:�-� G�H��ۑ�2r�q���� �|(W�[�$�j��,_y���{�k�_�g�h\�?���� ��;��*�e���������B����G��L��{����xZ4/m�6�n�����7Qǎ���
����g��b�ʼ�17�M�C�II0|��ؔp���<s�]���`]���K�/����{���4z��{�(�H��vri2�[�PX�@�"�dtօ�Иm	rT�7o���U}yB?wU�o[Ify���_��������^�u��g�7��AcWa"r���s�%:��ق���/vq���K9�ۧ}���������Gѿ�1s���ws�Bq�'^�N�����X�6 8\΋�*v�;�6�6��-jB�5%V�Rټ����Mfϲ+g�Y_'(dc��S��]�0.��b<�� u'1��<8N��'Y����c�z\	j��ƚ�nI(�Ȏ���hy1�V1��F(尊�F)��a���P�(��U�֝����~��l:����]=ʈ�ܿM_3VL}��ɝ����<
� n��Eڳ���		�:�Y��&F(���A�%U����.����T2~q�o�_�騄��z'��,3�:p�k ��HL��0
��W\���9�zՏȨ`v$��#i'�B����R��=���/�Xl��%/�W����b�	���r�iy�D;�;Ɔ�I9�=Rv����U�IT���"��h��J������tI��x�3��ˈ�ޗ^�jdTD�@%�����и#B;�t���g���	�p|�>�A����E�dn�N�z�ӈSl��������5\i�A���~���۶�Z�f8d��� ~�~��n䚛��Of8��fx�p��T,�V��D�b� �b����!�ԼdI뚞'E���S:\�`
��;�����k�fM�O�U�"���#uv�������%�=����+�04�t�Ƣ��&���E��՝�¹q1{&D�I���DB�ZUw�gM�M����rS.��O�Z��ߖ޴�$=%��8�#�~�u�B+O��󤳬�*���-��1%3�|��tU�c`�P;��|�JK,a_�0~�V�˔X�ЙxM}������U�zm���FQ{r87��/y��}��q-'e���Ց��Tt��7���ać�Z�b;'�f�ď��έe�m��n��@n�cp�Zt����D~�]|���2Lh����g	�ճL����@h�	��4~�#P~d��E�L��L�"�n�9�x\,b� ;��Mp^�;=�x�k������e��s�yd=N��
h�E����Ŷ�_7���<Q� ��7�G���B!�N�c)򒶂c�yKm��A˪�.+�f�R�_��4��G�)6�؉�q��
p��d��w
��g1���ƅ6�)�ډv�Ud�T��o�J!�L��ػ@���W�O�Ǳw����ǒ ��2�������!%�S�W�7�uX�AT_�m6J��@��`�o�DA�p*cߪ��n|0�v~{���=kȬ��N��T�daMSi��D��E�eo��MԴ�x�z�D,�2޾kz�Q�g��$-��G��m=U���;�D���p:�%��a����z���W��o��������"�6��;�:K��3B���n��?�\�5oh�S�_���y�V� b~��5�¤���M����N�v͇��ˤ�ή�L{�݌~^���w%���~�u����ԕ��莹�˞�$��ش3֪m@�-FL�D\�z�L�6�K��\�����֢,q4c�Q����ua;�E%���_�_D��;�;���C�M�*K�~p�pm=ǷYMK���N��nՆ��5,մ�� kg/N~�_�!����<�X�6A=c�t�\t�]�d$Q^$5��q��*�O�����,�'U�.ȥD�f�[X4�W����jǫT{�����^���A��ס�)](�h֓#~��z[{�K�Rt̢I}WW�)L><������� �X5ޗP�u�k�J���*pr���I��$��
�X���fP1�� �@%1���=r�~�x��i�8&�eD��C���ъ��v���Z�X8\F�һA��u4�T>��!���|Y
\Ω1�Z��ۡ��tW�6=϶��֫��yL��F�K��3]�w�N�r��]��-{TWF�EF���.
�뎏i��#J7����'�M�ˢP��ifc�$CS�dj��Ű����S�[)d�e+ү��S��l��~T�s!�!"2=ą ,q5z���\.ya{E�57W��XhH���	�qnyςͷ����#u+���#�F ���YS1R9ޤՎ��T؜���1w:kwR��pq>�)5��,�d�#�b�GW�����v���kk]��ѡ)ia#���d�2�0fd���`l�m$�=R��C�f�a�v���ؑl4@�gP��+�"J�����Jj���L�ɔ��e���� }-~��	��@� I���m��0D7����S��V�0a�`3_�.�����-�NI��GA0�Z	E�}�s�ބ����(@׽�A�yOaJ��`7M��b'{���l�k��QGkHVV��4���E$t��7a^���{�xn�!�
�"��� En��� �f�-eV�{���`�P^�6ъ��]@M�.v��.w�-�AeK���?�VmHJ����v�r>��vx� �s,mF>�2U�*��,]`Ot|��͂����a���sM�.a^��{,ۼ1�Jrk~�}�f� �����t$��¸���8z@�Ș��5V���ں�����pN�u���b�V�����N�\����i:�q[�<k�NQ0�!��	O��>
w��&3m�M|H6=#�o0�UN��U_XW_��~F�okX��������Ȕn� ��dx��W#�;ĕ�5��@iރrY#ʼzS�m֜�d� �>���E�c�)(�q�ռ��'qp��#��(k�g��J-�/��9��jx�$���k�	Nz���[�wCK��"��8nu,�֙���+�����aP7�.E�m����b7���i�n:r%�jJ:誜[� �,W8(�2!{�S�\̨U��m>�Æ��t��� ^��ʶ�Z�6��.��}���n��4���#��zHQw< ���?m]���F�S>v���[���z�����ġ&"ꅆת�ãUv㝹�)4V��i�����v���G�����m@�b(�;��"z�}�9:%�g�=&hg|u�m0o[V� -4�a�c�h6�ӵ���f�׈�&Y�lMc�kKe}��\G�*T��st=�o��w�^i �#��+Q��R�-��ԕ�2)C��T��vu/j1�ɋ[��a��'P�c�N�&Fs��E��~d��˪I���G=�E��f{�(�$��J4��i6��A��k����u�V!=�����|����~�$����Z����
�~W1&gXL�_��O�yR��:���#EP��I�R�a�0����0*�`̠�o;i�i8�'mO�r��
�?ީ�\׵=�
2\ڼ$_l]�yF5�O���*�&��Ŗ����\���_��{'�����5TVjVz�d�^󋒝a:�Z"��;�s?Ows$�Jh�(�JFWj����7���D'q`y䔋«��\96����#�v��>�����q?LI�	x
ɟɆe'��&���Z^�D,b��M:�}�Z��1�ү���?3:)n.�JY`��q@�Ny�dk#����wIѥ2a�i �I�O����ؾI��o�g���e6�="�@#��y�_��Gf�h�8��А
��P����礈��8
���~)�@��#(Ǵ7&��FIo��һs;[��*�
���}j5�kS�nϑhP���ae#tQT��_�����Ke<˵	�ɨ�W�ʉýlV���c�|�}sq�l� ��j��u��)�`�pB�w_r����h'�f�A3�������4*J�8�,�~���pYtV���ɸ�qO�� ������v�!�s�i�dӂ��ɸ�z���ѫ�C!����R>�DԳ<�J�Zڐ�箸N��Ѷ.(X�=�΃����\�2rn�L�hʰ�T<.=?%l��Ma�(��[�:�G!PB1 Z'Ay��Vq�}���WJl��-��1���Q.'�C&�A��i(ip��
1�=!;����.hy�-�k���)�$`��̗gj�
��ƝfOr��O�>82�ixB�gwN���oB��� ���+���d��Y	��洫�u���C�V��޲�����﹨Z���\k����i��9�\Ms�����ɓ=����@��r8qr�}fl� �[��ȥ�+'�V�֕����vhߞ~�����
�w<m `�}?��;4�\��S�%���QW�4��*�P<lR�����ל�_�;x�G�y�8P0 ��]��fy$��El:��òP9����"E��ؙ���V�5G���v�"��,����F!�ty�,��q� �/^�M����[�ZL�s�����t� �Y%�*��A�a^3�m2���b�V�M,��[5L^��G�l���&�R4mj��R�0�F.3Ɍ	1�!>������VUJEV@�(D`?��R�7�{l6j�v�{ �I�Wl"g$.��'{-|W���@� ������ī˃좒�i�O����(]�Z�"TwS�꿸GW�|���2�r�\+q}E�����=M�@�1���g�A�@�e������3�ɵ�FF,5'Rfzz����o�H����lr�T�s����ɖtٱgI�88�B�r��R\j����:,�3�xn#<�c�bI�n �����
�=#�z���s��}1�R������M��P 흚�ڌ���"g�VJ�z��䋨4PG��9���@�U ���z���S�H>��-�����x�A@Gz$�8=�yj�\y���2��S4������
 )�Vt���r\98�uB��u�}]�V���̥����;h\Gpou������Y4�+�+���,n
�tO$��6�g#Θ��7 ZcS~��T�9�n�\�l�SQ�-JխIϵ��U�QR~�jb��=Ź�u�o�9�I��οe3̄��晟�TY��1ˆ��@[_�	�H:Ԁ���0T��&" ?:�J�ɪ�:H����@4�`(�5��:�aȂBw�@�(s?����}���(KD�a�zq w�8��ᝅ>�@�Gށ�V���U��{g]%B�ss-��/���b��޴<S*.��S��qԦ���h��&��T>��?�V{E�Z�_g�����|1�vb��:�d�6�'9�Q
�/�cB�_��f��/��V����ԺV%��t5��_<��~Yt{�]	��X�����"��
s�#�S�����:�"�]�+h���q��`��N�lf[�"&�"%��]�k-�g��f�X�a�g꿳ќ�� 1���,Nd�ۓT��������{4Ω��.+SR���n�2C�OAW��� �h�yM'��\�n�E�X�ۺ���7(Zn-�����L�xS��Wa�89�cm��ئd�S��0r����;f����[��ƕ[��_	qc���r]h���JP�c��W��T/���}Vk�D�ј�����TNCD�_�y�����3����m�M�x���X���ƀh��i�_d�m�'��P2,��5l	)�Џ����Yh�#���oE�(�>�ՏS �RXI�\�q!`���&�!���؃�x�@P���7��ףUVM�3�|���������+c~�h"��o��o�����5><8c�k��M�De����s�ND�q�f��"��@~�Gq�L;6�t@�fH�O��dXu�
�X[j�@B~��]��ė�-�LG[K_��J�G�jf~�&�W���Scb�O������t�+�{1�Ha �p��Y	��q"��:�\:3���(��(�N�Bs�SQ�ή�9���_���d�A�d��������W���5�Ʋ9_��2L��=/E��������82�M��X�0ś�2��X�?����@�����^�u_|0ͺH�����K�A���V�,x�F�����^�P�� ���]W|��2��*��C��zC��}ן3��ȗ��㛩G�>K���;+�U,��]0,�ߙFX�� L�x�Z��?���H���q6Q�  �-?<��K����,�^�4�s�&����&`q��}�1�$���'�Ϡ[��2M��!��_5��h��*�VϛOI�xN���S��,�@u�X�%~j`s���LR�RO�iH�����n���vv� ������mʣ�u�	I�ab�L� ���9�&=���7GC1/J��l����ί�eq�i�,�v.m`w[KM�3;2�&u���^����(!0x�ȥ+�x4շY��'"�׬��_@�Uɇ�K�q ����;n�H%�0�a׳�uleO��Z��
Ci�#��m�I-
����
i,0�Xpf�$���Ĭ@�WU4[�t���[�����,,������a��u8# B��ʁ�,퐵-��O�A�mT�����(�m�t*�TPX�nAFcC���eO�E7	w]:����]^�8��ʴoDI�`5�Ϯ�t���I��=��Q*c=�2�t]* \�궳�2k��y|~��"A��1n�����fós�N�hj!n���5���I�]c��΢��/P~N����2G�حbt�B`.����$&�\5K��Ƕ���8�vr�6]�������n,���2%XF����]�:�	K�fRaJ�&�U|	Ie#�"�>���pvO!l�������+l��Ն�P�*հ�-O�����@������T7/����3��j1��E��F���*�F�]����'�6_�ps%/N�YP�7��G�p1�~��
�+��N�N�y�Ș�@gjP�.�"�͐��͋�����dS���U�=�^�u��g��Zn�'~r��VBX�B��)\�������][zi����tLno��ת�������*��ZQ���͜*��Ɵ����Ȱ{c���<�ŵV��N���T����!��W����
c��&(A�|)s��E���rvI�G��m#�	3�j����=Wf~��F.\[Y���N����wS��@z].m[#T>3�e=� ��`���/ۥ��Z��XP�jM$�Q��P�z)���d)AU{UgP�_)}M�h�1�Q ������ݽ��Qt�B�dZVy��T��v��-9�S��d�Uo�vI8�����G��o"�_>� ��j@z�:��JKTgC*�6~�{h�nq�
���þ����4���U���<�COpg��&Z��nD˥�Y=�z|��T�.�u��E}�UY;�9�������4绉��4��h<�ҏz�u������t�D`	��~�Q7m&��9���.v���RD�-1���k<�����Z�� *M˦�K����L����	����N�2*��(�!d��kv������������Y���ݻ�(d���y[��R�h���{�_t=r.��19XН2<;���S���%�����䭸�� ��ڛ�ᗃob�M������R�� �T��{�m�zT�[w|1��Ym��J��n^�����w�^�fȵ�=�#j�I��|�%[��l�Rƥ+m٣�Z���o��b�mi���N�P�ڌޛ��>hpZ%WK� ᑫ0���<�>l���K,Ż2f����5�R�K���(Fbj�׬s�v��ۍJ�`� �@NL>��M�R癔l`U����IgII!����N�4�{����#���#�Z�zDه0Da@�%�ܵ�����y뎁�\]�$8O���G�i�A��a:KK�ģa��D�p�LT������^5�~F(����W��h�(�iɯ��y��4��E�lY��q�B�t��}�b�2���E>�y!���F9s�����U���f�7��LL��Ru��'�s��N���ɮ�2�g;/�Z�X��r�ı�1sj��e�oE�z�q%���,��_a O��c?�ٓV$.#9��tA��A)5Er.�GlQ�����*�O�� 뷻>-\>�@�F�w���GX�ǣo�zΰ1���k!�����(PAQ��?k�L�{Q�����D���Z���o�>z��jT���LW^�<�����vԇŲ��d��=���aNA>��E��+pP��P*?�,�wYp�D`j%r���b��χ\���g�669��RQ�ƛ�[�OW�ՂV�u�\|N��F�}���&�K�I�w�]f���;�V��k:��W�lphҥ������s����y+�n�����v؟�]_UEd{��ȃO����a���۬�Kf��Lͣ�O��!�"���	^��@[O�A���!H�KG8�۷�Ժ�p4x�pD+2�͠Xa�ܚ��X�ܺ�z�#�P�.Ј�Yo!v�<�����s[��̹AR�?;Y�y?���RnRa�.}3.I۫�+O%�pP':M��/s>�bӵ8E'/;�*��̃���ˁ�R�v�.�1"�7\^�/Jqxr���>s������&i���H!��7N>���0�"���q�b���I��vE���a=f��]5��Ye��X�������[�;��(�ގVBH\6��g���\�	j�#v�����}'����5�,'q��m��{Q�sp@g���A��J��w����k̭��&w�s�(��掩"�^|�ܳOٶ�!�x�"��qkb�đ��k�������u,���D�\Ξ>y����x,���{�=�n���W�w�q��E;m7w� H���%�%�.������<tF�yiYj��w~�8����94��.e'�v���)�)>��� }��(6�Ҵ?��%O�~��{��j���ܞ]];�M�	�r�`(�+�gT�y�_S�Q�U%�0B�􏒼ѿ�J�oh�=5/eU~U$��E�bW�����H�^�z2�2�e��K1IyAO�� ������!�5���m;u�����b��@���R[����O����u
1��3g�e�^�1D ��T�����^EX}�A��zh.7"��,��B�K@�ȿC�K,�7����;�����bJ�
�C(�f��	#�W��ER&�VFudP`��=oI�;�"^��ǔ0Bx�r2�ց�����GR�?�n+��XLk��,,L����W������E���䀹�D�a�=�F���ѥ^�T�w�>��������'W�{��C�*���4�8H��a%6�r�M��
0�ЁP|��^��@��|�ͮ��@ً�V
��70���5��SXzD�S���O���dU��-�^q�ό���j���V��1K�H����,���&̅mt\�N`�>L5O�2���b��G�V8gG0k�@�\��y�Yhlݼ͢�b��������I�!*��<��j�
�5�g1�r�"�N�L�e�IXK'�-*:в䨻~iOS̳0�sT;�7ty	�w��]~����ڒ3d������y-f�v�ӈR��'ŢM�/��]�i��z.gS��&�Г�h��z]��ZӾ#M�"�[_���z9��mЂ�`�8֩H_�]����m('��wX��_����ZAH�G��7+>v�/�H�F�m�5��!Xwz7���1f�77����Ѹk�����>�|ߞE�W`� %}0_�r֦���p,1X�$�� >��|��Q�E�B��EzC[���.d@٦��h9*�U��8�����w����{�V��
�3���_��s�/���h��\�<+���	+^��X�xȖ눇1ִ`�.a-0�'HE3�.�by1,I0���aaM��_���6�e<�)z}B���o�,�)a.�������;��������B��3����oy�z"g:
"bn���[$jǶ\�M�6S��)qM��=Ã$���B�N}׾]��\��c�=ٗIV���	Di״O��&髠�xܦ=�LN����i�^_�r��b��!9E��
˹Sf�J��ޣ���@���>�@�
��aFѰ���;r�{X���Q�un:b��nu�`	缐̗��v"�����䊦�o,6��aV�{�u*�w�b�o|i�>��v|BA1c�TO���f�u�y�Fc��iqJДW�?����e��L,��9/p#6E�6;	��2��є��#aSW
�-ʙS�}|0u�ɇ�ǩ�K�~U���ϻO�KOu�!�����9����|t��O]ڸ�Dȳ�C�Gn=�K7j����$�3A��*����'|G�O7�8Z��y<���P*�"D�k��|9mӣJ4@�֣��{ȭ�K���lr۩��E�3+��
�Z�0@���ξ�ȍxz�|�C̳5w�C���l3��$B��<�m}�f?��*W	W�ڥ4�nO��<�s���O���6n6L��%&F���f���qA]�i���LE��-�P�Qk�,w"7��
$��{�5,�,O��4�VS��A$MQ��u��y�g���܀�f�p�?��Z�RΡ���vz��K{ǸX�s@Ga����7pl� 4�;���;F�U�B��`P��ݒ9?�1�b�A��tL��Hc�]y{r7�[�����S���b��f�ˠ�>��J3���/�[D'NjJ㎑�ȳ��+cM]l�EU�Hc@&mV>l���s��?��!;���S);[��r6!޴ L�OC��n��,�=�t��A����`���ʟ�����a���I�m>�~&��O+���<1R lE)��[Z�����,K���(����6J8�2r���7��"'ہ���]ܓ�����T!J��a���eaR^�!A4Q� �H�~3��L�&��G���@K��� \���8b�o�����sv�e
۬�2�RB��ɀ��%�0\j���h݅�A����aOCL���T��]�,֡�
�	g\"]����Ҽ"L3�0L��P��vV|Lb�9� �ɷ�§*B�g�g����8|'�OKc�$6�UnK穧 '���૱t�X����Q��p�apB�)��K��:��}��	����ǫ�l4/�NlĦAf��vA]<x��v���?�g�����#È�ۖN���!y��}p3<���h��W,�#q�Ꚓ��V�Sil��";;Ss\��H(��z�R����9���q�R���Mq���;ٿ�\�-��E�#:�����[Lģ
W5B؆�H�#ɤAw�_�a� ��*�5�7�؈��6������=���Y��Z�94�!��G��"a�?�+g�voؘ��r�QF�{�Cn��-�q��JI���G$�
����b7���s@�Y��Q#��g�	XQ�P"]���O���"�:}Y�M74C���|�KݧR�tz�R�"@r���2����Hi��W8u��1�{���W��o���pM�;����W Oj����߹���ʽ5Ν�v�z V�0��n^ޜZ�#9@^��Ç�@�h�xmO�j$>�L��&sӨf��3³�����B�SL�k�H[tbm�Յc���Q��YЈ�Zԙ�{.�I�'SAl�_��"^��g�t3ܚ\��|�i�fE��,se�B_7��?��$F�S�:� d{�+m�)\]�nch&�ط�$��7/�GH5�����w#�p=��i�
��v�G�w	~����!�M�D׬�zr_������\�E�K��ze5%_T�7Z�?:�[q~gj�N����NF������E{F��e��@���Ig\�M��&C�2Ĕ�.*-��=��HC �����*��د�WH/8���<��^���߹ή/��5K�׆��<��!1��-DvH1#ƥ��(�[��ю�ŧ䷹�J(B\���ɝ�d��^����������Fu*hȦ|A��Z9����y�x�Ш�y���G�V_��h����'(��>UbF�h��'�h���ng�[�i���j���$הnK�(7Ph�*m�.b*��l��VGT���x�(U��m����l���d����~Tc+�r�)�4�c(J;x�{��@1�ST:{D(�� Iz�>��|VK:U��LH Z#�6*p5�Q�@��12�2 �R}B��FT��g�0��|��
��E��`����,bkج���6m|,�bl@�7h��za�OQ�wlÑ�r�̠�t��ۖg��H=���g��S��T�F�=V��j���W���Ò��'�	O�����Z��\�t&����Z���6��Rꔢ�!���(��N�<�_�V�N�Aez%������+����)�D[}����1�6�3����ulnl��4�az��tWy�&O��Ȑ!���W�T���$�#B⭾�����o�&�|��?He�!P�r���W�퓪	R?�����5Y9�A��P�9W0�����E�k�<�ʵ�fצ;I|'�4��Kl%_�u��"`�QRċAy�Yx'�b'�� �~S���u 5>c\>�v�ٖX���9�5f�.��@�Е)���2�]��\Q����d�%��=���fZ����,5=�7�@�.斃�#��b�,������4H9��u#u���W���`�a��a�Z���:x�0K�9�T`K�,��*[�RaP�kT����;�T���ͮ����Ӧ�[T琣Ĥ<;��0�<���Em�,����ö6�~�;�!�a9���1f`#��v��K��'jY�3�@M)�Fa��^�{$�~E�N�Y��M(�#�sli^�i�D�\�29�3>���Ȍ'���φG�h+�wQʇ��QJ�`�o�)�E.(BN�RI7�7�Lwl�#�D������:����D��T�c=��d��ε�>X[kO��c��s�(��U�N������O�ålǚ�;�:��'�&O�]vY5��7�Ī���w�A��괅��@���P���)c�Y����O[�O�>��ƈ9����UU��=������)�Hh�q êb���곛��_ߝ��O"TP?	�����=���{BSj�D21f��*�d�:ac�q��R�bȰ@@�.�-�&��D�[�/C���w��U"�^Et�-��0:�e�OP
�k�:��,O�	�f���U�B\�zv��S4��d�m�Ӻ��ӊE�`�R����B�7̭Z�������tٮL� fOB�s�j�jw�&�C�ס��'�[�O��
��KɢB��{�]��ݣ�}���K�UO����C�5�t���	�nu��l)瑋~�$ ����Y�~r؋d0�{�X ���}vU�K���T̎�+t�ˀ�4�Ҏ4F��`��s����i5���b=w�t�2��<T�D���y;]NO�yd�s��\t>Yi�|G�b�Pi�-~/��}X�0���O�1���v�E���.�5�'�"�3�����4�k�r�I�ͱ}"g��&�z_�S�	s!�e�V�n_�W2υ�u}-J��6$�8q��ҏri�ԿJ�GR�X�w3���<3D.r.nҳIO�5>�������p���!1�ރ/~㆟.g.LF0_��"�D(��K�B@����ꇿ���S!��Ϡ�F�����_�fN�[iSH�(����t��|��4S"��.�3ؤ(ᰃn�C%���I�� \�'�����7��E�Ϯ�����>Ì�-ٮ�O���i=�c��@�(�!��h}x���bw���^�l���ʸ���%J�_I��YQ�
�f�mnQ�`��v˟��u�ՐxY:�lY�^�>G1����6;8�$3[�}�w{d >�IZ��
w�?�C�t�m���'�'�Q�1�߲7p1;>��3a��G���Yd6ǟ��7�;(�O���K"��ޜs��>W�7��Z$'�S��D������m`���,�H��*�v��T7r��G|��S:Z��"<��mMX.T��S�W�M4�F'ڡh�S��9Q\q��4!b#�L�ʄc1����c�x��%��a,�>��*�zS�̵�Y��u1G�����yb�R�<!S��Y/&X�%�t��H_k��vd�7pȱOce�z]���Kn�����p,��7�J�>��=��*l��]@+�1���%.9�Z'R�ܖ�d�7�+ۂ���r��:�4�����*�Z`NH_�;�@ؘ�Y��|�H��=��dur�]��[���!�G0 �����+<�����ěFKJڐ��]����[0���]� m��C!PT�`9�}�Q q�/��	{G��/1����?����c�5�D���~V�(A^�d&��X4�P�������gU�L�u:��I�h�}K'�;��xϙعRq���Ssf���E ^[Ŵ;��	��1b�����]����^��\�H.!ƔW���K]��.�Jɤ�BhF�-���=�gj�\�vձ�UPZ�L��
!r�k��u� �PL�
K3�:M�4�*�K:�Ꝕ�Z�^�!̥�����ic ��[6Et�"rS�<�[ɿ��+r��䛝oR@_�5�Q��7�7mӸ���hXv�6�[�DҌ�8�-�AtV�:1�>Ŭ��:М��  � :T�j�{��|�L����R���Kʶ�]!�!%�G3-T�*%qr�.Ja
���f�x��>�}�g��륃�"��?�m�_A����?Es.��j%~���J��͜jS�B�dR#���W˻0���! Q��\\5}N0ۜ�*��̎M*�t�L�ꄚP�3K	��_��`��������B�����i��J��[uЪ�6�y�>��S��5(��x�F��W��u�q�s���eȘNn��t�%�֙�9jQS!�	���Nك�D%h�v��`�j�WGxx���$���ө����[�ݳ�Up��ct���C�W�*���11<�M��t���W�����Y���F�hTt�W̸}�|1A��Mn���ֶ���/86������>I���g�I�f?BNd{�xW=A�}��0PK�X`Z��)�8e�0�����+B.֠�A �ۢr�Z:ӎ�P��8D���f��{�Ӛ�]sNCx-�,�eB����|�9���1_�]�N��-*b�~���-R_,@+��-�jK~t� �=��d�F��G.�FձS�86���������[|�����Nޤi8�j�N{En�t�L�� j%E�p�|�Y��t�63C�J��}$j�+�e:M!+�Q�C}�[$�����̐��L�$����߳&����h^J����Ӳ�*s�D?\��J��:���Z#�����O㠘��W��c3ؼF�G�%������Gi�ٸ�i��g)�u��J��T�$A.����6�tj��l[Bp"tL�48CT��9����%-^	��n���l�r���7����1��^�����L�zrp;��ߞ�qU[^p`��ZR�8��@E��Ej�Q�;���]25k���HN����HFۻ �ut�/ ՞J�E�;�����Ѯ4p���hZ�Z^��?�h�����?P���ńAf�G����x3䟰y�G����T�Vj�>�]��	����yzŃ�.��ZyWj���P�:�*к�dzT}�ɾ@l�՘�j�ԣ|��]:���Wk�J
)��#��Iy�=��6w3��B��;ρQ�`W� y���/�^���R;�}Ӊ�Hꁘ�HS��Ь�8S��ʣ@�ͦ/%�l�z���8��>*�����75Y�sL~wi��u�e�������|i}@�a���B�v��!�N��u5`��vd��_b#	�l�cp�:�0S�T��}���~,ag���8M�=#�����ASO���ֶ{���; P	�V��٠-�I��m5>�����pSC ���N2td�L_YJ���{VW�hxT�Ԥ�T�f���&+�X�s�$�g���.'�
�q�8֑6��y�3�yh��+8��Ax}�r�Gl�:Db�)X|���9���h +Z*���C~}�
V��=F�Ǉ�c��ҭ��%��s�0�r��k_�0�����B�'��� �������
 ��Gkh�F�b�̵�>	^nW��'�U�6��d 3vH�t�S_�턜7e����^�=o�,�z4w��H���|�o�^�.�cebB֏���2E��]�����F��H�2,f��j�v�ߍEj֮�й��-�~�ٝ�`�c���1�M��d�I��I�]�T��<�1�����x��f]~���(Nh_do�..�_��GhlQ: 0֦.����o��Ǳ)�39��)���D�8a����i�`#tV�y�c"zM;�J[�ʅKk�a/:ು�Rq������}|�kS�m�=R���������٥{)-=��%9z7J"�Sݱ~�j3T�|�=T���CyN�jɎ �K>�:�e���ɞ��NYBm.K�M����X��'@��U����0&���ȴ�ޜ�w�D��R��6�v/A��+=�=��=\� �����mM���c	dEٴ�a��u��7��_�� c7�l2�����p�����|0�l����k���/��ŎRe�	'W�ա�ǆ�q��CdQe����a���䎿"���;�^T/��hƑ��������L{��6����xB��am�W�T�ᕊ�Ϝ����1��ET�xZh*�b�bA!4K�ȁĞ$Q�ORϮ�!0-Bu����/L�`��Cm;��Tf�nl��=>ku�ɌM�5nvъ 	8�A,Y[������u��(A�)���_�іkra~y�CU�Ѓ��-�z�?�[�r;�T��E�p#{ڕM�����ڬ�WD��� s��h Bh��������8��c�����Ŗ��&��=�(�¶��U�>��\ˣM��uc�ۢ&��V8"��xV��3(�\�?�5K�Am��1��g���j_���"���<�&Gyr��]�EEw�ֲ��Å�'��=j#�¥���/�x�=�$WD�����y�ɳ�A�.��������ve0��Eo�Ӥ��&3���EʌS܁�v�~sV�P�M��'��lu�|�%���z��O��''�X��8���ᰶMk∔�EJ1Y<� {�V/�%@��sv�Q�j������vN�� 6��Pn���!A}ض c���_C[Ӛ�n�M�I2Fe��dHr�E=�������)�x��R�]#_�+��%�c�Q���U�CID#�J.k�!�O�q�@����O߭����C�5�����D(����/�b��E�}8��"���x-��P�t��7O薠C��lyB7�6 
�'ڇ�V����r �Z���i�؂u�j�(�3U�챒���@t�p>9��8u�f_�X���l��&G~���� ��3s0{���~�<�:���� ��s�f!��,��i�\��S�}O߃�q�d�Ͽ�� q����Q�&T�O��?��D��M)�	������ȱyH�h�Q�M�J�B��� 	�!��i'd�����MT��(�5�wA(autr��7�Z[4����^�T,[��Z*��nK����Ԙ�'�?A2���&5#p�3��� ��1r�ds�)Z]5�Ty��9��dU�0�R����5�U��ж nc��I�>��fR�f |D�~N�����]�ހ��叨����퇐h�;�V�����<�S#Y"�!�Z0����ı�"���k� �\��	/��n~-^9���uR�p�)�B�zp�~��p^�8���E\���8UK?JP
5#^}ԩ�[���;�Uo��IL��`3N�F�ln�w����%�lx�D�{�
9���=ݣ!m!��l������m����ڨ~L�D�վUk8:��1���S����LcYq	��[T`��#EF�4A+.�����!=�AE�W�ϋՇ�d�[�4����U�<d9���z$����c�e 
H�|�?���/=�hz�y��0h�DM���+0yG|�ڀ+g-,�+�7����s6_�_�ħ�T�c0��"�H> N�W�R7w8����7���V*��H���R��	*-�LVr7E� >�7\~�:��Х��P�c�,�)=�
�iX)?m�������������,�aDEX�[~k�蛄�a�&R��u��l�����=����3�1�V�!0��4��A�N�aٶ��E�4ݮ(}�	~Wj����6��ճZn��\�nD��R�Om�5C�{�l'9���`f~-�pt.Q�(�I�� � ��X%���:�`_S�W��!��G�ȇ�2�p'抸ͻb��.px�2������l��{���%Un1W�DR�2�{5x���3���б QTA�R�l����!�
��̓��С��V������ o^C�=x�Ǯ0@����,(�~��͎&w�/�h�UM[rn�>��q��H 4�-�P�v'.z�Ǟ��<��/c��X\��G�z�QF��z=��_����Ni�7�,b	��b!V���s�F��e>B�Ǩ��;	��?���V�R�G�LxUВ*�C����|-I]]��O�Uc�o:�z+�Il�r��,=\��}������eۤy$�>H�=�W74��*��'2�o�!���A�	Br�,��!+�%��� ���n�5�Dss4���2����,A�I��d1Cϣ�Ya���~RlO���z�m����&g�e�p$e����?��U����e���#z�M	]N��hG�����_4G��� ~�5j��S�If�?D.��i@) ��[�,:T��A���	�x
tA����H�|4��^㖔3L�8gy�C�޷he��:�<�u`H5�)XI|�|�;N��K���߄��U���X3���>�tNo���J��"�Q��X;��{��O$E�v7#���Qwǥp��������ЉD�����5��f��i\�70g)Sh+�\��T(���������>({��ɘ��/�H(�jcd��� 's��.��,�������-�"����%Ό`�ቒ�����p�T]������UfŅБ��o����wxm�VW'��}�R-c8U�����[�w��=��Z��Aq�fy����<^��e#�{�Jض�����?Vy����S��O�N,tL��؛]Kq���:�-�|0��,J�/i�߹�f�5��#�ß�4�
���J�	�,e+�� $�g��1ܞ����=0}�G���`GD��x�.Ɏ��.� ����4����O ��}�O�㰬B��F��I|�b�.�%�)%�Հ4��9o�q^J��������GV��,;�.?e+� ��,)�uR�y�D*��1U�磊,�Y�]��Z��.�H>*,��GF����T��!���u��'n�g;^��(��"$t��w=�f�VvjD=��ť��UD�&p��&�6���Wm^	ƚ��-����I-��u� J��30�M�Ӈl�w�T����xA+�X�у��zz�l�4쑰��Ռ��H_�'��pqޯ���_��zW4��k�5�l������f|m�l�X���ЛQ;84�=��C6c�MIUx�Ĩj�_Z$�"Hתoj�QܟqW���F�PI~������SI7èP�$�%¡��U�:
+�W�l�k��'B��y?4b��@�����������eW���Pӄ@weIbW5?*!��vxk�[�8}x��3�x���]��^6(񲢻���(���+P������v�M��V8��S�o�(U8�k.v�8lF��ܜݬQ��ې�\|TN$�}-@g�<��Ȳ�&�q�~�G��_�2b�İ<���ԜpU�S����}qã۟X�F }7nI�{W,��� �A�z�y'-��ϫ�[_�/ 0��>�z>{JR�L`�,��i�\L���(�lt��y��O`���ۖ��+�Ӏ��A`��Fnd��>_��~��x�ǑG���OB�.L��:�k�g��*\�É>�nR����0C�}������ ���vk��� /�ʊB,�d�p?m}lg�s���a/�ox;�a�ԍR*+�@�/n���3:_�0���1��Ӗ�w�s路�{����6v���w �z�$vx����nt��<ҭ�d�-�ܛU0�$!���'ލF%�t�9 uV��2��ׄ(�p�\9w)1�I�T^DH��Ļ�q��fh5�`5erC�2��1��Ȇ��3s�0�vtt�#>�G�0��t�N$v�6��v��g�0zHV�?U�۟F* i���2`��'���s�g��5�IPf��X�ݿl�s��OƬ�����ػ�R &��;��<f�$�M�W�Q��"���_yg�;J��gR��Mҹe9;y/>��$��Tsx�^��	�"{5�%��a+�0D��T"�f����La�KBHUs}���[�x�T"�f�o�c�5�q��3ܘ
f7�8�V�f�i���#:Nװr�M��?��n�V��OMၴh$!�4=F�XQ��ꈫpe�w��l�D�O�1����49�s�`�(H�����1^-�	�����G�M�����s����)J8��eB�U!�II�_ˌ���g*�"�4#���X�x �N�h����l0�H�g�`ϵƲ�@�JD�37m!��^�fH�p�{.ǳ��|�dIjy��Y��li.��u_\)V2���t�WX���P��DL�[h��z�|�T���|D�'u��;l�	�0xl�GuX�K*	 ϩ�վ�#��:-����_�/�_H��!�Hk�H������0�SjS��1��ͅW?�lc�v��X������z�O��W?&��v�}�E`s���Ȅ����/8��.WtQ��W���KK�$�d�8�Y�E�T%�W����:bF/|v�xU�F��FC���YoR���JONġ;)4>'Ѐ����S\�6�#&\<��2�K���p�ϵ̢�#������D�R��pY:��`2��Ğ[mIZJV������8ab�,�=>h����=%�	�]��Et�:��n��9#������>5�l6a�8D��v��)om9�:�v$�w3���a�����ceK�C�4S�Y;���E�q%� �=2��R"��Ei���vǂ�4�M�I�}[��dfs��/��b��.p��7�=q����z8Ҍ�#X�|�{����xmPn�}[�'2�z_�f$����1�dQy������Z�KH~����x/1%�7[����W̶Uz������Q��J��uܴC�m��ܛ�<�L����X�����B�`O�˹�nW��7���$��ń��YX�e�����.��e���e�ʪ��:*+Bc��TN�xKy'���q�0>�\!��z5`��X�z��Ը��G0~	���{�}��ʯu|�2gL��<^���\�D�n��	:�������|
�l� y7oE�j��۝����C���S��#[�M��S����]t"��H��QdE����;>�.�Y*-�����������v�m:���f�'�.�WG�� K3��|�:�Q��E`L���A�|-�|<�xR*X�)hu�'�13AUY���o��&v�$;��~�q�b0�9��To�Hw��gW95/	/�]G�鴷����o��/�ʳsz:lMZ��u�=r�e�F��j"�Rj�%Y+бl��+ù����*$Ob&��ع[�@ftv>���:��~�;��,���R��u5\U�an��m� ;o!t��<b?~�.M�֋ů���P<C���Ug���n�n���d���Msp��|p�>Tx2mae���'�� ���0M�7!l�;�X��a�V	�.��Ƒi�`^LHsy���]�zb�+b������f��JDs�K��F)�$Z�ő�1��/p�B ���NIL3�6Ӭc9��ww��8����I�t��	�ﰣz.Z3��ڣ����k�iy`_)�'K�P�-���Z�Ð�>�]D��k,4�»��[�A�R�a� [Q|9��5Dsɞ���tS�/��N�@>�GY��
\�%E�!�����f2�=̐c
L�a��dJ�{o�����Щ���\ŷr�~}mjm!�|�OC.,ԑEbt�UD�ר�N]��8�O���������J��ْK'�8��ܬ
ß�;>�Op���X� �v����Qz��q�0��T�?����1>�V22i�\Do���_�+8Z�Z534��/�q4�k#WH�u2k� ��}TC�26�P��#O���¡s�&A� �FT�p{�+�f�^RC�t���[�<��v/ǽ�M|��� ~�����r!�a��B���vT�V!��?�`�$�+[��%Fxgn� w�h�Mee����	-Q6ys��s+7�1��V�Qx3���ޝ�·�y�OW�}.�3�ΡH@��&����K�઻��wh�g�s����ꌽ�s��{�t��8��F�:������Z�Mƈ�nظZ@�X
�����A���e�Ҫ["|A��gLW��R�V�s�Q/t����Ͼr�mat|�'�[1o�ÅbC�e�3��~��2֠�Z�Y�*_Ppl�}�p�k��S%>m>�*ϰ#{+��d��}I��W-�e=�qh'�R����2��H�Y��V�н5�lu(=���&V�髸7.K��՚�f1�����g')��<�3s�O�nO�^�D�ԛ��T�򱠖�mB !h��!HP�e��=|��3IX����4���������M˷v|�.� k�}]k�������|���I%��=E����0əޫ�q���ܓ�X+/�gHh/s�<�ARY��eb����G�Fwn�î�]��s����O���aP����b�CC��+�����5<p�|al�	 ʮY�C�AM�u���$�T��#�3�Q}����ݾ��Dr��;W��?�+���]K4.����#$n�(��Q�.��1��΋jM4`[��8/��t�t�}&Ŧs�r#e;HfS�x!���<庛{�6c�PE��mo�_�Ɨ i��ĭ~����C�.��FA��|�$*T�ky(ء�h��M���A�=�=֫�sw.�����%��+]�K�A���TbAߡU}p�q�9��=X�mQ�QFu��,����#��$,��t�;戧�-�������
�ĨWyo9�;Z��l���m3K�fS���D��#�_O[����p,׾@)�F���z���%<a�C.�."4f��c��2߄�Q����Ce�������IJ�Hn��إ���n"(}��&#�8�
���e8�|�OL(���z�Cъ�Ɲ�x;cZ��&�V�^��u_�L�,F�ǲ��@V�J�,���(S�T���K�U��髹eS��>K�[�~_2��"<�m�z�J�!e���6���U�gͦ�ڂ�Ǫ�[�?53(��?��y8΄�%Aď��ճ��Nq%������3rS��F�$dx��S^vM�%���W2s�M��}?=!Te@��3?�c�t4��>ҙ��q��G���;� � 	���42~u� ���Oǌ�T��FB��"���^�Z���L���c'��>j�`Ѹ���[˩;
�P*�%R��o��&��:�ٱro��Y���:�=�L�J9\y
dcP���˸Nl�&z�|S_�]����dH�j�U^��{"�O�c�B�|Z��`ѥ(l�(ʛm;R�m�w+�<Qe�$�.G}��2�6�y4�?��H����b)$q �����z���J�=HE�t����=N��𿭌l� 6������`���!�������Y�a�"��P�w͠�K�]����C���w �)x��ۨzk�x������S@�W���hr������W��Y#�G��H&�ʠ4��T��5��B	�},�s�>T!7y�S�=�I��R�@����2tR�v�b`6�-Hş3/�FҎ���gX�Dx����I �y_(�O��l�=���|}␞��v����ݚ��ɞؑ�����+ �Ȅ>&��C��i��;���K �`�
��Q�����XuQ�҉1#�1q}�3�t�2�*L��}ݓ:H��@	b}�4G���y�nh~
$}Z<H���\��Xjѭ���Z�����#��mUc�A�=��s�)����}O��-q��&5�k ��\�K��:
8	�[I�Fœ�M%Ti3� �p����V�����W1�6 ��a
�ڰ�-���0L#}ž�`B�G���4�a����#�E̞܀��U�x�IY�+l)�vf#S�D��C|%�Y�9�Ak�{~��|�I|
��w@�a��/ƚ=�m8��32 0�%���,R��bȑ�Q�6(u<�O�I9��$��������R�ޘi�x���`t�)1��
�p��d�f��4�C�}���X{t�oZ��Bu<X�F���bo�[���݈������lW�;��ovrw1Lx��Zڸ��9k�e��+E (@���'?���8EA���|�1�E��Q�g�rd��""��ȓ���f��@�x@h���m�r����,�z��1[�h�n��� �?n��g _�{��ZY����B1DoG��M�xwŻ[�J�E&a�;�����slv�K�<��Uշ�:�b+���ʀ�=������m��YY)����D��ʸdjΠl����r�~��^��[�v�+9K��j�F���B�����P��os2[�Z�G��8-�\v1B����-��Ұ������4��3N���[�S��ߠh\5�����h�b��kP����zi�[�c�l�E����f���Wq�"W�ݟ�`\�9�wO0FY�?�LB�\>Yې�I*5F1�x�?��Ҧ��	1�ϐ�'����?x;��`t����D�m�b�Ep�6�_Α!-�Q|3R�m�ɷH�`����%�V7l#�D2���[��g"z��K�qj���>Ǔ�����۱�L��呪,a�HC�+����g�w`3���{��䐆P������c̾����n�$�c��Q�~�V�J_��N((,$H� �-V	�Ap�I��s�"rl�-s�=�V@慱���@���HW[��^�4Q�I�=���(��W��1����з�`�7g����^V)b-%��MA?�>ն��)e� w]��y����j��>gs���L�C6������Ͻ8� T��\��!��k�� �k7,��:nC���xa�{r���ţYf���Q:K�	/�?o�Y;e���)R���#%g~nN�TMe�d���Q�o��=����rN���3�=�~o辠򌜙�#f1��Z������Q�7����ׂ�9r?���~t ����f�R�#����WG�"�i�^6��ڬG߼��:��Ҳ���Q��#��<3D��zs�w
PnD�N�^`��`�~}X����-Q���1����*�3�ڡ˛꾣���k��Z�&��lU`�E���Ԍ�(�}PϜ1��1Ϗ<܆/���?�Ѩq�!F�@�()q��b)����AMF��【�
0� b�z����}�����ZY�[�2�QH�}�,��w��)QL$��EN��=��Y
�;=����-��]bbu���5���JUǩ"�p�S�t��gAD�ڶ��i�Nni�ӄ��̡����1Ӳx���g�QB��]�}�Y.��ݓ�7ɓ$�l���T��E�m�Od��v�Ab<�ZJ�_m�4ף�����k	�Ɏ�О!�l���B���m��[6��	� u���&�*� �9Ȁp<�\|kd1�Jx)�H�X��u�|�d͗�/q���%1ĉ�LG��Y��H��9��i��Ƣ}�=��K�I�d''��a�˯:Jv�C�sJ	q8�@Z����e~ٙ.K�� �b#~���S����	���ވ�zP���L��]0�(SdӃ fnu�}�[�v W�z��@)-0��>}�4�B�g��ǔ��
�q�J�v-`8�{��t�*Q����hC�/�.%�e�*��kv	�,�/N�q{�XI�aj��G�L�z�v�%|
�`�A><��~I�&jڜ��-���H˱-�Jkz��fV�#��U>o�����v��Ty��6���uu��f�	`��,�&�� d<��� �g�<�?oͬ��̱)��z�����r��5G�v{>�>��.�?�m��Fe��Y�W����Cږ�|���t��穻:v�9�Ɖ���$Q�k�s��PQ�_�|}V$m������ ���@��t��jV5E�ѸY?:�T<M��0�ǫ�����Kd��^v��q�0�2��B�*��7fQ�ۛ8�(���҂�\G!,�;��}iF>'_O�ؽ���D���r�Oq���޿b�!���qԨv�<��`���?=4��!�	}w������R�����x?5����W+#�x��o�^c�b(��1X���,}�5��N�k��bT$f�`�̛�P���,r`�Y%�6�>W�:��o��.��g8X��C�^ѓ�Nty��"u�M8�V��2E�;�e��M�/Zž��Vti�dٛ�����������z���Y<�*������<�$V$�O��,W`�^��^W��9f�k��c�������B0�*���%�qQe��6�i�\��~�	7�mx�xxz���H�%�nbkU[ї"�=Kq���wP�(�����uC��c !l�%Ҁ��X��yzP2u���;����|���~A�R��CVxzT��T�EBXO8u�ӱ�,�ez@�j�rE6�	�����ywH�X�>��~��o?pע�݋���v[����w^�Ń��Ga�g����Z1�,�'��/��]A&l����3�	��I[:�L��V�1�BEs��r�R�ζ�0i0�GZ��K�ߊc����~�I�z��^i�3�Vۅ�%[�Z�%ݐWM� �&��+�n
��ΏH�-|�B@}H!�b��g�A��X���'���>���KpX|S-�%������/��kO�?�}i1G�&��	�,�SbVьj����>$�0T�1j`ka��?�J���I��lR�K� ]�noj�����Fg�MAfKs�+�D���%Ǧ��8��5���^�3}	� ����&���G�ϹY�Yƞ�i饛���ҺRB��l9�0d��4�?@]�J�����	�ᙘ+�.�C.�{8a�Vj��wd'%ҳR�2�_kx���SeP��Q
���ͭa3�J�#������ē�)�
�m���)��C`?�hT�
�*��cp������kb�@!�IY
5X_��%���]�jq�֢�M��LPD@m���C��qƨ�xZ�������hxi
��ّN5�d�{�� ��Ko�)T�����z�[}�5�p��om^hW~}6�<������j��֞��T{a:�Bs}��S�}�!�`h��4l̮=8&��e�M�ȂH`�'
<�	�K��
?�4U7A`�ڈ����H?��R�t���L|4>/7���w������2Oa�k54b��l��'��7�v�B$@:��D�i^����7|N�!���˒��)~:��:�V]Ş��*�ʝ�b��=��?����F%Ν�/�+q��/-w�������q~~��!Ö
��A��!܎���w����.��8�1#��wMm�N�U�K�p����5_��,�O�.�����4�����@$1ꤢ�r���X[&h+��I-�U-�����5p]8�ى\�%i_���j;{���rUQ��'��^`Y��p��ب���T&)E�
�_�,�pFo��ؚ@V=o��v�����J��$ȵ�H=	�`̺o��ڞi˭4X0�w��+%Xb����x��m�<���o:.�oy��K��qpy�U��sεT`ԦO3��$5�8 ��k�����C����r�y ~��@�
*ѳQ2$�H����q�ҲA�w��chAë%_��Kٷ]��.z%anح��A:hY���<�]�q�=*�a�_���x���eX�S�ޙ��ؤ��#	ia��q�M10�QŽ�QM))�Yt��I�=I��d��¯�u��U�璬�h@A��hY_C2F��,]w^�C>�`Q�M�<	��X��)�d����C����`��^h<�b�H����EC>��b:Gd���}�q��`hS���($^�`�b�;�4����͖�>�)������T�Jo�HZ8�QJ�ఖĜ�Q"�tS�^�i�Dܮ���%��\<+��D.Ǯ0R)���a3��3�5��y?��C{K���������HS���a	��_r�F��*���{�A��D�-��t�j����g�M�!�)��Е���F�v1���'����5\��vN�нP������"H@�ԕa�j �Ԕj�j�7����O�.<��u>���lX*.�S0(.��:�5%/4	�V�*�P�򐘐��d���w�̶������r >����ݍnе��F��U�%{���M%kI���F��h�I#oMuR��h�߫�y�JS��ѻ���c�����dЫ>o����AX�����MV�?��;�wWT��S<Z���ʒ�8��)�E��֡ٹ��F��{�p*e�#a ��5�����ҡ�^�|@_*���dk�x�k�k�Pk��LA!b'��ܯx;�����2_[&��nTE!�9XT�YF���s���əgRq����L��mD	�m�S'�#���<����ʽB����M�9P�ok�|: �3'"PL�f� ���e"�r;�n9�ƲqBځw[��Cn����^�lj,]�d�НI���������6!�N��CQ��d٠� ߚ��}�^�C>fl6�9��c-�M�Mr#��5�;�]�@��z�����";o���뷿���R�`�a������R��)@D�����V�O���a��A��xAv#�-i���s��?�����*X��=�����#��q)�O5V����,���1��"�N�@��q|��ύۂT�(^������(��I��
�~fRD�m`�)�؍�q��ޱ�'���\;Z��Od�-G���Ӹ���|j�Kx�$]VC�i{8!ރ��R��Vp�0X�4/�9g��Bz�K�'E��&c����eNB���_�2���7�w���q��� ��2M;�M��NB�|(o��՝|��5���o4��3JQ�)!l��;w����*��Y!;�-Yz�������m�Y�G��}a�yeݓ��|�X[d�
��E�~����E:���*$��FX�F�%)ǸF�a 3Q��JG!�����K|8����ˆi��{ʍh=@3!��Ł2�o�O{?C��Bw�ҳ��@ty�?C]�� ��ϔR ��`���v@2j�������L"t�{�l�D�|J����̵}\��u.���B;�@���JxE��DI����������(�u���@KA��f8b}V,>��TP�Z�F�i��G���r�HZ�W��P��0''E~#��zԾ�y����l��aˑ�Tm�Q!��p����x�00ȧ;2�g�9s�c:
��s�d��|�'0=c�z=PR��������Wt��@%�)�l�R��e���y�G �"���j�~~q��O��v0�Ik`i�l��U?)���f�[fkX��'
�
����qg W��=@�;c��݉��l� =�2oc�y;��Z��*"n�v�$g����FD�D��"�6m�]*ܫ�L^�.��R��T�?�9A��5Œ�
��t
�0.�qa�D����|�)z4��X*ʪ�R�P�,�%��p`�� h������H����#�@����?��#�L�>�]��:yhW��:��d��ή���SX)��Pxѷ��*�
��wݢ�����w��P[o#�d����_ʈ6Yz��n	���$�������)>&�v ���9K�F;tT���	��ٕ;�ٽ�j�۱Վ���C(�������`�ua;F�UK�г��1�#fWb�� ?����m.�%���N����x�A7���$�YIq׽�}�%Q�ZLR��%��3r("��(����I'rWa���&k�ٚ�g�_�jy��	�c��W>���'��A��0�Kz9$��VH*0=	EՐ�e6��������<��h��H���3�+更����,�	M'�~����.�N�E��w��H��.׹q	r=�U�F�U�\c�n������w� \ۈ�Cr���Mղd�5��k����L�g�~�w�7���B�Ңyf�j���Rd�O7﹉�*Z�ќ�o��j�}���;S8ĦC���7�5�k8w����и��q�!�}0�ur����k��XB� I���v��15eV���uk���H���1������6�CY,U���x�v$��
J;a�P*+�W�T%aN qUd��A�H�y�B�dmYH�Z�V�H}1 a���
-J��S�y�s:��۪>�O$hj	�����j,D�ux���< ϹD�U�C�M�;'��Т�X�O���8I5H���F%|>a��S���E�,��H���#^�>�2��+��	X.<���b��T��d��w�ߡ���m���34Ρ9ŭv��Ug�T"�kI%�XyO���U�[oe�a@�����_4��cF�Ǿ�72��B�EU-���N�Ȇp���b4l�3~kb̲�Z����o�¤V�9i�m�˒X����փ�v, sF����!�e2������V�yfϧ�t�x'@\�$��g}�&�UK��Y��i=oA��g��.3#��6u�;��t�?9�?8����F8�S3H,/��`X���鍗L��=�^<�T��s�X A�'ҙ*�@v|�}�b��+�\c��իU���q�a��C����yh2(V�su_r��њ�w� g.�k㒔�
�k�Gns�ZݤCF�'�9��>H������K��{fWk��X5����H���[J����	�$�LS�#�E;k%4?����1ibd���L?A��s\�r2&J%i>����o���܈�P�5߂+�pN�~�E`��,��Tj2lN-P�mt�j��'��3ܴ���D�f�L��}�Q���[������3Ws�����/��4�+E�����v�^����l�_��yΪ\��P�<, ��c��L���T@�i=j�)�ĭ��E6��	ufE���8$ ��&RM;|�W�"���)`^E9���LM����4�)>�ޫ����Z���Աf�*F��t"㞰)�})4�xn�d!�w�a� ��WB�*cCOoğX��E#�d��R��c/�)w��8��W!p`�;�RLZ�+n�V�{�8�{�=Q0TGx�t��w��c�b�U��~Ww���7�h$��5+iz��F�*����R�$m�y}�`D����E�ځD��zjUE���xz���
SP�q��ژ6{�`���[K�YS�*&�M���ʶ��N�UP�Uc%�}6�e_�K����=�	��<)�u�ew<�YH��N%��}h��u�Bn���e�3<�0�c�@U�0 ��=��?�"!-/�!L�ۄ\z<W�,T�6~�7*�������9�{����}���;Gڃ�U�R��ǜ��loɠ%���*C[���g�����A!��(jT&9����S�I���3�@���~�A��E��-[�b��	�T�4,0���`��BD=�zh�<�Bc3�� ��X|�O����7#� �B�cQe���y�tp��YK]�@��N�|�teRǝz���"	�����W~k��/f��Nn�����O?)�
�$ 0֒~]�kL�ng͇�t�n!��!�(����b�e�y�o=�F�B�CK��R�������-�� ��-���3�W0c�vlo�>��L��.��}rچ=��K���-
��ZDc�!�����LD�(q��k�\���u0��̟NMF�k��]V�[�ZW�U]1�3ꍥQ��8�T��+��/�R_���7�~L�4�?W	�Z���!]�Rh��e�?xYV�S��|	�|��>*�^�9T80q?F���AQ*�����!1MF��uKR�{@�����\eF����Ta��H_���+�C�A�&<6e��s���6Q>�#V�uz�G��p8סހ���=ͼR5^��Br�Xn]8�%�`N����+��C��$���С@k��Z��
��Ϝ�(P��^)B�>� �wE��W8�6����60�v
�?L1���g��ݚ�(I7�#&>�`�r�2��7����ސE�(�[Fr'l��ɧ{���8-�]�fR����I�ԃ_Ӊ��:��l��K�Jڪ:W%�?rʘRD��YA�O
p�.��/\þY�`N���Z�Z�.^�13;t���1
�x��Y/��F�^��!C��A���l�H�pV.���_���,%�Y+��$�n���3��Y��hx��8�g��kom�]O�W��G	�xEth�:5;�g��Ԝa����O3-����i�nYkjAu_�Ү�kVLyu�i���{�pH����>?��ێ����u�VL��`���v�X?�cfa.�i��ܙ�(4pφ&$]E����R�**V����W�Ն6B>��~��=�[���L��(B8"�)�Oa���^Y�JP>@��E��9��^��e�:Z|��n+?��s�L�U���V��D�J�1�f�I� �M^��i_X�t��.���Huo�޵aie �1�Bl�Y��\JiǶ�_ʅ��V�� ��&��or9�҉I�~�KAª�ְ\(n$-�R��v�yhR�;23����jT�t��q��mܜ<�{��#�ي�&j2�u��w�^�9�%2��&�
�q_ k���u��r5���Њ��$��}��Í������|zq֗j;����v}��lig��L�è�	fn�;ȇ��
W��+f�^F'+�d�l��ν�5 ����H٬�x���ͥ�@�cvXB�R��7uN��I׏�>�����9��\�#�-5�﷬*z�c�aU �]� /�b�;-u~,8c4� I���6���O���#�f�eVx3�'z3;�ǝ#�~w�W\xE���Ƃr)� 8!y���Ѝ��F;�k���s�J�����u�����"֕8�^�y:�%6ĬB`�V�^[�i3�G��K���|��LA�O�1���[����R@���p�Fq��< K���>3�4yDJe���y����s�	@��T���ˎ��EIk�s���88�f@�f���U;�E�'p����)�	�+��-�0kȢ�&�ᰧ�
�K�m�ni�Q��,j$���3=V�R��wB�����=��;c��JrA�68�9)+ƃ�~�[����^y�cM��\Y�tR�P��B�>����*a�����BZ%rA��R�C�Ԩ����z\��z�"����銕8k�վ�O'g7�Ճ�w��$���~��wݩ��/�:;>����Ɩ1Bé�	
�f{��}dUG��?���6cO��L�(�u)����m�TX
|l_�1���h5ǍWB���@�$������m�;?+ώ�����P���w��E�������0���;����m�a=��i�B�n73dAn=ZK�Pf�ls�>kR����Ȕc�5zD��8_4k��X �^�o�\���Ð��<�S����tH��Wz�����-�ZIV�;�k�	3L��#a���\_:��)��

: J�X{�W�3�u����|��*�w�W�1D#\[.��ﱭX�ݩoD�ݵ�J<rܞ�7�wE�?%�nř�����֦��@c�
���dQu����(hO�g�W��]�(r\�t�F��!]��'2͚��-�G��i��p����q�Y������;z�����[�˗�=Vcd�.�G�t����O�:�ML&ފ�Wu��Ou�C��˲��Yv���������09���W4���h��Ӱ�诈�P�#D�Qsi�8("/7�B��Ɲ���Ŀ9���.�#;���Tf?��=���R��C��h�����v�!aŔ�Y������b[�s��O�\�iE��/sL��!X�[�V\p��>�7��T��I�Ce�&�	���Yd���R�@ޡ'Ub
w�O��Ax�c�$���I��ur�I�޺�B;It�U�|]R��k~TY�~k�����)�&(ٓ�N�KhZEhUnu�+�w�,�cQ<���,3)����6�;���ٯK���9N�_u��'����#*�z�f�e>e{K���3f��U��н�5<ςGj�}f�PU�9�qH��;�}'W%�S���;Jѵ�TlV@�	|4��U���>\��GVR�+/Jq���m���/7�ۺ�Ю6d8�4���J������5�4duF(��&��pa�7FI�'�D����U��&ޛ"ĸ8�v�]� �^����q�_R� ����_��@/�Cc[cK~�I��J ��}�i���`� �b˚I?vP���t���~ǋ�X6?��d�ӵ��t���ֺ�n>�y$i�笸w°�+�Q%/pҮ ��t!�8�P�\��s��w��bgFp�[���s3Υ~���U8�?i����R~LQD�ZA\�4~:��<���1�P����[��e�\;3m�Z�O�&���L�h."��OC����8�,\�m�h:{�z;����DfとxQ_������:�K��҈���r�����~��7-K�Vt܇Q�>S��.<N`�<��k>p�0^�v�t����������V�Lq���z�q�TͲ��w�y-�~�i9��B)L�x3E@Dz�,�^�{�wv�W']%�I`x��} �a�{�6��u�ׂC-9w�5jFH�n5$�)�آ�v�
�tr�_��zw+��J��Ft�A�������t�/;�\aC\��*���ol[�.�i�1#CZH/��;�>Q�Ǯ�]�	��إ[~�����$3:32R����"�����`Ą��!����Bq�X�^�{Ґ� "�9Z�`��`��b��b�B݄"���ں�(/n�=���I
�_��;\pW���?��]�dw�@A�����[D.���u}G`I�� ���P��zi/�fM+]D���������AL���#��o%H�F�W�P.�l=��9�2��O~�	�B��S�S�K�1RCx])�ގ$a��*8~�'�i�W�y,r��ꙁ����F�\�wų�x~ض�
&��ɴ~��#9S�0ȓ�Q���a;�i?!����Z*�t�����m���-hg���,K�*~?o�5�R�55hޅ�������QUx_�B���ibq������xŔh>XfՃ"��^�ž.�]�I����C����`Fu�5���É �K�1`m�2^��1g@�VJD�+1�Q�.�` r���-�j�+1�y�#�� ~�T�2�Z�A9q�Y�$_B \�,��c�Û��l�;o法ͷ)�OQ�'�}�q44F0�w\F¤J��r55�Rw�\�T5^!$yZ6��i���ZJ�!���?y����-�In�;@nrh��_�]H*"�_�����[@'�����Ŵ㕁]h�qh�笑M?��cL�^��/�c=���[�������H�cP�{$�	[���N�P��t�������oņ,�s8�C�v�7%\A�Ό������2֖?#�;�{E����D��q[�ţ$vx\i&<�4����(}$��͛�/k�|f���&�`i���n���f2�a@c����Lџ���oٴ�?���c۲GJK��X�QQ�������DIe��-A�=I� �g���x�:�y�`��w���.B��&�
7�*0����(�R��62�SLWH���U��:
��L�����ǲ͠�$%ބI>c�Ks��RC�F��G+�������E3�˜ߵ�� ���F&C�G���OQ*�љ��4��G���+S�Mq"��\g,b�h	^\���ɚRK��S���pQ31��Q�zU��X��[��]�3����l{CMTp�+�"2�|�s �I��r��!A	G�H���x�f� ;2N��[C���.����H�ȒsDG�r�5�;�����|Jyq�[�u�[�U������2x�;DXv�G�p��fY�}�Y���LE��43�+5qF���J����\.�Ff�����<�yZ:i���r�j��`n�����_G9��8�O��L����h�K� ����f�4u�m���C�g�,���W���Z�Bq24��B44Oǖ���M���L/�ʡ���g!ժ�NcV�EF��,�hF�ȣ"G�$"^9���t���z�ό7�B�A׸E!��̷�]���\�\q����{p�|q9}���]�Vg��SC%~]�jt���S������5�d�����|dSZ`b�^�����'5��y��TN"&��'�q9) �Z��|�@=�՗��_��V�4��_�<ʟ��0���,�QL�:�,C4K5�7�)���*�� �E)�/�H���S<Stf^��f*�J�ew��te�� Qf9�8gZ�L>�a�HF�B��#X&N��;�޾-�KKsoLUZ���}�!8\�E�$�Ϙ�&*���*w�*KvtQ[��g^d�F�,ùp-t����vPk]�8��NF�t\ڀ�Y����%pΉ�m�5��j&v4
�IW���ܚ���a��,�77%2�����}c�"�	w���̵�5צ���<�$�Sv$��s��WQK4���&����6L����Rɼ�ct�t���s_y��.�ۦ�]>��@�U�G�� 	x�v����r��||=��EE^L�VW3>)�`��`�"��T!G�@���[Ƙ�����:�D�&t�e|�C�������
m��бe@���FV�T�r������OO|�y@ZM{�����["�����Z�T���ϲ��	�s�
��3�b�m�J�c�i���y��1�Î��5�%G���h4h����9�9\y�L��9��(�C��Jn��CJ��������Ʉ�)`��>Ǯ��W�����<��/��r��q�a<�rQY|^kJC[o���*�N�f.<����v�K�͎4��N/l�i{��aM��m0��vճ8%��AT�mJKLb}[��D��ޮ�����9�0�S'���lH��+/������ŲJF���*�Y��iF����X�v�3<l�ʢE�l��nj��o��U/���e��g����6/�"�S9��l������"���iN�}_Qt�#���#}��
�^�\�B���`�]��7_��@��$�������i}{v9�k�@c.U��1K�	��+��QD�M:@�&0�=���Tَ�C�c� ų��{o���q�q�����۲� ˍ�ǈH�f�55ף��R���i^K��Wk��a<�W�U��ؽQt܏��˞�%��D��8�^���.�s�U�1���|p �Z"g\���KE�(� !5�r�9s5��7��|�W��w���jSat�1_a�Or�x��f������U�G8)���G����hx�V�#	���ܽ�ޙN>���yċ�,�!���7
|i�E���[�!���1�ZVwy�iXV�K>0,���Տ�+��,Ԣ{��Ru�=�s{1~9��̸��33�߈^Z����}E9�d�CG�
�0�x��
`�B��(a�O��
4���@��X�f�B�]+E��)��Jl�+$z����y!c�wA�����ȘU�F�E��f��X�e��9�,n_	3ݐ(����,����!
"}�Q�@%#̎��Ǵ��8�IKO4D<�>��@��ս�`�7[~n?L2�Q��x{������\7Hp֛������.�Uѹs�D���	�<���\}���;���K��in]
��W��tw��4�讁�~�xŖ�{�]	�dθ��mIg���H���]�2����6
�_��J�up��DT؍�Ջ��J�i��� �2��H^�d��� �8�o�"j�"oRlFѽ6s�E�Ř���C�h��Ț��Cn��E�'nČf=ðJ�.��g;���L�`)���o8���EuɈ�<S�zx̳��:wr3��+�����A�(-o����;����|�hV��Yi��7�ݘ�Fr���`��|p�>����Cs�ED��sxYy����Ld�J��b�踠9c{A��A�V��&Et-f|��0��	k�)���K̼��j��V���s�@���#z���O ��MӲ����<�����V�z����T�y�e����lѮ��F�]�1O�?Yoߕ���Ń����Q����S�����;��f�2@@*��%�`��kM?%���[�V%����jit��Έ�Aji�6e��.+:$(>vY����8�C�q<$�#&��>�搿���EW�Q�<`��?�s���B'ɞ1z�%�R����p@ܤ��*
�p[ƛ/�rKJ���k�86��yh{u4(���q�R�Lswy���G��DC����_<��� ǣ||�E�'4�T5gtش��5}d[���e��M�n.����`������fs6��	�����J��Z`O��Fh���v�J�+|�F5u�T&K(#�y�d����E7U�@����}IG�q�T�L�|��|]� ՘����4���f+Ŏ�z;{����$��e�A�&.����WhJ��"-�%ٳ1C�[{2�P�ߺ�p�d��JЬ6���0�����O���P�I� 3_�o��������W��\�����H��l�/��K���`�$߅[qN�$�A�`��,�3$�X���_�3����]�����s�d�/F���������z��I����4A�h7�Ю_���Rʹ�#��9��JF��%&(rNas[*�����p��o]�c�7hh��4.�B�vW�c#�<B��_b�;������������|A0���H�ב������^kv%�[�'
͜�
C֨�ܻ�̰H��K �PgD����a���'z`�L�C���ѝ`��\����E��k�o���z"�٥p�Z�v�pZ�$q��gf-�c�d/ ��,<8��x��6V�N�S`�R�W�j�����ck� ��$^>���{D��I�k�k0?�Q��)��oV����i|����Y��R��x��Rs���R���4�J]�5� �;�q!A����t�9U��v)9]��$ZU ��E��C'��2}{����7z3��\�1�	rd!\�_{��X>&^��y0*n�+�b��.�O#g���c��ٿ�C�h�=�Ό�P��J�`"z��/�C8&�>p�$e�C@DR+�W��(�0�4��A0Bq�`�w��C 5MLy��$�hf#��� �M��i��Eyd���fP�ċFI�g���[�%�p�������w�Tx����t92�p^N�7~�*��A��7#+Q'Ɵ=(��^p�,b�n 3��T�t	I�Y+9w/�M��X�C!K[oq��-zG���=<�^ȒΈ/K��6��R�X���7�#U��d��.��T�ɀ��#47�Q�A����?Dx�Ќ�̉��i.��4���5����=M��Żl��@���by���p���LkH~:��ߵ�+��M���$ �:b���F8
��0 �`_\|k���K���u�����'��UH�Ъ��'d���!���G3sn�0�%}m'S$<��p�3��F֍���D�H��=�~��=�IXZD��;cϝ7��Ð�q����X'�dzGϸ"�7L�_BFH�^a�U��%�h���A=�;͘[�B>\�Z�}�:���\���'���[��4ܒ������ ���9�*�Kb�牢�,�0�g�����uc�A�V����Ȋ�X���>t��Eߴ�� 1��q*��Q�DQ��
�����$�n�"� v"r�%������ҋT��k��*þ��!���+�eH՗®G%�L�K�|2S%��F���d��F�%�(_q��T ��z0F��iN�@2-%��3$.�h���,��S���?g��	�����,<������,�o��b��w�^J���~���PKi-��J��)b�g��D�T�s̍>`]�I���u��:�SQ?��)R	�,���R� ���ѧx�m;��spݔjE�V�A��w����?���l����#;��w�q����	�{��q���98�u'�� !l����5��y�T��r�Q����C� s=ו�uӌE��.i����'�y �i�K�@�k�+xV�v��8ӌ�QF/&�m��ۈ�IT�p�!SD<ߞ�&�y�:���v�0�'��c���Y��
/������~4"r��|*VQ
MQ1 u���x~k;��<�1��%`�fcs��A���d4X�'�"�{2y��\��a6�]׿�;�m6�(	����/D�<z&�fRW�V��|f#��:����������&���C8�U[�Vl�=c�$94$����+�}��Y1�RQ���Ghܩ�mۖZ��t�aʕ��;�|���b^ڲ�e+o���Ǡl����y����r�{�BEB���흶��N��v%7>�
��F�:�ѣ��S6ȭ�Ǎ�SiY�� D��'n;
��}��G۫��'I�W~E�A�jcU�L�[-<�rH���k6��P�r`���[�WNC��f���T�	����m���4{��4�aK9������l\��{�Y�c�[���E �*�5ϐ>L穭�] ��LZ+�thJ�����_;T+��V4R�LO��d�9�����l�����p6�Ts�h�MҴ�и g�����u��煆�j��}r#|��"��ĸ��d$U\����l�8��d��ð�7�װ�Hn�e��z`ˁ|�T0��<�p���sצ�t��L��h����-��
�Xٶ6�I�*�R���g�K�6��9	�T[�Z���l]���<�[=��QB�"��?��]7'�E�Af���=�z�c,�GZ�DQ�Cl��bo���R�aγg� df9vi����W���'�AK6�����LP�Q��	��^hWNh��li���\����_4
k'�Y8����rTx�;�7������!o��[���(E�K�9�c���Ԡ�~\�q��fPWY9y�R��7���^̖�X��hdhy�T�)�o���\l�/����A����I��L��!��=V�U�� ���j*䳁��Q
��ǀ��XU�lO�_���<�°2�qv�L����G�EL���I
��zN���@�#6Z j(lVc�5��d��Ԭ��B��
l��e�&���k�|9o�̢�"J��(�'����Ϗ ƪ��R=胍Q��g����X��T%Q����g��	:�t�͂$��p�>0�ۄ�7"Z�+��`"i Qe�A� 2�=R����?�ٔ��J}b֍�
6TZ���{�7��8~p&=�j�8���E7f`r� Tɯ9R���d�=��B����#[ڳ�Pq\�ԅա��P$>ֳ�@�]�b�+�:��d��0,ؕ�h�u�`�Nh�%7� [����wA�C|���fJ��)GP�ǄW�p�9�M�QR�J��2�R�A#�_�7�h�q�J��y~���K4�[{;[�%}�W��39A�&�Q.�ء�����:��韔-(u�'
�O�F�ǤUu)˙TK=�V�����Ŋ*'dTůޥ2#;. �Oz�=����ҳ����4�!�4�	��~�E�����L�I���n~��Ѕ�=Bݖ���T-x����I*=v�cY�)Ƀ�HD�G��U����t<O�x��D�+���z��{/tr��j�I��ivD������.��ڡп�&�?B1���^�Y .�,�?F� ��6�>�D��i=�g��ׇ�'�e���[g�-��T��C��o��[R:ྱ�u�0����+�!���0�I��_@�DT��Z�K.���{r[�"A�b����p��:���_�k�?
+�l�i�;�
�:n� �'�>�i�
g�p?��+ma�5A�/91�&a7[�)�����@0?�d_�2b,��b���{Iv	7��M�����$��R7��k�����uE&��Z �ϡ;y�=ǝd�7ƒby�5t��)!H��&�F1��Q�Э�l8z��x^�/}�T�KUʻ��)�����4X#0�J1:2�
-��=�z���1�����pE�����F ����z����uP�J�I�e�qCG,28���r��77�%�Nó?!���ū��kb���ˉI��D���{~=�/ር��Ұ;K�.$j���E�@�
�iqgyN����-�z�FC���NR�'?���}��^&�j(��Ο��(�o*:��I�Ԉ��ә���~��w���Ǎbk��*�!�S� ���[�X��!7y#��W}!�����_�����n�Y]�D���Xn��\���3ޢ������׀UH;C
F'Y Jj�B���!�MU7c�jJ�g��z�n��F����h�Q�@���=f%.I��T����]~�9�Q�.S+i�l�%�műO��Pr]�IeNuReF�t�W��!ӣ���^M�Hz�w�s��J��!�"�6.~G@)��O�G�:���}O�{U� �=�ޣ���3�:�����7(���Y�P�����;�����qp���;D������l�+�`u�/�Es{��㙦�x�LI�,J<}��r�f��);SL����d��I?1:C�vB(q�Ce��`jo���b]��1�M�����-;��a����dJ�C����Q����	PB\b}g%	���pC'���'�zB��`J��A���_�}R�ji_8yz�o�BL{��|�A~�Mԓ��mF֤�<2����da#Y�_�l��fJ\�����Svc|-�}��Y��o�����ė���i(z�E��
`~ގn�)�;���Q�?��hA'�F���(eó`��v��w�{NpˀDX�6�_�5?���.eU1=�lM�� �w��$u���_���9�Z�o6��X(�6�F�H�	�<Q�� �1��W����:�������k�u�qc�kV��F���J6Ay1�5��/A�7�f���͹���t4�p 1;�P�r� ��}�����.�/o���#W�������FK�?,QB��J�l��b����V�%�LH�7�N�N
cT��&F]7ټ[��I&
:�9��@,(���Ǆ����[,��o���U�c}�۾µ��
M�0��R�l�����d~`8��9N"�d�'������j�f&�E7 z���,F&��C`�����ߋ��F2��Q=?�Pl�z����,LwB��T�FD�>��Z}3�OY4��^O@�b���b�������~Ϗ1�E}�-�Ma���a�,�J�td*��ߩk����&U����1N=W��Y4#<=����;�\.�P���\�`��%"4��ɯ�����ZF"�E�O��fn�U��H�݅���A��v�z%e0{ŵ�Ҵ�Bٸ+U���u�N���VkP�Y�S�o�]Y�����w�P��P׫��L���=�a��ڣv��N��bg��hA�����r���p���ޅn�ȇ/����\3�ߌ�Ѣ�l�%*��m�5��O}�/��x��y��W�%�!(vVɡm���c O��r
�Ȟ�IQ�'揸X\ �	[�a��7Мoz� �Ѣ�L��_��3H_
�C|����*y����";�.�F�˔բ;�c�;m�&���uk���@�R��=��=�)��N�eIeVv���x��-�C�J�޵o_:U�c'w�E8��|�v���R���!�4�D.9ǝ0���WB�ɆJ�v��<6T�/��~=�+^FU�j!"\]d��v0�q�A��yP7�ܗO#��@��c�<����V�2���~VD�όRE��~jwi]�:|���(��IRŀi�J:�������UD|�}:N8qG��05\�|PvB���N���bpzpn�����0������i�����lF��;�+�-� �>p�BP~f���2��-a�-df)NJJ��0�ó��g�	1����ii��\à28|j���pd�^�l&�"A� ��'=s�E�}0��_< �=3׺0��ڎ��Sl��Ky^|�O"�Y��t�
Z<�S�)�LѢ��h9�d��3V��3�hqв����wP�<{���<�d��4�.�*��=9=7t�S�%3'�J.��,iz���5Q���-�M\N_~v!�L&����̡-�Y�'�����S�Ut1�S�ft�j��
�0%�'�B�ô���ӕ�$~��"���t�M4v�=z���[�0Ը	����N�<~_��arɝy��̵�="æ\`|A�:d���W�a\���DH�4�|�WJ��-�9�P7�k�{k�"_��Y��pV��D8 u`F9`�@D&.�㿹���[_ԯ�%��Zp!G>�T��އ��&|�s�ь((ɵ�i����.⪳an���9&�H��űhc`�p����R���wt3_�'7k;,�%��̈́�߫��p?�g���|� v�ۣ��Ko}ܠ����>~v}���X�0��R���$Di#N��}'������o]��ō����*/�?��<��T|EJ�n
�_g�Y%�X�7E�+ǝ��{�-��qV�5�%������V��0[��Ӽgl�0��V��ل;�+R׋���`�������}'�ɤ�c'c�54B�dh�����8ۛ�t�_t+�2�G]�(?^�X7���Jꑔ�!�rax��L�a�W��K��٨G�zևO|*�f��=FIgc�	��{�F^; �U\��;�V'7y�����]�x�q�T�ߘcs��͐`���rBSV����	 3���J)J�`%�����#��.A�����[�,/�Z�w�cv�B������x�3��>�w��(��ZͮhE������Wa�?y�جY��a����\���-LH�X��E�H�9���}.k�B��q�v�8k��B�ה���r���j�$-6���=i)R�D�R�G�}�j����T���|o�l�w@���铤0�[đ��"q?#�?�r����Ǖ��xd'�E����;Y0?,7�3�q�>A��G	?m7nς����viG��y4y�������gб�-�pC��� 3`Ry��肕�:qe�ܧ��
��T,����? 	?}qt�g��Q�r��D3� W����H ryx|�dz�k��6.~s0��?���ɳeo�����H��v�����r�V��D~}�B������ ��@z�������E��qv@��+� ��ٜ���S=ȫ:���>>��\N&m Q�cn$/0���/�=E3�ZN1��G���E�R��'���4)i�>�e���
Y��txI��'Ʀ�����J�t�H����AL��Ӈ�5��PV!���:Hsv�ǖ��R'f�:?]=�E@�$�
Q��|P	�K|�
�5���R}'*gB5�$�n
r�M45C�xp����"P��_�=t�^�G �%G�H�A����ނ��z�0��ը��>�O�ۈ��qw"�rQk�Ъ�|��f�nN�x,ϽCO�Gkg�L-�*���"j�C(%��E�_���ek1���e���6���iL�@k�w�������e�!�A�.e@n5A���T�+9lb���G��67}	���Z����V�M"�ۍ嶠$��Fy�ƌKE���Z/%�����3��ϧcI��aŤ ��0��6����so�;3J�E�\n�tI����цc�cJ��Cwh�^�A��5�7���65Iz3�E�ȱl<�ׯ�n���5׾��\�}�<J&=�k��0D�|�t!��歈����}��VQ�Z̝�I�._y��?�c�6�7���N?�$T��{W���t�A�ET�o��\�Nع���98�4���G���(C`��,B��t����R-6��Dq�%�ͻ�1��G�0Q��R(�ɞrD?߬n+7z�z���0}��f����Dz���>�H�3G�"!�VN-���$z�/aQ'^(#��S���/������Q,h,i�C	�c�*c4��.�H�z'A�7Z�gz��>���+Q�(��s���Lo��,A�(�s�mq��a�h��5#�_E޹����bNR�J�/F��7�T,�u4y�~'�e����IK�-�M���{�,��g�|:=��F{߱��;)���"���\�^FE�c�R�ȊǞ�e�N�����q�E��UA�W�����z �2����|��s�2g�j����;#U�B ��Α��v
�ȕ����5S���D =p؝�]	���}Ǫ%x{V�3_�ڲ�3�=�u"> Ŋ�P[?��hY,]�߼�f`*R�O�V�e��A�PN���8��*d�_�2��N�.�B<q~�ذ6��S�N���������1<�!��gH�ۮ�
��������[K).\.ݦ|��m�{��#yl�+D߯B!\�AW^���z�5��WY�֥>�O��V��&��n��p�E�G:ͶTnu|��#�����<����GI��75C3��"��0S:�6�0,0���D
_z]���N�2�tV��Z�8:�����{O�9���Yupr��8ӏ��� �(q�Լo�9͵m�f{�0&��b����t�8M����*�������m9���rq� c��:�D����@3�dҜ*�S�(��89�봔z�-l�z�4&�{n�W�R�.�G���D�%�~c=s��8 �"-�:sи6O��WD�qev��� qr7����Iy�J����mŭwE�L�������S�=Z#�ֻ{|=��t��$�FӶ����b��Ȏ3�����#��5SëXi�|L-"�+���)=rqF��W���?'�	�pSL�����aK������>��O�'�f���K}�=&���~\��]�� �+I���9<��X�a��Hf����u�T?�F.�Ѽ���EY�;�O*��õ+�F��y�	�h��rU��k�b�B���)	)}��-�a�\����)�koqf�.�Fv���������o�m��eJe���O�N��QV�d�M��V��M�;9cޙ��cNe���oo!8�K�q���L,�5x�8Ŵ��|��<Mm�$\�#U��X^*NA�2�g��^�[q�Եq�i÷<[KRx'�����6B!A �<�|#�Ϫz���Ȧ�;�kWz.�V19��l��G����' :N)OK���b&k���mDQ��[s4x�m�#q���#j�-�� K����D���%#�V�^%2����@s㓧,5��m�D?�`2� �Ω9��ic���j�ejzU�}ہ������,Ί�@�*q
(�iQ��~�ص6�������|�t��_.�1���s[�F-]����o���9�W�j��=[u���vTN+�Y��l��{+对&�����E���n����v��c9���)
��҆����k�Ekj:]�m�36F�^di[ �qm��ʀzk?{M�e�K~�~(u͘^$m�FG�=��V4�.n�'1���?�y|.�@�a� %��$;��$���x����~3`��ȗ4�!%6B[5.|�M��ś��:4m���E5`��������.�@�5q"�o�����	<s��)WɴaM������������3��J͵c��}�2ϋ�e|��p���6M'Ec�(Ns�L�ǩ�\��b=��~/�2��\XP��@�d���H?�m�9��C/b���>�� v�j�����������\@H�@l��ې��	�@��B��X�ADj�'���clf���Ԫ��	�M�С��# �4T"v�=�i�,�v��p�`c�r˧���_p�Ѓ��;�Hx2!�YQ�;+!W�2�Sem�#��LeC�Z�W��E3X.�2_���M`�lVie_�6bw�x��6T%��ĩ�u�낯���WW��i�����J���P��i丗��4m�`���7އ�� 3�6���*���t��*_J�˘:{`d�r`�ڞ���)%��s^�zz���%�K8}���:m��� �ZT��dMX�Ko��}Jy�ԢГ�!/��V�ě�q_�n�ڤ����X@���1��Z���N����z�ֵ��`_�"^��K�%�S��\�4��jN���l�km���ޕIG2@J�v[[W��w�&�����/#�x'�unH�6D
6�P�TAm�
�%`D��t�W��8���VT�kQ�׺����e����p��� �=�2(<X��LĮ�@[�A���ـ?��> n2��b[`�=��(�Sap�ó�ke��ٶ�����skcA��Ib�ވ�C��1��s8a���)��-�0��O5j*����sQB��jܽ�������TZ��������fߗ�:�7v;�8u�ҙ�9G/�4��;�	�����W'[3ۯ)�˱���W`�i��nI	i9�T��]א�����z̖}�+�a���:*��}:�����_CG�h�%-��j��;"������v�k��0�7K�%��(�E�����^;_灞4IW����)u�^���W0V�.u/��oC���Tt]�����#�^����X@W$�}�zѪGK�^kPp�Y6�;
A�A:�N�5���R��P�V1�;�6|�i/G�ߞ��>�<06Z�#��b�g�(.�DbЩg�&�K�4ֽ	qb�:�! �O8��vE���ԉ�>玧8�P���T�����X`Ew�
v�|TP<!ǈE^5O���Q�DD�e~����:J�=���k����H1���Km�KJ�~�����%���%�������kB`�,N樊��u�����&}�nߣ��W�b�!׬�WҲM�SVS
�<:��C��r��lao�Dx���{�3<���fTO��OVo>KI�{T�o�NJg�vw��צ�h���GQ�uM�/63EJ
�`g-4���4 ��<F���+��I���J�M�X��l�SJx����&j�����_�R�$]{%-ڿD��_.��F΀��~��b������L@7'9)^!b~Լ�$��
Uߢ��6{:q�M�h��[�*�K��0��}9�2u�ڮ�Z|5�w��Oe�f)��X��1*����l�YArA.Z��B�r�#w�:�W� W�;N7�v�m�9h��zд���:�7
(�'�R{���b�4g樵C��~�0)䧻SjQ<�$���7=Y2;���F*����`�:�LZV'FT���+�ld7B:�5�s*2��b����#܌����(يB�l�9f◳E�@�g����J����Z@��(��Ѭ����$;�\�׆IiȯU����7#�#hz`�v��T����͓ŕ�$[��(w:|:�c~�gsg{�Hv�q6�%��=�W;'�|�a�'4��!��ㄈSe&�4h�a$��Y��ND#��|-����Jh�h�)3�h��ڌ-�]���+H�7�P~jk�W�T-Ħ��
�E �iz���ņ
����W�wXWP����D5f�a��>��O�:3?��A�~|��$��U�^��m:����/�\>Eu��!����&�W��aEе��i��5��PD��ƿ��G8��q��t{ �!.����֚(�����}I���764���X�I� �K�e'g��|����YMل��Ep��v�g���������� ?����-vp�0�o��=w��T���u7?���ƥ0%��6�I����->�#�
 �r���=/�uyd@�� �uvbPv��.%��kN]��r2Ef�w
K��)c�<�g�GΠ�ƺ�k�j�`����g#!ڎ���
���<��	MC�%8��|*�bg�>q�ä��y��#~��z��܍�����a�d�j�7��
�4��B���d i����5�����U���D�	qM����¿d���>���4���׻�ٔf��H[��E������w�o}�:��� �lceآ�h����iX*=���#2t�AT{��!��L=�đ�8b���zy�!u	˓0^��N��թ u��̍Ì��x#������@����Q�����4b���k�`s��U�E�AQ:Zʎ60��xS2ƥ���֯(�K��=Ҭm���Jۊ3<�WH88{Q�N ���?o$�󐖙SnǘyK:�ZY��mk?g����t���"�yL=��c�A��|������a?�?���?��'W�mg�o>莆Q�����.n[�0<�j��4��� �)k2Z��#�<>�ӛW�_�~��iT+�����=��q�;��
��
���\�.��v�lI�}�M�����c�׽�9q@����P���<dVӜQ�z�8����p�0�Y��܈�V��2'N�F��lb���CYb/L	�/�tƌ�{zgph���[��m}��V1�@&K��,;,5���[ݟ 8�d�H:��V�����H�U:�ȄUM.Z�V��п67�(�Z����n93H�)?ܼS\��H�`�{$.� 7t�ﳔM�M�}��nL+������\���U�LR�Ի�Z����g!��M����L9��sg�3԰-����|Z�m�\��,�a�\A�Ĳ_*|h@JL��c��U��U"�Q�s�˞�aU����:	m��q���y%�w�.}z'{��*B�Ǳ�C$��1�`/cRԩ�׊c*En�ر���^��2�[.��ҟ�
�091Y���QQ�Y�P�[C�|sN$��.Rqc�gil|�@����J�5�E�u�o�/���؊8�HYL��e���V"�k�G6��P6����a�&��V˫���t��1��"b�m�#����q���z�L�/�JB�,O�5�@�6���	0��5�JB� ��̼��V�<GY��"	��sR5) �Db��d�>p��h�""Յ?��^.��t���}Vͻ��H�	퇆(�&��&�w�0~4g"f�	�$	0�țȸP�E>��k�$%��H�~��p�sӚ�Z3����@=�/���7����d�� (+òZ $1J��\����z��Mwɴ����*�VK��D��!���z �UB��r��D�ւ��,"�FGz�O���G�)y㇢�ȋ�J�kn^��T�M;����,nv��}��w ����5����rB����,$�J�l��������'�[#R� }j���u�1���Pw�� R�GD4O��{Ҍ�P#i�Qj��r�/��wrXK��,���]<��c����uSo��AZ���oU��x��E���y�i��X�����(ش/�����
���Hy�ƒ�3���g���O{�xYM��V�i� 	�@�-����.�յ��uA�!5�E�V-���!����@�3Zp�݀��Ί�Fg����I�����|Rƶ_��)ѽ������� Qfh"m��:�\WD!}��`���|ʝ�����!�x�:�d�(��/�O�t�|�}!5c�8]��+��.aգzq����7��ZD�즢O�P���?\WޮC�%�C�pH.�J��A.,z�OoV�������wB� x{�R��*��0U��~ ?���D09U۳��5��'�Ԣ³]Ыm�gO�b��Lk�?���)���^D���D?;YWcV�!��'3� �8B�wW3�Aѯ$F�/��_η,�䞔��%`�%�u�8<r2%8����E�i
�����HD�/)ذ*�B��Zﷰ@�������� �����!��sQ��H������k9�fQ1Z�i�}P�eL�� D�^DQ��������j��<�����{�D^�<�ԉ��d@b7zG�&2��;�@^��p��n�@!6��$�����$e�ݠ#4
�߷����CG_�}<�4 ���~�c��W㡠��k�ݍ�;&�椉�v��t�O�s�d��xo;܋Zw�ЂQ�4�����"s������C�1wnb��}_4T�;Qł�1++�o ��$!�$��s���4���+����Q/��!��xKC�E�p̀���J\��na����}F��?v�S-li���!2f����2��xMM"- �D1���(�l�w�ȣ|�=�{�'�#�M�T2׼����e$U��dU��淌$��Z��u$/�zW��_A����Q�-��穲�;�����w�?:t��}�9M%?�Y�#�?z��<G��7M*� /��|�}h8vѷ!ˁօ�Ք+?�Fضu뵪x��H����
k�^
K~���K;N�-�T�Z�Uu���UCQ�'���Ƅ��ց?�"T���z:�+mKPo���q9�;�2���(���t�)p������B|f��]����t�|�g�9&z�eh��%���o�W���Қ6ccλ�F|H�G
5�~����]B�7_8������M��(��GYJ�P��-��g���{����z^�X���0`O�Vr�>!S;�F|4�O��	 >��<�����w�ǉ�F˵�3h�7&�|C:�e�q���X��&��\ZsLD��i�n���xj���A4	�>5� ����=�߹k� �<8xOa�X�qf܏C����`R���}�
Y�?i)�6h0�M��ΐ�i��eh�vg��O}�=�M$⫁�*%�"�9�(L���h�ݧ'�˓^�f�L9��S���^� iff�{��WM�x��^�\.i���w���2����?�%_�\�.���2�O���k�ڐv'*�ؔ�`������d;��?��3�q�P�K���n���Jw"C���¥Bb|p*�`a8w�*���\ϣ��6��sᓗ�gfQh���e2��8��D�z�|k' �yѪi�9��-5���`�ݢ���b�;���Ռ�z�l��D�H�Չ��A� ���F�u
˞	�Α��Q&��c����M�4g����j����/���\�-"m�#%g;�{Y+3W0���i����O�rl��M���_�^�	'�p���?��)�_M��c�u�>h^������Et�	Q��@�`T�Ё$�."��`/W���x!��2��hJ�D�z�Z~�q���(��x���-��,Ҋ*�W����������a���w�"A���j������<n*�<��m�ŧ��.Uo�R�>�9�ҿ�,�f�������N��w��ڇ�[�y����%��Y���S����#����_l�}.d��3��칊/���m�-K��)��2�^��ׄ/�ji����|�t3��w��lﭡ?�)~H��[���/�q��.�>�1����~�,*�N'0x��<EŃD�]��{)��(=��:L��h<�"�/ W	�β�����>58�0r�ۮxws	>3��W���E��*G���v����1�s�'1������{Y�C��w��וF�y&uOj��(k���=~�ݝ&\X5-@�[x0"ܶZ��3\�ǀ��i\��T~���$�`%��{�!١Ҏޅ�+��ˮ$뮣����;ў�A�T��tu��
`�((��4��:�l���M�"�|�v:LW;�ɹ����:���wV�����T��]
�b�L��BZ�dC�(&(.ˢ�w���t+�0Og�����R���L������ݜ�|�S�vcӦ�A��7l�K��8�&��O+@hT֏7��=��U�=!-(\�}�+�v[��9�������^��F�����s��V�VW�,G���}ƵҌ;~a��;��K�"��}�P`��q7�����G����"c&о�5���A��ר�n��f��[��U�.�XY���u�_�t�&M�x���I��fEl����?��.��e�����j*��o�����v�}b�fUD��d�
[�">ܯ��07 ��;��x�����xW�_�U^��>�����7������ǌO�c2��
�1�b�{��kż��^�4hP'Jd�'�y�WgomW5��a�/���{V*��f�"!�������r��c+�j���C��_C���Sl�vv�n��=��殰�j��P_6����x� ��)f|��Do�l�(q����-��D�&�)IB%���Pn�W��x�C���b��˄u��IQ�� b�����>B���F;1~��!�K���F��9k�D�L �"	Q�9�n�I���x�1.�E35����7�j{���������b�4�GQ	��"�ʽ��|2G1s�J�m���\P#ׂ�-�����m�A��[��W�`�o¼�N[���t��5-S�^y�+%41��;�ʼ����F��N��9 VQDK�5������+}���'��AB�|&9A�~�L�{J��P�~��e68�D��͙-�T�_{�um�!�/�m�:� �fg��8�;�Or�i�(&��n���x�<��� .NH�/��=S�="��P�j$���U�ki�|�[ʐH��~����=W"&�0	����tg�	��n��UqH���G)��?X��O7����FR;fq��	WReY=��V�`�r/�`�X;?�(G�FTv
� `Y�P��6�,m�uLʖ��<�kyn�����*���^zh��>pyυ��yúZ0y�[� H��y�C�W_��m�qn7�ht�{ɍRbݧ���xjI�-�9l^dV�iȦ����I��+G$�����#��Y�#����*�r�w�H��I��i��~Q�s�v!����
�I��4�}ݵKSM��c�����]����oG�_;�(��?1A�	b�Od�\.;�ܬ?�'��� ���dQ.:�۬�IY��>d��������@�Dιn��*���,v�3��Ӎ���$���?�9T���l+9�,�Ղa"�^�Y�߶�PA�L̘�e�\1r��oڟ�}F�%n�R�E8`��d�hy��U���6q��ݫH���Yb������\2��ڳ��܏�t],���ԝ̣.zdn�C���G��Ǆٸ��N�S��&�E(a7�L��qHJɾ���!��!$��P�|a�5__!Oe6"��iN6��:�@���;��%���,�t9��7Ą	D��-�;�Ǚ@Fo���y�˷r�a	U����m�?�����Fʮ���|Cb6�W4��ރ�	*U�w�
Cy��x��u�s�Z����*�Ek�Y����B�g��"�hMa����!hMJ�.�#�x�ks�6a�v;�c��}O%a�>�p��\�t�,ʽ��R�^ct�c��8y}�9m�{{�J}w�<Q"'�zr��L}�*W2	��e�+�aЦ36}��%�H]@c%��h�z��0�M�ɜ���z�c/?��J���W5\�q[_��4��]�$'0�%����b�,!jX!����f���`��x*��G��U�`h⍴Y"���&"��e�ފ�R��>S�/1��t��� �Tn�����6�GūL�S�u؞ֶ�h��k�Q"�K������{��QH(��`Ŵ����c4��\�L��%'���>�BY�.�W����Ȟv�D���qn*j��9*�7h�;A>�>�;۳f0I��S��`��u@���X>�!�ĝ��:б��"3hn\,3w��WF��tM�Z�y0�G�����E�?8ڙ�8!S�?9r���+�uj�6�ԩ���v�����)�I��j���S�@	�F��S9�|�t�|�U��/��nO\��,��e��LE��z3�O�*�f �[�M���oGyffO'r�:�ό� n���?�ը�	m���fo`�	g�� �!n�8u:Ti4��a��&�>���!FO�e�OQ9��u��Wq�|e��PCdJY��U�.��k�-8Aw?c��©\^2��g.f��%7Y�@K�Jd�j����h� }9�/�魅$���l-�xf`�Y*�����Ѣ�5��lg��ʹ�=@h�&�kVٌ�=��-�ܣ��f�p`I��U�2M/id~i|ň�n
���"V��p9�(��;�o	�I����R�H���H�Q���A���a����#��J��_��֌C�:/�K�=u�`^鄱(dA��9,��~���x+����obi7ҧ��'��}�X>����Q޳�d��$�6���<�����)g�ǆ6d<]�xZ0a��$0w���p�O��ΗxA�ȇD��s��S�yM�3�+$�����h�k�z�x��5R!we�ȉ�N2F.w��ޠ8���U�%����[U	�
#�Ts�X�~���V0�����/�$�_��)�S�A�JՊ���8#�e�$�t����{W�*(*L(�� �去�5�n�b�w�O���D�*������u�EfA�@�'"�ws��
%2�ЃHbc��H���!�%b� �~�U2�H���*}�j�������~%� �.q�wM��O���tU��A�2}��N N4��̸E�v�4:�x�!��/~d�E�9���z͕ǒۭ��sV(X�.��|�Sw�P���J%?�ꁸ�P-��E�Q�+�>��<�g�r��D%�c���xw�DF�߈�{�K�'p]�ǝ�K0E��O��K�BuL�`�vc���[�͂�C^,&(U׈V��_2��e�ח�qN5�TT߽������$�4��w��x`��k����x6#��7��_q�-��_�а��ILA��~ޘ����5:��q�=	tQ��ro:4�	h��DEm4z'����_����0fE+�M�2��	7,6�t��i~���I�O�G^v�I��M6_����������xlMtu�m�v=�E�ա��xi\�������Dr�@��K��E� ���n �.�s��ԡ��jt�0�m�Y��g|o��K�ҁ��c����>�����?��i5���3��Q�?M��47C͜QÉktsΔ�MW�OX���cI"/od8p���x4�Hs�/成��"����諻�y��GWd�\;����d�Do��*Wo���i>�ז=�������<�x���j�)�nÜd{�#���\�+ӳV�&x�m����Z^���u��}�ߩ��i��5�qQ3`��1�j*��ޣ%������ȹjz,YQh��-e1�\��U�T�Q,���p� ˣV��4oKPP�WѸ*���C]���dsS�qC�e6P�J�Z�}�남���n{�U�cXo���I"���U+�hHK(=�u�V<�;[��wg��>�\�ꖫ0I��u@u�fɀ�|�B��i�x�Ԛ{I���2+xF�M�}i�$)_�h�,QX0*��bZ��:2�j�v��(w��h�9�R������6�v��������3���i�GIz������_n"���]����\8�-ɬ���6d<Y������+#��15�l1����{�`���㊞c��$���})^ ���%�<L܃n���CdQC��W+�j�G���%s e�0�w��+�)'DpR@D��Y���]������q֎��%��{��'`È�C�H6+���A���4?f��Yu���D�{�r��Kb�ɰ	3I^�������/s\������|��2l*,EpW��#]Ȑ&s)������!$5:LdS�z{l�O�;���E�z���*}�Ua��P�;ș�_�����LԺ�x4�TP�:����p��Z�fR- �G��O	*�X0J"0J()��b}��5'��$�n�yj���"��ke����tw�����"~�ǽG��# V��.����e�.���;�[|n:Sɔ�x��_ ؊�?�x��m�d��dև���'����մz�aw����lQxXZ�f�Ɉ#��Z�&�6T�� J�:�<3�2�� �qmm�0��m>�cN�M.��s�����E�ˣ��2_�Vr�B����� ������`���aw��bm��%�TI��|W�ߛ�6��@=QMԑ"Ӣ?�+-�t�v�v/� yj�pז'2x���uvGǔ��KGUό�j�NNt�f���0�Jd^��DW�?߫T(*�L������n��´��j��Nklmm��𨘮�>Z��8�i� c{61�K{�����Rךt�D��޾Gp�ۅ�X8�p�ˊ��I��уԅ���7�s���f����a�����=�� �f[��p @w�e�ʤ�	��r2� ]�9��TO���ɗP���D��"��}1�Y���=�vD���T6�����n��DY��\��<d)F�ړ��h�ձ=z�V$��	+�s�������A�'Z��0D�����sS�MG)���.�)r��FȊ�s�^���c|�Y���;���s��&����Z�.E4E�%NE��Z���Њ�}�"�pW4�Tl�L{!�g]��w��I��|2<ʑoex���{B׼�wᰈ�~���螏D(��2�Û�'���˰�U3���A[C��)�H+�����# ��u-���,G�M���v��EW7���+�F%-I�}�D����I��>i���N,�	����W�X-���~<���M�o#�-�����8@,��4�\�A�4��"yN�$X���ᕾ�V��~���՘��ӂ�k� ��0osw}|���������ޞ��I��Z�!6iXb�z*�\�R�IyY���n:��{6�ۑhp�ܵw�(@h��}�硳�C�/~j*�*JW�~��t.움 L��|�Q��s��w�����)Hm�x�}�����3M��6}����6Q�E/j ����6MvǴ1�d>����������9,˧��d%Rv4��@��u���9��l��Z��Bm2��̓Ӈ�2�zѕ��������k_:A))蛏S�%�M'���&�Du��7*�f)��13��S�LT<�V]�[sH�(�M�؋d�%`�ʢ��hΩ��%�c��ޘ�Gn�`�{y�<���Ǝ-�jdh2�8���i@-��V ��ؙ�s8(oĭ���>�����'�]���T\�+F�����΍4i��3��(B%����5���`�-_�|�U����D���&6�d>�+� �8�u�YŨ��eo����kI��OǓD�J}JLGݚN_�k=�z�Yv5'���X�\�\B���XKmd��	}�7wn㝥�&�Ch��{���xB��A6��HW�