-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
C0Lxgn5i5/sKdBdEhTGQwIdmImDhCn4v35bAs7AZgR25xVHfYfuhGdWL4RG+A6dc/7b99h89xtjZ
NLJFWBIobhPuGyKjpjMmnRv+Hh7QbYXK8e8w9O9K0VelwY/6BnQgLjbVhm01HnWSWPu5I4Cj0gpX
juux0/vRiWgZPMcXR3BQZTO11+BWR3OKTyU28FVSlN2SBek3Ff9MWr6NshMc3dKi1YXHSvOkD1W+
YrePGzPdMQGNPd4ACEUQHPMvtgPVO5MHn46p4w72GowkPYfgPbNcxiz9UgNXzZmKC2CYAbox9Waw
okSXP4mpvBP/4duUBbrGjgrLq8d2cAyK1NuwPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
emARQvhVZbzxyxj9XbZ1ve4WqeFY+YL2aQ06Ev3TczE3FkHZJjp6Z2anmXf02DMdDA09HmNwZ+mM
ECSchwjpMtqdrX9NodsPLb4bLhi6sW57HbGSNMW/qWWRfjh8ILO7OXO258gHywM4SCx5iLV/TUhn
4MA5Gcuxmlb9jEXkzIge/Uwlaz8+ji+eD2kF/eheetk6J1nCmnlf5dkFt6f4qe83ugbKACupDl+H
xo7vStql2pQl9PK9W69mJck1nImn9QxxXQR+s/EnaBXgZzbFJScP76dYN59myo2PExeXyy0R7SR+
HNog35pSL9CKQUxFvgHwZuCHXzWUg5W0eUbG6TU+/rX40vt+uhYb21F3HUGTI3TUQD77oEyKyI59
NCJqIfUnr6gHMxU7rqaDru4ygYrlDq+3r6xLjddu8R4dGX/HIVZyGzYlFYV79mrJ8A33VV3E+Itl
B6zWRW94a/WN6MevGN1oLh5Ge9i8FO0PBuJuBXj2IaqgofAz5sTBfm/jgW9+k+f33ZoryDiZKC0o
IpCrGkd0LJZ6Ivo6TlLgOuVv/5C81Yr1LMsDe0y1nTnbH99dNDsJDWEJ5fRKTfZV2aB4+A3CEtan
ycmFDoA2okA23ofctK/tdwE0lPq6X+qF8zgrxC0zS/XT+VPsh1dPnQ3Tzm1plnAUmffeo0F+5903
Uj9/TeRX7G1PNPZXgPVcdamMJQOGFMWKA/KYfq9I95DcD1C0jhrNY31LZgEk2DwdnaIsmQg50qEm
k6jsnUr61JXSFf89NBLNPgdQDFqyAFoUzKj9qWdqE6Mq0nmyfKY9fTxsdi+CyzIs5LeQcK16cfPC
ed0CrtbKGWIvsXhRTDWfPPhyK45SDsFaqHaUwApivuBdoiZj+mOQC1EtygD8z2ArhFtf6nkb8lPH
GoTRHT9oKPSd20GY3qgGFJbUI5WcuJr0ez1UDfMR2Z2g3DHE7qDP27uyCUvOiM8NNXKf2/dvp+7/
V34nj38pDJZnUIiORYROdBrqi7kIDqQlnayhfRo3h0gnM3DRzFcL/y4lGGHzJuYSeRFEkPI2+TVd
rkXKal98/QwvVma0l3BRg1s6TKrJTME/xRvFEXks9MtVFL2+BbqjBwUOHjeNDpi6pO32GC1g4ATZ
KQqJBg88ve1dyNZK5iD/gfz8u3uCOYLJ1fFF/ZLBWSOHx7spxGlQwgzy0DjTmgiUUSyZHBtSL9E9
1pMc0vsqxWMUA/BKLn6ySaWbphN7+MfYRb5YMGgwe6lO9JY/yY4fgeRQRQAcYB64FakU4tbOlT2q
aBptuX0PY+v16nXL4du/0N/YPk96jsFGTbfJj1SCm8GarZgEcnxBnKEgR9RCSHMj4mO0lRrZm4pB
9l8FEuc5KCvqT2GvUoVs+mBllF3lHVGTMHZF5ZvJHx9RZU/1eoRBggs9nG8yxYNSYgvwofKpDyy1
blO751+3rLMGtDY8z/RfKQjnw73VKww3wp5t1AE0d5m4RAeu+KkoS83DwIZR2Erxb/Wcf07kbYQ1
m1VU8go2p74dhCbDpugclrtXNaRIimoF05oT3S5EsDgobBXcrh5Jh15gK5G2ZgjQsTp7JTvhOPnZ
84DYBoenwTAXRMXlUCvIlU9CeweXnZKBCPLffn9tT1ytR3Z5YFMNhEC9I2km8A0biDH5sG81aDpQ
P7DwrkXQIAWa/+gOdiuSFFXT7ev8dGCk1VQd83ol4PNlc/Lp/Q4AxLSxso4KivqcLxqDRR1VYSTF
OE2hvlLp9oKOt8LbGB0lRjRwCmbUrK+8n+UQ7Mh9xQzDTyaZ/ysKjdeB6Z1ZhCSKLvUXxoVQkbML
rarXmg7o6dg4tgac7lJoQN8zFZWjCR6kmXBmyB8Gv3j9UbKbteJt6ERytgFXHoRBbRXWQZewbhxL
IiVpcjEfoAptbBlKdn85cOe8vBDkFOIEI4+oF1yQG/I6dXj+GSXQA3/TyGu3Zcw3Z6Jrkaj8JeHY
lRMV0odNm1Q02/DOqt1v/Qm/+3eNsxn5XidgP7NZNnrUeWfkMoi5A6MaHVEgdrrWixz+TVZGGI8V
z+dCH188TrsPRuc7pBQdudF8ZvnjRsqOfSZN/n9OlySwtA3vXbabZ7yHOujSM38sgKTkCMKf3cAE
8WVdqF9j5c6tUlDhbOVOnf0wRT2XFbWPSKWeTSozfSpGe4mdL3FQn/8TKTTAo8p0AUFcVFl3H01S
ZUv3aFYdrGDPAqx1lUsT8wCI6S92NGS7w5ooB3vnwD4SEN9xUPCtsXi15ohfblbjbCcSPTm1LwL1
q34IXr9yr9dpGN3eteckH8+xvw00fjH/cR1BBeSEkQNrEUV2CYZp7eyLN6XrltZiRY1fKiIUoBND
S4XeV9v2F0O6pvE/8jJ2sndJvf1lIyiSTGuh/TtWBXiuNsDLSkRRUlxbxHJey4aIhVJQCHQTF3d1
TUjpuKFJqHxI0gAn6gF3fPYXkMNAA4GQG7ZUIi04NSebmFoZxwoMX8TXnZQetX+Dx4OWfO9rJRQ0
9x7WfsW4zxnePBMpVNHUt8hexozcHsY1L1hbEIgbCtBqdDhiguiGRB0XyoOJxplUAX6SzeZWdYfE
oZai5Z44I9Esv2tgNsyOcFTIX9z9YyxSAY+yOeECpomP2DejTRsn7IZL5rkkCIQXRXPTEzs/f1LA
Hcq4XbeAe3ZU6EMDUsvwFtr8cwoeN8G10RV9YIK2U+i8sTEP4luNozf57cZ6EWEFWL/EMUG7YnNW
wWJs4JCQO3kKYoq8n4mkSQzbDg59bPIXPjEP343RfwQcSeYNgAr7nk5CyF82bUdxtBmE/UcLorPo
kyWTp0ILpHhzHkbdTf5lANMdBTlN8IM/wPvfn6HBORa1z/0ozTRxeSkzYhbvj+VfxqiipiTX0km1
UzpGGvyuEBxsbUJvFUsr7xqDQdRAhyE4hbGyaLKkCrAQa7jL3UR/dmSrd94h55vbzIuYwQjfx6XB
l9zYw6IDGQedzgH0tq+Zv1PpsXQsMfAP2/VafGehBFrOFUb64ZHaRMCzezTJLVxDG8oDcWjEveSq
qkKg+VqHYJ2HkC5S9mt4vT59fmfsGuCP8prZLxL1Am/YFLhVX3GGisa6mRN+Wi947vIiZsyrELG1
+EzZXJYZp2U38IDZLjuop36RYFrs6pHMP2fDRFSjajLotVNiE8AgtzR4medRKILLciZwJc/Qhowx
rQW4p0Y63dOspfR6oWqI8/wJXRgqqvdEx/B0IZ5b0xKrQqJyehWRI1RhADgDhO/sOidFakApxaQJ
C9vATTUWDy2puFAXfOogLObMp3dkdJGRAFG7+HPY/clGZ4M8gucifyqAeHeaZtxYx+R/f8+tNtgO
YQcudidG5kdW247ZmD1LgJuoONeTzDHiFGQewgWxXScj3e5HJjob/sT+fT4zeB6P83ZEO/qvm7hf
7/oxieVy5T2MSYXtvw/rGFO7dbrhUOH5K2KH1OPpspKfrYBbo8rI1Z+p9Q/mq3La7kfeLgOJ0JOq
cce8F4Iwe0pW3nOZm7qxU50SIMEmOnSW6JgS192mqUNW8X0xwxrfwtWwpsJdnRtLlYKdIOjyFk67
e41/HMAYS1z5t/vo5qoYnbNGiRviQ8m7DNinLNA0FlvXX570GK8TBIC8uK8fe5tnByI2Uopwl+Rq
ArJ4T96P/S25xRWhnU97i2s+Yt6V6lF5WoB5T5rH9XSqmELo1aLu8TuSSoGJ0DsKjG48HOOY744N
wFhfcIl8zbX+bTvpU7hCq17ZShdnmi67ZEJ+41vEL6tmOrZRklKN95FojufQfPIZhNgNQhQjiHkO
HQevjvpnYQjDCWoz3CDVKOdstJf0Ny6vqj8G7+vgS7la5EYlCXtX27dZPgFz47iNqWS4x+r7KgwY
DAXp/YQMcQp61TU72WruAHChQgiEHFu3BiGdusJ3N+KbLSrNE1I+fLq+RPhp3QI6deRmHCAkp8YO
M3cisOkvuQn/FcE7M0t9ri/F1lfaRJbExJ6r4xadi1TCtcQB8A+QgXiH0o2KZLlTBviWt8MFeee4
KibzaRJ4TRokQ3mrPnUIC6DOjn/L+rqqSck127ddGfALFHE4ulgzSvHn/yhxkfFNfy5Rw+f2GlDV
er/o7vtXAPN0Xf1kRRmG+zfYClUKkgtyMjojOmgmbuHyZURTS2JcqEYGxEt6Imi8rOT6F2uyHoBh
j5IXUtTjzQMdLIaA0fbVfkDpTAALq9GyZklwp4io9NytIFyA6YDWqbgN5O6xdgoYNWelYJXKok6H
8XwPyqWhpxCapFe6JuJq3/lBtAcZu9f1YFttWoxDpxFflw3QpyAmRz97XMGW8Vo+bF63Gpp/r5cW
7Gop28iNRjkVHUa7hcQn/BDOSFui2d65iioEJR3ecd9RfuQpvNEqy8TNtCDjzhGzbZvH/3bEYDqc
R36ws0ckOt4rqTrfVZraBjc5k8fhztZsTheH4uP42/Ym+5Biet5l4sCq/slW7123X/xKphk5K+TF
uB7oHRrjlHDAO9/JxBg27r1MQhqt2gj4W3ABzP744A5kKcLaNKzg9X8/ssGVUMbvk0ZcsWbcV/ZD
/Ta+8twf73GSepqx2zu3+nE+JilGJ1ASF2fKajVzFM2xeQE98nuqlbh2sa75UE483oGTD5dataVg
fDf3PKOWzXVXj4xBqQaaKZ1ruWd6vl4e4pHkGMRe4RBYfdJbRGZ+5kvv/4Hofmq6OtkWq1Rl1QUd
81/yuGOhe/xEhpqxJfQksqxR/T3FJEwnRRpp/NeJpNpv3EitQL1upyIVHGnHOLPFUSMKpupN4hUM
V+0NGpizNdlWhPlGQfM+qsmc3/3dAE9H+ecrraIqHwKVOVpimw0nrS6etPOcDBb5J4FhvG8WouUe
df1EbHnLpFh1cWSqrb6gD+pSD4p6B1p4k+LEfDMddHNVuMul7uutkPFHlLAqpBQOS3p4REJ9jrn2
NqlzqmwcNFq5LCDMJH+b+Sqvr0CwJM0nCkBzfSAbFd4upq61nMVin75Cs/ZfFgbP6expB3a0NytE
ZDbUZPEfW/6vJwDNPeITZXAiTJwjI1d4eolid1pCreFRFTEORVxUUfvqIJyqtUyWrfROYcYyHvGY
uOWJhiIYp/OrOG/imOq4C+jzNvvKI1ryunF0jNiKiZjBr0T5xBXiprN01yMmTLyGk5XCzWeM5dxz
aVGL2vdeLPHpFNMMpIUhnsg113KpPChJU7QxlEk7HiPZ9Nm7yz//DWlgbC4NEbYNuY9Xp5JzsbXY
zEhdgLypiYPpt0yAlPTVYxbqH9fwjWH/iiJoMJ16bN4z42LTuX+LEFjJwC0ONexuoB64uT884LH4
NUlOCeQfWeuF65m06Gd5ve/p41WK/EYw7x9q8051O890MlIMtDTAwluMeSdrjxQcbKhjhJVRet+m
t7PdEW+bvAZW420jUiVRXxHKfl0t9++1UFMiVyvhrglM035Z7EBucLcSo0OzdWhV53HYMcJ9xYF3
ezLom1abet0vZkbj3CW3yZnckWg6PBOiCYujzeAH0JcXnwfK/+YbuajFmm+BaJiDpTk+zUsEDYys
0s7lehiS4PNTJBDfoIviVm6FOX0yxaVSm/AWeWo9f7o++2IfwU8hqsK04PFVhTKJKDDf8Z2/c4ge
H0HiD8xWeJbaiNHfVgx95JRqxbWU435h6yl5d0WIknKOqEZw167hunCJH19iGoiYCjmmdg2XPZOy
aUHgqrchX4mBpta2vdq0IImxjEgeX3RNmuoXRR+ddkITRsZzKld5+T8uBvkLiL/oXVf4OB4UsPCJ
RW5ohU0CzahNmuQXz3fMTNVxTK71ZFv06XrWmpR2M1RrAKo+sYcEm0GJizrSzRwo9R3CUJhDRgNc
DL/aq2T53mIxUkdXf8IYOPuFKblStwx0SRVMR2hhtC3ASu8X8iIpJV4eJGD27iIjUWDTnphnP1gi
UYEJ+3EMn+FfAQJPWrUFvUB/vWfNmlyvXpRpcGCYjh5EXQl1ozVQnFTq865lVfzVqTSHtgIyQ2DU
yPaF5OBcvPtyGAJDKz+V+teZIFFZXihabhJeov8frsrZbWWFilxIQTzeWz45ffnRntDhQ3JrDPLH
U4qv3frNsYvMKgmXqilgNcees/RMp5mfS4mqCmNFe5niR/kBNZkUNkY8vm8NOWPU59VwN60sBFY9
1b+lrST41Pc7IV6VJB/+FBrLl8o2+d1kdrXB4fhwud36r7/IRAVtof93InO3GiRZI5RPFszMtZSa
r85ffNujGWOn7m7Hz4+KexBFHXGLXQ2UJ1mTugHw5NUQ34a7x1IyyqitAlhU1UTJhneV14gmba6f
FxMkLjBAkSRmZHpCVnsFX1TEfqrfyucFToiFHM+kPwu+xXneHd5i21+wdU9YaRvr/tnrhG8VRYQ7
a6abfep6E7J5zmIWXwUZ971YUYZ+Qo5+xAmIB1gfCwAdlqos0RFfqenMxMCE89r3/QoYZDAUY1Sy
gz4ZJ0BCzrZXjJlfGOfjXIaIsUZjW/V2WRIhkfCwvkz23ktjC0d/fqRTpCDlLrcjC9KCHw5O4UQ+
WOyZndc9wiGlne2aD1jPe7IU3xfBaNNsgIrXg30OTIu0fi6mLJEGIphkpHezC7eGBHJp7sx4I343
xjy9/FXgVav7+eanPC7NTl5dKBikxXiAJ/wKQavC0BS3HrIj1wdZRQuk5ViBTHP6aVqMkcVv8zyd
sF36aVgKZvhVfqzWV/VY/q1riv34P27IB/dQq7HKyQGezVS28CRmsF7B/yRKheWquNOI4rU6rFh9
cxmMTJfPwXNI7HiAJSyGj0jdt0FF9AFrD6VSVVjuAeKHBNnrE0kyB18bAoCzxDaBPuP1MFeszYnX
+ukst+a1Ght3jyy95mlkJEooMGeOusc00fa5NgkvBec7S199L6y0vs0uLcvHJMrXQDc/ug0wqM6d
b0PuWNhF3UJT2YayJrhqBaYbS4kAy1q5DG9QHlpB8w8hqtMphgQNQw5zTHaxygjV4sr/nUPApjlM
5KxypEfIB9sE7Za0733j1je2+auVTptVJtm+euIBAeWoP1AccIr/UXPeHzZI39pFRZ5i0REtsAxZ
H9/HyPOctF1VOs01kDL412ZS+HsF8PdiWdbj47QSiOqOomsLk+JOaguU8VikTmZ/VdaQAme++DM9
dw8N03tUzzgSiFaRRn/3EoBve91owqcDVDVJxzUYkhTjA7/yX1tqrC88OCDxeqyZHOuTdBvIAtDO
wXdO7NegDvSxWaQ6HEoW1nQBClJsUOv1MYBhMkTY/NEdHvLI3KvSiN+CBT+s/YVWUHmuq+Y1pvq3
Jz5TzUUrQBIlWAuRNaPgSEpHVAKKrSv59EXj2xRmccYxg8fLbr68J/5y8/hqNUxz9+9gEjOkIO0K
qAKE0Qgp9JeN+wm8t/YvNTXc2B8oy4kirMh9iZNeGvnb7cRH9ozZjJZpCnzIGFEIBdO9Vl8RPoVq
8O6bI6rbvge8otMCz1K/KQaK9dV4anL/uUy6OcJtYoW7LS4K7LVC371NfBjSJNf8HWvGPFcuhRsi
g+MIjzp+6mo99nA/rkMSABsxbdKMJtgPAd2T1NXX5BZ/3JH1vwxuKGnoBQDdLjZgMM4EArQ/VKFE
Otfk9KKPwz3UFwf+IVSQuOzjuir9M6CErYcRHqqJ3GhaJ1r0XFV1B+yS1IbV05aUJn8F45hw9bOr
oWO4elT/zJX5NVl6BzCYBZ81Kot/E6A46buJ7YFE9fYnDyWE2WkvWBYN7/1XlBdOy/3ZB40euhwL
E78D3SjULdGFCuIaITRbCsfGOs9SCiL0/W73DRce90uyr5nrthD0RJWiwYDrDjngnwZT5f0gQa/R
P6YK7hzgfTfZOZWUD5tHt2tpSURbFHBJ5vEGhIpK4DInJED/d/F1AEZ7aDEsbJ/exL0GukIJRZV8
ExGHCszUJAR/laRkg3ia4fXWmBLscWXeDCvGuP8CIkop/S7rAymHJzAEt3TdWLQbdgaPbs056Bmt
vfjd3dYyZSSYgDdvwnZHGSDdP5kO33V2mSpoD/sEWNJDTr5X1ke6TjRF5iFs3QvpBp2n+Yr2j2LI
NVFY+6xWfI2qsmSMkvPHyft8U0xVIbyra4NBKmeVPhl7olSAdIJvK9Kz1wnO8q/QtedoYu/9EtuL
ajeuSbgBNiPstwsp4UyO5+NriMqo9c4W5Bnsva3RQHHUi6/WsmcTiBz/kmsjKOtBK0nPPz9qavk8
FlPl/u4juyYLJDwde+98ZhfFpPT2fFndi6V9n1SIcX2fe5T1VrVWYAqH72hhfDaaM9geYAgo/d+v
p7gMvh+Spgkux24HoowdEdReR/Gzen5MsPxcfhp17sOsF5hmyqQyBPcWA2FstHjTf6VWHQx78l4W
1cgNBNgHji6tc/eDGl+rbb4p5rQvq48o87dQ9LORKMOx1hXGoHaIXpIcEF9leE3fLdhWj9IwDhap
aW+h09JLM4xVDVzIEgTbzxN4IGEeupANksESEm2b47UL/OOVemSfDyDVXwODjVgqcJYSPuhgiSwW
x+OEQpzePP/OROFI2fbLiPW78dNjJZHTHOjxcoYXX8ga6vSmqGogCG//O1N210MNUcamsD3vddNc
Pb+bV677PPvadqGf3cS54SuecyUcDQUg2ovrWnT+9whKOpul+z1hjKc/TmyTDMlibPRj038i0T7U
dNbcPbywPNU1qEgYtbGA4jDcvci7tr830qEXH4R/DeDyQCX8/LgO9P/RnupSLAyW9tisQhZ+flfM
hgDOuZ13vEHveMCUPaPkbG/CyyMa05tNQTMO79AzLrMz6Gcz7eLRoKULWowhbYbT6LsLpGC5Gxjj
htI61vcv4rwnxXIBOe+htNdSIdL70jNDpJE1AAWUnaNxsesjjUT7fYiuSr59UgO/oQXJ+pTdeLBn
8SHPY9f4H6xX/xEOV8WdeNJkGuwZnvikS1QmAgxG7KoCHgkiLbloZrwmxmH2bbQZ5WU7h5rI0IKq
ny0VWa9jXMEohQRTUI85UvY2rvt26VMuajjkD8gwAwDDnf1/0LUM/0N8a+R5/Bb15LnTCmR8suMn
BbSmjkhie8jy2VR+iFiYJuvzRGmOjsmZLSBSTAFiQIWbL598M2UudbLgOMsoWw86khv8GJmv3DsG
Su/ksI52pXRfrKFnudVUD9Q8vVZE0OEZMUZyNeTuiLW9CYK5XYaO/R32s1FfRygMsZjO6CBNtWJ7
8EusVxTmoOC6FBQMW638IF2XYdt4Qid0uWFJ9oqVtbHHCWTMFxzfRYFidtKmVa+6lgPeK37VAFTv
YhyiRkfEIAZXwbVrMHtU8zm9YaLgwghlUPJqM5cqcy9JOXynDrfyC7HPk6A7M3EjnXJaVOlOF6mN
/puPMAPeP18ub7UVv2wtvr/sOGHHIIx5Nq9g+zfx5fZuvP7lo98JtnOXUTL+5em1Vnioc69HU7Bg
OECLyx6Sbj25m8Qhe9mId55qh/ABk2o25K/bk4JSqc92KnONjtK6JhKFFDTI3HiZMhy/o/1OJWPq
EvNJHFhXs2N7DLzYRx+KrIIhNZHqx2ivOoT6RnlXpMWV/AdELGB+AfcpKcNwI28ldKHGKD+iAdWP
VlzvYfqzMrhyeo7wcKD09BtdPWV/UORSScTU2qqWSIKq0zdqlj+FSOjdHPPWbOe2OjtaWKHE/WLF
c3Zo0dj+DKlbO2aNNya553VZWn8aXhXNUzF2WxiPZakPTR659k5k4sn1fixYO3spfXYh0fjHnPwm
Zkj1d4qD8shuVwj8Od6dW+jWvVuVChbym9xpc65Y2vgakjxmAnx7QoioSy3ajpykxHFBb6vZgZnH
Jmf2ojjELh5N9J5nOsBwr+YG/1qBUIuiXNecwt1tkT5EpKbRqfYCCo6uQNTVrhDPYVpzqOONjbi0
WrFhImqpbgQLf8s9qfyssojymrRIhbk5H9tsaedBnUWKw0tyxDnqcTAfKKJMhM43K7VBoanIcBhc
ZhXTaWZEVo+CTm8t3lmhlWXerNj5BJrh+UPoDy9veAIgI2mY95DPupnKYa0k3TVrPOTllKoKEEqt
GB6bT1dvvkX5LJndwOj+eLHg5/BdDo277+9Ywp+Ja6wn3R+cbHe1soyhVAt1OZy4tLlzJX0qCoWn
bwx6g3saLVW9gyGADWqJ1UO+JWE7inedrRhkdnb0zhuZpXOM1R6or64x9XijIdRqnuoct7UrNsPM
P2OKCS9Uz3FJUwnm4AJrytqdWJhoyQXrZKq02+rFUNr1ev/AwhIMgN5doB8zG+GoNY4eN/pvWqEw
OU1eDinhd3gy3/pZKpbzklGwUA29Hlz6xv48oCkEoCcfxdSosdkx4v5625jGgZeR1EwY4b53TSvJ
t1dlJGFIxCpfU0ZNM9JplxjVjE6/Y2Qcr4g/EYAJsD5SeMg+DfGA/H6bd8kWaUqFamlYf6qEN217
PD4su97ZGtTj4C1dqk0eLIjju8EvyyPPxr2SWZmBPvhMcja/KM4ZgSCiLnlW65mtntA/HHz8/0oX
5sXx9++m5ds43rfuyrvkCweEqBxDoDpDoZBgvDF8b/yVEDLEt/+xXs4ftp4A2jMdAGVbd+ek0a87
cGobr3BqDHXb8nV83kJ9bp0cDbWzAXmhb4VPONlj5wpPtKiT9MRWiuxic9kZNs1ZMRTCzgbQtuhy
9uC2+Sv+tLP1o877Gt6EAJR4uhqbwSzUL8NVIGnCG4IrnG6Hx5ZAcuUzsIC38eJfaDXOHnDPktUf
+7137SUVudi+aZGAx6o8pMhesLuZkdaYeh8vf/WpzganYfR9hMhZg+0w6KkDWPMmzeT1UjDtpgOM
tV7nEmrGA35q7BqYbt6essz1y4e+wK2kqAXmcCUAxpdXIYQaRs5H7zc3LxTRIYMWaF7Xl/ASFNfz
WZ3E0S7vRYQQnXfmxMpvfJLmbNLZ+Gt1v6q5FT0z89TaxWULtWbGlJEUjWFb/ETmq2E9g2skZt5c
Hkv14jCkCmWEFA8ATM1TWVBPVGZjvtnVvZ/DYrNJ+VQ1Z2yFBCcmwO4zHp4eW+BrlnovSMpLgmqJ
JPMUNTj2X+WDMASmI0NGeaevhCFj90KeQSH4fu48iXfWfODzqSUxbSDfFWpvUzmk/gKyP6CNWWst
Hf5XrKsbu/lxwy1RwP5vuQq9ozsym9SyqNLYHKo2xt2RquGD6zLh8sbre9M9TsxGCs9PRCYv0WIy
MXCqvI+sVjC0cbuZvyssL7ULcQnlY9rDNQZcMnN975z4KkGho7YS96bkg6ovLb3LktyjiaavedLW
hfy4R3Pv1STODfxWWE39D2wp5XLZA9fr9kXHeZkbLTeM0UZxqt3WzI4A0TfdxOxoR0raWt82abfg
PFkG359g8E8rltZPWLx/91Ixm7Jxr+uAItgb5Kz6/k7gpEttSmufUAKhZF8Bs/3XjHBsY4dPTjgV
4+yDIdZNS2kBthtRUg9JJKIm2Gbshf8DLsoGz813C+8GF6FA9QlVKlt06zJjxcXiFG57Gc9PnG6H
A74/fZYhEdgkp1DYm7GbqcGwooN5aMeDuP1YPz0KiNPZRxov0L9x6ujBXBZgNytRx99ClF+PD05e
pfwQZuH4Z4oeiLZfRamKarAngRpwZE8RXvW68IJzGUgGVPWQu9Sn843gTiuzaNfEyyC1dyob8ElY
4eUSumSqMULPsHcgnCZU4Xb9XcjCcgTznwEjIXoLEi8xeLqwLJgQr9dAKgSSQkLADvmYZg1xavOn
BrRtoAEsMUhEMcrM+yu1RjA4hC6HKzHUVofRVOoncxjiYyD/Da1cQ16yjfjwhj6CATj1LCs5Uulr
BsbcBSqUy7XXn7ZJJ0HSM472sxzIz/w1KDyvm5luln5lEpfnrW9fkN3K1oQxlAEdMX+Bv4RtU2u/
44X3QG6mzbZrcLMlRuUstVm8K3BURl8VW5x50K1IO1mZ5gNky7UmqvOhxG1fgcwGHPUcmdw5lyFn
zPgCWlSXuLSC8Nk7FB80gHOHqWVb/NpsF/5byKkZI/t44EfWimR3JLZ1DhkQDR3o88yIm6Sm7N57
kfYemSJsmVt+D+20YRQebnNoRJhY41EJ8NAiFc1lC+z14sS9rjfK95FhAmfISNn6WgwHw91X8exq
24Ti0vc0Q5oj/TFhe2Eyrcoo5PIzxEd6frL7p7T9J1y+lf5dRIn9urDb7XRBP6lsDMPeOSABmD3N
Fqqtv9is3RAngpvaxPPuebhFr8xi+xVKEXp3jYuPkjELmTJQljUVrdshKsIOf4hEKWwxn1PnRRUV
H+UJ6of4p5Wck8fDAwm4kvPB/fnVFIfTILFssp0QjlW3Ha//anvldylSO6FRQwFTi8iLuaN9eHuH
GJc7QDXytedCv2QbZHGFrggVXs1iHFAz1VgyBeSTezeYj0D8kgkU62jmcY6ubEbMy00koFx0SuZ+
Lm5ymixUTsaASLJPLww10B/KgTBG5OXxFQTX0Zl/CZXKjDjpvlNzN/jyaHLSw6aV+ePdn4i0RHXZ
IpqdAbtFnX4CL/J9KOykYjC2P284lv++PRIyi0s4LRaRSvQst87o6yLsfyICaUCFh306PJZvAbjw
5ESIdtt6wrzF/eeUIoqyzdDBMoXfCKWCCjtKuO0gRAcSBt1NheQNxSMiP6zOjc4i1f0iGkgtzZ4j
K/feftQaQaXEtOyT0jGmgDoaE2aF0GJWthN3SMY2UUwYgxVWipvAPC2OK4jh/kEAucX4vacM9UV5
U/hzJWjx2bbd1iv2Jk3OQ1DssPRbE7roILel8d3w9ECYqM64KeI2uFq+aAL3smUOhbmhPTSt6bGU
4FrWUi/WmalxVz+D+mXom0GuQxNlwm66e0xx/bnXFPEAlK9dSi0eeVH66Aj6wRaQ0P7tNreGf2wD
P6JbzIA9SXYtXkKmAbop2I2D3wAq4ffMsDZrnFraX+9C8M2ave0UvD4ENf9ZkSAeTjOoSXHWKESw
XJMgJzK64CmfIadWvxvNrIkxf9fHzfSvo6SmvkhfMJpWl1+milzR3KE8nfBdTWY18M+s04wmz5yt
E05jKlSNejqxIvOXimuquR7UrMMGVU9/oMqL77WThpk1c2/Jar+64nhdP3w9cXEYFUR35qUCpqAG
hoDs+tk1Uurlng8YRbRXO/pKYtsEtG4LykMkEJ/eVhQ/WT892l/Z389AKqTdcWj9cvXbeTV2QVjN
9fnuV+VEEi/osZX1poOwbIBKF1BKbj0kKLwfzeAm6MDCUpeQfxRjheDbEDO6gNjLxKYjHUX5g13y
miF22SQks/xIIOUijG27eXfgbTEEjNn5h7nNs03bDZqGqlxFAIvr+Ea6J2DPU0EIUU667X+GqPhb
5tDc8337lXt3Vvjz9Wf2K9SknwIdk/MnJ8Nxb299LajXNN2b+kpTDIra5LjFjihqjt3Kc6vgPz5m
Y+7yybTVWXBtjxwfZXWrcqQ+75y/zUwdp31O5SOd+nD3jDO0J0yrgsjmC4+stkiW5mjzUh5llFnX
PA+zjIGU5nTlIJkKN4XJAJHuQDe6kxPQSj7IHk8zRI/W2d6tZoB0t8N7hs4TBo5/+psbq2pC8Ygj
hoSr5aW5CyOZweGpJdPJ8HsuLD5wlrT7XF8k7X+c4EyixuTUPUMmjD40yWUFe+sBkvvLF8+hAILo
AIzcB9LXics3nHU19rSDd9EDdSBkj/Yi/Y8kijsAwbjTdKx7nc6blS7UexqP3PK0YNjEJ4E=
`protect end_protected
