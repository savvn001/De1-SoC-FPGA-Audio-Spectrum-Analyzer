��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	�u����j��7|����GP�����|�����sm`�c��.�K��U��ܧ��N{����޲������Q���dH�@��lt�9�{�%qɁ79^�>�*LoI���$z���n�q���j�\q�B_���g7o�,���?' �So#�k���SZzЄ�^�L(OP5m�P@b�[w�W�s,�V����u��5�;T7k�#��ٛv$���Bv#�ns��Ң�7�b��M�]��A}Y��,9�����:ލ�##��������y��ˋ�=w��^��gf|F�ͺ~�Rf't�3�v���uaN�໥�ܧ��&�N@��Ʒ�������_��\ga�R�jez�:�Ͽ�ϖ̙�ogA�u���ʺ�99Qĺ��Ӆ?l ���+YX�D���N<����݄R���d��F�7�������;�k���<�ƕ�Y��Ʋ7��He��g��dp
��'0���RH�J��因7.1Ϳy���#¼N�_���#��yPǲ�#�v�k��lX�l�r�%�:�"�N��M{A�I��1	�ϓ{���W��FW&>Q� �Z���5ˇID���B��|�"#?aaaU�2�i�
�4�^�"��q�n9-�R�-!W$�ʨ��C����!aj.Ǐ��)!6�V��v�3/�|n�:��tڑ�c�̎�=Y��:���U�b�x�_H�	�?#-�r��~r�g�̫�3K,�FA���s�!K�yg�٥�_5�Z���H���K>�G�f�*Rϡ/&�P�+�HI�v��� ��+�e�h�0^��w�x���Ӆa\�����#�G�[��e�R�d�Ԁ�6������'AeP<̕�X��Xt�n�˖��[�V.b�-9�S��J�_�B��Ab�6"��t��ւ���|����������� Y��T�bl�j7�yO}"s7p��E��#VL�H!�h"E�%�)�|h}����zBA�E��t�:>	Ȏ�,�~P:64ך�'Ї/��;J+YM��K�]���D
C}o����V��NA���a�><R���ϧ5 ��?��󺅍�[}�$=/�@H広ФJ��P����w,41L��C���s	_J�Q��v��t#�Q�,��d�h��U��E�Xv.�pn��إ-��]s2�潡�_hڿL�|�!{߾J��qwBX'ȏN�����<*�*
�Լ�L]Ƙ<�`K��i�&��{�R��"3�p���`E��ח�| �C@(~۞�ۛ��Y,FbK�?$�P��5H��ik�!�M����}2�)��u,��7�/=Ç�Y;l�u�{���ġ���G׍ZMA����Ʈ�^����T6�����~,���>�|d�hTY�]o	��������j�Ø�}{*zC��Q����ee����.OЉ���a-��r꿥qs4+�ꓖ�y�&�3,�&�%�W�Mx���|�u�	�ػ̇^\�����i���j.�]�a���$d�y�����r��`j:�59����(P��	>1��!9����R�)��z��F�h 2� 22�<���񟿕�E�H��U%Nc� �2_�i�f��{�	)��w5r/h����3�Zೂ���a��ј��F���h�-|�yԜ��c�țъ��|D7@�Qխ�Lr���&����O� Q�#YG@���|�~�_e@S݄�[�|e��m���4@�{C�Y`Ҙ,�Y��ߕC���7�J��v�ߛ���wQ��!��%�ކۿ�5C�����P#����m�t����F�G��˚1��~決��H�(v�x��R l�o�y�.C$��i���)�U�ĬW6y15&ޟH�8�qA�C$�d�<4�����20��et�T@�ؚ�jj.1��/�U�F�׿�R)��|8�W?�R@~?Z��8
x��I���k�}��XP|\�f���}�"9��͒�#Fp?�Q1�+c �`)�K�譁�%���.lCh��C���b]L�6<P��quC辔�K���E�����Ÿd4�&� ��	�K�1\��n�RiM�� q��/iTG��tH���n������FZݹ>v�eN�����`�������z�TD�=h��P�����ߜ��}r~���5 3s|�]o?��I����N��

<E?o����q�5�6&D��?�u#�ݪM�p�}�g��ޠ.݀]�.�7����{?F&�|`���p̓��V(�����j�{���p�N����O�R8�E��Bl�k�ICl�$�x��	Y���T�	�8E_��py�٨'��[.�{�!sP)�؂q�䂛w�N�J�^����o�-�m�gy~ʛs��&�F�x���SV����rۭS��F[M�V���T�)�㋉Ngk���H>���}��ip�T��Q�RcG�H���F.P?\��4�O��U�(�9���zj��sw���5�����|KR��p �P�d4�l�W;���`5I� ��ތ��12�ˣ�~�H���vv�����罀oISt�C���#)Oa��b$��%�7=��{��V�������C��I�:�Eq� :�j���v�ig� ��U����3u	����01�Hc����+���7lk0�)�k�ٷ�o�ì՛Cq6�m��:��?N(_DA�?b�X��� ������0���J��-�!�o5�o�g��o�e齝 8�$��b�<N|�eM5w�@';Ҕ>��e:�ZP���$������Pp�*d1��X�e��s���[���RU�y��5�Vf�д��[�b�A�,eJ��o�@[��f�?�ݨ���C2fA뙻M�ў��l�ܾ&V������H ����H�P:�b�=�=��FH8�ex3������=��\���1����b�[ѳ1��U�E�z�G����L�}��I�1u:~���,� һ��0EM�1��,��qԩ�nӾ�@=��k�V|�X"�1����ى9�l��uV��v��(��ap���=OG|�A�YQ��:M07����ࠁ3qNwjײP���B�M��Y� ̈����(S ��2�Mn���Л�
(�t��3�IZ2�@��AӚ��q/*X��bqC�̯���S'���c?�C?ݕ'����1*�G`>� ��'<���4QH��̭/��h���yx�[�z��ݒGK.У�� ��.����O��z���p�`�j��5�S�2����7�U<��E��ϧ��q�^������\�JǾK�-�{��;�<j_q�1����tXz��C�Y��װ��@>ǆ����˫���,�G�%��OQ�t�}��'��hE�����X�kc�	"Z�Y���vy���Ob���$W��kݒ�w#e��乜,�2Km�P�3w�o��/>�>� �r�y	�/��=}�(�f�q�5�KЭ���q�(K����l����4�]�{#K[��i����C7���Taŗ;���5��x����^�a*D&v>R�>�Y%���|�	�S�Vs�a˒����d��-f�E���E�(���⊒dx/>�����he>\Ǹ��L)�J@"4	'��˜h9�������z#lFRS����5la2輕�(���Z�OC8��`���i����3"�sǲ}׌z��J���&_}�m�݌nQ.�!:&�a,���.�3�>V0��N݅��3���OY�2�2J��ku����+���Gf��J�	�{���;J3�� �T�+�y��x9��Q�Bi��@����>��:�j�	�e&�?�w�4�Ɔ�{<����D[���F�/8im�Q��������J���9q��f9�������>cc}�_5���Uĥ���-���������`J��E�����P{a���S���"�߲c%4$��.#�	�Ȱ�ɍ��bתq��� M����Bׂ�:�L�n&��LEv]dy�K_b�0��w���F��_�`"6�Fsz$�;�]�h���:�xp���](��-��Ǩt50���}�Z����K�&��ǿa�2h �łM��O`���+���]�~
<RnN�a�Ri�0��\�&�������z��-�ۂ��5�=3���0��{�x�)H���Q���V�]��t�@��cjƱK�=�ج�����G���i3�����&�
��
F�-x?��f%�
�+�L����
��1rUK�
^a�<׿�钎9���!҉��|LA��Y��mU�8�An���RϨR���e~���B�Ì��6�I��8��^���:t��P���dV&�#�Kl��(�N$V$~�_���Q��D&�"E��R����r�`Um���/ ��V���y�F� � ,¿�vm�=�@���:O����eJ9�0.z�*��#i���a'����fv�d�\Sr��f��ö��c&�g*ԏ�/�ClCD����:$��/�EY�L��M	��FI�-��?
�p�_�Ǔ��o�*���	�E%ZW��T��j�HBg�r~zݷi��Q��ǚ�Xe�e�|/��u��k/r[�H�YΓi��A�(�#*�y�����+3o	�Q�ˣf��7\�wvnZ�;��-�rt��{��EF�Hp��y���e	��O������0���V��@���y��F 5̝�	�E*�k d��6���� Z�no��x\�Zw��bj�S���E_}-����wa�/X:z�s=���륐�#�a�WU��Ȳ�ϊ�L��!�����/#.X�Ŗ��W����Jt{	��Ҫլ=\ƣ9dHZ��kXv���(�"���N^����P05
�Y�����ve�����i<�RY�=B�j��O����#���n��X���1f"�a�˭�[�aS�+Sc����=Dr���A��-�����x���>�P�o;�6n��չ�~�`�F�cðxF��2�5}��f&��} ɣi���;*i�~��p^A�4�5��R+�G�Z������Yhg���8+`���}�K���`����IцO�򬋁���^��}��c�X��|b�fJ�e �,p2���uq�Ia��&:~�J�@�S���]s��z�A��7
i�)��\�*x�`f�.I���Ɓ�3����:�8���ANtvޫ>�7|yW2��7PY���k��HߖVϮ�ol{�>аb�����ЕZ�o'�S�&�=f�w��DdP��1���c�����O���s.��.���nu6QK���iEO��ʾ�uj����`)'�.��E�S��� 巿AًMS?��X&��d�:W�y�~6�ʄ<���K�s4�=R#��{�`D	� �_khU�
[�\i1X:���$DqKsH�!Բ%���n��2vF���r*Xy�s4��?��|�_��}���K�oi��Jx�����M�<A�+'��������Ds ��hp̀�}�'e4���y��ݕY� �猔h?�!j��S���}�[�ץ<�l�~�2��zm�\�ge���"E���W�ss+\����_v&�4gW�B���"��z��)(�s�nMٙ�nL�&Ua\���|���*� ��8���J�r��H�oj�w�_'�*]������2Bs��:�^W��v��Mkdtf��F���)�M�$�)�r�?~
A����L��Y S���$�	7��
p|��V�} �����$�b�a��/Gc���hp����(�Is�E�y��C�i��3�2`Z�r��{8\npՏ1�G��G��iQsD���������}8?�X�P�Y������\O-N_��Ǝ��Ƈ�5�	WhM��ʇ>�i�6)�e�ܟX%���~��|���]�)���vل����\̏@3�8�9;&�/�F��A]^���Л�����^�y�E�i�	M\{6���t/�j�P��%�s���1axVbe����j��Sy�,ⵆK��Og�a$�#��gr6q��K[�^<H���'�\[��q��-F����٨���-ե�`Y.�UU�qzNNԱǕ�>����D?ƕ"n��3<4�TlP�����1f����c�K`-�.#p�Ef�����(FV�!G�)��,}��O�K�&w�� �Y��
]����U珏��?W��/�c��R�s�[<�!b�9��ݶ����Z�C�<'Ә�7�S{}�yX��3��h��{�@�[Eo-�Ϻ�0�WBϤnMX$�'h
����E������S޼`�������i�h��#�@�f$���%6��H�^w�R]���3�5�K��������\�խ�3Mu�;g����$3���Y��^���x��j����.�,f�0x�H6:�c��f?���@!~�"��J�P�=���Pt���6v3Y�vX��,���sY�]����� �O�c������/�+Э��0�/��t�B��o7����ܑ$F&�E�!, ]�g�Q<��򜺆�z��KY�Ae卦�O��J��N �G�a��&D���9��V�h���__�1���Ev�;v�~�̠����%�QVKɫ��j[��q�pkޘ�&�ǘ$-ڗ�8�����hD���I�9�����͝U�h�������D���Q?�1�> ��P���Zq1%���3t�����P�Z`uE�3�w�p�Ft6���)W�R��@��صՄC�3�>�1�m�����3�?;�k��>n�������m����^��QT��x�6x#���sŧM#��v 6�- ܌�L|�$t7P$�U��8`D���Y��<BA�R��ך6\�k�j�����?.�\��,b~-`Z$��i�����?�>P��L����>{۔&�+!ͪ�������X�	x��c�u�&�����h�3a*w����b:VK<Cu���LeN�2�7Z��ÃJ��r�"��Q���^����݌BERwUU��F�b�:u����?ɗ�B"�ϳ/.��D<8C ]Y&�T�jZCD�ݗ����=�F\�%�:2|��*�_� 'ǭ|�";��� [��Q�}�Nq��'I��e�v�����Qj@B���c^�O��<�~|��E��Z��/uU�q�c��#�6�-�(#[���-]!�$�$�JLͩ}ηS Q�gI��*���>��zm;�4�#[��,M��3��x��(����+�0�t(q �I������I�D���	N��p@��ߪ��g�n��'Թ�Q�a�/�	>��.+������6�`U��+�ܠ/�U�~���!L�ߍ2�����G?�Q-ݶ��%]'F���wxW5{Y��L_Yڇ�L��U�<]�N�>}S��2ۨqG�;nͻ�#����ax���L��Ur�1i��ƀm8�O�=�nG�}�&����]�I:�k/�`��)��E���9U��w�����cCӉ���s)W7�`���ݍ�
�oj�8���.A�/��p�ݰv��0K\��W9;����"@�v15HX��B���%�D�eW�6Ժ���*>i�J0��)�����@�o�n���ѳz$d�U���ah�~��S]��$�Wy���� j��(�$QRȬ{��^�'̄{�)�V�C�q�Ct|*�ֹ�s�q2�ok���k'�.�����3��J�ޛ\���9�b��?� 2�V�b�����Ѽ�� �7��s��~|N�gg�'���/��� �K�9�ҭ�U!^N�d���f�ߡ��VH�E-{Q������ź��&Z���:^<����6v#4������'���D#�p�T�&��ҹ �N^c�i⏇~���TtZ�j�A&�Xka��'V ��`l%�+	�ĕ���U.��)����q�H�@�U����j3�
����?�l=.�*�-L4Tm
t��٧<���� p�CR	2��z���u��Iݲ�P��Y}�q<��oYb%T��� *�?�c8`���ԍ �	v�e��=wnԱ�^ט ���Hs�T_�%C
`�;O9�[a �� i]2��k��cp-�!Z�K��HC�X�9)�"F]�JGJ��G.;���^��|jzd\\�`�e/ݵ[��~� �nn��� �X=���V�{�SP��!8�����jB|93��Km߆i!���M���l=�`ä�:@sG����X��;����=�|8��a��@��o�������7�_A�����|��S�a��H�M:ǵ�m�?2Yx��jqC����L�t@|G��q"�d�d��ٺ��t\0���#-`� x��[�,�7�%�A��AJ��u֡R"a� c/�/,z�^[�')#��q�8x��� ���S�{��ڋ��to?Ǯ�H�Bk4��O�1no�$��,s�vA<�)����0���8xg9�l�.I���&���SD�{.�x�/�x�A����y_o�o���f�������2�0$Q0v��x� �����U���0��l��i��ͧ�����;���\�����i<F��$�aoUc�v*������I���s�+�Z�ʔg�|Iv�_�Y���9��W,Hoy�M�@r���\�9�ݴ��.G<�8$�m���X�>�b_�a6����z�i�K�K��_vf��@�?��k��U��J
�����N���ɇ2����G���_7���p�p.�!��TH }��(�9qJ/ۭ����q�.M&���
����) �W�ӨKnwXZ�TO�ig�[V3��dӪ��Jki�^���-��ټd�z����JXL+l  ����V\�