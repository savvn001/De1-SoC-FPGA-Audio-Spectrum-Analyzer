-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
z1xMz6jV/3s8uevPw03weOF8qHtHUDAdYDgLVf/7NRu+ffrUE6Bg9ziawo6xoEyzJyvRdldnjBD2
j/xxvDote4haFaAIw6XV9ZaZOYaJbBN1csQZPC/Kr2Qa76GgjO+/ECFhqu9lEE7hPCq4tbxYphDW
Q5MWhbtxql3QHDpezvDo2ST2Sw0s/p5k6Nkc+L6FvjQZXQjMFeqe78stZ20TnPlWBkeFFO3frQxQ
f1Q3kV/8SS3Pi3imoXwrva6R45TpmZW36ED5s3B4nUcumT4DdRRZNo9eJqjKNw7atmKOcSGZNA7X
APLu4ilmd5OCwP8QCD8ut73LaHZHLTXDFvHpAg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114400)
`protect data_block
FdYfVBezc8rk84RqnV1JFNOlFi32tBLVBu5P9cjG9xrvYuowscxaK93HNRI5IGOy7K+E2Srx+sDi
fB8DvwgR3xbJ5Fn67JD3MeHPWf+U8wIEGFYtgPsrRZ5RWPULat6+JCBUUBxdgshmB4IaUAowN1qD
aoxO9S8RR7G0tJW/9cVf22tjpfRz/da1Hg+dk+QhDgMGdYO/ngxNl9mLdGFxTT0UijHXFDLJTQSG
vWXIGRWxUcO1Poei93/PDtmFZc4BMezav3GNasiIX+pdAY0pZE6mdINlqA5rdMamZc1gZXp4A2Qj
0vUKWjdmhx0w3t48DomJoLKInK30X24aRECme29BgCEzGzOQIoxR0Zc8PUqJkgvnz/Ns3FKHfF0r
NXXoXD7/5rMF8DZL61C7zSp7gx9uDcLSxSYcP5or0Jwxa8+fOP/bW2rLV7Y2gz8wjVvU2E1IONea
Ni8m8eS/oZ4+zSuOe08x2AN755rXMJij13I0KSJpoYFpzrpy53HqRcmf0MTwJxjiICs7dUKvk45b
27Uya8YvZPMRFk8s5/gkeJxBy5fjz5PgNIcLt04kkSvgsKtiMOeg1BEDuFKQQpPpzbb9IMioS9Aj
05a5uKqUlo6tFxFYfViaalGcPG0uMyKiGKIyY0D3xdzcb/fPPI674L//geLt6zZYZJ6yKYW+14Uu
oIMq+R28i6I/HmNDA3ffxfIgFNiMUJfO/WB9ZSoyJ38VPAbiaCaTuDTbjrrWTbd2Iyud+1jK3wdN
IETZk9YuP7U/Pq+vVZ/G2iGy4Web7CZBpNZyyQsoy61s+Y5AV2U2Cvt+qfU48D2jU+PvrRYJgqyS
fLXANybrVPVgGXazHhQLeraKvc9LR07HLH4DtZkGomEHW2f95FNt7yhe/zBqXNzZN07rD7FMaqpN
kx4/Q+XlZZfpdazEy9RS1gW8bu69hk5tB0E2pC5413aLFV+ji7CpfQcFjulFQyV13qJQ0yuLN/hK
+6A1qWbheRPdYG4n70PUoTY/K5JyNpEgwmaryFnb7p+fT8Xc7djTouTVPFtFB4DkvCxT5LSY3nRm
Dfws+emGVjKFNe8/AKbeTVAE/Bz/HCJ+qVBC1mWmDLrI9IpR6aDOd4lTvB+BWdjR5KntXd8n0pPd
rmSE46V8zcI8vx539OpySiTUkER0PAjG4KytNZs8dWao8f2yWre29wIwTLXxQQd0iUWAaPYb/zjX
f+UZBA7tlishy+pKdDxicDygnzo59aFhyTfV0mCG/Y57uR8/7TXE4NwpL5LoriKmtpl3Iixhpc4r
PLjowtPRWcTIhoaXFANTC8zGRXvywAx1KVOcrQx0Wy7Y389whSt9GuAXYW2xjn2rtQM8eJcS/ZYc
FBhr5rQKunVEfYuCEDyAk2A0NQZM6K2GF5OKxWzTkXFqbfVfeFicSuOEOVYv91T2Xwp6llI6t9vX
kZxihRRAluxa2BSa+0fkT9VUEvSd9tZokIWq2gFq0MbJ2xhk9aLiR/CnDeiv10fv9byzdeJF5u3B
9Kv0jCWHT3cVR+/NL+sTCptqg1IGRbLr8PaWbBXfVZLndz/SjO9ObpTQ+6q41eC4zuDKOcvf9d7+
zAqE3x370wl9DJdai/nVRH76pDOKi6oMYHKTCWeVq1Lf89Cc6trg0if4bHS1mhhdKB2mNQMBkcCU
xjtR4YcTfJj4zyCT8IS3+qWDjaVpnXVd5x4ma5nK61uAHG1Jir+8xbo+cWCsNmANbRQG5jBbhBEz
chmS8WD1WT4u6EwAsurzWtpYmYmGX4Tbo+hV8MQNMWJBxTTkrIEFdZUkBD7CWOKUeXey2OBBz8Lg
1hYAm3eAFzYbsiwGaxacbrCMqVPdIhMvCqK913ebfJ9TFfq/+70ico0Tizsw4skYlTn+JC1KAEYi
atBxfdYtYbu8zpz0bOjWICyK5ksI2pxlADfZD+pSxuxAk8N2TP854puVblc/MA1aiY831C/BC5pC
P7cRsWluVkKnkF3/syVbUxouSG03RtFGXfdwFJqGeWUvsA0rkDK5SyWtwUl+z6LOQbvaKS9I9d8i
jvJXDh2jm2mds9xpKQtEKc61oBUH8nn373iS+EaY27cXLMzHgJdcYcJopzLlAECDT1bl+7S7jygl
JvQI4MZjxPMKlEfJKINSuhlnnBI+dMFLc2naBdYUDOzSXNuk25LCXrhVZkqgfynE19dc5N5Qa9Uj
RA1jm6J5O83yJsskG9P1fx5/G9BJrbVmL11NriogHR0M7J6Y9VDb0/bfnhrs9HX3OomKvX4uHrXd
lwx2y0HTl/8JAsiHMYEpDZAGW9SnxqpM3wD2ew7jD0WGzCzb68TAk82DWUIxe093gx91jBWvt6Oi
rtVrky8SbhdMqKITPdkpncHUOccLFKLqToIomQwRwaKKkiBT8m/UKE+1twTPM7rtlJ8KL35kny23
ovChGB5N0oR7n0PvXnns8GQEQ21HWe7T5zo7kOQgvwt/5jI2KubCs4c+exyP2iLoiT5Cie3bNch7
JoTvr//z68O7UeD6ZYI7MFDpWx0pGBFPQD3ekSai5Oui3k8N1AZCjvVij0V9WnMIafofCilsG9EO
aaWNxhyxIWzBPxRFHfiWfXcCpxEnONROIPfLvvIbucKnE4xMPEi45bQh3sSMXkmvgdj4E4Z3GSvT
ec6euOYrg4xjxFuV3J+rBWJSnSlsT0+hNLG5et3xZSsSgTqL1jo4c9lEUwXooVxPYSvLYHqEGUzW
AF+N+PJZMTQ/ohT8w0T5AsOpNLJaxSybn1uHYdWT1AxOxuXjIwQ9CkoA0ZYiVatn5tvP6mN9GO8R
c5AcnzY6I2UAEfFUNh5DxZNWWgz3+0bcqfDI6QTDUmdt5MXEi8rq8b+cqev6FjGazlpSsuLhEvT6
+8Ug9eNlKeiN7PuIMshtg8SZBSv3fpPTg2FZUyk2WFZmYMJLUieUDao08vKjLeN0HDymYv1CZXXF
JxSmBZc+Gem17MEWWfF1CO2IzBs7YKlIp341sCmVYpy074JNC/VpJCYV2noI1ulpmJbS+lvhvngw
U2SsGiQHQ8fqvzTjHQYSKm8Bivq4Qvgztzb8vb+Yks+MYSeDaUxUHgfsVecNX6PFgaZi/gx1XLlC
2LPKO7YYNYiUDJcxG7r0GuwdRUVHLNCWZMBszcjj0Bw4an+pJU4MWA0rM9GyyRSkSO5DZWZvkSZ3
hg6UUPtpcvqnR4NytPbg622TLlQxpnObfY5TtsbRLmM+DI2WSt0eA4ppNzoEMfK4JSjRkwefTABD
J9hV++NmT5tDLeVFP+YAXn/y/tdDQWeQUG5KDIbDILtDNYxIWToL7MPjES+7CbsoBqwl+CRbKYbv
cqN+6gWhGLlY45E/AWfq1d+NPB8fsrYt3rpvD/9Lzydj5T0Xy/njpAd60haydjVCY1syUfnfMz1I
nQch5NzN6ffZrfd58o6sNr3gyCoAblSHF8J9SuPsVorfisuHAVu2+AW2vbR2IQeElIMfDe95qPxF
VSDRr6duk0RWseef32sAcnIgWa4qxRp4DDV/DU142iL72dz6KYsAVfJRKDnW6hEqYMRSe02Nz+cr
UG0i36fN5hKX8+h/YGJ3AanfobQoRYlnIrO/mcuErAAWVNbtqtAKx/GuvaMiBCyL3RxOHLUmoyFw
ysw36jt2oNXJV2OUoPUYM2bmHhVfH91Vp1msfxekUPJn8eQq9+t+Nb1Yu+eOzVmWSANzMqGOxeXY
drSvCbCgi7ZwiOjlAQomzH3lKTz+/qZM4gxl8cmWk2J+UseNdoYeepxI9Owq8IkAqfYdJHuFyVXi
vlW15At10Q0ODuKTtBYd7e/vRRpgrMFMhDQapVZi5KQ1CSFxPN1VIgFdQ7/A/CnQrxZYJFG/ZA+a
gWmdrlUA+ZcZ/eL9VjD+lQ0Fj9I/nGH87O1/oblJXrEZkGj0TguQ40JnaqYgytIO3rWAe3NhpVXS
t5OgCv7gD6lpOrPBW/tgBNFnnWG7QHYgTzsGadL7y+AEsjbuWqn1ndRAq/kyyPYvqbUV38PcQPE6
TQml1o4GL2ba4sgKH9JrkzgluJC5bGmLZY07YQ3q6H5fPHstyV6nltVFC3qhfdVpDqlV50NivZVc
XPx+lRqHEAgERRXFZ/PwXM4VH2W1Abjcqs/zEtlFMuY6cKlV3+WIIFypYf063v735WU9musGT1gL
BPl49v65PIslnkEgeLZSvSXPBL+GURIPSWxuiabW5Msh29lEc49ciUoSWUgHEKrqeI1w2hA0dLLE
zHKYwHsLsx22am39CLwE/r1LjaLI1TbR2+gDJ7TQ+lXr/e+bmCa+ASqA21puvRrpczX7PPxP/iiQ
nZtrcSlMo3IaRBUWs3YpyMo/kcFljMmGB0pm+KFBWvtcMlgafpD70nLWj6q3rN0O2Ls6zqNp95Rc
wYRBqXzB4k/Ks5KLcg57VqoqvNUp6LdEFGeorqpgUpBSCYc3ESJX8NP0IBcJEqf5AqWjhjpfaiB0
LrrRkMvkZskUiVHFpLIl8TSWNft71INQMjclwU/bZFYzgs1KNlasyD+B6MW2tSEdKzzUM7W3rzw6
HU26AYSVUHJya+wrnHLbsTW7MuOIqOw4rZdgCC2nTqKUqjmmAVVfeJqcSHDYFYA24kVkrTnoXriz
maChD3ASZlUBSjZGXVHpWh1umv98Yh410kKXChCeN4KPqH4ajfH96Df3NUCR+OlHOaHezcrMeYMC
keZ29fculPHUGt9qwQYxss1PgF+prOHyzHmY1Fl40cd1V0M6F36p6SNG3lP7LiOneRnmWGh53Zxr
kEdoqHzjUCsavqWJgmaP18Z8b9evWnixFYXa3BcqTnhQFVQ3I8eszNg0FSEoQrgk9WbZ9orUlZGO
KPknwWhq4azKsV5qUttlb2T2h+8gGzAWUq2cHwRxe/W9MqWuCtP/ChDG7V41U/HiBr4Rkh6q0Lj/
om1OaE9/fwyZ7DQSnM5Gd57fARYR4om/wDbCJ0IWwI1xE953p6/VyFtpsuHE0qkAe3IEXKtdXOsf
qAbX5k+7QfbKdNazuwcuISOIVDTTQujtPmyUO/3qO5Z7lgscdoj3hVenfonp/qWtFWiP4WePeyBj
viNIVzDG0z3w8mEE42QpMQcrKghM+eXUpdbeY5yYCtJcFTLMbqwkoDmhiQMFr3osrgqVctSZRxqo
CV6B+w2yfjnzIyD1SV5ed2hs80AqqCw7rpHCtj/yJYfXMrcYiFzjboeuYx3w9arYVTeaqUNNfY7n
ksxBXJ8QwDdlCRi9oetu52wCssphncHBsG9cplqL2NeB3JDO6tD8UlY28KgRPeLUWb9HJtvt3HB4
Xr74GKVugVcjkwEQKHzWhljMNw0VCfYekMx6e/PpEQ9sG+MLTVBxULxinDgSNAdJymioPJhLkpVq
Cei1hwRahlpwRPSeBsus6e3zfFIEf0FRVoTmOHmYWC8N7XtlUmW4W2xmklHeQQKYEWCTmG2/0Mgm
1RJrLk+fbcwPGNe4K+Q6c6wYedY53saR25zBb0YJ3a26ixr5zhVw/e/1oUaOT3VEfhkDjFG52fxw
OV4X7BPOWskU+DVjc7xAA5y8qrCA3Fq5KF+gzaYyDxEMY93tX7YfV7EaSG4+GDzcwHRcVvVlIUK2
lNMNEtl7728RenPLvEE0xYVjI6qWmlndoZQ+NY+Tc2Zb4Es9TXr/3KDy94BjsATCHrg4hS0jlSXD
5k8MUn3qeS5nH7VMIhzPoUiT4D/x9kp+FaGM4kMSHOaDm76SKZDtufVHXVy/uus4cczPw1HVtAwo
4IOKcU2fb+piTRr8dJZCWsopipsbMnM9kr5lH6df3kOOLNCHY+2pHVddFV7b5g+rESwO2pAlHCT9
vaOZeVV8fugc8Ad93rOroiDCAPQZcp+9KmjA59M4lN5n08oLRuK7oI16tTqiEF8p7wmSCodmoC7g
q9Pnn1RXROETuaP+p9XGx9P13QSN4llRAkygfU/jLgKWzd8elgDAX5x0aVuFaoAuvo7hoADChv+c
o4KXJ/jqMHac3/UKepKhSOgI5fyjqDzZAQrW2jDkuZvyRIhLXMnDpjNv6gDXdn6sx5s4oKoOkMxW
iAbKzlciP/SIxhMy7vu5LZFNGqf8mSSK67ukhrcNFCxEXLleLUGTPO/DO6wvJjnqdd0OtJoPovNq
EdmevYyz6Q2Dwg3TpBC5APKnCHDl60hHAYISfXYSvP/yZNpkT8Oigdct5cAKbTLCLO5kRfrxONdy
qZxBE6wWVZ3Q15ZzBdtqERP9YJHvNkwukxEV52jpDTKMiCndwjmM1r7nm24UrQwjvTaKiTxU6iH5
wrK+lIei9iocD8oGeQI/4U+R6LGH4Tc1A3DIfSJvJSud7TdbsMg6vK/FsxnX+SFsv69rB8SVzHyg
DlVCVUvdiksIfDmmgD/FYLFEktCmyKexSpd3CbldUuIG+TmbLze5n6GE16q5gcckYPQBQAM2p5Io
3n5mLCPs91CQ2mOQqh+jAU3dXh9lriNtFSL+PAPrFkehSeyjK0r+LD8XKlvplAxVjHHoBSjnHMZY
zWsfJgNANQ3n9yH9TuabW23EwBIN6FWgDCoNMAioy/mO0xokQKWdtwe9QOh3EfyySCnAcbtGRyrD
atDPaWRALK5CDBQFQ7z+dK6BTG6BubEJtvizRcB4oLadOABE0X7jMdENMMCSyZwJufY+TeGqgEQt
Xi3byA6PGwEIypRc2XGBQ5mRYrSX75AUyJDMxv/4snefvAMMKNRHgfi1VGZippZMOVeDWXlc6jxp
oJa+/1DutcJfXxWgwttnT4z/O5NvRHAEjqd+5U4ewX0rBy1cKhTIDABLNAgVADaIqu6/Wakzckeq
jQAsQ+6mie8VIqRhAjm3yrSgvsuN4SC0/cb+bmoe6YwR2QkvEGJHl05xUVNfSEyinvweHm6quMDj
IrvaR9CTvMi1jgUzBvAB04kB6cWSBCDEOA1QLZLLEibTGeeZhFLVIKZN452t2WKpB32uz5Yh71eU
SLw/C7zFSjpQmE0njdGF/qEmT4pu7Zw8FVcuTYHyTShgyuJHND9NpR4Pw2T+IrcYUeA/zwyJBhny
Bjyy6ki3Q9Aejmgt4oLZsnPYi16kiXQ+dCw1od/w4RV/PNGKjp5L9UJF1L6+nb4pbJTJR6hwhSyp
Do2IOnhAYdBXgtW4j25dxdkO2AWCHTIqtbjhh6vueJOeyWo6O/Xx5w4A4nXaatX71duAgHsfYfnt
gwX5emCKD4+oAxKxQbQNyY/w3bIrTvdwqWq8h04ri6fNsNSpWyzfuvN97YP+evRvpQj/zPa2ITxM
HXUbacVMCHergk+/Z8pgV79Ol32cJ367As9uBOmeGLmxwvMpr2jedSLfbJ9wa7k3bdce6OiP8NY1
eqP5rKunEZNy4dfFQn751rFcSp1C807p/olO2B0M1C+xDBMlAiZgyMK0cx2ydFmTK9mNmDKrXehw
IWuCi553iW2/NHYUUyHzwwi47g3tvk5pu3CWXHz3354Rw3fJHKfZfXZXEIgIUW3ipazgcFpcJJgp
GxLM1pWFoJD34Kg5Sjqj/l3+kmNYrTDWxKy64QBqUpiPA+wascMR7/RfKIfVKe5aD0f2zC4rYX5Q
JktNIVq97D8CCxj4sZVkIfZ6Uup8kKYOJW6TYE9nGq0G6DjynSwfYR18rwypxKBQxtSTB825DoWZ
uw11c843aMswLhYwoq3xkUU8EPvjuPnoXqTA9aQumOPLO5ms0UIxsHFlzEFSHrFM9VjglpSJB3ZL
wLz5Vvil+7KIZbjV9UIoswWgYOmr/Pj6IVXx+GCp2zC0Oq8ahedgf2M9sef1lCXZmpLcts6s2U3N
tdLf5CjT/b4uooWyuP/4Qtt3NGBOFQjDrVQ8iNobf+/lOlluW/9vOfrLhjFikoXOoo68SOr8LrO1
0xWiBTY2BduAW61MiMeTE7+GOZ1x+YBWuq24kEVtM6UnVWZydjiNS5kTTiANpdyoZP6SBLzxzlvR
uO2rFcUe+R+RYaNi8FRzhleq+khHvh6amdo1mHdnkmTohMAIxvlgqzjrmOOiYNBNmUqjmjcJTcUf
Uhj5jiT5GhhHQN3p5xwhWjtvHloCgLVUy2rJYBGf+9V7XpF8Tvi8SJ/EJsR0MJXF3Ziax5vunAvX
OPcwUPZfv4P+Cxvn3G42O1FtZMEPjHByKGEgSCNnlMUn0AdaEZvtYFtr1eoAZvXNlQ/cz0J+dzOf
GbH9wyA7BdTsfcCsbRoXEIIxsAA2W6uBpy6u5YkrojwiNMjwWspBRF6t7lOlq1ek71+kf3tfLSVI
v5LtlWEy0Xz8m8AuPY3EoIhNSogeY+ancoFJ8YNWTjsGk+RpoofTEDTbQV3tkZJwmXS9XBNc7UKw
L3I5YD/KFjsoauVIZuUG+aEdUiF6hexdwzsCy68WWkyFEYkipAbMjzN5ecxrc+YavMtlN9HsB7aD
tZO28Sy+CvnsLJlkFVkSoVeXGQuMYzCDibSkQp9tc4RncCq9iqI/M4yT0JWF4Spl5el65FdIm2dX
2G39e6xbVO79P+gV1bT+w7alw78JM6tOwf3jKDFC1gKa5F7WXetuSB5yGCaryhzBrdVPvNp7UPev
ymoSIueuWVUT8lg4uL4xT4UMv3eVcrV8MPZYR9Lw8sfX83AD+By0ZnKtjNFWzvIG4WyoybDDHphv
Pwl649xPn6eYIVvdWjiAa6URifexKvLjmnG9sKC4nt4/uLvtwmPayp+qem6Qd0vRN1h8bUErA4lo
lAphs8EmO2Z/SXO+HAPB1PNvbhMaExpV+SCdc5NL7TrpIi/a6DVhGt3EYn4wE8QSHCewSfVb+ZJ5
Av6qkY4wt+ijbdIRLVr12Fnb5s7J+uOgQizeBj6DIILEufMaaaXIeZv3LT3i8upHyQl0YIZV6gqy
hpoOuV2G9spdMxBhQzR/w/orH76gvivAdykjTu0dDmQUhv7mbJar7pN3agMeh8/bnNqcP6cgEI7s
mOOQl8pSppIz6oo5wJtznWNz/mTF6Dkt+kEPHUPmJbISuH3bMHGIbhtf9oZkoOC8HK8Jz4dm/CvS
F0eBliRLRHnhCDPsnKKtvwb0fImc6qkvpcn3tzQ0kYwObawX/k6TZlVMgHY0Kve6sCcsCiXUgaG9
fUCoY3zrF1GIMkdAXEkcWOqsSkjDlLerdoRO0RbFdioGv4kYRZMdeskmqx9LkElRcEqIsM47HhCV
exntchVgldNR4D4v4V9T4zQaBVyovzb2yis5DOGRpauFooHmSPzRuV5c0YkXQeAxbGDxCi5vKSSC
BGfPqSVdiy2e+V/GUsM+hm1nEteQD/+pVrxLPxGMTEtmw8CgG41KnSslyO5+uMCCzpdtS0s1J9qD
Se5imuGR7gxSfrtxje2TERm9rI524fXQDKBF2hKmTw2eT4oY4J/TkGAhASJ7XQ4xg+QEOZhl6gdk
KVDRW4rd+7Lb6hFe4v7XTYfB9ifzlzVCT0DrE6tT0/aPtjdbLb95QWHdamwuWMas2iDPp2swGjLi
VzU/wix+ynRMbAwKnkbVnLmzP+thmKqP18YiDiAiVMzABVGvMajISKutyjit7bLsXj7rghG7EYHy
Y5RKvi1aVaD5M3lUFoKkBwgIyI5bV3WzkIpgzzSTh8jiwRfDWklzlCu1XQ3sehY76QCjMEQdoMv6
kOqA7eXAtWysJlAhNyta6wLYrJnf5AleHgMA0rgOBCQrNJzb1SiTUkMns9PDEbFo5ePXESRQamzN
1K8wlqs9H3Y7vQsPKfmD+hptsTY118VNjWObxVK7EEWF6JxTOOMTZhFZRGdnix9A91FB2lxgw5XK
s2beEye+Xfvtm68YfVSItzQWXylDvyZODXzaY7FTsE+TGtS2u0g3F9spI6Bztz4MHjJ5878msj1K
yYssWsKosP7sQO79Yr71MND+V93QObWgLM4rwei/nwvBH/JSKbxW5FD8CFAQd1Pla0LxxTz889NN
xtS0tAw8fTAqnMHJPGzDydObMVo9wVIdCecZak2xRol6rokHktnJeB+CkH+0iJ6mBpxbdACQyIns
jB4g3GcOyq/vw66lkqoGAnsRkzGZ/is3LWQZhMXtVC7bLyqB0FYjENE6HymGrcdo9edDkgewn6be
aUjFxTgjs2NPgewn725EmzDg0sV0B/z+liBJ5EXFzSLHZDYT6kRu96/vTKullr1tWytEwJR6uhEG
Q5YlbkFIFO0HPnrta9LzxfZiOk6KRjwO+BI090NqqPNKb3sKkKNhYDqixl9g0q964eXCTxfRzCR2
0IK7j8f1ZvzZXYT6VQgTX17O2rAsxIjIC458Al2dFwJ9V3HJOECG7MpxruqJ2VC1CwRzNZgzBglo
QWHqIvY8TxXs+88ExC5MPZduE5mtmGlrNAIPwnuDg6GKVDCmMZHEb+OpkuZ8tlOk6vM/RhlXFR6v
cOnZ6mkQjbjeK2uJMonk9AW1dZMfKQ1hJfmGqviTx/Hkgi+9SxFxl65x/Ziz+2W6La25TUxqWQlA
nZL4CR+KhvwTahcceDD4FV6vkQ+Rkk9aHNjat8V+P7Cf16EIxaqxW6u4mnHY3mNtAyk1cHCKTlzG
NvJjs6+R/byHYmUapids4FzRC8qVpkQW09p6Qo1um4Onq6N1D254MevsTTfPtR2i6GK5qpJ6J14p
lfdN6MNvK7JdgYMt2Vmyj6ANRA3rDnuYvJoU9GXhAlKffYcGHps6ByXECeUNyX7v4R3BNQzarahx
00qCFa+ID73IL6MgawzdJ4uZ90VEIp9Af2zxlH/NJCIiXUJSueh7Xg19KSNDXut5n3tXKk6FSqY6
GE5/mj986Pq7VJyQtu+DxH0Z4DW1YMPJogaosdo8XmhDQy4fdMUFaQC2ruNEtk9uL0T+dn/FzH4a
MBRpz880llyftUn1W4hZxUH+lFsh+7sFxLojXx3opc3stYr6dYKBlrQPVfVJoywe0G+qLHj8qake
dN42zzwkLmwX3zdSPDY3LCUorA0yF4pDG8QtoTuCkTwV6IctCe02DtgkQQmzpmVxeN3DaeKGN+4M
sprrWpz7ltbCyXDu3s0jBmSl9vbDL6u7AU5lcdlUgyYUbca3fwIRLpR2M0MInQqFN65cZ4KhOrpp
QuTBzb8F37UxX7m3sYsYl6dr5dA6IcZCmM+ztpzjRyYXkEDZOWHIJwXf29EYP66ZIaP0Fc+crA9Q
cdQ+FaHzzZBxgoMPxlRVEL0zMobpt2OFk0Ds6lLLnbhPDmkRqV0p/qbKZqFPQQLi51c7jB5aDmMs
QgjUcpOzK6gtFYxshjJzfMLbSWXlpG6HJt0yleA2wiZTdsuz2JQWgMB+jZ3f5lt4S9zb4a1ONnvo
SmUPIW9KxYjYKWIjNhYISlOj/uyKU4IssZ4beyucJL3bijXS53axep1iCYgUxVFjvv8LWlyR29BE
fgaQitoL73CSSJR7jhCr0Ke0wyQy7zQO+7LS6ZO2fe9pziaPm7DhvTNYpiAUc3bJ1rNfU1oQi1VK
/pp8N/YwdhpJrAVGbIMb3a8jQ8AVyDRDRdmfwPRxjpYtTRBzOSoym2Mhq/4uA2bThGn244axjcAX
3xf4AFh2oXZjpGJsHku/8VAhJFTwzBrhDCr97ve1f0eDpRvfy2jqFMp8JRwwA7b32Beun3mIEoBL
0A0/YFEijp74q/mekb4TeaOU6XQDkjnN3uqpen3i5tl5Gza0OiQ40juO9j2ELMJko13egjkgckXX
eDTLH+Z93eZuKTxFwslEI+4oRfsOTL/BeVTpbLJUpsM28c2ISjFiz1kzNDwThf/4/ewnwtlLzXoA
DqkW1pW/pB1giA0DFkeHj3IVmquN3N1Np1c0ppisazLGCSHYs/p0Rm3olkSxxp7LywZQj+sGVQxp
6RJG3N6h0wFJSP18dbhbIVhe79te1kNZGrPsaUmVmcBGz3x2SbMXMR50gs8/Kicaot53cJgOJ0Ic
UwzX/0QDsInqSYhHQ5PBWA3zvZ/w3uqbC9c0kvq1urC/I0V2Ev7a+F1hlwgUnXp8k03Nrn6IcJ/n
YNi/MFkmLQp+leOUcL4ZLTx5mr88buGq7i0NjgHsB1H92LSg2SXU+RrnuxqyyI83tRw+OE8r/xhz
RyabGJ3BGbfNQB+/AiC+1X/vG3kzW+61zXK6Sd+HoW395YUqS7iwn+JXT+Ykddd6R1jQ50+G595t
ulUmvM+E7dNF/5yfLBfh5IcP6YP4AKpefl8QuxFcebE+NojyURFdrJ/5TmWjBOtWqSICAGlwqoKn
a3gMAAUEFXB3pH+hCkOiCAY2xdL5V9J8pOcrVU4qb1dXdc5gJ20/ZXIr/OMlt2qPwzkX3j/PH/l/
zE3OMSBBjnInH4JaV0xApv6O8DOgb4WhRi5vJmHQXSZCuTbz8b16xWbC4N8dV1FcUae2/Il6BpQu
sreuG1ln0U9lwjxF0FzYrovF29ptgTCS/QBqRHYn51zQEQxmj1zm71YLmV3mmBkxdgfZwZcW8FjX
OY1Vwy8vQ4ox0sS/C0qnZEfH8RKM4hg3ENKS7u+0JIiR/epqiOrW5aXExzN2L71awPiONsfit8B+
4xNcRv+gbm0BRGBy6i5cvHGMf+HXExBhEimCJv/XqmVKZOWtDztq2HJIt83LtSx9ZnDXnrhvHh2r
g7TduTquc4td9Cee4kl+F8Bz3WoIaH9990IX3DCuepEqu8ACpC5t5rUs3SpgUYjdbGq2pRq7EpQ5
30TfAXXMo9uUX9zmTM9n/znhge1cUejJEJt1uuzk5oQStV9EHBzICTuueZkx/nrOTFGsAzYVprkQ
2HBbUlqyKdhDEHmN5zQP2MM2z52XKEVLrWeDbOacXyTpgF0sKWRuwaXaN258wIIj+o5Wl8AuxsNz
SbqaZ42mvHnJMqUI3u+pCXHCTW1wp7ewhwL64SwlTteILy4ZvdUhAZSo40M6BNTgPXJ3w3N70DN+
As9qGYHha0e8WrvlpbAOx0aUcESSp+q6kYUh8k1W31ifki4RhOhMQDFxJz33UdrfD3zMlkmbZoUl
Dri3PrqMKq5k1vdXCEE1QeWob3A1xoBIhS5+uq3TXZC+mLW5x85sF+fP6w3Lom3tbCkqadHuaWIz
xk5nYEjzvYTggBV4yCpX0qTozw4Ne1MdPuEbR+xiSwx46jZSxnGhjTziZZtoDauSadswjwiilc1j
d7vP7Z33vSctroGXQ2GGopzqb3HDsrr68nCJclyv9X+/tQXHgR7T5gyT05NmQnaGz3aN4b8yJIOG
lBU6/va3f696QeUQrCcC6wVrhTzghZn4Iiz4qTBKoB/WZgeH2lGi94rekjjHKImXqf5UWP82I44g
asJpYT8TQEE/4u7nCYI7AMOMnaEJ2kIe9nyF8IUDKJ2SNgJnFSXGjFY6O47IMgIl3Ratl32pT3ea
tUb+d15Eq7zIexCPw0QB3wSe6XcBFHvCh+SGVXbCROXhOros+9X0WIS8KcS+ENeWDzW1cZr+6cCJ
wjxdYC8VyQ3EwTA7vypO210Ftp6Q8EAiYMNsyv9RfBnR2nW4i3mUMoEDhWB3AHPoymgLiXPJcId1
aC5NgVcYSDu6b0Cl3tNGeE2AZgJyMgqRU5C5ME751KJY9DZ0tdsL+g7pNodPDZH17kMoIzvCr+0j
OBe7O/7ct0GmyYNe8X1rBeVjkN4tqSvHxhV4mdx07UrQnZCpjwjsyZ2p5A5JIsuBvrrhRW1tRdu7
E2HKlCwt12D+izIO5VpOy4uR130H6PpmyivZvfWWSH1dsuToEfSbmLPGXLbujkS1dQHdfRDA2WYF
WOn2PKWq55fCyXrgxJBAuLSKpdDqZ7ZACBUn8BZJZG0hKk3XAcqeMOBo5QbmbHLX9CVDNXAIRHxg
4axCzMKDkDJv9wHNVkdI33cWywJ2cUHDtwjaPkuBQ7R1sekZj8hIq9mNoJvkQ9G8C4Qg9vN4x2Xd
u6FSyL9UQZtaM8SEBc1wLsl0yyZhC9Q1WqUn3ic6CLWubTVLpcB82zVXe83/bNpwSAtVBMazaTzm
Oo+XTNUsCqiJ6nDw0XEJMfGUC8FdCLBVQGkc/FrKrpCLwJrIOOaOTu99y8VxveuYR7GhPu3O4gcU
O9dfozc1v39RjD0zORq9A3YjqFUrn3aXpdfsPMmt6610sVSGv6GTXajsKvEjI/CgM3Iix5vMz5OI
gPYEodQ96bfK0lnyXdN0HVukDSMxV8qgqno8afCPaCEmybukoZbGl82J08hz989lk7JrXTlgJmgS
Hk9C/J6qgbrIXn2bVJhHyX4Q2zRmB4NwbHiv5ML41Xq5tgVUAyCk+qLxDvlrAVWWYnkBVxfOYeSG
6NymGg6SuhRzuxdcVx7mhHspYyFVktgrIik+9mzeHViNzLNjnRV/XPouq6Y+IVHvjgAn5rRDOxN2
atCj2T8WFEIULZAMRsewZvdI6VafA7EKvPRJIFhmwTILxaJYzo9ayoQb7AzGnf78ol1OCFa73073
uVsGs+E+RWnsz9+rnzjpHoG7gjZmaiD18k8Ofg25wPV1J6aTEb4Sav+F00KY5qMrLz2Sf2MKr2GJ
O+MlyBK8jpE3u9S+fJ6nLgcMzqwbNW5K9qUV6pSDq0EY4XwQhXYwWc0ZS2/Cf6m1QbDdkJZKbG77
bivnrV4XkUlllPjaQequZFPDcTEfRt0vnda6g+XDS7Lgm2Q/zAy+oZ0PULRG7EN28vk18Lxc6kCS
pgKL0gB6xC61AkO9ObNl/IXiX/o2JpuxwDAHRueT39MJOQ1GyVjM1LSdLbK4S4aMhVH84FwWhH8g
3bfYcP3KyGt3H0UWWp4fzrhFNZTXa9pSKvPNYPxxskuvfu/ifdKn/cei9Yl+yumhZdJP9eb8yg2A
VKKAO+EsBs85vcB4Ehtl9sWsegJ7REsJwUkClxx+OkbHaq6r8KMU1vjGACd77VsYTtqX5/jU/8Fk
/xA0gaLXXfC5sUOHLtArvtQutgENVomJXJEiNUD0SQ2GyLiOO9WvqqdXqtqVl3DNvFR7liyqybdg
D5PdonZ4A+lXI0hmgVm1vdT9zaJG3OvJAo8ae5y3qihwBJ0slMVTm1xd2K4pEqo//HyW9i2ywgrl
QmI7W7ARY5VoO+ShoDi6T1KCKap5M6yfcPtDuvG49UtLKcOpQsYfWeOMDu62E7ItDq5gDQM320Pt
VIL+8RUNhgTEXDep9dCChdeiK0jVpiYk2O3WtACuR5hvmDdOmXKc4GZxb2Xm/fRCU/jVwyJHXlt5
ilkkOgRFcwEKTmj6ObOQ1ac7EEHgWJ2lEEoWd7DQQhshUzbdp8w5+C7YU8riYf7EmWyVgvmAewtv
htvdDukIfEWrGzj/dahf3dVLCk/vGHdvjD8igjdQaO3yPJp2TlVub1xGc7rcqqGumZ2wVrpLLrmp
s8CFWoFHqMAR2nExLF7+MHIOKgMglfX3eJazR93BRTX4tz0+caH7ChwztjtTBT1duGt2kInKhuUn
KYP/INNNvZAcsn/vjwuoWH9E5VtMQgXEXiHjtzalL0ugP97qnDv5fQq0NkLuFHi2S23D062rrzLP
fM/K0zVW4BIKy6XU9c7wo4hZsQ9goEWSYzFDE7y1iYglywoOf3OKS2cZzO+HUQAp5iwkLm1ick5X
tpWGK3hQw+e4z8FLV7cka1vqpBkYYGFMHalgfgWN26w062u6q/02vs35ri/6tzVF8HEMlbl0GNyI
WHERqwQ+N8nknQn3v59IRDDtpPS1EDZmfTDXwyizemo/w0z5GoLIXdQfB4kBS0rEw7ggBNZi2hj3
dn7ya9Sc16FHsmzwo2023b9jCVRhZ/+aKXY4G+aWCb9/ByVr6S7FNKQLiKogScgvF03FC+0QU41o
76ZuCD3kovqClesDRt1BLwWAb+ARczHGkNv+qiUnS2RgHS0cHmX0y/VoJZUWp4qo3uFZd32WRqrD
uQI9x/GYZKqVfEyWSKDF5Yn6mWXklnT8IWeD7IvXgTjOj8tLXXw+Kr7MrAK7vs6PwHrIAbvHHM7+
rJZxZOtEs0+AUmqnAhMhkGwuoQnKK5RRcrKNjSUjjqs9xo8Wxi56ReVPAfM4C2M/XwapGguGv244
y9ybTRSVQ6oTsZRyTjKjVMhYRPsCt2jPC0fHJlXyQYadvVP7dgU9ppzUvSn42P8QEf9AV6xOghEv
QF7GogumKAzZ7E3skQeeUM36i1LKSvs1KzDGEFD5WfnRgNnSAe/5RCyBTaENKD56pRhLGH4i0QtJ
YT9eocSb6uPJJBxkIz3U1a4r+D+7t2KEi/4EucQHGjXsKbvJLTyFuxDm2TNuzX43l5KsAvR05Zpq
1PpMFIX1LHBiK8bpJjccVEDKN5zvwASsjL542iJcTSykso+scPKs0hiwmLLBoqAwlIQinLwToyos
zuJTYArf9QhBALqXB8bGKuKGyR8FmVdjyFmuEzrEKPGwP5VGxIaOOx5QJ3EuyiD/I8VL2zM1CkdM
tituiy7wFGsRMuMitF0uMPJetpeVsyCNZEk2CTA/nWugg+H/7/L60ZMyezMPxA3rMlThc09ISQCA
HQkW9tJtMex41AxwzryDGMXTlOm4aDnhlgb8ndFAXd0060IbOOZ+Z+W5mU4Iv/zDmtR+XPZeWEW4
KSEfdp2kJ1rdgdg8ICOHXs73ddGAMesDJwvUBIJOyTGd9Qsen+c1IKkbePgI5A1OeTbZgoYMmgUZ
C8CK8t995eo3gfacBD/fIKlWm1sCy1ZH0nsfiZ+j7zVVRO6pL3TUQ3JL/WzF4mUicJk6Sv2O4HS/
1ayBBwXoilxN0aBX/eXGXHgWgIhuEUFM5qdkEUg1wdF5kjwlnYJp9VtlCtGl3dvwyPbStnF8IHbr
46BOzitglgoFxO5J9H/qj1n9aeVqVCmoFc/CQPptf9TTDhClZ5zB8bJ+h0xjVDc5LcYflSuC0zgq
chB3S1BZZ2/vQzI7/wbQr3w1xsvjmzlTzHvsXFRzpkeCe42fGpgeYHpTp/CVZLRlNBAO/e5iiloN
Uow4TMVtPOgjD6czDqG0GtMU7RDZWruWxJBtSgtGMnGUqOMG7VH3hKZg+IftI5FvD7uDg2EAUkyo
YgZduccJyeLzaakgkZH1BrWR9b4X9kagMRwGn4jdqz7MbBn4FORW6iqhHnkG14jOTJk4MSYFzRUe
q6lQS8gdMR3sNABuJvmECWggGLqrd0+emYT2I4GPKMN2hpHtjFcKqUSX4FsJ3+6wzncecdDryvBT
87P9fGHyYb3D+gNE10H3dacy/KEvuy0yFNRJTwWC0G9EYUyTGlEPE1Oc4Xu9iLBlTap7PjkPdP68
lUsCq+Axqeg3QxJiN74P5Q0YbVyTOJa8HHG0ol2WvwxAUyXPeVwNEIlcvrXpBPB+zoqzoBjcCL2z
1WDQ58UAmEPOtaf7tC7qF1wbRZVfmitq+UXPQRfCOF8dSw/aXTGvH2YxR8bDAeGkX+GtkIgFKAQ9
39/CUiRLU8akZB/zddQsy3wPdOImrCb8M1T5+HsQspSemmG7bG6ILvtSJWjQNENTijDC9PNRqRm5
Qge0GvfZm3TVDPt1VH5bHj8JelAAUHFDxBcnIVgaUd4k2hMbFo4i15bEgAfynyz9IfugJKC6/YN6
ta2uhql+2Uw+ifLOdyAJBeb7zBvp/dmtidJmoRT0kGZOyOGWETSVCE9gkBxB1lAF+gSIdWTyQz5c
n/b6viVGdhpbXoiAoZQ3x7wURpeIq9AnZRBTPwWKXs701gvfnybQIdrgYeFzaAKqRHfpnfMf7R7J
y8p8njIDsko8HPCSU28W05Ve+dQajuYRR1SB4wr+SCj0CMaAxKbiVzXFoctYZRgu+4Rdw3jBYARy
jjanUQWzXEcICwGNZ6tc4mvWSUBxD8d0Ls5LIuS5DAWUPwvc9pKe907TClzQv1ZzgwlWGDkMioS9
AcLH+hvANVot1VPqFzeuw0QnqS5CUid8+b/ZlpxHYHjrJVqawLnzUraayW0KFqR2JYGaGVP5iJl2
degmrJzx0g3mXD767TY3fBCfSmPrCZlNgxEY+ASBsvgFq8q7lovOcxZSnIG9UedgvcBFCETEFAiv
rc/KMhsS0UlnkkQlo3AfZhP88biHZ9v4hXgkURlcRwpRuTT0lrcm+2VhuF5QfMSRiw3EJYuLgJAE
Tw3QjWxYqi0tPs87VvyHvbJD/BEGOzJrx1FATHrMpetEGhTQDMU1ydnYdseemvg+n6trvy0GbXqk
XaMORJwooTdOfhvNIJoV6BQ6yYhgmdIYFMKYtNFWUPwQxV6OG/UVcwajiqDWlW7JaggRkVh9GnLo
0pnf3WaHXW2eXVwjeRI89HMzStjIlyn+qjDL/VfRdKnhsZjSqwnWplRy44SxDIv3IQ32ZWRurF2S
WLR6Ok8PyRg9pCmWK7zWnwu00o3YyQXISuZ58DYVwPo1gnSa/F+9EFKiajtpE3mov2ugzWRcFjHR
f0/B7JaRdXu1ZI3huQoUjp3i8CEt7+YhD7r1yUWrbIuURvxz18cufph9oEtYBFhDhL5NLW9LWmjO
/Hubq8iioenpJN306t1NYNzBzMJDmOV5gSpXQnoZcYuU9rx82IRhhxifI3C+Uxo1ravOBrBWpYMe
t+ziJ1GMbVIcpg/7/AO4jfIHWpC6qAmf5D0WSkuaay17CoOCy3SVILFsWdqm970B6owrN83OT22I
2hYvGCLZIy5Zyj2tysSrmZ9oxJ5BnaobskLWRTa7C6lEx9ME+4mbzs1Ag5zwhJZXjRXccb616XFQ
7wZZkcGTiuE9McpPPu4UVyGpTNoyOKD7YNhhM7Bko7+ZyLIgJTYNgqcYReYTTz8ssh/ZqRO3O/V9
VQeLPw9Enyn91bdH89+KokOUqlSUIYFDQcZ0Sl8KrBgSTFIkM34TI1tWdI8h4EOMkXVST4IOs+S9
4busjLpOndWAEQTGKtoEqyc8mnlOPoBFwfXIGbHy7ms2WjMNmXSIIccRyARCIH0JvacsVwmWrYCP
JvxtENo8KrgHMMgoE5xe2exiQMf9pBZtodMTWPtN1hnY5ApTtSRTX92KlzpBsfRv9tiFmfo71tG2
Hy/jlYrR5AKDapM8P2eSs692KXjzVfgNIwcifiKOdFfQKYhfrNMJ8ga71jB4m6dojzFhgCm/sZBU
6YFM98sMRMsXUr48k2ttgnJ795crjICBSZg67avmAnwiEWWfkLmVMt/l765Lem1Vb1lLZDORAg+r
nKAgqWy1zeHjC69nsSb0l/6Rv3BYQ0/ob5wV4AIlhonv0d09VjEoXu/S9x8mpu9nM36WvZWZ9N8D
1AV6LiCZ3H00H1bY97Xg7PpBCBDeeb80Biqr7HBgN3rZmQ5KnFhqW3WsUI36eoyXsafY9CmZBA0F
+mmKcgyC8MpREP7ulMmv/sFqJ1xdI5HQT/gbd8jz8ryal1bIJxKt0YP0EHah7rzGWSXQe2B27M6r
OUffqbe+XO1jd+v19MCedZIdRzSGc9xqtzlGRhnZtsutHkxap897slg80H1EMESchBKODR6TFSz5
oSwwtr93yqY3KtcZaBHkzJMrFrWDMyh3aeC5hs3bWR5EQVS9XQqzRtYHRznAoDv1fYl5oRVOXdZH
kUtloHIWXbg0DV7qCftIUD4Tv0HqeFvjykAcvWbTbepT1gE21nBJMBlAvdCBhNgxwTVbeN7WdQc4
ZC4wyLjjve8U1sjKWoGQEaCM1wxkU7V7T64XEcTWX4ZVqWtdiQ1GufyOjY4Lb73sgGOnkwAe3IQt
jZov7Yw1wQ6G6xspLOqnHfYQGDeI7fYCa5hsbULEjH4JqDTbujzx9WnZv8KGEtA2H+o9naonp9BF
yQW+pqQNZOWiQa1fmmAAYyBviJIETC01v2sOWYb/95/3zxCvG7kb0vPX/imhSh7+Y3U9ee1PdHfR
yiTql2gCIp0U7ud1tW2DADQzIipt8cDZEhpKJZku1xbVVp7Iom839WFmkj3A0WAPH2MDqrM17f8u
6qcl9BG4vdbDrfo2GW8RukXGyNdl+qyrsvdYFmVtbMH67Jb9FEUuDo+me0rcwmlxV8rlumkXcIwX
kp7RV9Tz2UxnnctqHeW8YWQT9XxfJKhc6h+e2C/17GrzLfOvSVhn/QOsiadVaosotJmEATshDKCL
Thfp0b52icj89xf/QfuyJb3a+biploe+zwdcWc/bAmEDwcXQg+f1hRCvsSDFcJToRmDjShehc80Z
hpNlUmoIKydJ2U1rDO63kxM/PjsqBXbPaRnrgHlqudpdsPBLCJK4ZlJgKdNX+CQHfCvwFXI5+6ae
5vdY/BdTCRB82EKYKb5ksXTBqhdG5WCTHY1lSq7RMEFRSvT8AvS9VHaZnMXaBBIPO2OpCnVFNMsj
geF41JeAqqTTcuFkTXYroA+t/lHq1ATtaTMVMcjnTyI7lLQunt4KAUxGWmXSt3yHXFxicOEVwaIs
OVxozHkTLjHnVd8n5sXymAdZfdXhAJeM7rYPEPYJhI8buTD8J0Gl96E33UqMq6q67XLF2n36sNe3
c0Ii3nl/9ydE2l5fzb1IPnu4M/h2VF44tAScI+G1lliZe/Uj16Kqyad7eTN3FjiK0LF6Y1mvAy2q
su9Fz9+OTrhDHpxzs/KHCqP5h0ehsH2rzhXR3N6+6OxldcC1R7Wuh1G4l+5tShbBV5OkRw4/B1e5
o7ZowTdC1XX7fIlv6oZk6eu75sRuTXq+u2mA4CQ8QZplIUfTL3daTBfpRsrO4OC7uoD/wVvw9Qta
ToVLl3+Xv417Fq5bFwwCjvWAbprKJAXWPfSKLhRtztN8q4nSljQor9+SOnJhVTEUCuqj35OtB4Xs
HCCjACW/RJZ6AMJeWmwV4K1YzFcYK7AWsYqE0CosSSLQ8HfEHKPBxTb78awYyqq/4l/bCB9g73jg
afV+pZbnMw8/07ki4E6K6+rEzg1+f4PReuUIsDXfaRSeiDZeEUp3WbTSPhPlypJhmq2OeCVf3mQV
gAyD+FobgiHrvjcBi1Bt1r92opA7sAW30UShARWT3upEe9KGj85MWOAvtAhsXQI1j1WNGv7PovQo
dtVDc13c2pQYct8R2j5UoCNJcJ4OjsS2COSsg4r6pl7CQJbVGdp+kzlht5MXrSaVPIQ4rfk4QKT5
1zYWiCqwvsBb48kx2Ab3Zv9CcrFFvZPv3dfRyYA8gS51BCXj3Oi+jEm2i3TrvOffGZsCdyJ4C+iZ
sQBFCdya5DXkGiSp3h7bjLyeBEW2d2/w4kfGHBBxYnjoPtxTla1at+C1i6YMnuZ8W0Yp+d/d7xOL
DMVELPris/1Btzrp+sT4QCcRcfIf3+XiYO4NpV5/Ufwo3D4czT7zxBr1fXqEJy/H8CmhHCj4Xyw2
8GvSywyR0Nt0lHhTp64gXKNsTlcfD3ifFfiXPqOCzXqja80egFHfY45pafqycNkaa71yKGx1ExQT
r6RwzqNn/fZzj/skdaTL5bjLfdXP/2SzjwE8O9nUZXUt0fQrhtP/HA1OsmJBKKSCCTE0WhXkIA0g
Yaz3w5cyEEELUcaSsR2c28qpMKQgn2OhyP834otHRSGScu73TNfDITmpJYXw6jPM84HuJMMYhUEb
ZruNh0HR9rdw6Ekn7f6fMTdtFoHwSAIqYv2H2GOVfiZuxiB3bt8t7A/gg+qHzeXPZ2lDlO0mDpkS
u2BcRUkFMeCBRewWRyJqPfzHZb+8R0CTYE7OHFuPsFXr84CMvrNfvH7pfy+6nll1RijAM62L2dGq
4AMf/tSOOSQ3tdc2mrr/8YOjIjww6VKJ3cmNduw5iWB3+bxpenR1o5nglsQIFK+rM0Mz5vjBhFqk
+bSFPRaoyD33zn3QK9JaEJsWgdnfDoxwsvVl+hfJqHUJaZojY43rMyYm0hecg/n1XCj3qsmmgrVF
0dum/V2JW6k32rUzQUfLqcVCy0p0EBuGe+rjr/3DLGNkMnxG6qnmzjSXloVvU1Latrwxt095VK0m
E9GjsyFypo4QKWsTBa3W4mrQJcEVfevnju1wdbl00O1KS25Z4m4eelpBSQhEY3PvSwAP3MupFnX2
MyyfaKhs2vXV4Fl2VtG5lKli/FBzPCYluZ0Ml8mHPZMfYkgYpZPUERfJp2rpy3MOUm/LaxQvYwf4
5v55lAn0TczyJb3dUq0A7aik2sZa//oq7ry06Nd9KPWWv16xZb24nEwdgupATqAKM/o/MsRFSbd5
MCL6QrWFi/ibRo77cSp9ZEN/tYEcXWxAOCQO2idqc7/XsJIEnOSjM5AtTCCHbmK2SlEGa8PUgkQV
0SX9/8MDaYxTsC4C7FlTblpvo4Upniu9mAy+DU7VqFo6W4VmvLql+BGNsQxNdkM21TpNDpEG8uen
73+ZIBw5r0Bbh1oSgC9rRujAEYRAs9QgwKcE1A4+I+HZ1VAPgd2tlZ20Zo3HAcMXADlWfNSvGvfz
Wud+H6lQqR+lmVqmnacAwdww9ENubJTsRQBAHxd+9ly65YeqK7xEMn8gWuwtOiVqe6vjttvM/mKp
TuXgzf4Cps0k/xza7NOXjeudWj8o+UJrSU94LxSX5SINFizTVeQNUlROeHWEtM/3KApo5BD8hiYr
7xYl13EMYy3tgltCCvaWtTjcZMjHIWVi4USt6CZwaumNumFlQ42leW3mZU06FPFvrxafqC7ZAebO
vCJmKaFSv3l/kOms+RnwYPytq7v4yZWADOxgyf5QNIMfgi4Tz3JxGgOfRCCU1mn8X71ZJh6EZuad
ktWpPr+r3K8rSKEp8nkw2rjSoiowioyXznwq+DqC8n9Rs3LvfhsfYmBiJ1qoTC+XW5HuNGih7dAA
nJgd2cac70pYsH2iMGJP1SM02VkNYfMErlxwy1anvi1hS7zdWl89tNDkoLk8XBM7XbYwcIY/nrey
97VNpNwZZngXILe8TZe6rcM9RVR96x51pMR5sFrwqaUtkdLgO4epQW+dMXc6mJ+7jxUxJACGztf1
zIgAtLcF9lCIEkt6/f2Aqygu8vZOPYbuhLIXf0RC+OLdBhZPc7b0F0vSVLj31btygq2L/ZrNL+XC
AWrO/z/hyQRaxyZ+9dYSZNX9PN1/sgZsA78THOIRCJqV3gNQjyRuKzelRE5ON8bzaUBvb06zH3hH
Y9/LS9ItHlD1k8SOKR8i/108KKZ5EKzc4/qD58bTznWazHdpvTKlpqKJNfplnWLyStKDVHJRewSj
uCgxtZnKOl6RATP++lQ5afxbXfBz8u5bsMpGHauldx7EeJ3LHgpiuOJgPv5uNBJAQFHJ/FOpWLhU
egLwvB7Tiunfz8mRsIP0KdQfwY/5S1OnOuLPmFA/3W5Ab9gjDmdyxJzRR3G8YzY7zbzsBX6CUyGR
vUsPo2nNvZoBtTbehME+zWt/Jj6xNC+NFCXgxdYfZx+kCpybxfay0QYfAn6uvvsEjniL25pB2+S1
Y3rKNtJAeN0BxVYkjfm6QMKijxWjqHAszy0tBTwPiphTvR6SACjxO+8bcSgP7bDo2fiR/IejUw2a
NiFH8yMWBM+P/9HnEMtlT/9ebXQUxcxEM1bEAmLr2FA9xwYv6Xi9/Bz6JqBSbpe8ngiesH6u8Sys
QMoWc9ATIk8EHJqK2Dyzwy3JEvAU7toqyrXZii277UHRITGSULr5xOCJ6QRYdDDeAOe0Flettuy0
dYEtuAuAP7ausqhJIFrszpLrSxaWeDrWU780+UNO0TO7Z4d71Bs5lIc1/xzDR8SZ4D05C5fObOYC
l3z0FRU2ymtb2gJuBQUP+5Oi0qFFeK04kDLEGeTFipDbRtQeZqOlZsyp1guDbsvZbgbFd8nAy0YH
BTJxIZY0fSZ1OQuoyaZ6FmfvEQNuuICDf0HCQH0pHMe03IjDrHtbE/a6uPj9M5bLQpKjvpTrhXAP
dgybf26CB/OfBrSG6oEJdSuBh6UhPsAv5PxlsKTXmF348qD+OyLxvo76r3zIxfc1m2nLMmHEHgRr
CeEu3COV8ERD1eJxb26ranUHgBPWH7PRyXa2IbmF64UtgTq1XCG1clZhpgps8EiHOL3+hlVRsFSH
tCMWTzf4UqAknuPiS/jvXI+1MmstTvkEwsOb/i6zjm8HSvskR16EnRBNHRwLAcjTnIFXDg9XqFyX
uE6OOABtEoJl5OJXJ3LIUNIwFny3WCFjq+QJeYbPdLou8fdpEq2JMFJeOX6OChnlozsRqEPCldoA
YASBjrZpNK/E6k+o3I1AvFmGkVoBokmjdjdVhRaycS+ETKf0TGrwLbcNQth1V+jNPOWKeFyCzN8H
lramDNeDRz/ud3p0zW6ng0T5ULGCBm9zU5KB1HKiOS9N0C8HfU6JOvbib8DBpmJHCnu6fxFnrY4z
uM1HWF6kD9VFqSo0+Ia+qOMQL1kEY5D+A6MFE9SY3/YnkNcZ/lhrbFO4TG7qdvcLDZwBtN4TK3Mv
jUMsQXmlarLikCZYPqQWchcFNljNJN9XAYg0ZZbOScVNa0zxwp+7fH+q9XGTGQp2C85dSs/wrPzx
K06uQI2ZcsRbrt2bgnaf0Y1KJwx4g5svqSYrX59ef8qnYm3Pqt2ZXhndmpi4SefzczihXpK2WtZj
lspkA+Wl7gsvs8ANvdIEAo2NJuKSRwDEIxRcBQ3HIxY1ZDjfLZgq92v8W9ujzzM38hSVDNL5a3cw
ym47ObMybr++0Fym6/l1tCOQ8vq3qKU4elZnY4FLUp4/UcveJjS9NFLJaFqGTe6bkx021k5iS0j4
J+gAGznh3uO8CSLRVlboyrbUshpexHn6FV5CY2t2UkvpBFOqqVfEsP4DPMYUlBzUVynM0f03PiBi
bstbzVMZVWAv7xZMiuvgQ8B77f9XMZY+mgz+liar+U3KOevzZ9ahfX7PMtaYweVpFPk7noBJf3vU
Gwb3uHzy84MPtaO/BckpHi90QrlfFtQlL3NK3qx2y8R9EglqicI/bOqhRbKvjRSvzaBpbigGEUiC
QdLqysPz6wThMHj5BJvUcuUZpnmrwkbkoE2LyrmtDUCqKwxTGBSQDMhQeoHRuL7cJLYASNk//2NP
P8NMy6WHvP8Y1agLe0Nf6zs+t3flOWf7j6yRK4CEV6L8x+NBP1wLGMJrl5vC3mFVxvO3dxn++/Rm
fQG7Yeg4l35wzFnR+MFoFYqH8tRwZtWbjWYEJ3jQG1EaU7Vg/JH7VMxbyUn8lICdAmLjZFo7YqES
xw0qWY1Xk9PPpoZtbdHu1BtuzKjU0pM0hGUIHfcwhTRZlyv6Q7D67tRRx9Y8hmqtFrbe2CgoOWBr
oVdfNh3tkyoSnStiV82CYQxbX7w2TjGawJQdKw/LLr75qa5a/Z0GncI1VSdT9qih/WG/Gq79qhOG
EBJM+wV4x2ddd9xnEFtSbig7pHdEIejnDVMRPcjZg6nIDOwhsGU/qYB7/ef1DqRkYNCrgj5woWbf
lcouMyx4CEKH7N2FXlvQtrZMV4RyLknHkI+JxmZRDanSpjL7FnVXMFEBeVn9SyPciX+oiZW5wgvI
K6J7hkDUYnEpBz8gheEjHWhGKsjuSqmwJvlkEY5R9gLY2ZrWe+lvP2Dpn+SkTYPAVwehOyZAr6k3
55CSXF91s1ZHLjwFP978vPIVe0ZI7xSvlT7iis/sxzTkO0RhQHIKIJ/8tavAmV1pTZj5BRoulrJQ
sT61Cy/+0Ddvxr74TDSzk4VVuRtGSGqMdcqfsKluE68rTA/fKQG1CXh60a5GKID3p6nKOTCTsbNv
nrQQK/3KQMrzaLFTLXBSD8EniosI2RKCCFzMm7t+BQvBW1wE6hVsLN89XHgfxH6Ynm5pY2JNxkuR
XW/3M0W/LfcUhe95swyEwQQhQqufU2gY4vfmceTVvt+69Scw0cbvwiOR0RQNg4y+sSAHL9TTXySN
FvqBxSZR8DPKlgiFfaZBq+VlC7hVp/+QXG7w3kbV0iMtkOCZ0AmHKT4EdbweTr0v8UbhlkuKAvwr
EW6NvolJldb8R8BZcvpo2xUhV4TyijLfkHfH/iygEG6MD7dHrdQSxeRly+iRSUtdYfpS+qDDQizT
6u1ms3yN61u45LZrDCcxqxo7OukNAXlCJrTMbWl0uQEGmkuszhctU79qUG8IfhdDTSFjG8RMznaq
0saKCb/ZHeqlNHyxdXWoo2ZmrsSnbwoS0HB6sq8PjE74w7SFRrw6eeFpwgSVwyBKKXmowBZ+41n6
GiGSy43hvM99SHPTArhztyS6bpa7EG0Ovcs9iDBaaxaNasyp9+1p1PEpEzsXbuj1XPEZ58bl7QDR
9xpfgKRLtCAB8dKm/Xu2TkNvm+q7a2+Wbi1Q9ZTpcTwqJqDd5kUsroYUd361zoaqlQ4FHgkdCvda
mqENWFx0JZEZ571hBHB09JjTx79HOv+RITlR0NH3FLS/DoKz+MNG+alFk2izNm1V5Turf4tBAL1n
wASaFOJJB10583SGHAoCXlp6yrWQYJvSodgrbYz0EXzvH3C0woc57L8noJ8brzOo25GUlikO8pzm
KisCpFMuFZ1ltBjUBAA4wbim1ijl+qKL+wNB3YwEIPf6aFInyECpIZX9IG0fEyyS9elaQXQ+Qixi
SztTZ7hY6KkiFL1spRNAlU1dkL+vcIEV8IYFY4Em6ticZzxa5HMo5xHvaeSmC6DzkH/iiu7H2V9v
FiFn8EvGu0C0w6nkRSBQNXWaFC1RA0Oa9Vses8VTH/N5vv9nRJfHdGemsRgqPRasbSMDNG+zW+Gf
nv8Y6wp9z4FpVKeMMjjFgUlO85NZvAnB/A8OOhE5DDPdEsKPaPaoFXNGKpu1jCdVEUwvYa8F+NVk
Ol0XnKAB8uMMXVp/wd2yJScjWZ+ZiKPfmRLqRmkzKkXMFXGTDZ0OkKLQyfAssb8n5EjRA7j8gPU2
EsVYxfyuGwl3t7LLrLaMFCMsopAaD/ZSFDqHEHmyF2oosVypVfCxWCkRHdqQvPabcPRmKAOyoyM1
HOt+j3tpta40cH5Wnqvl0kBzBa7dxsnHC0JP80aDEB9LVc04CndilOvjKwDhtvmRPIJAS0+3mqNK
VMZcVJUI4Ih/H8LqXZYDmS/lQadMCWqYhWI2zXlC4zbEzsYLX5PgiSs0KpmbCU/n7AAimpSFqyCG
ydgifSuWaZ0Fqvo8JYFqza382RBPOjS0ueXlbkbsBkwzWnL5WUQrCdrmMLhU4azoHgZ4ACSosb2I
irT36jnZ+hXwysMFudAiD7ZPjIIOc1GxfCpX3CAWKQO9M2J69WZh6qDJGQjuZ1qKAgKS/l1B/xrS
a8IMXsMkBWvgGMxkaOk7E6U2QeJ3u0lExheFuq/9vpO5fcreJwbkmJQxmlNCqFZlBqiKmnQzmaKd
WnBk1ljgFFJVmIZ+54nuQOKIyKAtqeGMyNImpZAVlzN3KCHVybl0ls1d48zvyHBRU098cC7Tki5c
owdDijvDzM2S1bpVxvrEeJf9W+0NB0tm/lh9kfIlUhumbapHa3uwo34EFODduZa8KuwrC3V12jH/
oPfOQAADhu2AwmqkNIY48u1EuDZREpF2vqmWSmRYgnEvYDG6TiL0M6BL8pYbSZq4sf4reZApiIhl
3f6EDZq3s2TvzDhbnQcmH477Y19Kwwev4fzfPmdHZJDweaMlcPoDGFia0inRpPG6xDs6oSyUyz8Q
CRyQ8h8hYw3X+ZolzUKRQ/UjSb9t1J5v+anlPmshHDuai8ZyPDvU8MWXbZ5UfWnOtroxxpBFYwK5
gBYkgIT7bz7uQM5WkC8NJtnIyXigMDl0doRe6OrkbvH9BxvrKWKJl62PYO1iajVQSahEnJb90CP/
bTFRcw4MA6yRILleHykmEBKAI+SfUC2jyknvdlpKZT7fy82FGK0K7UUtZga98gCk+G6MZ2SMUUJZ
ybmVQEpftg7rgbUCiFKaDaf3r5sC9aZFekbNOU+Ezv2k1Aii8jI3iGwxl8dMpLYZKG3lqlrANj1s
3aaOQDRePaEjNaMhVRJYed8r60AIZqekYldmskyIVSH9vR2pdZoMhb6VunOU11Z5YqnU1uth3HdN
frTLT2/yh99QRSf05yM8buWvGvtq/uy25yfK4lQQkCUnbuAczo160pZGIDadUy+nxLtfqex1KsqN
vQwbG5j5wF2GFxztmInnZaZFFqOprodmczDGWjYxC1vcezK8RDU+qLWOoGrJ48NWZFEKLtNXo5i5
mPID/Y3P5fqy2hkPnRix2bZTYkE+SJH/IMK9zuwQV7lq/8athId0XDHUaWlFiGBhXjkTvfM3eKPm
5Xp14IwjrCIwHWTVAo3U5zxkakwVmgHwYxKyyYVzwfthr4q3tUb0IPd7t5cexYikySqkDuL29ZUO
YJdXORCIyN4lX5mb/8d/NpIfCtrPz+bt4uxTd5OwncpcT2hpY4RWeioaew2lTaQuvVo2584hlEtr
I/rSpBD5uwJmF1dxR192eaXZMHXHT7cwWdh/QxVRtdcqJaRApBABwdHAS7lxT6Qo7ZY2U5WTRauM
B9jUL/GXEIggq6pJ3lEV3QgbEB37/4ziPQvkBWaHErm3mNZu61ujYbky9f061XAAb2zyDB8kleDZ
Mv9K1dhwSyOK4fi0UvbZ4S6GEw3hJ2EUJbDagnrKVzVPNxzF4X6qVR81RX++5ko+rHh+NIdaZEiy
hpK1swchZR1m4TDvNb4Ip+ZjvKje3/YLEjwg9ixA3NvNU+SreCKCfBYox//DRQfo9d+EhyujKmZN
930vbkWgwRbqVRdavG+tnJXUkxcIgFyzykQpA5DBCOfJxGT36ICA3wdyvSa2G8bsBDBkePP+k3Yr
y14e/UF158tFWeoZ5353K+x49Q1XtI5Wg45gC/GtR9XL0eUS6to7K7mnO28c9cEIi98IJveQgflP
dJxf4eDRilTsc1ziTzFxpGn9z8oF6mRlnUPt2+Nf14Gxp0F+VKECuNqzKv+yBvDwfmo1bM5G1ofl
fD8ZeV9ho1bGKWm53qKirzBwHGqdsBxYTOO/Oi4MURalSzhR4ytu4IF88k6DwzXfgL0VMTMADw8E
+rgPcXdnSAKRCUBWj7tPg4ec0Yb8598IbBfz8ky3AJ0sv4FRzob04I6PDWEFQSWnR0IB/bUsxcop
c9dx83PR/x5jhcozSQZ2Qysz2b7xV5BaTPHvQ0ly+VAdxHE/Sk8aJC6gjAozF6dkYzNBbwFKhoqy
d9WbJoRJxWqKKviYtC20YrqvSQUQ60LE63AMiVIIQkREnROSjdJREdpiSkkpAZd1DKKMDfDgpn3q
EBvbFhlg9hk8YF5PqdlbSKs367HGXfLXE2ZYSAB5QMHxL3CVuyLJ4nndjZaBgiIu8NWHl3v02Dlw
lyyoh+sIa04dkfIOVbB3AsOTBhAFASGVd3sZymXh1zA9W52NqvTSCFSzvba/wdjJo5J4DoXzx92g
ud4bVUwVF0j4tgnKfqAscFrj9K4UHV6C+/OczEr6O/AVQs6PLBvvyJV609t6zCk+cSnbLWIbdjtV
S8ZZW12G8jwct3CVEbsjh5PgrYIiXsFe3/C3RLHx9hMN9t81Mnsxv6KVjJo3636wFtq3EQwRtoFK
66xIoROBq7MmSyaHTB8/gbxkYqd3wYmW2kHCF1XqrdlH+1nAVJPz7W/y7LgBBtY6VB5/jZDWdtsk
D7Jc98ida9vx45qeGlF7dppcwPkW7XzHf+LmYgYhhIzop2FW19+nAptf93KvYkpWFVyW+6e/I2Xs
xP/hN7iVicUKDGJBgIqM8Klu8U8bmofsasMFPHsHgm337j0X/Zy2t2daDBqmBFUUM67D1h9cA9m0
DqSUpCCoAF1XzdZfnHeCO+QYD1iBt0vFJgl/M6q9jTd6gAG3bwZj3QqBasRUKGRKmHMJs8asLOlk
0p4HLSP2h3FVR+wi9eHcNVkc0p9j8i1lSNRZN23sStAkR2IDSp8yasiEWD5DS62nuzeSFcnwl0PQ
elxITErWlMqlFo7CkHfRRKahnDs6UMWJJEWNsSNxYKuXaTgaZRltrwY8mEl8igY9riZQWxk2XVwl
gzs01Pp9PM5YeXWYHwdVUm+l7YbEK+C7JcPl0bH4cGm+MXuQ9cJv+VBNgyl+1MC1C6w0k7vRSPLd
rQq3eBRMZvmlL5egVUdQ2JQRwyns+uGgiQIhDsZqCp8Zt3YEx28HsxeFDKtcf4njTR4wwb++xPGl
+gUb7DzTsr0d4kdA9xArWBkUfEnYI5xHvf0BtqLH9VDoZifGHs87Tj+48xOcql14UVfhOr8rLa3U
TQN5pBPdE1qWJl7Jpen4C30CNeq/m5u7HtBlpJh7kxLmcVZiJC4MuzOLPXIKzLdP00qcYeCuGlQt
nZU88B/08vRk4R+g/RX8o4OTPBPQNdrmehv/zfABAj7mopBG8uj3eRNbT0+WjkMYZ9H8/n7IkMwe
j4FDCkCwlFNlCRJoXWmxMwlh0gDG94yTx332cxMZ/2/AFCNr+xg0hGQ21RWI5nf99+mLFtBxm3iU
JZgKoE/MPOy9uKNw3ombB1VQ2QB/BleSCH7bPsg2CEX73YPSttfE6bF4cFsg1V47lfBcbbTJXFBT
sBljrZzlfip7dCU0NiWk8oH+jkmrYXa27gxrd+sdxRYxOziUq/mjzlaa6DJ6LrbmnFUSBjXcVbq1
yM4b/CN0ngt7bh884l8lds+5GRhIYR0YpdpE9oqnnbG7Nf5YXkK3sZ8y49QMAO1UZLlj9HuxxDlz
hgoNF/Nmn03PJc7YXn9FeKI4MUNCppnYKaInSycfPN1ZP/XZbUKWp4nXdokR/5sUaPtoHDjQguCD
ItcNzyuy4suPEhZeqJuSjN5a5J1n69sxvjGIhzDn67zuFavKpphnoIZ/6BL8OMgOQX1Ji36WhFLJ
2P1pAIkh2+Q48anqsa02+s/FR+cZdMv8yP8AjXkXuKHi8RKY/CGu1ZfmTrIcAvAXEggQQKcaOANE
apYn6NrYvcyy7ah6vxAMk3PdKtbjFwC9+AA6WfpT8p2exyePtg9V7POb9WUHWOj6eAkE6CcbDNTh
Ou1pFuChBocspV3mPV+M0dgi7iQ1fFdb2BJXtiOkAfJxwNOiNztb5QaGAsQ4grIHZe/xcV+5jQrW
cAEX2ptXD46RSRWsgf1bbRGD0DsnVzdzN7+FEpath1icTwIXVS3R4ef+aKPjEHtgBKh3wTSUOdz/
e4aeVSWvkHCWtAt/KfbyyHFsgDR+Jt7W6SdZOQ6ak3WHlpXZO590joopLGCJxD0agkbIIniOBGhQ
rRN91CVO9JvHuX64aMYPQuOmSFpWKeRxb3nI1t+4E5roRjK9SAX9qmt9puUp6y00uowJF+zi2NcK
g2iiiu5Ncwt/L2Ev21Wmx20Eh43JaTkCWDk6vUnhtVWxF56nPpAx2QcpPGKY+kGgOuSCUv/mot9y
DSDsNgmx3xME/HwpYbpJs4cHZFOlWx6z9RBOp9Jw7vKSuYvaMil8ge/RUbzXBwKoBmwxpPbX9h5t
aLYy0Urk4epTKHKd5fhq+7QWSJ2/o0biMioqSOrC+kQI+t1vut0YzThssTEgDvwbb0N1fgs7EvGr
Ql+NdAINJ7oeo3pH0TKTeXR2/MwALHGByjj8/ObWGcSz16oX841DQzJrVli9GX337cM/2Ch8cY/L
hLEo3b3IvDmXNuN5qNopFg/5ptEorTRgqrJUASP1ez73CnCcHOiAVU9TN/eqyjV0yzPa+WnKR/4V
MTNcK31FUmkQ/uWvB2yL2qtIk9ZsnkhC6BBT+Ja0t5/mRagOl7isYeFWUqPBupLdNIOi3O+TavXa
g24PfrgY1f+G9m6o+l0WKjk3T0Xa5gvb+EjORhiCJolhsHTWUTPrnmjaoDtkr831zBm4sYKks01W
0zCCQWPUEmvKmkBOFjU9lTkSjBqpacB8lgqSiaEtlV0RalZndsxvtGsFHX3ot07mynfjtKYdh2Z3
rtT76mbzM1v3nO1CojJ7SiTlhqftvN8uiYWa7wWIB3Jm0sSw/SImLAyndZDOSKJoWyXbmpoXZOGF
sWOBtnDOIxUy5WAz31oVEuybqGjfunvIJKLURahR7HuBlqYJzWgRlNbRifE1P4kw8XiBNTk91+AF
dXLpY9VqRGT7rfJMrIUyW/LH4JS9bKSQ6odkW7ReW673VETJoMD/9PmZCf/M6V8jC7sYBpQ5Zaye
AKU4f3e8O7Gcl5pUCexRm53i9gqiiUyMn5Qa3x1RVQJAPcy56wOW9g0RztuI8pwxwKuktbGHt8bT
GbjeKSFjJPVKt7B4fS3KfY+bn1jBFmAVTfkXx4ve4TUSWsD7JA9bQHDKZBoWjCrCEiccUrffDI/t
NuTTAsMlc/I0/oWF7JIDFGm5fMLmCJBaU28TNKaIX1TY/CEDQuEG/M88I96aCDeEfmvGyS6fvkql
c2vMJNsgAuQ54Je+isARd2tZORJGC1bx58h+tsWqEfkEMbae3BetAscyuldOAs15Gn7yUxMGvy4q
z/VPP5mV/fwklYKdGeZQ0MrrKKwOuHnWuACRpp62uswbWKoTnz5Ammui3wFtfr3BvZed8YfaKkIg
IRg1cnusKiNbhgf/m8NC+bemlDTP4jLSkwyxjJzpw8jKipv4/eN7J9uTKuB4g+hm/hAi3r+Br0NL
OLqAmqzg3FX1hZ9HKgk/829+jtCGQPztIsobvwX5l0G1Nrq/ijbZHMCgkRHR/F8/Jd5YKLqSzuV8
CMFRRT64TWoiQ0XzD5aS0x9sVQLiop1MSXnDZuVV+igVIdc07eO/YCFaJpQPRgECww3HaHTaViQj
DXPdcO1zEm8doVTWhdsIN3QfV2SH53Myf3cIOjO0JdN0H6jC2apn+kE/CQSygyLfLs+fSpTqP9jC
io00WwhSujXxPnjXKnThlV4RB5znGmEk0/hlXWnVXIu/MLkQfnnQcfRS8RNOULOCeeqBR3PDB9G6
ge8DmJEKXF165CPJiLeQxYVvvQagsg+MeM038jG+ANoj4pA7vCl+d7lTBJZgNX04JATpnbNhzW8f
O4syKsJzyi9ahnhp9nnzlsZsg6hZ+1hSLGNeQi9bceYnPOnH4TVSExXFdfRF/caYB5l1tMp3lR4O
nOry+N1lMloO9YaCBqweuI/bunFiMOmQlZg4EdDaVup3+WfmtM9biXP/HVWvxljbb91MeuEhapDH
nyhVgC7UUxz7O5ZsQCnyxhOo6udE82RDiZE2sYSvrZweLDEatqBpRDVzZMnsQNdJlSsTqEs5jJu0
zerBJe9K7LrMDInudW8tktgr/jXp0TIypDObimH3BCgC3F+dqjlHB4hcbiRUQ/S1wsgOd2VhLl8S
YDrDJsp4gITaBcr5opeanCG9+qx/xM103gzXCb8ZggwWDayUs/SZRX5XjHE8EMGM2J/+Ru0HrhD8
12DTGhdPNzNKQpX33TjItfX7cZtKzkjh7n08CpbQbospfuJOQipVYUrzLYjG3WVyjgccvkrmbznT
dFpC5KdITyoUHICkbnWCgbsTggjwF71kro7CNkM6SXqVD2rTMaV/kVhRH2tCip+vtgFmMm5eoEin
oc6D9bytacuvYuwAevynPUXUCGrQGgVSBoDV1kiUFVeAvu7WuzKV0X5xYiW/N+hhUxYAZV6UymoL
ou5puaTGalTOITctxugguknsPwYuQF8/HekfFe2oIEKKhytdDP58Fjsw3MsZJre4xcUxSKhrkZ++
H0DApzOkLGGpr3asUw377ytg+7uqiOhBLYwyzcQPjn3AC+Qx4cbqolRPTxmDLXcTJvnqOPKMlLEB
P74Yj1NpQG/uZPdC2hSCsneJ63bvwOk/D+fc8BstYzCuHzOW55YmHQCdg6EWpCL1/roYWp3HGwMz
Eih+YBASIWm1fPqA8cGPWyR+lA5ODSa8k9g8U7kHp/AbSNi3IarJ1wpgdiHBJEuz3wtnMGKttDAh
0WUUM3eR0mQKAhQUi4IXW8YMfLbD6YzB8FjxeJeWSDAPknRT977CHtFIMyAmCmBEcmUxTxwXznq0
LbqHPimeGKshCzmrQ18CIg8EJ+Xf5ytq5aDRSkHaJjv17KBezD5G3pPjz7CY+MqBnIWBhbJQ8j3z
uJUZpbyndEiz+1eUrankenE1Y5BoxwYAYQmz0UqmJepmCMa+L8NxW2mQCJLdkZ/4B3+VUZOLKURg
jCAFJnSYznDWFtDK0XgPMotnFME7THgxCGNvFT+bDEXzyPmeAVPBHtV2xSiPxhTv3RazQFngnZRE
7sOcxQw2VwcylW1ygk+H80TlpKSSBnutzH9g2Cd0T8i0jezyAX5PwyZbsSoHJAQIrRrntfrPGqUp
DxWE5AWpf3kiIpYX0yIliI40kYxhVDsSjUSctT8qdr8NlB//Rnp907oS5jS7DP/5MK7RSac0nZ+h
BQiFbSLbj1L/vjRYgZU+G36axoZe9CTAg+Y6WU9UnSTFG5GXvIFYiyOEFRT7nB/16MpzjvUCCObn
h3YSZVwQB4NSxSJIJ5BxhVWn0Wq9i0+dL9GqST42ApIgZ5pLOUboWcVA0rIyrVZKf4g1dLbKeMHT
xqvY4dhu6PeRGG3QdK9yFBFUYM0UYoysGXN2sNPrZNVNanZvxmjBX2ukthSMRQVIjY4L3Tn0HbXh
I0ipNl5vgoyNGEjes8cuDKjqj7Jtyx44YnoJ5BZhrc/MhmHbQUB+igGYYbkYvGvYGCTB+7jFFDhp
mVtaB5bdnHP2isztJ+yQwXrjM7OvwogiIcGFK9CtrfimZtBGWPBfPlvjHXf+mvfr+NJeswEUX2ju
xUSmvxJ1d9cmJwY3AaMx2Bup5jxIGy7QyXHCxSiZqvsMvSykQ6Lvz1lK4bJxyMw95TPNj/ShjxsU
2O8M0WxxkUnUqOhf23OxAzKOHPRPSYo8yum1kABSbQaZH6bqN9vVSnEuGD5jZs2FNxPFF1JkQOss
aOHQ2bEhVHiFw3TmmDvqjzqqI0DWhdV/T3XCg0G5ZLgteDszYNliqPEyLqPtGTPv7WgrFyKsw3cm
Y7El+2abAy2hqQ+pGFfRUQtLRujGSBKRFHoOMQQvvzgQobaQZQpdMjZfdF0obbYxb0asJ9bWa3Aq
Cp13UZXsG6h98MNIxKym598uuOh3sWzQETeoxufsYnkoma4qA2LlIqYFtmlJ5AQI4LfGS7oTKwYz
murRtA3JmjFSVfAm631SLyowFI57XfxMKZqHmW7M4qFWgPalCmRZV3JTmRJgzQ0h5Vkm3N10j7bB
fPxa0AjQ5480zAutRIOhO0wInr4Gw5M7qN92P3+ZD5lxHtJRKsr1IKbpRNYnu6VlAMBmpTWRVwbf
RjeYXuzdr53il00VCjxCR1Io7+Z+kdFDgw/Yp0aTng1t4s442v8CGRcY6BPwzq7z7polCWi1flfM
os9car3eE6bfELIPirsECirWFFQXApXsj+eGZ+GDhePOlntbsAgHPkIoSW8lgm4RdxY0N8QRMV9k
gGHSNxeVvDYb4wycD+5KbfHH7QDwQH/DugEse1UU5g5GJb82SvjZA0TuubqUeFZ/9aLy2iykefZC
FSrnY2CBkztrZwEVphWIsq8PBq9e3MbOLXzx5FboQKkGk1NcPwHXUv2DMhLvm5ofsQ2iMcVTORTz
EvNzj4F8nVGwke6wEI+1j+kBQUMQjF962ADXte3vJlG8TrZKPtzDngHj72nDzB4pf4nip0ct6i+z
7eaD81fn5FT6LAk8GECHbUvLPqhjm27f0yGeJNWkXR70G1QqqTqK5XyAlURSfW61RN/62VL+inyJ
k17E32kjiQlS1ebRrgrgkk84I6W60bDDuSNGuxPCpBWmxGaMGq1cRki9JmZ1V8WKHJkfBNBeNiea
ArAoBM5nh1IqeoomgIpy2Erlp5ZMclYiOjRZ2Iji1VetJ4mUx0X9Mj/Cqln2WYT6lFWpn/k8fdgs
CKpBNST9A537zsizbSI0uO99OOhdQIedU23NHh81NrtBImUPUmwb3uu16Uso15r9Sw8FVZ02s2Bf
VmnFqqhXp4Nnt/HILj6qGM8opraOrvkQwmDFPtfZOXC9ElgNYGZBUDbTNqOPNMI7I7v8qE9Fu8PE
QHMIdrh0ZH/2B/cLdNs/uLQMSCoJD/icctN/gKFyHywNzcOAJUATvFWQ+WSNy6SDE2xGxpXRc2dS
K951t/GLSRjSxLzeHk67UFhIwlIlqdddT6fJ/V+G7GMuAWND7gZG3CI8F+CFpb8fLkugnLnO17XR
84XSf8PlCVA0/i1jTiqTvQUUcCzb07CoaVAlFTMx/46EKUeiETitVbsamM/EH6/cbbi2u371EW5z
MeW5ltPWhm7hHJG/jWG4uji+AVl2IyL1MuoDijc7JmfbjgqUytUsHsq4qwTTVwKdsCpIE/0H9IJb
iAH9gKD62Ux1Nvs78RCVvMJ6Vhm0SW22RTuB20BgHOPCIYRNe/51G3ZpLAsn/vvrlMsMNNgqYLCD
UIcevxIKCpumuTewvMDv4PRyr7TcYSFzKE96v2WaHtKE9vquPB6CyLbFjFKkmzOw0Eji41/B7/hw
+97WXiX/HWoePRwJYTEnW2FDQJ+0xkq+YW/R4J3Hb/Oz977pWADc8qa2ELmufEHMaPEzUQd/Xy1x
A+jowFaLwA0ttV9s49RAKSQudD/V7zMx+xTfj52OcEQG93KiMm6jgM0fI/zzc2HnPcA9BxhwnsBM
i+Eb/NRJnYE2SIk9MZmxRLvzpgCVFqCVZ/MCWCw2H8s8IxLqR7cGYyvxC/0RqG16XmiYAL4v3Fwu
m7sfE+zegSj7zltxyY0oYUWgf1Wznelm0vnTj3a5wDdRVtjWsJQOBq2N3SoH15OjbO7lJHYv9iVN
eOnBnFLj1W92rvTiXF6+SRnGW5nn85aReVa1OFl73/NP9pdfiAjmx0sUCQQAGIp9648jbO/tMApp
cdPYazxh1P9zfHJ153PxJs7uZFQNeag0Oe+VmbQr5oAnLS4qHkesCUDWimgEJRrxrA5Y0nnTka1z
TKCLbRiRUlsd71S0TjTlnLf84w2yK+I5fxyO1ggomTjP/JtUatqvyJnsVRRCSyyae2Eqn/av9dM4
R60SHbtNPT2HiuFy/lDrAyCuhM/4GhwYEvb4KKocXFjvRp6MJo2anpdv84MOvf3jrIeKba/WAPO3
PQuvvU58dHoys/55wkqmfXLT8EzdsQZiDgYbqphzgSSEBqLCqsvqobkXc4/Q/IjSzKd3xoFpsIhv
uinpzMIinBu5e5Dyz97gGyKB8yuDeBMpU7dfX5tT+DFQvz+creJQB39bC9E6RMS5rMMr33fBwvEZ
scO8NfLDN0yA1XAjcJirYUTMOTbyftPDBVT8p3MGfDBetyFSPyOZgUnIHJfHyk+v1yL+plK2Sb2F
0wC+UuoxMEhOSzHBiFADnC10zx1VUty7VeOdCwUCX1DrIX13IWrSnoi95g67ehUn5W7id4x+gRQp
ZPoMMqvQnqq2wFYYJqas1FHBsl3qpJpFYDnzKD+kPHeec8lluFN5swhhafvsBpmuwab98wCzRhAa
0pLQv6LTcvhebLvL3pu0MdcMHyvjLlz+ixV721GcZKfTU7k5otckt/RIrrRxZ5D2r+UuZep3jZHa
g8PBH8Xur5wJd/mDDUBEdw4IsfEI1oxSrsMJ+X8DFji/Jw1B65b+WBMvZ++lzdN47RXZ10uT2e9o
9oxjM+KQIklyYPNfKsu8e8IUuNJUqLLNSPrSM1VzFaLDxZJlnWplbtyOCAaIqwZdVvF8xP99pYUt
PQJzPdjMv2WyiC2RoLDikjJm6yU5CdZ4/yLeI+nnCTogOoEKGtk+tIiuz1Lzv6JbzBcuGgSaPkc3
ITn7acEDybwDO4uGy+ONigTbVxAWVwz38aJJMYOV3lITCTGYwxJcRlql2htQ/qdy7Kot/7oe7x+x
9M+crPPiPbhIzIpTWioe8U1B1LoO5Am3y/pyELbw5YWDZRdYi77/mhq9Su9+xAvoUMsQBZJ/vQ3g
VtN7+qmO05r7gONQsoGvFPQTjCN6fZKyngrBoQkg2I7+/83y66KG47+QTyiBeg5tOiphaU2MpzUQ
dAaZQu28E9TTJnMXHE6dNx0WIBcD3+hYi/p6TSudEFIz0pTsn6KAyaFQT9SldYQqmCHsPCjBUCXw
Q5BZMW50PzJJlm2WPvXztr0g+qFWZl2JqQYsWrYG8XjDCp9LuMZ2sCIDrxkz40Gns6W2/TAZulTP
abOVDpU1cTjzV3VeeyzfFk5hhnHfaDA8eUmZuP8Sule0i0nIhc5G4dJHM9dKsMI1Lq9kbbBv/IWO
1q8Pf1pkWkvQoH6i6zIZiRgAIUNeAL117lYHM/0Dr3LIzTvKCVih8UJnuX1sn3OIAkJuMewQuOXE
SvHtK07BbtIQ+eQGWuT4D+VPEEvediLcfuyHZE54B/48LUcFZnv9jYzi/5RnsgROR1+ZqVeGvUsp
hh6p0VuwSpxlRV6FG1lYUV4q7l7yNsNl3I6mlZrIUWlLrjy8VG1wPSX5xV+M56Lfp/xrdqBO8fBd
BHVv/5OpDCGHkkpTha32X8UVucGTIJqGb/45N51KCJtC1ejPxvyRBW/1UWsnBE0QCJNHegLTzxWr
Kiz8awuST8EmVpoP7EsKuHBO40Rudnu79qkxfYg5K6oYcEb+ERRyImN+QzM+pgp8g1O1NUY+dbg7
3jcswMUF3GdwIBI4JlXmC3GWYUV2y+y0Eh5XidPZ85WO+UcTjlQ1C82+4thxy06A6WNPAfWNTzIJ
KQvRiEXLc48/hTxbnjUpeIhum2IPJkKGLDImkycIm8N4IVYf4nYxi+dpo0/EbG5t/HdSer6oUHLZ
UxyD38+wSOqZeZ9nLLCjJ2Lg3zQpbWcY0MOLwqdRhibKy/1rhHSTIxWNTzdAmCfq8ebZbDIJZiHp
/pmNu4A6m8Bw+B/c6MzafBzOo0S4ub7bcWghDs7HFTZp2DNgu5Dwj4w9dy1SOBgn4SuH/d1f91+2
jW9xyv+RCBRUmkvunQbaSxrX7cvo3deoRuKdehehUEHbA7b5l0/aI0id+V5ZFU50VGlODNEXPUpV
kW13R2dRUFm8J/VFdI1Od9QOy+dOCzBh/EYMUCETAxvulOqf5ODZTGOB6AZZBtbZ6fEvdgeLgB5q
BRhakL/0UKpQumeS19/69pmhs4KQgVSHELkHdjbirqMtCDKS1yU+qZ+1lxj3knt40tloQCldN9Ir
0WD+PGrxkQqEtUJU48paQyYxwzrQpbzQKgUB0GMKIcfUIxV246sMWSWi5jNe0ncusZ9MwBp2S25p
m2q0Ml2itdpI8TmlLBkqIMcL2YK5wQzijB9g0sHYU4l3LxqvSm7yuKxfO1dNc7LekmTQcQ7c1naA
5pqukFKtQn/UJmgg2Bd0tEeGY3pW6OzSjUX6n1JrnOvTAfqchdpNbeFvfdM53xaQEKJg4S+flFvM
NMdy0bzOFCILykWHOtgnuLVWRLJldeTVgMIO76fLzdNQyDPwmGyI/4ZHYomEC63HOg/B9DcL7s2V
sf0/GiLASWdlIqcMPnVccyyVx7aYcjrpf4sJNEnk6il/CbfuSj2Ja8CEZObBkIkg7+xzUFB2XdVH
mii6S9Ke0/vJW2mHvZ2foGEvcXQc2lrYNrHE8KtJM1pwX15D8xcNfjhU07tZ9XWkoVG1ODyJEukr
KJOP/QvgLAMHlRRR1j3MvPhcSj4acRrkN5cEj8fI8t9rdrrlU4um/TASuUrk6kC2VqdMo6/T1bNz
ObauQGhdISSe+pVKwNgZ8nbM1WgpQFOkHTXtA2bFEq3UCtlYE1qL453w7teCBnYMlyMdScXYFC3t
EOfkOcIxMdnjLqj45o0KhFTPpzQNRF9PslMSYdd8J4ksG6GykUoOJ4thyJW2AaVNylLB1ekQHrtM
CrXaqh/PO0N2EsqFKgQNpsD3XD/MhWMezK53VLaxpdwKnwRiX7cdqejVmeCR2ZJUZEXrEupDyZTd
TMNKR7iqwpkKwJWwqLk5UQwo9xiVJv8HJIhou9uDI+qzrdoxkuD44uJ4ATXxpmowIedQxgA208Iv
NyU6CjsgQgeIWpB1axNQDlh5z5T4KGiALBxSs57HgJ7dChyVsniJZFXIxjuw6g3sIIMeDJz4PzsD
99k1Ox9eemJQSMQs8PQV442PIUzeAUEssLqadeFkzQE5rEUAImOy9G5cszjqsF4eTFJpOcsuf7Di
62GmfyijJNH5KmVKR/e9zyZaXuoPdnapm68BMtF8ShnYXaY0jSTvpB5b3OowVkpK5eHCWxbcVkfW
gBqqsGJNnCbfYi+YdBk7gHAfR7fChzW8kG4/iywee/NxF4+qPDgCfrlJt78fn6ZDIm9c0PEc0jxX
NT/TLEJcL43D1unwxlsiO1m/YHn9QWqtS3hMrrlNHtlkOeWyu9LeraE/Hjkn+SHFQvNq1NJjTblA
lk3UqsysKsLDXVcHCL2zqd0EvvME1/J3I7FH+RErh9g0NJ5cetQ2ZbFhXb31/PHs/uKeFEi2a61O
MAMKC5niVvFtgeWuKgIq9GGI54rimXpUUfwph8U+qLqfg7fT/TAc4q2qtlkXr5bIbylURdQm8Sjv
iSP9mB3bDl0yNhHC8oeKQ6oDtsr5hL+TddduopKoWwSK/JI9sTZDl/ukcnMLCiBTzj1QmVgElm0t
M0zPkVXIt3ulb5pM+8xif5Jwuk49RsCTMyb/DyfTzz2hymd7uTc/bKNdyxtuLqy18qzLsj3RrDBu
eaZD1Cvrp6EMkaMM9PclWvMYmyWpxYCEinzfZ8hC1PV8eOCjeruT+HNtI71f1YnlATpzulw0rw46
4rOELFBnteUd25bHM1JyibCMpRdTfnhou6ZRoDL7BJqAPj/BP83qOLBMiohqF10l2sFvG+VyhNdL
nX99zbHdTm+W/EJxs54ovFMbeoCVD1dNvG9Z9sQdxhJqVCPviy9Hy2Sh29J8SOhp2+d89ZgIdilm
fxF6DGSH4X94bbNgKcRMZyvjrpQMATXHWd3W3VT7Y9FVsiOVBRIp08X633FWgYrRdRRYkwe3wnF4
xTWSdbnxhOGqZQhi0VnA/Bws0TCh3BfZ6D48eMdPddfsgL7mFx3PB79vOCn9+hK/r8cyFNO9mDpA
+oY3vf0Mz5pQ7STmLfmpJ+GAUheHJZ2Col8mop6ddZuqb4pGOjDZF/Jtyl/8U1Iqf4rT+jbDtynC
AsZAEckk3BnQ3eeoZentH2bUrSGMywR/o6wFnaagv+1f2VoR5mzOJeCFS+42HWplwUZj0LKoNSZW
ofpROEIcEobjVdbyWY0m2igVpr+C1JjnF9gAuhh/Ot0GH6yKmR+rTBAm2ptq9lP9TFUW/XQBgeUP
4MsMsOh/siEpSVCF/EfHUkgNlonFOwS+JBhYWu80cBTH2gAjMyQdf92TQB1BBl+nkfeSxX7rxFaV
IKKsvv+77wGPsMgJ2lq90x+CjGT8SsREIXDDJ+GJe70RJxTBFVDebddB0h2bXZjiEOfhKqq2s/tA
jbplPXW1CbJ1dJyFWDOGJhCAx/1Sb4jm6tcH1Iuwb6aihfohbxj7savv0RF0UoUwoP/cuoF449au
DMPfLmxV8RV71p2nXrftLhtSPnCmlsK+C/2OXDbKhMNit3YJHT6+kCnHdSFnlbhRwDobMeaYY71a
wGMirhRK1dTP7y9Qe1X0MXG9ylO5ZP4tjN3tewphWFW/W1TQKALuZ16s1slnEM7YizGQ3WwL23PC
WKotb57845l7Ilr09uyresoZxzMjU6vPqbdv0LkHz4hDaMML090jYKvSMepJ5aUZwMedQ+DRw6Oq
tf++NPdQoAwESI1fT3/ryoXVJpUuKxLMC+/gW8GGW1UotzvxyUQqGxsAaRXNtTa8OR4qD4ZT6TQY
tmkxo+aZggfmuMhzyMNA/ic0NFVeWgQwsbBn7KyAC9EuQ8XJieZPh5LW/f1n61qw+oucRp4pOU6q
1hnby3YelsadbAbAvoxuBHk+osPxNBUoOm6WPzuudYbXy7u5bLziYdoZ76FDvedxaZfkIrtlMsJ6
QYw7x6NA389LBzi0TyEkQJEq1cFgTsRljPHIYmHGKc3t0nLNcTRqqoOMgp7Xw+TLSNQtLTeHEFyC
Zngtam8lA1TfXxsUHUmpdsy+CAAwobwrcqje1GphZMel1W9hxyqB6vkDwTwJXBDKPHE44w+PzayO
gRB2t+CBMQJ5hmHJ8YF9KvweqaF3rryxt1LdVBTRxWigD9uK+oI+BIPt+THxOWB2JQQGk1+x9MA5
kuhsY21RModzamjHaQk/W0Qm86kmp/XYS4TQXBTBSwpDKsq3r14Ckd2+sjGmXaSV0ZwxFX5hlAfk
TSfvAfTmH21cK+lAzpkgKfkgrsFWhkrFbgYrWJ2QFdRVdorItO07SRZCp8vc/lrsM5zmCkwzFoBC
jy5Wn4OyiDDK5c1lXCY+VEecypV0bRN3te25zD3A3ZO0QxMg+vcw4HucZVN+LnxRT+ozza6/vGYM
vsXlCuFv69KUPZsy6yyRJeZfybKvJCqzS/ypaugpWyQODiVluSiLw898wm0GWC9E81O7bk6LIoo/
9sjq3l+C5sK8uN7awfh/TXURNJwXX6maaAgYPaKkmlSOMrAUGzRjfVnS5xxWG2SNEZjVIVawu9X8
nfGAa3jw0JWiZRiaq3taMf5eyMZjKdjANAf4xFjuvs9dOR1nVKQs/Ygq7zDZtWjSQnDEwS5xPkPq
68MDNX9b8uGTTDkc9eWbg1KkgW6hWyw1UoohxuBfXr9mKEDtOrZztpovHBPAmieXczSnHw74bwuP
Q9+TzRYBkgRzDO11CM23M5XoZSiKAQ8e9oiz+2yCaoFUtNU1X0OyojRjVhWc8WJQDY0NF+0lCjo0
trQH6GJtS5Jp2A7RhbQSKonCFXBFM3mOyNPHLCVo7k3Hxw2O7ayMfqRAa80aDyD2bp+2sDcO0bhh
H5wfxTgiZY/KD6KNjmtF6GLBB5wyLzDOLw+qp1WUtDx5Vv8YXfgvq61OHb7rgsHiCP083E8SQFTj
bADt6X2bk+A76ruAvjjI08zcFS51U72KWV2DoXsQc1wPcFEfRmxVMlRTyJlNRgYlFjYOY2DIfDT7
UanqjoEbMqIDzFBmV3MLcimMedUUrjFM1xXbAHyYktdQb2FS7rA43hAthsqOnjTDBFQnFzlrJJgU
+PB7ZjONgeCmgPc5CgVCVwntSvGbXlQxkU2Mr2lgLY59SLONCv2BTVKn56ImOV8IOP0AGp7GdfZ+
/PtsttXhB5pPwenG3oOmi3nvS8KGYksk5G1pV0LSxp/fGLNTh9RBRjwH1TiYvM6SKeO31PEsqZRN
kXX4n0Qc3CikMPnTYVIWtJCWgjdQNmQICXmW0/cVxuadzHOvSM0uBDHUIIjOfl3KxCaWits75hEB
ZL/RQc/dH2iSCoVSscMHkVz5EP76a+dGGah1yc4pgUV8JIp7KZJhfQZyImS94loZhtIHQKjIKJUD
cvI/txTaVGaL4IjFSNZs9aY4KuLOCnO5+VaRU57LRG9R88WYy3iWLjoHTgDwSBA6+2P4OghoB27j
+4rTOr2QEZjn50utlN/TKqkRD3vDKLIWieYj4aqLY5B1StOmk8Uw/6WPvRcsZE2ZHLUxenTCLxDE
XQU+JwzvhlUOZwQFcIka6U/SSHIw3eg6zXK9XA5BSwt+k/VIfm1GZXSRr8MbW6CtlpqgfYzVC3/m
cLxt+5kvYUeoERSiGlvOJytFxJIejM/7SdaSsTo/GMqJlCp27eKUI/x9xvMlFqLAHgH6iAbLGbiR
lylZzKc8Ndth7lprlyuMwqskQvHjh4wCwsGZs6cm+0k2uyqV2gdHDpbRjZdlfQCTfznX3HCDoDT/
h5oMSR/QYYd3FOqX3bEZNKZ3pYRSvxaKxk4Nu4YI92Q4Y9anCxXpHjR1xSZ0HiQTg9SYsKt6mpq+
vOI13KpRnVdWOzGLe9VVSGPZmUvOnZfHs/43rLdrHktmWqVO/IR55lv3w93qp5HKp60276Pej4fq
dmAQ1NBo8mC66G46CNUYNQjmf+0E2D3v0G5Sfc6dXrB6QhYqsrKr+x9tKUHf2UzZdH8duz7Vf2vH
4721WotifPI7J3d4eL1g9OKwvy3a5CMC9g4Ys4j1A2yuOoJp5EyyvODg0h1yH2/dfmAUkhSBpeiJ
sHBFCI0MnoJg2OzMOd7i2DBO5V2RUkLz1AevjpPqnGZWdBIbqXas9+XUKGnxpACdYCcn2uX80yuT
rgHP9rxpQG6WlHZ9DRI4FgmtzIkPkpghiJXRwhB5yzqGjG9bkZ/6KmN44/jQm4rCP4IzYdxXRjK7
bt3v3H6TpP4q96ej3f7HiuJfCrxU22g/Hy2Uo8z0kCfzGCZ7CkfIxu1zvpiCaBUdFAw2PoqO43QF
ND/S6AXroiSiB7xxoWt80hJveB1CKHmeaJStI1iSiOFu5Nl6LDdtlkaoyF59tytaECYY5UArbbVh
kSIBPLaVbHLqTIWDJUi67DozNyjFesdzX9ROvJpfj+Ww/T1xpPOP/ySuL5Cq9MCZyh0V9hXovwk6
DRU3XocRklNHk7C0IRoqLXbnoQlqpVqaxcG6kdCOrcuQdm3k4wd1pMVyIL5ni0LOOqBxx8C8Yi4s
2DrQrIcNK7KRjxpkaSpAiq5wTAr0gspWPvZJb+bLA/4qv15x537HExb+LnPM8LEzSvEijstNA521
6O7KL5lsQ08BPMMnq/ioKUvQDkr6b+RAcbtPk/bA992Xr8n6r0TCT1jp+/3nTpCpxzdrrFPq62mt
rO4Ro8AKhlXIFaUE/2pvskHJlJ5p/0bsgfeV6vaDlexa9f57XQngw3tuGg87iBHLb6vzON0Tmgh4
0OxklYXa5y8AAd1aQe+JKPU3DlcPesgFUloE0CcOY1R8V9u9dPH+KtdCXz5exkbnJg6pXolbG+oW
LK7V31Wp4B1hbv+MAvRDtN9Jy4OZO9q5M53X2db+v0XwszrirljQCqStFDgCNFKMjvz/hjfaSdE9
T6sgz3iHlppcrtM3gJlRjtcHGbA5RV34dAQXXRkv4hrGX3eJkAuF734jK7c4nGFnQD2i8i1Nr8Mx
zK1YnFyIVx72XX3hDICQr9RjdMApQNaJ+8TkS84i1nY1/zyV2R1T8Spi3Z8wcD3YdQ0r6NO8jigo
Ap8qQYtl3CpeNosMpKFU4lvEV/N4FVlLfNbbRtM+9+wEPzCShN8pqnzLSPmlbWTyKOFdNZ6HWbZE
av5XDoD+WqxSZBIXEkPjOTK6VZGKI31tZbYJrjoHfIUmnSJ/qlKhxtcvO4dHkwj/yuGKjdw/2wF1
T1EBB4tvnihd52WJ0U2YP6BZHMm85dnI+IJ9eyurKyQ8AjjNzDxUQNfo04m3Oz9CkN8Z3717zPlN
F7qjfoX7CAOrEd+qAG6tA4kyXKkFSmoYzPcqW9x0nJgsnv92YMIPk8AQ36SL5j4VSJnmEiEZ4aUh
k4NHOCNKHRGax4hafABfChW0aVdDqqlB9FJKLGDQx31lr9xmeDNamJCL6cf8Wk1+1QJcH6dwkAPL
I8db92djDeXlOl6uUG+kr5e58DWsgCEMLocyPiwJOtOsXqMrb7FweGaPl5Z7ssrI5CBZmcy2lOOG
TTAuHf8gKIEj/xnwiF0AqefP3ZKnEDsyBwMbblLe80/hPwE/BHNpe86ysCAu0AOn39Ea5sLvn98N
6CVuzdomFAD6LYxatYlSWFr5CJgPtGs7cUDPskdf3lJ12vBW1XtRe+1bm/mHl0YXXRhbQqi1Szve
dijqgoRusI3G7KI6cl6MRuTVqvzHzn9BkYpHkvCI+bQ6+fSMGV3EhW2BrAvIXGQkiSNfvs2UdxCi
wgSyfGK8vHNzBPpEwM0PKotFmvA9GNOAjr98yh4Fx5oJA23fNfOWrn3c+tABYwbQkTbQW3wCHSd1
oTf10iu8gYKpiliPhQ4wNrpbM6PFndnfl4bt3um7gccQ/j067TosVRqZtpF7dgPdAe7VJEU3PnVm
JENQdOg+Sg0ds97wedOE9Vup35OQpw/S9DPsAuYB3zLp1J/Hr1EhCvFbWp9zBBAGTcu0a0RtxfW+
LojdJbRxDL7xKHblMtfOPWAd8n4xrPTbCdqj2SzWvx8Ze8Pkpw+L9DVTNLHbOW5ZIONQ3MTFTl3P
nUEfYs4k0zvWIgnyxgHpdYIXW1fjjP7B43BJlPMHf8swTImHg4iqXd/IyOehtVm+qXlvJuC/RwSG
JRsBUtyFq1p4asAXtTksmrclgfAsb6lKiFWYMxW8DxNtvZlE1A3XV/X9c4cxKa6ab1ZIqROccK0o
DgR3xoqgcomcrM1+iv88Jsq1T/1nqmZLuer05C+yox0EA9jZFykuONQUo+8s1IwxqV8+PMCqY/zn
AkdlSD9pzqLuaJLkfj83NX5hTvyyfzo/4ZPmEkfMlS6ekD2mip9VMkiMZG1ThxRmyK4AVb1howox
AfAf9SUq7YBqjIUL7vptNAV6NMF5UNM7gm36d/tyohwtAMtBqniNqQYavz14IwdUBMmbGrl/N/cR
DxIFYmbcZ7FUt596VwqgAxxBO/Sskm1n61JHB616+cLjLGMKQaYryyVuf8cPYYy8jsNYKCFOXKHI
ZxGTZH+NiTw0rrJnqMi4gW47kCnJS1NjxwTYiEDQeJcKaZhgHXQ/DWgALjKzLST8MnGHcre9t+rG
XVeuoVJ5HwWxAZRqqzvf2u6yDt+lAqZT8LvrPuPwfA3Z+FhwclToOM4AE4v8LbmF3LTrXMldc7cL
mqwFtjCUmexb2pTOA+rWQMZP+tJWNB/y+SZmtbsZVQLzNFxpqhRXmAkN+r1PBNTaYMlG8CI9BSzJ
iXrkyHp1XXW37tdfoADIJEpaRaV3aUSgdiWA70dMiXhvw3OdF1ihPWUD3ZsfhOBzqazTuBdk12ip
tumSx2nbOCI9Q09iCKOylqjqQyUk1lx50n2rF49WCAp1w0cNyuC2CMpCSIalB++Rl4VCNrIO/uy4
yqB8YRhSj+shPZJz7luhI4CIhMGPUPOu3/NKkxttp/0sq4j7z12TN7BuAGuobv1a2VrowrN46fTs
GKDZeH8/sIINCHBFcW9IC190LyMz57NjnphcgXckBiqOHv4ZhjzRlNdM1v6+2U4j/W58MICjEQrX
IvcKUdsH3YJKVmqx0jw2eHr3w/ihEPgOqS8LywNiVlvhQUOhpYYIhCJB2mgkiLqhEF6lS7wtK4bw
N7SFGsUDuUuVWRPGhbJ41OB3q8Jqp+DvK2bWUMRU1FcJ+z7UqgYkhXxY+u9LU28HazXHz+XiNDuj
S1XqbKS8ZCL0K65c8T1el0yzzJt/+3Sx6sksG45x/RP2qj8h1T3tDYptRHQlgXlVrNtvNAqAwz2g
7YjXz6N7AVxq/BPiI98fqd1xongoG757YBJ/co6tZrBdFPOfjpOdtwFpD4rps7/4WmtJZ1fxlEDH
aZWqtrEmCvBUBYK9J42EaWyD1KcIRi3vT29vFgofllpRmsRmgyhyXHRWgk+2C2/Gtdhglzo6vDlB
SUZG/d6W54heEk05Fqqm4qbFgR2faCEhHZ+wdRUwjltk91Rs6q5cZhFPAWkTRuIiQBcS6zxKKJzn
krdi1tKHOdNutOL/ASS7rmKZsGzlR5Pl676nm9weHlqzRN+Tp5//9M1pdEvM2Gzsh51L+JMN8xYR
PZ9QNdfaWX4rD9XM5lXkHdKQGhux0bTceYhe4NExJB3w1A/Ur/5dr8CdEIw3+uAVC4nVNlEtGK5B
4bPYYQCSYwaU6f9QUzJSaDomg/wArbv2+IPtRJkl+XVc/n2cCDnc2FI3AGMBwTwbdn1Ndf+59U4r
MxRCygrj9zfSBXIBlrFXhrdl6utzD9DrTDTFRrEfJXW9OcXyvHBvU/FHDIVO3/pe+ySAQt5Ha4bi
9LYWR9aM0BYplCpPZd24Ftq9hV8by/7Mv2lKyHIvO2ynr2ccUQLMCXuMVIwxLexoYghfmLXvQN50
Pw4gBILdidUcaH8RvsY4Nk5Xe0NznywMy3mKlJNUnGZUKmf3cCGw1kANUH6KBWtrcmXEAuRawTNb
fHS5Na/TGCy2g+TLifjGYiWgDB5JXa3zChcq/cBpTMh+Jr2EMt+4Ni8QYYVr/a3dJFa/AsVFIK+C
cKoafSL1Eomwe1iJaiWP4nHPcaNZzq0Qzhopdi41wrMkD/VdQrhFoPua5KyNvnS8MfgfSsevT/ZS
A46Sgp3W7D0JBKVlc1fBFMPOSPlpD+vRumfWgzI+EPVu7DH865jC46HIbV9ZvTjW3M1lBV2x2ezL
uCykv86Oe+qdvkUT7q+boYHLuisCBXWmV7avhFF45An0JOWKuOf2cGnwMCsAmD9G3PE3r4lxK1fC
tiq7TXdq31qATZnac93Db50XWgpo7f4c39pPAgOMF7eOilMrga51ALzaRczTPMmuzw+AGMR7pzE6
fSZYA5k3jJLkK+StXg1QG5Fx7TKjbzQV27qC2PAOEgE0fI5mY2ASJCnfnx6LDpjOmK/ssNnnfcFP
g6IuqPxMBPNl5Go0QE9N9ZqI1dYRXneyYZLQOhZPpE2j33TKX3X+Q8yLft61QFgCmKkfHIEVb2xF
gcsyaRNaf5gRYl6odvbSDRPuxBCBKOIKPWqULIc6ZbsY8jN9KFPNsq2gAbuBy37B0j/y/7JoBkVm
BMhIZDeqisH1+fixUiWxeV/6j4pWbWADkargTFY20zKHcstOsg3PKYYuqMaTq5ACyoBrK6vIwLu0
J844VJa5W2Iys0DpilLXMG2P3i7yFB/HVpOQ6t1NQBduTWU/YIKeF7ngyG/GNVT+1GsTEwdJdDab
FXWN5HunpeUMdx63103vEaVuZ23Ax+SlgS2v8NrXwsU4JQ8NesPM5Zjcs8tEpyXoKP/1poxoWrUm
KIg5ShUFUMTkgPYnwonqtlHv8RYJgXmtT35gAoc/1XBwulKl6kaKcX+qttsV3txk2WGmAJYUonp+
TkOvmA85aAX/azrv39Nm91Au/7KzC7fsbNOdkfVcR6ReZx3xovSS708d815QjtbRbF+GdQEq3JVZ
pKHK5hJwFiuOZ1AkSKvTsRpVQAjqT1ScH4FswWfKZXCmebIxOJHnNRuU3PW3LafDN+AAuNBTxKxR
J7rvXSmZJjqpbXvHVpUoRPpugMVszhxecHjnWSc/nn87xpImfX8+dKFgHI3G2kH6BiaD+5oeEjIr
COfc8XCzPg3oWu6V4zSj1YTLkkCYJawOujhO3v8rg1UnyvMO3IbmWazPT+hsTkwn3e9YaXN36dTP
28RtbCM5lVXiw3oVNYeoOlBay2M8GFPyNt01buZshO57sAY1v+7TJqOnjgd1aldC4C9pNW+5UzT7
8RDn5UqZ0tmL7eQDjvuB3VnNnkwVlvj2VXQW1jaXyRN7W+rI8RR633WG97b+upn1IDczcXcqp4TY
jSkaobYpPHRj5tGZojW2ByeuDZjKW7B7qV5jn8hGzakEWIC9SGOC6mCwCqcj+8O0wbIa6hCGAUGA
LIA2jAbFapIOOm1fLbX18jMwZaEK4RDrwEnBng5MNKmk96e60KJ3VLDKRA6T40opM108UCyTM5GY
PvmZuDm1F//DmLosvi8Rk0ZEsuxcln7RMfWDiQmHJijPkoC+swrQU/+QcVMzPxrRR1SGyUyD1Xp0
MZAfVDW/HSmk+TPM6uZA7P4LQ/AwRlmwfhfkZKnDv3ugmhMHubvmHHM8ZviPRQwgT2gjq3lW/3px
H/LPW5YlQ6fDhGt90OsW/9OYspSupq7QEnGVkpUdedLC8tPXWYH/ym46dX/wJKuxElGEYdoE4ZOx
ehxlvMk5ubkzSxYthRT3B9/K+bW/k2PSgyqmegXFAPNCfY/ohVM77p+ud1bbguTYmoqDcWsK2EqR
kKbKRIRi6v99fmhEwRtiBx91vVYsaPWcb+xuzO9IZjW01yc/dEpB3O7bEk64FkyrDkvlyPYzqXDC
/7IQU7jMLa1R7U0QWzgoKAinydy4o/e9OZOBTmDEUHZmKIHRleRNey/FyO7zMlGxfEE0WK/tTlCc
1e2LdERrNMI2E7SaE2uWN0WrbnUhvhyHIvwOZ/G4xG8yPZVBOgDLESyokeKcc/RKEy98R8kfGRO9
/8MHs//885EIbVlF4eRF/2DKnqFcBcggJaYTM9FQ5vEWhHo5nFUhJ7y0DLLIc2RGkH/QeFMrB451
EGyBmKF8GD52oFHEKoaflvJ0gsmQZnQVez2cKbX2bopylje+ymt+OMyNq05fnNJ7a7TfUvcNyDS6
Kxpag/uWNYbyMorrEG5jNr46v8ULRnpgp3Co7MfwcgBXPAkimH6/c6E4ZOkWBqVZiX/dh92bFXIx
vSVleULoMJBO7xudL6TMQRPaSOWsvZPR6Wy6hxpjgSYX4xnjGGYOaV40wB/WqsOtVzSkuSw+GUto
086vReZ+S3h9cwbBPuXmpb5Z1yPY7Qu/k9WOoPlni3ZMPCXyBOv8G4FRUJSOfkXsfIxJUHY/mkvl
O5kJNmLd7fpBmXbhdvjo20DXdf+CZ0xnKmYAHfawi1tdKD/VXIFnVW2SwH8f+Y5CyfQat6l+Q86G
HDUKjZi10Ah71KzzBcKO832AvY2OoQqm9xOrlFc2CV/TsHEBJZaFRD8Clzv24Meh7ighPixa6ZAA
L0j6gNmo07X/eMZ+ilx2RscJ1qPCp7uImbnelajfDZrgmh2ut2DnnaGn0MWVJ8u93Y4w/Ay8kXJC
NIfEzH+Mfzc8DaGEmdMW55sxu3GMbUIGRbD+IfKyJcpMd6x4kQ3oMb5+p/37S+ZhxF/rVRbU05R7
TSs32hu+vv9FYe0cwKITmf2jaBox8KAqGXHIKSvHQFnhQgqXzQTqEf00cyQEViHp31Nu9T+++EOo
MdpmlBGPd9lzjsFoY95setJ6d+3bkBpfuDf0pd7LMSuqwYpAgfgg/Hkgz5yE34P0NbrBxtlrp3iY
kquJnwqyGB1B0H+M1+TNNVB3DEpjA48vOtw7E79vdIS0DpDfaIAk9Mw0vwC02UN6XLByf0ZUp28k
hi017h1fCuT9zIAYqbtfQ2G+Gdy1xHCGSTFPRgRjxUBr25bZDkrdmWRCsD+diNtpkxREHiki1/7I
loge5tsJnsbYQjBzjAM2r10KYZjpmohVpffj1kT95xnzmxwko5SwjZ0NF4jINj6Ii1y7EYvAdDF4
KqQUtNt76c31t+0y1MbiKM8ok6q7mjdawiSvM2I3BpxAtYVyIq4/O4wkNOfcC+LqkOOrEtWqPJBn
E2lowgZbsUISBWTlUbwEp+sqXtvpWramvqc9fhZF0/7o22mm+2oKamPg2zv5W2MwzbQS8YL7pB+T
u1E+yBStaEaae57kXRHvWJ1yP31lNOcLBOOLLFJmI0IlxC4Ut3E7vI5ylh/J6B4baTUBBPVCIKW6
SNbu7G8gfaD/9rnNZmB8YiZSwQ+fmW/o1dwO1XZi7MOvdpXYgeauOVnAYZN87bh8q5XZ8dbMZl4o
mhWzH0ISdOZrHr+Ee82QB/aOEIcAsl3vesPJVTvZnlWqbOFNhwMZWkGMRahgIcys73LWKLb+gSTe
XXJ25H/l5gWeGnO6ZwAVIfTBAc0BCkjSZO7y0x1IH4qBAmyaarJ9mgNUUkthN7Wjq4FA9liwJ3Tf
A0L06b/c2eLmUJnTvPsq5nyaE3Dv+qR5ZWchmMrAufWraudcIMW6hyDUzVcCh77oq6yrl0Tyy/ye
1il/20sdQEhKmLMGyxbGn/ciPyWaxwjn/R2eS8LpHuXpmdomw3Nn3mkUuFo3k/Fj7epGbns1GA2C
N9ldzdHfc0O70lFJ80g0ku+FwYiKBFYSDNberFqLhPJAFVBAMdjT2jxtttXOAJlgR0fWGxQDxoZT
tBKwl4skUEuwyH2Pfi+tbnUEQRQ5sZ/yy8Zsm8lU2kqAj/jRLXopGdGxK+sdE+1E7oLgcSRiVgYc
Vp7T8NLwdxAWEBO/6zyMJ3G3QE48eb/9zVFKGfcXr3FRu5e7DdCy2ZKD+Cm70TG7hVItL86q3xmy
3szcgv21Z7ec5yoCtzFjPC48/ADBleFi79TTnxOuMBUbc1aSHi8FLaNQ1cYNuYEjo2g4kRSNbyjU
aHH5PJxdr2XdflxDj9dqO1hm4i4HYpFGWEM5FekumHMFOD6o5lf3XM/zJilgGDrZe1SzGDde8ja9
ODsXLQQjI5O6BsUxUwInlRV3VTfrUhzqGsAt4/x8N+PHJNOfJpwOOyAyUU84jtX72of9Z2QQt6Sm
ZM4OlVf8dtcuNG7PPW77EvoAOYQp5Bg6Wd8qaEyqv+2Qay31RAXunR/GXUX0zVLkwY7J+6CZZA0g
5+mFWz2/K/PblvtxaA3XRG5XHnbnBVNDUesBnxW6gX+IXcLBVeqRjOU97D3b2sYSD8voLq3GA47g
VlBC0r/lZ4HvtdMDaHFHzj7OTJT8Xjjn6ypXEeVDym0Qvo/Llv5XHoS0VFoQyo17v91jRriIc/aP
3qODJmi6uLVB9dnrg3Vn3ggL6ecT5DoNj/OrU6rec13Gnf4LUxkC+y0K6SrPlBHdt+DG9jXzqXY6
+g86fNEwekBIqdV5a4GPEXsMH1Ay9rsPUvt70CXkdW79hzidxniYDzLdJwYrODtXZs0hsqrQPpSI
ENQrawrsNQCKjgiLqa7Wt0gEmNsoksmGoK+fCTRzfDvVWuepHj/QhsMusSY2CGOqA7urCHZiGJ0K
0+oaTioRUXHUJT/E1NvvKC7Umx+BxBQdbcWVcxMH28YsHFagb0jN6oJdjR9MHB9w8i+/aNiHZM78
E7S+cvsOSvQpVkRcvF659iuMzYWjISI2hrUN0Kurv8Vu6Kumly7fHObMIn0a1u9hfl34k62Xh2SL
Luz+I1CCJYMtxJ+t1JZukO4sT0GXtwz72I6upPBd0HerHZVvxitOu/kLs67IAoXl3FnfZcR2FCdO
IfW3RqJZCiNFqItX+3+u0px2/F85Un9V884s5dTDt+dVR6ilqx7KTcH2B2i0CX0ZVQn4z0lsnpi6
bgLZdVAwjcqk9LcbM+gTViqtKlDQI6eg7dZiOVsZ0yuTkd+tWPjRI9Go/Rfy98Hu6y1XiJ3Cw40C
ZvA+jo6VOlIye9I3fU0dOWeP2+ZhYbTPNKYd30SxQ9ZOg4GhOXlESbIgQsKegJLdKGLVDRv7/C7s
PnAiAj0jn5Qy5r7WEiSvr8KjHMAiu1bAKiSrhhPtrfSV3AjtumLvgzd701vYSEmamCTcRU32nxP6
nIh4fsHDrO/Jzuq/6CiKYLUB/MPHM8Aw8HSIe+gJENFVIBvehQwAecrFUzEvlBtCoDc/4XRPFKMU
Ui9ZsS+FrZZ7ReqfBWFQBdkSrIMH/eCDFEOVMk5CZ+ItRED4Syggro5nZMTfiJwKcnPyHJqgocGH
NksQsfk/RtqPlreQUR6dOiKwCl5gZYglhT+cizLgulVLPAsgMY7ogvDMgiBjnQiE7oyIL2Qemsfb
16Nk/5rsBROhS5f5KZLqBnzKx8XFV4a0ceZ7QK2S8XTktafrz6dZrIPkFGEq8nA2BEubYXi7U9wP
l4YpYbGTTQaJzb2G03DP6VOYU4w27aQegkcpFJDdnvFvigZm9XzjsOhHjxxsGL7L67PfQLX1C+6u
eI/nYMcCO6/xWgYZ+A52dJkvnpkT6sqY9Ntlcn1F1XliIfN7jl3FGjhHQCzmNUwrZ0jQrVyWW+dH
SgXOo7Lj2MA/s63qqtz66KezgJFL+fWqLTZxi6+g3sMPeDdWp8YUVmrFh6S4BUeenbcrqf5cvLQC
7Fc1mhxXe5xDv/IWOH/4SxotZGY5f4YM6Yr7TL57XmX/yluSLfp+a9wAVMT/vPeiaQGvvGflINZF
owj7PjQBVy+3Lm7NiUj6FxZVU54c5dELK+hwG8ORgopZQcUQD62f1Pe1BUXY9XOdbWltJ4AL9jdZ
Ff0kONgMkDwIKRVTj5hcAmYb48uuU10IKgqTjAe7y/wp3DnDkwANbDxd7VRe1IexNRPxk2ceJXRX
FA+ONV3x7EVeF38h4XFOK1/qAAMscKUfj/shhPW9FXkUvgFaXYJl3k0Ojhgh+vTYBP+MEJqQmEAh
WIIXsHMbbIDdlApkprlGq++xW0HalWlQKfjFWzcD9yzS1T2VuK7ls7u0c8Grqv3tF6oZIqA6tQR+
MXLHY+kRiB18IczAF47H1KJbwlg4OoWuc78tJHsMybM68Zf5GZ1RaU4AXxbLJL+Y8TFQA333/dcf
HDvXTK0SCgrgf4WWmvHcNwcuzN38aj7Ap4MTebHfAvC/6mCds1hsuAyghfLP8ZGUUSqG5tYehaCD
+MbW/O0Un28SZgq5grwHr5VhLZhoRjEIfkSAvopoFsTtrAjwLoVu0k8jmvZPHF4/OjqQ1NxwmWmp
bn90UqawXDJGaHIEIZeL0m3HyoiWRjQXPuJ19/8vy/bARwKRAgUCsMU7HZc0OrQpSb3JNGDJB8Jp
9LWRaEwpmTBmvruEzvZBJee7VX4PiSh4qUkQOEq9A3yoZTOA5r4hrYFXpqf4Wyz5ycXNemI1yI6E
Lfi7slUTReh9uAIdr2tE+eECbcZylYMW8RZi8lq7KdwluUqiWpsu7bOdgO/5rBAxJoGGpo2By516
vuQ6XApsirK0PhMq8QJhoHBazCyIv3TvZTrQ9fnCzwui1BGY0ZToN1+r3d9FxHru1ycv3p18q0zK
IoaSzhI5m5N84waarZivTaef0nzjvBDzj/9ce6HEN6fvnVUCKIix14StkA2uHA7M9xsrDvc0vkcJ
pRClU4jbdr+bTKn168sPjUPNED4xKCKBgFKZa6coWOKGWzjur7XFaBxR3L72xYZ4Ng/7ErLreOdR
MjljLHnwif8apTvub3w/2iImvmQz5iZcWCe4J4OrbFyYu8MhFWqJkGUBpVslpEHMnXAaPG8z4UYe
U2g0mqfHMtTWLq/goSUAfNZHrpbfLXZUDg5CMqVq1XsJZzunVv2v7mCDg+FEvtexeZhIqdW7YD3X
RWDPopRRQAWClvg3MY+2e8mqg0nIrZBG45YYkBYKWfgHR5LboItdWYJtaMb2Ki3aFvOFxA6dpoDM
mzkL2tCndJG8EQuAZJ5uk+wg/he7QJB/VL8RmicQdQ8ufmpSuKvJ2urGkGNzYHommnhQ+9dIBrIu
aNw/nspaoJ/AoeUAP1pTna85DgThfTSGqmePtfgTLN7hWGX8uZNpGt/+O78kYdi962tVoChAgVj4
A9LkhkDI38rBWQCpc/dCFewJH7+xc2bPjfaFWQeHLmUBI3LHmGLSkeNTc7HGprYJkNSoRdIwvfDj
Jy06Dstlw7FUIGgjhRVx9vAjXAWlH8PRulZHmO2sKY7NKAlCJ1TeVA0oIfEPV+tn/hzpsqLaKncG
3/2sGsnarjk4RfltxHKEkyZzXFHGLeSLv+rV2RO8Lzvrjb3ao5PoVQSthzMCvNMCvZarDJzgEtEB
DzSjQfQYgz1CadHnrLqaBfU4ICafN/5QBXHTuxhC/09TNA0tTF2LHGQb0neynZ1lHhzmCI0Jw397
nN/PT5susyMatfXRMMGbp2Z2puU+wr8Uh5WsNc/vucVPCFpTWF8I6DUqg5C+PCboQBxNgb10TVdH
zLJE3tVLHBAz71XHMs8flBsUHazTfU8ov5tSyuHyCxyS+4sjanAzzg1Ev/+54xp96PbaU1FYs49F
CDp+uw06ra6VMyQ7eX3A/Fv6uF3FATWZjOnnhjURiXRA7LqUmaL85JQpCR1I8h0ZZZZlyM9vRdmV
+xUD8/OcDar8OzdXb/5ureAtpk/Q3hKI2LFbm0fW98x/1MrTIUk01i/HKvZMwPBSPGnugdJPGcf+
Xzh/WnR+8i3NHwFGnViYhKdCMLrIPYPFErnb4gnxduN5Ri3bKh3fWQ2HyyfgvBAX594iCj9Y5RUn
AJDVXfQnXUamD591rbjtM9E1fHgiNyONO48QA8ltG7mOwuQ4od5ON8XoHB+HLvepKOsYq9jt8nSt
ySxycbvl/UqWTx3w0grrNKDiDPMpaNTKPecNP549+sqInbruhEgwskLBgSorbE8panlaVq/3WZkN
PZNpxf8YTqY2s09+fSltUpDhjkfHOhlckkmNrWVdUfoo0SHEMCi4ONdaLq+pLtNVQer1tmdOt+WM
BJ8m6lK+Tp11CMxlf9znh5RE2Qv91cz9jB7I8E240P000+irwo/vzw/7KRJ5S1EDUybz766Y9j1F
hgNgvgyrcG3s9fQHUZduYgAfpWtlTn1S4fYmaq6RXFVVHgWe0CnvPhp+McVBEXVwA3aOd+YTFmEK
0lUiuKIyuil5V77iUc3V7w+aefVosEAY+vjIIbDyq7pPg71j+MhPvh0XKyd3O3ZnIX8DTF18ToAO
1aFG66IqROEpsd8QIgJD+6Msn72v5PNpKctlSQZMATrRP54zehZsSBPnJwB2joHhHX1kZESYD6ON
Xqt9i05P6Tp22lXgXEfgKuLidcQXWP4ql4aluRSA126UUJDfpmAn9/bOnu40luIyVkPND/agA7RC
JUJIo3whzGGstHmNL556VAwsP/ExRFkt5x/7lO67mI8ZmvMacklnRIave3aH5PXz6A8X2MEqLN9K
9bzxthuKhhCwSU5m1Jh5txE0FdZrlMqdwVuntHbygVuZPNzXgy+p9rm9v/r5s0SfD54ROeBTtIih
3qotLSVcIj8Z24/zL9mDK8Rh8YnIU8CjVvhFN+F+tChmRLBUOGtdmEIkSb1w/Iy/PDXFfRVx4viQ
LaF+yng7tY5O3YB6cgx1Ua6/zA8qpIyF25p/8VnUCSw4jgriUwPHUjw0rXXaycwW97rpWgeh4Rs0
pVuHnf8MNoM/e44z/vKONCe+04XP2uZTlx8lhxlCQqIunmSUkVkVpOgVUZhx/iETGsMCAAb111j2
pI5tlDcGvaz1+gM/ngHxYlXEf+YqJoX8Uc33gL6b0SDfIFkwb7Q/liSVvSsE92lMBQVDzbNWO8YD
Dy3i95315wi8PGSnlAl4WSspG3t6CQ8RGDXDD2l+w851an7M8UJQ1PINfORSm4mht0Cj9LllPzQL
9tYzAXv1QH4gHvNLA94l0py0Bwfl8QnOh6bwdT4gHo04GbsSOuGFkp2y7iMd1oHw0fgc6NYliagj
LXT6My/btld5aZVXqomTwILyWjpII09pZEmxyc1/SZf6BMDEx2F0CRoFXV+f+DRltbhXhJVdykqU
WIidPXI13USeUIVO3OLqZqm7ZLM5hBWOnGuyMGSP69WcycguGWQfrpjauyPjJmTYfqgOGnT3MWEa
WKEFanyP5XrFL8ReSkXhgoLsko1uhIza4hAWd3eMCl3iSU0XCJgVBHVvH4SjPptUPbfQNZBBaFbc
tdXPssnQwcuDDU6K3PNrfzW0Jk6rBstoRWgkD0CDWMPzKgn0xKe5T6CuNpdgfApOxwwY5zIfgCcA
ESBkvuhmdpdt3Kmtz4aEKEXpfdWnJhredA1f78JOEYKhRxdSVOBstTb8Wbp7wSfeoRXI63r8GelG
nAibJy1QObQHC4SwoZ2cZ4IuxTV8WpomXoGQ+edYoKf3lbFlqfI5FXoOXbwuLiXwHPXeGvloAwxJ
BekiYSoM21N7tNy/ycHIto5Tk8NcR4r+aZlT67yx+Gyww7z696Y7B42ru3F198Iin7zAfqmaburD
GZa4n+qyDu0DOMsv9apQmYGf2up/UHJKI0m1Qrf1wHSXUthsr+lXiY8gilwH/bNVWaXDCbdZD076
A4WMOVH/Qj6BC4ta3pBI4DbwVsok8OnQoO8MByE/y0jpBhQ742zI+dP82CoVfuZdGnczQhCCqsJI
ACZVda0eWknaqhrF+6F+6POdiNHF1SPls1S4ZI3HWl24HnROfTYQGVq15OCG3VtWE1xZksj7m2IF
s2EYpCQUuVzexoPdJVib+5gMEOrJq8Uf5oIfyjAIGmyA08+XBfca2Qk2K484UhtZFbLJpXrRYHIT
sR6oFc0jom7uU5rGF+MYosm4gJOD2rKOmZY9uTRndA6fdOM7WoZRv4mw8cV+4+BtdNaMJyw1ME3q
EOfbnx3/O35Liji1TofmNXtIHhslbk++7x5iy3fPxKwH7IliIvaCq7odjzJ0PfATwCtJTM9hpGUc
l9S8oSxMWtYj2frvbJUfISmAtJvCKH1nGxlEKsTidOWRrFgaVcqvl5A/Py/6qopgCkSbsQQ4ALCQ
sZMFt21Ffcs6J0DdDWrKn7H9Uo7tgy0n1rDpO9MsC/VM+Ufe7EcnuXMRebGREuzVx/CfKxZAMqra
JYHlr7Yb+wvWdNKAiQlK1HRr2eRqNlzcvoK5pVaxQvgHqrS6r08K9Hixs0Jj1lCKsYdWWozYtv0j
3yNJ2UOWOZcgBfvGvd/goykdlPOXwf+zbj6YBcvO4T+20NqniJDgvuiznH0do+Lep8zK2a2g3KyK
+JG+qRr/ZOviI0XjP3Y2YjCgfEGMk+u62auNb2zlmaY5Dsxw0WIh68MDalXMm2G7ApxS2suWCTgU
dmd+2EMVbTkgztNvOAIQaI6drzkUXgguLsaUB2rFIOwEbs+jyUHdmDAkrby1ypnUb9n/9wYlMdSk
Ebk6XJwEJad6OyLKe0zHP9+UOJ3slhYwZGDd6ZXyIV5tB5ItziA5W7M2T3DdbuJ2DALTUfFXlH7H
vgQPYOooZ/72cC2d9AjAM0iQy++i7/NzEOVBPP8KEN1jbUKHIh4AbItvTiOsfbbwzhIgv5PGMUV9
xx0G9jkr9j2eQuNaNQmdkcOUh+bST7nCt1gNQdUAZcY8DQIQxoZDV23ikvyltTVBhQclyjLU2PS4
f/MgwbEBmP8mMBE0D1VnmxYbPMn958vE5OpYGVt4uSfngV4HfKfkQsUe2IauyIbHf0AYBMBBOMSn
VKghFX/h3HkWj6rGogJyvpvppnHHLCpNLcvxONTEr5uxATX/RtpXnHtiAEcJtjY4RNLa90E2D2pC
LSZng+NUMJVwm0Vnmw3K3bLpHk3kfjFIiY2p/meDjMe05Ta2LHIlwm6Q4EBNmADnty++zlijXoJa
TSEvEuoUvb66YYvRGMPxWNIYgDjXHmMEkPkplYbWXn6TV1WchBEhweNu1Ola8GijT85fWFI0KGG8
usFHoEElK2U1cku7tjYbGJjrh8n4WpHwgBTION0tOm/NnKPUpCFsutQ9B/i6V38g6w/ioqA01tG4
jJSa/Bs2SKTebV9NNQ9oQ8nwZ53eFNEbo08lMyiAGMuVoQa/TV1kv+HgrJKYSuGxrFruWF8AqwVs
sNIOrAimMTBqkpQ0GXatrZTT6XKacXyqms9cDpGtBznwBLs+e5NOdCcmAtAlYe6stSKBaRYs7p45
RE97XF4knbM49wMOKU08bS2+xeUK19U5n2Qgujn5d9bV26ax+N6lIRZwoC0kUFYnXe1X6f+dduij
HhzlQSGbnSDefcQaFJAnY76Uy7RzlaEu+dOlnXWD1jqwEuc41V42/kV5xj9CrWEDzOkD2Gwp39Pt
ir78eTy7XzPimaGWXh8/Ag/w0gBcH/e3RS5atGDzKXZN+m3RpsXasRGxZt6LQ1//6rbj781ZhOn/
MWWtIIXpQUPBx48cTFKSnIchjJPX72qDAUbop53oOUZD21luW2BTruBwiMkiXYbmNVbHN6+ACu9n
594l9qT4L+ijDcIY4qWyDhfbZMrpXubJVimz/seiT/PKguF6zUKB5uWv45KqjXxklA4PzJjZZ2QO
DkOmbrYeBEo1hndOqHTWMy7ddFrG/zCvQBFbi9tdxqnImzZaM8brVD94xv3Tc6D9J3Fab6qu6qqw
FenuHvyxF6H3pPM2R/tr0/CTNNIK+wMOn2wjPGfq0TiiFlcwCbofNLg5qfJXuFVUYWFBGFjPrV4d
fdkUJTimHYoONs2hrDf/MHca7VUT7eVWKWDTTRkQTMJhIpTKbkV7GOFnyQioYtWZEbMaPMzDf83A
aghDGugIqaJGoiUK2hvU3VbzVMjAGDjs6couOEW14VoB/V7EJP96MZK7AMG89V0A/YDnPcrslnPO
hpNOI6tjaqQM9yZbS5rbFLLD1d2gYX41Pg7XxA0jKjFLrhppt/8zhRD/LaujmdqkSH11B5PLAx6y
uo4QhlpJxgSI4alOVwVsF32VZGnXnu0jnO5hmnIImpjc0QOHpdNjDw+8V5YugUFXI7fNEu5B9o6r
4N0Wp2nr33Iz5erJErbAZmL1JBBm6DSq00VlvnHoAUKDIOs2bnxzcSne8bd4l3NKoXe/vPpIQDNf
TkmZfm8CWvb0HiuTVyZSGR6yPoh1Tpbv5wKHbjIRwjJyT6o0KoWbbe3VfJEsqIKlsyjTlQAGiQPG
Qqh3ypEAYfIYQZ0JJNvLE3oEEkh17cN9vt3Ghtbss+0L4Zt2Lw+yf87422Ej5YqGm9020xplhEAH
RCSzdjsCoEniCc1IRZx62I1PDW40sjhqTQZvEu0t1Kaa3SzT4zip/zdPHCX98wlxE3JvR3SduWVL
+cwG9jXzGBkdDOguKV+PxSPxiyw3Ko4ExpSfdL/w+rNw63mobh5jFf7yOIjFy92XQXcAk08ZflOB
z+ZvjkmBWt2eC147zdNKuxzGLm6vKjXWYrR6TmS6xs9s5AkzIOcc9MISswLpr2NGAQnfyh96k9Rb
SrkdZrq5vxQCP4sYzU5D0nL1u9jmh74lV+d7EkjZqcEori89qp0cECT1ZTVVIPq4177QETSx9vbI
VnV9TecHpekBWYhqSWa8RvdVN5H30/Kplmrj/8CvcAwdPHxZe+rlWpAYvs+HLFoNJUvGoZuupygt
cnTWXeIXFS1ek25yMqINPySD8uoeMn5ur6hUFkwiHtT81kh7uaakIiyDK8ePUnPGqfWzFWuuPS7Z
73ogymkgK5AbDjjSL+RfNSyGrMMrsCAM6dBJNzNfNHPbk2OQk2xfWw6hBr0cAdGFSloUErjthKiJ
230w8wP5PIeAcHviOP4ijPOk3q13O1z2dMFnwxNOs4119jetxPNnedrF1kQKPaTzXwOVxtmyBA6u
OvsNY8VOgY9XrMLvzo31Tm+4Ui3rWj6sXlS6ncCO2SLJLY+a2dSGiTY6jnMgGIXC+o1TJCCDg8VY
8gulybkYtWToMmRY9xP1+XtqoQdG0wxNr7B7ucqtXHPiB4IFReHmUjljDC22B44fi2z4OtCBV7YB
GKf7J7ooON+ELciqItF7XT35aF474S5BXt0GoFP355jDEJTwG6zn3M/Bszy1uKm0DaY3tmZ9ypl/
4cH6yKsZJRMaQe7x6M3VRoyzGDYS3ay6P8A2FaRVFPfQU1mN/rBKsk2bKVWc3NwoXZIC4YqVMVt9
4MaFIz9LtZYXvgnkMurggxmosV4Q6CuB6FsuPqgfkxTKjq/KGGafNuNUpOFDP15CVG7fvD6fb7dj
I0CdkKRqi0UOaQDxaz3rUuhTiJZDeMy6RSkyMxiDGR/i21EZcyuS6lKRE+QAf4j9UNPoDhFNdYGB
x4+TI0UIeKzBz++Xi3akxECkh5msRKyxOcgrEiPWBHhmhfK37iUT+K7VX9PjCsqmRq+MaY8VDH++
9uOYsIC/bh516r+oMXzve9QhTiwFlJwBypP2Jpw1vwQfHCI43l/1bqKVH3+Fbwsi658+XJV9JBUC
eMhv3mtq07iHUb+qfGGCq/v4OTOmf06Xoz5k0iMmVXaOH+Ucjt+My0syNoB+AHdQc5i8oOZ5a4/A
OtEfEECcG4/iCjkTvfJDlBCMRC40ecJj7EC43ILD7z0rbUYfdQZj8Rzsf5blL4UpovjTgElWxr4b
fDW0OPmPN4oZ3I6yKCHsengYfWS/nTst7HO5iKhlMYHjHId9GfmJCg01PKglCJUtNyPuUw2WBK5K
1G9sNUoCxZGWgX2BYIDKwvKLLI5D7fQckJNgqD9auWKSPX8kkmAcXMdhdok6KmnwzVYePq6zWhNg
ncngpP1l+hl3sM/4XsxuzKMfDoho0XLgjnWQDc2kCC7jAUCoBWGbGEIZLQMh+q3W8CiSU7N1cWH8
zb99J8h8PE2T5kS5TpXYOa8+BmMcBBTdqa6nzK6ZJAyUPsKywxAUNdirUcIxxyhnkiDUy1bnMvkH
5BnM0V2on8t4F5Ipg/GYlNPjH/6Jp9sVcHWOmfrVUmCNP5EZeVmGYVuVz3DH0mIV6tTT0iX9qG2F
dURHdD/nP0WJ9EG7Zqs95E3gQ/xBbtpikvCN7XOyibHJ6SFkBL4R2OGKmT3iYJz3Jqs02GrgHEMX
lDN58NsrkoYTwQ4DnQu5ufjDDlSLEtARhHtinn3ATQfu7SFSbzVRYrShR7KeEE4YIUcIeHfkRntX
XESuulFQ8pHc7Hgw+xSsDCHvzQ/tFkvacgC65IDMGq4xPxsJgXDjUWqZ7Sv8pfcBYxzq2oFFZaUg
0dee8gDtDapTsqQdzQA/NdW8P0C9lEKaRl3dijIc/6qlsGrPJ6gMgTgxVAbN19bhe6+KzZOjoCCp
cV+6Yu4TvKB/UTSLO4YMiJVJ8Rr+ltTuur+oSwyyCARcDg+TmabO01G4mTZUCyK5KJCrqMWui+mc
np32vFbEv9oZMthZ+iG/aKBKbPDr2EAVSy2CdpwBaxgs9omrBw4TdSaBVbr9NbtcMcY9kZmKgVV3
InrQjopQVhQpIoGzlF7MAgawbT+w/WUyQLqMNTE9VGD/60FTPS3fAMDuErSGfyw5D1q0gLSHLp18
8u/yygyxXrAj79KPUH59yJYXruv8RVdBA42Kf0BTH9watO3CuxeIAJ+EB/fVktwii16Z7pHM6os+
dQlLHnc6BcHz6kjflKJqlgT5Bx0OhzpYSThO2urUNfxVb0nrBmNftQLNq9s9YxcXw7/MNhTWtlOY
4MsVF22owz9BgwsNwGzOAVeOuv8JD4Hhh7kybjzbzvMUucbYWGhiQVHnDH3FdtXtq+7NhMuAB0mR
MCImTz0TpW8jwkdgNKMrvozlAaC5zAYdthxTX8W7vIDDsfJfI9n3NYXC98V0qoYworV5UnSmfdHx
nnQBCuM5zRxscn/kh4AUXesSF/JA5jo7mZjq79YBp7y/PIGKuGsxKUQWuKJP7x1xXsDW51A8PrBF
7ycZPrMN4F+hQ8nd0CGXDJEJXmzvywjQNJl5yWfY4/ZNEne1Ku1TYgr0ubraHHdDhrzuJVnut7jL
vQMR8XejLOM9ZcvbgSl1Oj89xvC43Q8AVnyGs8FFz8kvHhrKopPSN4dH2nJ2GBdjta0/e+RRduo9
kTglt23T76of3ES1C/0xLCmKaSpem2hIQnqw6kt+b1hV83OxQjB+LNc5O7EEVa7u7pSIP9cOoA11
VmMyVL3TLW+O7WX7S7AlHXKDN0z57HMXmMGbx53ReRNrFfJgPUdNSGR7S1HJ07XfH2NKI5f1Cj5R
HijelNPhkaDyGhQHwp0OEoHwCmad9S2MELyH2kBaWSZ7IU7eDczidtnnTZO7GZ8jlV2Cw6tyvPk9
OaErsbiZHOCc2SoSQhQswBMYcr3N0ESEY2jJn5xqUAuflAcxUQL+HTnEmVXUR31yqMXyBmfoC6yE
cyGHBYxH/+Bi0eB0T+fbyDhQXxKvV3Yi1eK0dFexfXZ9/TFTugKGFoMVs3OneP+lYaCHRfLYaq7l
olX/KeUK9Nx/Yp+u3rl6c+8oW8l2gIWj5tSwf+qvkQitck0RWM/ObS68uUtVDhUe20sdttyCR1BO
S+FnlYgOGHPO5EmovuSfRMsVRlWN/64n5JChZ2OKh8M83nf37pStYvQcrVSQgdUPn+tDE1DessjJ
K8kyYayRincTUzaNms9/bEpJxKZxqt6bWZjg6bD/kkhLGZdbqE3h7ydBbROp+cb1/1r20upO9ZVd
2uQI5AoPvWuCC4Jy78bRIxc38oIWGBO3ZbneiV0XBgC03W8ijYMdZbNdp3sp1GJ61UCx1dELmM91
2S7SuBhBp7UMMSc9l1lzE1/eh9QuOPzO3mGOtkbFmL6SzwEVVbcEl39yAUoGerZBvyI8pdmTxXXE
/ULFYjgU39mJId17xEBcHmvMr+fQgq4yiZ7ilwEGDldJoto2j67IksLWcC4WpAx5cNXl9TWF4BRn
XHYaqFhwNEn58Zr/Sz/9bsDA/Cj07ivMxVWdQXidh3yvQ3LXl/zSLmftILumObnDkQzkitOI65Mr
ZTx3OLky60oYbnSpINnLklEgwprA/relHFz6nQ/vkvN4kHZB5HO5Pv/vmgIRHeMoXSSXHmyCm/2p
Togr2MDnmPyFyyDdE3vpgcxnm0NSYK/qJIvxxd+ndwfg7pLuoUwe+Ao1skcwRZ7BcAJGQOAJCAcJ
8DYZ5X1ILH+GI2hfZFvd55x4cv+z0yEBJV6O7BKyjLpPppIWbvKd/dELKc1k4oZUn5XDt4CFq/te
sr2Ebd3T0gWOMc3v3kQAXdWq2mmrjiArbpAwdru2FX1ve9bPiQZ7FDDfG4Qo+gGbWMcZ9dVeunnJ
T1WJazRYIS19CozAUwzVeqEWLK1B/qY1mdE+uF9EJNOQeFB4sYH3WylYpCk89kXGzVUwwFm2FnKf
Smrccai32teLKzKd0slSnyqMi4qyU+Ztn0TXrrmgw13w6mlZYLi10l+5QyMzrJnSP6xAqaYM8HnD
exBJjDN+LXO3t2eLWodzG+e4uere33gtS1vIDkg+YEUiwPkGyYgjFHY8iSdmIcEnKeRkmUK3tIIe
xmI23vU57DZd3yJo+5DaXpYqNoSOSr2HyRxm88dzkLPirCF5EQg4iZhUFmZFncnZ9ic25TZXm8Yt
5lpbxt8NIQmaVr82cl2EXywq1DS4w7kPHXFYlwktegpWhut+TrRLthm2USf3JQ2Gard8iwi4/N3T
Wq9NFE0R4m1iIjZ3LdlY02QkxRVbMcttq6/FS5HQKUjuQEWuhNtvjEKMoX8gVB/RDsqRBpsf+FBN
RcUDRrt0J1yROTPSSOxxIZq+shzexPm/ZcqhIwrWYCdBMCiirX+/qxIWijnzT8GMXM85o9m4RIGB
Sx64fFIGoFXtH4++AvyL31p/xtTFvKsAPPSSBZ007wuvBCR73TVaZirowDKFKjSaYDvi5drGIxLJ
h5G73Qakz0w5Y8QowPo1KfChtUhXsKShhheED83/g/ePGNqLWwW38NcGfhduhYQexVjov1A+6kL6
QdP7X/5PMCZhWMYmFD/HuDz4qrREOvxZITQGpEGHdRNRtwO9WFtoA73LBjVQtWD/zXZZnBSPx7FH
LL00wlRAGwvRsS9VX6UYcnAdcuOW//OX+IPEAvTuwuTsBCJsggNPfYHrIIzS6jWwyR4si85j9vGJ
HzJtggG97XhGx8QFjhQ+wdc2SR8EhQ/slBD8ekJCv6WpwWGhcwZ9rhk4/QmPO4EpGUrCk4NPgMVo
VlQ3qNFmNDWatGhfEa2kJTKB/VqNR9ouC3gQ+CxpgT6EoDwIVt8WxK8+vNDMWECt6tBseJahMqhf
9p9NuoXbmjixAzEYq8MyyIlPOOXriogQI8C0DjVfix2liuTA61hhMrozaXY5lzo6knxBeYRbQbPf
TSDO03xHpZ1hwsB7439rN3x8qdC1PwdZtUhCDuH1p3a2b6DNqhaIGZn3YuNwc5aOrGYpru+7CNx9
x7da/TRjXC9DYaBlUD4Ua9Q7N1W3RlgO+8yULN5aeQywQhcLgcTQpRsO6VXDAYyKr+pz4QuXOUsD
i4uIWT06acbpbZAsHRUky08lXOcq7krT+FWEW8v53zrgyMiM4e+qzfztBk9viyhf62/0KFyNmht/
YV+qAKaasoprOiMs4OBTxdp7rFX7hmBVsTkVqspjQyoUfrkhc8j0eor3bWbbi2bWaCRxUjfDWehg
bqGh6jkP0ukIe7QFHN0C9z/OQjQ831a+npzlB3seX6CeuE71/eou8cVetze9ryup9x9oJvTZDI00
agGVAUzDggdX9HgEad/GEw7QwGw9URWMHg5bBftZn9fgHoC/IwEYxZ2gTeMaLmSOraFMt30dxWTq
3c3tEnoneHb8dQvJ8QaoC4gh4geSjXX2UhKMUsahLFkJXp9XQRzkVxgYFtQibloPD1sFa5gpDybS
rqq4kdWbfR/7EgQIpUJudW7GJzD71AHJ0A7vYJjGQsX8IPb8NLehtkDhAxIXARXe7plOWMDJfTnQ
EIs1cT3Ztw2Zf7luTBCmkDGHt4aUSb4s8Eq7FsNK+TFHY4Crr8GiBJqUM66bevHstDQxTkO80WuL
0tTcgb0m1W+fCB/S1ro+OxxGPo8JX43lLbS9p6F0HsyjIFy6YOY8qoFLto4Np+ZLoDfulyWMFJuw
ylZ2Zn/oqN8vTX2/kb6RCn6r1J69sqRLA/4zS3FJMH+6kvywzG86U2WP1zWRqKwCUGEtDHP/8LEd
mIfoF5Zsf+G1uGz5bo3FyjMDw+HcAzGTC9KavJU4gjsJIoZ2YAtaoJLTrIDmDBesZR8O1HIllos0
OyqtT7FATU3LD8YShb1tJIh6DRUsdDZdFSbGO2cK5ukGL/OkPkaSOKbj7XAgDKrZ9bY60HuYX9Tk
sotjtPN4nemZpXifZP4huOCrmRBs2ZgCxH+jfGBLcb49AQByjRW/F+yyqmVmICmCnTyAYqHS0ZG9
gCb+EVNaJrYxIjRqZ6OOgkgW3QbIOIKF00Lko7Nzj/wugBfjIyVK/MBuePtUJPhtxAyg2APZ3Eie
EkkDDeC70xpS182xQPEOPmqEPqepwoTPTEm4Gj9U2NJmpu0lkAsFh8T7Pec0qGVZb/OGOMfcp5Qc
+k6RCRrJTQLls/hUZFVUx9TGiwLqdLRPPvUyNvZ+JQfWQmBB0G5C9hk3QkbTZvmeyApK2nu7Ef7s
OdNozioCmr49AVdHz8qL2Ws7ftDvthetkaQjtMH6Xnu4nnQOkNOvR9mlSvLAzhZ0V7x1OnZuE5wy
QJ6NvUCOMi+i6Lq0FPDgYJhmxHsETnp5JnQgYZlb3Fnado3Y8zqGKB99bmNKNNsxyJlEZquJQMRL
c+An8HQnhQ3T4xzGUZNebs0whxmLVw1uJI+tGIHKi4Nj/rnCeT0V0E3CyyzmJRhbuo9r6cnnrNxl
O+QGDUNDPu0j+wDRLGvJG8x7qyRQ4wIBMSDFw/WUvzJxlfJw9Z/Kn1xld+SB6rFBdOIGgjiWDh5a
nc/fGkgVwJpbrjAnJYdqLFg2vEYSQsc3tZfMiF+d1RcaqQcZLSdGp44X16SQp0BGThklzutD7Atm
O8kNXCQjLqZdia6jhc0DECqZy0Gg/8zIqesSVdnhPe/x4YVYBTZjC4ecJ7/vmHuFmyAzTgBY2iIp
fpEl1ahE9Ax4rGnvnRFCUUp2z6tuMgbgxZiBhHBqv5YQQlki6M+0zN4ZlcaEF+VAj7dglikmb2u0
m0f+y4xhy8ZIWCteYpu0gbSWbI6/2N52C1Vtq3RBvYYLugxnCVDrqAJQ81L78My5NbbPvcMum9E/
sTmtPvKcXmlTbGU7/p5xkwEbT4yt7hkrOaKtDKKHuyx6Pq13is/dUULfX7qz91n++VXnjQ03SmIe
KBge50kCXMynOCW7cbRXo//X8DvBkvO3sGBN3FoTdJOCFXnqOUV7lthE0MqGGBhlyZv7hKmuEAuA
e9Ye4dE5ME2sr/fj3sheW9pM+LDJSo7Zc5cDePTisQhk1FjmuoNqjPr70V/bc/HMVS30JKx2+DZ8
hJrJ7SHPtPNsqRVgqZ50Q9999f+L51sI/svKxKqTwrwq2VI4JVrZlQ+o8L2oBO1fP46IrrDfbdPM
TinhEcynHHwXedcAaLIqdi4AHO2fPzzSXgDd9mfye3aZJyZOteJ5tt7DPaJZVAh2to1mRR66yVeB
fFlsX3Gur9pqRUZweo+q0hNOf6EzlCmJvbUEeGIJz5Eb6bNuSy1BqI7cfp635IR7Sfo9Da/oNsEE
iPXzWaPgyW5XNy//r4eeQlidVThRmBwkTKD2CL1xGLjr35Dnx8PdQy6qGSBxCw2SCkl0kTqFFzId
xsYXk+W5zGZx3VVP6dw9RX85EsQYY476pvEr0pEhjnHBvq5AEojLj5oUyKuk8Tt3p6uaxF5RqdY9
u4BHOM7DQe7fvBMBU48le3eaGjDJttMvM2PjD9qSzZ8UnTXe/rHFp6g3cCIKlW/9T6ptCnx6y58O
NwAKijXa+CH7RYlH4oAtXt7h/2H5uPId2GQPaayzn2peTCyfhx4yrOMdMocwAO8OAUXT49Kq9KCU
B8u586NiADqNKldp99aT6LGf++xhzInKi2XXuWdNUQRl0jDpJ3bk8BDXOMI/go3eSq4+Pfipwdd+
aoAqT/o85fP4fA93CX/9uxP9snEVnMPtPpzVFTwMb/GwAA00k+qsu7yctV/5RRXrPBIM0Bj7sUs6
WXA7JmPwMNSuQwYiJza2KXgyZo40HExsgwyNDHHMqDnKq9RjAFWnKZ6bCmYzB/puUDRodETkRgQz
IgxX6fkguXchPiNEThdC/T55AhyLkxB/m/FuzYCPyyAL6OcahupdCF/aK9UbusYZQxGnpVNyEjnS
gq5acSAPEh2JmWECGval/L0UIzNYrDRmwlNBgbkspOrJ6rGdG9K2t4KfA+PhoZVJc2RxvitbhHgS
a7PYTvuJ2nC4+G+B8Sc/K7rUa6CyLNN9ReD2b02wO/WPvS/BRE6zXUxQRIlABNOFRsUVIba+ed6G
gUM+UF9szUxw8bm3vnnmT6qqlxQBJFP3ONjHP+a4/Br8tzGhAQunrAwVcSlZ/dAGsSatOBfXcXDc
CLMkxyKc+GYZR8mwjBwcwwbV7kiA7r4hRPfqBjOFpiJ/C9fOJm10QDlKrT9HomlDmGv6KVYTsPlT
pIH8MgcCPlFcWyZRTVDp3hipfenut6h/dTFkDNjs2Obl7zdKv2bExNlYg6Tof5g+h0yDbgsW82Vk
D1ihFkgo/lRONq94VLVwBKsg/+HTWPptmUvL8yW8YwBEpl6Fyy8LBquTOyo08lEqKOTiA2eNu1/E
gTl04HV02prIGj0bX9I6E2bo4EMZ9nm4RY6W4o5/rhcOhrS4NJyKadFYFPLAN3t9sc7zB5v7erwM
02t8t51U3baXnxNTq3ZeNGYEZ+v2hD5Sk/GuJjjv3MdypD0eHVld89l7sk4frB6+2IW0Z/gOIWmI
LtlP2mIitWxylSxi495NdbsIcNsTDTFRROdysMlmpId103zhFigNFFoRySQk9GhC+QDs7P6tgXPr
IAPP0jNARKpbC+6G40J+5w0fbdfmUDrLg39l9C+AtT9VPZibq3N7+2l5X5YBHJhzgxWnvEICHADd
ariD4g4eEgvgsKc8imAN+iv38S7NBecA9Q55KMD3F+SwzQ1EA0Kqny0DaR9fxy5Yh0CS+YW0+T/1
1RI5E/FpUNX4kauIXUeUYqIVx9djYOjRYOybjbdDckKcd9Q7sQhmZRCsb3/y8S/woKjhh3+6bneV
RwHvG+vHHRDA97g+3rAVrqgczLQFYlaKTiLwSoZruu4g1DwlZlmO+V5WikZA4cJ0oupj9jAmT9kM
U9KnzfNqutPPm2WvbJwu6060yEcsue/3WXRPmzBgYcVz8eyGnyLx6pvLX4fYEFJkrXF0jnssTJ/+
LGyezOV9In5iqBNkT2LLujnKzcFVYMFFvx6aVc9TayFpfoaq5FefAgJR7MGbqNHv1OYspT4Dq246
4kZswyJODrogKa+KNTVRLVPrv3t3+pqxO2YBH36vYy9HOunWaDNsrZRO+SpHzzqHep2NUyQxCaVm
Eu1wcvi16OmCE6AKqdlqc+YTOdVWV4oErw17ZTIPrE5Cp+m1ZLXARe9d/4dSdez9l14gBRiDYPKW
RNjNki5FJciS3Ls2HrL2++d1aYP9WpPCdbjLUmEdDfGfBk7NCktczPyYbLMBJgKxk17z89Hh4FzU
A+9hYPj1I9PTr87FM1m+WK8RKYWZGMtTyG82bGKH5HlUNj/bm/v+eGYRmnaOLK31vd+9UOyJp3qS
xx2x3bH9twVgIFUMlPREqneBSLwC9WGfByW/evDCM+NjIcSGZqfo2uIHF9WVco95eAwt5DBF4AOZ
QxBoD+YD1Dn+7NGHyEzev7/UjyL/cL1UCpm5dTYdeRM/a5fKpc1Zsm92HITM1FL0wTEmpFdgV9+A
diOt1CMWOZukY/0QqU6ZnvdNoEQEhkIwDcEheMAZ0A0MMgH16Bb2E8mpxbwAR9I06yknLsyStuwS
cwwL9C4KSTf7GwG8xTuA/msE5osqDXAOKlsWPoFqW3oe+H5MZsdtqnpLv+ljr97XFQDkDcILySMV
HUpTKXZjM9yWIw97KN79pgNLivflJh2fMFi2dkEIUCcUrFFfk/uwSgFWrSrj0T9eFGamD1k6Mebm
D8oeqLYHqZtkYNZPcLzhRUvc+tPdA3Y+2WeuM/CjSm7QNJ1jIlDIyOOpKTt8RDSGgYGCdWNs06Mj
9RCuOPvwd56kbljJoS7m9AhyU1EUhPllR762tWDGlVLjrNyo/1mg6uGzfPefAoANjJMjldqZ2QcY
vCn6v7UoU3AQkeKT3a3MyQHKdnE44L8oHMERAi4qu1r0A4LkkKJwSIg9DB6C60l8hjOPRZ6xwKrK
7avTaV6QcMgB9UlGbv2nKiUffQ+9TNCVMo/XDDd0p8E3jUwB30/Toro3pkYFWkpebJROY1FxD9HZ
sG1iEFA8DcUGWHCqhUd7t1RmeuRZpyMQjeMop1rWB7COf2NWBsA6fWBNSZjK/3UyYu6eegcEyh32
7LlNVzb22XK/VK+knad0hov8HXPfgZwIjs3TnavoWjzrSQrI9EnCQigFK8gPXq+G/ePZVTDIDlwO
edB7HfwQuicAdXs+qxIidZozkXHiwrfgElMvQFKhkPHYNJ3vfG0FdMQqKsAEJ1dKRNDJpjq01Kl8
qEI5fcBVYqCnKAPS5BaVpqTICn++/qRpsy1yorRgERePzrtsSm/FbYmjU4jjDydHenxFy9QKeGWf
SS4m3+fOiXTBzZ7NLSDzlvFJx43Hahu3PerjhAw3+KiVTGiD2b4Ugybc9ASS2+em0ulY0T6YTYyU
PRQ4ws7CPFAT65FSd8+Lep4efTFImp6nYXTtou7e6TGUDUZ8B2OCUkteyskJf7B+JQ1ZIR8p5Z6L
XjcEK3XYe7sA7mYkTZ3txpJTv2ogNaG3c007cueqz/wG7oAjMpliW7P4odeMAJz3uIZTp0QAffrQ
Igptgmyi7JRLce7te/HD9hVDzFiEnbndy36ochGInfXFIsoWvWf73Z08wH45QChj7CnUK+xSBiyz
Z9YYqzTJRveWiamBMBuuEsn4w3jdosUqlZXgnr42czTe5ZXCisOERZhMkwybm+OgdavpUhfJi8lc
jk+oFwOVQkuycRIa1E7jJvhUHyCdYDBx1JtHLJ/wHXAPO7EcV4AZVMr5/uV+Nbz5ExMP5GQ/xmt9
pnf7FjxqSnw2Afv0gGbsRZO5QwbWDHJZpEbrczI6SmfmVwMR3uPBDw1ALcdpo+/aduhErvMZ6tdU
29LMFTiHvXUae9JjPLJOsgODRKvBGzRRISqhrlsEzx15lDOUo8jP1Kz3ZzMIovjZS0xNFpC/R7dv
j4Bp5eysKCqxi1hPRSJBD47vETV91LiiEa0KpL7ekvj7zaBFQ4TZeUqFG4bfJZCNXxi5FXpjLPlY
3eF/ar3cILhfgRp1zsQ7goMALsq/8rAzR78Qnzq17QyVZdL+VZsx3A3VEc9w0mUIGqpkm/YZI98V
t2x+oyMNaT3CIPxyT+lLHDhIzlLl7e2EpLfc/NRBJL94w8QmYYgKXCReDTkQATUiP9KE2/U0xTMz
5VtpS+qn8I270dYI/5Wyf3O1EleG5HX/e8Rm07xzow4BZIFPWUJnpnFiZMLDyUQXixNTALeIVWrA
wWB6F61ckUED0ykFL3FqtOF5NOPE/cULLBYdt9lYMSfsHiRV+a18HeTozIN8w3ov6RJwiFYW8n4a
75UVVkeSvCOCB6/KQeBCz4ARKslArPDahNEOWDQdajr1bA0mLOvjfF8anIOtfNTq9aU63STVOC1a
prJJkAG7WvyHQPmQmu3XtbNNjKw/tbTqXp7JXAtLRpU2+R7+mZsu8mrUUR+3f0X/Sy4HW1QyzagK
s/W8S2Ja+Fs9skpmT2SkzWK2090NjnWYt25CijhcYK2OvYjv5FcRGkE7VAA85HwKG000tnklDEjS
PW0dOIR7sthMz3hrtN+9LdOAj5OYpdbNg71DqTI97eJlnqvMnEBSPSSdOmX8+KFar7oP+d7OSpbd
AcwLgpW44tbvpR4rNp6eMuKBzXHCYI+pzDFPqE0ObaSQb7zxj3VmiXrlKxcMxFaFZmbCxmYOGu/B
9suSIEWodzYlqTCZJSB44xZALs7JB8jadin5bmUxSmZ1u7bxBOYJYLaon3+yPBAbjPxfPlMZFDON
Op6NGKSZYPt2UmKMKO1v3b63cn1ME5kFPCKbZF0qaCOXxSHKGg4LRbifZxTzmvGeAfAjQaDhuwDZ
xC54w2xfkr5QjUQBpKhuqxvOnHLtlwPYXU1hP5EzUXZYNxhcNRQMkEMhSSBcHS7J6kTbkTSECSl2
pPoGwP+EsK6mayGF378SqzZz9GXot1wF8aS5SdH0K/d0Jevi5zBzBdN0S4BK1zjS8sFyXMepXzli
iHSyGdzkitZnub2gVZ5yEQhVoUIF39J8N+TE6WvCzRIH5+hdnETvWpsnIAQ+TJgGSiEu7Hb8yG8k
Lpho780nRwuRcC3tW81gKNVsWj4GGSjp4DO69cV16xfViEv9wuUbfRQsQWtBkK25/CbGXWnM5CNx
UucLUi9xyckLJoaxtiqC1zv6DM96cX2ap9ZLmaBUakrZEDqAye0/Isp5j4HC50bRffcFUXXoMkhm
iWwAXnw5Zp5QQHQMTsDzhL/sHZ1TAlL/pkxkKP2y8D7NJqk36CIKzHK7YNq5Vb7EOuIKVRQmis9r
kKRhJ6oamF2VsYe72G2/kMTpx5M4iXDPmpP+pzxq4i+uaxYo1a+vxKUS0klioiMdG+ivGiIE8sQ+
xKoRr9nyiwVZFOMRVaZoz+YnLMHWKAiX846hbwmQcEa5+a6Io8VUDw08ZX/1l+0QP5FNmBTsxRDz
uZ42qsJgdhwGwnpeuXg3hEE/pJFhpCIxzTRQcv8A3XCvmZpCVRQ6iI0OqFwYUPciaaH+Us24T8oY
ufXNyQ0N7gcNTEKuyvxK5Dox2vNgpds8GHMhB9FXJUUd5heLN2TrVsTzIynwEJjoUDaQ0l36dzHw
ngJKrV7Zkh9tfxUdNtZnu/2h2OYFR1TY7XDuFGVeh6ZlQ+h9eP1XiqmMZC1sARb7Wu5EC7OKHTuG
jXzotYFvYpRXlrsGFQj5Fh9Y1MN0KNxWX0lpb853JAByhxmf1wYA0mEoUlCmoe3+Y+K2X05VxEzR
W/3F1jyBUInRqKuhZ88hOP8Y9kNMkYYYGv6a+iWAutOgYwCcJBgmccB0MZoaGl0sZFYowc3a7+Ot
GJVF4wcCQsDdsj5gp0HElS5Qa9hgrllVljJ6R2XyJVYoJz8NkzPX3VKu4b80nveewE7sMGIHiUoK
yuGUyQTgAJcxwa5Dx1M+gpxEXDWaRp3s0euh+kO2GRTuwY0yrIS+UzkaP20YJippN4lVOdr6N5RC
dID5wmMP2gORJocv7DUCGtHEsqEDnJxMuyp3gpkkdL4lImDqm63tyau/uNCkMsypxUJyJMMYTPnx
yIdo7SoM5LmIhYjLrLoN91uA5mdPAQaNcTLclJ1JGYkqqE63R8V03PiARSN+F2IRctPZ8ufuqJ4/
HJ2zCFv1rNzpRjKLegk2qzJ5A3/EC88ht/NbWnixktfthRs9xd9U+x8KY4fNcSA6slPwHgy41pa0
s7TVqnUGrw8ek/90WDwtGssZe8sYd0+I0DeO0C/setPGdwHXq9aYIXPH/SLip5Sv8vGGyquGp715
zkV+xJKzRbeExV0GMQuE3RX9yN8yK40TInx0h1vdDD6/I6G1YfSFs4I1jjTNUWujm1rcs9ht4IS1
4YYRVAXSJgB1pGyRRrGblCR/8oK0+myIZFyuYc/pVppSfaV3K/enib1+XXRCuIW1LIwLS1zH3rxn
6/OqNuoNR4hnUxO1MM7sgGM5ah18p4iuz2IJtX5Jg2/flLUmtN+Axr/VO5mbfny6zuk3CZ7LeaeQ
Nwl3TDLRLl7xq0SMd6mOU8Ng5rqGESErGtSaRuPdDCoNMjuW3MUeUYpllJlw7MlweHyT0lZIHuQF
/nsz/Dk6lQuBgwQ586PHshdfELkZSI78ptxFiVdQ9eevzu1lSnW78Ze3oliAdW+LiPRIfVKQY8Qc
MQuockVo/zoLIzWh5TAP596HzoEJSQKJsbrO+XIPaTfvl2S0Ur1kn7ULEIFis43QbaTZlhxIR+Gz
NBPskbrTviaFmcqNV5z4+IfQ/d5ahr/mMn1WhlrXJJrz/dNMz/J61Iugm0eVZcUh5wW2wBJtmman
M0La38P1KkdJ/7YcAnepbiJ78+wxqeq2/g3qJghlQAQZBwicrRYixEta11B+Z6EMz2oXQPhGDzeR
MPT1D7ggHylFQAdaizyIJYh8OFXR3yuPRVNWm5M1NmAfbC/iCJjWApbhd5Q6gRu6ORtdAAuZOuoH
okl519L0M36H8dtIMyeAO14agtSXsxfevRp7oCIL2s7qbsZnLRjfjb6ZamU2fWwfldmsGEu5aqw0
tgN7zwmF3QevbUU0dAtzVRy1Z9b0/vI5fGySPP+1IDva+Cm4TP57jh7XDN9kFn+ST2MhTo354i44
JfxBfKUVBpAQdCZLZV8e3QOhwx3KmUSQ6Q8wiIvEAMFKtxW+2oihKy2h4xPsWKZDvO5OQxzTo6gF
p8764r0vbEKtmsL7ASyyGI/Lv/+tjSWmWq+YpYR7cYex/OpSOPvgpHZkdEowRsUrtypK2aBKyRhg
1gLzdZZbmV4OEBvEDYototyOz9TAKSLFMCg0LWr6PmiOTJaqgO+GI0ulkW5L9SkyiH/XnOi2nwhP
Ar7Lfu75iUjmBlaTuptC/kPk1ovDluG6aEfWXI8UzQy4box/7xn/7NbVryVCZOtNxOKc1CPakvQ6
Ek2xuAb7CNa2mUCktLzwk+I/X4Is9Y3SQ23cKHtj2ONqtcTANAl3f933sB7aMrgInxLQ95S149Xy
K8nJ/LISaOjeoaYTCzLWEZ5p8DZA1+1nSMPt1UG9tkdu2XQ4/oeU3KuBQvQG/WF6utxktMFBWKiA
1TAAkiZsJ5CyY0ROfEwYKIgXwLJMSDTQga9eA9coTYltrMgCbBFhIlYr6cf7KRy8FQbzR/KBxaue
kloxoFO7K9lhAe9Z2waVIxzEYPxQgOftrJFLA9lV4wHhRt2M4LuiFK1/QeJLecdkf1PGf7PdRmX2
Y2MtoEm/ZtHUEB2ZLlhhSXg3TlbHSwhehQElZOqVkO8EetGY9i6Ldm9vYHqTeVa8dI4nqvvB/KW/
pkneoBxqcbnrlVY/x+HE+DSjNUy06rFUxlGgFpZRoAml1Dpz0MTvPrWiaSe37632jr/B2O3wtRO5
4xW8N7q7of3gj8rztTpeYLM61wQ0hPqB72iPcRdnLHLENZB4eAhOXh5c1jdtObyjcoDFnhXiKSDQ
Z13A9D1DjfURFVVuWwzK3IQKEervCAI2bZ6LFtV0zqpbQK6MDXezOxBWcFC8VvzUaxRbVH6qeC1e
Ouhn2Bpn9yD/SKrjOPY1esGL/ff7n1sSCT9zoUJparuMbTDx4ftuM6npMzMQehZpJIba+4XvjX8x
A/85zlltETI2C9jnhGam30s/jbITfASzZsnBCCqW31eGEA1vnutHASIJrXnKOJvFE08tp3QWZP0Z
uCHe8B3ZAtGUppSi3+7GIslaegyH1iMkD9G4gZWPpjOH78hp6YlFYlGxxpqHKLuMRSBCYMESmZH4
FVPzlTCAmnlwkvTDtgKKEwMn/M0kX8yimrTCesO4ikbHHkSi6VJn3Dy/QQmzi/iG+/eNGJdcAPpG
i80RGYtYetSJd/2W7mjoPdmgNOPXAaMgNCNny06qO3e+lgQRknTBUBsYSucRPnFO5d+6Ox9kjAtC
kjFs/B6ctD/0D6H86eM1I6dL5Jy3Hgcu/yGifYXOb91raoR2J8fn8GbCj0KWNR0ZFAFO0xwJcOK9
uCHjkw8mCsjexb3NvqeIXsuelMwqSLPNQSvpAWZsoHAYrPU1BH3r+4IM12yRNJ5OjUgYrGbwkDhu
qqPdR9nGd0KTRAmVrDw4GkMFblRrRja3Bn2i1hpkFRF9v+OcILTp9rnCQZpVMaFatM6aKAq/QHum
1teNku1+qvl09vc1lhalaVOqscrQZyDVqgNw3wSZtQYHwHcW3hKQdvBhp4OX9PEz7n0fNJlWGyVY
KZXSIzusFb9a2yjqE/GBXwalciu6phA2wKIrTj3+2SslThsfOld3d+yc4EdfcfJ+0WB6K7ZgsUW3
pr2sUjoosb5dUEL7Jr0hzSbyt+Xpj95Ds2AQsJD/nv3m9NPnRbR1WzZNCbQRkb/qPQwnccSEg/l3
ygvJT17w1B8p4dLBHOu/ikdNryAZcuhaFbSzbsV2pw1fZWHI7hyXgiG6zSLb0JDdDisEw2iJvHz9
sVb7Rw8SSXyXUwGhO3BkPoDbbEjLDHI33GyWmhNoig+Pj3uR9zbdge7MxmksmI+eW5whdxEPJq3k
6K+pCovJRCYv5dZZXXseM5qzLgwJnTfLzcY6tr2u6vSQXoSQdZmt/3Kd8pDLRzxrsKnxisOx2wqw
3JaxHmQU3St38BzW3QrB0wjqfcqLZyyPkaxCFhzALhr+puqCJstIRfmgotqnebYqhvztch2TS71l
KwQm08tPYtOzcrmh0XX3M/WIu7+VA5d3FWNRAeXhSH1y4rwHWh90ANF5uSUfHluBsjw7FmTsZrxi
GbqJZo5VXj+Kzv2AYNt9xa/R/8Y/Qo4+K8vCTDINDKKb/pVjNxBAUMhJd6LID+nGd8zehc0igXhK
gEyalKkFbRRt6NOyf27uhXaUBjq+nL+k+w21YwzaP1EtFEwYO0WK/pr8MszWGKV/Nj+OO7I1gpPq
v6Bpi70PPwVAVVE7ZAT+aph4N/JWh/EXqjQxzhXSRBZSd9ZRH4l/kqtTviEddAp3dwvd6ONLAmVB
VZzs8352GcjnbG/m4F5VAfaya7OWlvxtSAJR6Bhwkzkom/iyoTNv5Nh6NBY9hMg7UHjXX/TGfvEV
omxXxIImIznhUTWqPMOhV3KoJdekPOJmxM0RqLouL+QjOiB1NAD7vRTKkay6iauScx1AuNbTD7ZV
hq25ozTQH85ojEQPuJ4acimC8esP4GJPIgkQnb55UlfjClld1qcM+0krCw+O6l0+AGY21qCoWCmQ
vf8tV9AfBiTqn9JODNwk5WGRKf0vQDNAJy3ZhxsHwj3K/XUJkp1Jl4iLIJCo/dcbkWIE9n/MtKYR
IWM3xJfUlPPIHEdI1uxnR/AID8QJAijdHGMwE1bYBcI47ieAuwu8+BUHz30x2lBVUZ0JUI3cf7QE
WmoAVupJhxmPLPRhfsO64sGDyhLk2doksRZI0wyxEUE1nPa07RCUUOP+KYI57oMXRdzw3bDPQziU
BBPQbH6CDQLADNS0IEEQBThlato0zofF0XfJyrPfGE0jwEk1AfjkWypvZ5lXCtQYzA+Khgr+l988
aj/wVCtEXl95NOIkrJKVN0WwAP0QjRzbFhRyXhKJACeiMi8vQw0Y3cRd/c70O7dLiI2zl9CoFqQj
QET3Oqyfx366rW/yfG1uBZJ4oFIyRYJT/y+tVS6fG41ahqvaAcCwiETm2U1cPIFZuBKt3UcmaRwH
GYqq5kk6Fv7dC1z8sVDm+Lb66bPRTvzIUAeBHFlH3NvwtUL2l5NG2EsQzCtaRrmG4d9shbCIyik9
8tsIrEuzZ1DBKIJmmdr+2KmZuvM6qRNAIkqqqnsMIw0jBXgWiZy85Y0ikIE97MQ70AS5h6o4+dVe
n5OhE2JW6/5ZW5gbfU1JCpiGaRr0IHhCj3mO8uUssqAffGBzr3EHg2NdrtYG7sA9EJcAMV5zTIv7
IdPGxdhlRXhlfIeI1WLyCCrB96aShDUZwMh3A7/b+Dr51sQWchoTEjoavgP7c0UiMR+yxAXFInKT
mPKUv38v+VQJgnSCVCqUaos2gWIbNDWBFAySgllU2iYPE3fAb6cd37K7g2d4NVAF0TuQcaaKLaBh
Xs+XqFobEuXkfwWlD8xGDsoAH6V//vFhVbKDs0U/3uEws2y2D6vuDLjZH8G/Otn3vL6PQokE4E3s
DcrIA8PGSBT7OTvu2EauItgn7VkDxZNQFPI+pvC7EwxGWEm0PtWemN8C9JV/vifJrbKxi8c0SohE
DG/W1iMCWRcx00BRrNhCdGK4H0chbEHgBjgy1KImhBHnxT9VRw761mZSSVZ5VO/PYk/iNTcCgfC5
v+XCAbqrySfULC393psPcbV+VqkFhjbkHLTeaJDN+mxbtsawSvqQW5df2feelj1IYZAtFgdjrFGr
Li9UI32jqYdloP0Wz/a7mBy5wdykB3tw3PLw+7HX/9ysHsH8TBO/7vaDWBWVEhLqgdLnIsGQBcIc
Q+cJUfG3fo+e3kf0dgCA0Lz0wVTVhEG5mNcVYuQYxMnFIuL+c957XWqO8I5iWCXxCg6WCf21Y4XL
858HfvjLpERDanib6FmWndDyJgeFa+zKzBfc8qopjugzcy+2fGaP/46Zo3qAkgUqIBlKqaHmI1yO
QCOkBF1657tGEA1bswDoN+iVt9J4SOaxDGYabBY8cLI361BdQ+mEHs55dYufskXYXuAP03fuS2GG
FkJkxVUM/uXqb/26Z+2DtP9jkSzBHppzH6MDHCI1FRWVxom8Ha0EMwljYmFyfNVI1MmkxjpIfmWX
ru3bqsj2ufl9luH61gjZF7ueP6BD0nh9RuyvmCnNN/Z6SQb6cmqQbVaqPlkrTw1X3A+aI3eOxSSA
9I9naILgtQX17+4nfS64mdB1xPXqhxWj3QYhgU5vDs4bDulA1Zehxpwryc5Y2UHLhDvG3vgAZFtb
EjM1oMAq+aao4lenmGu32PVTDGSIlB/utYCpBdKeOz272BE8WmD39yMcC2kco0coHCPLHgVb45L/
5O4sZo/J8LX8LjRDWh2MK50TFZeEVob5gNrDVnrw4IzxcQVKuqs5t+HatBtrTuiAKGR9AevIsUNc
ZPoRgMRFZgMr43Uku8oOxfRw/kHjdn9oLKpDIf437BTmcI7uTspcxzRgLQM9KNNqmxp18ahY8OAo
+QkkJCQ8Jdv8ZtS084nKvH/tiqysOXePpgSVO5kwZmQ9tFn4kwD6C0SDVT+JVbFMPbT4+iBqQx39
ahIx1wwbsFSNfUwUYTCXIVVI+ipbOGCz7flFbGr2zPFaZ5yZkA+ycJ8KRyBKchNjQgB2/lvVTESU
3gnFS8cmmAvIy3+c9cgc2tQhtbEXvDo3xPKtkKkmArRmpj17U/ELvontnKvrk31ySoLN0bULVgAQ
5iJcfilYt2GmoTVClPKyVcOA05r9DXWNc3g5UclAl6VCajySIs2Z/BmSaFvv9iKiDl0z72HvtohI
peyhBr+uTZv4uNkeQI+4lZPD17Mih5PSIwwfTvsazJ9OSM9xyZBa8jV+WORFUn5zapC+iKmvZc6w
04XwRWBCCA8x1AcGD4Nz/atqnpCNvR/HzL/+d8JPr6OFr7pLyUwLd8EUQp8QAhqINkdHUbGAc7+5
XgiPsOoM8A/l4FK6C+FfSlzmmN6EX7KBGUnRGcx5n7j07WiBuyoKcXf852r1jv7VnGdK+Y/na2Fo
lT/9+Ayx9aC4vBfyBaaFDv60CY5T3/ddG7Lg8FIkm0BFnuvqkcgbf1xizCsngSg3HC5rluIYC8KF
f05sRTaL4TP1hQ55mrf+osN7PWBFGK2sOBraIsNk1q7F8t444jA4d2Wq8i6YpI+oX4HXZ7Regcl7
LWU0XCw+keChj43hT1WRvb5/N8s5QdabDS8C88i5ZsDhJlqHOJbb9Txhj+zkhtsjKMSiG8WOsDAQ
Ds4t9Iz2qpvqTIWxhmXmLgRXXs51EBsvmRgW5Ho+vnOMoRFQ6lZZCo+op3ydjdzLTZsAGnZA+euP
X6gxC7VxMvGwVj1n+LP7SnL0XCEUapegjDw9hXUa0tTtsMvVXZp6NUUDG67ZeS6RGIBwyjeP3efk
yguMcDXgnTwKCNZFsU7vgT+g/Q3r50RejvCyEweqoamLEV2HKcJwlk8ScvAuriXB6/IicINEtl40
NJsvBhEO6ex2yB/5hmRMUsRrqvfj/SUZfPO87SBvakmTTG+Svd/+LwqjgnHqOzVYqM8edFHz/CU7
DEE7X+2GLB1zuV87Olcqu1LeyiWoBmk4r0a8elexEfE1Hnj91VXNf/sN5rfuGHmI6JrHNhEzQuAI
WrxeDQjAyfhm0M+ODxA1au51XYVi23wO5rxyBBTTcrDTNU9bQzUPIB3txhXLzj2beHxwbn5pTERr
XTxBSHMiDnyCYgpqiO0zpWh1dUBksEDacFIuAcam2BZcyqXCHMnR3XzjYlkPjSb50KWLzcAvxB5F
ywhYZSDicKjbHE8NScGxVoyBqIYZ7YpasM7BO2VRgwYvlK3Mj7aTNvfkNVEQZuOHhnE/2nwdSGog
uJlztNdl2GqZePo5463MyFj85YNH0uGV71ZLoKyQkm3FAlTabho19VQso5fMCS5asDge7WxIvv4F
dyJrcTeuKfmCwK+X3Dpp8ON1PJEt8otcosx1lD+NedDi2V5p5GRo9IlrGLkRaCrIYSs5bJ/lDWE+
VEY5k6Eq56kB5C6NAmmjfJ4uZznQ3Xe4g6k1z1DVWS2TF5cPkghLizrntH5AksxQapjxV0CEg8xn
Zh1xq7a+j9YOwYBfwP1/aeYFzfZXQmJtXIom8gabjQ/3Ynf2En2DFuO6HM4ifP/IZxtvhVK+qtUK
k8qks5XN7gLyrXamiGouVxEtm7ncVwIMUe44ReWupXnOTGOz5KocZoZ4SYdWUX7to7V4L5/f+259
8/wzWp+DbmOd6DiYM84DKfkjyRH0A9AEqVbFGXYjnFJ7wQ9TGmsNmNTMAp5+EFllNQrhe86RanzI
wqCeZHUT8hMsMv/eWudg0dQXTO8cakOh1lAswxKtjUBjJE5BkDoT9WN+SnZApOZdz6LtlfGI6kHN
sHxchmuO/KmPNTKjkhXbpyShBd89l0gipqfXy2Nx1cmVsFPnJixoYHnq9dE2pnaxO80IUG+AYPmQ
gPV5jKnd+Vs6QAnDaEkdNqGRj9+9lSf3DKfStTtfcLW2r7B01MsjbqRiPrut4BWPIpzBYc5bKtNF
r7iZmA4ewdLIZfs/TliVV2dlYjiSE8u2OibscsyaYz58Lz08N7MRmECUgfVDww/FZTeoDb04Mact
dq9JsZfRq5oEG7+NnTA55hq3wmQRItLsKM0jXHPRRbcN09mUDUdv6c1DaG6Ce5OixVFIo3T5BT2C
HpEUhYb4xUysK3y8m5XJ4yX2DQmIhYZFvmbxHI0HQMUh8umQFxJSE3PWiap8lttlbV8fZTsxlxTC
grR5PepI89YMuPUqDxnYp/WrWbuNfFRxPf2ezlXT0JAP4NJV3lA9W0G5XMMVVsnX4Y+IU4PvhngL
Yty0oLlQuFyfdZmGHm/Pzxc7EtHhhlutCY8UN5ssL/oijOMyuhe1HZGwk0NvGkHaKQZw+HO5kmoj
s1e30rfhs5Hqstttz5MhjjhHA8lDzG/TD59LHhakl7gyU17lluoz3wyBYoi+EG7U+ZYTgtb0Kdgm
OB/82paVQ1R5AyHyOjy8GXLec6lkVO2fAfzxTWpUdlPnJHK8TUb3ug3au0m2KGvO5O+uLrBBN44+
dueoCsAeSwLCJrmYZ/N37E5ICGoCf8CpWAA1bDPyiQRS3FcKXSmmTDnxrMOCoeMlCOGXzk+OzFRE
/mhWH4shEuP8f5eSycGAIPfyP1rBW8Y+6sf0k1D0vtZjlEZmmhCme3x0EXVi36iai+JPYqIOm2zt
TZKnzodwIO5Bl68wypTG0dXIduN0o55ffnNFHbOmqzunmtTo84AHqr9/ww38oG1vXKC2Mw5z4LUL
Ukb8hmfaHOyYh3khVWhDwo9L7f5QGRwSdXqjeJj+oxp7Md2cUKUYUBACDsJWjP3X/Sp3bwqazWiG
vrT06IJEtl8KB2Hp/LmzOKvgLJxGke+oofTvIIK8DHdCk4i6uiCFYFoaskvn9AWKtqzwaKC21pL5
ote6C7jfeU3MChRUoFCLGAyFw7caYmrGTLnFU95qtoLZ7w8Vtx7gw21KGa0FIw0igI3L/KZyjVWP
5op61OSMV3SsC+pnJEm+Jy8GJSMcT/T4Km+y248RzzcEAYMCLVRKosH4kbg68c09s2Hm1/QrJYd1
rLE9nFxaw813+iy5/uTlMgDnU3Qz81fgoNI1AqcscejXyEClKVRpZ7t+NNmwnmwKNCB60dqCLFUQ
LsgTwyL/xE2r3ZmCYzZSqdXF9b8J81zGIDPBBZ3T6hPQWprITkfJ1XHPLCzSWYFJ3d3ZF/73+8G3
43TeLKM5OxTY6tgx17WX1C6blQ4A9uVgVd+ss3s61j5kjP9cF0PPsmylN+C+9KMzi2YQ1C2Jozw/
7ogDyRJFgy+uhMhzkmY9siZckglBpvS4OFbfcGXEe+0IXai/G6iCHrCEBOzSKpcOrW6UfrllLYbk
nWFZoowiE8+f8PXcbVnJW1pl3wjqag3TFcuG13A26jMmkDWqeWPNBxuZNIsn2itJIpl8XyFxKjmS
0ep0du64rDik1+zX6x1qsyszVjPdBdszabQvFA74vzNkE2PJ+VoW3wvRshZ0wN0ulaPtU39CBIeK
eWWoHvTTNE+G/cMg8j2jxgeOMR+8vxqyOxBCOuSI/dqiYuluu81lZCA49jixjlh0Ku1HVQ2ogFAa
aScNNrTcLhf7rwZsGtqAXBelGHANMXQODfPnNaA3kPLn3H81PF6BXgTWqBGA+7nh3NKIyfRO+Rwp
S7dyJp27JDVnVlmceARIZkHIAz9D7ae7NNSK6bCcULiPf6qvb29bX51Wg9ZtGKso5X/qC2jUaU5l
bmFZZmSiDGuXmsShrg5p0hIBunScaiZto+uUAC4o/MWMGPCQesqIAp09iMDzc0Fkpg0ZM5ex8LW7
joGokl8fuZKRALyO6wl0d5MmiXWvQSQv7P3oj6qcrfpCJ2rbr7K8Aa/R3Gdh4YjjHZcmzhjqNhGx
RwobI3eArWgXt99JPa+ZHwvMBLGThyuJSdEIaNg2nnInQAv96FLR6qPqaLZFiqxb8YKcGvVCIVMj
OMF++Kuj6aGsDoguzOA2KeMrjtJGjhX250FUsyk4zy6mRK1jJj4s28k4GugtWacwM+ozvhfPUMqP
180+6KkmDBbkbZ7sc/k3ZpWXmwIj1CRp7vSGciwyRhjk0F+jQiUxsCeqKICMNOSbjxG1ymNS074Y
GN7glA290OfZh9u7oY0p60Qp+0+bnesRMTk3gfbYXPt25A1WU4alRhNlLnpA7xktYDC3MBsNBBDi
MgRYHNEU3QXXjfEB6zanLmg34Kep+jSz7Y1ikxCyVuEoWXDxw4xqdykASusuJLAlTRUn1WNvfoJ2
UWN3p7oOUPxMRpLimxUV33/iNUxhcnWMm1qvxGQT9bzXaNmKv9uVNN/IJzz5vSsfonGtzw70DBiM
LqHdtEB4CqMogwxoNoH5Yxrs0+IIn7/94fIDo1mBl9OKx9Vl1/s5T2PnRHIPH9mTrjxpRPjEqWTA
dsZfV2BXrSqnAjFoTsLs4QtnJh7nQ/MHvTji/e82IbyBpm58qgLsuQwlGj9Tlg05Q4H0UcFXMrA2
naApkOtotEExTeMkWF1SVzhaW1YU1CjN5CnVI9RLijjIVaFnKnc8YO3dNKEx3QBB4+/fc9kusNgd
/Y3O0dAsHz7WRDYT7vTOrZbA7U58fEc6eguJRltjpV8wzgBBuL192HQX32JyYSR8qIcYMV5IGzJW
HWCDKrCtmk/wf78doiwWzuGgZLlTHmwN7kBPJ8q3wEkc4zQ9EM1o/VH6C7g1DAsWYY+PPZmUxo40
rTbdRgCO9OyCRl+PAsOpP350vSqfs1uXT86yXcWlg4karFlHVicLRsZwWMK9olRwuUBZEZlRKieD
AGcs+txe7asFTARHw564LgXU/3ztZw7sAQS/iljtDuUt9Yl7VdQyYT79Fp03Gpt94KUDEgqOtKvW
hIugMJzcNhLTeKJL4mBoKO58mXmxuwuE6HT/992fWgy6NKluYYAU6jOB6hIDOIHXVyMsYBfcB8wt
lKetUfWe6fLSogbVwpuRfFm1+1Hhm5C+3IXOf+UPjjQLTUaDVgSlBBVNEOYW1FVKDANffdIHOcyc
EwpNybX4yMk0UZjA2UwAgBd9DykPzyBbRvHPQIV4ONpLhR2COBPZdKKke258MB+fdmjN+yfaWOtc
zbMctPzS1wJ8Jomm1wgUqFcp+BBw0og224XESDAnr4A0X04iPA8XZIBxhkHUHKQABbMDL8852BaA
HlNXphnVCpa/Sbe8cD0Se2i1xrVXruUfZRtA6PFjS1AXeE7eoAHEMWcbVkdBQ2xWpt8ROLqag+LN
pWeb147fs0yrOCgwcJy7YnHWR3xbs/+KPGNAJOTCuTiB17RhLUgOyJJbn8PL6CYuyVvG0lGWLfMF
0EYuSosTuF2BK7ZqidvL45zfTJ7lFeN5Hao33G2wGsYcsvVJWEEvywzwC0GIpqTvLakqT2fY47sw
nyhKWPBa/LkxxHfE1rbgr4Uwcw9yoVfjPVnmN/jaUw4JUPtRXGNarSTqFZ1Au/ehFu/ajuwLxcMC
Z2JcIzoF9i2yzF/TwcTaz0kHf5G4XxVf36ICoBH3e+kGs1HW4BxMDhl6rvlJJjuHnqbyIHUEZ1/g
XZfBaxqx3ahuNv4b7ppBz69lJwYp0+mguuZ/I1/T1KTqEexvj9HQYZjnzkPWqxllzQeSKTEMdPSO
NoOS63OVjelt5hhaVIFBPs4qsdAP7UDcfKmSq76jcuoPQOwUBLiulaKcXlIFhfPfuifgRVagbNBl
Q5WMYPP9TRYY4olJRL6qWPf39Zgxu6OGx00G659PsJtls2m9QhR8NOaxS6kFsPQDFcM2j0oaIB6I
5fcTI9T/Veks5bmHQ0T7AYM1DpJ/2K7f66N3Er0gpP6CzQa1izeogcGr65ZNR/AeX+4kTmq+KlEE
Y8gbXctEpgvKsTjNatnoaUJF+w5yUZpZ40quCDMWgY8exh5kVUZyWM0rLmWSdMZul4bUozVzT9JY
s1FEGNOtG5mRUQv14TlPz8oPseISguMvhmvUyxOQE+ETX1uZSITF/hQQJoOScEeQYXLdZAkhRrAA
qmoNGHCdP/tJWNyIn2uxfVZsGK6DidaHxMl9kzIQxSHrvogTr+pDFaTgxTjtT73d1UpAr3xdHDQV
YRJWjgoxW3H4KUs4XApUEBcRd7exqLKB7MmfWNtJdK9GZnPsgdMQlqiV+/kqo9pS9+UG4C4DQ5i0
S0AOlRq6kpvlmfErjNO2mBm8dpjMfX9um7CNqd5VQg95NZjuI7kTMozsv3LcaDXFnSPL3DXYYdTa
YfQTqpQuwHoRiJTqHowx9X4Hsz7sghpJWf9SZPYsP9RBNfCEkgyKo9ELWpR8fm4+crnoOWkAyFGQ
B8DYr9/kldSp7kzwgdwrIeutpeDhi42lKikvyyztB7ZjZ5UKbuPtMbONieI7xKhhhyyubrmpJpz5
OeB0lrcTAlM4zNbZ+lMIn1+FTAXOyxn9Ow3uA2aHX0q8XgQGEobAz28kxMIbiIVZTDo9fHkH4G7T
Q6YAgRpfsbvulhvK7Id79jilBgszmZ59oth2znhaduUHxIpNU5uB1cMJikU3MSl+7yKrtyRx3ABi
u6Z2W1o599kVFNIk23GOhG65TPit63KgP0Ksas3hcyr4Rh5Pq78Yrn7y3922EmqpJ7dng+dbD2Ix
710J5piO8np9AETf9bPN3zdh5Mqo5TarlU1ZF925Eks/CwE61xYDfTAc8NCyFS2z5yUJI8yjX+vA
9vL3h+PCe1HPN3uKIKq92/TrP5sViyhIeS4Y7ky6jR5Y1VQFtebdMPuDDTHEbRkfWCfS6XPqkqHC
L2D/Qqrc9HL65ofQ2IhSPcbyKxoQMlZd2ySaN+a8unV0o3zIhyWi/RlAwdQbmuOef6eKNupFk41d
wcDmiNsL0d9D2qu+YHDewbo7myX8WayB0UrtdunkflpsJgasAqJWUBwBQbjGTMV9PpfoQFCD/K5s
idkAW5OuJDSh4K8H/wwJthKISt1NNzQCWIGQo93i60HotJm0SxYeUPoZSpeLO00b1cV8u5XwBhmV
z6HB4iS0m95y4eOLqFj9KhT4zvtvauOElVXGj/p8Iq593hRLrTsrRlCJtahz4xSkfQ3jjWZqrCpr
I06NLPueaej0m/Q4Jq9aztS/62rBWqUIw2QMXaZKAQCDu9FXIcLIhOzhvD9ucF96CImHd6Fr4dCg
fzz29h/0IqbEX5kzEUoh6bV0SuPoXg340eTqu5E09Q+1ZqGiNWwfJGCtAUsGtIlWxQJj9XR19kgG
QGW6XQFP5vdPZzUW/GBsRoHz2smP9jRy7RLnp7Jx2Mj+uCfYL83IQUKCpZSR1iWsV4FJIlhdAdJV
AYx/pZ5RWOy74na6dbBZt4b0dnkX1b4i1yHM8vaUyTK9bbMhxiOv9I4UWlr+xP8pgkvFxeqSabEO
AJvu7MJITQKv7/VwtRbevKkW8P3VAYVqGiHRDBiIxE381/IjTJXcl2SQgiKXYYkbkboWPVhJ81sN
w8r4O2J9lCc4be+FCUy3ikhRFN6aljmOJQKl5r/OA7Sd+LB0ZTF2WZyS5YBgwOYlx3inXvzPvinM
LRXXI9b/tftY2kWyJglPV97kVPLYTJOv2D2c7J3njOZhEl9tfByluATYAX2eg+x+g258ZD0ID+eR
CaRFSIKRKMQx9lKFbMP55EMvOY5Rw3er1wlMCl/YubiMv/A/PWoGjInbwZGYfhgj58lZ4chzpro8
NPc8pf/SEGKZc7Z7I7Ljsyg7IDDQzyCXnjhoOJh2Sk421ahrqosVXDcfWP1pdC9z4fFUgkX8Lqm2
7CSy6iSqKVpugyu4xsJAgWDYWiqv/Z4aTgLWd1Bx58TCCD46+jLNTrIi+JVr7YolJ/5FOp3HsQR6
WNOrJpmUvp7XGiahvtyC4c167N1GJAcaB/bg39gXDXnAEF4dqedfnS+r2qpu7XH0cSOzV8V940J/
y9gqepgx0PWmcyUNXGY2jeyIn2zq2VNvnv3Fg/ftZf1LlhXZ75LxnDRE+vE72UPfpSdf8HZVr9/O
+MyZyo/lO4ahIhzOMThkDZdJWVIEI3vxZ5e6gUlpj9K/0umZZpTiKbi0+Npi2kqIVCQ5K9xwhAlE
3PhDTSfkPDMigBuOq1cs2jCTF6Ml4GPkQXwRbJeWwRaEkzo+KeS8zg4r1zh8BUBF9oyLPvwKtAOM
1EYfIbzfBMIZ3NE3OWrbjJY5q1bmasYhPdRk9BVjFj5x/Iag2ebjufaYfBBoWau9NFxOGsnBxnLY
N4+DjDe3sPRkXr02qZTplVLaxQvuuyHw0peYhO4E2npoleWvVo8MKTkw6HbGoBv0Y5Jv3yGCI3ad
iy05NELTHcS5i9eZYQpV2F2+zI/ieM9qeltbBVndIri2X7HsXTdU84rC7aoSXRCLt4+m9nx1eRBM
+AGFWICKDCJb1uFuLex9NZWJUc6LT3+C8gAoB7WCrF+gF91qWaegLbkUrx/dsSdgC2z5oVYpuhjk
1Aggt2u0lOAPR+mFlbJM0dzDgBFgsItjwXd5zWkviyjbFJk5+MG/mvVNj5p/35vRMkeg3PucPnk5
1f6f1FhcEkcHLpQrMYY3vkf57mUNuYCt91HtuLIWct1TqGgobhrzCzTcnyeGF1eOFLzF7upPeErC
7VmUA3tcP/Ki4p4tt5A1cvbBDw7v/1OOVZBkdSUFkv8Kkebn7y8Ni1OW1ilbnWShcdtsZGqPLOwR
BwqQsdulTNwv215ig+SiVz6aq2vJhoKuGOPCMmYZMMysADOFJ6+NLPKevtpkQ4mYmz424dKOciuh
lggs0P/XF6Yt5+HTVAfFdUiy5vxcK1UsIFXkq5T/Mmsdo/qERUTGQwJ/YdW0DlkN1+JEyc7QURJf
LO0H+FgcxQgJqI6uvpOul51rrRDsjo4IRAdscVfkgdTer0QKAfld2X2/F/6p+xuam37j/6Zx9qOd
5KeVOo0H6tuiHJQ/e3JPWzJyqL+/XLsOJPaAi1Wix5/6Zq+wjOYRP9ARK6rqRDQewLUFSAQySYKf
OPDPNO59C7I0P8B1R9CxbPwBJsITpeLEkc41IIr5njoYNGjuGL4o4LvqvYesFjE8FpPRocrJfSh9
1q82/z8tgswcnuhU+1sMvCNCdP4ibByJPm+XevmlbA55ST9OdL3QBDHjtd1ZPKIye5U2tVSnsTXk
g7BZWKjdRsBAh6uWhtS99YiIgdSs1s0nUtmd98QtCoTpfztC3NBsrMkvw4aqRAPfad1anNa6EG4p
tjh9VRg3P+p6IBQzlZhwVsphJyKCM2cWyyIpCKAj4P7d52enrGOSWzp2F5YBKEIuBvs8t5GBEZ3Z
ReNED812RmsgVSuRK5IJCZMYdgNU67sG7ju1m+4zpMieFpqtpEzsd0QFMZoEjmJe+ZJVMXzRjiib
A78tpcDN1mstivMO1mQNKuoJsSVGYRirhibWsBpUoF5zKtFwT8bVLLkPWcMOOq08C4JfE3CAYbJn
VYErqYr8nyiyMyqD8AXuXIFrI59rKs/F2Kvj4IsJxizlTiZwij46+WBTGqwFjyVxHNz3/tGMR6eO
emrkWcNrsjtCMXbkeaFhNROTPhH/nI3RlV3pp6FKEa6QzqJMrQFScQ69BCiLcVATeWlUU+dxG2zF
l/SXrJQM+cHP6cZbfgxPamnWWrJjgbL8W+SVNO83UtwkJhnBUHzM+9bMu+9WviiJNjkzR5sqG+c/
SdnSj199UDmhZ5yC3tFLdJ9Kz/C0s7YEPSfzyTBIa0X3KE1JPS8GZ4p3siZ+QBHymLidG+fYOFn7
x9XgRFYaKUpU1rDxVGDUI7ELf6hmqi+7YbBELVnWVQYwrHtcKqW87KrV1ne/4okDbLbo/OGCeSYz
crQICidQlhjmwAx3mebFJlc14bygojGVYpmOOzhMc8QiF9UMrYpPnDYvLtZNbzT9OxA6O1w8e9YP
7KpERUefvxMj1A625MgCSePw/Z6uqL+EjorB4tBOmCN4ZlnXXnnc1EYJSEzMWBJc4vjy/lCoMIIx
CZp0Y+fkgVEZrGmQzVxcrsaqnrNN5zlH6wqjawbDCEHBzYFWvEMO0WUTxMS6Rg4B3BTg9KL8pabF
E1AUzW4rxWB9r/GFPi4SC8yBy7U3/PNy+uIPCGJkRguwG9Z5hc2kIBMoG0bLG7fPD9qFyWlJdvhw
YN4ubw23Wy+EJGbGFesxRMxZoYHR0Eb2J7nAUgwOh+U+8sSpWPa4cd2RdejtMg7zOC1RNKAnwYmF
BBN8eDkE07f7PIJIcwlkJwLjMPbOT1ifKI66ID1mm9hkm3fuheeD8hQX/mpEr8Z9Y7qiR4hspMLK
xlHTtTA2955qgivpr/PjL9SX5JttN274Fwg1nMHgK+jrNQHctBIC4ub96C+LZ7oOMmtGtHc2/bkZ
yd69H4cODexHgEM0HIaSATYMl08Idgfw0Id+7IIu340tD0KsheSwBQtWa0K9rmGrPWnaieB3tM6k
mqoaDibBEhOEzNfVDd8uQRAb44EwEN5E4qiyw9lqxaBfe759V3DqwocV0aU7PzJYFW1WMzKry4ey
o/mREd7xG/E18ZvJUZS4dYM4C5UFa+a97S5CHAM9nEYpRX3QJwPS5QA7Lromvc6z4DvR8D3jU6Qe
yr0kLQ/Ch0zZKjFJLv1fac+LlR2Ky8W+18Ldue9U6OUH6HdYy/4Sokf3efHPh51TrzHCvtIpkTQW
/B50ufwUf5WVfFrf8KhWOyTDwy8lCf6OXOIDY0yXAYakBuGY0I/5XgZKyW4r9LNKkCUvI4HHRjlE
2Q9F4DsoIogUd7Y4xWvOdBSoPALtQJ0VKT4uIHZksO631322zYTJhdW5tlLr8+0plGOJwHnlmWQY
2OvxjF4mvUaKTcYXIa04k2dG2GphAPurQx2i1Xhml80Kcnj7+v5+yIWJ7XBzCiJTgB5MJp9ql3Fc
ZQTVeFvxrsFVScCAErTq6VMbYBIQ9qs1blhIjYugYdRPWYuhXDk5PfuoD1ZPj0dEDBp114veuGnt
661bPFasBkFqnwcZpNhCcC0MqExPT3yVEoQsmEig2bADOEHHyEmqvnih80mjt+stCqWoRwHiuRv0
m/DG2zrWbrJ75fFr6TY1ulmSiNyy90V+lxlzL2ecl8jeBWIWxYDZT/kgOY0WILoc7M/z9QrtI+78
209PXJLgOanieaOP5Tl/9gITJ1Sp1QbIDuUNRmjIQMR9/DkB2KU4qtSYLhzWACTkUi2XYVrF708h
MhzSpTjbLYO1aiIBXocoB0oUHIX8fJrdtQvDc4qRoCChkdY8WnJORiRk+pK6oJGbPMbAp7eup3+B
pDXfQCKzyAskgmw7jOwfjCjF2+qXBjt4vRhXps3ABrj4Oh2ozPVx9NquvsFM2Pk052JnBW+pNwxe
wpHYj/5DncJ3Q10vbhPWRc9pQkf+sRKckyrqWffHaAycKdLhfob/I0pPbMCuZB24Kot1Z2F8XOYj
PmiRbyVajLq9acvEZxS9JR01e48p0x8MeEXO0BO0hcp2s2+aL/U+U2lah5oXGVyRwTycA1v5QFvv
Km9IA5tROUULJdXoZXL8/8w6GRme++4ceI8iKtbmo3wI8xefVNcpBWlQSwGbva4XHjS1tDbV8ZUg
KpLsmUmRi+udpP5TghhujpXnwJuE0mvol6dXBcy2j3Z/k667pM0b/X87I9Bp8u6c6TOAk8KUtZ4R
xzLGV3pcYs5epBs6DySpauKBJyFfOhApYiUegY5ftCjiUkEoLCqSXPvjWqsEbsc1aK4q9346Zc6z
odPC+mJtuBMIaTZ51ybdOcGE4NniYU35zBS/7MO+O9VRkEZo3iOuqOHdSLUunFkRml1O2qDi0nhB
bfsP4w6XNobo2lFBPPTD7+dLXPbn8Q6BLaS+jYwg0bV4ZWoU/HBQIsvkkhrnYjRndMhQDCzgFbu0
pyqUo0O9xkXuhWBOU5UAQcpIORsICsxF+pca2QS58ovI7IHRj/nKg5tIA/yfOiai/DEZjD2K8wEQ
exYfAT4ZW2bEs2iVuheml560PBp5Fq+CP+U27q796WUQ9a1ZgEhPI53DXaIJ/An7NEK5eNz9g4Tn
xrPmX/sb+ziGdMjoILNjjZs9xtTU8ZBkExr2qUOI7w8rNpRM7y4DXrnG/3oprrNK6Z3Fc9RcorCh
0yZKpT3x7O52lO4tYe3yFeXa1owqbs3nCWYA5B7LSxBy2JBvyShh+Z9eXG91iq2KtNT8GzA9u17r
0FP51s3iFa9Iw+WsNBhstjp+JOPd4z2HwTNrnKCJdVkXM93x+MkU6WMNnF4T1EjULLufKe7Xq2Wt
DM3poRO7TFgCg5KKaQPRbG7llLRmzUyOhRj9dy9k/cjAYXtup7wfvnvUVFSW+anXJtKGbtyEpfJo
Dossl+zY0ORxTVP0vcO79kjWiXVhOsam0aaOxhn3aIB/e4V5rPxkY30DLDyZqGV1LMiBpEUqC+qe
xSpx5BPzm21xjpQfWNZ6gqtRWqM8Db+KViUrjGOV2gUlrPLV+uMBZCxdee4xtuKLsImglZsNF71e
JDfLHrGUiidJ0uL8dTFJanc432OTRZdy/7l1s6oBr/bBHj4SKO6YPwMwqdodOzD7mumqq0s/OF6l
EgR5WwxfBOiJhmSptFy4ewOqdSRvPe8iiWXBIGzS641mT0tfaVn1t76dAkdOrkQd/39w/GFroguk
tJ3Q+GQwIRXN2E51iqft5lf4xnxCsgA6lzlEX73mk3NGYjCzXeBDhfyCfD4jz1yGCTmtHSpRAT56
b9X/bueWXOU+9QjI05FPF/UxgVP+vBODhiaBtBnsowMirFWtHn6sZrE+uVjc6LaBJpxDzWVTKWaE
N7z4DTiLs0j3b2pEWDjFDiTLWcAVRVNgfna9vDEB6RtNXlvfucxUSSQj1Si9NrL04jWgFvymfAJG
wP9hYf88I1Vt0Mh/mQ90g2ffbz7xpbxsW1RQcMWFJop+mLf2MJbCBOIzQbmXr/d5lvRtrQDn0R6B
9bq1n0khOtC28cgjMw1nWJg7Lp9UrL89tGzK6HVJeU4UzYb0Q98RVvGKldNOnr8Kc8O/+0fUQ0MP
2ElBcLN7M21LTz48ST2JxZYQKP2PUtTw3CScxXwgwOy5f/29Td04GLKB/Y9/9xtQXSf2DEkawka/
eCoKwRO7sQZFnaPCeYeQgxVY2+rZdwkTDfYSPTOQ1WF1u+5JYsV1NXpg8uS1bpnX587qylOh2AJL
nLnpZ5tGi4NCpYZ/VRO3tgggXrK8hwvA9HNqT4EbbnO6V9j7Vp4NdOOVPeZAH8JOQmOZMPNwa3AV
fTkImiMs5qo1FnTacZSnraDKhk2Q/vhh7ZyERUpVvgVceMOctVJDiA+IPUFQiKpeFTzUjHPo+SFZ
Sj+9uIEE/jD8UU9KJNx6ff6JnxW2XziitPwoTS3yms4kYTMe//NmTPgNo3HV0bVG5KKtrkIBmvdv
ae5P3kOAzVIshDHMi8OsCRVhE0v5/xUuQrYGA09OUzFtKLH5FhFwwVdMKUqC2KTYugHHqJEcCvHu
H9A0sL9U/BBlDF/GYqDzHfaMBvO1qj/QWP+opZ4X9nfZ3l+zR2LtSbqZ0vCIsQDtiwXQKYKKXGXc
4NwX6fOujaJw/ORIoNUcxy1XA7yE6TcKMhQkw62Wyo7f2c30jwS7qQyP7bIHaAy4HFvn70wdhNRY
xjQ4EotcQwuuR0oGLh/++huxLWa1goxMQ1DEZ1+riUVmYneqat2xQEbDZ3/n2Al7QWZdVWZmAdDA
pw1dQkfTBAUfi4Dgm1NRT0yAkrK4Gay7iZRADyhew/SrDribYfTABNPrqCeYMYE4F8OJedOPbxdd
53DOSHWGF03NmQuQCdHrBcvVuX4yM+1/iLPdVAtXWO+GShKcoJUf6S/cBNvR5ZuJ8mtyeGA3ghDb
IfF4AG+ZNF6WIkAfqhQuSAdEALoOdxiSziq2Slj9Bc7Au2fCTHpWhCSOKMVvLG6SDWW47+y4trey
RFcGHaKHbVcuRu2NozfT2d9yE96kmEvYE3uc827pXO2G7u+JqAGNHKhJP9g7l4qE2QZsMxroLpe9
foNj/NOC9Dsju0Hx0aQWUqt5J8lTP5gJ722oW7vqmjjcbMZrydJR/cNNwU+SXp/pjuofsDoiMi7i
VkSiZuN7TDJx7g9zPTq3KhITC/+X+gpAKEtkLacAAVDP/qqfj+266uAKePBGJyNNOe0lGJRbv/+y
hYYE+JUga3kaNQdzjE7T9iYfuIatHX9+kkTei+H8USPaoehmjcoIKNyyutCVdO5LU0JTOIaAN1HY
zHQRLnxsq6JXbryqUyjinB+mNSfvHLUQ89AsCFUVTH+PNABAeGjLh3wPcdHMOSm9qW8jpwKEV/fD
bNZSO8Ydl2/nNk2cdSqazntMuyXHNlLmvu+qq4eTEWu1qpycLOPYjsiaASmvUR6RvVAn2jfMI5ed
7/8nUR4Ec7TduUuplrSGCbYoAv9JBsALLndCUoReerfDC6pQvZL3V4mAjIMxCnA+l7xvUMLqIzV+
0dc1EIv2QCPSYsjxfApyua7vxaM8lRGCziJUGSdYg+yHSV2EfnwraOGECH3mesNUk/8qpULMpVwt
pCNtHKNJUkLuSU5nb346lkLC9C8Svp68jpbamXe77ygwS5WLDUjXzpD9VY/SDx5kDAPOdq+X455d
0Mmi0EhwNSbz4sp2WRj4lRlFQP7gG8TJAOAOhwX7KMlxusCckXhXmQdbwnTJxITt66zfLIMoNJ6N
/94KyhTNyKUxfjGMBkEEDvog4FybkY/vXQ169sglKTFItIJ4vCtZbOMUrejS5kkGL1bBG0kPnGCQ
Yiaglhi5UfLMszAl0hJd7B/4RYjuNXh6ob5PVJ+Br/QzteCmPytUFozuA0HYNT4sLQJt05dn2uqz
KlkxNhuRKIR9qcrFPV3o1PKCS0Rz5Ryuku1Y7ekqKz2R3/u27URFyojY55+3Wd2RDjSEGeG/5vHa
Zn2mxVii+RIJecOTSG4MxTJkKmmUb+5jcwzhq+uyhjBtXHtyxzq9l7uSKOOaUbvd4wh5iV59HWhF
oyyWNFZbVekChO7B4gsDh1x4qBdXQrmQ/ttaGzemDTh9MrNXZDZpZgr4s+NUIkuF8y0lVhzCZcar
klN0PKiqJB7Y+jnqSW0kM6zh2RzAjB9lsNaIjKJXL+/6i/ehBXSihd1Qz4XPKOuEuQ8HN/SkpRSa
DTDweUsIV7a4YSdy69T9oLhZH+m55oapoEoTRCddG9NO9N6aJbgAtltd09qbQvV/KBbrWMuHpIJT
XnhZJMslMt9Ovq8pIfjRoGehDVtvzubdIuLyMTsvBb0m+C1Ss/9MbAgx084qWE/ts6niwYdvtNyJ
3++t7FS/6OsY5yNpVV9fSWGShr6yx1onfwGE28Ew/T19zmMrKkAyGSTgue1Wl3aGoKuBiB9vRSL7
o9Es9bFsJblcKR0CEXQfPyHe9jq6F1NdmJx3UWfae48LFRhcn9iuKf8bwK3TqVsLfM01dv1ZUeu1
qAJfOI5tmFB1q1m1xBBsiPeKsf7OBWyzwmMnF1UnOo1w9fpi5jWae0NiCUwJJg66fT3xqUzXnuI+
1zwQblJDKzYh+B7d56dxQcgS+L9vrdxcOxMhRHS3BSURx/VmDnR+1o8rxztII/yBZui6tASlV7oY
YMAnRTQs4jwMXp2zCW/cc+E10NZalmPt8JKPuttU9aPMZS2JrvJvd+3NX1vJkqXjkoFDcY/b35b8
CR7FeRXO31XBaXJO892ziCXZJSMnYPGiUX2obhZsXH7yOUDemBHchPmqL29tO+8ug96mFIanSua3
RN+B/Ei0h4sLJ9//CqFDU1S8MkWafOlINHRVJSEhDnUMbOxOcJ0vB1UcOV8OkgOuoATocHnsvZGA
IchFQTUXqOByeaTmR+zmIgJrf5iUwVQp9qc4NxSJO8QrCkt3Z2vP+xIyB/DsDj5UZi6uLO45kXNz
UunirWsKCdLTo/u9iaUGVRG/Kp8cMQlBQiP5sT7ZRuAN3mG5rtTxZ3u3AKfADmOKbaXtfuVkatkc
EGLG1v74PFaFahXHXFQPeu6UW8cOibwtdAkonYwg51OdDKSnF1B6IldCaL3wVY4N0gwRkpQqZJYe
k8dkgOENpkfZ5D4ZPRKV4PHXN3ChDsMx4ji3tWSeDYHnvi0BbMpUK+259zzDzmelUS+MLPsnKrax
Q6LDO5ZfHgPKy7smIlAP6qDDwUwtSpRPrgDobODnQjimFwzK1shq7UwuDnKeyKGmjNFEqSiAAeAQ
GLL0HOBVr40TlNUrdYxG+PVGfZVuRh/RIxq66QyXzdBhIG8vl86HEB0Aabw6hJKjJv1Xw0KdlvLR
WEeg+BJLIDHZ2ZzftertOjIovmYOlLfTxRcURt75082d5cjYh8ZatuDHyrZJF9SqhRwFNiVymtSk
GZgqRe+2bgptrzLpbdM6lxQUR3fj4UWofTolgEUkGMva1CexrYeBfLKP3g/S15xb+7LfnfS7UPJO
swq1/SPFDgRfyiCQo6yBwyuBXSW4v9rIxY2McvRuDp7XPw24NKnkRSqddeinDQ4AdlSJqnLytN7U
jsT6YOlY28ffOaHnp68/2JkprAItmZCUwB5rvURtWQilsfl7GktEIbwkNwtsX+KBW9cp190N0emp
GB9D6EeH6Whjl0BbqLQJ311pywNgCKhKntZv3vn65u+sIzrMza9QxHaxaNUxnXx9RD49JfF3Yvnz
JXHoGyETkSXclSVBR54ZYA7kTGGpQbMM2ehIbP927LCO4Itfeoi+ZQm/T6fe8Q4JhdWtE+CvKugv
GkyglMrRARmJTWKTy85jWFg6HUqXAkUrN9ZB2AUKuai1Zk3f1JhH0bRDifz3IZAQZlSCVtvpuddE
m5QtF36TirtlrhCc55ngQtiPhpNoNmeASUyTljDruKp1/U/hlizTqqa4mnmwb97PXkjZuJhY7ClB
m4uPUEV8zabH4FRcRIuQfQvJ2d3Xr+UfqgkyrWa7YT9/Fy7StCaHNGyUHjaGGy1cgEM/ZjgwQ2IN
y++F706lvPI/n+qvqmuWDnlKFVm+6y6bFhp2YoiUkYHQYjrzVybtqUFNSNikelQqJ5IeLJFs0zi7
qPhUNNxZaQeLzWndH2M19eNTDhnIRgph1Xnwvc3bRk3+RRlcIoRoLRK4NdIIkvNWGdqCaerwrVVO
e4Yb3/27oYVvjqEmVO9dQE0+7N2G61xDop1aUlX8vQd8Rkv8mLw2j4cqVuKadkg4Yfz2sh6JSIN7
2alCnGJn3+kh78jc7FFsgmO4WDp7uqIkZDE4AEhOwbQL2MVcev/eQhSsGbwAU85/SmnoD2JvFZoe
eBeuIqnJDyG+xv8PRZug/opok9wjz/3Mw1vqcRtDz9JVgKVYHWZPI2+0CO0AJ0gIxtK+7pzWwzq1
8t+yXSbjDMiUG0QYxgF0xt9s4dIr/17nmz5bt9CMw7iWdQ7gtDoj6twZ+c4QYtQhmkxVNPoNGd6G
74nk23xzxiuW1vd5n60lrkHGDPhkKDGUE3iQ3EUQfU/4QerIDytdbVxrfKo5K0qMEu/hCwOKcYyX
UsYRa9UdWPLQddTYZMTQIGLkXzupB8+EvWLUnEeAHo6ezNITpyID7pyPp3AEBjBHijV9y+cBbGVq
ml1r0oBmZWiYbrQ3K5yWiXmOTu87RDmvaaNXKD5RavUirFBYRU3KtksHEwOgxqR9oxWTt61Civny
hwe5QO6ES9CiDLmjrX7LkhQuEfRSF62Yp9IFPkU+QUWT3agGa1wwVuOmYWHqyz2qbepg25OCfW/e
BNQZYvxMGYqcNFNiMJDUQiBa0M82w4PqS6GPkopm+eFNsBOuwRFo7qwt2vBsukGBcsOhm1aq0CLt
Er8Zpcs06CRWjsFVEo8AtpLTfpfef38xfMzDwWOuU5ySh9mTir8ZHjIppu7lqa4+ihT/k5/iNTuw
VSOIirbGN0n2zGncKPQOLNTg6N1oYmMKwZLTLgc3UG3Pksb9i9+DtWxXPejILt1H9mYj++uxAqly
RsyOUQbg7fuMPbofgPWdIHiH70TN87+GhzEkRF4t9wzRiYVGsfLh6Bmter1C6LrCF0sLlh1HuzK+
K8FdddXu9pmm0saf7GAs6C9Xo66ihmlsCHrDQEZmR2hLFtJBIzF7o1cIev3julqk1h5/XmgL5b7u
Lns+CnxsXG/o9P5wEJ76uMAV+ainlH4iWGcKidScmpkrq1HewVO8LOlTmbSro8IwaPzSoTrVz+b5
XTTpEWt2U6TsY3s2i0cXX0inN7U0Yy1nPy0MtlB9y0qYSIuKItiqzKI5rkLJfy8T6i3ITRpyBF8n
jDlj40LGm0KgkvOEpQZk+LaZN0024Uc5OQej3pphK6XCHWIEdIUI9ELYV7o1a5b8lbFLrMFmFCPt
43cy8duG5UNJVL9TU9vUFmEx4XZ2rEW776fdchditJyLSS9mqDfZHcCpDQXF2B/Z+fQTP6mswJOl
uPBDrJyuyPgDe1lvNkg6LWRjD0h11jXBV6gLPyP9ITZJ8SGW3BjJV7a2zbpOp9od+aQeF+KIIKhw
MWhDcoMf/8YfQ9k7koNgCAPfOzqTdoN9czrCzPgCgX26Bb5EBkSwhx//TY5pZFwWnaYY95ZYs9d4
Ii3OczDFToFToqa7MLeNhlpm30pLVjteUIMEzo92zbUm+p7r2zFUqDnZYnFg77iq6FwfJZnzx5Vp
lOARUnsmPYIvXwWfEnlgscTVX6lKfzdN1WKf2VKUL/rPQI+OWBF9FkRUkJ278QEvGaowdOM+R922
jVdjsq6WrV3eZ9fBGK42E5NDkX4QYYr1MfafOjWpos2ylvtQrrwIGzh0w97g9uGfIekVtzQK/GKX
tJKPxg9rm9FSlFstmMjgxpDs4AIYuz5v9GIaGPsN70fpaGOjr32op9ihmnIY7PgvZg5w7jJJZZab
kJWrFsz2+fGHL652nqTJkVRHs2x8e16LMIImmM7puRcml7+9A86gghhLSm4VE9aFWMwDTqwBQBC/
yhb+iJFJXiKj0udnTSa95pFAShPaoRsQupiW0UTuuhcjqOHuAZ7JpdVV/CpNTbOdN4IlPwZYvmej
dQBoL4638tMP9CB4F8d1QlhabWHS8XhIOlUwF8rz+QEqyFTVUA6zu1SOcrN1oYwzHjgy/z0nRqhg
u8qG30+NJHNlFBeWr0bn8XoPvUbvpMCu46FLeTtB9lAT71VsRljtyGJky9FEXE0+wZRNeyd8Muuw
jFQfRmYBRX504xlUn1dT4XPM1v8ipQL8wqdx3DDGHeVZNZJC1Wr/AmpYCocRbvM6fzNp1vpkuoWt
lM45ANzCp6zTpwMvku+EP2gBfTaaH2bsLWgCGGu5ZWdEyDzyeQNzV5winiHEB/Ucm+Z7nE1P/bac
27X+LIehSbFIBGPHzzWgrei60deDpOL8voPMvEDrDNI+pBHLY+T/bNPJs2W7WINun9PI1AwTvFCF
DgV26Kx71J1TwmCPYf2ubHqI/5wrL6sy3hnuXnCY4UwgOI01EB/5y6Xr71qHKxQ6gCyYJSxi04QC
oiqLJ/ME2gBSoHG0i2x3Oa2L4eF0TlOBzl0Sg3aulOiFOsMpGixcN9XyGwqqZRF2x/bMbYemXp5t
VNRK6J5RmXrMZ9FpZJT9sqW9ccv53zG+7c+yfLAqYp0cb72DA5XBnabYob9Vl04fswXS+NbS2iv5
775FRfAr/ly4tARtYLXCVolQ6twEDCqvL+k66yrEZktn/6DaFITUoWOmu7CH7WWFPC6CLHu1fJOI
uKib2P4Z6zJUCfz3XA6BWfiy6d7Q6vrxlgAjTiIVLdO/LKbVC3NFW3A383qSc6JsDKNwMABeA7qD
810Ik0Gy6bRlXLzPRrBjkHA+3ICyVQbw62V8/ehhJdhmoE5m2ELEBeLDkvUHO/RHwhkCY5xTLsuI
nxvBZy/NcmO8hgDcUa8WaEzsgufoACDW4HtozH3OXFTCygklkDkeZ2VHFaamyV3mnZQBMK4Pj2SD
QP7tZgcHMct9GVIMuyZvav+XAkF2mmTwgIEhfrP3sUXRxcUpETxxesGCgvGSYCopN6ROtXb5Pc/3
ZxJ+xYnFTyCbZmDYPLCzOvVwsuPqKpn/r/dR8pf5q9OOhpuZDUeWlrZeb57ueIc0WqW9rITL9LSf
viqn3B+Pqyv2cRfiYTkq3ZwA5Y3Yt7uCW6RK8Yl54F9W54QN+yzJZk/fJr/eUmGe3W0qWMECJ7Tg
ak72c5aJR/K+XuSkcwvG90wihkvQPo5GLrpfqnP3dDt8Zr99kDA/pPkzuqerD8Nam0exp566NIAI
knFt53ru0ipYAoJ619BP870WwsRUnUBv8hOVfVWuNth/phCAtTv0xT12+JRc2cGmS/hZ1W7fpx7L
vSnzoG3LU5N3Bi0+BkgR2aLZJ6pTpAv6kcTWpoOeELIOfa8GvDSmtcz64L++mEibqFRuWRukOnSK
u5FbALM0s3wkVgsFJW5qdswVVrq+87iQCZXGfNPzTi2lxvV8UxBNZW50Lz8lh0AsdQrDAyxcQKUW
AbJBcKJwT5sXpawLDhEn52ZfUUzHdBghMxlmP1WGTZVK42AefEw+WhohQtOq3chae6Ztar99eLnU
yOnq5OmjeAIHgpJlBml19nf2WqSEHnaWZUJVnOZ3nTl4Hl6oBhpL15H5+tWgvTryJZZt8Jh5Kr4N
qQG4Bg43l1S2Fm7L9Y/YfYFG+k269B1nD+OlmGY36ydn2Pto5g+7KA3u8aushlSHbVjgXaXg21Cy
5wyiFlu27rQQwTwZWioBdvEUmGVlwmIjCgzIvr/40GXtwjJLTGgqIXlSnUJ0T6WFpB2Kus9bLpDx
f1bQfuguUQxN/KeRQHvuW6chEUwIzhKJMuGVxsERiauZ9Xdi1mYhGbneKGrUchksy9fer0mQRbzp
4VjgOn6ZG5bqoyM6hWReufGdSYoH5CwT2xWGQC+7iCCyQsfUoxfpOvnOFsV9wn68NLUlQnlX27pN
A467g8UajEARHDfbBwblC4LsL5KwaOZaQGzuOG5LnZtL1+eHnWAb452zRqV5VXLieZxEkszpCupV
p73qO8YJclcKdUmZa1kW7CtMFxQ0Qz5gPDhPaCE3H2Js0k3ThnZzowEHNZylybKzJxSXQnw+OsCC
2mjPmCpBWs8G3RWYsYNfPanC2VxQNkiWJp531Fc/0MvRz+dZEnIGMMNrnU/h1ANj3bkvpFTMXHny
PJ/R5N5cUTVulQ9GxzL9VBKHu3Po2AgtQya23YujQlSSFwkZ+c92UHvECiSu49Y6YC9yBoiBwqou
tGW41IXdFsoBjBoOlq6lWuDaWnzudLlOdLaG0D7n3dGeV03tl/YrKjLEbNjpQ3OOFYgErMB4MGfF
pGqPhr3tQ1DP7a9FL4Dcse7I1T8SWwhjv4+icnA6hUo+6vKP9lYjCkhqHuwJXBRO0tBSoER81cTF
aFyL+ZA0OE3hU6s6Hs1slOGonklLvG2c6LYWkxsh4kOQwCLrLfl4iy4bY3XgK0ZTLCHO6dyIJnFG
mYo/GRiBg/yfwPKYsYvuHYRUzD/psSocfahaDJ0QkYZ331GxDr9rP9DINNsj90YqajbLjJRalDCp
SctYdeZRQPRvTvyjQsMO2TPEv7mm2rc//OxBPk/lgofA2L+xhDHusONNhrGuIg4enqj0l7VfK2eQ
gXWWTuLM+UMiRs7P4rYBhYC/nMjlDP/VaCh2u0ABaF3fwizpCwqQ8iPJkcG82byGlZdVkpco4li9
W6yW68PY1o8BdXx9WDSKniwYefmxBO0Kp4xJdcbHMQKetdJX2aWLMhDFY/n3dU4Ru7hTPSz3K/Fv
b+Iadg33ueRAMxzPifhRkPaDEmxNYUdEjoZVHpp3ZRLUnUt5VsGQV7EWTVXuC7K0DSS1nStBA5FW
HpybnaCCG37BRvqIZ40SZ+pW1EHg6RBvavZbDmdXZ4/NU75YG0iPFv0xzNBmm0/JdaeLHAtL/s3k
NnARJPgb7vaYwQM0iqFtgobwfGZ7mI66w0Zfq0yX6xGO02+CIdU+bVFYBrJnkQtaeyGMYPeoaizl
gIup7S1Xly38P5yewgmbgXhF2FeQoIgWf0Ubjei5BP3q8AIROCwk7ata5IegGnle/S82GlN6Nnyj
TYbKb0xbcdi5t1FtPs6dpohJ9EZYOtiTUkqLHpOkP/h9URz6fjdxIpo68EQJpmGuqkbuSGE9POTx
tYzO2QbcqLjXjoBEwevJa7a/3/eE4lJmW6RTR0gAFBsUkg8tnOAYSXp+AQRU8xsWEi9SqJ1PHsyu
k7YPRhhv8yDJFgywBSILYLTPdKtFu3Xhlqn/Zy08K05dmCwMUiQhouzASHtV84EoypwqxJsCt6Sr
1q0OZ9vtBtodhpMTACxTprHRHHmTjb3Wk6ovYo4WWQ+bvxj4oIYWl6VsrjmzoKnTVB1ei1vRGgiA
AvTIyPDmEJZMyIGnMU5tKhRiUborp6/Vrm+Y4MD0/fI2cXtjMqHdDVMwtvx5WbPhRg9OlBqlg+hO
6MM9FVUByB/BA5XYS7vAU0WaDHgbBpLQxZY8zfuDdQIlCIL1J9gxB/kb5m5lGKLnImuos4b6je4R
iVzAUAY86+rECgu7Be+OEOMdSYVyLAl6mKAndycjeRZGybevbCt4IEGmJsIYfty+qRcbNSMnMzf3
lw3/l8i3Y67C5BtjKM1skoWwOfpEuNbREG9VBZJFTiwQvHarx2GXHyHJlJ1D0sHfhKFLjvhl68Ta
noDCJvkDa8uM65zfy7ycKtDIkI8sUt5REL6PrgoN2XmvLj/bO14nkQ8hOMUXVHJcerIRSCMKlMh1
YG81eCN6eaEPEf9PsqDgW+XK98u4vag/kJt+Bs1sf5H6MfQnVqjIUvqzhnQKbtjYStcI6bRYAc7f
rJkVQ1n7WRFm4SUt6n/NBfVg1tL/ieiOXizJIze+HrUQW70u8wM82xm8ieRAM0HAlV0wl3hwNJ4D
/8wpzY8Y19U+3lz4F+FbaI0Kr6+UEsTy7/+kQa2nSmlwmNv5yJGzIqkQxoRcNa4XtGrUQ39h5TR1
jLSMhF9sml7Em7pMsB9dupcafs/HtK1gJq1KycDXlVnexKqBlxICY0nM2U0p33+PtAU4MpIYUj3u
Yayb5Wx+3G+ALJP+eQ4CH/+vHYx4RB1LPdKfnPLQPtODBoZ0Uc7jwlheB1Mw2RTnRbyIqZXLrRJU
yGCVilU8heeRdE/J0S9RUPjNLM2oo58BdO8F6T1V83ZKXZOHLHOqNmM0jSdNAmvEiiNtTMlSGDea
/tLtTuqRz9MxLQMkvUOG8ACTTzAznfRTKcG+ou95E/gesJT4kMsYristQ+ur0T/jEFekAjvWLAUO
7P8xXMTMcBspUGlWCqtf7GXQ5nsrySNdrliZujGML/OmQIzxjOxRu215dPWTa9fvQSYr+AiHb1u1
eM09hDMCezncT0605mxrOe6kFMaDU8p9QyP+WQD9Y9+RZRwBtwbBtqH1h1HHSVE32VU3DkLJkou/
kxc80KM5KOTIfwij8kv0aJ97H9/KdK2s7jbkyY3EVYLP5ExOhFMvXgHEf7r9woAYDihde+7tdojL
5b128aCUM4AN6WwBEn3ITAo0EWU7urpxcmjmEEIcORwsofYGUTbtf2TtLw9B2HEy+keHta5DHegZ
ICLcrTHMU5JX11rCKXCugobhK6HZ7Chm9DQF0bX5paS0VNCcboRRzIoL8dnQTflnLxj1JIn6wmqz
jnKVlsTaNzZAm7EKeFkP/KMbL7ISvVbkNo5Uu/VSB8RGg9sHcSHS04K3c9mfeFJYCiEwo3gp7Thh
AtZWtoK1Yu5PkIvkUTbqbjCHnc7rcGZlpOn4GhDw11Jm7guYAGNutNfyieXWO22xR011pY/IKj9K
2oeTDlrIU+eTr+YEpuRwm/qzwfxR8hWaArUiDlb9VnJgExYPn37Elr1irnKc2AZPnn2YzAjgcznD
HhQ/YEzj4xpIwCyojxZITyMcFmnCojGnq513IbzLgXFJsFfJIes45hNZIJFTq9HMEgSIDOSnPEAS
fTEcrKvq/oMUrn5Y7ncwWidTMwmM6cGBrrDSkQe5j5gOT9QKu2GPy/g04y+RXZ+11aH0mzEOybVg
qvW39FXyQEEDuiVyn0FRs3Tni2IpfWR0T2N6C/TW9U2cv32Lr97V2DkUJZi1o3r7rDMr63fR/bjo
zJH1XYaJv0Z5sQGjtbhKqutpQtZX30rIs6C/mzXxAa8XrhGC4lqYBi3rfF6n8xEmoJFrYQnubLi0
5tysZc8IlIMdd1XY25FvCTdKVmwo67NsOivv/Szo+VJ9dJljq+MUKDdKaEdm+tGW1sSKPZ/3VHA5
H9v4uCwGRxhDCBgjLresGf5bP0JZeFrx1tSs+LOHpG7As8C2ryezYb3O/VxaDZSMMkdh1RE1C7sR
Ut8jOdzmp2t2A1glxejxA8hZfM7vdcY8suD4BuN3+BeFslh7hy4FvxAVN4WSKK1qJCznolQC6fur
9KM3nUm85BiTFJ+HNSMGFiyNRUOcYPH3Fm/YOQ9k6qu6b3k7m4QXBWcVlEvQ1IhMRaUwdjRNEh6R
WTeKOfMYcPMBMmUPXQHHY9emQLiP2eMJF0ss7irkY+RR/wR3Nl51wIiybYVu2NzgIjP8vDlV2xFM
6NvLc+yYVkco403CtNeAesHUXEXB9ZAKCvYkjTf+hKdcXncwj1AJiWg1el7h6cKn9u6kyktgphZU
13KkQmzo4zSF8kWWdogswh3+p+bX4osDjvx4kA6auqOnTVXPellf8lHCMaEQDcRhfCxg47FG47TW
wDKw2N0T4kFpvMGTHuO0gKi+1rR+fT0+uqeiZLmr0/eqzameq/jQm9xFRmi5R/W4Hf7jf5V7Q0uI
gL7Bcbaxz5ngudwrDQwXw+pQOtuaDPudZRu5EdbBC2UMs2AFE2j1+bXnHbpVXtWF0mKIrOPCHZwG
p/BSvOIxagggUR8sDXzadDTzPJlyEDRTpHxEO0ZY1w9ZQvujk7zjzLN3RGMfyjqk+JlPCv/j/QiK
La6Ll95yTc+mH1Tml0snH/fT3wYnVU7bbwQusp1QUs5u8KTec8esNnuqQhfmAEep7Tuy8hNyycpo
W4gk11GW4e23PUTJrptWKd/tvI99ymdXF7vV6FhEV6drfn+O21CTBSvFd9l/64WM9JwkuN0k57U0
it0lsBHOh61KXalQ6rlP2pJDTP3fy/CkkGOcRFobPBe+9QEaFK0NR+8iOjLHi9O7prDqv4GmfHp0
Tbum9NfjstYSZZjyHYlznyFuZKhzcjV/gVeiqqcuuDp5QFx5BJo5X+GFMlbDoTSCN2H1NNV+t3oD
80oa2FBzLrMcIL+0rH3iuvBlaCiboQcevaUqPv1gAw8Cx5GIg79N4iGJVMoQyV2rkvfAauC4UeCC
Sb+NII97Ia53xAtASFfvMke0i0nt5mpauj2+Z761gb2TKn6Z7DvQVyrd1STjLMhAzH0Zo6IKY1NT
d+OL7tO8J2ykKEx+9KIGxQHmrE+HFfwWc3aw++tJ3A/r8MEE6sPJvIogVpfZzC2BjXvfDV6Rlwuc
TCif7rVG4sPTytgJFrJkye16aR5/02r/xcvsQ6zxhEnCZKUL58ebbzslPSZo3Ynnj57W1L9DjJxg
PR5493x+JZNqBnX7CSb4kaX31G/eYT41ztdPWghgA9nSBCKtp60RELEV06QEUq3vek8cTTKp5rFf
sb4zPTPU0aCG4HAZk27w8AJ3pIPy3PLhw67Opzp/e9REqqzfhbTia1HWHSYWMKZ7J/RWG9iTinan
qugs4nl+6Jrm6K4vaCPHqtBBe/muU46jFByat5mzjhXcSluwWGzHS5ohj3jv+zDSs16S9DgMFxf8
dK63g4k9hIrE6UTdxG3+l/VqqlytvEbE0MW6HIIQ3XoMCFfg8eMHedTC8ul8dr6XJ0P09EKTHcQh
MiqmUyTi2FSzaESN2lOp/6BKIe73d1ErLslDdSciUYLxyTshNZWRH2u6gPJnrSARTm8JnLHqsZnl
RUGCroZvw/pfHSDdeOsDODwY0BcTwfCzx4BgHXUovw5TUYPwdcBFcKb5lXchur/xY3wxoVPPwI2S
KV7mqzs2/eShNJAGbYA/UT7rNNttJqrOqsqQGGHOOb7x6kQ/t4k1gkFeurv4cQ/7apLEv7XO+jU+
37SJGuSraLBGzDAUXHl6RDWIdJNuhzBY41gfpejsy6ugj6esKW/9KPwKUC+qOscNoDa1HNyqXw4u
ZpkqhM5ldZRj3HECXJ4PXMNiSYIVK/Uab+keGwFpw5eNl/nl/kvGqWfDNQ/8XT1JtwUa++NCd9gZ
8dBusxj9H7pNF5zxdP++YUxyG+yb3hjeWt6YzrabkSF+0rOLBTu7lcS2fuLGJD0yU5u6DhDWVLAr
VDVxYCj+KP2J4bJ7IKv1QGlQTHwH820thhxTaeAuNKillibRliSo53HCdTmJcfEIPJTpkd8fwU8o
dVFVMYJvjYSNST6vv+5ZFQQtmmM+/yqEL7aJDQkjlgjNxmO8pP7sN3MC5+UtzYPJCtoa5bi75oEX
QQ3nuZ7d4rnxV03/9ujmhLNr7jhnmE95OaLuYfDTgRKiKkitWzidlMPjjJy+0hesfEvuFdEu5Fim
Fg6FM/kUke+YI9YNqvORs9PkT9lGevEuWC9BqMHEtd8V2kbQRDePssQ5RDMX0MaA0IAMZScrs+1n
nGyM/id/BtL4xfCjJz+WJx8a9dnddl+FgOSgWwPsSR2tjp7H8SvAcG5YBe1IR3mPXwE5eVlAVyHy
AkZMYi2dEI+HTsD49ksowLisqXwtKuF7KAnNKYEGMe/gLdXXyW/XSf4eMZry/F1+pynzblz9tkM6
UnJHHH6UnXrJqZyJSZGCKRWcMu9PIv7mbY08urrly3pe09AUlddTJiSxtqDzntTEwg2ecpzJvts7
Cx+foR8zZsaJlsw8rPoJCUWi5hfifOIhPzoswTKXTgdezG9PeyM3nTCv6MQgZUVhxwg8HdCvFi+r
ra1MxP8LHHXv7qhKoC9CbsMCiLrOghcKqnaDBrEbiTfRHGqidd3WNtn5WTqJfLv+qAp71cCDb/m2
xjhc5Y1fZqHJndY9NDZS6AEVFVHadP4lO55jraVl2tACKFWlAim3yXt601MFH7oG9bHOb6dNNi+x
BkAaOsE4S+KUvPv7czGi132a3bOr4n3MtUwWr+o/JwA1jAbopu2+ttipQUFO5uXhnuhJqhxSIlR0
sI9rFGW9wlhyBTUkO0aqbi8Rwj9s7dUGDlI09C6AhUfCBS7xeQIaZlFGMQ0zZMdfzRbAD27C9clx
xuDKc+JjpnIYl+hxVHJ+TYdjaauUC+F3dGxA7kOu2FbFmXbGS05K09PSOU6CjGwcO50lVbiET+DC
S0UvJEvzd/wPzXLq0Kcf91x3aV3t0BBR1kstp3Q1MHJOH243cpmGdp5hk3R02dOaj//jlNMrx8hC
NkJ8RcG8BvjwM/U2doKTGjQBXU0BfIvgU1MFrgiKiMFWv0UYJrOpCQeZ3BCMP86YmQwJSXsHMHvN
7RqX3vyN95Jdw1g1Ky1Y220fRcCSUnkQ6mG0YKaVFt2i46kyKWDOEob6ZNkWiGHK4JkpgBSQt0sn
RrmHYqecgvwcapqvPSFASXOCAcxqbtWiQwACXABuUsLeO4A7d9XAxJuXd5J/G1tKVM67PxHbdebW
zPVRtGkd1iz1KnVoUVdUGxgoDuAb6zes8smLbQMukgbuTbYvqMNx/ynj2Skzt0L9zXhf36PU/ydG
rflau+XgRQ+5RCAxgFRDpJk0/tIdUW6bbg+uBtSsVMS/69uoXWtVphWSpkcLAGlZbtJ44VLNcp5S
j1OH6BGtp6UG1NZsUBN9he9kKAuluRBr5xLUSXsU3a8lX66/2gsFxMhcfjrlhbvrDYwMsVktRxtE
ArMp8g335vyEdAmiejEr47uYaITryR6NvCVa/q+heL1TcT2fUwQQyRNOe16ZqRU6+bcO3yIMzkJY
CWIlo6iV3vs/RhqFVy1l1K4rvAel9n+KrALoJC2OKoVBf3qaIJTrywr1a1YPnVHfvI0YdvbEqwMO
MNU7wZXOm/ygZzCwUAr+YDScufMq7YmOb4Hj16fhd0mRtFn/AhLkeD2LXITdbE2+NNb4R8jwtt1/
x3EQAcX/uUeWscMDxeOEgy7s+xxmJV+XthAaWG3h9Aj8UwWoet0KOYlsm5l43CkPxgFLM6OD7VVl
o9P2sYroFZ2ByScd1r5MpCWDvPvxjckIJBfto5tL6db188sbzh19q2LW2oACjgGn67saZCJ3h3Gl
y4qz73E0Py5jUwggcoYFnjmS/kDiDe8uuqMOoNd6csBstlXYunnXasu5IepnI52s9s/ZwWOJrg6f
nZ0nhyRIrVKVXx8WM8kJVGeUB9CKdCxKO0wT+IimEAIv7gCmPdYkbvyw3mE7txuqW0sU220cyPlN
/0bCOdVoRrnm4Uc2R52nUsvm/Pl8dCJER6z63zBSixohVqV8GTTQsZtBKxvHAKMKVv4VuUD3Dvri
jgLPuLHVKrU64MgGybRt+Kmm2bwlQkH6HR9LNLWguBaUAk4PeEGchNSvyVVtAF6+NqjprVPP8gof
6HMvKE8i4plTKIZTTl4No9UGv5LO6XQNdBIMXow1IVE/pjStBy26dPqRIs+lnLPXOlHVjv/KdlXM
M8CRCeDfkT5pOdyb2hovmkSOyShZ7mNCuIqOXVXdCZ/op8X24S0XbN1Q+udr4uJx2m0vm3fFcALH
FPhPLT/lcyzukLRW65s4aq0mk7maUyzURPUxHOdeu0F9OriTSjV5Fyt2l90zGUxwb9s0mqAbsmXD
asSAvzBt4fWx0FiAOV8k7jGpBJ7/dOPF/7XUCPDTCQl2l0OZk7Ru+a8GTjW8EaExWMpAOaa2k/+x
Ib4siUL5uWi2Oc5uGTqNirkDYl8FETeEHfu0JfjU4L15F3UJ1wPyeemHu6UewuudrTz+VKQMgWKi
kKfhe8Ls5wmS14hxEPMvT86nM1ZtKji91mvu2YrzA6jJ++IiwbyO2DqHuhB2YSRNmIMAog+TGku7
shPCmMS56vzYj5XuZxsPNcl8kansoYvzVJ/K+Ks8E+zfXkUPn1ffTB9qyCpbNd25o7duXR3THjIl
ZXVeW7KMJO1kNvRqm6+pZHxT9MYUPH8dBSJKGnroBMsRuTFTWGzxIMgTnvK/chU2gZyRJOrJtVKf
lP1zc06zLqChsGHv7qni5tLw2LAr7Lgya3diHMyyM69Hs0YM09Upujy8K+8LVAtHkGnR0+6IBu2H
7/Mu1Yh/p2WIsHrlVWkBmd5YZ+SwWLzZgXxXbg7RFxe5ibLct0FvaXcbaFsDDRV1F3gfZAbhP2Rp
ZQSwuZpMEcO+H3CBRXv4aDP1i/dt3h2TkopivibEa9vtZM3chrjw8HYyidQQMYS1Yc60Q9vNDi1o
ftpQzdbVfCS90CIuv6BHUGfdq/64r9LmnK76hmcf+z76b+/l9hQJ2Y0RYG9ZA5lUxyKciNIgDx4Z
OSDceLWG/nt2KoDyjudKgyxjSoZxRTCv6FfkOBJir3YiMwdJEYyuDRpFQLk+rmptWYWmtY/RmRBO
sY0bB+92dzQx6gquCoXguxV+624ChzJ+1xG8WogDgIyNV37gX//z5pO0sP57xr6h4ahR/wYkAnJX
5MYzsUYI3lX8kSI3mr3+P4DLruHHkUshwO9uS/SnDSv3psZs+RXc1aIBp18vlHmpAbZ4kD2A2FBq
z4Cm0mwkZ/RZ+bryDzI5aghAWV4idmbv75CNsaGDB86x700sxM/ORjsp4Wcl4pHFJuH+5tiAC5fr
0JZZIwD/nT6mVQ3UALfxAE77uZlf1RoI6skVbq4m3ix2rDFje7XDI+HrI93Jp4AaokgKL+382fKH
WrnTZKRV2BGxH22Y6EEcP0J4lv8qIN5aSHSw0GYlRI8g2EOZMwnqKaaPW4hzJuTsOgv64+64Aphv
NMZy5LEr4A1QNsUE2oC+9YxrJOC9HtQ71UJfDPv7HQaL7Yf3C1rLxrCcx8U/TILw8/FaTSgbz/L8
KzyvVUyHwDhieaECooPG+MHwvTy9ifLbYcJeDJvhhu41cKQftrS23K3HYqSEDo7fwGn5hYOkhRGV
jZSYtXmVbcVKOcEXTJ+OF835YXdixBNtPg4OM3XRFXRZUno1gJs+M8V+hSxEDE6UH87lEtAAmGv9
eJK8VyBK9SucIQpHjQynVpN0A+o0ld32hKYl64H1wc/fX5Ql2x9mf3KNawfjrUY+a+8P/76QslI4
IcjIVfM5YvYQ12OG+ZHzpT+C6LUoavs9ZWRB7Sj30TwjObsf5IbpWt/+4KMHwxUOeSz1RM0lRZ6m
7FxPAJwiAdjSpEONXxIET+uliGIxmIx28IaoUtgBkPH/4NZSsQ0VZgdMjQaFolGk4KaCPmKU2yWk
ogyRydLXHoV2enV+lw7/h4Xrop65a+wvy5ZX89W0z0KU2h/mxRxZYJzKzK6HxINZO/Zz5VCgRIgl
uivfv1wmxV27ChnBkgePI4hUF8YGcmp4WdfJBt5NfLgmyKkZP380G1Aos0wNboiv3SGqGVQMQY+S
B22t/pgp7f/lF5WpwZBgLuLlWHsz3Xzjv0zOKxdly67mSTFj2Uuz2xIAoytASy86tIxG3/P8hTjZ
kOZLZcZ6efbwlZrPUKYWGf4UghX745YcE1KeKKXIjXlgdLKrbOQwyTTK9Kd34g3nXex+kELCH5O7
kzK7zHbh6qe4+t8Py4WOd9Glyhrn/Zw2jzctwiwV2XGO6ysJZ5bFr7CRd9n0V6zLU5zgphQLXe04
+lAs5DUZWQxau35suPOHaHI2rvv9i0nYeLXtOsvd5AF3m66yoBMtS73UvS00dR2kg7Fb1T6FC0B2
1rLg9Br9+0wxyoA3vzXeAjIxztX78AHhDcWHoerjDzpw+T9Lj2HfdYIN2J10WVIetuGN+QoAsTzT
nHaBEvqVvyV7iDF4VUyLgAWmEiKdBfSgN4gVTqwDnY9uGRl44ZR0DYElqXa+3QeZ7m8w1LxKdqah
c+eNksjW+ooXy1RacjjZKUMnLWoEEu8ecyza6tco5AMvRpZhNW9eCnhiV1QbT7DLqQIer9ppsGPZ
ql3hLhO4HkmOXNmJ+EJJk1zcNNuMO1KCXOBtNmBrQfQ6M5pBQ27HPX3UVRDeqjiO51IGSoJkpJSL
hjhvZvArP6a7dbuz2OUXj1dqUlVOg3fTqGUDlYL09l2HEN2PlpUMt4UU4ql9OUgyx3h70jYNQTGZ
Gg09hGIVCNUnw8EONozX0L91hIEHCDU4kFyaz5j8cRkYYJft+MFtS6w0L54eqnNbO1PCmLN0M8o+
WSzBrWV/AoBanAoQdv0K37Zap8UVDpwRgPLsge0e4TO3o+pgkNMoEW1fy7NReDLIbRDoislP/sNB
no9FTp0eygWvBJytGNg8wC5VtprTmE7U7lu+t++uY30ixc3EYeKAPjJD9jzmFz/GGcQo3HDD8Dxi
WbJxVF+qy4Ypdjcl8VmP+o0CCft8KG0p0a/XzUo70K1dyxB2FgG1i97Rn5bjApPTofTb59MFNYbO
96G4X2KZ8E5SvaUAQCZSudG802NMalkpAQamTXHDkzwH5IL1yxE61FQWx5HPnFbTT1vtZw4xQf0/
JDNO3z8Zz/+dJnSGkG9qb9xRmkp3mWa9w5ES85ZDAwesgc43LQTPZ3rY+WuFeBnnJwhkrkT9A0O0
fjm6Z22b/P24ORKyU5JynmX4ARymQwtWp2qBYDUpp3oZgGPP6M7RhI9V7gjqQoIR+uiRDnZpcCSW
YJNJ6KGK1VVvpqyo8GouQ291GLZyZNfi3g9ZjQPlUZiR8JbBlD6cbMF9GYNFVVLbHC9R8yTLnYh2
dMC1n56dSJp/BGoDXogqCH0gSosqG5EtlVGSPkZ5JZ3UTubtHwhitVK174EJzBcaIvXqsX/COwGX
2H4pNcioIoJKgXCA4rqLARq9lScX1DHA+iZ7RVEFChNWOsTEIoDjr5+DkrnfouSavPBjizthqQ50
/WiUGlHjEaNJFIddcU2KxrXWU6K2W5UpJFac5njE81RuO8uxS5QtyTL7tpdCYP4QI/Ju1b0ghAbx
qlj9SnjTO8L1zJW9gSx26QKfZFZ5lAYgHjT8kkIiXxI7l0MPlg9CG9JFrbGnsWBpA/dxNScB7ci9
92FGJbDUR16LlZf2RsvmfFXFPo24c+30Pc0/7eVUSjz2P+dLLxLAFDEuoMvzX7oMtoUlOcDCu2rT
RTcqAAq3EozPutrCK8BFQxpFuK+gshVDI1GAu4G6QHkbi0VQ8qZtPakS6B+C9/NGjLM1/Uy3qzUO
Vcb1lwn5rQ8tIyaAFD/g3MiJE9Rxs0Gtz4dWK5lsHI5VI2uxmPOrmQP/tLpAnsMiQYBD9dQ0YenL
LGaSFdECcx2ooVX3Iy9uYz5rk26Dq/BKxZ7tjHknvaRFNSElCeDpxdJAujl4fjVyBsOWVz7kjHme
GLJUthhr5FSBHuOlXoJWACpMEZGnFnOPrVTPG4H0wqNLHs33S7i0UCOFFeVMEblvAZHbe7ScYPYz
RbXygtCR1BpVoP+hwlm87O11IqmcBudtx8imkCHh8m2Mdg/fnv+jGz7uE1k2d21J6LHI7KKC21Id
LH9+EowrofGqj2mPEcTELFWGKOvAzCpuXG3Z+rLrpiOh9hMRhfbPJMF7/GgIZNBYW96HrZVlZVud
e7JrobsH0H8lUc73XoXCaxyHAW2XW3UDSdg5Nf4GNYy0hNRKT3A8+G/0boRT9EWWmKcFRRUBCcb4
lY3LsNYv237H7rjswwK/tRVJPevHJFuRrteCeNuzeozpSPABMA3O2ePkNzolJT6LuvDvoiynA5p2
jdsTgF/hOn8ze22ia592dsNQX58FYY2pmr/hUED2lEc44RDCdnkHjw3UWB5xvlhbI6tr1LhLcgqL
MXxV3houC5UNzQ4I19B2vkehYqZfJEqGWrz/W9eY84s4yBxIvzmgndUgNP+Ign3PoXydCN4ArWfB
9nU4X6/9xd6d5KIBm9tW+gUX0LbMcWzTxnk9EslgWo5UzhBqmscr0wNpdjprbj72zj4WFNpghiBk
/k+gSdhXi3kSpwEraxGviBwYxA/lpZij3QVqk+6c38bTvTssbStlQ0NhfKuSb8d7CRRc76vBv6Qu
HLy/O6LM/HJn484qzeVn+5w+etD1CBDD1e8fJi38R0fpZEq3LwpqAQJjBstJSJ58P/H4X9P/pDC6
hyr2rLnJ2HCoe3ot9lpwD//FtL2y26cGuH4Fe6zOB7r1PXJSmcgEgOJAxxHY3u5+1XvFNsGskndQ
p9ByOyr9MCKcRCCkQH6vgOAFJbEQoO5D3CWvONoWJPc3MgJgXRBleP3yX52omQvX2IKMuAFOZAOp
2HFFTXCe70+r3oqpnDJ+QqjYT2BGuxqMBWOvnkKmqyOvS54SWkKYu/vGw8O1mO0jKaGjOeLXBpNl
fWWlRD93x9z1RcIQ9LOJqIrE0zBuyiPV/rmCQPOptm5xXrg0zgHdMW7BZmfKG3fOM/dBCEE5LglI
fSf9CALFd/3opI4q/5WJgtYlgP84ii1auM3ZeaEziVRDP462VnJU+9Es83JqIsoQOdDf63bHIqGm
fHFZdI5AqmUuZUuxGHHN/jo54KHnWe7wQKlzV2ypaW6DxIizf5xFpsmDJXsqR3DBLUjziCIcz7UN
5rZmiFcsyTrPSsnY4iYQM2FpUDSwETR5ajOnmXq5HLX9dLBZp4EZJNEgTCDeEBTuZ3mFTH/u+tmn
2GZucReMPyreuQQyDxZ8w92EWfW6Jv4CTQgMCbmLSrnquKDljd/Nk1eoPeLj4wy10xlSes5asO+G
5UKfqwfcDe61cKFds0W3jleTnBenhQ7Uxpua7RaYbPjwWSVHThwrrhboM3yrhg53TzjrbeNSedhG
foeFVimjZoEBYxeyAB4o7yQ5w/x6/NSHekJXyd0+uu0DJCA2453C22+GFzlVABdo8Kb3p8fSlz6n
hrmyXGMl5OHI5RynIDliG5s/c3XkO6ed9/PzgI7NX7r0oPdqvNIWcD+UcHG7xOYS17LyhpWNsupk
/BCsK4Kh6Ya9A+2bjSeLFwzu9ZhjXt6dWASQYlIvJbJT9D5zMVmx08ptM2JcgoDFWzydPzpB4p7f
DchDiexmr7A9i8JTrtDKBYBL2vlj5Sdqa+Dw+0Ud9Zz+Yk7jq98uck2QsZueI6aLe40K24I07JOY
7/PGo159GVkJaj/Mv1ywpffaMTY8mDvVii17GuhhTuan1IT+XhtTdcWq/omoN3atNglddAGs53KD
lE60Z4zMWqh5+tZHPAPGDVylBVtOxbqZPkJPZ0xq8dL5lV1r8+dUNnxVZebC+r2/5R7Tf+ToFCxm
jYvxFDVfbFzDxu+5zf6bh5c+iGhcAZw74wrhWqy/4V19kVazNiDoRmJdhywo7mQvydwP6CpGkiSN
LNkfPsV8gL1vQB9x7pe/PA7dqm5fhoNa8CA2Hj+Gd8ISf5Nnt/QMNvi12jO5LgL6oDecBxl2kqCk
UlqyPsX6hDfyb7t+keqakDrs69ljc35A3JWDx7YVDfxB/tdSc9mlFUKfAJCOyDn2N0dOzzVvgx0g
0ayDcPmHWoHFlE3ZpZy8BvPhqVbMk4f59e81cgcyyfchsbrQDuFzmydW7QtqwSlUqwSg0+aZY1kW
dM9Ww12o4ewIxwIyRry2MONMtDCTJIGQEJw9KxgCtYXP7AUvDHZN3qGpTA7wjnsQvDcyxYCfb6xg
hDEWeuYUe2bTAOa7TrAlPYky5B0swKnUbp3GE2jAenl9Qhb0EozjGf342m6j4DMMyEvilUxPXeLM
5eez+YktwE6mrzmtNLCKnNTMHr9yE5odgJ3RJaQISO57s8fqxEmELrIZoNPmcqyRaHTaJyJmiK9y
KWC7MwX3hIxRrvFdFv7R9gPRAEs9cr7wsaYbl68FK/yP3cB8Erzqx0KGQYAeP9Tejw5p9LFtz50O
Zex62sDL38nq+fN2URTgtJaEc5Siq8XBOPh14snqQDcBHRWS7XmqOqwEJBw6FM5TobgP/0zfA17S
LNURiCdXXejIqMt9DL7k2VCD3zU6Omm0DaiMRJdG17fEwTMglpGMB6VEfmsp//upDlUl0yhJz9Cp
dRwyVjWYaoctH/X/KtLaPgt9coRmr8RNzOsO9n5avlGk8sRFpZ7rUCOYZyNvTYVKpwsAqEC/YTF0
12NYkdTMlV1tP90v9kfF8PbUM7aLcxrTM0Jnaq0nMUceRu2TVYKCnppKDTkXp8vb7/gMTKIMCdu2
PPGLQaDeBUfnLa1Q60/73hfaZ/rINGeKDxLiblDWoOcpquL8rXhbkD9VGPYKoo/34GQvQmwxOQuL
qfb/jX8brGrKbZQkGFHd/1C+xp5Mk7/xtG2JKHSBHXEuqUqS36nQ1qoJOTpZst0VyFStGMDMpEgc
oAZNjPmrD0RRYsSuOXumvHopR06eQcUWjExlRmYmA+Y5siT9DJXukU+ID9qdApNTHsNFeojQRZhq
E9FCrphlU+B1C4RychX6Xc+XF+9I9kaRxQt96MmSghp2kvUVm565lWepNK8ZPx2qaaJsYgRNs0zK
wKJ7H6VQsWhneqs1TWFWq7U0rrONg8SmCKzD5vc2ZlLg9gdrxyVUSacLnXW6pyi/UaPq8ygAjl7u
IDOBateZp7gI5jvRCdJKa4Oy+LEqBENovxXO4PpfF0Iu5EBeEUqasvN110zFG1xGvCTjntkdRnGL
jDlCbIxM0KtCiimZr4STlEwLQYQknVYeJOU04qghb/d2ASu9upA84Gdxsvf4vrYU4dbCs4Zv8Pan
GWPOyFcqzaOxmxD++ALQ+PDIsnMCGzUXuaTfDTV3OtSYjiHvF6HI89t6r7qoi2NJZMJh1f0VpN8u
mmoQPXwJVaI4yz0eS9mesgb4g5d9eJtzJdp5nUXyEA1bQk8KDADLpeqnCZnVy+Hp0BWIm53qJ3iy
2HOh3DD/wi7ayYrQzocmR55w5Y8IJWNQhUydKIrrnWLsY25QuzxWOa79cdy2/OUHfEilz8gR43Vb
bXK4X77VD2mUNwZagRqekkm24PKy0fJDqtQS2hQngFvFnMt+IGT+Yq1Xw95SLFYPty78N9tpi+nU
LKR2B4CjbLjV0UF18U+BYrJz1HNPRO4OoVfyca6o3zvTkPe18vjHPI3d5yZUwzwKpSjWLRg+g0Xo
f5myLqSSGnAiccHqD9chJkZaXDmMa7ugPJdiNl1yMmvhgSmBi8aY11TRdJMtjAh1H1v9QmNP9aJk
xgpuQnd66/FDTfQd7oVy6/VjPYGGZUNb3M5402KoRZDKSQJv21toKoKMwWezQ1fF1RblrIPQdx3V
68BdHDQxU9u6Ak2z5FxcS2I3qkOdugb+siVGXDa2CVvauQnBpt8BwiVjLILaCSPp3dA/R/c8YpRe
s1Uv5wgC4j7A8oyfFhBLqpi2wLlehBoxWdpI+UKReZF2TFsgVifD78UmyoSihHZR2QPxEJ+mdIrg
hzwxCVmdBTN8I2eSTsOwYaBccaZZo/cl8jBP9d1DsWJ48oAbe52Yfpobm+Ttqry2fWZtn+VVCwlg
tnX7dTDJ7QILmACQkVYI8oiZ4YigDylBmfllUL+CcaDM6IObDZBQYffp0I7VQ89apO7o26lG+Oc1
IJSFvcyVnXqFdc0pauL5IlR6Yoln4rdaZL6H520kLSttg6/lyoZ1Vug1hb0JQM4GsxFUno0RpvCY
V28pmXVV9fNCedyUWE9ahqBFYOoswRdJCAAxyK+v7NGNp9w5+SV9v7Zn8W2FMljpUd5aQPQ2eXMx
KNxaiQlxXCU1Q1TG+JH56kYCVD2BzO4edwQWBupB4kuebI1s1p5hSoxjBVBMZs1N0fDM8qOm63m+
nZQXbMYcz5m5yntAKl5d9FAPOI7AzggF3po8qJknZe/QxSB+J9vylg6i9BE3q03FA2GMvpAt2E53
Wz7/a6EuQdhY/XHQjybNI7dtH5upifa2N901mFi+eNsbCNOY5v8J3SO4+jC4soCO0XptaInlZRH8
If1FOLz3JyhzOt1RcwXl+TBUmzqKCgrDlo+sDVWdPcshOjNShPcYiyC29tGzSf6nDgb7lZtLN9zb
VFDYyivctvXtYkNLvtP+umqRuBqB0WNUa9Vk5ljH0hIJdrdIa5saPQ/NNampDNzl+TEUncxwfc6Y
6k4mI4JnpqKU+EWClT6PVAelxG0Yg10Oo7XtLmFTkYRoicghyemlHtpkmiSXtlSZjo9rkT3sojbC
Y4+2ipuo26Yjxhw3Uwloe9EMdO5BNK8nhAFPkHinEkf5oOS5oPWpI/GLhdDaxlmlM4XhhqiPIcKV
xmK2UkPLzQ+Sh+d8GUJs1iwJ1Mnu5HndgkPDuLDMBaz4A2/htcx3IGqSAGckEq7NYX4yfScxpdT7
r+sBr2KOHKUXvZAURaq7OUJaN+KrHD22eJ5jVQgwpHtWOPmCodiVoLCcojN4b/kOa6nckVdhCjlU
yrSwwL8f5BdShujMBV76G6NRPf/S3QIl5gXog5G+7YUHM9HB5PYegJKA9pirCXj08Ywh20ynHJBG
ZQnkItvgpdzKlIbLIt6ZnJ4k6uwaujRBxCEdYNyynLhy46hX7AVIgHLKzn8TavPPPQX54RvD181n
t1MoQOYJNNInQrkyDOiOWBrEhKgNPtuN2wtKZqRYDhYGAL9GZZ+3X+j/JErHHpLBokaLD4sdc623
E/TA70izSKI7p7gvouzEwbUqnxvMXyg6stb6xTrQDykn6B1ojq6dZQr02mrBekyrs1VohLt3r9vl
FnUOwklLVWlIHjEwJagDHB69UQ7ifNXUnTQxRHKjIY2cHLzvH/vIQ/uhTL5BsGODEjKOxiQNuyRc
SdmaPbSejlctElfbYmGcdLA6YykUjOhyW+dnnym1Sc0sMbGljatDqDC4SzC+TbEViLc6dJU2qt/j
Si6A0ecZeKOijbEzowFKREY2KhQ5paei/fDuIWPXoBenDOZzIf4/JJxHShcvcXW3y+BuPAm1GnxC
q6QmhK0iZn0dO2FSZ7AYLRjZnIyLlKm/sezXkMHjpKnlqfdQgd0qn7bgxN0/kMNU7L+x2aW1Ps4A
KvSzRVdx6UftzwSTfv/WP+ezTHnhJxHndADS3Uh3koKEiuikeA3PbXi3MPzytQjg/yTI8DkNgh0f
CwTzoqbHuarkGGgDLxdgDQAc4WQbjRTnU8sXcBk6QBcQBAt2ZkrlvHT3aqyFrlzBlbSvBpzWN3Fj
PAIersplujxHzUWgSi6QmLXDoznJ6FBjelYIba0sOsP+buRymJQxsjf1Hzb2w0zPBNaXa/JjwlR/
cGZ/IgarPB32cIuguqlzQI94A+NHkfGXhypWcJuL1ZxI36TAWBhViImJ0j0iM3fa83YDbbtiA/Hh
wszr1VBY/xM1bYNHP+UkHgef5ke2jea0pILaWBLH5rMTXIurOGqbI7AkV7SFaN2kj+dPMTuJ+n5k
X34YXg/Z7GLEFqh8rrspEu6wNe7sc88te1H1QJucdcAxTK+aWBNNH77wZR+Lcua3rmaBsEkTwNGX
nIfB+klDPGkOuI8lMNYmimqRrH5R4sJGLUG6YaA3glJdw9kEjf1/p6SOmWeO7P9aA5ngQBtyMYSF
v++RhqkhzEIrGm4Izzb42bWf1pflbTFNDV/TWafbZ6b8x3cJ95le790KP8UUlEgXiHSMrkRo/P4u
TjT+YwCuSdxHjPz6EDIs45ELeBj2g6qFOHtmxcVOA5s82yZ4exskA9srmuqh9ZaPSGmtUnhIGSYU
8NMCkvzV3dKAhzAgjduhZszs5v2dIcZd2hgrX6/PvERzTQ2I0OwPSeyrcGtGnkcs/ggN/lwCgJ4p
Edzo2MFnw71WftrQ9nhfVv1RciHpQqEGZhSRCRYKyJEh/yAwEA/m+vx/1fwxCw9qNHAlQeM0otZv
/B7SGaaK/KwaAdabfizbqDdmAMcS9kPxaSBWKtHZC6mQlRZf2hcBRs1OIrMSSaUCTn524vxY2TsQ
mE0Q3yc67UkFH7hBNG9M5BSteUSzJL5QtBbS9iPIdDkXzQYPUVO8mKLSXqq55w2RZSsHO2RzBkMw
9JEtFZ5+mZl13Uouks0QiiptVvPZ+SeAp0/hL70HHVjEw0MbTskDiQx73hmjaglhy2PJClMB+Uu2
SEt2XyGwRk9VA95sKKoXpdd+nbwOxImvIIXv5wxIfYMwdazKRou92no0H/frLR9Z0mTA7CeipYXz
oyos4FI7gQ4DlUhxJfPyn4pjHkOl5zbc0lfPCyiXirDZdSCMBfwBRuJY2UJKIOb5U3jlSrdHlbda
ZXn8oddtiYElULY3QxPqsVS0UQufQM4c8eJYZyPb/mC95TzdmJZbJ9z0x36tH5/hVvWsL61L29yf
BEbzb/OFdEpQs0lrMmwg57P3Z7BncLt9tUW+2FyYsxqgc0qMjmJpoxMjvGr+FX87oS6dsKHtOCe3
0hoRqmw8QIsp2QSDk4KHrcUPXKE26EHZLseF5g3V4I3IHNWXHm+mOtQc0Q7REA3jjIYuPsUYzeTQ
BwAQrDepLJwFx8/LdoXKoOb75Io8xRyAwXQo7xYni/vXjSPyHhLL2ARyZjrj+OwmWMYQyuf1BGMd
oeHhnEqaZERrdlezBRhgFBogVeq6UoVO8lylbyKYjldc42OVi9fKPAQ58b2Hc7fJNTQT6fIZQhUu
7sHRtwC4Mll/sCiMBm1Hzt6rkg6rNxs9rahXUQQJrl7mzkFXoeVQhiLp7+VfgYt8JZPxiHE5XjLT
5Bw4Kzplh24VdpfgjS+5kvRP4Kz7PJK6NmIboFHFG01yerLjQOiLrTlInDLNXj7XTQ1hsShCnwlC
iKlfpuZ0oKlUs+PcM+5mvtAQsvU0/jf+zAbgkNBMXOGWYnCENG8sHYqYyaXHVX2JiwfY0Dcd8voC
r01R2f/C6csEN+FA/cCmLAyzrqr9x+AYXNUVYaKNENx1otlm6JQ0nnyH1KWMmWyKn3/lQMJR9Qt2
6XGoPHFa2CkrCSdKZ5ZbbXLBLIXzp+ScXAC3g58abCZFM/XXHR7RHk0KsyRxKqItMzY+cYVVEOpK
MY+MEOqjBCufz47eMaNT5zbzN/jK1vQsNyUSAAGzCem161AFINiGmcx36awdAKuOOUeUoT/zCMy1
HtVYHHjRPCWUgn9wvVuuUuwRp1WboRI+mXU4BP6CwnQcy/PDUufriyq0QBnpcVvPD+kN9FfovNKa
4Urh/1BYPMMCqQvOuJJ/sN+KZcUQtwH1lSUv8ArCNHBS5oGFsni4iR8DYLhfZcY8Tiep655Rmn8x
X+w3+ejrqUdLsGzvhFW8TefPN44Ns4OgDNocVrG89Ma9gDVT0yXCkDVeNi0yUnruARaqQzl91EON
IJQqXJOwmtNeJnU3Igt6V81gKaVGqCCGOT+Owz6ECdynyn5QigDlg+xuMDlF20aL86Ha+r2c59Zh
79WmtXle8rX+jGrlt9aLQPpdbuYlb+GwSQZjc30xykdIoJQrOBMEewj0OzJ+6qENmL8A1f8kpyVj
vn/JS7bVl8OUy7QaY15DPkOTYwZ5ZXk9umMjqRIGyHd86oQTRXlwqb2LPFNHxmBViDGE0QewuXPA
8Z1t4HmIztBivt4JZs7cn6+5MlTggz4nRWAqr0o3aY3qt7Czhu5yGXDhl7ncXFWyGcLncqyxfqNp
rdZiX977hvlwC5ogaNd0S7JWtGdSe95cnBxd54vK9pb0TIosHmkxx45CITcWh1MzIdLeLvqYf159
QmHbihfRjgA4YtJsJh9xXNYCW60MmiuRK5wgxpgWuW5HwB4cSg92KA9QOmMLkIcm/9lnwBEojlR6
UKsRv9wdxVmuimHKKI6+TSMzsfLHk/xkCcyyWgWjgrNvES/VfOdf3+cSZvBv57X6AuH0NwqFja8f
3aUuidmkEQl7uJg8b0LNC0NZAxs+1LyY4WFc8mbIhj+2Jh9TlKBeMHyhk2fZc893Er4cxkbqAZj3
m6CSEY1FwXgOCqGK6+hhm/B1R5etrRIBeJrfPGJmOOxYZd6AWlRBoe1VNMsW3QqIfKom9lDxZEqR
gi2LgWA8ZEMAFc34qUIB67TY0Sda1dYF7aKisnOcE5c7YtCxkhVmYU+7PEN4tpKetRxtZ7SDdtVK
r3ilrBkWgo4J2mxbpkb5YikBYW8N24+u/4154sudyqe7RVPbu/XPpZy/HgxlUwRUdsUdeaRJdTpn
pdW/QlPuaR9RgReDebt6DuAg1i+GmtJkPrR2OHEWlRTQ5og2vO+turMw/O6tLM1lKrg7iHMqVy52
t93IQeAo7nlwysLsUKZ2z9VwTo9j0JBZrVQzIjhixtw5OPGcYqQnB7iNSIvcvQDEvGC4hSBjZbTO
or4xAqJIoA44HK56ugfVPSCVxmkHoCrYuMkaMXcReBfEnRjar1YfpOxhj6S4Lt4+2JCiFfj+3GX5
3+DQFFJSpLiQ3ilggwzb5yW/0Ls2pU6+LUHmfiC7xi930WbhC8Q7ddO++3RUMIt9nXAtwQxhbSyp
00OS0Llkci7zfZIXDjr61yr43Ja9XNn5DZglznmfZwSUBCYq6N/bc4RGyq/PMRnaILBv6GaM6ArW
Dw9qiLs7lBwlZg9t9ikSKdyhW2UxFQQscw2QCwZKURLOKlvLKO7bwqyB98SNpS7T40sW9Hw6OudV
/IF7GrM+Exqpt7GoAuZFIQylau3PJs3rgb0exCUgrJapmCzWfQfJEO/pCDz2a5b0f5eNNfu51sJp
KWzWuxFUxJkiST2c0tzkhT1X9VnuGbuJR1NSWLu2ZahQaz+i4JN3Xvhi0TUf5c5HR+4QjxkjNIMk
3j68nOCjuRiOc9nW5VAoii9SGgmJu/+uyXTZCrH8DBDUSFKpjqrWhJ2Ghd1+CX+NLczjHlXtn6tG
cT6fSfvmiGEFZJbc5TGC/Hr/WyYtvW6pgkqUA8CZDZZAl1W71MqFQYo17w+gpQ9kv5ixLzcKO9c4
5twSDnALtQM+gu7uX5OwEVR+8j4DEvSxpHAQwwlBX644Aq4ZvHSZppMVTvpYjazFlzOjF9rw8b7x
xgYoufQpjyqOf70XD8NWIjjspPwW6W+R7DOzBB4zPZ3IxJ+ahb9vZt36yC7yzLQFnpwG+5XuPb04
X1lsknELNUTNWEEFKfkBXK/Wjfqk0y4dJJtPBqBgL+3LaDLMOt/nWhoiGAfGHv1W+r/yg64u68+h
zp8guc0VF3b328Y+sD2J1DtEjPhomxZ+nJZLQLvyUA6cS0SXA08lFrrE14VZNhbVKGQxcgUbowkj
ItDUTjpp88SEgRi6O2G5JTb7RmbMJPcbkWNp5DSqbH108/yGyvyxPjdzxaeeaLpwFUj+SX70VGOE
amIBOF5kbUlF/gkFHqsQ8EVmkG6Q6hvJMAQ61g5hTCoOucx1x4Lh30fgdHXXf7uC71jDpV26KZ80
/TfyxBI4O1WA1quTjKMecw7+xe/q3qGb9UX4VuRznAOCc7JVOAFVZ0v7IHJi8CF1jfw6LcswBmoC
5Qu13V6P5XrLQyUDBZ1sTwDmZ3nC9RG0ODgb0gsJ42mVhyQhjLanAvu6kGyZFnj9zqJw19F25Dn6
S31Uqa89pgaYC/CSQ3mQKVJke5QOjwF+E7BKOlvK5PtJhDNVqGg7w2J+jOH3AoB+n9+kHm4knivv
+0ivr1fpNfsth3WiAsEoLAaXgjOs2Vg1v+KrmUb7ZFaQDMKM9aTYeZWFkV8fWK+hXx96aU4uCcCM
5qRvJiGBEgM7WtR95xpAu2qTFRcFbYdF2eX+URB8ZUbLXmtk5gdWaOaWFfKxP/RPxsPWTnpaTk0g
/2xvPgz+ZTXHTzB3xmuSNnyLX+aJfWRcgvRA60St+zVtk3oo9ZPVS2h1nYzjSsHLBB3T+U+rVNLv
wz0YTWLNoPXqoe8pmBcmPA+DKasUzrVMp73X9EUWvmyMfCpj28d437M3fSRzSiTD8sRRNECEkNBF
dpLvPSmJd9koQoOH5P2CI3UfXvmpkTG7v54GXpFlBGrNSdBbq3okvglYXv7RqKNOiQxUH9l5oVKs
bw/V4CXIxaogB6nCpRZQ6qysuYjcSfNR2jWpAKiYTC0Q2KDvcHwz1vKqioRp7/8BjodoC3md5bgH
NU4P9NEmAS/oHKJSl1N5156im6CNrl+H8ihW/bkXHLwyDAkSoYgr4tU40T2wuGWsFHLw7cuP3onm
iagAoR7BRfSKCxlTwtip2sawGiCG1om34vUV8PsPUhu7rgYOzJt4MJIPr5Is9fUKmvyiialxMG2w
lUzxlm7IO3B4efbxpkjefL81ax2AV93ZS9Zf0lvF3bNky/1T1GRimcTI1eAcDP5GSBqWomt5ablZ
pDUJ65QaCqqgChFiCisb1cSTj+iprI5b3YXbIkBkdgoOSnVaq+IOboD7Ec3lgZiX9ou+Fd9RvcaX
kG2+cBzzT3zKWigRNaoOzW5klMezkCNQdH3YnfSGG8fOzqe8QwhNMqAOcqO71/Ovte8nFy1fH/Lt
X8qwBZmCW8G2XNVB+Gco3tvkLaC2+2sgaWlCSL1Nsi3CtpIs8CeoP4N96Hje4eD8eWgX/bm/pLr5
Z1zo+1iZdFBxHu/nWaH9XO6V0hIxyQAG9FoBHes+XEmGm+R68Qn6buaTeVu2QrsFW1uiJq3BKpUD
Gh7OJ30bSoZj3O2wg00GQvNnoE/K5wAKEeBljSpxv2VURHa9TmGAr+oiEUo4QPyaseFnFs9KR661
2p0MvZvT2YjeXArXdgDzTdGwVFJRlC5RklIX7JNjgdKizsr/oM1F2RjdPrWQHGPsNlHWun0FI1Gb
Vy5yuOano9hx7wWbRZlB+1SenMU+6FDFp1WrnoEiRxQQIxfjrZHIwFjVMn/ARhCOeoZZ+wtilYqg
kHVCvl5T9UulKux2NHK+K0Ni7vZ67BVgEAZ5Dt4xUbbJNvXhQwkig2v+/Df/3Vd3NbsJdEiztLRy
ZBWYQc9s7nmLsObIpe0hZOuJOKn+ncJ1cYj1zaHuBozL90ImSGU9S16Q633MJcBG6+FLp7m75xrE
zdNNUssr6q3DyZ5SG3DCWnOsTKQHYpfNLyDg5wfgOWcu/GSAdOHS0m5TvNRs7e/o9k0N26JyAkxt
hroeXTDdPdycJo4alHo8BtMgE6v8HpOBQcj097Ywhknipijd47qpIt+/3PrFEKQTIYcFPs8prOJ7
xd88f4qovROZ8GdTonxbcKPevM1MtRdznAxykPpyNK0t9iCxfKSa+K3f2aJD7YprAp4Mf2CTpuMJ
11mUHMIIfGnWXUP+f1cRAggrMKoH7QRqlb6PNOF+EegG62xD1tZDpUSR/dslYpmnpuD2Ru0HINCZ
z0mLjSSvS6JkwgTB0BGtra70FF8kgGVfH1c5BAgKwzMQu+u7RzTil6LgSnvC4wceVWv2LJewKZfp
KvLUlr2gtuwIeRSgA2bTVJrRuaHb/WK78KMYsB3DJGh7Vjp0UapcxYmGXTEcpcWGmnCoIiahZcqi
RzEtu1rTW/5JlAGdJ7+ga1aFEfjo97CpQ8C+dQ7FceF6FZItwAEKUbcNONCyNU1AMjMC/0RPVMgV
pGEXliq5HmTv+k+mFm8dK5A6beeWkxssjfmm/XdwmZpFdfIfOopZVki8AMcQz2oGYAW5gHjEl36t
S0MaYR0LEgi9+37lzUbusV7oZkKgMeIShAEoBbyWiVijgt0X3+B2vNZdVhMPo4m2JaJFIJiJVDke
ECq7Ac75DITTTfIbe8VEln2Q/x2cfumTxY8xQxpLLlKmfQ6HeEeDRf/29lZvKy/cUh5XLR5pbdj/
0yD/YOpahF3TVKEJN8R+3urgaaD7ygjEGAQTrqavU+Q8A6YOMwNaqKPA7Fru6y6cZMA5H63GUtAP
0yZzhy0bU0zRUjBwijz3lNAsWm3nZQGmXhGXxlXQWxWqLRd4PPpA7tcfSM+BPRk/TKioljju8vgR
Do68wj0NnU8qqnVtZW0zmT4H9H2zYkecPzWzr0hmG/keixrUBGxcFLI9KYO/Sv3/IFr7ueLFPo/R
I90NIZhqQYm90YG7I7n1K15BQFCrbzWxBz1ML4NPZxYHubS4WizeP/barSrOOol07g+wsoj9Kabh
+qPhUX7FLxBzPm2vfz7ygubGyo5fXbAO3cSQ8tex0fg8C17hkg1jKR2n63/pdbJpc2ymfPNou+67
PkCdvujnWkvlftKmK+6kSqZwc0/g+dQ+G6Rux+sCAC4sUhjat0TevTkF/CtYRO1Jg1tcUnONlpGE
bqw+qANeiON5xKWBbZg0LMPZbqBujw7UW4P9u0Dn7pnpSB98YE1Hd7dOSwtoo8JLb196NGczxVaj
b0gPowRkxZxSV0b+XmDnGIolGM3X/eEm5xdn5gaRZ3MQ234v40o/mkJ6wHSb2xPIrLqL/jw8Zuns
Wz1RHl2HwLbUhnOftkYr4kOiYYDq6KZ9j10Cq0aKquh/qCq4WK6gZatPAPArKiX6ynz/uhxOlE+g
lfB+UrQgoVyFnMV9z8j7Q+/Er1RPJ3eEecvNeSxYanry59Ev/CvHnYCau8UJncFS087sXIZvj4ng
0a1kKT9NYrJKOYTb9xSyuBqrWRh1dIFCXqN79d3x42zyuhCu+FBWUEaqtfHpit6FNAXbWgDWlczx
0VSoKkn3Ju5zFXpYhRqCKhAsGcYyQQW+AuPAop2a5UG/U3DhmCmMAiohZNF8n9TncU9/0TUWkCZM
pXVr88K4p3roAd+MMV5M0y6nqhym9GL0Z4vwOd2f43pNUOMcxOuvwpXOxPkCf7hsJ6Z3vvCVF1+/
7/ffPVdyM+USpncPUsIVRG3a+U9q7HleFu9c2VlCCVNMYSPhoUmY9a4XAnq2pqcpQ2EGkBoqvp1Z
6dT0QOqZ4YvlQg+H5DuRJ/bEp6g1nIf3oyXKjDINSydMcTLF5F1/86pKpeMz36NHhxA/g9xSJUSG
+n6NmcQXIMKbuMVYbG7LRckaLGi2adcFjNqrvru0JjqxbgnSw5YwSC0j2Evp08kPbvadIKmdzIzj
v3vN+4OAedKqpX2u7M5a9n4O5mW/UCEdFFfUSPf/xetmoYqVIGUIZUzIxYyzZk6NiwNrB4v0BeBC
fPWb6Dxl9HFImtyfqaYiDUkuJWm8cvQ6V0zeDtZFeXOsQl75bEGZULJti0lQs71BQKFQ4ibtsV+T
24YVEtODuzZeA4IcrJjTu/TXVc4tlvW1goLcA0Llmt5Ne297lxTZgLD2HuGfW6SyFGc3z6P99ONQ
AccsGN9+B/28YHh6g/8QCY5vl7LeAr6YYpgs4L3g9rLCZWAMqc9vkq1oivg7roSX/4Nr/u3TNUuD
Wx88oYi/PSUt7YTKcLrhJCRER68ypPtA+PhMVdiNuhBf/Lw4TbFV+YaB74qaifEzIU63lxct/ZIv
Bc4YXEP9dBPqdOGxO7+wk+Kcd3UCoaXSe48gG5dFsYewmxgJkQ5+W+3f8DUmwjcFWXxS55LiHHM7
ME0RMAgLXJot7kYrnr6tkUreapZRvv++bXxzSdJBhMgzD4eXJb3wtYgh9E8hf0q5PViGN7+UQfUC
bDVFmZTBXz8hheEzUMl+ODx0OqySWyffGHBVLsoI1mqMXM5XpEkLe/wpFf3cmXhJYMxvhxj8vmlE
qaJ+r3AX1M4F4ohn1hIka9+q9jvc8VrMHbbi8XNlSTOcKyGzGcB/25XyFf1QBjY8aKLhFOrIPHn1
VUwYwbO3eAZ8hZ0amMSN+/f//1uCF9Ra2qHX6K5jffDLmzvQdo1mNdRjRe4M+W/Q7paIilKOLHF0
F4o8tnthcAY3tuJxeWtkM0WpWE3UfOBaXQQQcc95lrQW+V9SqD7xYs4BPy54bFug/3Q2W3wUUcwV
OQaxwmkbnXdZV7yqNKfU8IM9rBUOQRRMSD2YST51xAd2zo6zuQUlNHp4gyQC+53UQji8Epibu8yf
q1iFUWfW62FVvaM09/QGTBpFmNlfLTYsM8Wo/NzGzj9XlFInX9ei8R/nUndtDoSeWf0vb0W3yKhJ
nwNCgy7Y/RhEoCRlJxPKUqyw44oUgfByMTYQHTGoMvoUj8kboEXWqJbyneGHHxhC3zXBWo0lBfTo
tfhMrSlE1+BuY1EbdlVoQnMWofhudgGI3lSUjkZC0swHQhBc5cNpkS3vVDiDrq8HnSr4P+uFZBoH
zdOxQDEg00tJpxLvMrExXgkvFn0VdYibLKvNpfUmwtTWgdCxh/OzZ5Bb6R+o//oLRKngJysNhhPI
QalNhrJEupoRWMoX6MTOzUmqhjNnEeZl8NO2joBgyWn3uPM/1EAHZRl5DLEOqThoy/AOXjWuRKrR
sRybeIlNYnpZC0IAaetOMHD9P4YpN4vrzW0Is23Zo7Ie6vlKYYyouuZntmIe83T38M+NlLw0irCh
CS6cQ45gLrGujLjRn+k8P8R7BV6WZF/UduWUuIlKIrxkWiUOfFn89JUkL0CR5wkkmJ8v1p9vL6gy
q2Z9po5wAQbIZZR5r+Y5TRhqyB8Bx2IUwaBsuKg5eDarEPaLYT4DT0gfMkCscQXB0MNWDvtSsnzS
VSTznw+6c8oTjcmwkSAOFCiffFbZ1Tqi/STBkTNnviye+R/ONNeYWgjSSxNwGgE21t1bbWJ/6/L7
eKMkc3s3bKPoCsAcv7girr0a+DA8vCjCXDkBOgq1LgcnGsHjb4biFmT3auJGgVxIgHUxHkiAqaUi
/Iv6CR1BW6nDpMpWyA9jiH1uSu7abCgNyaB8eBYQYyVamj/k3lHDKgHTuoQ7eC2Ry0N+pS2gBFLN
d/YtytAIByH1s6+OohuESofSHS8JEPKEAWjdJ+CXGoTiDXgGTyoQ0VIwM6vosVPyn6KQIqsgh+Md
vq+r/6NLOTuO7N0duWBqi9y6/7F0Txmtr2ajJzJjsWH2R7NeedNP3qHnTJxbK+xLKL9b84614D8M
qleIUNs2zPmUK3CHPjgxugO+x9L0fXI37y2zVrd72ATp7Uxe4D5ViUlUsweJXVxzwuUceqBUKZh2
5aEAW9wETH92daEeZMDCuhszjhRO2VXtVTqz0kEmy48VzGWYwNX+TKSK4/vMfiOOSv5Zag7yIynY
zALeir/U6qRvhcXjEvPEQxpoObmzF0yaRK1BrlqYfXQM+kiPSIQrmS62IunleHPJPXaP8tETANfP
GLzHicw2lgFyWFVhgqsI+iw9lFFDxZjHXLSG9u4P7vSSKy4j9feZgyPfKwdURjoiKTn9CzDN3SZH
dz2QQVlFl6MyHioS1EfvSOOEjM9I0ZFFIxyHjt9oj+p2Fnp87/Fj/4JEnc698jRiczSKqOkEs+Aa
JjbZHuJgo01/4Q4f0PmM39pkxa8tWBWD+1dubsjbe/pzBf2VWWkaOLSDEYUJDpY+zO781u4m0Rp+
uMspbc1jNR6Sz27m8S7kiSZ0O5YIXVeFi02upjjKftDphJP7iqXDCfcF2QHf+yM58TQ+zdWGt9EU
qGtY9vz7c5/OlhA/qPtqV5zYHQHA6C+t5rCYOwDWJSWsD0EQgndRwqe3o7eYroL1Lt486hk4a++F
1M/1f8uehXDb19YHWAebQthzKudifx4EhtFYQ+nELSbFJDBMM/WE4qjc/YZ/ogZJRsM2oD1tSIn3
gq8w+cpJtczNSTWkzvY5Z1elBCB2y5adcw/r3oPQGQLDBJO1Xx0YHVRsZaZvJSbI0o27igGZ4uDU
a3rTe8IagiATkEwE3O0W0pCvbhpZ2LzGveRRJ9fRV3+umTtV4nn/wtJFBHHmnZYmf1CtaIbuhSI+
ekTrkaXZJFQuUoVw5e/qyHXpldde25HZzlIoML9DIna1HxCqQgiYju/Scc6KX1fE5rhgHr8guGF1
8J9FP19bGlrofHm8oVvw6bUTg2aP6VHDcLbMXf3lh3hYQbrRpxOLgdI4/xLNVpP83dg1DDmLMp9I
frXoMxpjMAkZV9sawzTgjIRkjB9Fsd4QbzJ+LDB70G6jReZF9jKMt2oa921KQW7MS8tr3Xp0f6AW
Qy8TNcMxnnI+lY2I1g0mnNVSINo1Vqj3Ci10dGPFyrN7xqSQYj4LNaj70pAsWMLSbaqtUv8bHXR2
TiuXOqT87/Zhas4Rl/KrPCJceAnTBcQQZKfAiHfeAWTawbCTmbHzkkWXw6hQYiPxbIXH33viSmV8
yDIW5y6h6+HZNRoOmnjFoNDQcR6fH/vPIjUzsJgBvkZ0ucC1TEOl3RS61O9PnzYP1y6zhPNUl0lv
2zZ/IX7Rxy/w89mvN1x+OJRVCygqxJRc+zZcyTas8o8Y8TaP78S0Dyew6HQtYdWzZj52tIgUXByy
s/w95o/tUoYSTjLeWgmgHXo7dgFqtl6jjq35W8qRw8GoADpx0wjwzMIhtILP0e3qEXwa2aEIpkct
YZQjcHZGtwIfJCxQn53toCdjsi/k3nuJFHZl9ZsYdZjFhljgbDwsnTR0g/B8yPwEyc0+jZXatNz0
AIycdPGIeYrlvdnY+8BdbHR0BBTomW/owJvjOtH84RDaIDKnczcA3aVjay70RcuRi7Ziwsw3WjxS
tsWbaUZk4SE+3fbuj3V32bCpt6ICh3X17K1WszNLFpOJaKY6wfzPMH33CaGYckzJnvswtX7EcMJv
0fOz0qQQfbvuHAMeKMFMW2uqRqNc/VUIcluaAfnlwacKRch55GHPaJriZQw1KP76KvpZlOXIMv0f
Qid1ZjZ5imltVrdvduLH8L8M93LBvrmIG5RmHqtv4Q5etWd1m4tTHoCrUcRVT95K0e93H25wCEby
Gml1uMr27Rg0poD6GkzQacQFRBWMfbiicggz6iyAhHYm4e/WFyenHdRdR4jpO3Vb/fPbMLrDh65E
xIB4awD+MvC0977onI8Ov8/hboS7WlGA47AqbNOpEjjVer7Hg/+zqq4/CO79GIP1Bz+JjcmoYvbr
2vj8ksM7LtvocavKfe8lISq3Yb0aESlc6K1h1GZ6afPGZsuj+hf56cz/RRDVkRYJQ/k2l0CJ7Zb7
jXiwhtn5MmOOl3MQdomT2Kx8HFoUmm7SHdUasV2FNAXKQ8NSAPtTmCRcgYXVrb9Z2IUs080BxDII
+58hoHvRpHCZRxguuqhbqjWJwtYZqrgy6AdSLYTiNobd45eQPCCSeglt2UbTJs1uTsevorWWhzEC
s/57tFGLjA6R69za1BploN4Pn4wCuVR10ywpDKzM4ypGED1ZKoOjMSQe54xrQM22LmbsjjPZnWwr
Dbp6y242Hh6I4csgs7tqPFwpVL3V890HfzWVUG5AIp/3eLBp6K0vlMD2bWApX2mxNfSSB60aGkDa
0qxn/Zf/osZHPqygWLAxDL3adLuLU/6VNtcDUyor13+uWRO7Qvd1DB9FuX/eIjooFEBFVn8Ba+mm
aoVTJ6XSXMVpoDm1nxmAeIrPKM5YAgJPwv2xWJTrplix1BXUjwaIs7acDAtpZyCNWfnZ8anp2Y/X
KPYKV/fkopKWarTBVG+1OpvyerCQ+shu7YE/PYCyANaHwBRH/rTz8L4UKWKjbXlvE6JtBqwTnRj6
AgeSWPaSGg5JG/fyW+CRm/Tv5lZ4E5M1ZC4wtRXs2fFQTV/6B9DYGbDkxNnhXaiNX+8N5KymqWEF
Xowm2PIirmWz2qf98LvEdNXudUesytZAnTfidPx0AfMH1vqzF4TVS66BzsB5+Ebc/Gl7eaV1+dlY
gEyHD2fEWqgoOg2oNfN+ginYZyhPVAoAwKM4f+/3G2jJIf9EaoAcyr/emmWP6n1XtG5rW+QjRX7j
G5hI9fAQYoBtvgib19mqooHhFLYRzFIlsjC3FS3OriNuR7lY9gadSTM8wlgn360sQ3I0SeKrAvz5
uUHQInX+LnW0RM1tYpJcuNi0w6rQ6aSh1qhBnb2JOL2L54uZFPSDyPraCMR6d3jZDoz9H05Lb4KX
+iTIjZOM73XbET5i5MXIC8t2wJPepYOMwLxkHugiLLCwqhd8NwuBcsXbg3t9iO6vtG6fnCu9jyyW
YnF2ND6kTN5rbMxbWte8V3r2lkzyfmRhVd8gQFo+o6Te0b5nFCFvEkZcRkuaRHie+/BUPTNIreKd
4ssf6qH7kuH3u+Q6AU/iOp3vJp179/Rug4H5hmP6zN9W8yeQ/hWYuCUObqXjAwSEroJTggOvK75F
nvzhdSxXo4coyGzUWJOb8q3ozMpzftJbVPmKAFQ1IFQbv8eSxSvSlO7aLXPtKNOM5cUbar+9Hixm
fXGYJsQPaMbqD7WZYxaL76svBgbyGTLGTEWZpvqreXyiH5TYVAj42KuKgwLFbv9Fjc4RfgWYMSA2
51XwISzaOq9Jj0IJ2OHRGTKE1lp53t3cYriC3eXS07m547CjtswwVZCP7KVU0gqTYruwyGKVwsOH
MVc/tGRgo3KMW2Di8uj4tErIXF0Uy3jPVgFa2nUfx0Bs9KS0dfPO8mZTmJDDstywJ8kIN1JXMV29
eVjnEWDoMcC2tvgz2olVB24cFXmXcXobWBnrATjsTvOVO6o1WltlWuE01LHX++EVbTvobWbTpyL2
g1XrdeTPnMPbsY+/il8CghlskRgsPjOIaiCYdJkbtJ6WCqvFTxtqYeFgXLZ0GMpZ+oPxcPzuIdQ8
zPi2YSLtvhSQ1xh19vpm9JpUDBcDRliMfYzg+ubTuEiw4ytjNHDXruLJ7I5CXhERothLTaB8avzy
ZaxlKGEXV+lvaDJVk4Hp4r4RcVwBZJ84A2XMA3xlu/1R1tsdwGSX5g6yFO4nfdTg95bbve0+4Y1B
12iIZFAAWfkhqsYYbf399Xk+Gex/uRGuZSiSn2mpWDMarSGQn7PM/K1vIj5CbqRVkPZHYPAIk43R
zUEjNbMRCRoDPm3iuTO0kvvpLE6B4S1KaX4+qywvnN9NHcTBdE2N3/DlI/Du1TPlcMOd7XGHUoEE
8q8qNjK5vsiEKZwHPEtrWHUp3pbbTNlWAkASHhT0bC79tmYhFKOd1dmBTrZoLHUZSHZScJFhEPY5
ym2MLTTka0T134yd8ugSv1URgXjd163CFVjHDnASEWxrUHG4apDraw+PkS95OMOMHI2x7kfAqZsv
OKYeWh1+/29Lc9QCsPkSXex6eVPVkUlXjyFN45B0kKLPPclvqlMtK3kj1gmEhc9dChMkMkZEhIF8
JDUG6c8K3Fgo8I+jvk80PKIAhMcrMb81r7npAASRAi8b6+p5UhZ7N7gTiLDGIE4ke8xUwjJq3LCu
C+atSMI/GpECykWbR/pKs4qhQhC7KJzwqlTXZrBOOrZZ9KJNPr1WktwXx4+4yCNK29swF3LRqdWt
IHMjd4jbtY/6kRN2HbIYF6VQkvejxbm5iI+00i4LGDzzqPjrrgNQ8DMtoLACTDRwxdbe1eZI6PkY
uteXQMlzc3ReAudwqvsjQ2OnOWOFvlg3I1cldg6MxZgHPgNN83hEWN1Ub05p9DiXg/MPCTDV5vOF
VLjLDPaeOqY7HzfgB7jUOM3NH2cYmV+v18bgSoH7TUjRasZxsUHizVhza5P9J1mRxtWairqk5/f2
yGCh5GJtMUVe5rj0Vrtu36YV0bPKOjB38pKZ4fN7Y4L8K76zmz7+fZLNEu95yXnaaaBOldU5DYF9
fEoa/H84ltiYghLvVQwtdk/mKKVUZtcVitCuVFcNnc+0zvf0uAxPMDhbK2TWH8qvg5YNtHI5YpxR
NQckK8mdeR6IvH3RpUROElRMt+bpnjfJsLY5Jk40kTbo0QhwoBiq/UoHb20ITljiQ+nJ8gv8VDzJ
GhS6g2jmMKz66CdqgVBLXCcae9fJO93b7iUajpvjC2DCX2gp3hrSBO8pHFWCS7dyQGxyd0vzD0Vc
aMHMZT0SrPISNsSJFiz+4SB8E0/pa9VS/nOmnN2LbmKLXO0130VQIZlTwNmJgwuRlh01vJd7/5+D
dKYkuzIli3oxxrxpuOhgAOSwQq6rdo7ZNaWawPEpSgA33kxzn15s+bqlzDQEEblkNVOKv4546xHU
MnbTd9lVN2e2MdykBemkZrJsVzoyyE8owlAr7+/tg4zpYQu1FnjL0qr3xEHMzwrlzAmQMXZVmIU9
G90nctjRx++1WOZcmZMyq7Bk7Dr0/iXfwmrIdg73sGWV+2tLvENrzgKKpSEQczxt8td1eeL+3Jz7
J4CMxImEOP3S3ZvY59c8qUXJ3rQTsX/F4nzTG7HIAFTFlO3a51Tg6gNu028qR2DYHzcZqo/A3qp3
jtGZGlUYMMdljawA3s2jNz630n6+ERka/ofNBme6gCXCw64I9PnqVE68FuJz7ytbMjmLRM5tcpvJ
wxueHzRAVDMmhdyAk3aijPgYcWrNtIhyOpXjw97LXRujh5P/jwp8z6KQtGr0kf6/DUeRDbIK7iie
MxHB8nex/oTboWhNEiCQBn9WZZN2xv8jd+/IyGGlH9oyOzWJ0fwVR50sr9kgyH4mEttVwYQ2Ljh9
u39y9GzJ1bLtyTvnBbSyJl11IV7+xbJ9a9TzeT95gjBBRrMKN9uEmjn9GnoggK37t8ZdDfQ6o+dS
NZGNkrqhdW8RQ2eO5k72HamQrziEFZtwN04kFO4AFVUiU1xYiasg8oAzRP6yz6A0QQQhbkZGmflE
WNfYrSYVX/KaoxClcyDlK62l3ewn1Kt+iBsxnkV1b24kZnQxobM/jyfvd98GoU5Zl+EHzLWNrQS1
rZLcNpeNHFKw2EyQ0QJjwsh0U3QXPuq4TXd82vgaNtjTrx0Y9gunrOtKmblPsm9t1n4pie4iSKqt
fjHOwOKS32twneivR3uJIP7nhDGHujoLfhbiNvCoxsf1VEHtRfJqr87qJXSZ0+edkRKBL53cFPop
StJVYCujJFhhurIke1z/pIXQz8bBJgsySJ42ri6/tqL2w+SRxM67BMxRDpj9XGAils2pdMIdN1ND
gG+mE56mSuaAUZM3KXCr6UN0phNsALs1NqpU7rnak8FzekfeFgXrjDBIiX1YpSF22CSrCvAR4s7k
NnAQMJrA/FWCi0QDprQ1xuOWIIId5eSSAdId5uDneghFE4s7YZ3I4K+nlQneHpeisjll3ePDlmxM
0O8rQLagCJSsS30uclKUwbnu1SyTrct2jRs/uHGskhXRYeCRwVoVQKMY90UfzMHxAUJT6LgvRRV4
opDMR+9Vm9bnp7ccw1NIGUPYIs5P2FUIN78y7OsVROFGSDxLHMHuVomLOfSFQf54j30DPgmu6kxR
1z4W9DlTF7l6kT2w+aUgB98udJV8WZ0yFh0RbrcVIDfOZRe2fcIR9CPBP3FrCTMGaUvBJketQFAp
S8+d6sIWwlCCCTQdX6IUnD/NdJLJjZssFnVSX84CPzNfsuC9MKVqo8Hlf5dE199o/ZN/rZH+J54g
rZsYLWUpfktMOCqVadjWFVCWGpd+7A/1PMX8z2OfouV53UDkg1OnSCPNo11OiHzUdcN3hMfLCoDF
cI9HkyIsLHNUGGgAQsEIRZGL6RWwCwYi7z4D4yK+8gQEAqjO1e/pyRfer3Pq/7Gi6uo8LT1qo25T
2ldSUr9SJqj83l4Ym2UBaiBZji3G3jHprHUUZZ09QhSvpN2OaTeixoO1O5zyZu52lcHoTwQhy88B
Xp/PxroItgHaXg6LT6OjQv5o/ZpFaljZMiCocGC0nI5vvcTxW90plzeGp4JVRa6oCrdbN1FVSdl9
PM4xivFU6U1bdSJSTdbtkODyM+svxCK9gtaL+sJnLn4DTzTqLfgbTVlYEboCdWF1Na/k9DA2vF4g
eg8oU0QbB+uT15laixVMuSgIQosu51dfg76ejpCAUzZwpMNQPTrhCI7H1vmKkhJJyF9yKVkNE9U0
bPmGEAKDfFaKmqwnBkRF/59wIL3610R6bp62wpHTE5ifOjGxsfqZqPVf2474W4+rj9yl6ldvXjoW
Guxd5o+p06U+GMhasCoi0gT55y1fjQuzyoiBXnHObMztavEJ8OwZ4/Zl79258n5/HqWFHbzWC936
HcjxIZtRD77vt/lEPIb+zUMEqcIsKiJSvT8F+8TsEEpA79YBFx4uGlKfxVBozWJejjm5+yMMq4jn
69IL0TpDiFHk4iqlkalfSeSXhrrjBU/NTAMIMF6TIu2L7ppXPMHcYfYVXRKLZjrgPg6H4VQNujV8
KFRPkL0AH9ltKsyeE3OyKxnDmcio+EAZxmXyQxNf/4EpcR5E54iMfWMG3jrlXkpOvuMAlnlNGoMf
K/Ur9SASRJUSFApp3AzIt7sj1QSyxC3Y6ZiHb6mlusyqE3I3def/pPh6R0N10gVTR7aRXi7/yWhz
6hXRwtdEU7sFrhpvnr89vNECn82p9zNc2sSdjAAFxP4DVEFmDN0ogoCv9XUvraILTO6kQndRnHUi
L7N+927UtGbzDXwDdsYHtlT4YhI3KdSDfqmh1xG+ki5lEak5vxf0U1D3a7eqLPZc2GAzRFI4wia9
JZYUERrpph/Ok9pzgij4La0jY0IAeJMxBaX2ABEAGWo6YixiYmkZA5hg3TVJXsFHOIvHofO6WG82
JN5vj2NYVHADOHjcyckpjX0B6i5lRcF/t0bCNtvyujfbhuvVB0JDubdqT7pGlZEWk56BixneB9Sl
DUKO2HkrpYW8DHc3yABn9l5NPXbpy+22KO8+fyp+6WCOiY8smPrBXuA/9FflgWqAQYfctkWdF0b5
L0oyt1s2yECtQ1M1W/64KaS241EZ8s5OVxxIJdpO49vaencJGVwQqkJl56GLnn0Nj5Bpp+MVBlEo
wKBbGRFHrF19+2YE0L/+/iqooSxgceMA0cDcv3h5TihLCBRUkuOYcKTnkrPJisvcKjvKWbSeidnX
0idelIolDBBYunSUdp1DKQoynWQvVWBi2tpOr5K2tKMRxb3Zmr+LEB7kwlPziG09HBKnZll2+2Rl
ul1Q6UDteJHpVB/TPx6cgtgc8IT60b0/60oPiN9P2pJGzfryoYe+6kaIOPb5OjIOlhg/51VnrJp9
HbFMWWu0x8v9ke0j3DbIdMCt7S6kUwTvvAtHifI3GR2vChq8C7gtgl8p42QcbjmbayK109pTc+oA
JVePn1HOXUH0UteEhexs/1E+hoJWFiXkhIQTjELAbpqP8SCDljQxkaQk9CW66SXaiQe7LddHzset
vFr4617KeviNeqK3ZvMSjH+yxEuP16cncHTAj47XQb4zjTHTSHKaLPxTKS0l1ZvS7efkX9MxcW7w
GH09q90KLhMWWvd4LkJuB7OIPj8Hd/pCB7vhTTb6ZFog6Qt0qmbs+ybfHMF5USxZH5K1MYkNOb1t
fjUTzYIw11ZSt4ycdSaQnsgd/ryUsTfR1Eqf0X44zVCnABblDSJbTfnvRLPGLqYUimxPCFpTXYpQ
4Rm5T7wSWmwOMaaeB8g7E4O1pCSv2q8GjTQXJblJLSBCor1cTn4Km9hTPBCDvgjHqL1yb3j0VI/d
z82WS3Ae8ZwnXj7jDbriyh765tk9MSuZ3LGdCh1p2jR5oyIKFwnB09s4+4MRFP2FY1l7f7Z/sFH6
cOkTbS+T9o0meXMfHezVqaKPEoN2TkiN1RcwVqLbStX+89Zvoe7ZSOmG8fs4iCEZVVO/x/bA789k
UVvdeMXaCsrlpw5SkYhHAW+cbJ5kl5VAxrQyMcYcV05/LtIhdLgrCYLvh9efbbaZqdFMRXJwvHjj
K0AYctY7YBSRq/ZhvlpcmDvRs3la4Q4yzo7MwehuQyjGZA5yRElSajL+CNM4T16qdH3tfFZ1yEFK
/fRAr7B2tAVyRK+fXXiyBBDm0JFQdd7VGfiqk/PJHwJFUn4WtWqPQhkhUvEAMSOsgdY14OcYPTns
JcCz3Wq9DV9s0odLR0C6hd+JsrtcHVbP/FqFBhnxiCUqisSpHyMx3/TXTojbSMsdAvapXZ1YcoAu
yL5RlAPnXBz/WRWXte5fEnrGkmlLCLOyuAxm5/JHpmcwj/zMJvT8/isxzjmcE1Vk9/WarQVBP8hN
/53CbYIAriSU5/qYv2mwnbTnvEtHBWQsjHd/L66ZwCt0PKE4l807mY8SzpWWOj5war5q01T7kCsY
szUs+9aq1vT3akVMT/b9fOTLB5HwePzgiipB3oBYYhvoEKnVip7gMGzVF/J7tFsdQo2K+fkQhu5Y
LuUpZb4fRdglvYZNYfqKmhz4Wh7ilLZ81uflh3gTmM1GvGeXHUU5HZyxAJZIC9tD97jjuM75GpUk
3vacLgzPGea5WAkRAxewK8VSL6f4jea75QDlSgX73ojc7QgLTylQPOsLoAz9uHUxOwSKQ3SKwStm
KxnXpbZROr4r/g6S/UlG7SK5H41vwrTx1hqCXO3nJOVVDhgKgHGvUbmEVyiYn/WIWAMqFjueRgCd
Ry/SzycquhQoA0sNq4CcnhNEx+9Mv8QpYyen3UI5+O9+Pf31/psXe6WlzsgSZ5VTQOwmXIt5B3sY
4/iqojwlUCPXzrJUO3Ad5jxurI8rKPfvieYSFvRRaEHfjo9B9HArjDoMfieNutmsbYQ7a7YlNcad
8fAjVEjLVfFT/6afG8uua4ZfC3JZgkByB0QqBP+96R239DHgkaekn7LQOpRXdxz2p0F6gfwIpBKH
PCmah6Sypf7tpc2dFRdAOLEwuRDh+wFfRcUAOAjNTV/lMAEFKZOcNnGcfOQTB00BEN9txfVramFR
5WUMN0+Hw7yiatpTSFPmim0WpfcOh53bVQFNGEgt59+1shrKmwTrXU2/buHQLTirXldKmvoDYdAz
PUG3sDvrLjLvXzU+x+tq99V7oSk3ZUlbEST5P7c3wJmQ8MNZLyss5SaKI9C0KfJWE5Is4Wd3QtAK
xQGWmNEN1A7WhOXQmmgFkgK1ntxavvAaInT5roTHL7yfdP7Y0Q+PulAe9xG77aJK3HL+BfFOBeMr
mgNoARpnzT7+e2gkYRSUtPJVPpqGv1L2lIdJ89pSPqM1U7XV2H/6Vl1z5A5ZEvg3TvMQ8x3LEk9K
FwnaCbBrXESxk3OawuJisWYrAks4pQHVrHbuJdAACTSf8yCWjz9cxJTjGAVKtOXxwiHmuLBkNYP0
CxFNs/OgbIJgFbNS/AVYnaC97E5KpMrCf8tw70X9oyG1iCilp4YGGdZrSJk11Bk1fNDgN5OjaUtA
mgAzxT8DsCl+Yu4vDyZjPf5w6mfsNL+4NSwh+sQSGon0SlYBKOdWqfnne9JZvTapqWJLtvaC9Fio
PD+TFW/bwgBj+tIP5yWNA9KeFrI1L0GePKbAEiPXIoyR9R/prIeasnluyHLvgRbeaaaLuh662h7P
55xogLBHg6aINdB3znBnko0ZOAInMm88n69ge/2eRldLuIDdRaxtDOULhc4q0hTnYQCBVHpbpsU2
wMcaILn9KKXgT0TlkS7GtAxOrRZvx8nHrZCvTjGwtYxLA7cYU9P+cNH2nceqW65o7uVx9ZIy7TpK
ofsaQ6FzrWHxoMd3VYlWRUtj3Txweztih5u+KEyJ+aEbNUv18mPYLQzvKoNsSl89NTH19YCvLTkS
bcubgygLEWvJdohij6LZ3u6VAz34KLAgBWV5Fy3MGFnzZU29biQGeYhHdVyp9AOw0XZeowB8Ikt2
qKQk1JQQx8qwce7aXFf9qaZccA0X1oHifDowz6rfrN60plmasX4NKUzuxlIprvHZM2lhJabgFcq2
F7TwFddLCRv/8EQOOVu0cio64AznnT5Sv/ddmdYkacMB2uoHX5x1kLoTl3kZdhQktfGgSPKLTS0L
UioB45VJK5JAJlXHrO2HV3ACCOb0dwNa2nAva3XrSfIVPZKXm9joX7wv1AVtcX0dYfS+zRuUyd53
pjQkS7SDxuOsEn0jLoh4qQcHrgoZv1OI4Sdf/b6zfxX0OMjvfWvi8Ck9pObUx6C//pBlVMddEHLh
5gbNdV1XF7B4JgxbnSZUqCKdvfCmrBIA5XtMMjXeGhWS7mrUSJYNIb3figC7fDCM8j3yqA/6aJt4
6pzNU3xqtgVvQ/g5JaV9FB+Foztn28emMV63F3Xca5CgdemcT9PlhrX3Ip7OiwmdQ4/nny8PF9b/
i+uFmGblgBxO9sOLUVUNVZ01OJYHF+G0DWjLcAnOGyaE357mHxTSNy2Nxcg0T9LN8DCz2nyShvla
0fbZjMRLF2cFaQY+bRMujJdLlWVCL3HhFZg6LzNA7v1eiYKBogRvfey4FJtdjFRxhYNcrgJy1WLq
AjPoeFzCHVJ9yIdXewkHqKCiOrV/2S8gu1j7EwNyjnINI8Bw5EDtpsXIcpZniTaD3ZkG1k0ZY2Fd
bOyUp/SJYJ2zykPIzDP9nj+K8XuDzelFix84uQr9olldyQs5FkLK1IEwq5EXygt7udSIQ1s7ck8E
OaIk8oYZciLgx+/AjZjpzwVriKLpYV1EYThwuUHa1W89vgUA9NFxzr0KY/dLT4IjnZL807k+vnCR
SV4B0ZIcKXwJMt89iP1QavCtZzkWtCYlVL/B3pOsUpCZ2U5YRzEj3PEIvbUTf7E24FGutgnklrVP
Hswx0mlMBYrfPW+FHphS7vKrllla7/huUUB5luFwWUCvJikK5T93AI5oFP0DpsGjLy/vLLQMTaeK
u+BagqtsGxJBy1lughPWZHDK7+7Dms3NUaPSdvWXT8RLldtenTRubeE4ffla+oGE/6BO/r0KKs3w
LpBobYkvW6gwEIKcrfd8SJCfCZVgRFbpBEvfg3PhnYmRjUAa0gKMS7Ijtw7kW0CFYC9P7f24DlHz
rV4olwWFhb/5rok69AgSdU+79qp6P3laoBwEExgYs3jiLmocJ2lV27jjXs8ZslQz7JKmUWqbve3q
2b41Q3IVd4dgM7edCUFmWN4AOo2FaAQ9UTdsNB9L05Rmzo9lYqAjLhrczi/7Y2XoVgUQTXuuJjG+
hUibCVd2DPBFepdW0F041a0wEeTQoANLeeCaybOiGASo6xXxNXw7Tfp1o6mmjjubaLCvIz6Pa7k/
1aijUDjYVINXFi0viIvRh2+cFmqVG902TwuLQOJ6yQHntKWhxEcq0FZt0w5yBCiWehD4X6wz+ej4
l+19zplhuGY7ScjUJaXCKLk4wMgtsAy3GQ4leq962SphvN6iw0Eu9KYob2vCZVvKaEfNXJeIfKtr
RQDJAga9dcWvOXA81+Rq6qZwVC+YDPJvI8sPyJOqLpVOTsD0knmQ5tqhzt4uonrZmpza9+RmntUl
Y4zCrO0zpXH4zHPWepo2ku7md5jpjkTP09LUd5q/rVCMy9QoMrtOJe9vHvbgRe+nYyg+unCeHhsT
fcMiThr1ad6LnJ9STayumCYB6/zh7fx+QIa4bIaDpbA9L8WYC0Z2QY2H44IEzKbjiutdpBoo/+po
PWmbKOgH2+g6SuguuHX0mloYEacg/lBUg6thTAT5OdlRWn0k5e8nf9/1R1L7n8h02NwWRhyZKmSu
j6HuhsZKPZDLoVZLy+5VwNoZZ3t+Buefl3frCwESTo3vsT1hm+HXX+pE7oZVV30FYcjSwaZbTJp6
BZP2c67rfBXb3riDsqWJMJagmhiOHsoMQm8Ta9Nm7a3HxOgYfA+uAL5BPKTcVGN+8pjULMTIpuqr
TVFKFY2YZGWSXdZQhuWbgHa4KhAGnX+HELVRxbLg+RG1fO6mdDv3xdaKfSfC9dOnO5BWavLWBdVa
k06uf594mMaq+l9Rp8Rwy+YUR0W4hrMVTRKN3PNWnUNSzICBLa2R2+wSWWvoQty70hzFA7BIPwIN
BufL4mXa/u6n4iimKKlyiKtElMumVuYPHCx3J2m6NVDZAvr/RcUxS2e96gXor+LwBae1L1kC6bkP
hsXfpYA2BDS1hQhT460f1mQgpsHG2Z7ED9kHR0t1m+L/lQ8e/jty5va/LExEwKhPD4cSZCHqPZCx
SuzgS6+WotaWeQi86+BFz3/cEWXuTX/2Oc0q65LvXz5E5cZ1nWvGLBnYzP3IdrM6X12yHAcTeowR
zuFd1neuVvehfmBR5rYn1PhrjnvI+7Lze1tb76zvS822vu9PKQAxOWhS1OmKMk/c4xjPUmqitMxc
a2OMCF8Sro81Otb99wkK52T9mV47t1fxShhda29lBGe+EYFx0yQBvLMfWI/qBvlbq8nddWVfXE96
8obW5jbBoaAnjvJ+1hXCYZMirLayeOzcN+cUDt4hi6gemo4TC2FpoM38lQL872pl9TKZ1jpipCOg
uZOlMNOJenPON4rJiVPcdCchjDXe3HsJXMhCeD93eygBNUl9WRCWDpk8r6OataMHxs/1HQ7RC8dj
CPd//DHI23Hx/lQLCzBuz2h0cXNevuAxhDRQNqhIlWcRVMzS/zJrHRc3QbYXFMosFd3GHlmUL9wQ
7pe8maJxC0huWa9fMRwH54F6bOx/eQfuuH0fVIlzD44qADiLH6GBzJGdW/M2H0Ta3YbDcQchpNUz
XEM9EgiBhYomuB7Ys9bFbFeXQEmiBGdFy0ezbDDVgU230xCaiRbVwduwIky2SMySPrNBUDzeg0wi
/fchkuhC4MyXtud4SA5JcfkgR6ykmcyNkEA3OgoOyTwhnYkdH0jtqs7IvftfaBpe4QxmXpCUNcn0
1PbDEB7MyBQXqorDVzUSTRghROf0rfoUKzzXREyGaSBwl9s8OjQOc11gSlua84dp68Ogr0VEdLZg
uwcRnnc3OYw+MfYKEpMUviQ/gBpsMK5WIDp6oGzLnVq+sRJ9jPVseqp2+TpfEGsCgl4v/pVYceJh
2A6E5o9xGVk6axteIvaFAFcMl3xF+JEd6ESzN9HbwE0xpUSSLBL2Fhrzd3c6FhrtT0UfWqetZ8/W
GzdtjP6ZjfenkvLnkS4KFgYzs5rFJ5Teb+9SjcmUYUaDIB6pnZhOKINqAfvVgsK8HawC1YRNeXYI
FOT+9hRKFKtCEpiqh8IXzum6LXlQauJ3z9B2nYEwHSe0VKM1/NAkNZ8dzAXQxwTzGqaBY7uMAHao
OowBj9D2T9qvUTaRd57BTrE7xn0UfMKE5BjDvIbSfC3Iq+U9d4NTSR2KMNPouSA7XTXu7sMH4I/z
Gx7AenRsOE/yLHsRIwfPSE65DnV6prhrT0y42G1od1vnrOGDLUXpAH2pXrIERnWM0T02noJNZ/SI
NCquhGzMBwghZHU00ASJmVCShf+i/MvIUExftJpS+vjEsgt0rzJc4ot0vCQo+dk34cXltb5MYnkj
XTNZ1KJ9V05EYAlur6FTyR4SiWe0MFdVwz7+cKpFgyHtySnrvDVTT8sy/HPqc5elZf4OCWRIEDRX
afDyN5pGQLVAvgkM3/rHzLbAMuLpFNFDVFNhdqBbKCh0TJ83kcqXfoF8TIvQqb+6Jby0tGseWKP0
Fe9+aX5eC1LbY/+1AzKQsl4iNxsR0ggU9vo4Tde3ZzpaPjii4BGQ2gdUaS3Jk1rJ6aFHzZRlaqg+
JkA2AaX0U+ctoxLdqXbVADnv2YMg9LMPolPv57rmCg75IUlKRz1vo0MGI0Mj+6+gr/A56+rc/U5I
+Q7IGjvfDoN2gKSsx4rql3Rp3bJIknjNR8TPxdCRaWFcKDINQbFRWaH7mvekFLMVvNT5f2B/iQ9y
kVFnG3lFIRqJuzdBoL9MrM/DBNYioI0JIJbEZzBKoppjOhVH4LzRUMlZ6V750TYo1gmXour+WYYN
QmTlP/N2ZI15pb++LGBTSLvtrj/jbn1E0ZqSRuFl2uFYrz1L3WuybPuSvjXWiF7aX6clUax1bTdF
NqE09UhnUOTDd+58QeHIpDIwXO+yt0PthqidMACgP+tGCMU43sfeLpW2Y7QKUSCgPgykhvz/40nA
3MydWtKYQ3LmweG0ZIHFupLM37YQgkAipLhb6m+RNJpRt0557F6rkHtOO/ZwbB/V2XI7bhHomNJ8
FREt1uZkZ2AFvEuQLwLHXmggomb+1ATaL844nnF8LFnCKah/Hr/4oKvQY30rmgknXRZqz/nGienb
rxMmiGGRlXq+vpX0N+63ryAa0IZiMSVvuPB1BvA6vtMadqLSxI6XaTJza2yzIS2Gt/sHFybgbU0g
fNFGkJnbUDWIq1zoBgh1zWeUOvPKtEvZJtLb3RqqTywwGVJcl0aPZhPlVpuSznwDZX+tqlUkleDx
0NNJhMdaE/9+kw1IWdHh0LTjZLX2cjbbKoU/Dalda2FkzraIDjW2RqyfXJnywQUQxtfOZqZ5EWrj
Ui7oOm8oFkzGovA40fmwX/CdJFrreQYtLIAytEt4ejyD+5bLAlgeWzFYwE++yCo4ZNx0IJZIQwU3
SGpwhgxJ8NIWTZm6ECL8oscMnLiFRnV8VXXs+gP+kHnpVXqQzz1PEotVJGinnlFNlnKCeq2Yl3Ml
ITa87l668txfWY3ekNTgjJNjn35qS+t6ktQULe1pymzO0qnGXkCdhpgAqKR9gehjsvunE3BHTGse
VT44o16bS7ZCLNdvjiqxXVdzIRPdoZZ5prJqzLJoioTmxs6e2AWHCYxeusPbIo2Ne+vkg53h4TGj
MG3fIVM1J3p+IWCjxVCCxoCoNQA2KNZtfJiANUHuOpX0CEEpehBbswQUMFqGkcw8Zv6ZhkQtvU8K
lAjc1RxK+READmTLek9UixVC2kHkQScwo5CJGooCTKOgGchjj3B7UcKXMnm9he6kNJIqdN+CSra6
0lP4kPpIVLTH9U9+wyrokpb0HRTgGZ1z8+3lt8Q6hBlWtJsZM77FT/PHYPc/JmppvMC+gruK35wE
/6zgoNVjJfDJTJ07qBdDMt7/Pwmc2LZFfBEb/uFANjauBxn4CSZSgEdH9Fywq4uwU10VXT660NMX
z6vk+fK0D1KqKXBftysnbm0axM0+JQRHvMLdmT007bssyf2oLmNl9Lad98OS4cASXgvh6YA5viNH
wqBzSHoJtvbtjD5u9p37BQZeutk8XGgHjc6iIkWHmSwxxikbRGLDKmaJo8pqPpdv776bUZkqSNwm
Nl7mBYqJcH+fto9c+mw+ifIlviMZqlbRUzkYPo7qAYSqPWUTKgIx0uPs4sWJW0KxtskoJ01PSFfQ
qPbZK0Rg8/UVZu9a9JTPBvlvn1rwEDZHCWNWs3lTmIsrmr53cVirc/NZ7mfVOu9ivS9rElya+KoN
PHgpMc0egvZBXwI6/O4BUdKFWwxPt2PTOOKj4roknJCh5b9AG4EgOV9r2wMlKLCxTHbsQM+i9iQl
rBVwkGcgN8n3a/CMGcXYZBMdSmqcvKTeUtYioFktPPPNxr56boLbfU940Wx0yZP5nqKHzNoSgbxA
mfDX5/+IRfRBFb4N0/BD2YOThiabqSCDuJbhbrounGrw8vWMEGd4Dvi4J5rHuO1hM5Yc6yVf/KOm
Rpsa4UaKYFazdrkkt242I7S4jRMGfo7eW0ie6sXV65xr30CXzapcqlvmTG+SUJNRaUGXa/OP3l3u
YetDowP2sgJ3/v58ZzO334D16jA9xrkgTIBOJN8/B2uTLdFHpI7/LXVId3tIf2bi08YlRmriRAZN
mhoS3alYugZ+UNaL7WUuR05DfEcbCJrdIvW+JKSca+hphg2Pf94g9DGDgC6RAYyAvBYYtcCJ5UpE
urUvRGM6/4wZFauSO7OK4fa+/kuKDHKpcD4LM7LXEHDWTbkuslO/95ujkcq5a6/0MB8o0D5G07//
uLkLvRUsuED/zlMCl6aijAW27rEWaaqZaDx9uaYTEXtZ/JIMAozrt5ViY0SXcvdTWoVCGBE4X0ha
Xq64kp1jzcvB7c3fb1mST4Wpn5U3YIVckcUc6nqs/B8a/xDoPYBLNCeqhAEsydxXSzNEbbluCALN
HrnIP8ZBKW67tmVwB7KawEPzgkriND7u4wfKwAyxyaodX0ydmnH7B3kWVLQCwRHlv3R6/AYa1RVY
MdQWWjVxYkpPuJ1VrX2brA4CDwbts4vLP9CE31mchaoqmgHfh9nd5Rw/IhRbrPZ7MoXgO3yFAoCC
3BujQEcgfDIQfqF0YBLkjY2XiMZAVocgo8hURxlRaVOM58s9A+NJkIKpHLYAJ1j85S0gbv3Zdh75
0HFszU03r8HFnJioFP+Zt5F3t+37J9OL3q7ruAOX/qx6nqJaUd7eSSkTAeBLUA85GB4L2fffhc4V
rAtauITB/YKY56X89LVUed8THczKf2EaW0JC8urIvyZJS9CzeoczO/HiUJUvvNE9WoTGYHw53e9l
EQ0P7Y7E0YLuJ/Ds3to/jbU6wyZ6cL9bKCKDwCWfvs2bVVpBqu1TLkEwQbGpzOY7oEID6y3EL3zZ
eWKPlXG6PR/67jstrPOnDBReIgaS8ZVau62PcgMogWjWbdg6DGmqjaFn+IzihcsTw+c09LZXTW0s
ByYzyWGbCUPj+0FVxeQ0od5nv+5T0P71ZDq582WaCa0ipJS+NXb/cfuiK2PTcB/Q0WOf15Lq0XDs
O1PDVeSn4As8au8pZEMXjgCTgh8PztClxqscd/AxpwtLoxuh+7Kwr4u14vdjo7UFr1kM8+YPptnZ
7M8w9Fnhqd72I9cRd0vQ03PAuPSDvW4wzkbDcTEdBs8HuF+osISEJN4SjXQiNkgSXspl5HT01Vo+
T4U32pQIzJOcBn7izMn+QDmNAPcncnp7M0YzpfNm6eHVpkvnjeS2gI7JMh0W8sTr6zvCARlr2jLi
AhYuOIk6H/AReF4PxKni7aMtwB9TZPyX17Bk0Kk3RI4On3aZzPSuhuqDjRvXWwESH1Mge+L79B2l
v4EkkIZfYIy/V2kS6uX0m49Dxxp7jjAvsvPVMyzwhI6qr5ZPsREfAc2x96xBGPPOWZR7pqRnVQ3n
Tw2YFTLrBnFX200wO0ZbZH2GXXJmTwsj1O/UDfucii49tk/NjKhPtcGGZ+IGw7zQv1tG/Hu7ZSgJ
eKMIxB8m4y5aPolks9d/2yrPO59Ke8EnAZSqko4JiEOwljvFrO0vYCERpgMFmo6yxTeyMMCu3fSJ
Q8ZjYnA9FY9mmuz833YCK6g7PK9mcCWHJy/QxMMIGDl4Bpc9CkrCdlTMvPxIRMBlJFTEciXHjlf6
E+WcRqXvGcjEbb/ZgP2VyG/P0t9aNUfCLZiNr8TvWrXZExt6tUI8iX2UZjfUtmnL4ljZeE0OEYLH
q7Z58zKKCvaVA7FJtnxY5+8SMfrd555+qozcmlzICiinvz2Nzls7lwhSy1f8LefVEXUFqmaSxqoZ
K+K463kL72c3yDNG4QwD9pSTcayFZ1U6cFHHTtKYA4zdJZqSmWZD/8FujQxILaz5XAt32fKvL6ij
8h1NHjZpqfKTOQHR6idYUX1RNnPMXKe2+tsNTncBGYtwydIoocEE3GWO4hwMET7o5qP8voWp1PG2
FUEoul0ADVe7Q+G7OzSMPVbb/N31CNi4DdroYPz8V/WrPbfvIOIgu2ZCI7enTfG94ZonI4jXzQtD
Y10SvvTwOVvRlDr36TXUZh6EZatGUF1LtUZbKKNGwphHa/CkUNn0cSVw2oPGft6d1bLKvwN4p3vp
U4IpvmvoOpue4V+VC8Rlg6ZGk8ZWvyk+L/zGfkq4tcdn/PQlvldABwmV1qz2j+dMMvFlBYBMckT/
crI0N4tekV1m3wFIQz8uY+PUHRzuJzBj1NQBoGnumaKWB8+2YinK0sl0jPz5Bk7aaGleGiwI1x0y
dl8LNT8ySmrstWs4uM8Vauc2iJ9g4TgGH6I+AKFD21/DqtZiyaCCkmlFyqkmE4crOrfraxoL0WnC
4FAl9qduZyfDAqaqnc5eEwU6kXu/5pSTpVddNZFwJz20VtLWeH+pxGCep40CoXBP9TYJQuV1ZmK6
9/qnSwJnSXVCcInyMOKHpfsYJLPOsjNISsuwXVi/i9PQq2bFonFTZ3Gkw93Cg61+M3ohbKNCDgtz
LCG5S7PNrlOjOqbYO2iynab2cuAnsTzKNbdcTUQzEFJ3t6RGksJ2zSm+5GaEk48zjB3U8jb8nCel
MvUBXZkeLms/2bqgTIwT+yw9louvm76e/kn1wjnUJ755sLOtw8OB+UdODrfpjLBLMIOUW0soq2cX
N0NDIobpASXJlZ+G1pduWtbz5izwjTF92LYnplFXALFq0kQDSkc1L5N6/ZynJSb5zyW9KRFF0Q7R
+wOj+v8ze9DZ5gwrxxXyMntAGqd2jJDXGS323DVTyGTeWjtRRUZPLUVE9UuIFktFp/212qSwJ1qn
tB04ZDqR3Hv/xE+WMSi82XUgfozxhX4qf03WypnkY1Rf1GhPvTV4FO1zUqhWliejs9tnzcqVF81I
XUlLdIy0bdGsAG9KyDGTRhacjO/wmiRnUazE54YNFyjIBLythvbTA7mMSbGxFBQdEhLwdhHudN2L
WDDQ9ZfBQXwv09pGzZ9N2klHIhraEvoknqy7h6XoW7CbjJn14TZ+NeYkT+nOtJW9A8MK2rsA14M6
jma+q+BIT//Q7/MkwSr4DJ9heZd48JuOszg5gHdWn1pWb7Ad2owruIddtdFmDybqCjSwQyM9ke5O
nVoGAyuh9OHy4xSR/G5ZruImCKahd8+MmVgfbs6+Zy5IKzIIOsKBOILEpryZCn1/6bXuc4TTucOo
9c/t4XjypnWIQMp/mXx3KpwC3rFRiQnfvlA8YDOlYAa6yT+D454yxZGYijGwUu2A1Nt2dIm1jdyK
ISm0B9NJGDAec17DPxIiFgJxXI07NnItiEs+CG2UgGX/2Lj75MxUFZvtM+UFhfBFVTmCrB8nhnQu
9v/mB7Qto4X6H2QCDDxfGRxBYlo7x++wwHp0lgkoLqXVuKCoVO0dDmvOJBJucrNqQP4ytZHyHBvi
4Sx9QznWJrtJVz6yGNyGQoE5REvBxvCUU6fwFAmWHnqFuVJrYp7dXK2CiMIlA9v2QDVDLs8M27if
+yTr2clUaStb7bVfUiu8arsLiqktmGDVbdiGrG1/j8gYx6MBKdpj8kvqh76G9yqwf98S97Uhy4E7
5FIwttun9WmYwXlcZVtWLtDyygtMBqHbgWPhHTKCOoYD8CB2/C+t6mnAScKdq9pEU1PhXty4+Xyn
JoNg/+DXoxafimmnQ8/ZZcyMW37A2AtLtsKdAJts+ycoOPQO2wpDANMfjjWL4CvfCjX95vtJVkF+
jfbIQ+ROxI/XMzgGWhT9w+9r6BYOW9LLc8lqDF3x54nP07wO5So59t2NMCcvyJt7d5mjTipFXuf6
GrhoWbScH38a7YpzFV7pU9l9pTpSQ5qjocS1jrp4BKKHzyRDRJv8S1KfXhAw3/Kl8K9EvZO/qB0N
ofQm3wEP4dDZCM/ZlMy0huvT9RGzo6eThLoh2Sm1XAAIIYt/qQg89MWZfOqLMkNkmlWyvGovh2Va
M06Fsnv1FCep81JsxXCMqqhPIDfk61HwATtxyZnPwrCGT/i3x/902t/V3f5KiPkjiNUn5CWFC04z
zETmqem3K93A0CD7xf5sjZpXuKQh0ffDeKClHTXV8Y9iy4UHNcOd8AwhUiOluBWh9I2CE96CIiBN
VY4eOcF2RMyySY2oYqFpQpboARf6B5b2zhbxGl8916YpYBgM5kWXkvuIOTw5ciQEQE9n/UlFdjaV
QkHp7Z9WHi1EcDn8XfERVO0WBL/nMBfW6pPbPb5po2UzTkMHITELE/Ev6/ZlBRR9L3jiehgiDVmP
det67+npBIMMxgqTqFOsmLBCvEg70imku1VSJe+ZhJMGdJpSNNfncO5Ftm942q3NzOGgyxUq9UB1
SnSZw79IH6vFcU2DfF89vxpFERCQTtUF11UcL74X0R207NC9FubZ2XCAaIFJlXF13ePozf8O9SP9
1NDb5EOntZaYR720ejSWV04nEftNKE/WEcLCOoHvX2aiMjUJP0mYHCxFR2gQg2e5hu2J03lSwVDM
kUP3G2y3qY+oC/AcXs1SRyojQxWJkkyCKRgRpltmhdvOSptHviJVi+WjSYhyUxGY5vmD/iDg6vaX
d6lrc1ngZnNYd73ZZVXKsxSWFhfWj7ho/PFTiAq81swjtZV1ChDJEB7bfMTYVLI7YsUYnLMsLcoj
s4zU8D4349DLM4ob9W1qcckz2gZNcfOn4kPIaQ9JRxaJ7Y3UvLE05xusmZ1zTgaMDHRAS0mzIQi3
sYikbtgmBzR9DTz3IqJGLqGjFde4luodyMq8jT3aNScZadgE/xtnfz0idAAun/yvZlkvf6sz73Jg
jBm0pKZckQQAfTg09McvXNS19tbrbDysc107KNRcoN0CCkMq7bdyh1IPoSTikS23heOr4y8qbWdo
qTBezNLdZwmcS/tNr5NPeKAE3ENFVQ715twQ1H0++W5PHIO+l8nZdKs6PZS/lQAPSVM0v9N96wOR
XkRQoEMlcnCD8qKpUiakBFUyhURaPxWv2LMyPwLc+vf+QI4xRg0Jh8J5AnzMYUyiksMTFglcsIfx
T4m2ImLwk+IER+71IUatumkYFB/3pcbiCxw+15ZfOlmkl5vQFqgvwFJDdYeiVmzSAs6BEmzwvjqQ
4OkjtEEwxhyi/EGaJA7pD8NAvY9uhMuKlMH9LGN0brfkCzlDjmbE8MaOGojDR5j+OPgHDvkx/3hA
gQCgZVIezsQ4O6u20Ik4WTjKZ3P2cHeGCShiSZzgCBZ1D2y6U+hBSq54u8FXWUm72GGEhFTfQXLA
L7yFIbJlkyXSeoOXkWlpPOpR7dTs0M47SJLnlY2knXUeroLs7zDliT4BqO75Wdfm0HB3IeKP1laj
YQ9EtYJCHtgssEk4cR4zh9tr+QtI/XgU7qLUP0a6lVFyWg2uVKMziwKqCkWRJSV0Bki6j2mF9jJv
nxiO/zFMoc5tJ8E0KfgHH6d22xyNmaatWO3zow+97RMBKF/BhRFaCc7vvaGU9ewJx6clDUbT8/hQ
kknZdzAukouceSzdPxZNTy3noEkjAiNPUhoOwBzQdN+QGwUHRT/clSY3RQB2uzOm6EklSyycte3q
0wwO9KJa9h6lb8dTp3CF0UFguxshI7kecGG9sgja61D9m6CE9kJtDl0taTa86jDLdduEUoRVR8pg
7caem8Bb3jv9dvzNoCd6zn931tsIfhwgKfWhT+O//CmC3s3M0eBvHqWS9ADXfTxVkrB3TWYDp/6m
bn0SvHtbPn7JvsvE/VX82HZ39xMUItRIJlwwiPrrisqyZAG1sVLyDYvq8SrxFnib77p1sKjbqJSy
jYr3i0P+Jof+LZUmLw5xagsea5ncFIo9K1L4FMMPUjToBoVMGK+49TgPk2q9htg98RQvGe6VpFqo
fEWHOmLohG900Ci21r4yfy6WV0yEL4aXtYw4XRNCh/VOOmV7ceaGReWDVu1ucDEUBgP6o3yFDZQd
pZHdbNT7R1SkpimiOZk4lm0dD+IxpF6YzrFzZi3umlSeS+FMBl/teWsknAs6uCYYCYPoJqGGbAUh
2jCFmviDkniqCxuDsrHkCJGkdXg2lfYQQIOy3mBnLNrSYLotvWKYLsGIurXq2IxXkqj5qgnvbakJ
K9xeo0NXqrqD1m43nYz7VhmKWOS8l7LOAFiXPTrXwq98X6asQwMF7qM0OeSzpZrx1Sx4ypuBHxRS
KQNt+4x66+Icun64qJJb9OAboegJpL8FPxzQB99kudFwZfO45o3J53hpu3KRydeMTERNJXNYj1Au
pWD0TJ945tNrS99KeSHQJi6g3Gx0J8mcO/TfOkENRtjLlbOqMnRLtC7ePNPUGPyUrUF5D94Pcolb
dWIrGTzf7f0IpIPCw4crQsKzoAWChShcnQVywRhL1dzO1msx9ojQ65tmM2rjJVnbvpLWo/c0cgP2
qsJDmTONF0oFFPWEuJVPV/VgLhN0m+sAaDo8iHpMClsT+p7bcSHrItWrlThxHY2H3Hw137s1tRke
5yCNLOCxvulrU/NNj/Aa79AxZOwZL5QkAdGL9aEsOHQzO3HHP4XuS/gSQJ+xAe7BHY5mjtl0F0nQ
hpajkR0Yxnc31NetlXmh5nQeiRDxxf1g1FfSKaMkIHEGfPRIfT0Ueax5r4T2cbQzRbmf/vxfGBuI
1oBZrupVBzlnQVsSbdkGIDEEn4hxGL+xpy0F9u4zTMFKypvgn2L25hR4i/S6PY1XAYWn5cO52bx1
Ih8UkeWBQODVnn5K8TngUeMklA9UVK8Dywy7Lpxkiw7DU1RcfizmG4nBSpA2npqRemKDEOHHwKm/
OOwsu3qA1B/sVp+TwFWTrLxqh/t7pyFUOt31uWBdFwmpXFZB+fzfzm8jyB38uNwvdLEcrlde4Cx2
rPggssVuwuCBUDkDpggyEgdZ8hz3BFNR/YTn2vcyXcdYCmAk///PDCbDgzj4joqjasNV7u92zEHA
PeQhgwJ+VbPDABcue18s1wNUktGRp3hfgorEQuNUBbMeJ7kSTLevxEJZkp1L/BoD7M3pC6kI/saf
59WzygHG1Ho061QRY2u7HXpMs7U8+Pe8MYGNucfHkHkQ/09i8njJGQwWg4fBEKCjpSbP8zjINI7K
FtK7p0o0+jaeIAmFfHjoCIfjSv4OA1KZb2koy34yRcOODX1/B5JgVsRJMsV97t4sEOADw+pzp84R
VZPjDbsqn6wexJEWtAk8S9jZ68ykQ5od8WAONx+cbeKwTszkVHIJ4tJspsQVFZK8qjPp5ZRiOh9t
F1pilDzfrovV1+cwaTk3SJw1qxmNCkUrTlMhPCYnp91IBuLkkDPxORtHDmPYSGAcehuns1CsmpMv
y8dsQtXaeMUW/TM4rHBKYpRG/YlT8NzmCRWHEqky9xQ6BgPEjjHY9kYjTvxmUXdRtxgRJNApAl6B
OD8EwT6kWpZe+ZDU4qmOQVKL7lAB01Wy0PfEFWA60dFIjU/IwznkAVGZhhH3YdPrmKS96LnuYiYw
TFyKu2SgXvQEPYwCCCne9H/DoAjFeX6JDNjlIkZhies1MD9CsFzl75xELDspJm9TAKid6G6Vds7c
bSKkun7q8AAhXs3ysoGzFJKhECRz781afThoaR+M/6upas/cQIoSRDBRjq4x4HoYX9lqciUNO4o0
jGYlafP8AUXAnzhom3cFV9Lu2AJWxinxbqflxhhUbF2D0Q7QqJa7kX0pPs2cWQ0mBeS74BKkah3y
4eA0w2H7ET36anbgNmpso8D0HPLZ1RjektLwuO0VpCUhwJtWiel/69SPDeTE5/baFChRe33Rt8iZ
ol1D0QfFUYZgHHAt7/0YfhwdnCcpsIJO+3TGIBE1gRJuHuepmRrM8f5FitVMhTKCbndNmjW+MCZM
mPV9aZy0q2PE4DOZC4BO9CCUS6DElFVteP9LBmy0GoVKT1tGrzU0jFJDiFtrjm5/VD+qFbB7BUVN
VnaNRXg0iZIrJgtIsC1iwQO77ByOeK0vaUV39WGRT7EkyG5/5SVqBWuV4zvlxMSEf7lvOzi2AAry
zl4qn5b4RODl8qgOIK0j1yZNISZBBX7OEsAEa6zZlq+lKbguFYxn/4Zi0lNsdM57U26DOWkDHxcL
ntTmKWKv4nxEY+H8Kl1opA/V3dsYKlgip7acDIm5hjI0l8QbuOwzQP98KBRL0x8ycS3FTEuYKACf
zFpbxJbFVVCzyIkLPH5tAdB2UBb0LTdM+mQ4b65Txx+2lrQ6hjwQMEtkH+yM4rmxCUnMBIZS+kS0
UQTX0jrHrZBD1OFe1Qq8Hqxpucy9MDnlhbOk6fDYzIVT34++FprYMuKzKXFcW15TRka8/7/K/1qP
9Ff6uKiXYh77o3RRmTiJEJWc+VBtkILBmR00nbvk9KVR9Tz/RFooYVOxi7zHD+P05I93WpCLdA/v
Yd4NnLLSHYtgDbrb4+TlBub9BBbLoqahn+8oC0+P+6kDaT3q7iJAw/l+k3gt360qSafrjs2A3dn6
GWRdzBWqAwjORqE2cWjSkwHrbOdymxYRL7ce5/WYLcEBSklNh2wVumInf5+WHmiygFm5v6r2w4Zu
cBB0aZW47i5cR6xUFnWCXjf3i/iyPar3ZJw7Kddkw5LqxBAVyyhj7gAlhG/8kmQCqVysrn1vLYGo
r/VbAWXd9H2yvyHwBqQG45keArQ/BCLvIEg9R0zUvx85TtV7lleWgwm24dVwyKlBLjLNQnOZ6iiP
XlWPUKyq7inZB3AGwjGF1WIyXl6iLyR3gYt9kEqeRz2fRvhwebF/MnkSg3/91tfsvWoivGeRz041
mDV9loqu+3Pjnh6Q0qrhMBAAZNtbTMxPakjwYJMXavWYvs3x+xCILURKRu7G7XOv4XXBGkYn9DPG
qQGr8A8nQw1crREfijJVVr6YElGddb2STNG5T0EsfE2Ackyd/bJ7ca/U0ZrIZ6xpIjnwubnABmCo
kInaq6tZbgFSlgpo4JXxYk0OHmU96bikOAncJO+H5ja6B/HSdeKYd/ye+XfFhPPaMSKdgklUVXBl
Bn5Qlgi7tMMc5ikApGORsHWpv1to8AksrDdqtplp8M7Z+bkUCO1B0SWoYu8Tqp4sYpNK+9VVXVVr
OuzT+jknGKK3akezz2kwrEb6jGUIQ1kpFMllmD60tj2rPMO19Vn0hrOAZqfOJjtF6SHg3d5Z68O8
5Ril3DdD8a/WXaEUQCMEhIHpxO0BLjMbc/j3QjicCVyRyyIdlGn7jLRx2SwiHL/D/NVmcdVRGQvZ
Vq8oOoIrjh/XTB8inUqKzFVZ38l01CpMfhvkvQzKtuUUgLybgWUb8c/oODO37pPI3JaD0nWf1Xmm
aiBjBjW9Qh8HB3wYNAJAfR+jPR8SzsDlFwOfvLurO4k0dbe5qJAnQzHOP58m3rX3gyAGHoD9F+6a
ZtXBT2l0MTnzTAQWVyLAprWeYhRGbSbg4Q4gtYExUH5av1NEDQVDJ/BewBU0yKeasDtTVfbMAENf
f+dUPs64z6Egv/SELjlwWRK8a+t/cyHNSnJ8IxUNSQ2gIzpf47zOEb+hsATlC0xg3biU79Yn5HhR
kA==
`protect end_protected
