��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl8��M@�	>�Zk_�j�$������#k� y�B�I�5z�ӊ߇��>	)3@�מ8�U��ѳ8����1c�I#q9��5��<
��H+���
��=5��a�(A���{��I���S�j�X��_���X���r5�ď�=Ubh�� �p�����~��$zQQ}�+�eɶL�709����|&�^w�������=�&�5)�N�`%oL9�.\x�|.��0>����;��N"v���]��0;j�.�j�[@��9R��"S.?�+�pM���Z��H<�0i+
U��'�{g�n�}���I�!��$s�מ�T�k�;���z�jl��-8�v��Dz��6���}=�UQ�ų-�psz/g�S��~g�^����dЎ[qW��Lְ�7�RMr��Zٿf�u�����M��^���D�ɕ����	�ʝ#Qbq��*���{9���Eȥ����	2� j�Ggܷ/QtJꠜ�;���'#ߊc�u��d��]�Q�i^,dB	����մ�n�۱F�e]C����M��-�����y���wUj��2J��*맏���*7@?w5�t ��M�&��4�[1�܈x�"}�Yv�=N�/Y��<������,p�U݌@K,Lj��Y��������{�>��<�1E��@�J+���
� Ο��>J����
W�c��̥���*1��(H��j����}��?�/䣡�� *踒����	H�띥B�w3F݊7�`�<���C=��&�&�) &��EV������+��"���9B9�]ҏȡJ���4��8������P��]�l�&ε������l�]� b�:��zw�z�1Kz&9;뒃H@�C�O<d�=�}v|��gׇ�Dd�&�'�Β�6z����B�)CA�`�8Z�C�51I���瓮q�~Ge��[C6,ğt	z�G� L�iu�B?�������X̯��~� �#���՝'�L�	4�}�� ���Wa�-�~ij�R�u)*D���A�����C�pE�3�;>5~�F�g>'��ܢ�����V�B#��-/�\�kԻU?����O�~��CI��í���m�R���1����3sͼ�<~����w��Xۻu6UG���AA��E�'���?�C
|��\	�c�F��Ge�!�
�\|���+����ԍt���U*���D1I��X��I�@@�̵�4�]̓:e�<�[�0zz�����y�����[���aP��&��$��b��b�����/�tb��rp��ǯ��ԋ%c�CeOH��y��D���aļ쌿vwߒͧ��f)Q i��b��Tؖ���}J���&�߹�X��ԝ�|����B`�3����9�œP'����s.,��M������-������z&3�l����J+Ɣ�?X-5ߋSϣ��A��J{�	�U�-}�o>�Y�̉6��v�z��럑`;��}�q��$yH;D3m	䌮Rf�M+��	��/��y2�)3��� ��fB��vB�Z�}A�u�����mH��70u=<Y�K�6O$�S��{�@��Ƴ�X�Ӈ��h�YP��{iU J3�MS�pQ�p���땛Y�>�K��E{���ty�`u�~i�xoR8�$w����Y������bF����[�S�;(@NQ�q	�l��T��a��u/RϨ�u)r�A3�A��/~S�YGm_m�Y��Nԍ�A�!i/�:���x�ҭ)ڊ4��F�Z�^ڏ�T��ȅRe�}|��蝂�@�v�M�-m��2Q
�Ip�"n�mC!�Ϊ	�*�XY� �g8�V��'��r=cS�@L3�} �BKg�u}�	���H�v��ĉd&qT=IS�nf<Xh S��=+y�0'�:���n,(aՑd�A�G;;͆pXYv�'%D�e��`C�J����z\�^���%_x&Ϛ�.t��7��ȹ_��;f���qL�!_"�3�$�-tV	E��������D��oK�4��M�in&�>�#Pj�EВ�CXA�{�n��,3����-_R��Lʧ7�/��ȹ�X��1`;Zi���[GD�ih)��A�>���ވO��c>K
[���-н��� ����D}�h)G�ȃ������$:��h$���Q�+1�����.�~`l��=�e5�]�K�u�M�Y/�?=B�Z��mx�֮��~z�9�I�Z!��2HCu�@�$����W��~+���28�h�<�u3�*�����<Ӯ�M%'<�Ly���F}';0kB&�L3���~�+k�~�9�ldͼ�HF|��vc[^PO�3��R_���H�j��c�p�ϴ�o+P���Sןr�R27��REt� (�C���ֵ%���u�z{�������;����+��`������k��b���L�=ñ%D��К��9�q!�8�x�/7#����K^7�����Q �)�u�[�-�Q�k�i�!»yͯ�?4uC��~�)@7i��_l�'#+`]|=c4`�l��Ox/�>92�0��C�klZ��>�r@����r�p�N �~�>� ]BU�mBr�b�ՠ��{�`�_3�k�̦W@��`P����/�| N��7��g��F%�5����#+��q��S(�3}�se�k���T�.D^7��W�@�"���÷���az.Tw����?�%��ݢ{JA`��*Bû�{cv�0���Ok��Ȱ���-y�N~M��qJ'��\JX�?t�a�:U�G\�Nl��Vv=�����sA<[���L�W_�_��B�S�?�s���q��%;)N�UV��>I?�S՟�#fݓ%������$=��[�k��h��1ؖ�����Q��������ڎ��4s�H��'<X��$f��*@��,Z�c����T'	D�FS����;�/b�:R`4��H�g�K+�ͅ���U�'$v��pp�(M�OmM���Isִ���
/���3YϿs�0��)���`�{�y��#uK.�Ld2r���fTˋ�>��ԁ9Z�;���:�=wQ:����	k��J$!,��l}��=1`f�~���
G�5$h#0";�7&K�o���m�����1����O�FZq�+Z�x��vN���E�UUV�N�?����[J�]�9�4��>\��F�uFt!����@=�@{��Nw�����YC韷��i]����`��e6`�ɺWQ~Y�� UF`c?���+��N(Y)-�%���(V0f|������6x?�@N��L+[�o�X�螟I�C]�aC�w��Q��9�6z��3��;�h����a���л��~y��5M�����e�\?��;�9Ϻi,_L6��v����?oۓ?���G�x6��������A������ǔL�Ah���/]�P����+ٶ ��>�ǉ	G�T��m��#�M�������c�<>`�DS�\
�qL��r
�I�����*3��#�7�j� �i�)�Td��.��*4%L2�R,%��"����)z7TY]l��		^��nn���)vɍ���ń	������U�2T@o�aۯ���J`���d�m����K~9�9i��>r�/|x��N�H6*/zK$�"�!_8�";�ڄ��@��B9,����'Tܚ3k�𶙹���J!���b�ri\/�a���0�h�K� S���&��d�q��F4�u�������k��K��CMiUo�=��V�#��Vt�x����J6�''x^��]=U;��[��q#� ������B�Fo�	AEV���yt{2�b�#��*͌�<S;���V ���Պ�Z,��[ܷE_l�4�+���6�f��_b�o����ɦ�w�у���d���V��qŧ$!2BĚ�&v�}h�r��;�+H���KB�+<����_Iru34��r��H�ae���{��8Hx R�7�|o~oֹ x�S�h�'_"�E`m�y���9�W�%��&e�ۦ�;ی��?<3zW�����BF,�����eT�g�*5����y%�G��2�Q�[|��(� ��Z�$f"@�S�+ٶ?>�^�6uґ��>oՄ>m�-G1�[�!L��h��./�}2�d?�y�;�˝+���B����7S�@0�~*��p��� #��֘R��զ�I�+����D��oʃ�;Z��'���/��eO��VJ�~����y!ɟ�h��$�v�n��*)��yՕ8�I� p*G���$�=��D���m�@U��.k������E��|;o\�iL��zX�l�4�SաܬA���a��N�Z��E���M��Nw&u���4>����fO,t.Q� u�69�"��$�Vp�IQ��A�1�����
�����#F���.Ngi�7Dn�0�Ck% Q�7E��@�H��}�Uu
X)epG�B�|(&3���]�j��cӱ�_��7 �{KF��<q�g"�.?���'Q,�Ny`�_�iJ@�u���s�V&�otw*A�]����W{v��Va�2�	�%�T8� �����X��������W���(c٨1��ܼ=�bX9e�RN��D�!	��r����=Z�)��!�
i4"��߯��ܖ�q���PʓJ9ff�"`���]������M�{�xҵ�;d�P녪3�Zl�~�jH]�m�B��_5�I��C` �]��T>(2���O�,�F�Z����&�O���j�Y�4͇��,������T�Ee%u4x��Mԫ;���<P��p.��0�ga��˄�B!�ET:%������˄��2�_��8fM�΀��2ų��!�qr^1�z�5g����[*�C:o��'��>�����j�ΤؚV!�U:޽fw���x��z�>�`,�,��� �\�Y(�cQ@3.=f-6ʆw��^�\^_�<�����z#vW�uEAʀK���޻1��TnX�F#u>&kr��r��q\?�t���(�(�*��o��U�:��cWb���Ο�J�R�F'���H�S�X|���X���v`8K����h����ۦ�!&���X:�	.��85y�Ы���ێ�_����+���Ԝy�t��E�>�7��S��bRtj��2Խ�+>ԭ��%�
$�z�i�ڊ��������O*d�AY�r#�)d��5��Vg��uB�|���x��뿟�mL�G��l�Z�2V��w�����]�� �m̈́�?8z\M�K�C��M�ng���T��Q��Dt���R�cÇr�@���9t�7�
)�����f��8rOl���a���0�;{�
[e�H��I��c�8�D�tql:��0���2��e)�`(�Dq����C�OVBo�uno�y_S@�_���#���.T�����q|QS+~]����ms��\�fL���d��[�D���L��.�ʟs��IO
}au����A,�߶�ŭEfs6�]��Թ}�neh'v�J�Т�~YNP_tv[ܐ��'ן�č����C��>w�$Ri��q6���D�k�� j�Dh��;���ID��Λ{_�셡���s�]t>S1<y�u�3uҐ�n�B�S��n�0-�O�4��Z��E�v7�B#7��	���Vj?i�G;�a��,��q#E
���;���NW����y�g�]�]���M��~I�-vAFF	�s�.Y���N���v�R
���u ��YqO��K
۾)s�d�*�C���C-x��#M�X���5��J@)=���P3m�r��>@�>�I���n�|*���(��9��AMj
���~0_����*VyA���r�2Dn?�K�٧w����a_"{������S`��kD	b�M���3h��a	� 33_e�n�de2�ĲQb��Yʓ���~�x
R��l�P��d�I�=��N �-��%c����~;�#������+�swo�FJ�}8ݰ�ks�_�Y6&۩�k��X� �ػR;k�5 ���ߵ��駥������B!I�=s�Č��d[im��o��o�&���/�$��W�LI\z�;�+,�X��'���G�u3�芖܋�0羥#edD��ϔ�gf������-����Q�6�5��5�Di�R<.N��\��J�V�]���I�#T�r��N�@���2�O=5wuj(\W�C��k@�U��^H���|�.3�{e��r����d6���-S�#��!��S�q�m�\�n��fyB�p���+�N�S��k�fҁ�L�Wh� �#=���,Pn�>H�@��4>�,�Z�LJ�}�R�pY�)���F�nR`�"]�܃���v �(�|~BZ�Ȧ�6�0`�J��Z�^��3=�ަR�M�T1U�$�g�e��n�C��vI�R �Q���R_�i��N��6$�Q	��Y��[[���m�����Ĝt��I��o�d:��գ�s;Nu���ڀ#�·}�7�2�*�4��v�^�X�Uѩ���9YM%_�K_���p�J1��&��\�I�ք��z?��	�f�ؚ��{aE�#8�ݔ�q��e��?��Pm��Z��s�sF29��t=ϞQP��L(+z+.�����5۸��#�B,8������{��v��C�,oXD���N��q��|��Go��f
N�[�[�_bSϺ���_lL�\w�����A����!��Hd��~v1�0^!T:#5���L�夝	צ�v��ldu6А�5������'�8��;y�N�������`>>R?̌tS��q�ު���f�Xn����W��`(�_`�jp��x�	�D���}Qvb�%Z����6�/$�R~�ռ4+Һ�_���$�d�u�#����{ĳJ�l됽25�٬�s�m�8�Xp���µ�2V��%넨�T�}��։�"�o�B�5Ԃ|���L%���-�X����ƽ��N����I�� �r
�H8����1`	nY�=��,5~���ؾ�A�0(_u��e�	���{;��El;K�U!MS��x�ZD�B_��K���.�x�l���H�r`��k�u�����TJf̕��Z^s��Y��8l٭  �_k^�v/C���`�2.9p�O��1QO�H7~C����ѣ+����vJ�N6�<i^@�e5<y�Z){���2�Z=�AՀ�s@����`U������v-H�0�2��#�� /3�1����FIؘ{�!F#�Bɝ8D���E�ɲ��F:.�O��j�=�s��U��%.9Zj���s��E,�qI�W�҉�O|���
c!90D�-�W.��C^�u���"�R��F�*U����V��i�o�Ic�n�v#1��pT�W�� r|C5/��#%��f�Q��)����X?~�^q&0磢p���%Ob���
�4{M[�:�l�;Ր2��sp�
qƻ�����E�>��$��K�� �s����\�c���o�r�#�^�'��t�*�D�E�"(.|�_���@Ε�69�]֘ۛ8����!9"n�k_�#%���;=e
|���px� Twҩu�8Yg�!+����OG�0��a��g��f�ݔE��yy�h0t��<
���(�Q�܉ӫI��Y07��kO)�I4ͯvnV�HBb�]t=&�H�oZ`�|���������8Gu_v�X|%���=�!��ܫ��o�� �uh灁r��I��}	��ӠQ_h�*��Z�s�޴毼����&���,+T�����>�;Z@*P�h6�B��i}ռ"���q���*]R�k�@�o��F��R	8�":)��jJ�����R)�zϖ�Ѐ��(�̌�j/��ԑ�-z�T��[��J��ߊ��������u�[a��q��p�Pߖ���?� D7����k�5=i��w���
�q�I��,[����C���B*��F4����f}��W�I��2�'��j��g����������Q�r�-�rs�w��$I�2js�Wy�O��#�`j]3x=�
��T����f�(c�3+M�t��H�i	;l���;��������V��l��%�'~4{[�~���v�\=h�*Lk��)��UV0t~˹8� WY(W�O�ќX��!�殄��e�k|��]e�&n��T8�#w�VxN�$��LQ��a1���
�4���i�G$s�֛@ڐWb����ZY�w�z�8m���/r��&cY�7����Ә2��U�$䖆��^ծL'�*��6홃5���w��t���wbE<
#�
rm��n�+{�ń�<ZGm��iV֤���;�8xqFf�nlt��ҩ	�_��b��!�yay�-���^��O�%ԏ�fΣ�̾sߚ��*?��������{�'c�-��R��wy����'�qT��:x:xF�4�:?��iJ|���?�@Hx��ؒ�C(���+���ȸL�1����3����S��zt������&%��<A0�ܽh�O�nO���r  �k����`FT�@�H�����-G5�A&vS������@NS$��v >����V����+b��*x~�8��O_���-�+#�����>B��'ϒй��N+G�H��Q\hv���M�S��)8�4�'=щ-�nU���Ni��)DO��9.����� L���ţYz�^ؓ)��8�l�W��nΙ�10'��)��>d}��Z��~�V&?r��<}]|\���,�+a�!���ɝȏ��Yfp�%Ӗ�@���(~�����l?:���t��m�5E�1��:�(A�ԮFS]�&S�GǺ,��)@k[����fvM��^S&��-	�=�FU>�[�Y�K�W�������`PR���T����l�(m��-����
�=�ͅ`�f$S&7�V���>TԈ�7�s������Q��[��E�\y�5ޥ�A�V��u�nB�>��":ױ���'����o��u�v�J�B" MMy�Z&��@��k��5�g[�{C^��Mo����
h�y�"��r	:�L�Nw�s��Imɛe^;�&$H�x��Z��(�|��A!�aBC�����|�(��@��{�I���%`�И��J*�9LX�Ee=N�2�����bFccyA���#��&�����5Mr��Z�U�w����Eh]t��j�~H'�p�d�l�M�~�@�5
�.���CO86"�=\�TziA/I����4�Hcfg��j�G���'�퓫,&[(���7G�u�����>L�� ���
0 �u!���Wh8�B��Z��5^�p���U����+3.]"J�/=c��
Mi��@�?{��[�w�۫�M����w��pN����@�f9�����6Gt��
$ڢ�{^0�a�q�O	3���:�3��,�Y5��yêȱ�j�Uǿ�w�
ũR�,�x�j};J���&ny��7��Q��?�;G�����c��eP&*GAğE�~�P��
��E��c�Y&)�暴�)�hw�EopäaoS�V �SPdZGP����Ұ������Y�e�
?g�{�d�����O�<��5�≗5l!R zCzƝ=��0eګ�Mֆ�>hP)�����߱{���/�Il�ge��6_瘕��B���ujA��	���a�Ɋ�C�R���ڎD/����P����ަ�����drVhW X�#I#��+�
�}�z�S�j�	�5�[xo��%�O3h����oW9p
��^:��P|ųIAT�A��!�n�#�W�!�'����Ӗ�R��R�����������`�t�]���������w�z>�מv��+�io5G�Q��ZTl�����ڸ<d9�S%�w$.31$����e�'�J�A���S���,G�:,(��󯪱G@��((�Rk�M����\��G,���g�B���S��i�㠕�N9�}[m3a�pfU���sqz�Lׇ�,Ъ��ż^8\.8*���|�"K��	�y
�t2`���"^��9�L�,�bB%J�|`�e� Xx�RHCcݪ�e��:� �蟨�� s0�b��l��>��c�m���@�:�`v���0���7�凪
��Ot���b�-`w���ge�[eKƉ?2���Ԕ/��M\r��ɭ�tIp��H23�+��P�}S�4j�����L�v��DG���_�/�f>�q+�Ι�dYi�[�ձ�tc^O�!�S��Z֬�V[S��h��Ņ�E�H��2u�0�GJ��7��ˏo�np�*
�~�t�:�`�����u5R���&����@��t]'W|��<�3g�Yw��b?=�÷l&{�
11�zp����gQ���#0�h�p��%���4	��4P@ۤ��߿�rbH)���"���P�R�|�Fe�w�,_�Aqv��:��w\~����fL�G8�����> f\�>2M��r�UҲQ�N(��B��j��� Nx�#������+�]Y3t�;�551��~*�$.���23E���غ�3�z��|\ɚIϕzK3>�D9愦���U���Ig?��f� �7���O�SD��la���ĬN��4�?�P��
M�g�ͣex"8.��z*`�t�aC|����?x+�!=_]��=���݉�γ]���g�~;1ƀ�\�/����Q�gQk�F}� �Rq�cEE� ��V�r��q���䘧��l�ȇ��6�*�̽_�ض�:��������A�JX��ߪ�Q�
v�5�' �����B�F�H>L�(��0�6�����ܐ	�I�zղ7Ν/���F��rh��4��I���{�8�Dk���+k}��αj�,��Rt�i�͎Q;Ԁ�ET�C��~�V9�yx؋�xx���D��-jտyF�;��D�7Ը��5tZ(:�<��B����*|�R#�1c�b�QI=��*���_swBK��۞��P3�X��/��LA��9jM��樹��l�ϴZѣ�̀|'���\�9T�%����|�P)x���Q,.�1X��糂Vl����-�	�񍧢Y��`������HM�'D�4L�{������J�$�'���� j$��ķ[�=��ޜ[= w4{ ��]��Y�T���^Oꛯ�5�� LV��;c�����s$�_w��3%5V��a-�'�3�)����xS�h������Pc��Y�&��ԋ��=Q�����u+48��~d��$���r-r�i\���(�M?h��0%���E>����� ��$�)=lm��<0��rZ=Y����X����9�yC�.�Tq��z唚�!e�ʴ
Q�z���D��S�M$퀁a_� �h�6
؇�f��I1Y�L�
,���*�"n��І�[!>�����c|5��;X�^TA�H]|Mj(�R�������8�po�=%~���q�\�nf�-	��1*𷂇�Ƀȋ���a�5^u�ϤD�A����.dJ����mmj�"UV�*f�}Y�v�'�����(D{ؗ�e�I�5	;��vϫi�=y,�e]g-�x3~0�j�D��o������[�XЀLN�no5�;��r�A֚�^�D-k΀�C�'xх?e}
~2/�6�4gPB�D/yr��r��ˇ-�.�l�u���q��&��}�/��Ȗ�.$�[�s���̎�� �k�#�6�I���K�)�g�P��Z����E�7�<'��(c���	�y�y�7��D�1V��$&`W*�##&�)����i&N�F������"�-G,��D�_��f�H�7	?���1<:�G�6l�N�O�p�Q���K�C-E��7�t YG�J0;�������9Y�Vy�Kt+yjT:L�3��[̷'�����re�>W�6�V���$�m��y~/�$�Qx���ed�l���2���n�>�R���ڪ�:��f��r੣�� JV,3��ఃh��ua'���
VwSoef��9lƒ��H�Ef�ڀ�	2/��"W`?���+�'JE��)�(��(�i�.*���du���ِ�y��H����u���9(_��
��Yk��ţ����[w�V;���X���U��z1���KY&�d���+�}��u�v��}&,>ʉ��~����(l1#^��G^HԚ$g��X��;ӈ�|'��ƺ����'��e�:���Gt[�X�^��J,lPUOu��8�i�|��[���l�56����e�N���|L��%Z��ъ�+�ڦφ�}����^�?�c��df ?��.��\ �8��Z���h��'u��έY������G�(��z^��sʹ'F�{GD������O$�b溭��@<ǭ����9�w�C��X���yHâ�/���G �q�9:�vnj2�2�KF�5�v5�&��NA���d�8�k��*G��9Z���E�����I����Gi�X% �p���w�����L�V1��(Ky�o�^7�La��Y3[<W��r���n��7ʊ=X��ٯ+�?�r���p� �t��4�q�}�DV|�����D�N��	T��`�M*x,����ׄ��������y����V�
cw��I��S߰�(�%����� _��b�w<�]��'�P(m"ƱU��&�LO�N�zϠKR��8m��;��:�x鍥!"SƵu���!�9.�ֆ�|��9���*ع���q��A'܁�(���6_�XCv1��W�nq)+� *yx�^ę����0/ϣ^cvd !0NJ�;�1	G���}�?�^q��G��|����zU�e
uW((�a�a�	_�p��$����$'쯟����/�%���7KdUZq��-o�=}��k�{�i˘����v�6�dӡC`(�͘@C踵�a1����[�{'�?H����Pr���˾��I��M�f��Vݘ\�m|����N��)Z ȷ=`�W��~��$_**����g�tؐ���EuΌ�W��'ꝊN+U�Ր%9o{�~|��$O)_`0X�����a6����/r����J�I�ߤu6?%����������*M�t�/U�徜=�f:�$̶����"�O�`��=m��|�s��u(PA������܍�J�Q�cVω�<��j�@���(��V�!�2g�v����GQ�.wŤ��̠s�m�{f��\!^ইr�q���s"j��r��)��ϧ{ '��?��K�q�MU���5_�S�Vq8�~�0���*-r�1��C`�ZNη.P� [�3σ^{��D���F��F
�P����@�80����ۣ�%�O�g6�b����HL�毈������t��}��8JN�CO�0���#+>.
�kW�%�q �t��hw�/3c	��|9�b�NC>�?[�;���Q"J�>�χ@s^a��2��;��xk�u&�&�	ȋ�{�,i6��40���	��t���P2P�ۮ¹_,Ƿ���+dw��ߐ��n�g�%�Y+#������ {\���H� ���-H����Π ��Q�d�B�@_��xZt�.{C"�ɗ��`��~�;���\ܻpZ����z��|`H~�]��e��N�݊������Ԓ�|�?2�a�CD�'j:QC�o��*�,�H�/dE�땩i����%�#n�c� ڴ��(��S�����^�	c
��_��:2�>h������a7�D�b��,��'�z�f��<B<�����ؿ`����
��ڷ#���cz�v���n��2H�1Iuy�p�ĝ(�>��º�~c�s�o�jb���|�IS��G��X�h�H$p�l!�Q��*������-�M��U�V�o0�|�ce!�mCxY�������	�;n㣤v2��]l���@g��&}%r�I��Ĥ��)Q� �e�?=���"p��`>Qf�?ǅkBk	dB�e����c8��o��=�gd�3�?��.��E!\L�Jgi���+/.	p��� �ЗH�!3�C&��
��3��I�,(7�?C%�� {���"� �UT�BP�:֓r� � x�'�pK��H��@��\̙�~�!8���]&E��!�c��%z�c�PZ�A��}��.����������|�w']���h�����$Ds��jgψ>,g|(+�{�lk�(���z�\sۿx3'��/K��8�I��Q*���̗�H�Nt\���m�툴�K���Q�q�1���:bX���y(�V�l�p�	g�P{�8!���7ü周���_�9����꼖��h�v(�&�`���L��:�^l�}�/)���O���\�qVȄw�u�7Q��eF�U����eq�h.i.ۙ&��Z^w�{T�x�� �V� ��X���	�Ȣ�k-{�*�%|`�U4
=AN��e�"�)Uze��$�����qZv�Œ�����6���p�K��޾J4�_�����8%����w��s�=ݓO�h�-3�I�>���<,l�A�+���t$z3��ͥ������,����z`�hP�m~���(a'S/�j���xO�y��HmK�C�s�0�N������ �ڒl(�e��Ű�dl^��h�q�����w3���5�_!:vn�- "D�_��G��d/n��&�MX�-�f�ˀ�U�/������By ަy��Y�=|�.7w�:sEI�����+w��߭��agl�G#�V�C&��ug /Kx(�jÆ=ϵ��1:��ہh�3M
��ݜPx��	���O�v��75�ײ�t2a��l7������+�m�%P�!^�_��#�S�B���{҉5m��M���*�Xa�i�](8���b�(+�ȁ�\Vd��!�p�Tn��w��\�:A��e�A��AV>q8H(���caxʙ��-A4�ۢ����! o���&��gu�j�2ڹ�L�#2��i����Y�b�`�%G��q� &A��ud����R�l�K����r94�+������'cz������,���@�+C �4�q?�{{ƌ�س��%ISص�/W������PC�ͫn��cBm!����G���l��3�StRM=U=x�ԡOfeS e�gEؐ��,	��e����i����H%l��}���ݱ�i?:'�5����&7�S��:�e�J��l��M�v�iC��n���1yv��~�Z�4��v�[AHV>Ǩ���1.�=�W	�p/D�xKw�������`��6������i%;۹�cc���`�=�*m_*Zd�G��?����vf�����N�5~��nrܢ,�_���*C���x�Χ���T�cf�q�r��oP,L&5�E�������*G�K4��	2y�x��n��|�{��U�Y\�T���*���Vn�T�8LT����g�ҩ��2.
� u�[]Ap��Ø2���dDa�F)�hV�������||B�be�7�!��t͆V�	�r~������q�N�ڹ�\|5k�XeF\��}(�d-�qd��m��9��9q°݅�?}�'��Sg�%�(c9Gm�=M���k/@������_�Va��;�^���~Aۏf:��q�-;����7Rv�0�4�:�S(
���'�
�
:ж�i���n�H˻b��!�6�hGG.�h�)����ʞI�Z�ۺ��#��_��P�T��LC �̳�UO����c{�%��-%$;��#���ڙ<X��1��r��'/��p2'֢����*�G2'��Hs4�'�ߜ*�ܶR��u_�-e�#Y�����I��i1&2hɠ��gkj1!���&��|��֘@�$�~D��R��}��M��zŠ��<�?Nv�k��ߔ��������,^���
{2浃�A��ޠ��,z�J�WF&��&__���[�u�.4�x���_`a�0o�ѐ����e�I	w��D�IZ��W���{t'WW������*A_ʊ)m�O(�������Hf�s�).�;&:�p��4I��4��o��}����BOE����y@>�L����2�vD�27y����AOGH���)H�e�Y����ϊ% �K>\
dG[��D��<|�RЬzܼ�m����j낣c��)g�Һ�3E}���b�]�P9:S��F�����ߥc�y�슭��������N����0�/zWc�*��o��\��k��[^�tA|H���fw�cT[�^�������a�t��QTE��4�)�q��`W�ɽ�J�(ߍ����zn6�v96��E�&j_��cP3;n����!آ宀A��P�@��E��k����I��[�|TZ׶u��#��U����7��ŦQ֧>���;+x��z����pr ��r2�wUI~�b��3���%�.MT���X�����uQ징oe��J|v����Kw��̹3�����p�����G���8��od�@�,1�e��ڡ 6����u��*�FAH��p!��X�$���?����2��v�J�1���Vc>$�]�o�F���K�Z��N��]�!��N?�$��>��I�	3���a�<TXB�49�l�5����~đ�@��jک"�a��x}��=�}�r��֘�K��'0��q�#g�b��L�_�����]���
�:m�0F>�M�{��7l�roEm��j��@��c@�>����B0t���'x��vՖ�>i|��mΎ���a*{�>ׄ�"�\-��݄1�*�3�,I��w�^�owb���\>6�pE�r��c\V�Ri�����)\�c
�y �QDnN���cʿ��8=����'��W߆O���F��C߼�Q�S��¨���T�{ t�N��T��#�"2Q

�|!���F��C�µju1!$�J��FE�(����)���X���Yf`���n�1��W�ط��I��-�\�{�hO�)M��C��$�i2��te����F��<����a��X\�����5CJ6b���8�kp<��,���=���������rQCD�F���~��O�j<�g�V��H��I��;�_��	G�T�D2�.Bx�k�xJy�?1h4�2�v��{߷�7QH=9��4��W�KΏ[�X��~�x��3/���1_�Z&W1m}YF�j��^����kP`cJ;�0Gf�C��ހEꙻۄ���0 @���
rOG9h:|LT�L������x��US��eU�0$;:�gs?^[
	�X��%���+�kK�����3�%*�5?I��	eMB���=n+91,	Ըu
@4��y����QBl�*P��pE�ӷ���^��_�����?H�ӳ�K��E\@��Y�����;,����7@ c9�i�������OB�c��'5Ym��Chz�����T�^��8�[�q1��:?km^��a�����rj�a�E$O5�%!z#:�V�������ƺĕ�K���'� B1���������c�m���k:��苇:��-ro�F�3�;e5�\.�p2BF�ˏ/�_���r����r�w���u��"6� ��~Ǉ�x�sq��ng�x_\�y�Tj�4���"�;%L�#�����j��Z,XI�]��-��1�o�>�/�^*`#�7h;'��0�Z�j܆�U���������U����M�L���B�]�<Aw�!�.��}5"�|�m6��ф�-8uׯl�'yG���t�s�8���E�<�Z̮�<37Ɂ�U�~7BJRD͚ ՛ PȬ��Xl�O���(#&�������|��1ؙ:�:��BGRM�veџ��<��z�j�D�絑ݣԴ�F��;t�kc��c5����9[V���j��R�~�MO�6źUΧ<z�w�͠/K�[1�%�Te�W�*0�(s�0}M\+o;Qe�L@b���J�e�ȕ�ah/R��R��}+�	�06�_G'�Q矍������\����Qݺ7��/�:�6� 4��f��;hf�����g��ɩ��]�>��6ҵ�W�j��w�"q$I.sa$�CEL�����X�'����p.�(H�.�?�i�C��CD���_�˱���AtQ/\���3��j���[~Op'3��F��O�ɱP0ԶD�^_�ٶB&���ؖ<Ӵ(�3p&xF&��~^����'���Ox�.G�|
�=5�Xl�l����>��7����~��Ӎ�e����5��b)�n�#&<N�=�J:� �C\X��/�����:G��aR��R���z�=��O�+{0F���W'M6o�R��y�0�1��a�t�*������^_�W�����RC6���l��|�IS-��N-�'(�b#���"�ݏn����rEk�F-�����)
O�E�z�X���/eι�#p{|�w{jv�G�A���] "T��Zpl��(e��^b�ƸIKj����#�(7�T`<V��Z�����ja��?A]�%@z�Щ�ݣ�u�+��j���k@6�w�$�W�Y0H�;We��)��N^������f�nU+�W���6��؜'���1s�*��`LyG3a��Ǥ��Î2�8"6i��A��ޞl�ڥ�#:�����vW������ۊ���G��m�.�h�=y��%Z��|�����X�?�*�ɤ%���
�rn����'A7�Q4���t�N�M�O�����LhKD�!|�?��hz �I��}�3~�Q�ɥB0.At�N�+r%61�cҥt��09|K�����l����9�`��敞�Gi���|�P5z/x%�(N�Rg�&J�s�SH��O����sF�tn04��Eُ�TZi��4=������:�5�cs]_��B��΅������O%���T/�A?���6-ٔe�Fio�!A�'�vN��A|9q6?Y!��p	-J���
��x�ⷬ��gv:��D����ĳh=�6��U�dR���X��oR�sF]��N�������[��*��ٶ���`d���P�z�}�2��s�xoՊ���3р�@��	YV��~H�+�	�p��A^ &����sw,s�(�-ڬ�T�pϬ9q�Y�����Ĭ0�|�SA �]N��-{1�`��
�>���o�cnW{����4��{C��Y�\Ͻ,`�d����2�T��9����!����I12��f����1��_���WWN�[��XC�B�=U(C'�O����h�8�
(;m�s��o�ԁT!&K0��E�s1Q#E�D��C���