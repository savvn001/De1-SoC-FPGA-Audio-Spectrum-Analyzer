-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nvp8DW/DoZqE/6Sq+YDpz0Jer/h6bbIaMDcfboi1jkaYOAOAVANAmG/t9uUbvcWg14k/TEzrKdly
ofD6HWy0qlj/pUaRbAO3KPrHtVroNo+BmWNqVREJ3m1UwH4ZL0oZK+OJUm1wQxOzc8j3W2TlDy3y
0aIYD0oNdu00MrqasJXR3/NggKOlGWdLrGyT1ytR455KcuAwautOOLNY1UJvm9iLu/XWlpXThnZb
Dx/u4xJoXT/sGa/YpKZY+aR8UAOf1Wm+MmoTz4/c0LZZzZJNMySf2T12gSEsxzU3UCLqPP2BDFJO
goEzrSqpH7RszgOafeyZ4COGEZQM+FQxvAj0cA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4656)
`protect data_block
6HBaOFlPuYL1B1v7RRp2I51oKoyxc4+6CV/UH7dxmscpwY0wewnot27LM0qJsY8+T69068DcCUdE
Lt4MqvUYBZMf4aAOv4dFiBl7xkYk7zLv1i18MMSsm3jpbLbi2mgRwHRHXvQq9xWVjvoaQZneeP27
a8de8IwFz5tzCMBDpA4XGiYJLvK/Mfb8PqUZtCCib1OryXd2l/0fRIplXffZ5DjGOCos54k6R1Le
47rQd84j7UZmav8i22qKhhbPH/HAE+Y5AtBQaME1blCCx3uWcjqWmGTsBwenr8TEL6S4itUkh2sB
oKGgIA3KlcNyU9EvwoyixWv4gYtZDaV+Zsx2O0dYXqbqfbE4x8b7YKAkxC9gQcBDLjb57r70U0CD
GtTlWSDAy2eO1RQTN+0XQrxfAKodvPZ44IV71sG2ZBmCV+KDB1Rfu1gz8nQ4MevFcpSveWFrO5wK
MJE8+qeMivnr2cnkBJUA+pFkfXSocYXskeg1IL72fs53RA92Ktwpq454qLs95uNUK1P6WQak+hhO
Xwhs0Qtkm+ZrAbB1vv6Mc5loW28HRQSBSgliVfg5Xr9ExT2S2Xm9Xtna1OKOhFmJb33+o9//gIoY
m0colcZy2UUktC1AIOkb57FnmDSfOCwkXlrMO2ecDX47UTGVqOK2Xl+RALnMDnfVrTWdC+EYbbxx
Duhb6yVR2liATglVu44/Kd0c+wcZZn4D+K08sUyES4zQAQ6OKdP4cD8DI0KCkLpWQxfmMX756m6B
oZgnXilU2yZol0fmK0vWZvR/1pg8gxnt5wcn9yC0WQpKiw31hJmRc9YqBO4XppBod1w/BzD8Hcc/
VqrWdb5Hpnhw4llGXGIMqzMVWxcxEDvFfxe36LXtnNfOjtmG7LGwru6uQaXYLzgQsEmoKTre6GKw
s6kgjBRt1oXtqUjXLROitBHm6OxFSYym1f5jvrAdXvlyJsb+BbAGpS0AQsz/r+8O+aTAmjBirex+
DsitbXkkk+uvzjKfr5OA2rjtHnRuu2wZAcN1gPDp6VVK2qhVAlCcs7mB0Zs5OxM4N8zRhjW8YwlC
1BfCKLsVeSOHnhj45oVNhuFUFsxJ8L1A7gCnwFcbbEFjXUNp0N6gX8kGjFZ002+y/uCVCj7pxXOb
Jrzh3roGI2PE/KGV8SmS9Zpau/nnscTTyHo9alNcnJz0uDsGsPgSymSH/O1hkdH8Bd6DZdPBqyWO
UV56xYMdNhEJwVF+4w6FB72iV684a/3gK/LpPF9fqF/vTgsISl9NJAWDo/RLXxsqR9i8EUrxgEtO
QHFoChwwHZ0wSfHHg85VIWqvU3d5n8VfuFDafFqtMmOuhIJ8xf2W9MLfXs/vp/QPCCFXQ8bws24U
871ok2rB9i879ZEtajldmPRxgyUO6G6nCe6U8udnwBZ759AEu5TBo1eFzUqkEDPMBDeFxlZPM11r
WSHtzg8sS1MMLRfzvgJ7WqOQRnvEw2a20cYjYx1n9/34rClLkbEKTe4jFrlA7fGZ0SJRMJlsCMgz
nWVFWP/sugOLeSe8nH0fN2eBdUamBnl5oPZiN6ytMfI5ZUEMY+OfIic+dxLpymlSRhJKAdFpADAj
5AyycyMBHFvtrccgT8P3U6TUKULpuADTbqVSE9vGeZXSRTXxbwYY3LKORSn4cK1HRM8HHqJr6xYB
DSLT3DvH0TLafmaqmmjQqshGG8j7b51HD3YfOrqiyIkQhcxirfwpKqOvmyVvhfdq9jx80HUNRHsm
Jj9yCbGggWQeslQoE9bAzp+GGHENaB75zPLP52wZENu9xzEjJ5+U99fQoNK0O3mvakRRqdeObI1c
dl7i9G8uB20Zl73IjpxEEwFlKiZxjHZJNWT2FjO1IWZx8TvQaJ2vKS1exfU7gjPDDK8VKd+zVETA
7Mx1Shx18pdHT+6VAF0MoDZybV1w4e0GaO4LmoI2zZhJSt2x6uMNu8do0Qo7gEdiRxLwtoEAJVvB
+CjY47qmo7OctuZe2Bjo7Nn1jpPS2M74rb+UB0XSFyD024DTC2C3dIoOFPUPY0LCmpY2ELN09bkX
sfF1lf4tM7klZwf4WC6Ox2u/vJ/L4/5BB6VUUuORYCXplQ2dgLD9AqKWNwakyr7mdCR1l66KMMye
0arezVHEVd7K1RzEauy/EZuFhEx6utY2bmuS0Kud5YjVmf2C6MhUkjUNmljpQmed6XT+GNvOb1T5
ALCMb4sHbbzsEJYPyQaVb3DWSu57cpXevogvWM7U2Xs+Pd3Bz2Oxo5mBvOEnQSPEfp1f4yGJR7w1
OjAEcyBYPKfiV0bFVDVkhoqr+mWCfIZigASfmdgHcXx/h/Hv9LUMhzx/5x6KkPypUPMlP+UB8cUX
hXdW+nuZQj/xCPTrZKNI2/q2XOMlUqsKZ6ET2f+WznRygszFNg5pw5gy29owGLuy3iNw5Bw3PSfm
SgDUIbujdKsjxqZNz5BxiepBOSrikG+eglACyMKXL5LTt8qgynetD41BSf/znnSGFTaR2TvygGv1
9XwZm9zIO2zj/osmy4FFPH7DBtKorHTAzR1SQhBJz++SasuPKZHQISTV9lqU73IjrmV2UFD8zYLl
/JE9fUuA/wyPCeKpqRpMAfQOXb+aT1fF20AkOrIaIDJYsoT80E16tvRnn5/FQuG7AXfyRyXGkIqd
xlERVp1V6vc54a3wXx1dasPWKzDtAVXI5XRU/yDVRNgnjDBLerHSQ+knhoEiTXoSv/BtB3MDmbr+
yrwnr9ifD0NRBKV/IQpU6wQbsO8HH9Llm7gI5gSuPJtxnecDUdE8C6Ds5wmr9MBGaF9MR6p7To1f
xXs6cYfSt/WiWHC9HDtg0De621QowaxwaKpAhQTc7cVV9eK7nTZCv+4bVqkjqeVeRKXRF2iprE8l
dbncgMvY8EyUbzQXdgEuIJ79Wmo8pGUyVgGanbdlBf9XVIVp0g3JbDG0ZtOnh/9CWoBLRLuktJWG
pTOsvnDfzgZmthW5H5LykquXHu1ek/dPLc0TtdngaY1V48ERMg9i5aypSA6t5HN/jpgDp8j0XpvB
KuabipRcENrnuDlKQ3ZYZwepNb9t+W5SV1NQKanwAK4NyATX0ue9IdGGs7QZVb0Nx+Hyvl29E64d
SdyCb9xBRFHmTWNw7tYS4iQyJJUcVqUW+boz/A3lLpNAiUAsmeAioKrVEhwxtTdAPdhfK7d2Mi8f
rxjZ1yD486fhO20XfLJRqVFiZ6ee11QaTMDe5KsQbz/fMuWCUgeU5EAeEkxDVWbPIUhFsV79HC6b
L0UUdRE+P73ODq6UfuszFzAl2poeOtwfq+vYFzqaXzA17ZVsszCKODhJwyogKevLoryLcO/hCwql
7fh7fSieRFQf05Ch9ZbQtilKZPy6/jRORlJ5oTkUQ+SjMRy4mgV3GXKanUjHVFg58s3L1gqKPTY9
ItrDK5R81BLVmw5T1bxAKyJDAGPFYxeiFZrMNneO1fiuirdalqMwdHkezWJwYPhfwBHx3B0Pv2du
uQHtUZYFdsL2MV72/rHSr/ltxgNdZa1O02b5J4GSeGUHqbkoNVVhMGf/aEFxwdcaq8kcM4ZdsgpD
oFMMHVHthlDOj0ZP6vppaZVObdwbvfcE2KePJ9QoRP0jtznzXjADNu7UnFhpYezZKPLqm9PSnHT/
tIOBjPadhtymJn3JiFI21Fc55BX7eSq54sB175CW6w43rcUfuqqCFA+1bWbnA4CiBFL59Gv/fsGI
LJoPP1ZOStTynxm/BBbF8JHawVR7TeHx53EehhJVhezz7DYTeJ5Va9iIbdsygKsvkELl83yVxJsv
3aasdOueZMYYhz+BouCCu4oQpA8UYIr2SKeWEHgqrtb/+0fWbhAbR90ZWKAky9iYSyLrAjAN+MKW
1OOsEXOC/nVXc1bj68FPAi/3P8nXcalvH8WJ1DXD4oTr4wuJS5PYN9BpvcJHJ4BP9WBPrnwteSaS
5Z87kpMeKn0hrlJUMDth5OWzI2Yc9rVN5hXP7eAxvcBtTvcFsImdrkqB+3l5qQQFKH5uMKUUgpj6
0AZQd1g9XcWiI+ANbdpxpmEEhvciqAwTh14dfJqDhZyGY75mqlO4IUsE+2ImT8ahohlfxSIqYCwb
omaLmG8dv7OIGkd2mgmogFXIyhZFJUwY4KMTp6EQFyV555GW/zovulkDvkRzx4JHXXQM1IQADArG
J0LbqC+jjdPk2G/lA1AVRjbdCCqZBARnOP5gG1bvbf6NHUCimFBW2XrXDwSAHF54RrtJlTs7RKUN
SiFefIeYArehxga2VgiNLyCZnrI6ajfcIecAOkVnJzHlhk5UBPjmjVkyLadPeIoIfPI1BbFpjFlb
ykld4yT3wARLZeJLoeiYCyFoAlxbEdUL/v4uyH4rMbY5t8U2g0MqG4RwnS+wsZu/LejEpKpuFvUh
GjJ2gP9br8ryJlZYEXbFQfF9UWy/mTs47aMNSJUhLgn0DHLpfEhgYAVqJ8rgaby0tEZTI0kpcJ7Q
fmRHiy+0E2xeCzR6kJaZ7ZEAlbs7p5rHsThCeNELZGIUEBkXKqo952PhFv5DK+XbLRtd0FqvKeOE
iYnxSL+nc3/gbcvIRx6fhFWANud/zo504wPAbbwUKyrdje7V3CBtvy2MzYH879MQHWxG84XcUiJG
crGQqZLHsojBjbd8SU02NcaXV3GbnTVFT9YPIMhI5YyevvDbPc+BMCjzQ2mTYAWeFFZKLRlBLXyA
KyYSPocYSqAvWM0Sh0zjrEdIObyZ041Iow8EO7+9E/M9wFf5Q8pUt2CQTr9nIgL2WOF1DRi34YJc
2YD45L7TfeMGoLes8/0P3HM/EjXMq+VQSU7CcEoa1rSmXKUlkn1DYkSdfY3Z5SPQNEnYHVtlxJPQ
qs+LLSmDohN32CLXEIo4qVqZ2k/nOt50xC1NOFlCKlDPrnZF3rSZu6lI4ziWedT4oSRiQHwrGtlF
yg3vdP4IuANJWf5JK7w3PNo0Smhnm9+2IJdN4iTKdC7bt5tKR+R4BOwdaHgAc7C0pEq+qPZewSFa
DT43o+mEXKTMFW6o5h9q9arR9dKu3ZYRf6qWCBneF0EhNawTlfzVhPqIDi9XyQSAXnlyb++O3TQF
ooCyEHL3iyT18So9IbK1vdA7/ZuCTbAXdueA9rFJVEvHWf/p/xows4uWKxhIYfM41M7rVMRPoEXk
QLiDNVdYkB/nJ8XAj19bDLEheAdylc+iT17QBB0VUnpn/SyJwY6GSbKmM/2ednbdh5JcRCog0moz
CPjB7zcXAbkzQHsAfvwt8T/S0j6tX5BImTY0lt2pxsbI3p6tsDdwkIZKUD8GjeOibzZavDWgZAlI
R8G6slcCcBFx7/RdOQ6VpRgnhMCgCh35MblwF0L+nqQBpmJlomMsWxAoQaV7W4BpszGLNueypM9u
QXLo0+plExMoX+08vY1HMwHRwqOq2/toZkrEleZ7GbFgyP8vBuyYzCDMMgD/LK2ljBdbWjg3iEtZ
LchkHuSeG8ILtFIal9ZNwQ42XjugSXoqqgqkrh07gapvpdz9uL1ZiqYY1GGk/Qw4TqfCy+HSDZrW
kf83LM7rdaxBZA1yy4yg45zQWQRK91FlzckonJuRot9Qe6YgodYhEQ85Qt9blb3egIzE0FBDQLsa
HqllbjBMzO3SWYg08TUcjtgg5Xwxb3XwXBjYGZ25s3Xvg7nFTG7CQ1cvqVMj5xHL2wjzGvsXNOgo
gjZYkxZ5uG6Lh8mWgFptaysGCm3mOrIhBeXeMwz3jGjPsxxCF/e/t5X9JmajG4K+/vdE3Z7BdKki
pCQzEocf+FHNcO0VNS3Aj+CZ6iyA3T1foDbkaaDHS5sRSsF0EAphxvHKkhn99fGkuOxbUKCz1as5
TcGJoUdnhs6XLkzV03ffOToQ+OadZiWkk5OjjQSG1sKNXQyYy9bQy0DmaWqY82F0sz4Tnsnm8VEm
y/ksy2yFkSykbSECGqg3TZZL7PvbXy6DdJ1zVf9Wmsx7j2BeuU7Rp1tFYEZVMrHRUcSHdd1iHzQM
OKEr8UX8EhOxm/sCoFTaP8uYk42BSGvemmkO5XXvNFqdFysJ+tXyqG7FAYhljm07OkEHxU1y87wj
pb+S+q9H6Tnt8MantIgV+VMS7i7JwCxgDYITyqnIY8ob3yyg5drXCcFuxmJyIXv7/XQMtPs2jyg9
ljpKVU++Yj0hkMcT9e+GGO4jOXTNFDKQHVOBQbHdPgLvdnOUgfYO
`protect end_protected
