-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A33dEGZApYuBR+pFbMcKaDPJXC9f+ESP4t8Ni7Btxw7UCDRBeGDJGMQ+yi+wj7e8dR74I4STDuH/
D1jTPTVDcSmNBSV4Ls0qg9fNKXhxrXTN6DrKvZDdOcZNCYvZ5fwhS0xnEvafA0nmoJkV9/MxX+Jz
Rl4EN2HryJ7SxUyswoVxgDqJOsDX1NJ6hXuQxJRb7bTMPHKGLVyWWYf+X4XGPzsLd05O0mu4Nim7
ivgyW7Tci0eQB35qoviBb8qMBMXmtIpksIC13+6BSU2KZFDRXzP6s/7RPBMazwgWx/m5KPHYuu9b
PoX92FfGLdLHBvf+dGsSZJPKgqTfmmNn5nM4UQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
cLVjPfTfmQCU8Ju4lhXZdiZjCop7s75F3UF1tf3iWm63kAu9hWFm4OUMlJJIy081IHkvRyTWt6xN
Lq/QVddTj8ZsMmn7rvONkbjG4DQ7V9KeIxLtS9Sr1sRdGNFz768k8Y8uMWx/RUoG92xx483q7eST
5Fo4S7odo9sjewsaRHrWEatgr2azEC5hXmPsn5MaOb1ZQ+LoIYjp7DSR6dZXhxOTKWEC4dsg72ID
dDleiZ0c8vIZRzf93DVyeYdCrtdB+l4X2Qb2fBxtR5hjyZWatYylsa8jlf11IL9N+1rrkvZiA2RN
OcBYlmXfKV/LF9J8cHciJ+g/b/jg8u1RhWJtLF6T97P42NHccLuCzt9S7qmrgck65jyaFA4IA4Uz
aW/9XO7CaXoQD68zqLa3k+8tljiQciFPj2zgNdMExTt2xDU8uTC4ZaaI/8pqqNbZTcbmGqebOYa0
/QpnY0k1k6WdC9U7CaEV5q+zl9SehET0BIbv4sTakACJS+Uow11RZQV8D4sL9hc4Pk6DE9cnyXeh
k93fGMMToNAXrI/NTZTOnDc4OKgTUKWJpnT01cSE4W+80k1UppB0J29C9KiQcbjXm5P+qfH0Die+
VFRAz+neWTXoh7MEbKyzf0uP28jYVTXpcHCJtxDTvfSUcAwWOWQoMBM8wO6xDkzLLV0RkD2b1q5v
zgrLHuyE1xccmmWRu4C9PP1PJ5YJIi2nzcyikZJItXmElQ12j88I1l/UdxoUA1FyQl80TNWujkpc
A0DciuN6IpYOVdakEZkQPMADy7zOi48n73h9BZSwJ/PhioOQKb6U6GKuhKIP+crvGDPLMCwIkQcv
MUtuPR2mvWR8vjvk5hq0+tYq5tgg+id0V2JTT/VnGkHIXh2CLr27qR37kihyEEh/ZrTS/53IMt18
kU8cVS2meZpgwZSuxVlXrLqOCyOaC1xMyJdtfqUwod9stAxswUxguieOS3PWCyNSunPcw9HUf/OH
/HUZ25l59Y/TnqQPy9+O8aqgjYXc3lvYQq1LTAnJrZle+LdcgR3zLZ3Gwy6S4ytI4BnYa/lnLtFW
PJNysCCGlE+8OH9dYZ7lIhwaY6pUp7fR7zuaBu73qysXgf3ut8rw4JOxCv4ZcH4s6/yS0FMmbdmW
IwbTrisWki1TjQQ/cMmYX6Efb1Le6MeTX5ZFuDaiyPs39GY8HMz7T4ZvXmTjVyCuRwqDA1tYG7sK
D7E0fcGir/xjq79anPY0u3KBob8ZeWtjdE1yI9XoZFK1tw5xW7QziuzeqzWG1NTIGc+egvpOIVRR
5A/6XQvgUbAkFNjEb+oHrSWfrM8Uye90FaVnR4WQ3MuC6FDIVCF8RE/nDWcCA3C8phsW0TyVWbuW
Q5DF9OfIiRtXUP+rRfncedArYkgfK//hNJVXgo10wUrCmd2LBn/8ErC4QwlhkSeGSFE/8o3IfRvp
e9qSQ5sXfHAbdBfpfpg3aYJ97SV3FSD67le+3P67oI9ZhodqYSoUGMyXbdSUzFMDPm2SfI8G7//z
h6f8jDddN8vnYsb7bkiLBS3+UaYG0ril7n3KQ4E6dEmOgVttZJwDqmJcufXAIHONZtjZPl1vepnQ
evlIEwBSkMRcV5F3zfyZPaLNLtOxkJA0Hgey2I6V+w6EaFtuc0FHmAXBYdMjjLDmxMNIQjxRhQe7
SvZTOOReZuh71pmcUg1L402th2kB0hugWd+bUj038mijzciNNjWlHcma2D6aVO8koIP1CpYXxphB
vFEP4DEHAlBYrklYBkAEzo74YmeLhNx3OzYeBosRgjTnxyiG2i1qf05txKGdvHoulMkOEnO9VDX5
21+kYiLYuxovITOhARAiw4HFYFzFrhWutUtduqXZc5CQzxbw9vF1ezVTWi5ms6X+IyqLxUId+Lt6
AJF71wdxrSuyUT2KVFNYrwgTBbOBSAt5pIkNqSVvFEh+lAoesBnOi9qLXmDNo/u2W7i5E6oWrxL7
WvtHKgOBqv44Zizsw1pHe9vyLRsZ6z+HivrssAPGHmdHGxd4DlRkqeFgLefGme5AvMRDmLXNmxzA
mX78ewEpXbQhC3stQcwcLxcGcNlG0t3TCnLjSTrE9UEw4uhgQBy00AYjeyBSM2pAcmb+IpzOr4Lk
SgfV7cXQhwUC+/KX01GF0qBHu3UmZZbRu9QZPWZFVgqbPHbMKHeOZxvDkpWRkU8MSSRg+eU+2fMU
Q1ry8MuszkSFNnQO9XbdLkNybqI8xsV2X9u03zv39D/4hdARUafzuRSQq4GYcVNAjYicIm2Wbx4q
huwdydDMq5MCeg8gnu6QsLICWa9s2hpk8uTxZ2QZ16x+noJubr7nEX5SLILNmUld7QKMmsmiq5Gf
/o1H2DaP8WWfL3t7nhCwq5xzcfoRUV7xE4zft4v+i0MXGfjNN0WdPTCYyb6TWJT/EJG6Gjjk+SSQ
4bYHGsFggnlbUSFUfWaPz3zSYKgP8Lzo1mHdSMJ1e5k/98ZeHtwYYBgFviWpRa/bOcMlkAiE/g5O
18NNlYFnBwwzAL0gFBoiV+MdN4vqThWbiCKrg4VdBhLDVvUQOH31UMgnDq2KoMVCzNhoFMhFSRQP
Rj3F/xSidEHycN8qEj30LttEIKj4n7llfnPpK4KyO/FW1wifm84TTdzvzI3S2If06nyuwKlZvcMf
/MhpJXepAoIV+UqHuAjfiVT4MlISzkuucgqXtay24L09MYxp4iqR4WSQNi90hP9RNFiTsGjYKQO8
rbfSlx7AsL5jWJzI02vWx+JvGf1HeiJcqgBZI5w2RnxzHU7YGIXM514yZkWJhnAFgt2MnzzOxMTy
Va3xDK9yMlIWCNQHkwAaprLNOi9ahBjLphhW3Rl0uCKRulHiZpvGO7Vjko9Om6J7hPMBvT14zNLb
OntM7RojMDKAmqUgYqDcRiwoRnBLurVQKZfVtB/C6CzJb3gagE/tpzX8XPf15/baue8jcTU9BWAa
0idgD6Psr89tju0IpBkOND9Wpz4HXjzExIeSfV/6VUCtikazQoObscMadc+s9/bWpnW8nC162TO1
toRLcTNTH5I7yyUphw6szFRRfAcgituzygGiN1An75Efwj9GpPIwtGrdvdvhAxGbZViVgPlQKfZ7
vDOR5NAsu/UKOa20UGQbhOUau+3k6gZpqRQBvG/bwDXgWwPUSwh6X6991fn55Yzp9XYcQxf9+wrp
qo83lP+kgP3vcbIb8XDaP2dt9rZIYEmzdAuxJKMnQJUr8+fb3SeOTh+g6FO8WFybk6/Q5msCLIcZ
pUUdlAuyps7UIB1uNDQRtcwuBlo3ViIlFw4tBnkLVTUPdXR56SKx3pcX9g/jJuqTMHjn+4GPRRzZ
eA8sm4maWRXdhf55HDbTYj+XN3GUUX9DROlMhNMPeDuuQtog/B8MFVl2YIigy8POeyxmjuQi0siN
fC+P8a/FvjeBUWLQb3sF2h/oCxk5n9WnKWXxAif3CPCgHkXy3pnOLxO114UM+bNhqjeB4PctF+a2
Zrt+zVkaMvTpORjMhqOo8Rb4JXMv4skhyh2DOJNPC777LuAab1UXorPZ83+C2Kf6zS1gMFB6r5vL
TVN/nYixOA9Iq2Z6CM1Xns++OHYAIOmoYbmUXNUjJw0ktHyb7oPAyRNTR5CIXwNT/D6cCxAQ239B
m+jfhmMxEvChXGJ/1IfIp9zpbc4G30jJ4w1L28VvoHdwD/NDzBBjtSCI0mIXejMwutha8T99VCF7
z4llYTtIi25UDi4ta1A9qwlBKCLjFViwqo65DZGKNO3zHs62iU+rtF77k1Lns8Iay28dxIyjNk6c
GpHQQ0L7tFILQWGB3uRrPiucux5Uz0CeLtdbZxW5f35vcOngtactosJXgQ7CHnRucuKIlyePNElN
32AI2jcRPFRE/oCecwBbzSZbI8uFamyrQMbWSn4KTQAyom4XyBIvvdQe0slg1dIKRylyy176ONN2
u91qV+JoAYSfi3qUMChEVS3Fut+T79W2D5QbYNpTLlFTG+5hu7I+LBz/Ge5XNnbJ16QMA4M+UmHd
U7HaRGwaLPKSwgRsqA1MPg6+yUenXQK1ewRRhumJjln6A9Mk/O7ldAlU0DGmBiR37wJc3c/j3ztH
hfbXPicKkUladJME9l8qwTdtDIWaO34iuSc/dx9dSrA17+g0+vU5clLNY3eXxaoyyX2cWe1eGrfM
nNQ+t9iTYOqFJBU2iugUW9773bEwcvPmRMrbItEd2lF3TwecmvBijaADHoGZ9R9d7C6M1SZVvce4
Pibxca5Z2l6ksqWyirgwwv1EAqL9tqltrZVuVlAybGJ6+ZDXnoZ46H1W7tTdBcdpenWAE9BugFa9
1p9k9W+Dy/z63zNictbi51NXzoOZleEBwiwc0aYPzUYUrgF+blZWSPgvUfMxL3WY7faWp23b2AhL
CC9R3qc83joKscjnokDebqgWZ/U03GY5aLrTCypWxloB6Pb4WzJjWWUrAHt8tGnBnXstV4k0XNNG
JkpZXBFXEWqGG9G4EBzONEeWFy9ozrld9X8PgQabaY0ntuSuv7XYOtxXUTy0FJbib/3ky/qkm+sD
FU0tZtFYGb//zSot5nRF+I1hnApRnuPRjb5WwymezYxBf++a7QhwpGBIszg+FFYr6jPG97Sng/hu
Uk4GPWJexKCM0M321SY9hABOW3nCL41Zl3vd2cz2MsIwDkgaUt7HIElvv6X0cfDvExu24Lh6cGR2
eMimzBtkygmvMHYAfNXd1Dqn42QTGXoUfCFESubCE7okLxXfEEBC4Tkp7s96ccYcP8GhW4zwNtkA
dlSIHBx4OK+4amO8veYmJ2x7WG80f45nUaSGlxgdBMAGhThj2GZp88rVv1Q//WQZtJJvPmPnfa0G
e8DgiQlpbRESdJBPJO/jZwZz/jihs8VZIuC6OZPzUrHscP6sFiKcYOh610pAttJdmMOOGbJ1LOMV
MLsboDPBkPL74xCqWhOJCh+1qxD+MMU+GfwcAFzhpChBlIQdJ8N1BJECInxsfqqU+Vnf/Xd1WPKK
IZNgOnNUPxu+Vs+ssYASZ7zELhOHx1oyE/58ztHZhpNjJGJ7unZTKGsgAPFTfO8Rp7b+lZDQNyXG
2v0/cfSblDMvBt0d3pKF93LHPdruQWgqIYOuKoCuHbxJ8kwt2kWw9/8cNYHhANCWX6Q4nn1dUrQM
MMCcx1ol72Rp91c0suwovoHv/d2qgZaxefd9BF/T1NhC5jndFSUBFJ35oeRUzKKEk5awpuef75ON
oCzw7D7BIrMx6Gg2CkhGeSQdCJh3L1eJtAY1Cr8h/uDE4uWXeIJetVjDHnDppa0Z6CU3oVetp5ob
0KMlayYvT3M9SMyGimDUy90EarXBSqo/h0pElhaFZbn5ScFwOHhl2Y8EUoh4HYiocrZUyKuF1/GK
DjnLfW838BqZ1XLYhdqxcZO0cZNaJDlfHT74PqItgBQTnfseEUpeZm6oxPdVZrDBZ8k7pkfBcqa7
yldpQh76BUFZTCHmiQpRMegUSYMKEnK+YGKGO4L/1ygD1H9dEGy/UrsqSnJqK9bBfvTsegppjq0E
aBc1YCGhdERI8557SRJEBoyNSrF8zEKOA6w9xv5AoPHNS5iRzSfs+/89TTErAF4DvNn6E147MaSq
seiGG+X60lmwec0nR14JzxG3cBIYccarh3wwzfxV9lg9VKGXrAfi8Dxmfh0X4voeJx8SubPrud2e
B6TZl29RiCLzcXUjVcKKNC8/Sd00shmMTD/x8YbUFZ1lmwShnh5Oiz6lums4G6OjEvdVR8823aJ/
vNgcQT2nSTGoT05lbXYAz7BNxuT8AIBiCZLzZoWAuY3yXezQHWHxOHDG2eepeOZNJJmUO2YSXxtF
EjH2ABW/hdXluZL2ItJGBpcw/rdIQI4Xic8Wm7FsUXO6kUodEJK/eCIOZXP5IVE/i124CGUqSoFu
JJpMG4T4xVz5LsmdUAjwhq9EU+vv6+mVgt+rw+7ZTmPs8MmcxGmHXLIjuwUbDcbqZBDEzCw55x49
5b+/b2ooPc6CiPU7Ehv9IB5kR1M2eERp7RNQyh1VNfGLDXRKuRquWYmH4L8ZC/ufLHar3kypbKCX
Xn7+QKeXAbyp2AMtT1KwZI1F/UhE955hVvoUS8P6i6Wp2ApgysbsGQLlBruXzgnIfTqE+bFCyozI
jbAAVF8wW2BeGI0pkFJTCW3Ne/KJXqJBJy8EyPP/ZmcrruXwtqqnaWXEuus1JLNwU/+0qf8EpA==
`protect end_protected
