-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
r+Hi6stulRSN3+4zPCMMPTk2OBuGoLXCjjaIg4viuEhTi2FBPswJjxqdeLQVu3+1jSeWbCZa65V6
JulR1Hb5d+g3IhSpfsB8jcDntYFEZcXNA+ZMnFhkWBNMAivzkBI4EGGYqYiJuQlIWyaDWBS3vID0
KMH8uOLHknJZnD5daL5ZJn7BCfcOdtNRgme59TcgFCmnexKcqsmQWMzXTn+1fmJtXulga50DC4Rv
eM+zWxzfTci9JNZJQs1sdRQzOPaxajJn4Fornfwe0DWh7XGBuEM/liegiMPvX4d/8bnqYRqqVb5w
T2rea5yQKbecYI/ku1dTKHi8QdtZ/ektdSDDjg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
ALFDQaUZ2amul8zH0Y3vjKLHWZOe3Zwnx+w4GcPSuwV5QmBlOKs236lygZxrp1ZEWZKs/lEZGyXH
11sOWsxdUnX2Cn9aCC/XbZDW+aJ2NO8aEbMAJ9pZaG2CEIJPPdgpaFjPwkjnhyPCa4YdPEJ6mxZX
cvZNtLb1/JoQb8klVMfoAh609gQw5J7Rt9eVvUolwrfsC0DHFHj7ldc7ExHaUMjJWme7k5YNxXFn
nbnKOtm6/nPEkfiDvc63C4vPN8xKkm5UhY0NSHsZ/gCZ/nALj2ZQH4wCJ2A1G/newa+Jrg8plFhE
MkyULCcI10MDt0xt7OfZamOPVrfLA/TL5yz8xEtwEofNlAgpejacqvzFArWgGhW39gTaFrJkmZWM
CMKSEaN7Y6yldSdzaLSgQwk6Lik37muTNmO9l5JCJg0DZ27xbiXxBAdZKhmZB9gXishGWxKOwXKx
G7zjecR59jp/xdVkckbpZsPO3RRNod5rTJwEvtn9uV/uhaGKFJGVKYfhJMYkaOpiHFoZp4GAarJj
k7z5LyLMSPO0taPq8HwMIjT+Zi4m0lGsf4buagkaQH+fwBFUhFrSopD1hhRiHHf2wsHD/cJo6mGr
YMpyYkfoNSRAd/vB2n5q4N+wOeM+CHmGBvn3le0Z6dsrUYR8RqZ0xYG9Ix3c3y5hsUGWkszw2/54
YrRtunixD+Noy7k02LyeVU+jBuFPsOpQkr0sNilCVJpF4nHz7RJ/OU7hzcy/IS5JltWrMwyqyAyX
3iHQ4vtoJWt5GBe+q0yQG0vDHR9hsXDtrmUNNE3C/EuwNZYcAwApbD0miYuBVoaMxI7k5QJ1MnX+
JewwLbGY4Rj+PTfj13gtWX+hK54NyhHw7lRNEulSuetSeSo939QterCord40LxTZ+DL+DeaVTaEE
X27db4JUudVj6fwZBwlx2IkDXsMZLPzyhMwHi82NqvNEbxW1laXb9NeSrXMpe39dYUUfFOoAchUA
jV/MN08aVFddNb8ClFNTdX4nhSCTgEQMPj3gsnrG53wLLgjLqtr4YJjhjp2Fy5clDBeVvl2CKHh2
6nUSqe+vZvrXPJu2P5jHTbjYYy8UC+T/XQtFdJarVRK3yljuwG0nG7OlHuA4NoJTDgkxehBDxxZ6
gfs8WQIfLJxaTUcdeY4dJ+PkUKPk/Zjbd0LUiE7QhBas/y9SiXwxcqzcNqJRNxI19QcrDzoFaDPq
VfhRU44NLp2rMysFNhlTCTdEKi1a7r747T//TNruZHk+OJ7LmFjlK3H/bfu29wG2I19kEVk69xji
rO5vQ8Gan7aWU5mZs+3s++YtJVxGbEJvJCY0PgL9iC7KPcaZhU60uTZf5Lmo+vjO7V6VYrf1v+yR
6L2ZCj8InF3VDdnIxB/STkE9zDrJMLhAy2siElxSnEYyr+kLi22lL5L18vDDq49t/BWIp1JluWMT
BJm13WKUHf5t6BOrkbrsLcwduLL38r3BrYQ1AUc0FV0LG7gAW3dDCJFEbf1QFhV2b4te2C6EZ3QN
28wH8+qrNJlXOnAwY0o50dKIwwgTG+rDbuunjq6VwMCZkREbaznWVpaxgmJ5VmVhQd6MkAkCxOZp
vQuVGlPQRxN1EdC3hecse+Be0y/m6wFwvLxVMh75I9ZaMacECNh+jin25GyzGKYZYf015tE/9iHP
8EmL9LV0c0ZiHhMPe9sjRmfUO5LWKsTJBsRDpDgZgbdTbfTbw7VYtPYwCT3XS74eAG4YzzBaaGdU
D789gsUsETlo9+7I4T7p3q0by+bGPjYwSnvC/IMpPaeeywG+Plev7aaWuHdsJxPKnpvt7AvOtLrN
JHDYlg1jczDc6zqFJInHvNiXhj9DOvZO7rfaai8nNeDd1/t2AoH1w67SGbessTI12HVWKouedll9
zAo/LFk8TIneE3sJJm9BCUsGLMjTJu6rEx1cYKslP8nCdg2q0WXT9W7XRl3FVWjkexiXAAAp122H
Ad0ADTJnpmTcFixGJWQzjPJaIv1JTbm7tRvEnGlF5Wbj/ulHCQs/wOQwIm/BleaQckpGzl5lPrVz
daJdteqaEC1Jl1GBoTXsR2rplvrPVxUkCoe4CZxVnL7SACIgEVJBloCWAJ3viiql7K76nKe92JmT
5j/2YAPipytoQAtbghJEKG7i7HE/5MlWTV+R8yM+siapc+Bk/dERUJ4Pjm572t8e3wAX7lkjkKJA
wC7ANK8yqgkMtpWSAFBd1m7vLHypmt25VgM4O1W2Uk2+jycmK9zcQboLABKygfzIFdagZhalAR2k
6WD9OsnBUHMyK+1chrMLwiThGtIWN1FbI7KaK2adYv+wdyro53sHXEsln00TzCOzLe3loXH/S9ZE
t4hf6heqMRD5hECNJ8fmNpk35fFWxceTOut3ijfZZIzyy4F3ArTyc9Nn/9HvlYI4R4x85Doa1Jag
FWIxpaiuVpLeYRkucF+f7VQ2lArnYtCBUPaKlmOjdrGfNL6TEjZVBgkD0r3SjXuR0inCw1mOLXfv
HWa6TiyZMu9knh40aSRjP3fWWZMcLZ+kPHjsbyS9GNEnmeYQGlwpG7SB5GK4ubDjDn1lnUrXQF5b
Mqn8KNoGbK9GEW4CYRTzgCxeS/2eYmi07Txr2rkBK1Wepmv2Y4jOwHN9fdW6VKBVCyy2MmXTiVoX
38ZV7OIYVnve9aAviKY/gf/i4mzBgImClKoPvouDZ7ofvnE/0BRkXfkbMN8E/Evvsi6DZOliLGXY
FV4wV71oSJLGLSYVLjRWPzG9z3GPE82O/UfShTRKHQjnPbBMhPHofcGmVxYN+1gGeTZSIdUScQxX
HIIDY275H/Z3IHVxMvlGYK5/yPGj6W8RZkxWT/IW26FJnyRcQpPkGDc1GzD0EC7AaMpJToQY4PXm
+YAYubJWM8f7SoY23KbksjEuFwot+OLHtWh1rIUcq0gEI7NoOlPq+D70Z1rYXoRB0xkqMdHF5rHH
dBDYMueMLFfhAkuB1MLw4mjvt97gLqYQDKs1muYhWJzoyK5zNcjjA/uxEEjtX7doq/BBhGBfWJwO
YFkCL874AUDmXzpdHmfJHwy6wePLQLqBz6/GtdmkK0SMlOnViDklW8w0mKWd/kcQasocCRRPQ4xs
npa3GXXeWNee8vIa16aqvPwQwdzH2VdmUKQ1619Lv6UDHoIx4l/WXRIn5oXkpjWtSQzTg2e6kWKL
6A8vZZFFCQHAH2fbd22g7CFOhZh1WJ6lgV4lzpCYy2K//IoSSjqO4SDrOGpC06Fkw6A6S1BcIYKu
vXqS6LcnM1l02l8XJzib0t9p/f3KqewYUHdaZG3ZRpMTThkb1l5+ERmyQX7sKgGhDmGlAs0vMFA8
816tBEw7Yj4XUxx9dKFnq+WdGvOpubzKA7vwlKuD0OiB5bspbODCZK6h87dhmJI5rl0Pm3Pb155b
XilI8fsqdk6gPiQ3MVJUaWkM34kpe1mwAVnJ9HVSiegfFHUxwyJckAA8xe4kVU6HkgOAsUzjcWQ9
7JkB+GjiLPJYz2RtfLoNyHKVvWh600eY1Z9ae/nivXSbjdD026H/SKcapOpcnfnL5Vhbw5IPVwa+
MWQE4nnV/4/Ea7IoxcUdUXc1Crop3/3L61Hr4BFYGzQy79pm3J3p1X4C/eRT96m7RPBdbr6fQxA7
C5FvKDfr6zLB1v0eLhF/wXbJXWjryWpniT06xgN5RsYaUgq52ATLYqr1UlH6LUpp+/IgFyOtbdE9
OXD8DCXKR8tCgjHV4LugZ6UstwpmXnDQWaCdGDHl7afNMoivMid1PNrTP/O9Wngmh4TqOo56t2pu
kIgaSDeEduL840sqb4N4xh1D2LjzeuGNzJiLIS16wNydEeSs82bbt+GN9xsVm1mPYbt57O8kv96j
L2ZSgZ2zievWljKtDGOJRfvicWDy9MOh6U67l9h6flt2HBPShz3LuulmNiD9JjJUn3QDlJEp4XBO
nsQ+T9SdeRAjSmY1CNykBHzo2fFw28CkpOU0Ijic4DBjbqR+TK9hM/4UpBaAyblgawcWZC5YOH5e
bU6ee7yBr74fUsDWfUB+L8pRMZc8YQtjAtaBkaKm9VzIZZZ1Vf6K9eySHa8egAH/U6X8GEQMgvAW
Tga/d5ils/w2T2Yyhc5gXe67MRhcobyKWIlH+MtfTKX8ZqK+8hgBCXif904Q3k4qRskV8w0pCO8L
8UPuRZTeFXgCLTWtHkAFRNvEp7TH0nVMOzXHmAw6VHCjMvYqAYVCFrScBMzeCD4Gmt5+vG8PTZlQ
bl091AFbh4tLcmF4Nsiynq98t7Kx4Z17YHSdGOD+ID1uh9Ih+DcIEtKH/KoKZ79sBkgdhJzHD685
6yGt26iNzqO2SLmMp1Q0swL8wisotn+N2JIMOjAZhIOk22e41ydfQN6jb6IDzGh06QKvC/o0a6de
5eUfAvBm4cEKckRK43IiF9Dc4tGKmW+oys0NzVaRtgRuKg4c2A9TYAn5iYpSGAUr5wDgEwC/0Byv
YVRH1Y9AQ/UjoCJFMeDi6ScaJhjq4J6wIHCp72hUeRWWbcSZmjhL1bvoBZhiZRH8b/83vWs3f4Kz
m9RwIhnxPCICuaPMBc5aUIXIqZ/v+H8eb8ZXN6p1XZr+R+Ff9xZ53M9hodstzv03rusMQO9+MiNH
fpmZcqomWKaZ1RoWxrF88kmupUlDFwTepELVuwI8KP22+9qRGrDGfXvWmUQq/U65hW9hhnZcfix3
Xs3+K7lkTQrG6YfjIzmPLDWqX+rP2NdxGFjsE3KsRzjKH1o1oiZ2dfu/zqpqmTx6AwzmgDMmusGN
AzjKB1TkRHa/14+eMSBNNtby2RQe3yK0j9GCbA95xO3xY/4b/FkpKPOk2LWKNx7jgt5SwIL/IYWo
vqThWdrw6c7hhLzUC/SY1YbjIFMPMVYkX0eqJ4SgLNh0E7syd2ED/ipw2AOr7j/jrC5uF4nIBH6Q
Kba8PKxC0ECIbTmKvFF3rRr92nsawiYXURIxJqW+c8bjpJiC8sKqd21GIPrfZbinOKP+PjpFb5aM
A6Bl8tPOzWElNgsHOcbpACE3wNd+Q5RjjDhIiUZeQeGpm8TRG+dwFaLJrGyIvfI3D5IMVt/Zx8PA
o+qdnmFntQRFYb9Jr9BVdd8TVd/ULDuqgZr+vIS8JVZWBhiXD9jgm5wdtitRbBAaP1pfVErLAQHw
AdBF06THC8WzxJx/a8xHLgQHCa45HLoneAUZyh5uhHim5TF0/Vs7dXonUC4wOHLlo/No3EB0bSjJ
FBJnFK+tzR8RfFPyQnuB7a/vWuB+pVdnbdhy/3sNcpSZHegfEyW2hjAKg/I4VIqbtGongrgvOSsv
qjleT8G/e8NNAhIr06S1pbru9gSo6c5v7SYvsqEOsZnQhnCHQGGv6fVkv4C2PLNEG22pyc8hbNbT
Yzn4DUUfkf11YUW9uEvve7cq8jHcS+1wrfWilYmBgGbe0HA9FYb963ca24edizO0dSjImo05yqrE
I7gFbSbj0dPJnSuzUXtvkGgOKFZAVviNX2OLSOqQRwbx9D2WKcOkKZ/mraYLQx9KXrs8jDS7st+f
lMVNQUDopCREKZWIqAdXWZV8P84aDSdTGetdYCoCZ0IljnCMxYaTi7uHsQX+dHHYjDxBmjCPokGc
SHRvxvRR2CGHGbycaauXNSr/vvbxtLrsiaC0996VmlcIXhfF5PJDRh6RSbgeqX3fqopNnVv8HINQ
Elams+vqP4+Lu1Fc6rmym+RY6/Jam0xc5Fy7LlLE9boX7kv7Oaay58qaJEfY8yCr/sNz3DmmbS2q
qbhOCufUGrWXx2NlGkxx+OXHN2om/2ICoglZE1qqqC5SWqzcxTXiqqrY0nocdvkDmppaaqKw8QOG
QxQabad2TCIoUDfDuGphW32bgSDcG1Fmi3JOrycmBiBwgGk1LhqJuJOOa1yAA8426WbQVqSEMFzw
WTtE5hk9/vsuP46bKil3/eGnAvuFJakEzv9v5zRCKFbRAsrpboyNm25KVxA4xajppdT6iSM2YDwH
zybyVHLgYGgoS08BywO6Ro9iHjY0LR31nSEVNkuXvadCl9+akmERAWnJWpF8MaZhBQ8CXXm2ggtJ
PETCX7dVidAdwDFJjYWIyDKfUXWWFerSnraNKyXD088lkpQdYpmecBoVg2TwDBkwglcYLH1sPac8
8CEtRc7cHq92il+oqN/MhDOu/PkGiGIW9FyXH661KbptvnYENoBEgHKCBe9xDzEo3XldQjSxwTyX
QP3j5Z1ZewlOq1XcWiRxYlCo773+6xKJvCbU1kswa7Hc7QWvoNad57WYkWJmYbTu1Ml6nOA/B+YR
yqEt8bmREfR7wMUA5EAKpXTGlV0K5Apr7fRzdwlFi9THj2KQy5fvRZwLdmLXJG1+GWA+qWwDG0c/
L5rkJSQOGzeZSZMv/CwfIEB/f21D71IjLX+Beko9FZ3uh1zBq6ygrLKUPbd0UvvvOdPQ7MK3kJQo
uGWyaZl2RpK04/zxq1a3wrjMwVkKsLS0wF+SwLByXnpwlk7wHUHVXU4wZJzJKVt2Aq3eupCsyjX2
WeNF6a/jpy4fbuq7nsyv6zecF+wz8Hr73WIpsLMLL24mSGiiW6D/qtUF95hyOv/Po7EHTqKs2atF
6akUf1V535/mKwTvGf3nTvoqCyxfTtFB0lcC3j+/zHQ3WsoOih35g54vWGIluxS82fCIv0jIRWVe
Phjg0aHkN0zYmN00/xT6egzyu+aPNYuAj2hP7Fvc4e4gUwclkqJvOhcJY8ul21MzG8UHYjL+c3E7
dlP+L/E0AD487dY0BbA2gWQxw9f6F/tzwCqYNhyLTnnfiX2huwz28lXiWKM+9/ZklO4ZXVJ7PRan
z6m++DDudVPO9s3VS5G3uhiX3Z/5Q3Day2bzotJYH3HtozO6Vh2yCkgvc3qAq5/ek8XbDZBrdVlf
ylqmjFK3GcC9Iw2oEq3FTBULNyRIGxxgdr6ebCSFoWnsmE1Bqsy55ygt+ZhShMdgk9ew+IBFob+s
IOo5zoSLwBFHO7Mz/gJgemAhh2SeZlQX7w3LBbjao5Jr43bBlZz2wLAUS+tp+C5soAHdzDclaENY
xkFJC4LEIJNLhaugTGfJ6381+atznif+RDrm9PDsSe+ajCzvjHZ7smo4erxd54o6He+3lCPK8cT9
0G0YVaubsnGE7iFGI549wO+gsB7tQvY1+6DC5sICGedDVRGUafRJKQSnZuOs5xtOy0oaLuTMN3Ad
KCWlqniSuLp9n6nHM2eDN7TBjobKFyEABmix3bX1skm4sz2AeflvFxiD+e9F5ot1ex/D8jF6Sspm
TwLgavql01KjU2nHD6yAhVbW8iY2Z6jafYEMIsGjESC5Jtj8U1U0ZADu4zAx1nlf7nV3+u0WT4FR
UGv1F4gLhJmk7MxMEV0SXJYahZDaXlxAWi90YbVzvGqYTVuLZIFOLSCQj3xIwp7q+1tiSzYqpED6
M2x/Wltz/Gdld+8QUtAiWtjhlY1I7Vup/zxALbNBfbFFyWXQwooyPbfR4viS2XLda6NevVDeAU9J
vYzPLujTM/5lN1cIozZQUtQiG5LMCKqycWTJZwX5mn6Dlxg8llfqaepUvgCIefWXaGVeEd+T7AJS
6Xay4xKlVHet8p0sFPtqaNI4/zeqvowTFimtUnaTBbVxMQQMiS9yIFqkKiOCBJ/lz/hErzlL4n/R
WBpQjHTpC+bsjFVVZF0n3+mAdJ3NHozlmbumJQNSDD8e8NLBrZAZGp6LatgJfMhb7x1L/EVWswHD
nWbA+CBHeNeCBCqDcvKFCXI92AiXEOqCiDz9h1tE98XwBv1nGbGNFWJbewty7xIQkT4qzyB/iIs0
BnnYOus62R/nm5vJj2k4ZIQhHcE98/xU/Oz3pWcamMVPeIQYBe34bTZX+mih3gXr47ddkCDxggqr
tp4gwmlq9OT6MQJAlJClVMud2pI8mZOtTmYEkiRMlgmhtNLNCopRlx+XMOQPElFHNErRxf7MtDha
th6GGksUtQhCMaT9VBsna4Vtm+zWeMjqBukoLvVkn25LGG4dR2kiBgNi1gezzm46iaJbF4vqtU7P
3HdU+Z5Uk/Lqg6dL+3QQdnNestEj0GwVHR8QhoV9tnjC7O9qetllx8/OW8i2vjdDt75AYP/YeISK
OqF/ohWDHBsxuyQrHz/K8ic/dPe7TeNud+Fdk5Dj+jraXt7L8JbTvwNFHqpqrnCr2xkDQX5f/PFU
zbJCO9508lf+Mj+s3pBGbw72E9R7aIvKSFWswWT8BbUURQCrfGce22me2B1FeRyAN2GrqcDmZ5m4
d5fSprqdhxnpyR1MuuCsRVTLX8l60v63Y8+H/1yFM5b2YNsBP1JN3qz0ouMC/jtcuvVfjW2BC34U
6u4O7Ac3BWqvGT4f039Jc0lbuNAXBsViu9riyytLlce8X2MswUj5a6dTQr1gw4AFTjlk+mdgdnQF
h+DuMoUBJvQBaLzFzXBQwmNv4udKBVs2SV49sT09whNBfdO4a6sH3MuRWjcv/Kc+vNuDxoKK4Leb
BceEjUuTvNxpY2pnP/cObOxrrNMrz0q1/X7xOyuzysDxitnnwmUi36LjWPbAWdAe913K5QoRRbUN
aoyTG3OaloZkPhRnJ0QCBOUQE2s5eyfZeYEGcqF3Gqh6shBy31YFBw3P0i3i9XPfk7MUxXwxDUWP
xt+v+nqM9Gl3xTP4KoZ6h8ltUyocxTx2K41j8FHJhvMXZlEG6TWa4eW550CPBSFSo3sEuL2lPygu
6h8Z12lWhe1e0tr+tOgXXoBUiRaHZbNR0IHQ6fsQFVfC+VoIYjenzwrxXsGoRCTPZjswRERpfzd9
6rEzyTKdX7YixZTtjNEoijOZ3/lV0Hhoio4eV0kkd7uQ6dgkEZch2MGRPwUBdAYWWieXP6y/pnU4
Ec2+0ZC1LhF3jWYLLCvofDLXCFz8a07NpNXgHG+UQ/4ia/5l1HCcTh/WfpqMoCpETbN1cb2d5MEX
ODldXCeTzVnc5MUbLGQj9UMa4yw4hwgI9+kTRgjr8Mom1H8/jRHFh6I+cktoOtW2O6XgEbslOMfu
CNT2e67BFvrO/CTVdr2QjeCUZPJzwP7znHlsoZDLTlaFr04d0oEjsC2I4EflydH5oGG4b40liTVf
PV25liiBL7gZaqDbr8vgeY4ywpB/OS/2RK6QlpMOPxkeTxC9Oaf5cHtbUGoF9ySEQhUdenvYgnM7
pV4vdDDWjSoMgY84aToratCBJ2C8VBb6S8H8kmCPLH7+hk+nNg3B8HDzXhGkDNshoua8RS0IT2Lc
6tWnq4HdvMMwfXxCL1VIROoQcxh4PUp9/kTQnuf/ozIJFyCtso0TVENw6Yq3YHvUNssfpOA7DvTe
ZZbJ96TjWsvOxp50w+yBnA7BYPZsOnvFtosT22FOW7qoldtlKXO77LuGDJQBDSx0uuf1E9OFXNKB
dfEK+CkaMzwHoueunbKp/JYDTfpW59VSJ0CneLuqQoAp3wRlcIY1LHlFr2fvw8EcHnQhARIxCyED
EziT86CuScJbnNWn31aIulpk8X6OpDtSW0NEN2N7kwkytpIvC+v/LQqlnyHZki4dwICnhdP4deTE
26p18cujUmyPQN8BRSz2xKEsGvUwPr8q3NScfPWISOZnH017+gbqJKtXmxawn3FU/e9YidOp+qme
qh4Fssq5lB0krOS6JA1Q9pBllZYe2Oros31wQRJupJ9fS8cNMHPjrYB4GreIXYlzQ5qAnf6htG3/
9fmOGjcbejZE6Pq+Y4/mAFy++Rx4+bGnPq2ihTs5mL70Usth+pkreXn1viPllEyOK7NBn2gbJAaM
5nGjlzM+4GAzr/Jg3G5H6OcH24D2wavsLbZEHLeU5f+9K4mM0XylFn1eiWzVynYCVcJ4pTT8yN4y
pnJhhgyq6kWugDj98teTYO8mpHTUvSkWECM5pFt+INafBfv/QXV4u49Yr/1VfQt5ADIwzfI6FGF2
/OJXkBoug0WFC7Pk24yxn0mCEuH9lNc4OEsNXgexqrPPu3qEBRtbQ4K7B7Fkmw3DhjumoFqYz9eG
dvU1PFhjT59vUJ3VPDp87DXrUfkIZowlpoXAjrmvm7MXnTVT2mO+W8vzqEQG6FRU8OSmNl6V72Gy
aXlh3WNFu4feqQR4MCuU4Z8x8GuoPBs8x5ULb4nl4fnIszfTVVtM3oFH37s0U/UjNiwYEWzwZ/1l
vSlyQj9JTiyuwr38RDbZkIqcE/qtO2YHitZeFHF9WjrX/jjYFBf0gaVwy/JE1ziu91k7aiI2s/Re
GU1RKzMyC3e29CtOCbpBRNGLdFeSmmbqr4UQcVEziJEAP/KEEoGfM8wNr1i83b0ouftOwwrdDPH1
FxXfov+zyF/8ikOS+UcrgpLxwh3k1YbGPHHgnBDw8eM8nGm/S1e8zWKMgocyeZ84ohzR35wJbxqE
BtDKSjktkPHi9PaR83t9z/edUXzerdEQlAQ+iUu4Fu1bc7M1zX0pMXwF4z7uE6rUxqKn8LI9lsBK
sJ/18uApH55LBYMzgvs8RZwgZFr437KdjD9bsdH90RhHbbPMCbYExesSik0NbJ9O5jHT0RxCoISr
0+6p45YZP/QAHQsTnfLQGI6eb8gSUoa7+VZXyPK/T05fjJC3qdwRgG0P3AAVi+g5R3mtjFvmr1/h
iPUoHOgZMFAvGoXENuqM3ltRlLY8cGp5MXvSGeIGsoLTZicwTNoFSnrRIpByMY7ogHesFiQgq0fx
QTAKJegtg2jweENQWXhtgqYCeYApj2fKBH+YX6Wb3CQIP5bRjPDmVer27lw8KaYyGTiqy/ZO6yL7
BQRlwTKsB35OVykDw13xsBJ6QzXF6Bay5Py8RezEKDaUepq8oZRv3aHUymEigKBVD32/G4/NFKDm
uHv5WQNSxyhEeQ7CZ7Tj28JJpqG3uYdZnZFTRHRiE0Eam8Z/TDD5SuOVC+9zW9aBPaVi+q7xPwfa
2SQT1Ygqud9215ahwAnt8H7bq0wxfnt+bOcJj7bxESOJDhud8v9GElN+fmSnihwE1VyWW6DXQ6A3
D8kOW1gSsjhfsOt6gcP0EemLmXnxwIW5i+rDRZD52zKIzZPo9sVGSFV5hz+3WbdhnHX2kUlMTW+Q
N5cGS2el6eaE8jkUz1JGxHafI6LRnqIsSt0qfMmeh2wOHKpiYy28nI278a1FElIF8uBoXOjVEIyP
+JDn7v3M0iODugJQHo3f8Km421rjQ4Cm+l08qgtoRh33nldSOooa8cq08hPcrVZ84FQBoqE81ocq
xwvkRCyit1zshVwVT6NiVEjVGKkN58gf8UZrvTNL7CsQUs9kpk1qU3zMq3MXLwU66eZimW9kZ6Ro
H5TezIqjTsIGhlH+8hVGiZpwEyo89pleVe+9PhhdhEicghVbGOxZpPnBqTSTG2G+ZaJeXJ3OLaQA
lXXWgHmQaUB/ah2pK+EaVCmg5H9nuMxme0um8elIXLDItb0ESgKNxiaECKuAhB4zMLUIWjmWaPjD
b7FjBtK873EhRPPAus/WSFpeelzRybSBl9mhiBgn1RWYhQ/mG27Uft4LMKlQ6Tq9QL0lGZure2cN
7HCOq/TxcCDR2TwHHaprS9mSRhODFNs+naVKjnc7mFHAtlqEboD+GR4fNNQQXn5mYI29S+ChLP1S
W+14T/vNqfZvNdE0Q/JKFtMypYK4uLv51ZARqSve7pzYrOyw19FR031rZKIJltf91q0XTDT5VAjo
kGvswkOjTrVduqCs156MCiU9XNdyh1PFIlbzWU24deNq/cMfdixn0xdeiMrA1xc6U2jlcdZ6TVKl
iZhU3AFiw1oMg1tJ9RMKwQpawcmEAZ6IZWjI0aiCRtkYra1qUGzoJzIeXBdJ3ifq4jXJSSlQL/DT
eze0KSBH6q8Gw9YqLO0Ua/8LeESGf1+t6wzwU2JBlNpmJ4F7JMDsdzTWOC5bnkhA5/EmT5KK5XJx
3liBjj7W0M1n97EgDKav86lxRKDo+f7F5+d/N027LxFk8APBZT7crqlR46R/U3ztXWyGVuSKBuLT
PXleX4r6/p+8+1OXs7iEbQV02M7kgc68WqQaWYTgl+bkzRZn/wKA3Mmy3G+9DACxeX3oNQv4J8bK
1d7tVN7YXBh+I9S/4eFWINFFmJUDF9NPKCpTxdoB6uT7Lj24JvPWq4EbqmrhyONyB3LIMZquHTy3
k0sAOdI+3lTqQUmtUaeqkRYslLzYl3Fksa8/p5DNUWwOfIeVG308uRAt/bX3/TJmU0dBMh/piY3B
bwDTBMUg2IE4A35HUPsTNqVDoSQiKb73Ycb9+i3bWqG4DlGVFCa45XerTs40Od2lc+FK40AXRoDf
gbMxRiNC7QUsyxYaAqGw1JDyE/HmYDzSvf30cNE0dknvoW5Gs/hHK0a8FuXXkglMjwOXAO5uhQ5b
Rf3l99ExjDzZ7c4oMKzrd8zR7iLjti3mpX8RFDzj4Bt6qgQcH0dv93ldlQ6OUUGZw1aGEqj+TB1C
JfZ8NiWKZ1dJPKe6etqBrcF1gpr/y7gkIjzEsahWrQfKV5DlR2J9PQ9yOVobsOaXPRaRqBZQfGg7
QMxd8shS6124EesroPLNQbtTtZvWesDsUrhhGO7ftCcdW37M4hKT/TvvnQwCoxWHgrKWR0k3Vpnq
BIANrBheoOGoKQ3doKvmudzhinJcYORK+opHAztfN3Ap260id8IWdurFMTH1LhqJmPrYc/C6h7XT
aB+7BRIvqmShByhEbeVlyDD6YLmZjkfBQcWObslRCSC6cZDW3J+Y+XhF6XXKlM3J0GEK9DuIMAlt
wLDcCxBw/IcgHYNlKoQtyshcYu97FYomGxHM/fdsVy6F79FCbdC7LMoi2MBQ2y+0Efc+Iffl8DQX
RUwZ7PBhyUGMC3ZcNczvqJLK5lsgdxx/ylS8KD0Uk7boBSPLp4Iber2X92O2f7FQxUQt7X1ttqbk
tCBKJV73y3lF81GSJNT3tFFRihKhHzAPzlRwQXBF9S+Cv3F65QjU6sEN6nYQrkxicfc08KcJZfcz
cX6ljD06U76A76dYVkwPXBhvmYILxG40XdjsivajWFgGE3bu8KvV1ExuFMsxx/ojymPpNgqMmb5O
zEycoVkR/Js3RdzElDvwzG70FSlCRKKmskQA9duPxGcxk56w2UXDRRI8sjNKNT7skRlxjYoqDQke
vqDCuul46nCCDqpSclUy8wnNZzW3Dxf0bGfsdq6eB+n6t1c/IL5LHodENPbyj9f+lo0PvZrZ0pWS
IaL162zgpLWbKtbdsYEoASRHL1L3lbwLq/IeAFcBw5Dxb5gqAmluyFKTtJHqH1ECXoRiKJL71+Qt
/BSDgnmu0+rauq5TrSgOfCLDtyzXjBG5SxA2UdkUMj1BpWiqHG+VCsQtG99EjBsfGNHISMHVSxjq
GaY+ZoJXovmiL6q9LYR/YgGdTswhKJcrdT3XXVQUZAuKxJM3iIIt7JOoB2IBx+kF0Q4jw4vwqS13
YpFJAyQFOKJwmV0sD+ceomzslwbeSiz9fBJvdMJOQvE6D0m0gizNtKNTfHyK5kTLKOSShKx5QRDP
AlOZe4WHTiUEVIN2J+obPPXdU7x5tjd2YHA1d0tqU35HPe4xD/pmzlOBg9zG6WqzQZjxzWYcGakF
KBxEwg7JjikuBdFHAOOoNkTExokrzGbyE/jb1K84eeWkhpdNwSjh//aJucd0gSudUNiRxo/OnkWL
tK/vm9H1KJicEeeEW3lpipr1UuDsoqEZQI5mhONPahjuoMqli8DX8zKAud2/nGVtxI23II4nMw+A
fmr8Q5GTxQWYqnm7HdeZb0u2ZrxO+S1jYjtjmkkbUpqZrvgTIFjLeIS+vOdxo+nQbpraK3bAJHSA
m0Soh/uZpEBfc1AjpF3KdgrdsCLgjdA7LclkFhH9BR/OJc7cuYxO5dv3NMRaFQzy8TUO2OWPIneg
bqe/rCnkuKfA0PfyUwz7kvvxJeMvhvojPoxw8KOyFavSFnXSU33WwErRBH22fJOn+1Z4JdCxDeQY
L/YKlFOc+5zHW7oAIniroZBe5AfP/8vDUGH97bj6/0378vxYoQ8/oinXk1a1beNKa1bJNdzIymDx
K5mnpag8iCco1+HbwB+OMWyRraLklkIY4e83f4wBmcVsxVN2KZxHXKU2fPKABZk=
`protect end_protected
