��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl8��M@�"J��=�s�7���K�.&��G��]ʅGj�A��F=�E�bpU\-���JJm�6й�����R�g��n��%et��}#<*"cd.6��3�%��J6MX�7��&Ҵ��זT��_*�n�J~�(��Yͽ�^�<�]�n��hZ���W�ϵ��c�4��M}*�
b���E����pt�^Î�B}�+�����vU��ո�"�nos����q�B�82������lZWS��/�������o+�
w�@��T�f*��fԖR)������>�����ڻy�'���̨�VA���2�Q��;홙���}���� �ƹ������8X�N#D�FM�X�닌��;���Z3�V�Lw���vք(6=���|�]�A#�����tqd�
a�0���q�%�����U��rLט��p�G=��g�$�B�l��%Ka�0��N�n���ӱ��ͯ^ڙ��d*�t�vnS����_��U�;.*�L6t\��M�s8��}�Z�Z�wƫ��$�ď����)�2�y<��e7\;r��n=�K���a��]�$.ϙ�r��M�M��
֧�Tp�L�b)�5���2/�.����ƍC���"��_�<2�:N2Oi�_��+�io챩L����2:��wCtM���Z換�M���Ҁ%��"h_��ͧ��@=�������6��3�S=Uk�4� �S�!�ż����ak��Rf�dP$i��Rgmx3�IcY�hG�p�����ij���s`��z4��3n�]s7[���5p�;(:�v�>�nu�����n��36?>mD��R����*5�hݨcl3���h��)���|LVW���I�UVw
-�u_���`v�rcG���P���@�_ih�i$�F�~�2�3�KC�|���S��{-#���z!Z�#��nE���Y`i�����usQ�fM���W�ⵟ�*�֤����)v�R`EK'�`�E������O�Z)���'��m/Lj{�e1g8��y�H��"�[�vP���u��1�����!�JD*����mt�,�--�����Cj���Ǉ��Acn���qf�źkQ�XN�J�úCof�fc����z&�Z���k��J~�'��¦o�/����nZ��u�IP�gY��aؒ�V�=X�p�j�p��!����%[�,���oq�$�l�hQe�a��f������DL���L�V�7L߳��0��#��e*N;>�/��q��ձ���/�`�g2�*J+�2j��I�HIo��EBsv#w�Xf�{��UJh�-�u=�߿���^Ft���/��GW��^�N?v�X��v���n�22�_��У�5���Ϣ��K����X��q�^�F�ir��@��ytm���~��p=�����Gi������e8,$��@Ѭs�}��r�\d�Q���4�`�1L1�{{v�H7�73Al���n싫�/:�#D~>r5k%���-���ju&�+.��qK�����x�h�]04u9|��ZLS�K.U @���srȘ�R�Bo�3��W�`V���,���|W����C���jRW;e$ꂘ[E��{:��M�l��t�vn�Hv����?�7k@��R�#�����U��$P�&���iN���+P@a�ņ:�rʪ�}7�|���3��i�U���1mC_���4��3���E��U��d���V_w�������@:�����NL�+Y=�wt�#��j�\���R�e�Zj���v��/�F�|#���%�@�Θ.Z2�V�	���X9�_�p#���B�Ԏ�4�M���;����	����â|���s�q�dq�>��d�?g�7���b_�ݤ[�a�>�P�v�Lo��\P���^o(	�����\���������g�(�
��n�H�c�<��tc�#p�TJgp$ʒ��Y6o�Mk���Xi�AX��Y�!Z���T�G�Fn���s���ͳFt���֚lpa'՚�l��QNt���Ƽ�5
��Ʀ����&�l_`� a��t�n>�/�j'1���c�-.�X G���~��d�4E��e�"�2QS���"��}m�1#S��#d*����f�`h:�X�"x�Hw��{k�X�ٌ��	��_�n�B]}�!���#ƍ��N٦��&�O��+�~��a��w*��4?�z�A9���<uE6�C�orS��7(]�?�o([�Y{�So��m�[\�$x�s�K���)�g��C��@ua��zX������ ���/Ae���]�cΗW\����L[�uj�Fp4�s��rJ���w���_��ڊ�5�D�ߦOB�*��v�3��4S�i���㖕�� �+��Xr�i����Xn���,�{��aw��"�v��:���|��M`��ŸM�NL� )�θ"��g���Th���fƭ��5B�mr�]Ɨ?�k8��c>���jWyI8��j�Q�!�vOv�؝���aF��nr�����Q�E9�P�2}��2-�6�;&S���Z/Ք)үl�OK��f��2��u�<f��׆��֋�o3�H-�9&�����`F��E���$��G�.��^e��#�'1(`�)�	��T�.�$I5� ���i<Թ��C�F�|�.doR���ص���n��i���*U�Z:1�,f0�5.��<�3�$
�"}��w`�ȩ,�e�c�/Q8�.�:g��r��w�eQ�)�J)���y��J�Ա����R�/GA-$�������j�F���;
�4߭�\�ͽ�~UM����:i�Vs$�Q4��SD�狮�p�fv�:釐��#��0fK͙%�ȃ�<�\��S���?�2B�]�'ۯ��wa�H�0��<����D+�I�MݦG>X~=��ݬp?(6���h��X�/_"t͗5��ӻŀ�5��R>�dU��}cn��� �N8-�w���v�&|x��29>�VFvC #h9��Q���#[�x������N�U��t7k�����1ZW+7�X[qOV��Ñ�9JQ_+�|�	A2eJ��>q%C �2�C��������,\�=c{�c�`�&��x��+38����K����6�K�o��m�2�T��n|��D x�{�A"�
3���@�pػ&^	:�K��B���nr!��ߕwc�gT�A�?�l)��5.��A!�����m��9I�0{��=������b5��'،�����p�i-�bA��D�堗��Vֈ��}�t��פ�XG�IѦ���7����E�<���	�.�����E�@��)3{���1� Ķ%�Q�ۉ�E�U��\c��VU���2J���3��x�ֈ�\��m��kT�A��ê�۟I��q�O�lND�S+s�'AN�a7/�S˚w�%��!ܤB�����,V��LU���0j_Y3�Ѯ^�z^�'�T�gp�?jh��`8M�~淘��+����#Ȩ�x�vz7�%~B�F�N��Q�t����c��}<5�=�(G{��D�85˄��ϒ6՛:��$b�.*�M��`��
D����L��3�c�җ	S�])�m��w�+D%�d�c.�ˍk�]Mۀ Q���cg��4�Ҹdj��☄:R�4��{o2J.�ɗ�%����X(����#�����Z=.d�p>�ƀ0���+�|c�찫����(`ڍ�M�s.Og����"3nK����.���9F�Y h������g�yD���
f	�b��V���y��������"����/�����mxD$�nP���ތ�}9-�����bY���B�,RlQsk��_�`�Z�vGKJ��>k��5�D	���6�&F@���o���`o�����G`K�#�g[!оT�e����H��[Vb鍟����{�ю���P��.]>�,_\�L�n�[؜k�'��_�0ݩ1�D���-���F���!t�3h�u��Bo5�%1@2"`�͢F�_^�W�O��V�	�	 *��%��6�5C�h������@�y�z �˙�[�'�D
�>S���z��s�83E_B����u񸤣��q(]�s���fm�ǓP�57�I�̞��f��
u��������JaQl6TiG�M��cs-cQ�y���'S:r=B�XV��|�D� �r�`��6�a�1ۘ�i,��2����� ?��R��M�����+�z���No��@��ƴ�$e�DPuü��:J�׿�:�������YF��Ō�K�rm˚ީ�{����JuB��G��l�儜�K�3^ª8��{��m�Ou��� ������	(��/�DT�}�	y!�8�9U�S�gv-���M��E�~
���Ȭ��]�x�>���q����*ƪ�HX�MmI#�;�c�����ġn�h.�8��-;�Ò��@�ò	�E���4~Z�$���qc|�ܜ�4؅Io@cX�����	[��xš8��Q���u�Q��h,Ov��TK�L��/1@ �� a=�W@S7��:^({�P�<͞OT��e����vlA0�ŭg��L$_�]@���v�_/x�2��]м3��Nn�*��)������3�ŗ.�.շE菈}U�˱����������'Q��+=�&K+���~��c���V���^���ˋ�64J�n���V��{�k�rq��P�Q��jZӑ�v\CwM(�+���[-�j:��x�0��j5Y�����{�㮥���r�h�C����uL:�Mz�R'ȍZ��pt
慇n]
h��n���2
���d�ع���  �F2Z�w��A�R�_*nT�����Ѝ������r#��R�~�������쁲9�����g�9f��W�,�.3�sj_� ���]����.��Fc�Y�5���m!4a��n`��u}48���9�zͭ	��c�:��Y����w*�KⒸ�oۓ�RK�߱Sl�I;IAxKI^��U��%�ص�����6�<p��q�X�R~dӐ�l.�;�C�0Q��Z���b��V�>�No�TT3�(��@��[�$6�X$Z��j��J�'F����u�S�aϏ6f��m"�*��׵�V��GXi�m	���9��C��-��N��_�"��a��g8��7�����zѹ���K7kc����[����]7P/���6e�W�F�$l_�d��()ƥ�@b	e����iҰ0���ܻ��~�R�c���ū��CEi��I�s6,���ZR�l��4��Z�N���r���|�S4-��eM-��Hg��ځ�׆�!iz9�'�)����p��d�~B����~M� =7��ڜ�PY6�f��[�l�*H��BJP˼'�_��lǠ�:�`P��O�7���fo�[A�l�L���\ۭ��d\)�M�z�pJˉ�
�8*�C;�v�e{���瑷�P�X��ÆS{��T/��6�C������	ٯ�PVq�4�.�S�6E&J�.i�㡄�3��yk�F˻ٞz�)��#t����O�h<�p�<L`���4�o�KF��7.׫��*�M8�}���x�O�]RV,\���{�l?z9��\�����#qMb��T"B`�fW�����ʰ�.���g��M�6��e��C�j����p�k�vq)��q�\o�!p�|�BRstY��&P�`�*��7�m\�����
h��n�!�}�G ��I�s:`7u4^iޮ$t<�p��@p<�e���;d��{���U.����;!��k��>��5q��\��<�<h7�;�E/�
���ܞ�G�2L�}'H��D"���Xo�`��E�r�3QX�.9�����oh�3�z��u�hEn���su�w0 d��V�x	�����_�P��5RAKA-��F���g���MiB�� +Ѯd��]w�|���M����ل�U������}Ӂj�W1���gT�����&�W�ox�¼(�^zB\�����˟�ő/:��=�=��f��|�R�%�KY�⪓˯Q�n��j�K�|nX,���gFz�}_z�d,�oG��4o�6����{����V5��^3.jX�i%z��~�xL{D�	���H�[ݚ��o��=.�ˏ�ll���uܞبO���ِ��=��	�����5_��U\�9"r$�9?�5�����i~c5@i�����$�O�+��SPv��0��R%sz_oPH�FR���`��L�H+�iY�"4�2e�ٛ�c�(bt���Ԯ�t;`R�mü_�K
�IM .ټ�`��2��e��Ju!M���D�l�����/�U��o� b�?��`��}�YJJ2ý����?n�ۡ�(�1Z���f_����	�����U�ó����'�V��^�mx�m�5�k��l�mt,���N}1�`z��K�l��2��s�L��i	������ws�{ �i^L�i��S�ף	b��E��d��Q���9'K�-�[~z��;��0 
Q��ǿ'C�v��ȣ��Q����e�[�!�'��t�(O�V�j�}�iR�����ksd4��y�{z�*��J޹�H�"����ύ��(U)|>(���#m�2z����=�w�(�����%���J��r�9'N����U��k{oA�KY�A����\�����0��n~�7x�E���(�5_���CP�oMPG��uοC?�aR�ĝB(�5-���v$��}+7�1D���RPRv���;���r)��y���X��k �|D�)&
<�iT��R��Ɏ��%� �Uok�y�Ewu�8��PHW&-Z�~��� N�-ȇ�K���ӝ�`K�I{>`�P@�57d^앐S]�b� �U�%}��v�k���?Îehn�ؚ��`({OI"]cjR�e
\d��-ڞXx��u<?�Ś��q���m�;��s�R$�w���ݶ­�IQ�N?5��2�Eh鹝{���3s��JX��C�A/H>u�N����8�����L'���j'�GW�כ	O?G*���g�4M�G��Yr�]�c��!��H�lÔ���� 5�/C%�e��!�퀨���F���&�HF��rq<�gǓ�G�A�K!��s28�7h���I����hY�+X�(�t�8)�9��>�����p_&���Ȥٶ��O���(=�X{�3�s
k�#=�d��^�=�rj�4\/��y3zKL^&m=�܋H�Nq������3F��e��֙%0�I� �4<T�����J���ND4In&�wT�Ğy8F�/��z�'#�k6֦����d3�2�푅�?ۄ��Dmf�F�辡�{W���I=����	Թ=8N���L��]���o��[.��*��5�9X��B��O��";5h�a�׾ʄ��y�>��.��oT��  ���h�$J��&<%�}�ѝ�촖���01jST�� �&���D���2۾��PP6�s�waW�RTO��+jJ�����nTd���P�0�Jf��5��_�nL����@eu�oL�]�5�$)�g�'~���o��B�qenx��?5���^l���b}�^Gh�M������k��<ݡG�&s0I�)�O�	�tⵞF�j��ӌ-�^qu��j�g�̈́8��)�`���]Շڲ}vj��n4SA���A��e�P��׈�s)���1�Y��S_k�'Ol�=o�X*|u���34gf�3}���v����m�	y���T?R�Z��X��eS��~B�N����RC�r���޵�f���ޝ�*�����l���p�_H�Ń	T*W�ŧ/��Ko�3͝eX��"*��J��V��Κ�H�?@^�r��lNgw��; YDM�����(T#�8GR��ã(&����eT@����b���G�Ӄd��i�f �M�'j�h�O�x-U����RJ�o���ӈ���֕'��� ��,����0,Z�� ԣP���(;c�����y�O�jX�@#s���Z��х��T)�a��*=�K�y�mqZYkS;(�xNLǘꇨ�K�s��yҍ�Zٸ��W���#��ڈ��9�S�p�3��x��1��-ۨ��Z��),*�B�Cb��L�/���b�+y�g38=#J[x�����DtK�4��X�m��`Z���U`�,Y_�[]��$�,�&����+�a��V1��濵W^ �%�|�W[�8?��qs�S�5�oUXc gʢ<4�Z�����Pc���5\s�]�����6�|�d�+�t5}�4k :�y������g�ofW����g��R�L[10N�x�|jz���	"��P���@�G�����y����ݵ��UT��rϩ1�w��{PO�|~43�$9f- �Ҥ0p%��qiu�)��<���Ѝ�A;#���YM7����2mh�rk�n�y}����K+L2H��{@Ü���؟���|�Q����RzM��$���s��;�r5�L�2��3�Թs�x��i
 ��)AM�򂻃y�ʝ%��!����^g/[����#�gKH��{OJ�Bv�0T&!dB�o6Jq14��M���$�䲾�ù��W�����.���:@�M꼔��W�r4S<PAWe�B�.��p}��n*��LaIe|�\�^���m�O����m��9���}