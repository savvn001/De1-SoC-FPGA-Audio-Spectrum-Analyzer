-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SioPacdWjfV+yqnDzZgEpuMSLKXMmRPw3fKgwNzXHYzTwB9YEy2PF4j6zRsBFikjdPM4H9/hVuPf
mcrd9isWggqegDbLdz3B7ISrw6mYTph+FTgoN0I+mbDspdEfcBBreR+CVq05wPWpckMqDP1tgpDT
K8b4HEeYACq2sp5PDvyKu3wt9qiHeF/cHFHwbe0RHOnTHlCGbrMulwo4xD/YTYGUJVR0Id0/Ve0+
YDy/46H2Pj8HqZszQK0G9EDN3BQQtJ7zAKw2V7cuzVGYWxv1crT08hfQnOKKoZOXm+/rYaH/R7ia
4DxrogvFZAgr4x17PfQvi956M6jual3M75AZiw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
U0D+52H+NfO1WTDNLM7JIlRhAVKMCE31IFUswyqJnVkdm1DoHOsc9QfQ3BTX/3deoXPNVJl+kCfd
arFqLALed+uhlOhQTb6KLO72eqrJKxNxSzuvDi4aovNZyfS997Ru8oSfHLTaGy1DA8g2j9/0RFi6
2XnbpgztRoM/4Ghdcyd7IBGr++wyHqfM1D98A5NXs0YRsDN13pHKZfhFxBLIjBxtHgpf1KHaVd/M
MQ0+mkWzqhyJdrdYbmwYiiWo+KUMYF/34CJ0D8qjyKB5126GF+LZbbz5KuzkEMIkt71JA9EBAqze
PmqcL/z5JFRlO3zEX+lLpaLkuNzQzqVNjzrYkBiwDsHyQeV+X51XFr9Dm8jgRxQHa1gVJ2iDneW3
3k0pNAQ6Xb6W9TLMB3MzR8WuN1WW8uPeFp7Jk0gNmAv6PwY1HVOb6aF6d25Aqe4XJ6JYLSoRABJg
BRgSlEm/j7ZsWLdWgdh9oO9kcHB+cF9Hai7yz4QfVxH5PAMkllalXR1orlZdc/CJUEYDRq5grSoq
VaiLU+lqx7aCeKfSYjuPozkzc5/qpiKrtw+FYwLF6lEZSaiWgj933+85mmFZ14NFR8y3slBl1jwk
UEPkCRVV0ivtG5OL5iNwJP2D4H2/GeFcS9OwBjsm7XIvIU9IPoWCrlmPYwedCaSUQIY4P74Z367B
iCmhDM8PjO6CqN1CJ8MGWAllyo+2/2nXCBFcYLpBHly1lSwaz1J00x0LZhOIhrAEyMQnMYcrcFYx
hLmJsn7AWk7mZl96chV5h3AgMXigXwXTlqPADno2zFLKIBYDNt/0BNxqq2M1V2GOwWqC0A0Cx21v
PNdC6A6it3OyS0sh+4F6MO6E1D0ZPUwD2SpgmmTHPsdZzeLFez6MCmyl6RS7QT7vCLzZJ8Fff1Eb
mecYSw7iQmEwimADWwx/f4X1LKnTeBQedvGeqWwUXm2WI+xq15uIe9wMOXKwVn6sxt+bLzBrms7q
jDtqUoRaLHdBgVGokQLqWAND7gKXAqNqZbwByGlvyR+4K0N0yBbh+rw/HQA0huCALm355eJn88A8
d7zohEjiYTob9D/M0ngC/Lc25XwC4pUKfO8DmAkCfJUv89AFyGYkEnUw+FeRd8bUfZ4MP8C4SC7c
TMzyFslX6zgCIzou97uUPxXzwVV+g3MV+uGKc4GQpsCXlATsh7uKYuNlf11psfYmsXBUoim369MR
ujh3qJWiBsy+HGKiIJJjH9Q4lMX9psrFW1O7tFMgtbpJo2BAy3JtHuh41GwS/o0Seu6ATk/Rh8rW
AhblAwGM3wS1SxnHZEO6YQTzBsPFWmVLv4B4YRYGfv04kFRAJhC2B6Bukf2ytRytY/VoYfzmB1aw
H+pSFO51si2ohX1ZAQBJUKtzGomcz7FVM1ZeWkuungKmSKASEiu1svzopjxjZZSlQ16XCEyLpt2o
Pik9YUYgRyyOM/nXr9axukqAt6SF5er/4yAXaJ58G8Wxp9k2FBEhEP3iawhaypKf5lPhYdma1PZ2
liql0ixhZwqfqLTsUxikdxSeK29DDT7qw++SMoaVz1ckHb4g59SHosTy99gOxbrTc+9DOcRIDgSK
mFST5j6ioBsUcyZkxwaBmeJ+DIRKCsZHwKwA8vLCqZjokIX/2CFvpTfqTHqvaGrcNfA3si2mQHyT
xNMfzGJ2fS2DNJcvW97beFGsmMVnav9MY0ZTp0ZBn3EshOnUHRxzfXb9GtWH0fFX3AcLoUOsK78c
URPL98E8IeABd2n38L4WQ3ROlvi6H0a6GzK7kaNF23++fP8nio+uspVPLMYh9X1Gm6eMWn5g0R9F
V/LyLGynPL5ryygrWyqzz7px8A0CPx3sxd0n0M8rlg7UTbBmEG+iNvAqe6VOxfdCFDYbgQiOlsgM
DThhl5o50N+Ohe4Juyswg8tcUpUXv8mmxWx0kdOOxwbpQae8totukMsbbCCPvGWLpvqg0ovLkY5w
5aTCLOCJOVHXAsdmucbO7B6up9qcDk0hvQGavjoZfsycu6ewKqYBTQX0EDFe1orou20UhLgTjX/d
ma8BDBAa6XKe31s44rZZUPdbR+08sL6I0ttOUIRxPCS4vsx0B56fCAL8tbmaYp28ap3lYKCv3Cof
vG6E5kO1euSLMVWvMuAFNRcjn+PNnsAp4iBSU4l8pqUzy+Rn+2TzHehAeBiSf3TThTN2fpiwJ1W0
7o0biMZq9mPbRSn/edfa53oVIfJA+vzaQF6eYk4zdiv4MwsIQf1MEdV3IP8h2iaNAaB5hJFVEKLk
uQgyahF1xCfRZROXigKbCw86/LK1SfbBMoQlXGdC76Fo2ThV8g3cl9HT6sRjDRcOP+OiRf0OJu+B
wpvnMHqOi7HNIfYiMu4b3HHNCnIGHHUVn1MuqJejsIJRuAhwqZOsAwGoJ74rnhWVao10Xj45L95r
+s+hK7eN5fR7q1NuIvj6AO+5tF8T14Kpit0gA4zQzDuksAJ1uBfDgc4MSWZeb7mf4MRyrvmIv044
OaLtkCPjUhUONusEg4TDJwNeTf1C7YYvwNwIk38ckihTupGBD9CCjC1D8TzkwvZZ+G4F5nxvaK1/
+5ew9aWbRCk0JjQySH4zv4vvJ4Ey+KfZ8/wPZVwZOFAaSEdMJLPNZBaNjvoaSq+NZMOMT5oV8xz7
TYhfAAUJpY8u5WzfAIgYN6/vBWo0pd6kN9x7xNteruhIhUbzUWK6xfLK+v0AG3Hj4H2wrQToRVhF
G1P+/c4hz3H0DDdt7aTjqfy1oOgwNfgH/esVh0f8z0NcNaM6/mEItyoG0djeAc4JUvjXsci3fAMm
V4G7G0XDSDXfUSoiZeUnDCYIlxQL0PVWDTwztoXfBu4QEKdOJUGAY0qqNL2EpAt71omhxsKZwVYw
W/JMSZEPjXqZGHYYiBtsGCtO+qXBsWcziy1NQBp7yfXmxHG2NYqfLFpi9GZp124Mg2isVrCseDpX
D9Zcrbz0GOJcQI5JuwPxkmoCve7LPtzAfgJ0k3Bruuf7LDvUaKzxTSerR45ycOsxsTcDokeMa4lM
c+1iZsLCQodZPpRQoiDWtS7TxrOc5eVMRHhLRNU0QeggoGL/lXaeRueMW+TnR7IFKwOK4F2rJ0gO
8P3J6UjeiRaSUCqa4OPgmwzGM6v7lMkwnbpOhKmq5sQRaBZi4e20xKe8stSG+yqOFa5Cfm1WcL8z
ELKZbYzk/MqufrxjFGUJj6F2ojN0nJmbRLBCTHPwwYnbSygL5hdmLzouQ2X3sEgi0LfV9AtcxlWM
N9usOokDc/oZpjcfv6x9sNGxuKN5LxyATpBE3mhx3/4d+EKdhQwp9DYwHNb7O0f6aVDDSImrK41I
moj+EaU7oIpbwpRxcuHg0hSlmDQqV9ftmLWO11CKsxxllTYPDqMVf2Vahoy8vKolzVq1ddWfq++0
YDfuqW2yZl4UYfISFVO1MtwxWQeBTAWPx27tWnxlZGFdh+PbDxdH6QeiiP6npOuISNxVGCGFDV8t
CcKy0Puo5Z2GDzvOcSjQ50Asch4kyilldyUTpst1Briwt51kXUzqLfNwfHNYM3HAs3BJKR+HGBXU
jakoANAnl3nuyxfiRqCyatN0cnat3GcH5B9RzBdIbo4KnUOsxZPNJhFAVg/Wd1wDHJSfTjL69aW1
n/MhfhZAM7LIoqWXD8RBE3tATbVMISc5xbY5KV6nb8eNNsLJRH1M9/0kHDUo394rgqNaN/J9dLXi
IjmocKGcgAd0jE8Pv+jT4ZLsEaHggsa9fI5qSw3QKjmWxIgR/2CSdDmgtd9dgYp1Wo0hwg7YEIYa
d3PO7/mmxaAhi4WBCBaD8EO7/Ke9agVKUpj/EsI9Ao1mB2eaTK/YMJOfUt8q0L4Uvzo+TtSbiV/l
HUIkZGOM531CIrZ5Rx8QmeiXOGLX/Gs8mKz6Gkri6T3LKE7W2hOK4zke2sN/pRUBsAnq8TCRRuAv
URW3qCX/76jQIfHerdfCX6mjvkL4nkMwIleCs3FhaUMOfbFemQMHtYzgZBopU0X4yNn027FseTdC
RCR3dLD79I8jeXgsJD6Z5V2SuvH7l94W2vkmotb1yB1lJrH6lRYA0uOwhBOP29jS5+aetbkPbivv
niKbAfh1Uzgf9FGtTFpgFlvObp7rQxzGHwrEa41dnHqQwV3rFj+aEUkOLd6DYwEadejD9WNRVbOt
fF3qeMQ6ocpQqNa0k0zXvqZTjZtoyEQQBFvzMB8r7hOp1730bVCzRgeagxlgcPVdkUde+OtqUCk4
cPKGk/y3l3lZzDn73fPCcnR3ImYAzcqB3KfkHq9L9VtVHMOhP/JVfjTb4UrOWE0bqpbG0icPTsI2
SP3Z2SRtz2T6QNMYhwt/hP6hPQ/HPUFDiIlHZBn8oDxX2h1Yj5q1cm99B5UPsncw+XbACQM62Stf
FayEkQSWrtWX9760zbRHJF8TKmWBqUbYwzoYbCauryp1ATrnreCzISyDrlcnia/74XF+u+vDrmN+
2+/I2/iEubprtqEE5m9M/3vFa3b8EgYdptm0533WNdqSitIcLNqjokmTl6A594QqiaHWhevjRVgN
bPE2oxI2kRVMq+wnklPtj5N9MI6But4FgBHP0HC4r5M7DDCMNwxR324EUrSeHtTnIHo+9EEQWzq7
IyvYKkmH2DVDmFkJwTvGWiKI1WQIrXGTKW5UK8c3X2nJZlYT/EoXjle0q5QuclJkAUz3/DIesskW
FZhP9YvV5lolC7g/hhvnxqDadFGDe4DEgFtMkzgxUCPUp+IU/n0qZHf4LrhLsweNR40Ry4jwZ4TR
o864oWpZ9hxLRc2CJ8rOAjVdi87vdxZ2otp+vKCFIWVRbjAyIuHdMXMTpFI1sZRSRLbEQGi82i5E
X78apOzJn30ex0Yu1ObDWWDfguahFq+HOPhyFssMi6o0bzBw4PNzJu7dEOfzZ7eH0kH5SG5hfgIc
X42esC/t79PfsM80AjXvlfPdon3VGyUkI+yJx4ucTcY5H98pzdCDmzn+p5mKztjwKhnINaGJZ+5W
iRrhXVfnN9GSmIDrbaYkwpJqgu0VLtRDn2q9tVmGVaZi5H1LHXHppIWLTMenYzWCWzV0ElNUpjnn
5e5AjOUw87fugB1UjEh4scxRF7JJZUdiwcVCcnDqfuZEjDtwqiRV+niMrSvJ01LZmwgWmT/D0q3e
VhKuzZU0Yw46QMtbp0owxBakgqOVmoEnIiqsZGsB5kc8GVtyoXV2miaeSg89Reg8QVxoekf4XPBB
ScAaXSo9PQjstgnCqFu+xSzWFyRaf7HGw1r7+Wo+jWKttD6Z9E4cTuvULQ0QdqSrjWh8tIv5goT2
gm7fxoyqEMH3TSLu3zPilexwmsQ4kEoP08C4MfEXu7h/UhqmO9zlzpQOB5HUdcl/4/o33d61j3c1
I6HKQ+GorloO3U7Ki+xpktbt71lqXxHMsHayUU3NGmUEuuWJXyy94gt4OVgP1XWqGYksGFRHt5JM
ojrgHscxs5jlMMLnWYois3J7zqlL3VNohWP6R2Dhx0M9OKTFeLMieGmyAO6twZRbPojKEYheNeKh
dpQUbmSPDxq77nQSSkZU3UQtruJdkKf3k4LHjaycmwzotyVuB3dZ8RlbqEWdve4uTXIEGfpvQA8s
GfJfAreJCGyxxdm0K+5YTtMe4aDM+t1KuJIXq1Jq3PN7Yt8LjXC/wDLdOelsJWVq/I7112AZICDb
HJPJYwqs96BN+mu8jOUwC0HuF1YVw+L9hHhY99iX/EaKuSeJ0Z3w4sea3Ya5kerJ6VqAyShQG7ue
JeaUJLCIHvZLIRpyeWPWJFTM/ipA3H4fRBAun8VXwMuf7tdddx0oZ+2GMinBIgJMV7GpLlUeXg3v
CrTKeovUQnq500H/Kp7P7ElrTYOC5ZlSm81gRCS9kImjMIF13hrhnKMGfi0Q2h4RrKeBv/AWYtou
esNNumAcRL7/th855TpIBWMou9rbnooJJNBg8lM17e4ZiLkCS1vhUg+TTJK2xCD5ujVu0byAyK6J
HcySHI0vEf598un1X75JWS/NDDhID0pNSUZ1rzrbY/eyX9/C6UfHdkw0Y8P0FnGcbVDuaV1KFTfq
CARhhVgkHNDR332GCtDDWaxqUwD5lO9sVSnJo8BQeebs1w+67TFjeNZvorVP2C/lhnHskWuMeObc
KuLWklg/vq369OJq0An2i3UJMNOPpfa4Yvk/9pgsOmz5jaWe0OML5noCbCn7FdVWOTcQMJQtz/zd
EK/KjHe/SWggEXS9JryyrQCJf5j0jYwN5kogMev0rYwsWjgPUN8OLJuEalgsYnTRIPJfgw459Bhw
mPrRkH+ImbIbMbfsEnUc9wV+ZD5gDcvqf8i8jI8fn3CZLTmjAOypLSeTOD6+bkrRej81lzXsghP3
fqQ4kAYkiQkRUbRNIflsirB1rCsI0V7T4G9kHEwzQeqY6pFEMXP1uPtQlGiMqCQjiM+szsdlnxsu
qtSTC3ID2/h/IOxFDnEv7P0i0pVW7pCqNwtiESQkwOKY7SYrwB91scMObAjY+wNZPu7PTk1i71cD
qyTaFk8uaADGTKVAsEg2RTUb91rZKdB6wl5QN6Gb6DB4CZRYTXeL/tOrnDEXbf2CCKZRQzU9AATC
hLzoNOprmM3O9cG9Eu6DtKQimtL3xOP3SOTS7TEW0H9fhcX0MvhCZP1SUcqXehlgqolce1untfoe
TTRB87GTU4VKfG9mlMnlu85JZfxudMgbKOJB7UgpE9rMVh4Y8YktgcAVCIBbGcBe0K5RAvtdVjPT
L19ye+tta2xQki6PhTlM0yFsRfrDkEfbe0wsgMWlseCzfF16scSFW6VN+/prVLo+5i/roqy7hA4t
Wh9ktkGdZDgkLiJIL+nVJ24Jg6kFLGcVhIbZc4wY0pfyNaiJvS4M1o5KCk+YQr3gTTUCfsaL81Cn
6VgQn0+wWnouZQwLta0N80mPrkBsUpObX6PBcelmxblH86T++ULh/KCxDq3H1iJXqtZ2ab7S0GOw
MblUWWhkUun+8D1TyMIISYfZE+3tkwtjOymHlPul9zmC7muQDVATO5/4aEUfPKgjEeH4cgAKIej1
o7Mmv27UTDDvy5X6rwAv0pd2GXOpUif8HH7Fk01Ds2bCdMYT1fkYZgRaE3us0Ca6j/IZJjWyk7Xp
lXz/fqppkXJSwPgTnEkmCbMhL7NWfyYzz0VZrkhtk6jaM6iZwz+zWfNnWP0zZkmlbxI11dsGkYO9
bcBr23NF72Z1rCXPFYqcagYoLpjhM5gcQCoyvU1nZXdWBC05KV5uylSmxpyJxdA9x9ebAUPKkCWM
+mXdbB2Kd9RRRvEPbiqsXRjQhBqUYRJpRQAp5CA6leY63KiZ29mRsqkeA/JbcSL2GRl3MiLyhR99
db5aoN0b7ieAQXiDearuITxHtVFJD3+cK44htmULt2mkANewjIk1UIoJK45eDfgDBbES5F82Efpb
LxP/yIPpEOldG/W1tzOP3t98HisEAzSWEaPNWtdtD5Pn2mU6gVrK8AWXG+sm3/H8/rcLsyw2Z6n/
qKjKeaJ5q0imHsLuEvv94ZqvyWn9JdPkgTey/yUAFJVegpT10ZtEMPUK+xGnxrWQIURv9sve3ZVf
iKSRfocyL2TCe8VVIB0HmExN/4XqHxYGDsj0SE8ayKUdN29tk/2TpcoQ9/Ff+qI8QImp3Tfc0PWZ
mUKW3a1I4+zR5bMIM1H4KusYjMWp1/wwV0B5KGishua+csR7U5uj5j+miy6jt0+p0JnfZcvreTtW
LFXFYrKJYUp0YRQwj5iqWhSQFn7r0dFp7pEb+yeUqcUixTjf2/NpUx88DN2H5Ol3d8u5CIaRWdxv
YAgvWno66lT9MSL/eS5wcGFMunQHDUbN19N2SMNaZSjDPtzDGcgXw4K/s7w6jox1/Z78qeaF4g5z
jwxDBH9avLbbgxxvqc4qCBB0qDENs+OsSqA0TiI0KYi+I9osK4hjxla5F0Le9LoTg3aZQWIBZX0S
x7IT3+USO5pHmV+VpJJQAugFqPsTbynDrTDl840JwrPH6BAqHaUjcYaVgxvP6j/Zy2dFHIiIsXWR
YcWg0Q630uhmoAxC5PXvi/hM3nFLbpegdOV1BbZHe0L5EUqQQinL2X0aqEbk8UYXHsnV+U9XI0zI
JSCdP5qPileJwgCnwC5YvYev0We49yFcmnjx/LgrNcZ/QuP6I/uQ+NpN7naGpli6y3zV5fImm7ag
W+jKLXdO3cEXYaI+BzxB2sliR0WQ/bC0DUNI/wVD559P99PJdgFeNtTSVpWy3PdOKtvrdZtNmcFE
ukuqEpHBLslB/C+tSni+i2GW+9mBRROrguZwuHOTBmME8mftgrD0ZVaQluZWFckcmZN80wNpovjG
A9OHK+nn5eYfX8rTf1R/pm3zm3O2mSXvo4cQfE+4y18xIhC9H7ZyOtvE/H9rYRxxGLQO1QNYhaR6
y0zQWBixpIMrW2ONBLquDfHrgyKn5Zth11UWxDttaZP9UoHHC0J+alwrM4GvWc4vBi0+D/HRhfw9
Vqm0CRr2P+QWJGuqitXr7McBZWIiHVS+d0jIl9TQnSM2rTHtdJ1u2tGYwSYmBbDh/ajGu1J/El2W
gYAd9W7ZrLKtoZ/HpADRe+lLBnPDXjY0TXncQALBZjAzvTBqfkz4lUB8KXfxbKOpTCIBrDn1jsmX
186wwDNRf2v+PrDZ5awTuWICYGNH6GIIZZtciYlv8gdp8bJykLf6UhEwXCE7q+Fm9zEGCCcg/Agf
Wy2SaWt4i92XnIG4PuXeGMl1vkMQpoeen7unMMytw3U3jE+aQWsI51qLieDRYLMzp+TX+Cko6i90
31zDxB4idiC1j45OzF2n0I8OznSgXLRMkbiXIBNWZyz3ACwxHpg2oqThJ7z1urAzgGmXWu2Z50g0
BihBRO4K5JQpwTr1iisLiQe9/c+0yMzXmqE/6cj6m8CdNr5yo+BIrLSP8AfJVG94QO7WF7zb0PjV
DOAlSyUa2ROeT3jh907SYUcqS8E+I5RUYoTabKuGmL4YUUQ8KwK8FZ48Wwwt2nJ6DHI0CLH2S7wX
WCrvLtmKAHNDiPOxi7rxaV5hBRIyZGr/WTSpj2viHZ9nTUjR5F5j//+hsKQEq4e86fb3TR33iYP6
DPkmlxmKyOQ4uiXrIDvmiPuLsrQJYDK0sity0XllmNBgk5+RpkKFjGuWVgtOAgJPo2wo5SJ3UVP8
UAHvRXpjG2k9YLa8EKa+wq4o4hBk4L79sbzTu/qy5yjJaOOrS95ghDxOWpH4uHoar/Zps9lc7IaG
7DK6G3FMcYTdA2IzFlqKFuQPW+Ho5LFBpHBH9GP6U1kM2pMgUkIOjPNK9FY7YBXgQxpwB/v5xEre
XiapVAkaR0+BgwMucFcHxTf/QBPJuQrlBUVqYCNzJ0cUgJo6KDtkN+dbTcQcwZHVFHRUjLa/7qXC
gBUuFxlZNH+HSFs0JUMeuE55M6V53Zo0YPlmxT5HGPY/CdrAi9RiAEP8ES8DKcn51viCYIBXfxLA
Omm1/qjpufF2b/HRVT1EnYah/8xuf+Dl4q8ZfeOldEURLBQuqSMUsskaoRB8er6XKqR7vkpCV+01
UtWZa/0EyF/92Q2aQmRuEIGIiIGCrELrq5CTQWvcSr1ur5qAMJFKHcePkZgYEU30SmfYLFRWt95m
EYyzNP4utke+4kh4NnG6vpFWX960HSSHK2Z+gfJ+1iyI56YxdVsREX+zvKF5CyqxNq+DbRsO/8mc
nIC/X0P/ysQ8DWm5XHgKQCwq4Zb6pft/C/rzPctwJJxiN1/srtn1wnoACt5/xqLqdwA9zLt2vYW/
sFXqhs5orJLCPUnBtrc77Kw8xhJTYCExh2Vs3aLQhawoFKDOLXFAWBMnoRoTKc73aK2zf8q2Hx6q
YN35w341NEzQop/0e3s0cNHhx669IZarrgetP3z3C7prgtKN33z6RmWhkewJip8hQbh5fYcGZZVQ
rOt4FaO9+UijviCGV3yNfbl6tAyHUxMs7dvH7+4BC42KR/XHTES8hGVAEIwP4oXLmm4OyxTJunkj
eJInsNGVv76ROsaPRlIjfg3rMbtA+MFVguwJf0aaVh/+S/EzgmP5n5MVe2zoXaaMJplPU1qlIy5A
FojjKdVYlVp3VLJvwjPINB/EZzoLrbC4Ozg8RiVNsdYOHPE4glpb0yBkx8JFAHSTIT+fFdYm2qvR
y+W5Aimebz3KU2Boe3JUioFUX0r7cvmxrf2UcAUcoQoVYi2i+7SWA8ic5RIp0+oxXSLNkCd/a1Rp
hr7R9ee5qiMTLcyn8tS16sdtFad74KagcLMZMALq3KKVHO2eMvBLhA1C2lQcHnuyyeQ5K+mYy1AZ
hRYjClP7SKFUJN989gIFT9DWhufvFMITebscv/k+2Zdhkn1i8ovFamMO4U2pTe9ukWX2Y2h+EY97
exBr1bJdrVfTg13X3B/DJhmKkFoizScJw+BXfD9n1PVLs/ox9QZthfjcgf/9nvDAaO0j9+MN3VcO
dyx3f6QwV4V4P7TO1A8ItU5t2ytQTP5IDjl6heJm4ht/MUmOEnxZrWlf/OkvStiBFyfZjLHjatdp
ueaXMYtrriKiPl/vdszl2c6B8jeL/NErlybmWP8OIVNmJDC2+M3xTuecFdrx9csiJGES0uKjul9t
qMjq6OVvIpc90ExhPPk9HV9Qrkk4KJvKi6JHHCfCWAgNBJMrbbGA3Oq0Hvg8LZCV3QAg7hHmhhkq
WyXFAKFqo6xDh0XuNYqLpY9F+nzIGwtMfOd84H6kk0K181OGKZBOWnzg/KX53nnClFji+glegfrI
/pskmMwlCFKbxEUKXi5TCCvNdMe5QniySrAUUbcM0oVPGRS+dPcHjIVKY9ICtP+FHxaepYnGVBU6
cWkYPAaDZt+sTpvrAYJ9AjF1Qgz/hVCV6pmaaXJmEJdKol0tXRFjfsymDV5MjvAJ3NLZo+4mwBff
XIWJbvsdjNgNcPSzcCg7iS8eLqLUYafRzyamRLr5JzeET++69XQEHm0yqSpxdFXOeAPUrPk/DVcg
RCv8Bh5E8WKMrVlOc2OetsGRK7TuTe5ZoetWdnZpkiZBs+l/ZmeIknY5creGwCsi9uTv2x1hs2a4
c/6mugm7hk8d2kD5IUvPLboFgAt8gVuJ6kX5KN+dPegLr/c2tPGfREKzm0zgTMygTdTeHX87A5U6
zkRT7DOVilG72FaXbKp+QcSHteE2FbZwEvbiUYWHJx5cPit5gLcceKIr8p2g6o0SEjlgw1NpaImY
HXxkY4I5xijPO9iIKLKl7iQhZQWqoux8a+uSy0qSO6NJiMBf2BSG+EEsEh/sXAFXAdnFxii7/Kpt
FRXbfx8hQj0ah68FKcFJs0RW+EMqmhbAMjmSpU2bVA/xIFBU9rRfWz9YW5f3m9XwPHqhle+8q81y
9IE/+8wR0CS250gqTwCjPML6VBeTW8QE+iDeyeFQ/RCfN25gOOlZnxY50s3wp6LunmM0kTxToTL0
DG24b+ZkL0ox2ISE3PJWOZMlCCUlofIQRuXKjssU2LlbIe6vaNhkv2QJNh3AHZdvR7weYKM5XPhP
gA6HE6iUjZXOp5RvaCYjm9v/isL8jsTlFZ3jmY5HUfRGpK+vybCLfNrVAlrBc1xNqiWeFyv0dNAf
06zpaBN5LUpUl2qPNGET81RolNq8029awb0T5HqZM1jUCH7KJ+GfpvwspekrlCFBHAs+7vMIe1u7
kKEtWIOnjntIRNSu6C2auv63iE7tO1vpydsWXML8Z5YN9qbWhT/rxKeDBJ8TFmW2Uezc3ARdl2Ha
jxYUg4k3dGzzXDXwJFahWHsbxYcaedNoCW6bGYXthkBnJ2/0lCJCQ4JocHhpZqbYuRQaW2d9uJLX
7NrzTpOuop4iXv8y/3GBdi9SPAdPDROp3G07287QCzzbI15CIf2GubFgb6RMPVVZxTgr/GD4bVhs
EInN87mCtWP90manBHOX27vbZoFHO66S5TfAaoqIfXtUyqXFfvjGK3KAScRjLRpxJfVH+k7JghQm
laKPvf7dkaP+AMae91z9067japHCQUUvI6pp/1jVMc587XhERpEYPaCNvPJmXQ2BuiPlpquvDrLO
j29XF8MkzeXg/ohcV8GDM0NtqXdEbMEFcSudRxtKMc/YzOpgsWDB8dHQuV1zEiPe3IjJ6ThP0bJW
AVpAhBzj+tIiBtNdW/yDAPAlmAvD1t6ZlU0ywNIbpQOqZAxKMbZ6+ST+9L9/59ezUVXecr4THouN
ABGBjnLjhYThkUJhNQcx1Vqp6eh6bzTUUoIzyo2nELaygvXaUF6qg5QkWiDyq+KodMKXpzdWELQt
9NIAgSp44oSUKxh+26b1YCwzBYPLw6M6CM+0BnYx25tAXgPkKHoA8MzOfdbJ4GmONLf16UFeVqH6
mhyWc+f7gNV3D1QnuHvq87unuTY+fzpagEzvIlxKzT6qB2P4TSqVgWBeAaEAg7/RpfHjR24kfKz1
YjyhW53oaoXL9oCfZvZ+uTUMjnPBg+HE71IFhj/FT/SIbnjkFinRMCMZ5FiMYwt4hdJsTop4pC2c
VuLLiNnwTa9tm/xQrwzXjp2p2aPFWId5SYqth5QKSSigjUbT3Qan7Ziom3aDSJ2UXciyWifh/xHg
u0x2e+vSj5+6/jEUfH+TW66MK08j3GntUTx0bjnkt2/x1tlQ652z4n/4j5QSj4Np08npQSCOan1O
7Zh1DG5Hf3ld3SmcAO9pUP07w4KPP0akLryyi6ugjQSC69e4GkWcg7x4i7XP9BS0a45CsCj6FCIG
fNZZJ9GBgFP/8WbB4VwmvP67R0eks7+BU5NUfQjBdKMYfeB4O1/xbFpY3+Wfwplen4srfCfH25z9
3cvaxGpyH5AE8tKADCyN13AS5bd0acZtSifkdvDs1UniajWU/f8Ln3+TPE92fj7ejHUgHNLZDEPk
J6FLon6h/U6LYDle0Ot+MYO09QmcvMoTSIVqDSkVgCtkaO9qLv66NfvJci2uQ6PyZzdbDOtpnU0w
xK84n/Tlwm76ZrSCZGYFJjLMWuvVaDxtlLoq+AjVAYJW5wP0fvGfpxQZVyD93diHMCCiRo4yF/Jl
/hyi4xuWQ6BTyJqwjbj2EApOqekJ2nz4pcMY4cVQhucPtKCxFwVWFCqSiY0oDvXtkCE2mrsymKWS
ouzCqeKTAiNT2tKW2sLP9Ve8MHfA/DqQ+hrY5nJNEadCny16IhzCsIx6yr5pf8+i5VVkFOMeTJfq
n87TLIyZzryzgdxqQmMdp8Pe2wCGN58GcvxDkn95u9meElG6XfacQ7NbUNq6466ciIoLE0qPAaS+
XuMgd2LgcZ4Lm/aHcrAwibfLl6sPm+FwNwvHdAUzO+MO+Ty9QMOztHNHwbOv2+bbSe8AV6VNybCs
/KDhnHSX1VhJSgu2V5aDNc8li7q92Bgs15XtBg0gg0wLVuqV0h943Go0WFFhowbtHfdynlfA9UDk
+C5WXm6WcrKDyZ00wbker8ZhRJ6HK7HR5Y2iLgoZOvJyqrI4DACIsVy+D6NKF68auXlWR0Fp3Utc
8uvOhW0JRgTNPKo8/D7cxAG/TOjbG29EC2FuV3HCwJbFu5efuCycMaQ6Pu3TTooKkWeFt3IUrLYs
a6ris4lWeZAxeN2W70egxjbuaIhV9jkvU0kDxHXdr1tYCHAMvUZYBXnFIzoSjtT2VU1Xd5/hPfum
CkMU3u/Sl9OPDln0VwuWIt0wY5v/Udx8jFRHON1hJ/JCu22mEiU4qT5hJsrjRtR6KP4lE0Z6tUr0
I23Yv6Ph4V1Bf0YPQkgV9DAXQPiBybE/iworvx+u5MgZ7tw96LY9L/XN8CeKMiwsp7koMo7MPQ+f
p39eVAUSpF3HqvkO9ElOiWViEkXFYQO/AZlN1XZEmTqWdgv+kB3jQJ73uQw5b+kU4Ic9iPVmU/P3
1qmZY7WTppKjHkmdb1KDq9/PnyX06fM9Pq+6aAKyCicmyT/5raYL9B4zYCzYos/zr/3nDx8feE66
3O18Y+PGVNZ22TYfyd8/RvYJyHlbkuwtAvkya0/tKjdDp+U0i9iQgmyHmHVioVWM2iSrJbrEHy+C
jVniy5UWFNRkevtfvQ9OYbOC0OQyuzqdyE6Cq6yBUV67FOej1AO89H8Ww7KgcQytGOXSyBg+8Azh
lMge2WvAt4vpjJbDv8Gn96sAUu43lCYM9R/2a7XD/mqPh3XqtNHV3O9qHnswR2Ienwzvx3EQqcuV
htByrKf4XZtbD87FAVB2VeQMrr1EmhvcD5VuGddZl5lnidmPks9SmgpGzLSlrOm7cXlbTHZrVVTa
wfHOqwnbsq9QAl6CiaG3dK6oMX15k85FZM+W/ozMd05khv9+PRnxyycEd4vGTRrCtsJgMiEllvsA
oYm75gw4Lx17E3tfPEE86xlqcvTIUMnhCg5SgfOs/KN2xVWGzHk4XF9bv6HDg0i+Nvi4qNQviF9Z
N8L8KVCMhqw29klypGpEjlAp2L0SJP7RjcbhToQGRrdxVsrCPEcQP6EFMAFs74UzpD2OJwY/7LKE
SJ31IJWi0UCFPVfPSL9BPiSw2f6vlq1w8yQ+qkYG3FX5O5uRhJD3eG8cKzp3F7haCXRHsuLKLg41
c9CNKifKfF/4JhJRvHxc1KdGRLSx/Xw/1UxQ1zUn/w+Z+lj1flfJeR0UOdsfes1eJoan5eDDZb0t
P0tu9jL6Xoa8ZB8mmozUSpvmHMVoAig/4YKCUikJpkBRNhPRsWZ3Kwd1hXzTx0KnajxREtxOGPUQ
8CwtKWN+/hGCGreQaSUvdcbZIaMZw4Vw+aOLndWxLqAxFKZDZ42QLIOSeuYPfjXs2RdSznDvvJu3
shMXP9samQRFecmcjzbsdU+jJKLW7J2Jv7evLhRc1ksXQpuQWy88Ty7W2p1rDszOTs1vOKU17+nw
8x50ghNUTX7zquW5xGZuTWS67lelKy3jgzCLOaSOUYAnNFw923QPeNe89MAUgMktkZqozLFJv1DH
lBPqDIXK5gKLJBgZwn6V0xIs+OqoNYGWaz32ESwg2rhgXHfIBoHDNicZ6GBEstm1XhSgCth2DZC5
UclwSJYhjw0IeQtXjA+Jol9CKtt5WZ/5WKaUSJt4TmD0umQeFibhulG9UBCWjapMoqQ+lY6wG1bu
CCEz9F07CEIzjpRrN4dyiVA7xNtQUlIoKDxFrMqHEnbXlvEtA6s6uSaJzDh4+a+dvFin8bsYYtLS
+G8L4LND/weTxrsLE0QfymBYg2Kdk1pKbqctvuZZP3gAQ4Ktl0PTZVMh30mqrC8nQ73JJrbGMt6j
wjGfPpNBBisENMzRcMiK/0YEzBAVGHu9hlOV+zS8bLSFHP/N0kUYVbjR6IFTaTOK5apJm+1EhIeo
p7aFqnl0SSH9k7NcoFECb3jqr1mO2QbTMXve7S6tlGZPKR03hYzjpb0MgaYpssdXp4Kct6D3eps/
RXhz1HKrjSiz5JxYdxDApiLWaMiDL87izM6ifTM4255LItnqEhGpUV7ty+gwqTzwCH1D0dtz/XMq
PvRARBkGjZQDgYFMvXSnAeRKf0rNQJ8J2ho2w8qf2HXkj14fE6dgve6gg0kN1xxbVeKQIhhdA/jp
PXleunLxqV+cF013Ez1y9QQlSW0LzS/K/+hpcPTsCiNqt1CXOO5+yZlf1V2xhD6K19/kBFzXpEh4
96dKvLqfTvdF1I+ppi/o1xI1dauQbhMmlzAK8b6JOiuKvTcU8KqbC38LbudFjOpQqTFNGrOwpza+
CLpTBf0YvOP5kc09raYPRsdbJ1FHlje9qbXsL86Sz/zgB137fzwMlm8gR70rTAF7FJb5j1/to04Z
RLrbOugpPYvr4/caCVFfBrYmEFVagetTGB0F8z6RC64bkN4btqzaAASRT9MhX7V2seOUGsCrR9dU
GU8eAwi/qDWe2j4ommWTJxeoSUY3tbtH9VA3L3C2FVO67uFxMKlpQrJLDHWaLM3bW1QjCYzTclgS
3BmmT0JpbKqzAiJLFbluUjNPwIBMjUfZHv0tYY5yn8pULiE4H+H7/Sxs180Me64pv8ClIsAzCGEx
LA3wuqyW3bca/+P8bhY10aw7BPC5DrK9WyhFB+e81fMPDXDmsXgPiG+94Fki9+qj891cnD/CuqVz
Y6hW0jRZAkqdh4wW5vXkmFnUiOd3ED9z/upqHHD3JFd29sVms/LtzeA/Rn1osXTqAQm0WNfsNcdv
28EhrlRgwfomBe/9fXSuSE0VXG3KgVUO2ChKpLGSES8lfeejk1ARdqJYwLL1AafezdK1rZCj1VUW
2kuJs85LPvXUfdp/kai160DRy71DSaIWHbQocKXnwo4jp8N3YNn7JS2pDt87Q8upc1dsaXbDl7o5
51y9RD3MuT5lFEAnegpPFUUp+LOZtRSi/pBc4la2LrIq4sEZMrT4kYq1+Hym4aBeRnxDCCVy0rLX
Y+QmhoY/V+IQkmrdCuJZyMHr9q7HyXk78bCfpmG899cTijRz8H3tPYgpiLzCVWwPXq3GgmaGspfr
CWfkWHnTxedrc6oDZkpUxWPkEHeeOHiitiK21pbSXSHTl/lxjBnNSfXAE2p0Mx3P4/9jvo+wJbrk
4AKzVW42UBBd3hMJDLf782Dwxf5ycqOSjhQayqQRCoCxcPCZCdy60ZlRWvThbzXtH9BUHRiWn9M/
xCmWTf9W/GZ+aH1h9jqH9o3UXWCjL58/Murb1qy431l9Ncpkcr6WqoAj7E6cGCrTKaDunS4xhLKm
d81SWnIYGfnqCsAcY/B+i7Hx2XGSF4ff3WaH0hvW4HN5jQSxaaWYx3ENKiJbUa1M31Vzy8+SMgru
jDym1uTkzmVqHohRMfzqEQn2oc27dSmb6REk4aqbG59JyTA8Veg3m2ZJaJvhjrjxTvYdbLHuuHAm
XmGsbLGetWq3/i3JFzJdOXny899PbQk2nrKAPFq/EwE1wBFI0ZNWSy4dnImF8onhhuVQi67W0c2H
8qfHDMp/kNhziTA7F8TmIZphuszSjlLiKcZFaien8VBECYLduB6tHQOXyLxCt5L4AsMnLxhegD5x
39oANElPfRHWmaRTTQttfpuHPsApM+mENnH+iVQmT7Am9dXFMmYuqEeUw/CvXe1kdZgyVVX3htqx
iWhITTN5P8U+XsGNScre4l2AFyVopiAza1UV5VraMq1BHbzQGcjQ+NP6aEGI2m3ZMyiRPW6C5OW8
Hb/6Ffc7NK0VGJKZc/cWJhkO0oxsy8Phb8FBflGu6/fKcKAlDCjleG8wJF/u0qLKnXO0Nll6P3Hp
luvqQfehZO9mFqmoLydhrNi9ABi/maqgVIWIJjHcbEsdwLVFFqZTHQPtzHoOTQsaVgGL9svnhdff
01aYB7Z9GEbj62PrclITHi6Qy89k8Fee2jTqMyiotHnd22MTnww0H9qf2h6I+gwCpq+ouKdna1rx
1Y+XEaWbqgdFbnFEQEVEwzwG8a1hV1lErV6W6LIIb0+mU2hg8+aq+WUGkrebozBCSGSmILoGCFIo
Uu8g0jyw7Cje/5Egy93lkx5AHi3o0KrMRx8DurWJD6UgT9TdShFA2QVD59X2c2IRnFZ57v5MpYb5
5xfARohK7HEVGOapUOjTmzB3F7aM+pj3adN2LIZSGAaIFzsnxbX4T6AWmzQnaaEPvbA5PnkIov3H
WMWytdWPaVr9oWfnngOLj4/jfR0FN0l0RCn2J5Ii4XFZGkcLGitpe/NBBMsNIdLH+IDkj3lArrCo
3uJ/YXI/XNXqrkOUlbs+M4koq9mKCrFxpVZiGp+5yhwgdmBdFU3/khi6Eyo19+iXcKw5zFonE/3B
Jz+FfVjgf3TjluXW04r4Ji9gsuD2UzqVtj2ByqqPDmYB8qbov9Opki3eiSmcN13KahS/Hz6m8tCH
k5wTf02OSHWsSWc4u9Zc1RxVIH29qeKxY+T5EjrjvsYaA1ElLUNgV0Nw6jqn3lgLSGjqbcdT/bZ6
Q0k6zk5C+7Sc/BX0B80oIMFU2lI9kpNPoQCTD6CJFO0Tol1sMrd4uTIDUifBSQilMvRjdV+eglZa
V2HivAitQJqCa18n4Wh+s3AYLeShUqh4xH4QxPIU67HJVP8azL4uUXIGS3zLCcUYQxnEyJd4KMtD
+LBbiZVMj6leqShLJolr/AQSNO0TcdH16j5b4DfAt9yMCW0hRj1AVaU1JC/V5de5Lx1JRSdRqh6z
sq3cYOZdqBAFWouXCcVP30R6+nhPtqcFlkWL6hiqbsV1BLej8io0OoppImfMP+HZT9D57UTmKLJz
OxijVKFQJ1MMkwWpcY66Cu/tLHEzToywXeM7wSLwOSMqXrMKcxHkTKgJNT6T2MF9qTSRiUgzYm9k
NMEShuH2dtEfeMZBnoti6W2ypqYTy7SVqp1nHuI/mUMikgp40cFGVdx4GpDHMXAjSDvtirNeK+kN
TEuHzRYbVZwluez5d3hdjSxo46D9qSumpD/L+lJFdzaWlQqoTNYcRu44qTZI09uT7Dpk/7vivwj0
FORoiPY5PaNKZ+VlGSOMKQH7OU5qmIQZBPKG1HNxCBqfL1qRRiyyePiQEtpa3WLxB3HZZkc0go6P
Y2X9db+1lWS5zevr5uVIHly7qC6eudyrdZpjox81TbPbdYDz/I8yvjd+Kt6J2triTeqg6g51pctE
EHKxbvpPgIj4BCXNNiiqaFu8+pAvJCtkH6Kxhxol/iq7BUMSOgp9omvEOyehpgUapvqjEx+es2jf
MKTfB39OcYKwK17edJEWe6Tr5jB9ScoygCJikTauHky/+TmMn0KUahaCfGfkZnfJ7rJ3IPqr8qzC
ri5itb6zcBvmCkLssdA/4/h2uAfdaAHsHv9mXxMZkrRdYQX2EYpdjBXYCg4r1oZkjCinR6i9zVkI
rt+82kFe1vhOJ4f6vG43PePgUIYpFDnXD3B+zV3iZfI/XS52NNI6c2mSndt7LIv2+OYr4uVcRBLR
ayRTl1STw5R/kcwajUxc6h1auG7DHJ03ktAzVDXUmi52+xPjgrocY3fM1Dlfn0oadPNnB+02irVC
nifqUPnI2GhtOknd3tXRVOqWRDrS+Cb6/5vU8FeBjNr4M34cAtTvOiJYpNGIojD+giDOec40YG+R
zs6UfdnBxlir12UAxN3DYQ6CRyb89QB28/NGwHeqoakPQ3PuM8JWTaBhgfjvMWcrp66Ji7eHv0Fi
3U/Gb8SRDtBpe7atx2SGdrqSyzBewIITN/EjFICixfyJ1Ugj42QMDfeHiFNyDSI/45wnMS0EoS+8
4lgLjJHcVRkDk+3dZKjGv6LJoppN020DpCspGiv8IC6uZlPUDFWHviLAv3VwGa3igDMOJWFgBB71
ItpPlJT0kjtlIQ2k1vAv1epegdidiJy/Cpim/ropQa3+kmXVzom2uwt1pm5CEDszZAl07Q+9km/o
8qBvTk42pzSAVa9IIlcSzH3IiNbpNBnmjoqCX/NvLZqB0v3eRm96Ku0oCxviAw4IpFsbMqHg34tE
345d6Uj+JSUyVKdEWCCOponwUEnAJHBMHmyOBNEvnDpnZ31pYcVusi6hzV4RQ05OSaICroRsZbEc
w9MKBMfQleC05bVOrs98HMT6b+W2fZksZItKiYnVmEbR5XjWFGdKzY4GNg3a2ok/cSSlNeolKOfi
49aDhp3TqWnbgKhZ4+fUHzmV0v0KV/7id8KyRKVtnagbkPDWyZknTipWrR0H4H7MGf5QCG/zTe1p
+6Hb+DoUqvuKWfklBcTsAqWR17nPgvFasbU4fTYfC9Ad3QihuOpDZkEKkg8CwoAvxGXJDGdeZnFn
+M+rwXcGkbZ1K0s9n6DpG5PP6tRRREbc0S69T4EOPB0863HrNlZJmnfOasU2vy92qM9zeecCcwl+
chMi1pbsh7Umx23ttCosCVKU+QBAdG92wjjfcPRYS4PaBcK2EPIK9Am8VROBE5YdGH5YMLMuf599
IWrgGG/0fTxiGIFrOo/0IW49Bxc/pFxKFz5RZfqBIjU7m1jKuDn0oPrc+gbATJzJ81KZAuMqpllx
EzASbU7ztlHxrTj4kR6c4Kze/sX8ivOyClE5M2cbgF7s2GhLNlSrQJFsE/51YLpFcRsv0WBa82wT
xRQOyjvQijsahicw8YEECN4tPNg+EQPE9Y6aZbCY6DGpNExSM2FX54q5pv3DYDHByOg1kmBGNct1
lNkQdj0gzJWx3XYL7b5iz6K105rrmXZU13T/wtt+sMthiVALCPYpkbHC1zFxYLa6R0uoYqlboY/0
/RBPq/LwnVt+shQ7Ad9uOBuGxDg5sl9vN7ds4EZA5+9wLP5gJnkS090Ke+P7ApNOAqO1x3f4rJXx
9ILbif8zwoCucqQyrmFAjIQ+xh5sP2GK1xjf9dwGkNmcnw5z8rwHRWQx9/LoXysc4bMD1ocGxNkY
N76HUxRnNKPmaMY95Im46kraX+JY+ixzyZD9Ae0o135GQLPlQ3NdOo6QHTwaQ01vg7UHx1V5XW88
3KZyhTetRAIwmLAPh3V8yXqBuH19he0War8BGvex0o9M/ipJtypIb1f8bTEVADFIVZTsRvfiJsRH
QRjv1IyOD3abfNpIYEa43jQFArrkzyYG4Phz+3n4RwWjdKJ90ovnWd0IeoiJw2p3/coijApVrFhl
IRJa9KyLrARhzTOuS3paJziOox4UMnIvkbtTCcQ8z1S4kzh9CH6NsvYca3XT32tSfByayHegi3Jl
O5QavVTIB8mgdP3Opc/mFtNwjtLdOWvG3AIaKnHNhJhrkuOtxLmDZjRbqN7pEP1mCF2Z/uqljR2z
Wwp/R+ZAa3T1aehVNefr6XE6typdycrD6AUVzC8nk+WMeLwd557n/5C6xZZZviFhxFL2D8ZOvv1g
7cV57Lbf7tSsYU6p04zR++jKB2sb5r30cBZfbfxKHLJiZRbCMn23zIR+35l5iS0JmLzIc3fDqOLG
9ETI17CcPq1107IyUwkfyVCn1c2XCG2FIF8/YFkCS9ZKEDCuuNu2009sMxE9jdLG1uthds39rmJV
JDoJ77H05FdcoUkzvPYsMYgWMTon8QHUEkPcVN76vyVDQv+5teTqj/+LU3X84RGtWse5ZJ3rZljf
LAoNbq+DPXfeyW7YyJ0AuPLeYkjhOvEPzpYJqL06Tec1MkaxzLtogb54IT8LgvrGht/LHnLFLabu
G/Jyc6UZT+QKLyPOjZYHx5irr8BA5LJVNHEKxHKjqlzREC0ORBh9gYjAc4TWKgUWyoLPgedKFW83
o0vDzlDXt6lrQptTRyPzMHt8dywa2MXyfbGJUpHE+9FNzLKWrinho/HlqAGZjS4obLdddNGRYoHV
0IqUs3FTKBnqYlLTsg8zOfQ4Cp/dzh26a0Og+8Lectkv+k4jIrja/S2ggX6abv6X76GTnebIURU8
Ximf2MY+/K2ut4Z8aOFMy+y9NhLAaFdkg1gZJu1k5j7jB6MAJqvswzs52oIdu6CpHBWfQCQ7Gme3
xgaZH1KbXaCLCo19vtr0FXxXHo98RQepjGDBFr0AwEwgwNoK5cfNjKHSHwFiQSIwObTWAdjdUdta
4BaEE902zeb5QAqahU3/xULKhmmp9UTpHOF2EMH+1/nu+/YkXqfsB+VqEcO1OAxX6qEsL6EvrCJH
l/aSjQ+33l3zDWR2Hj2QYVEoy+cdGv/qTet/mOBK6yvL9xRxBPzqYACjLwAkkzDqbuTMXu+aFAKd
LEWxwCrJtZUJF4y3e2P6d+NM8uwDVEvfMG2HSvq/xjnpaQgHiKYkNWmQGQpMRgI7nVQDODIhFBME
lVZq2/6HaSja58SsO2cnYuaeYAh5MylAPAbE9J/QHwIzmeiYBX9394PYXDrEmkYNilTKCDkhRgFA
0vhByBwJo4p9am3SShSsIWyfzGzdBD7xmBKaI6zs616XM+x0F6fIEZgeQPizsy1VnXvkoPkVjoHP
DXX/NdBGtmbgAKWwF2sjT+jLK0YPIBmVJhei7zVHf+/az6fosKiTaN0It7hpOP46bFqYkDRfpOlf
kPiRoZrNlUSTH5/lc2DKYPuEFSwQe2L1qEPme1c7K3IshQ/CoQjHKf9kiVOcrqtB1xnhlRO3vk7o
2dZnuV+f4k3SSujHx7QGKcU+JbVqesW4GNl/wI8iPegDayymEjubhRFbh69WmnwjRvzk1Hkl4XyE
2QicvYyfW3b4ZZK5YqhyM8GYX5S8YmC4BggIb4P6MrFcW36CbryvQkMX2Ssbq8ftjnd/HWHFx+Kl
jg2s6cRbXxe2+l2//eN00jsLo/9c3hE5hkQAjXiWD89G/x08Egg4Xy4MQiBMuy7WnIctdKSA4Yyz
ppg5D4VC/5i/S16v5QgTS5s6r7v6xrosFO/EpFwZ7ZLoLIf7BepOJyJ+k5MmbS8Q8PL+R+YIa3EA
9YFK33wZpMNeE4K403DBO8P7vzTwvsl2HnBiRxt/40kuPyWwHjK9cU5RcV1eJeZeG0Sq0UE0GqoR
Ud0659w3WJKYlnvkOvyyaM2FK5KUZ8H5XZ0SzjSlbF/hRPwI7VCjBES4hxWqERSJf/bDYlg0ymxb
JVfRsy0Hm4qGgMbChTSOm+fwkigO3UhMLjkJzDHEmslGtRScb040d7OqjRxmsytheTF/pRoBlQ0B
2XxQ8W0J5AUQ1+q57pg+Qw0G2rMDWrjp57jO/m9EGDjoSXg3zpYRkSP7an9OgCKjGznrSIYgCi4+
f42ld3Vj1tbViTnd2XytdYWIappeqpWwzTAxq9IwbY9R9bEme0VYeH1sgywNsc6WEpcBEZtcbo0v
Rm8sf5qaiXLBhDLHC6WJ67fu6ed7e5al0ntdURbXei4V1vriIi8bpDR8bROappfohr/nG7AKdLxu
dIL/4WvhuxCecqTeUKj8XVgu2sD3XNG3kD4dTSy1QqZ5AyBlV98z3fzpgGXA45sbJDqG/GUhSV/e
1HHQM1A5NCN5eRKGsqMXIj7OVhppVjpNQ6EQcvWwJVds3rkEO9Gu/PUbBxZ+Rzr3B6oHUv5DBa54
ZbbuqOu0KTY2yrvZ3qeqghWscMu7YXUJOPJ88r1JP2frL3Z9GfWEAAb+QPVlG+ar7fgKOh6PKaqg
ByQn5kTPVigRwI/sSovhwWw9Q2OP83Et35RlNFmSeS53D0laV5JFTZQVTVne64NGPquRYuy56VVN
mGm8cKguAmDuNsLYmF+Xkig4gznCYHc4rc2IjbZ7MqA8/OcqJK0+EGBXAePqOT2O8EBjT9PUYoEU
o4PV4x0kkE1L+1VDnLJcavoIyirUL9J2Rz8HYjMfd7/6V5pyVXDrn6M7NDJxwE6LsqDDjrO80l3h
GShrB3aAbvU38WBmro8nNNZYeK8wKRHqACbLITKu4SCxUdUGMtpGhlWLhovVUTC5iw36QtVHRXNE
GLh0pQsgRRF9ZRsieJeDuzQmletCfQicPXRl9MDmH0CatTKCYCUz4LAc2FuF4ZrIHtd0Qqw0jSq3
UwtQKdx4mCEBqDNR7YmT4OsAUXmxuBATli9MrHzV/sRNEUOtJkcu3deVnUIondR9CR4+p9X/U2Iv
O1K/mixGh9mp/7/1TWhs7BeuUu6hr56gM/semAUXSXomgQKVhOgucgwlTTUYBMmyCta2eENkfoAw
PHtK0Q4JuMCptytpsZ0cUsLr14soGyiYySGnAmVoiGGmoyVHaQqIWYCdDdpKu9I2PoviGO6GZP/l
B/HhIFU/EvCpcMJC6SHgCKyncnF3ZSgw4UR9lfbBIYdUGjW5dzGdwJta4j24oHGzttdonbH335Zo
j7Lc+OR2I8WTt4T+hXogmQQJp3HyNPCHyWZaSaHQfGMRVM8RPCMU896ukFBUkWRudsUBOTE4z2AG
luffQe3CDp6yLcwCMB14aChmEFBN8e+sNOhVeYEpiqcNiL9hDkvtO9UQfAJExPu3heOzDXYc3v10
l1bxoW70otcwabJVxEIAMW72TrEHxmWj9vJO5sM7UVaBaBe024dIwPqhv2SAqKBvL3+0/HLYLCXQ
fUVeuvWXldSTY0idWgj7vIqlLA8Rd+5LqRk+U7FwYkxVbZu0eRoQ/MZTyBIG4esKsQhvH9aoHQbz
1zRM7Q2Ntb3QvVf3IDe735D6lvgK+oaSadyXBJKLUeM06Vhcl5Z4q0DWXrl/83gtIsHWj7I7D9Rq
mFqAY/ytw9tT18lp7rumkkebmrocdckaGlGC3pQGJ6HgCnx3C06pon8XdIxVetSyOvM2ISgFwmPz
21hLAFldmL751ZgBD4Ut4pdc5S3QJggCR4vj+/QZg1teIkCkK9BLZWTbWLEjRvH4f/RaOk76MI5a
B62SS5XFB11t3SYPKOpj8cd3IvlfBBls2jxmp1hHtUvuTuVOwiAgtP+MhTD47fD73LorkDzRUL3Y
tggu0UugyVB6q7HGExo4faYh2ycn+jVbOprVcMuynyQu01zyFCmW9zh71FyTQZvssp4B81SDJITP
Q3FmPpaBwX857/nf8ZkWVD9raDJ5D1bH7y1YL4VtB7TSZakhNkr8iPTaNs26wfo0pm5QGrJhVcDv
x0sVRup/ofGczGKUxRmuZMwq+jz70wEUQWypdzThbHdvV6iSH7Uyxh//QIkcrym8fenUJgDIZfif
1jwUXZr7mpy3jKuQe7frRUnZazXFSdQCDEWTCaATzjVm1QwzY/sTvvltIETRYWne2a4IgcAhpotc
D2x0XN6cpEMoEFmEfzQh70LoChq4dyXctj+DkMITc7jseLZROjDgTFVmRsIQP8DDz+BCUGKOFojs
Iz3lSItHkPB7UN0aCh4vPiI0ZvacEQqDHQoGsSbgyjsiGkOoP34rYTVtByTRvL9ZJVYiVOJX50e7
spVyNIXa5hPMGR78ehkGmIaExwTQ2XEtWpUq3uJgU/xnFzYiSwIaaRkYxWDOIEoiZ7fH4QMqfsSg
V9cpAB5+DwhtFs3tYuXCX/0t75XXx/HpTc6g+S2m9Iya++XySGoK0vkr3BvExmbhYNEYvtm84Xj6
q6ko4eB0tcLnRY5BbcwZP2FFHvuqJMpFkE5G4n3sbPVoqzaus59aqkkFfApISuT9SUbp5kWB9pNG
Nb3otQMwpHSpyG1U8iQkwnWWz5gFhQlVXTE+CklfPifyAALeiG43Oi7MvfomKuLjGd412Wjmejs1
zQir9mSo5+dPFfabspCNsMtYD9YENPVz7o6teAjEmYnYeBivRy4c7Dk7W+/W9qbsKPRqAqvUBSzd
VTHKD9Bw6UHAKpON/8r/SZQ+nO/CBjuTmenXGuaV2oFxsJZe1Yr8R/9FQyFSXWXnbxKVkP1bsewy
lvTVuo8vQk0hcgF7mcV8ppgMxIxD4UVVn+9et72JC2jDAMVb8bmCn1lQYzzFnP0jlJ0NZt+3r+Ll
pTKh81CcWCF/YzH8l0ZTYAGm7rKWG8GLbLKIXdsGOYx00Sqq5POKn9qDSDl1fBNvzuV8yqXT3SWG
cjeztMwEJRFTR8LjWzbI37BkueqUgqpNCVcD6xMUno8RkTReFi0FgpzGx6rOPhkiaB+GTnsVeiEk
T1RZhiHQT65XsaVCCW2RlGFSiSbDjIIUDniB4TKTlljep8FEHLIcybegXFnh8wgIjXnFbsrqGBk/
/DtklYd/dii6lzSPDIdEN3bzx6sF+V9cptgah78rdqkr3gvUKJwfw8Tu44ZvtNyYkT83zedMl9Xg
bw5yQZGqvSbz5SLDF0vz8fy0aAGHH+gdzWk//3DlhksvVfbMxiswVqPbeMv2uGGiNeiIUrZO0Ha1
w+XetVmeEwQJVr9ejN4XiEXAfzpC02Ma5BAWLY18OwCCtzuN/7bpng1ysdf/3lxEM1cC8kO0wsIq
qqGjT3WchIMf+cESvLucmOnbNfM/AFvOYx1RykZoZbyDyaRuksoXDW4bxF4lqLjXLmc4bRQQCbQd
op9o+3u/Qx52BlUV0AwT9uukYDt1qteMG98MtmFJWLohWdrsE8q0hO+AKO/qjB4rB26EyVdmz5/l
PApLPJvyDoo2Z1gM4RnXF5/whtpnH2TM0nAVUAozAgT0ewdinlbgX9mM8CSQA1KzRMTK3WkxCTKh
l1WZJrcxrZzYu9C0GOnBILFeKpg3UCk9itboSekg00ZIOGt+dfuMAdYs3F/c2Lb71iUPkv040017
uX0l1zjvymQq1WFZiiL+VhDxRIjJsHwO1Z5f4LYE7pifgqx6tUE9XVO7t936qGqu0opEMx7k4kl4
P5cIsaTG3iJW12jgVHZkLmxBV9C6B52sz9pwaMu/F7JDZovgsiGplaGkRi2hdtdOUCfJPXVHaPQm
9xRTlWvijxR9rIJQXQJGGZqFaVMRKVn11Q3+2gfN9NkQSGBI9KFg+/kGtIP+yn5JyaQm2YNCIDdd
pUHjxywpd+aHq9D8v694AjQ5X+KT4ruyndLilfErR/ohiTcd90pxh6Dxch8nXgD66xvEtzhsNX+9
lGV0pxJSCnwVZU91t0u8Us3ek1OLQcR4z3C/Wl+KYqA8ffNXPuKxtOmPxXB3a060pFWtLOywdErm
p0T1reof3O11tcWjZQbRPnWQcNuS+gkd+ee+op7jKKDFQEiILnm2eUmRNFyf7POb72RxuyQwxoGp
NMUiPtFc0Dy5Z9Oj3iqIaXVKjENZVZR7vjfqtRh+JIzlWkGo3wy1mn++cOlTvm2sw8LytAuT8zrX
ouAX+6MFtr3C5hE5mmgmx8AP/QP9Lwq3b0R5GGC/S3SamDnuE4G5QPIXU9k7jR4Pt0H0173Xsn7B
Eb6gDbuPyR/hW4Nmx0/ZPXIxcSxEvK2hDaqCaDb6uwcpZHRfV3oaEZtSeiPb7T8eqJ3BbM92o8hw
u06OySjeQ82tzT6iM/FG/5sbt8nhQlFh1DQba2TV5U3ccqGQ/w+j8wXQqSwbVVwQ42O5Lf5rPEFP
HQHY4tku0w5kPllk+AfL4JsVdOHciMqumGRuQRj4g5blWH9JQddekXbw3xBrF5m61j97G5F4Cvu7
FHVUIw/DeEnZr8Th7Fl4b0oO9AIQ1BebK/Of8Y0cFqUwfyvqddbJfdnYJMaMOQNXYOrBtsVFz6iT
7Vo79kb1a1VU3LOzu6HeTZYV1QXT/rgThlFzWHErVihuagA86vUY6JAN2Vu1Mu1bt/n0ssSZvRqB
Z8Zeci5MogObiWK6GYkZct87QVWb18Kxj+DyHtSNsAU0ff1VfkIB9zlV7KrfLZnL4X77TteDLQHi
6IbWyOH6Xh0mQhkhrSxKmxYsXcfMAoG13WemH7MNOXw5aECM/fTnpIBNPVt+cU77jtjSxvFDENxf
+MkREHXWVDgGiPGjoJOcQEgR0DA4+YUO/QQ17F7Ch6smpCzoQgBRrXlHTSbyZSpZVKl32SvEdxCg
WtJ/wsLXIeKvTHdM9JEP5E00sFu7PRdgw4TypzNrLeWKGU9X/DNlJTq0EKUmAhqOK1G+8sGwnZuh
Lzl0wCj96Caw/Q7Kx/t6voMKBVA5w49S4jdEzAUCJ2rBebR8M+K/OkFVME94MmaNyDU0q1GjiIhO
bm2UHuyK7a8eIYcU8lM57mgpOis86hpNGBsD3fMlLlhj6ZcRqduFsJeYM+b94/cRcttUIDTn7b97
ZtLwzyDmdNj2aZYVbVBoV221s8hHycvTFitC5R2jKG1uXV/Vkjy59KcyBs/dOGyhPWPxLF5jCg2/
ZIY/OmjDeYy4NScSyCuR2tIxJGTFC+QVu0Ds0jHOPtxzZLvhJXzGYWQpwp1l4Rl3ID5HhgA7777b
iAUS2SFYUJoLwNRcHeDJZyBsalaU8jf1ZfBTo7ZzBtBUM5aL9hvsUnQg9+HJnb0KtGEFP+Vt54Kv
Vg7K06pyRQ1W6a6GW8SsuFkFWNmtkYdE2duo3LsRs/boC7hyhvcuALZrax/qRPdTYRbTWOj+F7eA
eMdSK/Sr+q1b7PYReUFhGXZ/hq8FTmAB52g4lRPY4Tsk8kmPgwxP5cdtQ/J8IC3LGq2ISJoOKqod
O/w4IcO4Pc1EB4hU4HG1gaXuaEc34yO0IbB6g5E5/XKB7WuNGcBLAOnwppxwlXTK0/KgeNU7fNQQ
y11k4J1aobFhiE0rdfPY99A7PgoBT31J4GOCRMFlzsUEv28lynhQRM1N7q35n0ktuC0HNqzi6edr
Poyo4hsdQANrpORJ3LfNdxZCWL/OM/V9epatsUX7geFfk8/nBiN/7sTzVbB33n/QAJYPZoYXhoTK
iyfDuqt2N//jH6dKFA1fiq/8o5KKY2oSorDGVIBs1gY74L9IFXZVP8giNEhElc4rB60+8UPQ+bdD
6PgBcgieUmsiPG2gM/aaTLeNCnK0Q5Qc85h7nnzhky3GBqWPEUuNVbJt5CBeteCFMVaFgBPIq1YX
ll1Pp+uzVESk6QqN9DyRMthEY3LITV8n5VlP5B4v2itpBLVcPPSPfrlz7k0PpLLNaDudLvVLkTBM
oBu5ydwYOKF20W0A5Rvv6aPyr743pnW1vKqwTkRYbvlsopTtDI/6qyjJQLxUBCVsSAwLPCzeFQit
G2LtWs5YdGXv5Z7gyi26Ktmang4ZCsrfGLcn23da/30PaVNdrlXzRXPFY8wOor5x09m61kkPFdiv
YCQw3kqzP6Drlf7eSj2znBwfhxxt1A/Ie4R0Yv/9vYEbpdGaY5A95ScnmS8quqgyQI6Kmuc701NJ
kAoQKCbD79BWgXGccZNJkS6F5nD8T5YWT9svbPRt/3ltlBv4lo3Y0zP8bYnll3LA4M1mGa6rNcuZ
eMPTQU833PEHdp7iz/uLk47j9A1LTfpRMuI0bs/6826BRc+9rPxNBYvtLkvpYZOwIiYC8+TT3X5Z
ZdCfX8F+uG7rEHYTyJ83krSIDDAqARPdjdetbKir9irLCPwubF9W//tdIdfk6rcA9PB6wzWOHI3q
Kkgpw1YRC2kCQohKRltrh0zrk8bLXColKA2O6PWjGs7MI3gZLFSjpD5b52oRugP583+3rQlsI2va
BRYnwmlh/fqsFci2YlNZ76cN64PZY9QfnrKBN74+v5B6p9DCCO9YN7QbLNUlaB1glbkTR2uBrofR
6O24fkDU3cMlK2w43VC7frCqg1cZpeBHfTpU/c+/6wdDaC5rvnqyRn36zipWQZ+vot22kRPDPW1Y
JXzlVADfxvFJrv0RZMionv06wUAijUO7PgCk/2ExsJEdZAq8rAD0BvavztnLXvf9D9ECrm8+FZWt
GK0Okx7NEqHFZbPvzks1Bf+M97XGK3NnSf77Njr0aCZ+OMD9xlIu/H4/hvNoVkXZ1iqwAjMBI/Eu
OS5YrAuWz1iX6KBq4KVU8iIqzKtKWAUefOu4S7vNKUYn4aKw/0yyWBnkTdjkhi5GKr6qlBgue5y/
6ulGOXvs0VEg2+DnKxkf3IIkOWgSm9ROB781XxZ8qUws3tKmwihwLdxSVN5TeAHh6YA82MJw9jgs
8NgG/07Jplg+PrM+ejwpKsbjSR0+qNkspsdA4AAfwMvBZSmZE9WoVgzRaCeoHZm+pxx68zxI43vP
1URwTWcu4PFZnAndq/suvNxMH9e0+stQo3m9HxPtbJ0CYmagj5fu4v0kzQ77g6RLxwgnoEhxp4VB
wY8wSxcnUhy3TMtF0PPhLx0F/lehTMLz0E7ldTAxjMQY4arrcWzUhrLylOp6NjqRv5H72m8cBvcD
DFd6F6AH40Auavl2nTShd8IEReqjUohWC4F2TAEfywIGn4gDGbGVftcIshuQ+aafS5Qz9Y8JoEGa
iNvdJ0QCw82pVte0QFKb5py3F7iCc5Cv8EN+blEcwzcPS3HA4UaKA2qoeGKlWHWvztGZbhUiz5Uy
1fvt+3Xb5HPxrdRdmJtntd1zp1xJAczEow0dnDO+EdKov5f4OGUyBymiFhKyB5o9eNiWbRGoKCAZ
H+SNFyE4OZJCCV2ERpgS7095hezikXmCFYe2c0LR+TBG6tMOlpXaYr/2WdacNajOfekGaCZct+6i
2v25AKasbd7xq528n4K4NK+886Hg8iTaazkaHNq81sVsFd+7WdoMvSo2+7GPU4a4eXLJbqQBxMmu
Ahan9dd5yUS6YerEVjYN8JfBp5hYbKH2Q+SvfSjB7S3Xai4yTqzmIdnuNMflFQkWGEtTCuv00x4Z
OQC+DJPqbwllqi9fTYpJVSjwrFoiqd84pKTQvvnbTaEn03P7eYzls5g8SnIAP7uKDl2rT5XGF36n
QruXQiGzsnHp4rmaP0ET8fE3KW3VfQS+1DhtUeFz4i8h9BSJdvpIdgASJnd4UwPBvBD9efj21rps
lfrYEw6ZVkHwsfLK9o+P7S57EOzDSQ+gj/2royeRFzLOABHhI0tgwSZust0c218Trnn7+S2I26at
VLMs8OPTUrbn8GDo8lQT9VuRoXy10NNvD6/SLO3PWeveHntMJdZ7wbqHr1et+W4ifMhKprdZL2dJ
nhNIjPNHqgBOw0HYy67sovb4p7N8jfjH2kkj0Lqo8t3zb1e8eQYoD9BpbhNmy0FAUWQG9uXRqWdb
pqmvChvmxqg2hxxecqT/n4hcfbywOCpiom3+3wFo/GaDTKISodiyb7tfFYOKQ2Rel990g7Dp9H78
fIEd1SYkeymeVnaaLSD6q706rCY3bLhoYuRC8ula9q++J3068VVO1bi3OhDta4R/4NeW8oBVU8ds
Pnk/ncKARz0zDhYFHnYc9SlPhrfbCWVkC1PTWefCjWSGzrK/K+RT4p4PJc8Q//f4UCjLiz1LSBVm
ald0DHZCJEq3yqgrbWTiuBQXjR8ZCQwCazgi2GdteKkVITDFujKeLJcmhQ/0WhpifrWIvMJpiQ4E
bzd9S6I141ZJiutlVyIQICfUOtB+aeNIp29YNyn/xg8qXtzFPgNv43OYXJQFI5cJeXrKzbqlF3Xy
MBYNHvKvIRqkp3hpaaykDf/URVUqrxItkcqNIruRmVjHeGIeAwnVIbARpr9ND2KurDt1fog91bEj
/WSJb5hTfWzMXp+qV7FlgiXfOMTMn2n4F+c+jXeXK2UmsWb3xAmEjHF2W3mpBm4fh3eqLfKSmu/q
CTwy1Rh8xSUBMGsMQf35G5wABpL2WBf8XeGYoFVRP71doLuUdOnciZT4CTXexxNelKMVxFVmxdh8
9oi+vsjuYQH5Q1zailemLT1mzgEpyb2TaX99Xqk2SQbq7CANOk8UpSXhQJb8S6e7D8EK9Bpt+FLa
p9SVuOKztALsO6iTPc5HpUpn7rOMla0R0Sx8qJsPy++r+VnTHjXekJxcuFM/V4cdAYvCVsl+JN6q
q83ePlPSQq15iSRI56vbDBWW0LCWo1v3b0uZ9rmilfluQ2GNtxd++p6C/Pwdqhu+7Ipz3AL2RX+c
Yn7gaUZ9zQcjQXgA+EzN38MCM3/Zw2KCYjogGqYV+qUcLNfaZhV6AuwnxLgXNQbnTQhAvoB3T09X
j4fugrx+C9zpnr3wTLDYuc55y/9Zm8z9YEBmpE4Thxc6RbllCG+GWg7COOaWJdQvl366F+cQ8uvA
PUL4GlRa9tuRWW1kA/B2k868Nxzn2zJRqOa4P+8zEBGCtViwjJqmmIBT4xlJpJ1cPS4B7NCbmxEE
zJ0TQyEl4qOUGLCSRNIwJl8Wdmo1cl27yqPYNGWe2LEblqItlyLFRqObnOh9KxLn1B28l+xCD1jc
rrScpnKhdrIf/u8Gd9Aa0GR4Tjhppoa6ZOdgdda1YDIjSYsgFiJ8nZB44NXsEa/Gns5IMdFdsq0e
eYZZgYSNsKPakidFQ4UXjkauwNAOaGDLnoXs+akI1iQw6GZ44MjjglMJ8kFUUpz1dArdWELza+Fe
ZZIIKx1jASEp3jICLZWlu5xj5y8CrFsXpOuJZHW2h6z4jGkHDhq9wJ9ce4a01rOfJU6zGb7jXmTL
qwwI0KLFh1DHTd9uDO7vZpORq+aYrpsQFw9Jj3IsZAOoSJN7AlwG6AFkicw2D4pnQn8iZ7a7+j7E
7/kyj4ZFB9VUTWgtfX6sTgAkb/8PYIHtxZPnnbbGm76TcOKuOWkte7z/4HqpLQMPkd7qx2Q+VtR+
pMOovRwzESgUukjMOC+YLXydz1/9OTx7fSfVnujabIh1xKK78Ih2csskYhqO+bAJxOIWl+2hGCwe
Jx/9CGzATuH6Sk0r7fxtDuYXgdvtHzNvzznLHbS42Qn63sI9p1pObe5nD8/6vKr3eYyLCjBMjpVf
ke24Pgi6dPvA215uciZB7sNLjLKVkcYTH0xgwPcm9WX+vfhSt2KvpOy1H8GmfwCnBcNMgiNHbit0
IXPKMzxYQhOQRepHjxdk4/48GihL/p7wxm9WSR6Leq6XGG/ljVJoJW+lXOizjmOKLo6QmrWaDWPR
rWnTwA2b++g+XKgbuOcrgh3hyPTffNkUvW5PiX8IAXuTMfEZr/8bMWMTLm9XPyj5Ry5TbxehBtM9
ePlAdSNJkW+1/y+x0YEPl02kEotLgPbWrKl2fOOFW4fcOX6IgIp8O3h4bpFxGDm/ww0aaCRp0tds
cAst3a2Gh3N/hmykqO6/y89UrUxqQnJYpsvVX6UCoo67c1ih2f0LmlSgrunUkaQmJttdTaLYb3iv
B7ATeT4+GkhVsfyobw+4Fhcu+SCpQLphDN1Q2Obmzw+KeT5Q1zEYzAi7eXfzenyV8djSbc29dH4M
fxO995w2k9+vTGW8/5ks+M8/Rb+2U6kzhFuJOhslir3HW8OJmmXYVGDEdmjcKq43xI1HgQr6+23s
Gxy4B0XrevO6/b9/4k1RTSW63TFJi9vw4tZ6K8cjtRtkFL0F5BRaoBNuwIJRJdGeVFwEHQ1p5Rbk
XHZtERJo+EorAXyKJpnkTOPxr7TztMyxSae8uVKVQ0dfNm03URSYNbXPuRNQAuIqOsDJDMDVPTNN
AEQZVYd49KEiQ5uauNBa8auFek3zV/GYJCS0DhAqiqGjuaIb+hRJOPiu9mnswN9c2/ERKdacjuYS
0FcIOn3+s3tlL2dGd+bKdtxaF0tF0/zBTuhczh4mXeq4F3uTDdgcQZKocN7hBB0ciyRp4Dp4mk/K
1BggMEQQkgv0pUuZNoYm1zIE3oqHvheluyOkwlIG2jb253Unq3UVuYhjIpijtrRPZ+q6igyNYY5a
c3y5YYJ1UoCJ6ZDIhNbLrCfGuFNPn68ErIhMYydZ4Re03yYFEppwHrraL8Yo+vjEVj6OyzqXK2yN
VsqRtZczSSs1WMitj5hBHweFaOIaBduu2SyX8xEX0K+P8DqpSen7Bm5vfRcowMEX7wsplfWrd35i
f/h0tFmoyUfPyAMZnGIYSBLH0jJdoHZe5HIsmL5KHdTYOdNeI1RQein5UYSn364UJZiJfIQUDS4S
KKWeH0txU/OYkqqerrd6lS8iZMKUp2ErCKZeG5nDm3qXEnOXKiT0a+k24ltvNxu3DpADBZ7ZKbeh
Ib04M+aiZyS0mwWL2Rs0KTI8GEe6XGfx3Kmy+dCEhp6JaIDm+syS1+cl3WmXPyTcTWwrGsPAYhid
o9zFzYOOlznvRGaLm6g31ALKX370YJRaxL/3fi0XTgHE1n3bE9FJg1qA1mcT0KNtikddGiDCmhpQ
FAWIWLLOQLCUPdFtdRNmxTSh2J35DE1hHGeguXMv/dlJWVrLx0tEebvpa9pAHRSQNs4snoDej6iP
glAI2NHiee4YVc9CS+KMSaoUBkwEkKAa1IS5khW2CsFSKUYwURvHVSJqM4dbtjnZISdcUbCLxjcf
TWuGaBg/yODBHV2dX7TtF9P8mNmBVKDu6m8jKmcpdi3J7v/U80IyYrLQtg6KgaK1f3EEZR4Je26p
6DKm/pz7o2HM3geEY13MSgaW14gcvS8JR0sQeQr3goSl00GO3ToIgkV4pI77ZmMRgl4lBavcq+Mf
U+Y49GGOv8U0mfa11h9LXWXyHgnB/cvBMwciREmr4faB6qz2NMzJsiuvcaFkPWNWXM64JeIUW/6l
fe/md4bf8kV3YfcJQbGILzzfPO0nJZivDkHUokV4wI26odwSJA3za1uF9CI3MQT8zDNyg1hUpbEM
k4ZhPfNGsWBIt/h2ZlIp+WocRc4meLpSPCHJlh6KRvdjxUrqKmoPLWy64a728ucJXWqYkvIR5Jeb
cfrQc8G6oC45emUbLBSVkNcspn5HaJCTJc/Ojq8ClJ2sI/avAOHvycQGoQ8IS01HxJGuAZPGVLje
ICLbCn/Nqn/hBTjeBtcPtyCTopgIx/KoajrOZ0x1ezYIKLouzhn7b4uczCKQ/gu5cR7HjCEWHLBg
+Djqhl7R1H9COIybfhmHuebD6/P6lAdkc3Stj/w/R/2YRWiQ2dLy2wBo4L8LByYiW0e/HOx77OkE
2sVJ6p/uq/ZNcRa8NHIFTBSYNMx4a2xNq0gqSEJNmVx+UM2AhVF4ANEmAjQ2FQ8i8Ux5vAbMU829
XlrwsM0kE1gbidrzQGc8cSdBqR8zIyyf+IEgJ5izK2sZ+cKJAYM1OO4rEHWn9iwl6PhRqpWz3I0T
hjM5Wa8ue08KwlOUoPZCvdaMQoVybezV/kc1pt+Fg3GwaDuKrW22DE3YcupWXwmIaOf71BzVUcCj
s8wsePeChoNxzo2m8ik6WhrD4zPVgzZuL8XN2pk2Jw67SCCkCuCvEX7AkMUCMrDjHWctxthaiz66
k/oc4W9Q6hQKUcPHznQNXrMjj6VVVnrmdUbCtvWtmNo9r0m2W9lJ4eKojYvmhJywFgpGXtS3pOyl
5bSpiyHDCzbux5A+HhbQWQnWtQjhQaRBzEIgZiIKXn49TmJIil8O5k9vMRI03tuT25TbS2ZtGa+A
ofAFdFAjkU1/HAG18yKx2WqsrKS2DIPQ64vOvLkbnUvES4rMkVsYbcFtl9PUNd0895me/h9qlYJH
vOODqxKwobPrY+Ip8dWP6QG4WU6ezcPF2YVM7oZikvB94KfSp1L4P1jQ5Yqgu4Lk6SDPRmKywQIk
7UgbvZSB9i2jCmlbxdMknqxxHFy4lDyo8u2ZeBFGlgmR7vSoLi+wDazjXpjPrtbq7Phx5FQyXXVO
rgYuDiNB4DWED75C5+Fkn2KA47zyNROTz/W3ful3pHHfUNwdEghaEvd1/qt8/fFJFCmZ2wb0N+5s
/cwxz9qe/6yKeJScO3ipKgcLwYz+e3UWC3R7l3Dw9AKgoemjIjbse2ZjbA5274Byjz9pvnqKZxpj
bHm4IAXDD085UyCMiMYaN8YqUEDOxB/XdWPqjwoqdg2ISyza5r3o5BakRYZZ9OiebZPX8ZZKupD/
uBqRSGXXkbciUPQrgN/a73G1TD58WfSM9FzhurMZS/8/C6eQzqsEj/i+C6UTF/Qlc/e5RNTnEdME
1SyQ3t/SUqPIb3VrmQ9/zW80r/hr7GLfrvPYniI0NBUm9X8E5ECQfZkGdY18FotNJvr882fpPNis
8a9iVpwpzBKntnb4HgO1H6U4ndntzr/N+2G6C5sOctoRcclAACSpdGQ/nkN3EDHg3gYm6t6+GxXa
X2EszRbQ7FDjJ4sgNkoutNN3hLaZfuEsXb81d0C1ykoUOcdu/1LVTqo7jogcFEqATeeQ/BTXQABB
8CpkQX1n4u6sjer9cw7gQy2sI4d/OlCLa4BsagEwDHAakEwovzE6WYEk+u2lszS/whrxr2fSGzgN
+LVr0jJnkgHMbn4pb7tQ6xE+b+Uj0rcszTa4h+pHsaK1wR60feQ8nXKOjzFpEqTOp3NwglPmde8O
Isi/ADcE5VhLTjh1RXRke8eMTIWjCHk6i8tgwAyJkIof3De4PxR3WWGPQkA4tYUSitS9kYjbqmIU
G1GlOvgs8ig9nqjBTmqihqLAoltfkMjDgxCjbLr2heQBt3JcQkmNHzbU+ZhussAPH5YQYoO8RRY6
aF4iQaUwsIf9fKUUdD+RVZsLTcJTd6Bcer78ObZgvmKBPmTijtTTRCJAIw5Atl+S1+7OlhFMG+d+
dt6xtUZ/OkH/Aj7Mg2OARP/PKVG8dAeSH8V0hzuZW3fGr/neMvbsJqH5Zi2inPorucTxiZdgAv2c
CSLHST22XzycUKe7Fhhd5ZY/gS6ysRDPEkFG23Stwp/NCMJMDAuxBC0TzWx2d8J3OP9dJHSnXtue
PdTf/3z/v7MZ9vpzM4KIQzGrmrAW+EZOHyqAQ6hw5VoYzk+I/7jyrvAWy1bToi8J9055uLcLCn5D
OiJQinSDQ5lxIrpZTITYDKwV9/aSgfcPWsv22blLOw6gJuWOVUbxRD/Ub22+rnp780mey2sJq9um
1W2HpjgCFuRABHi+cNKG9iUldvWfHKjZT2hlTg0U4kTrFv7fUVv5buq4cxDPROWuTq4Dksc6R2d1
YvHFUtEJQ7yBAWeuEZwvGrzLeq7PRW05fY/O8Z2jh/A7VMCJdhPvZYO8fFYsirj0Xh9Rbw7oqmmu
c3Qnqljpbk/Kj//no2+X0rk8A/4D1UtWJ3XzHlB5pkIHDkgq9me9Vm7MTxaGK73W5HKJFGfW/Pvr
DTfVnsUb8KkNAOUTFKvYS283TQ3kgXowKESHC6/u7RSDZQA5VyQKGFsC8fWTxbYBfBGiD8N4xphf
dhD0clRgBMcC/Kzkq4wtKK2NZaVFO3HisCGSvh8Hnyp/CsVMTXh4bYId67nTg1tem1GBl3uQ7I7N
vOh2brmtXHEDXFixqy2AfpAmOQ9QQJKdEoHBd9P81PXQmbcwL8OTrM/Ox63E0lAF47GL1UlMMHby
cZjNR6ltwOQQYKXuqxiNRDwGmvJDzCxoOIRc4FnF9SxTRWKLWimW3GrT5zDmDvta3UJRk9uIchHE
D8W7LlIwYJ3D0LQAnlWHyo24N5mQ+Uw7jvPQov4F5pHDaUgeYGqKgFsEQrDz7PbNMcQ6f2/GMwbs
Sg+48z8hnVqMBBrBAqNJBC/U0QGGsA9L0sGIKC0ZTjrmBGQXL7Zxz1sSExjKY4tuqmB7/E5723cZ
TTzD9R8BAribO9y4dUwZgolEQFk0RPCCMjmD/sL215sZCbgmEEm4t7o7670Pjla4RAHYReCZ9CJq
rmtG0wP4xX0PeyJ6rk0aJVoUGRG/PLxiPAquhuCEeONXXSBimkkzUlkEPfwgSTJRgp6pHA5nQ1sJ
2urJ/u77pZc1GezmLaqka0Mwhf53/Asb573m2l7kBQwIZFzoeKga9wHW1DTQxm4JyxkQWFCzVZ68
cP+n36dEKbpcacf5MVb8jY7k3TafrnuHNAyeaHdFPo7t6riI2zmvbO6H6xt/H89bamWtoeHRhP+0
W7zvFqCVfD6M7hkJJ8GtkF8L3uGIY8mH6SlDLl7EyFX6NmUMBOycOFoTKO4WEsrxHZ+e6Lcnrzg3
NZiU9FiaTGvvj1a6ITxL8Mc+geD97AGLnIM16wTpzkz4wOJjn89CIop78wQm1l4oQ9vpdRGMWCHC
/EHOcQdOyT2ZdUnDf5ZSK0bfUwzXt0eBp6Oad/MY8jq/+6a5IkPUHEUggiDCWOS2pLVZRYMfEBqg
v+uZkyNodww62qzMzZBr8Uovq1Lz7rIP+5WWiNjtYEwEkiA3N/dfZpq0WPBV5jnOS1nYeZ8XTouM
xs2J/XDWKDJNrkQ9oPqOqCe+sCnDWEF/2S/LYkpUDUy6IOldR0UoESR25lEfiukMEg5U+2PmDL3r
bgKHmYhToQsBlVROSlgDCWuPCuqlVbokEMqkwxURElTg3JX50IF9NjBOJ/idihOlx1IlUgjvEmUV
QwO7XOIEuHPi5bpDauBUQLkF+rxfrQDokt6d+Wegyu2ulvkm+NQcZ2CYV/KGaPJteYNTMhRRCnZB
7rPMJbPKAHuuxOaWWr3lKIoRUH7CuKpK0Uiian24xHtTdJMnt5ALPqNLldy6s6HSN90AHI7ToQrN
3QdUTA9cewZNGDSKyGhJlDuLgo9d2PIIDoXy6HPWlv5s5frw1Rxw3wU98OHNfuZHOLxNh6JwxICd
UYCkvBPGXRrSuwSSKW0DT36aWekNKIVSMHLyQLDzcFJTtGTorBC62IqLSch4btN1+Oewm/KDe7ES
O9OjwM9uN6vshP/tdoJLb5VIuGfmtxQ0a2vV4w0qQ5lSRY32UBjE2tnz5ZfbwZJRZWabuR1fJdcM
80/ItwOj+9WUT0epthu0Uzuse3luhwUWQCMcdxX3W7AMwsIieOc/9Wj7TKP6npKOPOc3X2kiXKVS
r5xrMqxJSPWbzD2AkI7FGv4rMvA/hrJS8rYwSQ3hQlsgYKYywWeTGs/gX4gmpIawJ3NaKyabMW5L
FKmhMAxguPBP5xDf2h2kw+iR1etRxxv2hQN+I/ykZlEtEcPLGKJ8+4A0T7FrwiCfJAzGF3U5Cir6
hQd/PwrvATQR5Y7Y6mr3MFAP2xML8z72P4g6vF7x/BugvS80vV0wHLWdxbFPG9BFy3bynJQjPc4K
nASkCD7dy07VsemRhXxIslfATgdywTEWRAH4Ia223h3qiZ9jMCY/F6ZX/x/K3R2bFA/WsuiJEnOH
v08DKEiaA/VOBNWtHgE35HcNyhrZm8c6BOJmmYu1JTHmPcmDQfTl66TZfc40mlb+5M0YzNjcOyd7
Bj6+OnrtDxLbYhVrfL7drCYVUaEPMJG65gNPJXg4fla2v1N+jdSC2Snydb7in8XPwCYffRnoJsNr
YvEGw8oCmVY4a6U3CYrCW1tyDQC3MznWP0ZPHyrfn7LhJMwHjTrbtJNhatpaq/ewzdmj0IRx6m6M
EbzqExDHGCv1yrutitEBvLqC5Tam9QpKguhhPMEAvqRJ4qZV8AA4vqDNzI3JsJAd972O9EPriRqn
oTQ4GshpGUayERmUxBiAn4GtkMnEN/b+etkSKr1azSP8VW5gx/R0Xk0JDdYZUM2s08c2Ae7P8D/G
g9QDPdG1wNwmqczwTLBiR8MlvY2O6+zSC4AKaBH71rkD67RyWHzAmKxXApfLyDeJNe+miq0Z64ju
uLJaYFgqyCXBq6smphGVmAbyX6+XIpofLIh6FnlLaoH6LHQevdAweACFR8bWro2DRYA8sexWdqO5
EBpZXvSB62QYW4kMIzOcN07k8TBqadSshpfe+tiH1w55OvAzqW7cKq/Da8LoCTRIl/DAZLaQpop3
ezr4C5o0I5XvnVjOTHtZ4gZlKEizdQX/5nvIxOmsH5hvrtRqlqhrCLUGPWN2TFArIrG8Xt78Cgva
7MYyVL3Rnr0cTgHbd2mgaXxZlxky5rAmgWWgjaJfD6NvhYXdRVCoBxI959zCiPd9mMIfQpo0Eptq
3vqiJcDwIVJUzEfyL5BSRKMuXMQCjVsMnWTEcC9QC4V6xk1qzMOD5JtostsToh+KPyjG5WCQPb6v
w/B6QNicsDuHqurWn/dOAEEl6BTZrs5EvLAHopOsyN1HbVw4ZBqQ3ZOp3CFtAdD6rJA+eFs5rdi3
ZjqW9asLTnW/CUSqk0njdWnJ+ygpTu0/JeojuxjH+mqvA88IzJKjviCM5RaompOFh4aLcj2dPZvn
OwupqtLXs9zmJYajpBa3rW8lCbxk9TJqy/s36LADP6glLwwZVQgLnMBcEDxMO09H+wvUedqQftXJ
RmgnS6f34mWx+gzQ617YNV2T1gczxiwPV4Q2fbZsTD2fdnPcipmMigLmx5GsJQeotfDRXNOWO+qa
Qz8Hf1skzAgv7ecw0ve7ZF4ggkRuT/eeD8UvWqLo4pRSDsV0U0OGWPS8Oc/GG7apiE/zyDMnWeji
asZ+DEEI9RQzD9qAvxIGmHsvn9gQRw9SHdysWPFv+XkygjE4esZGItC5m4FreZ3Fkq2yuNAb++U7
794mltB7TpFHum8uycyofffq8ps7IzVyXm5qopCfKMBKb5mlBLzKw98GdmCOGfrs+E1PqQnJUtzr
mcQyqLx6+OH7cDEscooDoeXzRt2ho1ZeCj/7GP1LBEr+iosreltd6Q9qyS3jsmY2pVWEniXLCjE4
jWKNCPp05MUaRW/fwLocQGhMne7qxRycE5StpToxr408cZBnAlHirj2nImHttbQ4Ezu7WDCtAMb2
IMuJUhqgd6gw1vSk1anUhZkejxEGpl08mOrRHt1L6Xg+d0JOQRDsGZxAb6i/dOjOf/c3hExX5LxN
D9DvvLQmM6NTTY/firDEywAuVayqDc+XdBQ/mqjalngvEH1Vql0TdbPT1iVBoSuaIneGWdI49LfQ
iOrZb6uCmpa+HNE0D7OuwCfHJua4Q0EaKDtKAKAzr9qHeg183edjfZEAplQeQyx/DqTtblisKQlS
V++dwresuNKa9AWZI/e+wMHFrNxPktKoximv2NoUZFmktWOAgCalYM1YPX5HkgGkgn6EdzljCxfv
+kDBhvAeY8qr3HZCdSktmIwA431YGDNaNEAQfSvxWKn36FLP2s2a9dgNp1G6ETdPcUhIcRTN5TOv
arg6eRIeiGjZjwqrdSFK0Eu5LwjEb0Zy75pmfVRuOAyA9AcCQS0rZYkUdEYAn80WbFuCdEjEyIjk
jJA5Hg4SxVHL5IRdFnw16x2GT5x2Xc0PkHi/hiLHWaqspVb4MYNL1VCk3qB8k6dzx1GIYrcqsjq0
aRedDiCgUIOB4N5drZ5rJW3vEjYy2SKnQi02KKsV7isez8lTjC9/JY8tCmW0bw6oQXylZyyOjgO/
SOzxKi4OeuoMv2IwO7eDKS2gxTSA5i4K4PF4jvUN2KOC+PcRKfNsJPZA9KHKouYZOEGprFM9W2Fj
BTJl6r+UxIKdlBlHTZhME4AjcAxJ0KrQdWa+OxrfVk8CskwF6ouqQB/YxObrnPm0UncRL7qRe/7f
FVfeOPXlcvaMYzaGQdM+MRMXaGFpghhf/tRyLtKQ37qpHsR84xAZOu9uMgWwbtIWz4H3EdyHPVQW
qhcpdksJjm/DCtg1aZb7e1qlBJ50ducLAD6/w8m3FXKMSW0YXYaH1HFkBKV6JzXGfq7IpTDOXJNY
mJ5skaCfxLSBtKllFqPILRxJ+I5zRTX5Xq8bF1iQePhZc0pl/08d3t5EkKCRl7R0K2m0cqPjqCX+
xKs4Svxa8oMaddc9IkiUoVS9y7FZr86ZFErqBUyZKRf2MMY/jtfiY3S/HSY8C5MOnNJ17qNR5vvu
Lxz2JhVQhlgvNgkJO0+5gER2J4Jb+UyJ8tn1Gwdi4/IwMrNFrxxWOUxIeSK+PUEtjWqYuruZr5AM
9jqEyGcHOtXKUI740hXkDVxZThz/zIVw6CAurCclENsRYPLhFyYJt6Qr1tnWxBrJ/Z3aS5xAFa7w
gVIRD9YMhG2CKbepDMVhBRJbq9jPnKpkhtvpg8fVTKbzRTCLfnBEQbTF7+PjxeTzuMGKdn+GESwq
VCUYDh0/nFHmNUf6GmuuC9I+M+VBnIiDPsIsJfNo5sN2H11ZoFf47dZktxn60j1Oj6d0/tHLJmoS
TXXPGbodr1rtuPdh31gxL7bls+GbxcQ5/1C53/0ZSJIDXLyFsk+2qFtiQ+Uv6JMflDUBXkYdVIed
YmC/nVGFS0TKy1YK7w2K7Mv0NgU16l0gBNCYv/sUFGJkGvK947IwbR7ywXyjquc+tVVogtognBIi
CStVuTjNX9mf85dlNKzqTv+zladbTB56ASuVqDyeAlf71qyNY91YFw7LPUD/mKv7uLP5z01QC9kd
uYtoBOXqKlSa1CdP2hDaJOL7R4of2Rzls0YFg8uOMYOd0Eu4wE6Py26nQ1vF+mXMwG4zP+ufL1Kf
uMVKSz7lXCHV7YqA/pd+GcW0inX6b99hb+Crh7C1YWO1jsRUoAgi4I1dPJ6iIBh5iB2LMkY2p1YG
ua8ANKqfLbk37y+gx+1Je6ijxWhmBZEBoQKkgzmxVgdtT3pCiutuk9F5gCrqZa42bLdHAyhtNjyB
nT5m1x21t6ijJYMmWe6EK3GyfDtSvFln/QaPcWYCoSURNI181VLeT1zLM7N5oXFFKhEnIymnpOky
DQQ6XOihFRV6IXMr/xD73pxLoea+5xyzawmFelx/JiykO8XvN4VzIDIiSLjTTOacYuwaBeNu4dcY
7hNTs3JCgc5uLvlJ5d+7u0bKFSq0jwmtEdzoS92tu8Ly/hivS0/Yu97G1Nt81J/HY32FDnQLoDNE
r+ov/s5SrN7FworiHjF0JnadiOh6IykPDx3Z8rk59E4Zi0VI654kn1KLW+FvpfMQGtcFkdJ68zlF
mwWDN1hjhL7dsv984meiSRe0LkU+W2uWZu6jWT1ZuBCaK++X1rvZXru7eC0iVViOIm+sCUCb22e8
g1xFfxXWSOLkUbDxOE/EH1WKGlu5qg0D5TTCPPKp3QFnC2z+ZTCkczuXRW4FLuFCtcgJScUJ26o3
TNjf+WxP6gRdDN7tcOMYKTPAF7GuDGchOlODn8/vzJherCe0Is95k6DN6Q8zMVcv5T6b0BtA9vGb
dC+Tr137lFDJaEgzhwBd7Ee8p7n7GdHAePMcoHIXg6Ez3FJrvevOHiISC5VnnIL50QjMIHQsgEU/
e0dCM2q1Ah59EyKQHvw+m569g47E33/9ohbvZYxsOtUigHLVURmoE3D3RCQtJwBN7W2wDz/50DLK
eKWPKcE4kL1ajNESnEcdgjeyPmRChbaekrLhjVdf2OkQ4Z6pENpMxj78u3yZBNIocWYfWanPwqWk
3O5Oy7fxVhU236MBC2AZs1vKSEJKhvK2KyRgZVArepIyrbnhfdqbWKr6rayaD0ddEt8yddbzQOsu
gKLdwY34C2eG+FgoHHzLE/EdZGP4BkLODOp+NU/LxaiImsaXSsBIssg3KxIOmhaQn6PAgznkMt+K
yip8C4+tTudsnlqxUaO/RstsSvWwYEzmflGe6YXux8agHiZXaNoaTp0myIEyh5usJL+XrmBCTEpJ
7Y17vwwAG++vUilioVi+grzp/lDDqDYyc5KwLahQJC3faBWPS/0SsYxfX1e5rxVcHHZkfIsNIOXs
FUCURN721nm1nj6mUp53MHJdSradgPvakEwjyl4fiE6UG80xoy1AMU9vzJN8cJfmgu3VGRZdLtu2
OJKtMIk/8Ic5DG8jnehq4ktb/I4/vnY7zGO56JUccgiO1mOonIbGW727VLa+S4s18tcpjr1EMJeZ
P9uOjBDbv50UlHO6fju/wHCd/ptyK0eNzwsyITUveueq3BShcH3dSfzJvvwyNCiH/4r/243Z1Rf+
uBvBA9PABn1huLlXoTMFEQVSsW37/gpAFDyk94triAhKKyHDHLigTqEQbsKEa7AGK10dRhpH6jrb
vGTaQ7/XyONDnmy/IDwMdUkQZM94NgiERuA3azdM+DfYWgfKQffwQPDannuzTLyiyaYQbHXmUdfS
ssO/Npylyh+GpcR2BvDQkWWpX6mt+a3hMV0m/5yEmJd+HCB959Cejh6+o+WLNM15SAq+OENKNXu0
Z9egT7B6iwi7VLkoDvHWfifVS5p8mpLmHCQVBS0+wWbx3Yu4HS12Yol9hpTkw0sWAeoaHzuXE8vP
4sLraU5BaTQGt55oF5ULCCbL9sG0B+2siFFQMDmvVmZaPb3QoNS/1QwCTBFjdrZvYb6suGLrB7Ob
Quuoj22BXApYvdQnZqcZVxjmaOdsrRPj/D+itGI81FFA4bn6SwcR7JcURd62+dcTi94/LIDEj72f
TsAIayT7a5gz7eZiPyo3XvnILAmLOUXR/js8/Gelt0mlOwX16AUnE9D51jeTMtQQyShoExym0j9f
SOD43uDZpHybVOWBFFVSLB/XH7b+LZyr3eNUViq2/oJkJFb7G85PL3803h0odChwUN6jNw0VORCd
Zwo9tiVrK+jBpTXok2f4+Yg7NVYIzdNV/MxrGTLYtZIAUJrosWmYA7B2MUz90GFL+QIvWjQ2+9M+
4VbSAAPuFgF5gkXxntDgLOLGlDp7SX8f+8FyECD3hcG61npYqAFO7+UdfDw6GJ12nLnX6fh0U4Kq
yNGurenvoccz279kAArjzjVOwj8hWj+mhQkuep3Qfzh5/RZOyywZdPoUzXCN7crC9qD69fE2pY8d
7lDKONiIMuN5xS/7hvRGLQ6XjCP9Qp5Q8ZfA4G/6PwswRwkbuGsUSCRzwHH7vnMc37/bVzC+drL2
Lj0uhR089wP1u8HajoClz+wO3I0coJ8YYZipwsHTWg530QaMNB+lhzkfDGMgvH3r9IEkH+ULmUI1
LkUXcL1+Pw/U4wx5lQEu33sExqFqvPSDTxGlU6s3IvbQrqmB1HuQg6dO0MK9sUsKrwQ9PxEHV4tS
k9HxHy2euNalEpASFmSUxJJ5xPdfEE/nn8Z3UfZ3c14bDil9MY8Bo4EbkvpktfYdlUjhMzTGwfMW
CiDZBGMK4wS/3yklbXmAUZP30WjMSdABTaiWdcYBwAkZN5bYLjqk5VQNsie82vzqtWKu80skI1Q7
ZyOoP9+urxCHWhh4Dfxyplbk/gET9LzGJESN4mHxm1Z7fCEanf5vtcfJN4X9Mw+E8tR6B37Eb/Hz
ccGN/1G4va8gC0eqbin8A1IePLsEIdUMxOl09lIJdYac2SASsAwrLaTtZ0W/IqBDSogiaiq+8RIx
pcCeqy20ICXUgx/BJfZ6xZSVSUUMGM5TkOO+lqsSjGBXMyVPNpH4Mwk1Nm5VoPcxqzlYTY8ns1KJ
0UvvdmtLvDWO+PO+oyjgUmOV7ikHQfgZuEqKPXNUy6mLImPSmlFRADOfO5yLt+swV8U0xGo5fzjK
t2optsUzpQ8jtFGW/tZE0zjxXnLm4fj4VYI7idtZS364+V5hC3Z8YOfnZWigHyyk43wAuEZBLvpt
BJb83XzG3uXRV/0sUOimbdLy+2E8ryI8oLclUo3vLIYWpGR6eW6sn7T8x3JqPjosBHNqJaJSfqaE
RtIopJwJ31+O1HsIodSLGZXhC2ykRsivauWG6PhAxyiMyzllJdLoBACMnrpOJXB8rKj8osab+IJd
dyGwvMTcFgSwU5LhwmWpoqZwsC8gcBNNZUYPcv3vp/vfJw5c0f3569+qCVAohYlcmieJ0toaxf2k
2BAoCO4zvqsfh0ngJrCClRN9mXmrkRynB28jnbg1u4h86gWiSUMn556nP6YCJ9z+esekk9eQEHr+
904NRJEwrWSt7Qhby8OD1vfpXs2Qxab9bXGTJPqwnQ7wQOwf2+Sgrogq03PuYYgb9GAMz0GjK1NF
cXYpBjPhMIblm0InocKH4efFBW/1aJY4gagV3P4eL8sRS610AyKFZ6kx4CNmXskZSgxhlo66kcAe
hN5DoPZypuBw1WXwLUOatJ5iJVoEdTy5gHyFoO5UMeSR3UW2SFsfqQLNuiWBsL+UFSXCa3WqSDDZ
llUpCkHRiAix2/nINipoyW+QG0vCntAvpmWzukb4dkxVXm9EaZvzJgbR/401eJwCaK5Gl4Jvcltn
PeDDBcOfXpm/HQeeWDELhRzFJSXt8XdjimY00NaLnX3PBZN0gzqZtzecQfF2ioNivpUFxZ2Mzdnp
VcB10ty2hh8FUlKg7sWIWKgQK6rcv2wgU2ky6xZDquVWbXky5nAuRtslS73ylzM0bDXFkSwwqIt9
Z2kcleV7H8ZpaNbfxBsKWqClIkSP0Y7zwFtXy8xYca885hU7X/WV5qXmdHOStBEMX+uJsdcoISbO
Jj4zXNWKTfVtF79MBqSwJRvwM4wYa1RxR7qdLG2WPgfVrlZ8Cw0sAK3THzJjtJzCe8XZjRlKKVCd
wLq2lVbCn2RIkJOu8URNqOLHMLxLgLAZXGj0X+zE7L1KzcAj2mFyDdxnHcvciy2JESSi7CNtVSR9
72IFh6RdBRaYc1SareN0KkTwUDrPMkii1LVqC/y9I1eeYDqyxcvB/5gmOJ6ufu2es7z6xq+Bt7OV
1aMl9mpm0PDpKJWBQ1Gh6T+wks2v50qStuEst+96u/s6oSZd9teKu9AsQf1mqFBQjyN5UN1TI8xv
3SUVpUGpBSW+UF6AmeYP4parDG2dOpf85t+EJoUq5gJluqAGIAAtobzFRV1z2C5wbceFTqxZ7NdE
gTC5sasmT5JDiaa9Ogu8Lak43ci0VnL/PZFYYMG71O9WsLyHtCPRni2PWbrp+fxGsBALJuLi2wHp
zdWlJPiPNFqIZUitLnlQg60BlZnQfjFUETKrTc1uYtFfoVPxxkYTaOTy9Iovg+pgsvCckrIba57z
6CWcK51hUDhpGJ/Uxmb0kKRMxR5rflrsYbjs4Fh1Bjjws6OVz7TNHj8gYVxKWYNdjn/DDk1IDm+k
JGalDcx332ebWXnT7qMy64sn8hL1dCIFXPbdl8O5rgTdyHUomIpnKDvXF+Ydm3We66IQ2bqMoUj/
6z5b/We7xoT8l2YxFC6maP4TS8sa02zg1uTih/3Jzz9C7S4j68T9g4VTKldeD68sFoyDOkfDKcgd
yd+i1IrRt+OHUpQDQ23mRjohxx1Oc2Dc6SFvcTxBwYnlvQuRcfk9zttEZyNa59b3a9x/UyZR7TvU
WvPQ1RC1Axf8F4gbx5b5BKxN17v8ELB2uAL0zHdycPJApwFejjErWBECsb6fBmgb0tH6BzpikF/I
njP/DiMrygZKJbRgKOtGUlIZmTw9cldeGg2PJmrwZ864HbKnbV2SL57aQcnX9ow1N2bc6caeYiIv
zsRlH65Qh+zApPHvFGE3YTk/JVmpszF+wfE74SEqyDoejEDVf8a+QLnbwnXQbLGnQn/spfvHSUIO
XqJIzAgTHJiFVX8cpwUqcACuUztgbtH7Vxh6Q4IQc3oAfI8keLC8BNxO331SpVY7rEONprk1dwkj
Gd+Whmd/YHCOAoqImHVtoCuaEgjWIDuF5DsJ2OxPuERwAfusSW+O8+FjT52IuF0WLk/FCzKzSDqh
dUYw/l2IyHioyasSSyd77S86bo+xOazrRVwA0ak3XSiGRgSwI3doXBCP8EnnAtFTHzG/7K5XvtaA
BV3vI8JHgzJSbUEIJK39LQTSY2DwH5mXNFInRkTGQiIWNLTMjaibLNwP9+61Gi3zyDI6Q3TcqQ2J
SY86hM+k6zTyU2fKZnMu44FDItHSePKvVVkfZ+lEzv8sdMZueRrCQky9x3jlgnxr1WtEPH4nmJ3P
GmPyH3ZyefcsZ5m8/zasvs9BMHR5IUPBqnlrRGudMxSwcgjyjWMCYJifa/SLOFyfN3Zay78oLKoW
P/iZIfmePF2C0lMVGI64FaA3uLIfSwb4RGZKnn1spfNwyEodklGyyy2WtH5CF/eBKyh2/3u2/q+d
oeVImacn6xFOFGW6Ee1wWwgwVJz+f69P4YnAODBfidEUp/N0pU+Mm89kNRaetvOEih0A09aq4dKE
imHZavcXOYBMSVHrW0ogID6l1EnFU1oo1SGdx7rQuuqdvlGZjdFFNjFo4P+V9WmFSrad9YtympZR
svGDsO2jeRbhc8yTY63/e2riXLNi4YdXBtiNPM3WJb5PBtP/643e6lZx7xey60DqEykkUbOivmKf
2EaBz9yc7Q+OtOmv2gSMJL5JE6zhJKX9QjKVr9hG1GibaVRTAk6po88PhtENunMmhScF9mh33FSa
lJpSOn4Tva/GyTmgq1L8kzIh9hW7Ali94g7ZmpU6mK5DPxL/hLsxO1dbtuolBG56h7zNpVTCNNU9
9PUzjXj8NlCFNK/t1cw45jpGnlJdEbwas6dPlq5k4ljLjtESfaqYdJT6SNu6yNimtDiUUFfwXcWl
Y+hzmQ537tx1lOFm4eI2noR1bdNtdGqK/54E9FLAmhox9Na4G3F6rvrIzCnljDEcjB5l6FrMkuPQ
OZTh3T0hiowJh/N8IRjDP86vX5K6JQtIE9VWbuymNXp3dxe8eyuAusX8yMhxk0kOKgy6O9WHT9aZ
ju3/ozppNLqkYUmSVDJALQ68+M+2+tCDHmefxHvFXYN9Kr5fvS4UUg8pA039rzSS0mZq0NMTe1/e
gzIQkc9F8Sp79FnRJuLLlRG7g3Adk6LIGHLjwL4nnpNIPGx6oPhCez7B5MKGSMqNABjgX1D1uy7f
tU3iPgoaUwsSoPB1maDgNZK6hxdLgpyKJMa+BRnz1WZQxVJZuzDbiiYXbLZJvFNN3sKFTz/fUCSv
jftOWxJNBGYzDlYlhNKOlYytovz4hOLfIczC0n4HA32Co0R8XYw14JCXmGHnAkoey5uzk1ukeX3G
fUxEhQFtS0b8JGPo8/F60lIx7eGKTTazTvyf3fE5/bhVoa5jetdyfI+IYr/NKtyh4rERt/1acfmu
BGgE7ptWzjnKwgO4z1lMaa/qlvWXzvtbIt7r/bxgmoaaWFeYHpwjb9jtbG3soWjWCv/6JzonMRl3
lb0wUj1jSv9R8JBC6NS11jsu2PhPWhHUmk/jGSQ5vITiFnZElEDBpoiAt+gq/zWmZxZMvUXnUhfs
J4beT3F3zkN0GZm8SaTQKKzZK2cne76WE3vJ+bxNYMiZZAG4+wjAZCnrDfsDdYhCtTHcbFeEQq3G
XGrfNtLp0PNeGpOAgws1tYkDH8tqeS5xzk+GQRv+yIQ9MurCHSdk/f+gbDeMYe1+CtcYPLi0CBF2
uZ5aoVvLUlA+T1L/O6Q7lGndoyXOIzNWS/f4/fiDlDEueKhQL2U4YU04qQWP7GP43D8HVz4sGmnr
u+jBwkfQWn8OeddKmhAK3bz/lvjqav4B6NgCqNzat0tlgyk+R6agK/GnoXfOwaddHabWQnvstjXR
UkML3eeZy+yfi+Xq31DBPe2UfyP9SMrLcM5FX111KD0YGGNwgKQ6wF4PTsF1FAfO/fM/FHG3xHD3
xLBwNdpyuBCSsCAG1su/uIVGVOpgNh5XoowBt5zr4gN0FDBWdHtmbm7eUW9KO94EMcqbB08okPON
Sb3T9DyKdTzSeGS1CPjX+2aScBo4NYLQjUOxwYKc9V024fxc32189WTHo8ROcvqbhI9trFSbDGK0
osbmV9pVLx5XuE40huF/dayghYuxpUF5uixJu5Yo5oPv+lHhaACztWYjZIRDJ1G4+gdT/45oYdnp
FTcfCeQPtYRNNlMKowKtkqkoLzvRfkoyekZvrzkCsGo7IezLnnUUSle/wdhYC7LV8jiXz4eq18Ve
/Sv+JT9wgmwrkXKa0mMlrgxbj5L5wosaOkxtaRsy6yV/hderIqiB+ZXG46THkpb0omnn4FKTf59L
iC/ReFmPwZ5lZQmDh0ePLoDoYz0n04eFVtZN+7WsVoc2A6DJfTMMQMR28uGOz6k/SY+IQbXDtz0a
Xuox9KboeMAM8a2ZI2rXT5CMVcRZkieeQDpfgbwaWIm34yKwyN5eXV4LD2N9D1jbOMZAO1M+5In1
H0vnMvdd98VK9TYDV+wa2giZnYi84pi+lL5pQ5q+Y1Fbh8ASasYcOClSA5WrfP5bFybz33mdJFug
2W77Cxp+VbJAnI7fUQ+/nXMGELJ2vUmaOGqqm3JhuRq3heoZ2IfGTKDJ9gM/Fd2OnXRg8EHfWb4J
WMHsccqzmkqFQfHU134+HiEbI/nvlV3Gt8SryIhfT4xCUe1B/Wd1KgUZoJ2uWVqtII0eFLXLIEHQ
bShy7X9QyP/D/MX7E7K08zN3vsub8xtaGLLvQs9/LCyminm0oY8gxmwaYBEY3QICQQBa51b9IuU+
SmTb3VMrzHswKki1l/+eyqncbOE1JUxFVhSPJ+Q9S/9/L0qD/Qwp60zH82EMRdUqNaHNMkyTUMvc
pX3XXATiRYMNRkakFfBAg9sjVsVPUxxo39MVNqkzW123WCGzB/reYj/msu+MQpIvTTCl9FmDBOXd
k+He2mZu0P0vcZA5Wg0bY8xg+AJyJkLzYE0bdJynqIjjzFe02cLr4pD/YRK9gsHV7MSyMedUO2Z3
QFfecneSFrQSYN4c/x/v5G0spDZ9DeUR2Vqds/P2mfN2Vqsgzj04F0wyiVT9qAqkHZHKUVboY3eZ
b6Ugeox2d/B7JNGFdeYdnu1kGhFaVV74SwLq65iVP3qWAfF2tab7Se5pSvEhhCq14MlVT4sXJtL4
BqP6A+FZx5xFgEZnyEsUoiIbVdKiovfFewFaZNNEDs/W7b254HnoOdNl6MyvX9nmSkh4MG30n+Jg
j/ZVCaUGp3FaomoO5PfPV1+tlRbdR2YsJddzaY/LqA6XjtMvoUvJ9qWP8qek8IWqYppOemOtcEOe
8eg094dnK6IaFWrN3l0bm9IHkvK5GpYI+SRKWetN1oUDAK6iphb3bplvMQzd6W6vA28WfySyVe+Y
Dq42k/4NndETOUBLqvhvks36lq+4OMrzfsiOFEz8BgLPiYyf/a0QDkns74s1t2EIwJyI13llsrRu
1ee/st/FpUEIDQzdORmM2pgp/LdZYTluDwhzW0dh9itFKLD3zxohs4MbN5NhhO6BVMjPSctQRNxA
HdB9P/S8q43hnEGOQr2IgBY9eY/z6o6ZX7T0HH4TS2mPRiEn6CIvcy91mDXl4DEqHE04pgf0JrNd
dxyirx7NVHBCD3s5rajexAh/U8bjrqaOl5ic+9gkGrQOcnhfoPPp/N+jl470SEzS7VmK5qwUTvQZ
4txI4VE7vK0aZutt6lf2ZxgPUojgUx8qeys6PwB2MgaAJJDRViLWRh052Aam8e56bMOHqmV3ZpBN
PVVCBJXoYtZMHBx8k4nErTqrr437tKCscvWJ73V40LzAc/s5d1KiCSYfQ4R7peV+SYyLMmx1U/VA
7xaBjVso2RnasUJiOwEx+lWE844sJqRwnGEhgCuqNJOjA2IADtjA7NXVUDHZ/XWNI7fqZGb4rqkx
A2iYcGjPQauyHLOJiQo5RzirjFmYFh6e3IWDUr0iyx7bsPX9Ug0rM2iePgaJELneszSudItBMJP0
ZDEc5DmkxYcbLjV532/NRW8JAVPSVzhJSvCifMReE/a/7X8t5sT2H0kBeOGDZyLxVqAR3cBswXZI
hyawVoyF1WZ7DLxvNHavoSoamKVd62m2mJkrn2m0Gv7Wlp+LaQvKpfRsurp1BQFWGuhDJ3bQBXsK
RJ9jwvBDTX0yiZw7tvPB70ULT5eB2iJ7U4JkWG9c3lQkndayiSauBPQrIko693jKYZ5AC1ryt2Ic
MFMgYProu2ymMa5fMRjIK0rBSxX9qGeewWia3pWFPTHqevqDZmGjjlMY81n5Ufc+cn+3+eGux9h7
3bdEHTXjwiMVvC+GkqIfPpsn1+97RPFqvD2UZc3yQ0Jkf6kIEz5gFRjsYnev60x/6zKgYG6tSbvQ
O56dlP6n8vY0VqEAm84E2t0fKeUMLAoPJ4H8aZVLZVN1uoj81i9QDK3Iy6oJqwgo2VUdw6f+JAj0
FYbb8JY2B5Ftnwj/V3a1uL4NkYOTGICzqJpxW2ZFVJk576y6OyuHu6ae+jwrvxwhKbMKfV4Wmi5r
y6lWx5ZQz8fnSMkQrWin1Ib3g6kldnn0NAddERc8ZHIFd7OPrQXNX2RajjR9YlTKSyiZQc5QFtMu
tjmK/O4GbW3GYdbukAwPxoibchtEJieTiwqNap/d14ZJuQFv5NouRNzDDpZvAo5Ma54KgDUGPRz7
2OYPSKAYN01NOhBGe8OEwKR1uknAQJEsb2dJzj1ls85d7PDzys1dNvEGITsCtrrj6BewZZdYmThO
IXxz22s4X9TqvKsw6TMiUMkszOqrWDHy/Tlwcnu/bsEHWcfqeEYR7coUuZQqFEO9+fzJeHl7/Y81
YofeAr8nThf1ofHy5VSdcDS4o7WkNI1epDSx2doMFvai42SMIA4/xHB19GZzLSfstEp4Ol92r+CJ
3qkLecFRtzzwDdXLjCsyYuoWMiYMW7twsZIxbOupl0p9+SEhONNB/5pbBd7mPJuXgzOH52Zdecr5
7bhmA9dFwle90IYkPDxVUzzTY27MFgb9XBeOirXwwLm7ugaJAzaqGs+AXfg+h4iPd6Qoyk8bDDNJ
rCinKFyf3O3YzDx6FaGxqGkjIM5cKIJqJEF1pnWfC9KQilbPeUVlTfN0d2RlGJWtIL6/4o1zsq9P
4Ax5vBh6cXUODVivuEGiyI2bt77AsN/rwKr3wdB379yCY+xOc8aojaKB0hnYJNQPjm4DW3N4LNQL
7eZ0XX0MF08K7x0uCShNI6wYzglQFRm7YIsgVYI5dYR0FYtGeQzGcIbGjtKENcx3np7NoyKIv/l3
0Yc5QD1kaE2jK6oUClJ0ufymiNrzHs53max9vcxh+/yElTCvP01GrLq6hCx+tci9yrQ7IJ0CSZQw
xlFEUW1bAg/dVsxFGC5FtIi+KGMsX1H82gSDcdKnt+qmsdvq0dhixnSX+psiYaTgfzU6bfyjhmEc
ugNUUCBlOXW0JsLerbwKP2E43UNkPA06gM0dmAzbIw2t8M+1iDMRDtnem5Gj0tLcsJvS+Z9JlnMU
uar5eNtvBO7LDMx9JPofc67nDJqeuX4MFiJaMS+FQDfZQApXbze60g5SbmlU8PVEA1rczfiDmSuh
xra3DLbl0SjawMC/LTnN0fyenaO56xdJYhQ6uvFltLCewHmkyNHrOgYM+F36aTgSrdVWtSzp8a4p
vX2zVMhb1K+nhIfVwccONGxiphX9fYV+aePNZ+HIpPnwn8/RZsBG6BkgzlDyQhxbJTIwrRv2awlv
5/o49anjaP+dA7xpTgeODnmZ62uxJ2RNA0wKD0JGOSVFJYE7kZ6kZUAPVA7D/UkNHSN9zaaJWy38
d3Yu1pT2B4EoxdUm2GpwA+M0IKSWKXKL1vOCNXdb2vYu3Mb4fUBzBEAehZk0dUPDTQWeZ0NoOIml
Q0FBsNgDSEA3WrftRkAm09TZZdAtkLi2cerYYXwQnsDiNrf2BZP7ChegDtJwmDGrAp3pUYgjc/cV
oOcwF/j9SXvJ8qUcbDtuenpWgNgfg/f69e+8Tf/VaZknzdWlx/qNa3txZ34rcINtnwrwebBAHWPY
IriZlyCkF6FkBAQNZqyvzQXIg6f2sy9188hIwGDrAMbathd81GHr1BXuN+Ca083OT6npjwkAbsx6
ihfQQYZ0V9HOs9xVIRdSWoy4t1rFQ6d/0i5aZJZSL449VwN5MV3LesgLPOaPvapoLrcMQetGdEV5
h/7EROPvp4kU2EO4OA2QdQTy413NFOJpKEzAbRltJPTsYZY50wB5p9k20v/QQ2woDn+g3IVp7rqR
Qbwrtw4EQ69N70Hwmsa8jOJvruJ/5ZYn32Z8M2sgO+Rq+hX5w6/oRuMQuo3zoXSiwI/3WjiYb3NM
ek3eG7D7G+WIlT4FuUJFC+2tfv2Wq1tofPDgYSeYCXdyi2EYFUs7x7NKEqFLOSXQKVSM2+8hAh47
w5nwx/OlncCQxP2rdrwgugth68TmS69uVoIP8V1igFRrB8zgcfySc3y7Em9y0o4oQchAVBXVVQyc
oa0suNBnbnxSImUdairLX+vpjRy1g+hnZvrlA6zq08jyFAVrHmzJ9siMNEjIfJ8A3OYrK36IdEF9
V5nWdMaGs+okvcIrAz/KBp1jK7Nn2eFB5En0sk2dibK/URARvLAfwZ8VgIiHnNVFPE4fqr7SkHFa
aYps7gkLHVMfCuGH/jFMOxyA4GzVejIXJNhnzzQHMMt8BSr9Qg0leRn8R3xmNnGWAplqg3vHsUf7
YWItgcytqCBh6Rw4mnfRgLfiLnRlOddDUgHu9c6VxonwFgGkx5i+UE5cvrUmrxBc7PA8B/4gRlXk
QHDRaSqxAEzSPI+tcprLWSAJPTL9gu5rQVoon9IWgZFrE5Sbybhyk5MdjH3BCKVRiZ7DqU96qNkD
4cGDgF6pwqce5ZZbICFTmWNSDra2E1JweP4M2I0MoGc1x9h6r0HPtNUAb+R17qpbOFjeQN0BWEGU
5rHxhJeP5bahj32D/TcFmH/MT1MmXAtvM2qOOnYNDhq1/dkUBQznsyWAzTXuAlbyagJt4WZpwJCx
CY+LbzJnJjCCtTB9JW/fh6cavJiXfq54MriPdJMjeDVTNDapSlFW6qJPZP7XV27pVigpHf3sR4zx
6rrmdCOsgpmW6TdqPdI7dwGgNwJwFsSQGV1/hNqSMCfLrBqn/ci5/JL+5X+QunghnCWTdofrw0Ll
epNgsf3pCquhVcHmGAwO/gOnlyJT3CGIuGrMJ95BFZLsg5s+/Wv/x2Y/HycaGYSEXKPxCkZVNT7V
6lYeArM0KOGiyVR2FcPtJ8Lr7/7evJ6fAgbUgakIIHPpm0uM6YKuhml2tyocS9iokrBVdd5alR7u
JreOkrW+OGr+DmAtfnWgk9jxnfoFXD7eZx77ACoun2rQUPyp/eH38mOV4MLm1LdBi7aOfXnglJV3
h88zbefCM/lSyOxnlxSXu3hfsHizISpHuCfn7JMHIo67jO1WAPvAwqeoltYtLAW0enJd82LStR4b
SNxAygr3YhuWRwjLLl8pa5QWl6vuTwnFh3O/XEQNLbPON61r12ka+59MmGXJThrxBmguDHXX+NVf
E2Ds6AOCA68bHZbmPIQFsuYFb2N5TOHEf1/oG0VfgiC4oJxILP+pjVytLw4wqlhBlN/4qZeVqF41
d4jb9+mM9cxvDkUJyM4jsHUlcsLjdX9JCBm7tteyupdFoEViKnBe6/Iwq/IDp85gBE79HwtH4YLo
ov00rUIwzwgGAh+dDTkaps/dUI5+uePTEgmxyq4mMgnO4pOB+sK0qFdChxyM8c5Jl8aIVxjGQfkR
RbS4ZTwm5orIEvBge80bkG4Yc7VGNyet9Rkg6NoFqjt6NV5GTuhCz/LnN0kU0pGQnBaHprL0eXVh
41XKhiKGiorOSIWIQocx3ee58opCBmKNd9F8V3Uhz02CX/Nbz+o2Ru4ktXTPcHvgSJsncMPtri94
1Luzt8lkJidibyXOCbFuftzeVSeJ4ErsDwn6DEg6Br09ei5eIddIlrhjNPmpcEj3sJVOiG8ACaBM
3A50CKW9YKNTTCksuMBHcEy3LiW31m226riiyEJ1Timc3uV3cbA205PwAMMSwFBgA0WwbNsoL46m
SsU919spF0CwWj4vIYReGZUtwSW+JNpPj8zOnFtZPFpvmRtPWLoLPkPhr4n4Epfa4i46016NpbLU
a510H+M6aMZ0xCLeGrcD4KJGnx7+Rhyw7pRwqy6+VOIwaiuMqVYXi2IRujhiW2owUaq6v5OjUW+k
lNohDhbArWODDUdpQEA131hpGOAqOa+Frka3jrcrsz/s/tKrgejCaKup3x6u8V/hBXtTmjUCK8xy
FA+0ukm28fUQVpP5/Alq/mhtorDxJbSuJIQLqaVJnEqNoCcQWjaIxeDLb8Dbz1gvvMa44QvTZEq/
i5sxbFVTRJPm3D9NK9vIhGHMd5xAfqUR85tpf42brgQyGywlXTuHgDyfujoPXabc66ECMlBYU+zG
yYEPu5HwDhT11MSyLdqlTCuRsrSbzONf7yTFpbPI91AAfwRpl2bwEQjc+clDleC50SvsRkFEX+WY
lWr10+LYFzygMIrfFNLfp0IvMkuCHg8ykY2LkDL+U7iMhP4f+ryZIEg3/tCJCiIq3xvTqzyDJ2SE
XFnK6EW0nwBQ+32T3yP1Xyg9gK3/jPNoMgme0aKdxSTYRmFC41QlB0SvH4GappoYLyNm9mqTU6We
S2+ZC7jBfyq9xXGRUISCYK0kE9EM5MSPzK555qPiTxnLK0ih25oZCEIKCK3tNv4WwFMUCgZZ4FTa
8j3fW+J0JAUNl5eA8wQzhliVp28X4eho54QWQIEuToenAj6HAuiSS/tO1o7Wg9hOZYrweMRQKA+w
H3mZqs+dhRgOsw/7+IQeH0J2NVEHtudk7DxULM+1J9XJaOhUbZfBQpSwf9+w/U2jVrA80/zhCGji
BPUr9sX13IrXiymGOYSXck3MLJFKESIZEJHsJ+yqM3pnwrwrhvUszNHxqIwWVIXTFcRFgQ+LVj2q
E2xYUAlCEeHaKTYycmdcRhwKH5zBNP2QNCc7FBoBhgTfwlaqKL9zFq2gYfvtxy0WgjUdtx9iWiIT
7Ye4Az/O66q9luTBNowvD2b9/uDifenpxBDMsMwZqtkhIcxjXfs/fk7gtRWhi2jg5SWhAsLxwNwo
gfIqWwdt+G2SOSwYrjWXSc9TsGByzdg5u4Blm8zfkkRNuedZ67Oi1R1ufZFb/BWlCP6JKJ4f1oDN
NOKdGYlNaKhzAXi4K6jFYOAQ+tLR9H4JoEh/tF40pW2FSlDIckf1uUqp8euUxh3ug+89abZHYa4E
G2hurWsiQhBJ1e2Zo2tYc9bmiaMJgNea/mw24B+4B4fP+XQTPxzvFxxzArYE7/kLglsUB1zuxsw5
K60byTtzFrH12qpCMJP0ft2FEn//Ann9FbGofB0HttmFbUaJcnK7DfjwQJYZFyiVVDegqp0QR4cs
qeo2Npzhbi6nbyBDMugHBWblqbbS8E1UiFN4cwPmcuGUxqEETp91Fo/2FYBXKaAwpGpfucoO10Fp
8Op3jXHMyncIiN90QRaioOoRGZ7SBufK+S56vwF7xvLh+1knfbpWVTbcryCihSWz2HcPV32jEMEC
IU+HtS9fAmovrVIUqwOe9hb0G9gP/YWDnQ3/Ch6UM8PYsrypVVkkZUVMN3PfqHewzvv17Ldbysqc
XzKyAmOXoCSAMsNIbNmsmLlxwI6/5p2D0pki/RfLpc4WhjgCKb1nRebScUOqFqCCjJbPun/79zW1
Eg2Q1VYJuvfA7z7et99JY3BBlBq0ib6/uVu+A9kkBa2Wt21CmLgJRurcAz8LsEQ8ORm/H2wKoY1f
5y0ZzcjrONmv/5zPpOVr3oMn9jF+ZE+sBG8l0iaYFR/k6DwbzwUUMwp+/DsPcPn7t4YUGbC75gZM
01OiELtjXwp4vDvcnMnShsokvYN0VerrM5z6OtAvyxNnE8n+rNHV7ekBWqdInH23KlFxS5tABSNT
LhSNsJmzqoL10Xq6FR5rXcY/zAJBMenCobUZhu8y99tfc0PUFacXb2KvmNy6c7ATUNM4jKbibeyy
yHDYMRnEAHKK3CZeQjB05YU+/mbSy/cicsV5NJNxQsAFbJa152+1ky/4sz9K11dSpUaorPSDIZco
acuiYTyn1y8opgQPJkbtw+3JBFNNQsiUhLGMEqs0o/4hL8Qq6bIULMlESlHkBK2LcTVDR+PoMqo3
ShHBihA8qX7iKXgqf/zXVSXTeoTYM3CY3LPCesdZy5UVxNAcUU2xI+TtBdcEbAMg5qrZdkeCTg+C
SbQx2mdzQjql8H1vf2XNdd60nmlPBqbtyPT6d6f2RivKRkj1iMpx5Sd7+FK8HZppGRw4v58IkdHo
khKGlXZ1NB86RtlCqMQURKTVbFKcx+irLfF2NEYxQKwzK4aBCfT6255ciF5Jol+Nmj2dr6LuP6IM
wxUIAAwNY/f/Hq/WsASz1nwNUlooIkDoWkAxMfCxZPHk+DI4ebNHOILKcs8a1HO0Sjwp4Pvd2Nad
sP9wXcYtye8xiv4Z52V7+GA2+KkUBa5v1pssMTdzUum/8XVHv6mq6zZtRtFGBWz02OVHwsFusNtm
TGanjRRL7pp13kXz7ipD+r4tSZARQ7QF12bvzE4BkhrBfdWg0D6aC0VJNBFIx6CJlp7zGs4wFldy
NX+czPY1lHTApoNgbgMlaiR59iftW5TrLWje9Y3BVF46ICIIIUTVCoKQcvNxRtIidrTaIpLBjenk
6M27UfSCJYeEnig3gEvHvYIQKihzNJP4q3qSEhv2w1XzIQLtTIjQiDUVusk6sTgU4vaTbBsKQlhG
e/cgSL7kXkzFNe+wiEqsATxDXOEK/3AofIhjiJP7QAyridMyDmdSB+vrEoA2IxawhmFDQURzb64I
WroU0o9ZHn3foO4SlUM6c1kl4T/YRuFjPgGs8nrTfLtTBzyzE63wRH3XP2mJVU16I7StHS/hw3Ul
ltmT+naCAPkpa+1+wDPFaajAiKVJZcQCrURmOt9cc+uiRiB+foY0LHEp+iFxyRyhSI8VuT7LnTvi
t1/M2fycc+QaVukNInJQLt0BRvuXZIWRHvZBhVKWY4CM4m/Pso8kB7+Y5E95rv6wh9/pqYgf5S7i
JmrdKmv1BIavtdXlGzarzoE1ye7bCyKCCM1VK7v8sLFhUauOOUIUG1CEqSEX4ubT0187JQYP2Vta
3qr07vB3IrCcx+cPbmdMuRw5hIcZI+Wv0cYUS+aqnvsa5NAfHbaYoalZGsHdsSyfQSCDIjP432B9
3wkKuOHPDYOwMfFMQY9xsAHPrY+6X4db5y9nN4sratZMANP0lMH8feiYce8IKRGUZqk+sWh2tUJF
2n9I+jfAZ/B4L+1cTzMV4lGAbEKV4ebtjKRsUc40ESz2WUlIOGbXhaG7iPUHHCTW+abEeKQEdFWu
OEgq5WLOkPxVITK+uoZG6TH3nH4aux1N2RSpgBlM0KjiIl8n4LUDyiZxPeCf+RSSYs9QF4rC+3Ow
1CmJY906hDcd4QCqpq/CvDQZ9khITjQ2EzTqjHjo6pR551tzokmkGDNb+e7Cja1puOYXegxx0nhq
8cbvObPmGtHHs7PFvC43DgpEQGUqaO3CgMliVDCICMGGKowSLRPUeCY4M/LBpS5w5UoJo5DhCFIV
Es5xb8wuPKYM3DOzzT6Ut80oXYRbbJCIsWw3I6XvYrOjgFf/7qGgf5FCs3bIZpo6JX3xjlkgspLN
sXLcW59tECtBqfYkKrMGX259mtC8t0Xg3EhJPANH26cx0QWbNbrrVS6eKUnP9U9ezaoMsvp+iiX6
baFJmiKOGHoNKFSdofMDgLyvFKh8hV1PmqPbYIJBGgAwY22tl5Oq1l/aRAJDHewqNeuLQYFi984a
FZLCNjC7OgQTJLdvOhF/Lj0B/R76NSauYP5IPastZDCLDiPiIbgfUjJw3uxgHj6rnPswZF0vxK0w
ZzJmWStEYnsCuK7gs4E2AknSW7nAb8MalGnAR1NHuZ40phF69R2H4ppvm3sPhOpm4ABlNGdVD85Z
Vpi89zeGOnmH7Zm796AEBIkr2xl8UZlzBwm6ipXmtnR5QBjT2kbVA6B5lJvu/8bHgx3Z3g6kK71U
TDSR5RP0nfKTF57dN3rRDu5gxnJ8yz8uztcNHyJrAd3KmhkUmQWyO93AP9RY8EBkP/3AvFYeRzD5
gqd6IIh+RV1dqtP2i4md95/IflOF+fkNrXRdhtk9F7jKL+8hEtJ+Ud/GBWed39/fqpcur6hn0kq7
JBQSh7nXixSx3ocVpyEiYrxUV+WhsF7IaOxoK/t1zkRI8AB3NzhmjlHAX5JZwBuR03nkmwI0VqxI
iE6IGQSz6I2+ojATY1R6hkPifnM5GaMwCpWEuSV6sbDwTqqtZX1C3iYQMjJr7BPKm4ucCoVyOzya
+FSFZnt6T2Etzu4BkXLRIJZYLZ/EuudJ5XEDVhGk6CuIsNwJ9Uoof0CCGXbjM1DkexvQhq6hK7lE
Owt4RAjkF8v9HL5DSdow9UtzIcaSc8vfLl1fybjSbqRFYspeB90iTTEFxWncMVQcVC/pGajvpkmi
XzUAzB37PpNlH0bPQRBa8aGk//JkfJjLVysKy97VQYhNXhBzwXfsl1cgygjHPaJ7E9vSah9PjtXN
MxoZLx84bryejz612dLgoNCSbADZYyDEhc5U1vY8/3SrB7M4igQD0Uv+Uh/enRVGZwp/aqHaS9OJ
Nuwq609nsDRtWB3W9SZgC9n3guJq1BnXv2QgtFcNovyjXVXGeN3hOCcjd1Txj11N+w9JZRa0d5oU
XvkqmkYq4uZLeICLmYJGSHlQhtTTuK6cs9W4WL/Sh/An1y6a0sfWq+hXVbBOS7j5VBaPv32Xq4yz
Vf5WDk+o2uXyIGQNqlV5KZ3r+mdUzcUsZ3QMwj5nnNE+Z3GQx13loXq+SIycmFWToehNmKP7LpCT
tXTzoPECghlt/xB7nDGXTbC3bFTgwitu652pulzXYJ/WQ4gKV7AJHBFuYkCxySdvIPRZLElgYu8R
gZ6aA9aeaIDMgOpFKSjO0oArNnDGABdZlLaHifM1eQzqvpe2rNLKjRhmukGUP8Txf2lmT0CSe6iB
VLEKxYdyE4yj7PPnxDVIRs06xQj29/yoG/PMpMpS+7b3X6NDzkXKnTU9Dcsbp1Yfk2cVIFuOn7zt
lUy8vSs5q8319lL3/o0KIxrl0qZWsJLrslL254wNF8/Qjb8NCyJkhdFxeVDS8dL3OM7HHaGBSeac
2QO9O0d+FF4kPWb6ruOrCkeoJOZzYLB9s29shrWfN4ihPFMsm75vMvUlY1mzfOFA5T5hGUhteIk9
J7D/sicbBQrTiOYLQpd4rRPP0IHWm+ryQWqOxoTWIhZBQ7rI8xCn96ALuPEsaUv/zd4DdLmp8HUf
Zb2LAjPM95JjqfRWNL3zaODf2C4ejXzXm0sadk+pQuLLElXCZnmbxfy/Be/FFZ5Ol8TnclaJXuPG
0DHVeawP+mu8Pgm9rcAzPx+2IghuvH3Ak/cUdg+O/9smwkLIcAFTdygFh7Y+oKVlLwzZCOvP1BSi
HXs92nIbNwHGyr7JJEX5BmL7r/APFxEPLOTJj8LI3jLEPm475DU19A9EAwVtZc3D0DE1wqjiR5+g
QNzh1XLpZosbhD4FRSRaPsUS7EFoN6MOJcN6egfAAlAqg7UGJlCZER6iHQGcSZuVql8cWGn/rolK
gGhqDcgFvengj2Do7MrI3hORqvW9i2l4pXgwjN1iCnzaOGhtAKIlyMvrVHgds8T0gUMx9hQ8VUNd
4MH6+rVVByMgOdGAKfRSRynavG1RLtaNT7i8JIuvVQWh6yCFOhpqkAa2aBEjhDQUqsVCqFUxA+i+
e7S7UqhzFnVCsVm2bzJDL3frR1MSHP6hovpOnJymRycWxDh+SOwqiwIUpZjZefZSmm3KDMQTQ44d
lciLAM8yYmSSusYGCmiiaG942XVPM8OGB6a66+JiUhgfDu+yiwBi5jC+HRvsN6AxhT/y+voQa2HK
iklfKpvcO3VKgAMogr+2m6wUjxljGFVHb5z2T1T7yxRNVGVsZZiCci8FWRiYFu4zNdAooM7y+4QY
xHV4GsNKAQL4zsca4Nl8/Zt7pLc2UoExbDFmPmujo1SZ0pbeOGmlRx690ccFahKCennRJpU3BNct
92SVNmmBKOdiMkLneRBx3Qe3+50Jmjhy5sVAJW1v+SqJVKMxKilsCIT3KTHFAk6YDxVOlFSWXBkI
Aj0jvmZdmCZZTJN7SyNg2La2cKCiF0gvQYdNWtVxw9v5Y1LGbMSUYE29MHuF6ViibOW04+QcQHWa
OTsDg026KxYvTefGkItnfP3GWkpGLl3zKchO15khJk0Z4l2GOtF+s71mthjsmY1b5ktzjGUd8izz
Q3Ubx3q7XaUHZqvaz2P7cKWLfLj1zX7t3Bi6bgDjq0FZA9hlEpnz8PLPczIPyHl16lx83emVBTs7
TytHw1Uu+H1PABBrQMoQ4cPVV7W0wLfWtiSBYXTE9IUqOm2R92M7yFPo6fP7mfJjag/02AhzCEUJ
ObK9NqwBUUCjLwg+BCdOkiSxPp+a+1omdZA9x7ykKIwJJEtv0/kmpquItAYkPTaUWC7j+LEv8zUG
KxiA0Ub9qwa9IH+LKvyQ/Amn1QQzc2N2hofINf5bpeiwnTv91lytwscW8zj80Z7KJZu4gpuZBj7Z
sfm2GiVkMxeLv/8qQH+37xMJuvZfM+paA5DMsleza0LIR3I9JZJlme+zZp1Ak7sIMPjajrtkL46e
rVYyjIFvU6oPzbVoAqNzkDaZifYgiI+5IAirDaj1V7w2YIhboIQSjBMPUT9ZrQ99SHbVvUy86JGP
/Dpdsxt217NCakTKBLyJ7jMriFA0RHpwjMEz9ywPBTGY+GY6AgetaC4gEEmShZ11uhSieRFMqZ+u
OU/ioE36ZTX5vu3Ye3dB25RnB/PnJm9jkkQvWf7t6XadOUynudWqbESZQSbVvT/eGb9cU/gbtiSi
E6a9dwjX95IxPw08FQpnl5lNmCadm05iO6t54b+N+nIjGs4DhJhN59dkLeiG0sbit8Mls3eVyAmZ
A+kLD7wJe+MIkQsxZeFasxLa/heBuu1oAwzm4I9r8DjIe1SMwivFKyQiW0ZpuX+oYThhdw5qqPtJ
qeuIqA4nZqDGBhFtE0/jC+sRI8ivfUkp8qgGmn/TvArH1lfiASucxrFu8suIyEolA7CeeDYnVLhE
DqgmR2BnmVM6tQd0VYKN6gBEsCYbOkePua1DKlCZu2vcYUPbT2NnQxfn5+8xG8jOWDEGF4yVX0mD
jZq53p6uxb600AddTKK1GWxW392ZNFq566fR3LAKQQv+/NUquG0jQhJrFEjMo8TlWGjB/kW9kyeo
7UO/dslTimWIYZogwtKBC6D7e+jS3b1nffqGnWPmLePIacbY+ypN11pdgwoVE8OxdNZhoms6zgT2
nxn6qHfAzFJ4MKnOdPAimsCNfFzC727nYondiRLOq1ZXdZvoN8WKrTDC38EenQOiIW/sPenXyaVx
gj+OWR4ju1vKmSJrP0qvHzZvloHUDZH5lqB/FoNOgyGx7PmJ1c4JAleGbtdd7V6tc0ZIz6JGNnKW
hlCyxqwziB04anA5Rf/P9zx/2nCh2neHPrt8mrlAMQJysmDOn6aiJEAEL45JdtTqU9V+qDlQijrk
MnaNqRwOMHw2hVleXBkORS98QUNqmzHDn1YyKc6X2nnWlSuDSA0dD1bxwLxvvCRuQ/8nrCB22wu5
KAwSG3IhELkM3RX99SrJ5PyI+VYM2tOdwL/+th0dkz6iqcQ68yAhAYG3RRwjDZfhfcB4eeWpaAag
eaAL83m+E0V5J698gcJbFEOwPH8k8zIQlORLmG2+K6ZFL5JJXJ8fodemvqN7IS+pJ/QgYv87/2tI
mVhHJA2Ic4YeKPiR0iA4fQtFtREU0Jv/NhCGvzYaQM+RqX+nUHENbuide2QWOxNjkALao6i+04if
r1OKXug1jGs0vCXcDwFH7cHPyXgDp9xMqJbSdk5gw7NLnJ30J3XxkZjTXhEMEcsgb5clN4He2/J5
YHBJmby0HG6RAyPVY56TI4mHsQ958+wsbnY29MbCcG7MfezqBfqkPQW0+ZUGPHV0X3Py2t1g2PUO
sw4c5/jnEKp7xoUy0wckQr75cbu1Q44D698FeGFN3NtG1EA5f4qKcIf03UOlXkRkuiNe8AecTqxa
uaOsOueqmQKkwJcn/KYuXiw2hQRjUaRoR0QyiXWhvxaKR4Z1bO1rcMlOURy0OobLmExpJs66NXpE
IjUNOWlqoFfldQcUi9K1f+6OR5nqrdGSRNYZJcgTLAE9NeYuf7vf8JF0aecCUjgpLC8ar7GYkHXx
4h/DM5kW+GEbr0Qi9HEsVrTC8j+t0BOktDpJhljPWKzC9fA32YV+vlShVK7vQzny9+FvOGbMq+wj
Jga1KjxMSeYtGAbIPVFswBErqLjKGdfk/dQ4JQbLRCSRk3ci7G/cqb86jmzBj7XjGxDcqiC5YGb+
P0beYGml2SL0VCIC/DxiX3+nCvh9sf5nFLPYUECrdn5jalbO6kAV/kKffytST6zREppn0AandJs3
ppAbzReUHZl7X61VtookfrW+kFiwebbea6GZougQSBP2olgKRcb9tNeyUq2z34ZuPReJG/ODtWqq
J2Lb8ditnojJEfXkqzCFNhsYbJPiI9UAgATo1MzpPEVQdUWsjI/FqQN9a6dc+VQpMYoL+aeKMhoy
3HlbHiWcYFJr5LUGy77M+C2XjWS3YkzWaKvpuPMdQPTz5nGB7BaHpBodv9KVXgpBJOSGs0oXe4CJ
kwfV7LDm7vHJhubsn6YPPdswM17idF0bnI2LJIJuYx6rAAW37OYWC2AjTUwc6ynVQWNm8qzCxmwn
W/C0BlsQGaIDaHJ/zaBz1o9quXQXJmzCN44Ut0ENup5cBRnTNdqsvy6htmHq9d0lZlqDk4CiVvY2
N9pChC6pcibyt9AmqztVrQVMH9+r3pgUd98XtrZe185PrInm2xdI2jEBAt0rPkDNTM2uzp/zyvak
WYmKrTcopd4nS35pqlsMiVsBZAKBF3UVVoA6uVQx1N9mwMH6xXtiKWwMfCTkcbE0AdNYFDlsY/CS
5Bj3drvWknrNCTZtxiU3RAFYQXHhOyO/uV8wqws4/nnMB+8ys5qUDYynQuBgjw99IASFBVo//k5p
ua7GWilgaDP+qvk6z2T7/D4U+N/cFManOEV94Mpau9hqb/NOWI6cYtLaJ9/1yWc05ICVYOX7VAgf
gQ4PTlQEHU37YlJCoSnsSKu31YgRVKggL3w3w4LvrTEOo+OSI+IqUCv0f7rKjvWcnzdQ9o9ipac8
H4SowOXGh6sZ0hVRalJ5d+qB0iBz88bpJ9u9nzYzGd0F3bii7tteJ2nqQHDk9sItwBcBBd4Qpg9u
sj8dAudSkAnwL7d8Z96XC7Nwv37CfJuNUdoe8v4/kXrOfUg+WR+YVJlQl+xPQUCl+9s2aA3x+TgM
KT22bRU2pPiQc92mjpibuJP8evGaA7tWXBG8ozwBqQ4/0auCdhkB2v3Ly6F/r4UqXtl4rMuYJGKq
FgnNT0SrpDyAHUrIbA+GEpZGQAX1Lth1vnromGuPGSnplwRBVwZHj0wXjIEvHwtiNBk54PYc1E79
srfiL/2dQTSuNMYvmRCTi4K1XgTAb+lAW98dnMCccrrscGaPZF7rHItotqmRfgbiWegRTaCOXA6c
5e1bqE2K7euPhu6+Ae021bJZootWhTcYj/Rzq/p5P/cBDN1/mMC88/5YaP7cWWLhWsVd/dgyeNru
3Ms6/0cA2j51YIL874qaIv5alGzl1RkMlTl4cio3CS0CAMCBcGH+0QX3B9kFI81kG8uBVNg/xSDV
DvLI1LvrkGrnazkRFaWF1pxyj4hBd7OYMTQHXdOuBOEBYCDZ6f2619a9Ia6EaHAvhuKNG9ysDtnS
5xE75VQ/KMoQbkcWnlFwoTd9xjK+MZ77KyzsfZhsVfytm0ZMlIH38AGRpg4OWe2i160KlPANi6Ms
iFlpOBnUZeTxTIHAvebVpW9B4047YJWn3ejKIh+kG7ZgBQt8UBtQP+9UQEIBiCZ3cmxCFqRbKLXc
gu/qcx17LYLqEdhaNMxIvtIUWJqtEXL/LXrq59+nnrgoD1IvSpL/qpleqYXLYlZYJ3iN7G1S22nP
o2K6RZCim8u6hADvFi57PG4Ertpkusp+HerSqfhugXYpvCZRHrNTat+fBEYRr2eWMjZ1z7Oecykh
Sg0AW3VjWXUycKEDJllQFnjgTmzWxbsL1h/Z9ZZtVCpxMbegGkgQNIs11TNt/ABj5MyuRClY/qc+
OyVt/Ts2gSu0IUEpAe51GC4JVnmshggb8JoOd1O9TfHJRtxlZM5tPRGXBMVgiEevjmw/Ja20kAzw
OHvuNzYtjVPJTfVHdplp3yHs9pJli5ZvhxAmsRnk9Ct605YNxRn0yIu9Fa+vcY06jmj9arr0sPSy
SyqtrPPUsiBcPuC3cq5yPyJLjrmcnYBE4O3o9MQrmPnlk+Dc7uDruKfGwONLjSg6JACFS5SGjMD/
h13MUXQhQFttt+2vSo0Qw89CxOJ/omy2boXQYMfIZ1vBo48sDyCNlMtE8fePA59tiw6L+i9XGUyC
fgLYEDMNys001BlN5GnGKkKeSCGLP0RnhmuO7hIjmqQKKDNhCOhwBeaDCDNlgASJpUAuKZBSOlvl
ZreyOVIiu7Qo2dL4n7fFjHNq6jkxrol51oRQC2CCqC8bJK5kE3SpM6DlpzPzdWjQizVyN8Zr3B6C
fSP9hzsGRzBusT3vHt5C0j+yopazxthXDWw5L/ZQ4Sj195fBQ5k2uayIvJEvF0dBXFvV1AGBQKhx
mECJ1YW0LzBSa+RHNSMtNa40gHHD6GlzlTbp1FavRym06m6/W3HuNjab3Uh2+jL4Ut56VtpikTWL
CjMeMf296kDDn1xCl5yF8BEjb1DINozKJRlV5FgZVj5j8Jn1hPy+BuseNFI9mzSdEFkEosdYuFH7
qZ2KMPc8a1VTKsAE8WS1gawQjxSkvJjHo6mGPraR7SXIWXMnGCR3G/3JrOCDZg0iXnUGct5fqb2T
DzTJeTXC7czReGR65xcqfFRlN3e6Xf1gKDV7DTXVn+baOVF++9MkJL6NnXY0SFUaonwnLybST+2b
aoI7ivN9AIpH7wOpTRmhEf7aI/ecu6sceI5EC2B2fSq2sbxj33px6nGGMx/6LsXYQJeo1fRkpySY
eBjTppF1fJ7P7prh3PPzJEB2VlC8f4/0DKa1HTEGVWRgnIjHISRClkF6xc96sIc7NVJr0967+RVe
xSkfvoCacRll8p0V6hILj4c5pEitTjAHwK7BNt83Wyf+Bo8kDucjiO+Ndy9a0seVafl/5nzUpUnW
b+CJi9zTYhUfSqEAwfFrN1V08dloJ/9UI/eKl9oNKXGtfs492wtCeKYww57nS9sBU5qvAuyUToNl
fK1fbpm2JazcCl6mFphuacUz2lajf+xngZ0pmmW11N+v5WPcZDfOFCz0a4F8a36poaWQdcycfwB8
IxWDguuWsKmtfpoafou/msz81qMVt/UfREr9Ho3zxwC74rXyKgTWHdhs3UUfsbRBR1F8PnBe6uQD
ZDy71tFd6XmWdZtowZrh/orWdZ4tJOVB3RT+qKMaZUgzWM8UCblKY7NpytSQ3UftM2Zx19y55Brx
GLC9NCoe018wELgFmrQqoCsMRrO41COhdaFyCxThIrFdroxEmMoWwAdyC3ayUBasIEirBZ01+rou
fIK4tf5W5B50NB0H4yGiY9bYTSVrfGlY6XCGQnvFnDj9/HXH/FDNHEgQuShCzoxynEA8DLzKk3ir
7hZe41FUvv19CxYbsGtx6oNaJ34wtY/xMwFl18eM/FZmfGGOML1NfIWqEDMrbmjdoesOxks3Vj/x
Ruvrfl3YOemUic3P72fth+oZMR/Qx6lq5QJG5MoC0gjRT6UAGYtnOH/GIJ266354mSsaMPAQXRwo
jaWsxJOrp3atPS+8iBw4aNidMgKWznhgjVM5jbV9MDBcWj+LBvQbcOgvZsdWaB2pzy1wAYnuW1qA
SzvBisCX54hmMY85QcAO5AIZxbaw3xHmGV/LSMbv1a0iixVsZLxtzWHxARCdlLzd1zvkA5OxAqLD
DOBmWWm0faH2VUJpC/9BAKBu8MOcKEvzitiVgKm7dRacAo8JT0+5Sv7eeeuPlLfPl+91CfSq10Gl
FULR8xxBwqn64veeclGZuoy79yhWnWG/yqaZIZ2+EGA+Uw/RHtRz16G+7mwj9+n9Tx6wam9OB3AI
NajSl9lhCWydM4VIb14y9g05nlOnwSvC7zeMAX4KalHFfUSbcSkSnf4eWrBBQ8rgNCTuqmCAjWMf
S4BZkR4S7qskxLXtVGc5My1gd4ilBiFknMhh7Z1K4fvWp3e9GjukGk9POLKANjClt1Govs/W/e1k
xL3Tyv9JOJSqaa20GPYha3IcE4miYsp7vQUfB7kUkUtw5I81iEHMlPx81vJ8iq/43mTBhtWastgZ
Qy0xk1uw0m7Hm4OSl6jAoWK5PKxjN0PiC9XHsdKPeYBxh85pKp/gh2Sg6QrBWEwphzQwzNXkrYep
QkrSKFLVKHW4yMC6/z8mNIXWmlaEh97I9kvSeOrPouv5Q8+TBv3/Ojgm3NqgvVp4U3JMj02CIgCo
FWIqN3QHFAW+W9UAMq98X6lKJ9RjY416acxaB80qgBVApIlmFMgGMfe0BfnvIbVk0OtWLkU5cf0o
4eqP4oB/8VBqV7mm3u5orMVyXdlW4V70/Sc5sg3gPn/qv7ISg+m+glXxTPQbKg6AcRWvZi45pUyz
5KmFWMBSfm3di145lgU7T5U975Gbw4qa52g+SJpvbHKfgPgqLvhlqXYoUtBiZTxEaxcpEIgF1pfZ
fS9GBbPgORnBJRUZaXsPDL+eaSnnKq9h8MFsD7Nhl+hoBAZhKAmHFJJ7mUHYeZ+s5xtC8JNLeBES
e0G5ZSKr6GzxprmetMlv/zqHmjmtbXhsmO5Tg8aY2ci4rfL/gnq9o/zpd0r6tDsqCPaa1rUkiXRN
uBKIYTYyWiIv3W9v2WlAGLbZC02QqNgd8qLz9I9CAmFR4bA+68Gme0YlXb8zwB6BKz3CblzRoZyK
Lf7BLWxmLqELog/S7NwMW6rOj8QFB90jCz8mFcxJaV7fD/hkvLX0RPTtq6lQkKdEYq4wLJZWGOXW
Yim0OQtcScPVd1NRYPx9lW7f1ew7628brKx3fv8EyMpQnKAPq7Z3Spg05Pz1/yOnhfYv4ViviOyE
BYTwH3Ad0GKf8E5IgChb+KOKdz1oMzTZNiJeEsssSQ4dYAqG3emc3lPtdXq6hvMdVsJj/eXcaR5I
RSYihZE7ddJrwPj9JjKorAGgbhctWsLGBaobCc5IiIg/+4fTsFoLfU/jCJwhSNYb0xHGcSUBdVRX
U1Mxijf6mSNxutMGmqeN7uAQ3mPOn69Qs0B6egIFCzsQBsX4UfkdQ9maZu+wpGsmwPS/7ebUaU0O
ytQwfHnaPZTOGAWdTghUIQ==
`protect end_protected
