-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0T0i7nOKz0ie2K6llV1SjCJGCE+rjrR5B0d+IE1c8/l0m0qezeA1VfwMDldNLwMIiH7kDjFzTn8i
oWC/kKroOHTKIrlA7uWiNF47j4rZUTOiOFrRsJ7h+25TeJm8V1LuTTxRK+DNHhY3MSH9rwfnu+uG
o2oCLkKxWuO/yHZifCBJ3dq840QXEAeCZiLr23jTNaPceHnh7blmskeplcNMlKotmGRwb91aMcZo
u5+Lb3EtvE3Xbtcy5ESZYKIMUTI+/GCdCwnovq1LXQs41UBbgnDrz0nE4VitSdjtsq/ZkfENWliY
dF+1YHZYvJ3bNbfojcWiyAysyhwsdepJE4FMyw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
buY0jxLVTgSvZUsJc/j+kMVmDH/CbcN+NLkn3tLG6NfYuQE8HMKEjHmbm34iDENFWnWR16keJa4w
S4N7OmqHa9FVjxBe1aHPZw2rfxuusnVRT5t9hiLXo3XI5Srj5pwfCfzoWzVhfGf4HOM+0fHcW7a2
S/KfIbL95W+CY1bG8CZ/Dl6lfCsLN7DILZswmKDTGITII9avicHEuIDlAsmLwfxpp2yT6x5bD76Z
A8X3e56YWWd+qP0Pq4VN1p9jye9ijA+kqK8v0jp4F3kXhpHSVhJuijypp0myWudDD1DwDTvqyhLU
QWN4kaFIgE91ki/wqyIC33XkvxDoTl83/YeIQy/YMPVb7Hd6qAozertUmD8UWKoakN0YTQwB2XF+
/70ltHvYuRF9UNkh8quLdlwGl7Ym9GRJY0A0TlH6YsglXJipG5APk9rNsiL4WvCNdxX0iKC6rkHY
G6jFHHI1HYWSgqUkDyuDhxpOiNZaHSZZFtswty3LhrXagzd3JaEfdQeBLUEF/PyhtDmsN5wzhQYQ
VYx/jqf4kV9CsvMsm/XAuENyywGNwzl/1CSlq6OR7YJdI4CqkiLbKswBWwShT0A/JJxNKdXZyVks
LKRkTwARjboH9TsWA7sVJjDtVHgMOLm9/8fUhZPGhMoA7mEzAOnEJSBrSzc+v0hEHA65rP38YvPy
6np9yXKHq5fBTTigvrGUOXNWHLyDnMaGBB1XxmbaervN8iYPuZX2XWaknaGZHUbfCC+rYuMU2uOx
ikU8SF0J5tUpOH6ghL3pXiL3BDm5vI6+2SoS2qhqjtcpnPYwrg4A7PHpEe/CV7Viqy3Th60liv59
rkCCCbKpsTYj1/rD823iwtsReO0f25szn2zEL5iXpVgQbqJJ6ES0JDIIUYNoiSEDGEPOlwGuiVbL
iRJpH7XI/bAOZZm4RqCCAlk/2Nqt0HKv5OJ1DyF4MxCjPd2Ba9iJKJHhYVeq3uVE/ULgDeEBBXui
lbgH5px4W1MUb+3aUI1SUPhLOidXL1KnpAjfNu4tFnLGDAW+jEwuIP2CEFbkfyAlAvx5jrqypGVA
fHWBYC47r/65VwjvSlYdzCI9Z0xnEBb6O5ZSKiaKnjC2q4YsDRyHPWiGKzFi1xGJUeklSUDnEmFB
XfVUq+zTkD9rZyHIVDroqTl8w3v5NE9s7Qx30PyayT+Jn3fb8rl5CqMj1+n/xH1q20w0wb+EqtE7
rICytq/yVX7StgnXihUbP41ypzsw4eCvK9rGRT0AQnCDKKhEbXZdk5vfo9am0kP3pYSWhm6LVLpm
mixhoA3wpGfrdYQSSPFfaQhd20o4NnjMZPDXrZND279U2ip4m7Z+V2t/AeLOpqM8bR9qPAu6cQgb
hpIIZrBf1ri7DjDuz2+yQ7X8aobVjf8om3M9OtX39bNAm4b4RC6RiFDwTag0ohSGfb1l0VPmJu2t
Hme/iJWzASsl0JBygkqoHNYR4U0gFVRjyPjqtewd7PGxgJ63+zNJn7CUnoLZEJd5jIx/bjVS29Av
QvbFx9p4dXPD6JGsMPuKZtkD5WuvBxNssjMTz5OOSmutxjrfpGHav5qcSInCNA5AcUlHSawWGsRG
DABpDTqSyzfMcGgR3hN+VupxokAxhQ8xt7qZdKoas5WKuixpQ0cNAqaA1hHaA6ow3GdAKp23I2Rj
IK04dwc08KuzBHm23FtV6Mfv+AtelTbANToe1gUEkkFwycmVLc15p+eAVe29CPBDANejdT+c8DDw
aWHxmkF7CMyFxREjqSHOpEiFPtLGykseWPv13lLkKgQXQoen5GSjCsJbdTx62VZ04YDZeAMEgCg5
vsC96QucgsOL6+GxeVaDfmcOCDy4o08Bi0VfNhaKhK4P/jQyuV9brDxi8Jhel5kbUpTVWdqhvhmX
SI8qNm6P80ODiVQ0fCaut1cnT0iYAuGZ+66hUzi7FVrAlUsV3z/HGrBQjoR2DAmEtLgqTGjrOLiC
UVsKaoFAe0pcs+1OiXQyW60r+J70j/ACPu395mNMffuKb1s1ZjSLn7+DBzo/lbhv5Ma9EgJEIklh
wz7d/f7Kw5cVEc9aTh8b7BHDEt6vmusOb3EOtnb2zjLuAK+Jd4Nl5P58g/1eQOvehK0cxPdwacoh
PQK5ojXEIITBNMQP9oDhYI+H3VvXYweq5RQ8wTJ/2PiS41IRjVASQD5H+IfT3ysABBoyOFQmRi/i
L0+XFBtfSaH4x4KPwe2HkynN+ntcUZB/o0pxvshXiAFMfw5nIib0Msw2VXQ3yYaikCm/nXsQARgM
HMNgHAKqvsokopEJV8FcI7CrCRH4vDEOhNyLXJsbIrH9IxfN04szsx67P92hekiME79JMkXDwO6e
mZzlKF+GnHhthw0FrwuL+11L1nv2S39tA0f9g+2j+YMNgbgejmu0jGw7zQZ3jkMupqu9PVL3zRbd
lShbvRwx+QdHsZTgyrce8/CbDzM0GUjd7FeA/rU5MC3pRPTi87ZHe95Zt7F5inM2845kh4M/UJvY
y4zbBtfYpaeJURIaPhkez4RZaDFF/BstNxux4PgytD4rEvxxDLy5od4b+kSRNjWJRBh3XqERiMYb
nT5pLDNeurQpE16QXqDS3ZvP/0CqiIQ7AjxfU4R02SnzcgDhfjav6+6/JfxPKxW1IXX4KhpiGcoL
yagMDGvyplTFzEyPq0bgpdWq5zoGBSEGai35p2mLZ7nvUKSJZOR/2tb0OIII9T/pTH5qi3KZKlF7
gbRXeSRuUum+FPENE3uYbwRgnomlFXlzpZjYLFnorVrjAqkgUGBqbPF4xkdE5gMmkWw+FrHyPiFJ
Z53d7qfQIcZnm2aGuaYOgtqUjIi61QiLPgBmQQOArjiAmRjtMmCnAx+2b5P0XHo24zRtKom4aRL0
UlFpNeGVcHHDVxhuv4R7Ls6G/yfSkh+PP/CTwBoZv4rvb2ltprTa2U5PBRHC3Qi+O/CxSGsx3AdG
ZKzaeJkSqj/d/Sii7I/sN2JrfKr+tvQpY4hC6H3hMxKhbTGooIDsg1/eZzs4y2CQ6MfUozQ/hoHx
0d8NALPwI0KlxufJPIfWm5M4lgbwQX0KmGBZmDTMIw4r4wFZ2WcYF09o6LVVq60oBOSmezCLkLQV
Ri8/VnNwsARyM3+QkW1c0xGo0ZAKms7NpGEIZJP5qybg7FC6luoGN0uquifjZtPcr6m+qH135/ro
rySyYYUuZU5X3KHNhziZQ17AZOKntWNQ6FKhO+h4k/rOOVphk1BYvRypL71ABP4IZT7OokFyxr5p
s+oFAii991JKZjNKcVwx5mCMBlXqXn+DbmLlq+MF+7n0mwy/+0jNzd0rbPbuEX9ogGXNQaYS2pru
0myHQu0bKQdGyCL2fzh2MqGN+9CKtygPDH3lntXwzZ234j7PCJog6DKYofgpaoQ1Po/TQrYX3nD7
gMHwsJjlSQ0DHxbsZVaN7yGbT2Zbxf/9RspwqWBeu2P0XXbCEYGZeBmRnZbvvhH1B/M+ums+wySu
WJamYIuNosC14xOf16sVSF35KGWDovWi1JfXkkqJnPugUmSb40JGu6B8CFv3O/0ySXZGznf7Ykt1
fYYCuAkR2UV9R6w22TWh+Q1Yqnmjq6tl8mDLleGVYyYrDhRSfGoC2AnT795J0KOVMYohvB8b4KqT
349xiJIP+lg1DjzEdprkF/IKSBc5yS22R+U9Z+NAL5me+JtjocTIljZNZktCr5skx71OMYvAHxof
uxs991ajRH6YW7C+QIKFuxFoJicsy+bnthjGPNSeW2gIG0EmNsB93p4l8DUhULNXlv3yifNs0XiW
ByioEcBqbAxH8NchvpYzWvPLutoa44v4y19nVf4ieF3hwmuFW7xhZpMBzLbZUXX1hsIRJL/WJciq
zSu6nciWxa5wzxT4G5uAr5snySbp/e/0r6HomJnFPncNyeA89Jus3tcxyENH9i99wNEZlfOpcZm0
fIKArD7r66BcaSUjomXLQk1HOH9N1R33Q+u3FckHeZyqjtmgpk39T5gNXpLqTHVIWLWCygyFCEjf
4XcK91t481hi3jGIFkxmo1JSArXx7Kf8HYEJUgJLWcq2nokx9iFDekkqeug6GgD1/HAcxpE7amWM
2r+JDp5liAuAxNgzDUGQ94+JuECmUXwWXo1C2g3gx+3lGmbPjSbffaSx9gDVnKoZsP82bZjtmFnB
fFVIUKiR7DvM8WWrHK1xLb0Upa2+cpMjzWpdQsXlyVBi63YH2qGNqaSENmD9HEYT1Hgi/0y+RWLE
zXIi+Lyc6bimKlpoEg+EgSGHMRHs0i/+DGYxFRvBFRemi5tMe7BypAENjvpdxOcjSGGIpAOZE134
dIUGgvmycg5D64/wyQcklZ7V4QAoMifiQoAjm5qPFKKvhz4sc5X08k0pWnY22NgK+v44igX74voE
W9vA76cx/BfESC2WKFzBRg1OvH8ruBal9G/T05JM4lP9LkZ3AcC579XsaXacdMDbbvyiDnr3MNO1
ZSbyQuZNGsDSMz03/+nPeZ9XvsjyTU978EJcvF4mwTBTdaVMOoNjCop2AJbwv+eOehFkbSRvx3Z6
7T2fE0khAi7k2ZAp3ko/Uuf2hycd5d4LUQGnB0fN/TVvmSr81aKay/UiZd8Yexc/L8L2uuMPsPWv
9Bhy2pGK1kaGtks12kEbxi6THQruLeaURuJ4fHzekI1a5EuDXs0FiPRNNZvuoaVf2gcEO8nDdugj
op7yD+DB24oghT/dAQBfK7pWYtH9guWbYOc+b6jBa5z/6L73FD9Yn+y5s7rkqHu+gxp37HTKWUdD
bIJJRoHuqYXoPZpW1eo984hYcsgYZFNyin1UdDgtV6uVI4/Kkrp5XcPCxxLdsCakXutzDEduPPec
HsnIowZ/4sAUCTLPcuOcoPNh+kpCuSC4+oECZncYjQXx/TgEnbxTOrFeUatngj1IU/ojfibGN1vo
NHKIEVo/UIi7WHQHk4hOSkoj1aDDWVZ9hKUwaN/flMObWOuBKx9DEWgDv2QRY9BcM9u6yzr9qpG8
bUImYk/3ES9Do6jiR3uEBco4qX2dOIu+7tVj8pIIh2gkc95HHWh6Ahu7xLoNyg8ixxt+IkVPo1Zn
kGyyB/QH5r1NhxLkd194RHLxU72LoU0Ocg6jAwDudsSI1m7W+3VXnLakhzeJV+EkVxUdXUi/hnNJ
PziNSYpgCrL/hx+0dT0uMLPPoaz9DWKwTarPbCpyboxTKt3KtB3rYtWV38x5H5iAUtCnAbz3EpiO
tRhqL1MpTHH7qrdi4oKKqxsZQAU/0Kn26Dl64WXJ/3yAKwxhmZwKGDCXxLgiQqVaZVvH5toXKVyd
m29xgKJR7hIceLY2CRXzA0K3ONOQUMArsEPhkW5L6tJqy0N3uf1iCs0C3z5pdyYAMIlxsQVNco9b
26SQhycQ/2+K7Jsj64vAuRKQH7R3lVn7DY+ub56FtvXigsgQF2/K797jhRg+9iUSmAP8EopRX3iH
F4pFoWizyDLt/8SFRnbzCyk8ieYWV0bNRoWze6+8sFau5XlCGg8ld8ZgodkZkEx7ZznvmAoTpiDr
VhdLZ7XJ+Apmuh3cP8cEJh9hkFvEg54s4Z5x/EO0hn4HFu7oUy/3McGV8aaYE+CKkhslnfoMjADk
3WKfGaaefzp1yK2Ql9WI6RYM71skvF+z3b+AYI3nny7Z89VeCPPEhEnC/AHWsrrIn/eSkDM3b4BL
kfBWaoCC0FdxOL9ZIyEdipF6+bb05X04amcqRIEY9WhrbhcH/W/20ultkHm2znAWbZ97Y/sBeoWH
MnXPxNQLs1+ESevHQjys8qDY25/sTIVYKJnNNKLplwkEGB0SUPpkf2MIY/rx+Te5Ferk67IK0ROA
r4XEgDe4G5TiuqSbxggSFFw2REPdkHizyt8VsTjTx68RaLCCNIAPQHTJ/d6Iwpy63VK5YvWQfPFn
ENGy3fgvefRD0dAHbM6Hmoz38h8ur3c6xp+aRG2kqLHqniomcqKEyNCHSufNoSl/LG68WS7eCvYI
pZ+oVMftAJySUXpbjpNsxHwCld+IIED5H/YJKhopcY198pZLK59UZsQLswTN2xTevGA/IKsm122+
40rNGN7s0E8NqE2NRDWAbyFtZ5oFjMI7R3gWP/CE1uLbgaN9YTF2ghrpTZUsKjDE1ew9P9LuQZP9
izGn3tSHrm+CP88gqVf3yfNLrMNPegF8phTmngwQj0FZic3kwSKz3q8REvWezpGYDa6SI+QfDE7o
XXe1PjyVaUwrOISjwiAfv7K4gw1B/1tXMgnuB4+D7CziZoYGQGZNkUan6Yq48TftPR03rCH35qT0
ybHFojvlsoYH1hCXT3AHZBkyo2XEpvDD9u9KwtllCjD9/xz+KsSl5JjbEupBBVNBCU6rIWvzz27c
JVEd/HZYcNJI2w+JxXhP6xELYYqU7ameMWlbOqnlX5VhP6/wBrRByw/l9wweHadfAaz5Fdq0sKCq
5cPIQ4NE/JMXnCC6mnjubWLT/iBNIZxqKCfH7egMqCfV7kvgQQ3ES6KrMgCL4t60VcTeHxcAFFUv
j5Yj6IK/pv5X3Vlp4wInEEfHqVjWK/DZ3OkVlSdS0tD1lgv/2b3bQu7MHPiXJYnGAdRcHQZF0hLg
SUk0mEhhN9XeOQDiF859AATE+I3lwniu4bh6/X9RpwVQqP5DAagl0bH6iI5w79Yws6uW4oHLajxt
mYEr+4Q6pcJ0WarM5U2ZZm/DTdcHJswYvl2oc/+MY6yEv5p0GhqF4Pbwgu2Gx9fJVrWKj/y5dyTD
hkMx/h+WHvUDfr1EVTiwEsxpAXS3OJQyCjClXzdNHC/3YRHPHqnxh6DH+zXsGVp36UFO8FYxa9mh
ClsZh1WF42ctMVNySPWrNrEaaGVGFcohUYlC+cIE/R3yTRg0s3exiT8FNp2qOJvKtr6kCE1+preG
+dpwFwhAgbULXnbqfmvjtZQORhr/TxINrVNrFtqOuqr4cHhHG74WIsGE+ZGim9r8OwwEJcuptdFR
kyY+LqS2OX3Y9Mqn0VCjFNA8rdc+SNmcoAQSTx0G+cO8XZmoXQUfGrguYE6GbNMtFx6SQrJafPKC
nno+M7IwZqesJBobUHDpueNofxKtQUJYOUIY0ho29E7gDGq/O0Gw+gQiZjejeTkr2lzC79jK5Qyp
nzbzFbiBwroMARK0CuX6KR/T87Xcclkh9tVJI3bLGDomFNqHL8u+rK+rmKULF00hdbPjAoWzsBRi
2v/UWQr+BLWGDKuJJ/Je3prulQaeCkbtsXlkC20sUPzOdVvixDVFZp562BHbpf+afMJ8LyRKLM3Q
0z6beOcs8GFRSX0Id3eg9ONUVy0lpKZaKUotZ+u4VI3/I3ZPaFxbMC+gyMfEjv9kpjnVR8OWsAQX
YL/q23IWlFXsFkvP+xJS8aXEbR9FyrEZGGso/ylhXvuzaeFLOs3VFVvl1coE/fSqKAH2c64sN853
wXOo0TJW3tRFR8DGl25zMsmuw1aI2OSGIAvgkKcfcdH0/18kNnmZ2stmTDflIyNBYv/H7+VPgBFb
YMbOWcXr3MwkVh7uV3gDYe7/SHqsPyuBaBUzrrW4I7jYitS2l0dtw94u78WXTe2k4MKF6t/MIsLU
2B3CdcQNiSW5OxM/aNSF2VFtqNuNJ3l8jiVBiLMR2UmItZoWhkLBejdWDtSV4RoxINgf/7jdIoZk
/tALUOuUMOnA1aN+0pgW1poCfABX2ozEpzUkIL9nC8od5KRSr2TOmO0ulHMgyxWhtVkHnyZJf4V2
jxPlsM8prP5+H5sPUjQqcRkD6WYXuzkPSwU+fzrgbAfnBeBE/g6m8uSO3M+1Fe+qYf+p6L+HsXqN
tgmAh0GFDwJTbynKB4/FyNk1DfbugWyqSusbsbzITYkrbyE3rOv+5YGt278eJNjVs2vV+xJb3iaw
awto8mzCnwr25cNcTdl2eiNNmLIPHU6qAIymZwIesyncD8CiUvuyi9lRCFGtuyTAOUH6Lqya0CGo
w26mltYBUwA8IK6C2cbVqobbfFY2nczpyVYF2s9NZB0vdlehnhn5XlCFVaqWMYS9a39gGc/Rb7iI
epCBFquNbzzenH6bSrsbQWmYF9pR6pR843Z5k1iWErD/dXS0ulWdesv55lFY/by2RdarGczCAiXW
x+idB5Wn/ZD5AlrD7Eo3QAHj7ETGaR8oa/G5/tKXHv7UT0hPbkpV3gjc31lNIMaKwqrwjJpPRqSP
ighld/4A3Y32zW5mVmgNEWyVQnXUEV/8KWmfNme3vlym0uY7ZoFEAbw8r7EVAaWwiy5qawuMd3of
ozBfQjZICS+Udhap7vUt1lbsluBmhEtaTd+5cDInQwKGoS6tFJbL01oY9iyEbehO+vAPSnQ0aOmg
+a+aGJi8SLDh5NSV1Mo0qDP2rjYGtXKuQOqoIBy8v4qRg5+HY5fsyvPlTmiNDjkczZ1W5i5TSKQd
iKhwoysnSPk/HG2KdvXfmaTzXfuU+XK8m73K6p2rLz35VGV0wOnjFp0kUN9XXj85LFcVPO05ZvCX
KlWA1u51xEPd6a/sjUpOWv6HDX8ZglnvLhopDF8xvhu72Zk2FTLiQ/gTA4lWhO/rvHMAXfRf6h6w
B6ajhTJSVq+VGEP+1dE82akJeJORSYidd1BSdqJ2XDmbQVIEf/Hy8O7xWBUgeyhKNhvuRp9TpCkD
liKshUqOCXgcz+O/gZpINdDSgqn27cjb5XSZgrk87mWBayf9KYMPOTK7sRJxH61KY/G759WxzyJc
K5O+Jy/NO+Ki5mnugZ9dwt1c92ccH0aLDpKpmmdU9kH91bvOxBj/DSncYOYJ/+ChSi441+p3qYMn
W93zxrsA1NXRO2Q8ZhkPl1Cnnzj9cnbzfb2BqxL4iNR6fWlQvu7rkMeFimKtxA6064iZ3VO42tI4
3k+O20dftnHJKHdEsZxLi27Yrkq8HCD2MZYU9ttTTqyTIE1Kkx8DO9VpbCu9R2UsRtZtOJM0pZDl
2r9FhG7ub/aHcaCNEEWYk6d7dTBI1GP4tnW4vxYz8gBmKvJsWAOWoyg9Uxvptj1Xlp1aQxkSj0hj
faAD18S6NGKotMVRU5IkZiSqS2I9Yi7X1neF1oupWLtc+nxdbdofDofAnN0g24Q7nCYOEAvT53gZ
eTePlU+TjmX+bWYqvtsm5HF66ysgfivfNSSkexNW0qa7d6aUICNvYretMymZaWXw2sS8sGucCkAc
t09IOBoN62kw4ehAV0ldXTUCAWWzBMg4pZgKMUBIBaXZqw3w27EtNGQaPkFGgGyOOM/6nP5qIM7D
66uJvXdWijhG2w9AQ5CcZmlZ4misihkkrcK45ITXdmht8BOT4uNv6SYAqDZP2Xbmg76SOKYf7zLL
EZvyJPsgIpow26YhP7le9ONj79c++gnR526p8Gpy9+KhKZDOZw1HueUmD5AB554Bze00a74Fo5eF
pD4OKCx5MpAYrbkWVAHrplVNCVlau5Mo8lghFO7cmsJg9x79NOUF1qMULlBG7jtUtssKR1tor+P3
dND9XPWxTdFQsidBnWUkPB0osPhTqCp+UV9kzCyUbyylYYOi7mFUEI4q7sg0VIjF59aIKFSjTnJM
CfVRDgLxvKQsJ8qd8F3qel/7Asa/AS886gAGmajH92HuP3nsyCefvOh0UJHAScOGQfteeknZluMJ
R8IeE7VgeAkHqVNSSkOmXIeqacnJm3ZzpsW2StWSkSKOr7C70nLMGXAH97FZY14aDVrZwP4ob5ff
eDpXC9+GKiPxJfR3Pe+i6u7Pe4zXXZ4bPyAT59cb4e54qR+suHvDNHZZUxG511+RVZs0klTIjiMJ
yl+aQ2Ek9t0pGkMWcplsAcX/C2GktcRnQ4GA6R8/w8/ZYczXCFbXEwuOh9ALwW0AtKgdEEonqL1g
0UunktUL8wQORhMiIXvMJDc7O6G5zvQrRvPaml+sU5M293zKwlwprMbZ5vnHb/6uX3xi5l3CW5u4
EaK7hQfmBD+xEWEzoLx14+0E7OQHWqoYtRBvmCyB12hRoiNNSdud90ox0p3qd7M+PhuK+09kUN30
fkDB7ezmIlwoT6zUqnGVze/BwwRjKTuzEH7YHIYLF1sFYVEwH4hTKIsSsFjqMW5yP59Wd9dt1GWP
68TLghJu/krQI2Xo5P9Edp81lIYXi3piZ3KwxAaePf/zv8aPNgTddCZjVsHpAXE7OGd2m7KOIROO
Daon1SK4tcg/x1mvU46ICfFHzLbAygrhxaOZ/+4zkuTKTuMqwDZRdiQ/DJS7H++cOJRVwXs5ykKi
+jJ/0oxxpFiPPkYfOErWYiAIkhvzfJywmIPVAA3Z4QWtiZ+7bsq+eztQiNTTRvku1dddZw0iSoBJ
q+tzZsU1ItPPC8kn90H6oDk38L+V2aFTKW5JeUYrXd/OkoNFsM5SueBWjGw25xpomv2Of7oXl5Ow
mufVgivqsp25Kqtwr08m8juPYxcTkeBlg2WLS31nvLW4j5Jurv95cEsE1KbzI4SePfCoi6XTJkAL
xCkQAY8J23j9KKBSi1m+3ycJdezDGpADX7s162CacceVfGyIJkRFPulMC+Xvu8lJxrTHu61WMxgq
+90pB6NxUENzRvpCm4qzOVAH7Xy/M52WnL/ae4McIL4WouorT3P8BUfIqeYao8oy5kCNxlOf4wT5
Kd35oWgPFrGF59EiUuXxLQ6TZZ+JhrgkRY8TA8BUGQ4FyrDqpPyPcsmHdCEGVk9o9Zr4QXxd14sq
DJx5WVPUfhfk7Skq1KFOWjGzvrMoveGuCSGq/WNu3Oz9XGh1A27oLOJI1lJO4eHdJlSxy8slRfFk
FB7zdmUkA72/CMz7Q3dxQ6PMm49pxTTTzKnn2G8kfpbtS/D6a04w9QuUbzs/38E6MC3kiCXz98mC
FsQRmV2wSTGdzk8OzSdGol6zdwQHNTpDOVHwmyrDBhVONpJIEyx7lMDgqf75lTB3/77p0Osf23M0
erKUc8IHTivl0N46+8KREPRmTWZqSbcLwmm62RHn03cmJ64rZvbBQhNe0pLycwlFkMwme/0heEao
q0j7LEVxgUeGRIIfaKiGz8mSgu7nTX/FftMikUN076QpH+X7xVXHF92IUr+wtePvLOWGL6u1bW8Q
hmb+ZXlE/6r+xV7DsqowHe/uxlUjTDJ7VMMg0w+bfz7DYXaJl67aRY5kuG8VE+b+WtjeEB//U0Bu
/+8Ad3mb1KlTMPPCfMsnV+b9IaPjJBSc2hONIxRz9Fr4FzFu1j1aK2/sw/eDqX1rxsi+wBj6mY2i
8YDX5G0Uh3TF9In+bApnWCixa0TcWDi84+NsR6sVybs405kKxBN0e42GPttvcz12JScZfZP9iaXT
SqAlhwAc0b+Fbx4748cl48unBSvTktmpHd4HNbZM7XyeetlMeIrDCqfwMfId9orD3R+uYGirI/3l
3L+yRgEuhtw4P127Bj8CgXwCm5dSP5mV8bwpRGYlSyolHMEXCRp1bCrU63qv4GkDYMYFVrFgssIu
4yeUK/lTa4i6V7xJW1Kq7SWistJSdAZUK1mHpU7jb1qOxNY6OSeXFhlDiuWl8NJGy/a3bzm55TJL
m2sPHNjM+tcLoaK9zLYw3YcUtLk6TTsUx1baRyFbUnZ6QTOxaAdA+shDe/c7bt+GbqgXzFW2wDZ6
+zaCYiOVMdH5S/f/XChE7X4p38ezUYV4ntc+H6aQsg0bnZxkvplgqQtZ39qr8HAgvX3eCO1P0Lmi
gEeUCZb/jmn6v/jTt8mdrjkFywTjArMWwFa6s/ERr+MAN7Y2kQsplILfyJoVDCTBuII8C0+Rs5pU
9HKT6q59Pv/xU0bIuuuP6PVZDAjXJ4bFAfRpaCITVDUm1c/hrjP8vRZ8uO5/QtquF9tVwNoa/yoT
6sYLeFO4pyffmtvrKLil1tRdO6F7ihKYM+bi/Hdie+7vvXPbR2x8+4RPJxkbfqcRstwcizb5zee4
YBPJv5M+2hjPD4xhmQOT1MMq/cSx1rhVSGWrtmr84qpL/f5yfy11IHfHq/wtzysVNSbfvE+SvisS
DGVlk1IL0DD6If4Hs1oyaodeOR99Ejn79dnR2/K/tYEQBNnUnTiHlOYKXaziofUN0zcjhlP5NT4d
jKxW3SMF+qzzUDCCrOueggH2EVoQPJ6LzZXrWG71XFx+R9Ss/FDkLPJRV2mpgWHsOI9+TCMZ+23u
sg5mzdOL7+5jtmB0YCtcafJiZCUFsbeDkuY9FZGCXXaNEVCJDYmxt8qb+hE33JLiWoYI0FdiP3nQ
G3KUlKtinJ07ljrUwtqv5Iii3tjyuHcU2YgvWVUuchqjUhIrTaTWhobf87jy7TI+aps/Hktc8YiF
yI5YOCIk6vKr6OE4Vfdse5Ro5Txk16t4R9/QnMQI5ALJ80PrEq0ERUI0hf8H10ZbYN/5TkdT5Jxh
ua3wKC1ff+iut8x47AZlnt/3N41VIEoPcHOOtaaJdXJMramhDTp0cREsf5InD6LGOlT1maKITSKQ
pZnN1HikrBWPiOnKbfwH/PJ5C1+PAg5OKoARhTYWYxzfR7V+Bhl+AU73mg8X85W7147ZSIwDYNEf
RliGnE6MJ8yR6/dofuA0xmwg0pg+Pk8vcT4meJbP6at6RDjy6EEtopCD4vHt0mYSjFkhPfmq9EVh
iUjn9+Z4GplNJn6nWn4qia5K/W2ZGsdvOwx9tNvd8z3pItWGVJO04sKgu8mXq6GlTMd9naV9iCyU
iKPB/y7CO9GGrebRcoEOFGEi5vKeWAvNoRliGjfoKe5Vf9vW3V61VhsySfvF6NvRhvQ9THDHv7IE
okEv8DsFYu5DvBF4Yk7nBUFOgHa+P1laBCbSRAzNa6ocFa85u9JR/QzmPKX+gs4xfA6MZZA9sLml
DsQfQNQYq4sAThWGDqjwblO6DJy16FQ45rVCbyyrhYU5dFVrEXbvgsHm4i1O+EYsIxcNNrGSzBuy
8LWulTST7AxzA7oaaQmK1COvUk0U+0kErQw2N2gzvYp3go+ZjH+xXoMEhOLpVfJPLdSBT5DcX+OL
lz+v4qr6+crcPMjaBgDhl4jPGI5XwSCu/Y1esdfG5AzdA+y0I1wSLjRHJg13/DjxtkhnNG/jpKgy
jmw1ZjipAb/EmvN44xn4kaJuigJXNi674lghUkxla+0mrV0jWqith+qavpr4v7CJlGccSsWgri18
pXEjMM3rQMMxvIA2NYExHJPfR+sUIKUFTP18z4rj9MuVMiFhY5c7A0RPOZhW491PGSNCu03/gLpd
Awio5wtHLdVyr26tnjRsbBDfXChxBSrbKIVRDgGgzGcAwEWWETFnqJ209fGVjRzqCo4PJtjBzhUU
hlTni9JyVz2aex+7Tc1Tzui3n8zTQH7BMit5+1+33yZ+sumdjAxipEcdmQWFsSV8GM6X6PcxcVh0
dxV0bEP5vMxU/tSj1TvryTaVXi6cj1lPbB7iWxTfmbm64WVTJvcV1vc0mQmVc4b0nu/srdl/eBgF
aPnZ7Jfqo6n2szydYz8KZUg0FJcDM24BBvghcYwBd6b32A6YWfkPIzPJGvjTU9KSd+0tzmyA+qUM
U/YmBm8Q7VA3jGYgv01NponM1/8y64XDYABLIBoRX2T2k9go8kiLChITmQFdU7K7z2DaoGek42wv
YnKcdin3/258cprnSQoRaxmS9PUnhe3+1qHalbFAPV9hot6ULMQLQ2xZryPYlgnDKZBxYfxsk/uw
pkWCVuuVMjP0aY+1WbOpMVcvXtFL/6y3Ifrh23GH/5Nd7qiS3TPBvUQ72QuY3HfQ2F/uyhjSsZg3
5MTgnUbpoIlrEEDXIIno4fPsJRNRPioLIHmApy+6fx0kq+cA0iHN+soXtIwU95fzFpNBsiH5BkkF
BGjOOb5omCicSdYWl41yFQON/7nWcHCFWDY+4PcYSwr+sgJ0pvwCVS08JWq4S9cm5RVzgZrjJxiu
9cXYk40ECMC16P5aIpIe/fAhUQh6rAgbOZgHorn5joavy9ulR4Bo7ErIk4Y24IFon7BI5DJXg82z
R02SkvX7pJOU/3SbIaE9oEMxUTULi1mkIn8KvoW3gIeflnEVCqFD47nDej8BP/AiMMS0CbRI+R7m
ZRkilvg17hpDbWiOC5IjKPwsPkWWT3ZuO2IvUPyPQhhPcvMJKk89whZ8drv/0hn8e20/mdDlpL5L
pIiBZAxVVDMYlC1vwg1ElAmtzmyIA5sV/0/DiQJeBQ0SMDUYBnci/79N4JBjbR0aNXGDB1kvgVGn
w3N+a81yozUWFjmgbF14onBwMiMTmIopyUMfdk+kYMlUNpvifIYt9Ce4Z9gAtEuGa3FUsh5r/nQf
qG6jpRBPT35yc4I7/fGtZEORZuoDlSGDiLL61FATS0cH4LmaAl0qAahjemrIPEhiPIwgsZXZElLV
QtyQ8qk4mRKfjCHKLv6dQ6u1Y7i7LUYEe7jlvTNexKWQjrPLtlJbO4hZwgNc+/g81mY3u9/mVlzE
kWGay+8mUpdlsdTfwTgDoOKT4uM7MfMLrvxvRMzbW2IM4ELUCP+FPQrhTQwOhRIvzUX3+lGmYV/Q
P0xKkECZbCwo8F4FmUD8Vm/RkM8Azups1Vdpy03BbKCPKI2vjwu//kwXWyPyvnVjmH0XpebcO8zV
wCEKvyTW9/ixRr29wgy923ItjD9BEw0w9Lq5gZD5ebUgMsfMgxylPAMoiUcdjiuSH7+R3++w5dZU
mXiDRpfsEU90K5njPDyrZ1ANPrijx0VlZYDvkQt5Z9ktFEF5SuSzm2vkA9kMgfZDRrZ6Gh7uCtem
SKMT0N+t/w2l4f9YzXihkDiPrhx6Y+rIA3LG0oTSDU+ghS5wQbZQPh4rWVRYuteqd+C90/c/9pTT
HajvysNoHkxp+VoXzY0LeQr+9BlQIB3B7focLWbrzXmSj//+4b5q8g5rQyzWu9HtJnf6agj1zapJ
XcfbZyMosBJA0FNJXsyhumDDOqCyqzRJFrXLXA6OhJ9w+evH5ZjPXa6OowHBf3gVeYuWajj8wX6v
AUxp1vgVTbV82CAei/h/QRKoF/DZc0WSzkkfrEEsOQXjJ2Gm9ANYOSdsNSrVYx5AI/2q9RKyEyWO
msdDXT84J+4he6IwZPZiyg45REOuOBvMX73AGcvOZGa2dTvWWTLjsVj+w9akqIJ/gBbr6HUwd6Fc
ZplyxkqwwJqcZlgxHSwbaVAvIx6+VVTC5Ax2d8NkMTFbucicBXjNsre9TuUbVPkkoGhUIp2QbGbv
0uyFnqKZRAcJqkMdhCEV3TQRtucJYPNlBPzsEgnLXrb3iJG7Hfkg+B/flDVl2ugQ3j+O+hSVF2PG
oCq0wvDT0KhmP5O/7uISDXY2T8HKLI8Mojb3fs5+Ml9r3l/Kv3RBNFnFzrK3S5s0TaAYd2GGfgcj
lgUpAKhw8MmjpbIPB8QpZoHAElikZm17SHh9eNX3MOcz09bZxkZyHno0aQIw9ANNs9pCt+9PL+I9
dtErHfAgkjsKq45hyxS66BbZWDotoP9/WEvOKyTsOZv0rhDUkQlYJhhXGbb6u3fucl8h/c+Qk5L8
fYys2VzvjOOLVxcLOT6p/V/kX90qVECAy7KFqYF8w+dU63TBE8RTnv/+aieXkuZh5PwbXt9nve3y
BbsFvaoqnWCUM9Lb+Efghyx5vuNt115E5/sGLjDsF1RxLUb1IbwhSx1IVl7AJNzakTrvA+65SAue
vHfSHEEh8DKXC0K+4X9SNKr8stygq++yVuNFTc3cLiCvOV6oBX6ilITDFXg3iPHU5IJsxdmPcDBU
W7uWe9RzbfdOsz/Xr4Yl2ICTsFZ4QijJjIF2E8/OxZe5juOJtfppfHzsumaBPnp4Ob9GdQRkyaCP
QL6P7/mj+PerxTScq/wxn5fSSmCA+RnZbzAJ3SlInJ8i518zAu052A/HbqtGNiIdbwEdvw66jDz9
CNg0M2LiAjTfqvON+0m5FcqN7T5TYJilIjygOaN71DsVQMGuo8is4zg22zt3Ez8aT7dVIYEsAH6z
CyqvDHjbN0bXvL00g0f9ZmllS/Wr1pJfC9rALagxIPJnhM6HVbQCQSGg51zy2Qmu4kdhOwaX960b
AwGGRZ2TtxHdf1sxPx13Tv0Otmm5JM/0atKBFYfBl5bDdWIidfbGzAbu+4HVMOd4USk6U3IHoZOi
zAlF344HHvVy5QTaXeqme3JWxmYsRqJgfq9MCgPhnx0Q2io1Ya+linLyOqU8k9HRPDt8LHhccHnJ
HJlsrGt8vPCCh2j3BEcZZUK1VY+nn0adFsiIwpY4uMbxZmiptxmXPqEbf7UH8v2Nqunljzu6QjJ1
/H2Owu7DOVq7rndjoM35VxvgPqmXgeTXVuFnQPVGaTZ08AOGJDywEp0C6EDBUDRJwNxEk1SwZ9gD
jL/vfOI7aLJwDBpEmGaIAMPcQLX/kBrvzvXvc6DpyRNrr96y8sxzKP3Bpd+/3Od2RIzoU2PwDjca
IDOo+CjruA7bAbOQCl9BaGrK3SQaJHX6seUJE9B6bgrigjlw/Ig3f+zN/dr8ms4trRPuW/fRuVBq
4tHuCEBkwCX/MTdM8XE/q7vy/o6+kynJ1ZMio3Bn9IwEQpFI3HWZCOhv/C8U85DqR+PEuuvmvRS3
c1fMkL7lDAi9Hyz1vQ7W7ZDhQHixo+MwGkxAX//VJSq1QD9VN5TNevWCpOdKK5MBCTvPcLYwqKtA
+WWAIdp/LBkTTf26PzI+jzPYbo63d3s8e9YTiGh79ivCOzUqPDgazcAhKy9ifLE+hC8kAJiQy25r
G+Ng9Ot+YAn6ZXWy73gS4kLBnanjdL/dntbQwwng+WE6DWeW2KPc4ycd2Y2siSyjxn757gaaJypV
3MmhnxbZ6x/Equam0WwajoicqEnRXk56LC00pSfeI2ulGzLbRbe07iVvWR5RxOuw7V8c9WRc9scY
BzCgXtB2wpecRcxD+7Kt3XL31dG40mZXCKsC348xUlKobdGANuUL3qWIVRlvI1SoVy/pPkQonjNz
uqZJi4FgShRZ0q2RCoRYWYdwr74MuxPw5IwnvVO+swSQ7IT+2341zTJ+/QNyZaKyQh+I5XUaNGWl
i5emon0L+dbO6PP2C0elJ9E2zNNb3uazWecxsRkYDKa1ySg/o2sQaboRd0EqQ4QZO8pDdAiYAtv7
TNQz7OG0rZ3eZHS79gvGM6Hpm31cP4196UmwLYvQHM1cf+EGzfjRcONpobjixRDNCRx/AGElGwV/
78tqQRjxJhhckacTUQR97TfVpnnkulYw9MYz8UHwctXLf0FL9iMk5n7fnY5WYK8RO8tU2IDDTQSM
R98uCbLu8suwdxZRG77wfiF9hFi5M/Qt0P67uM/Cr7iiN3foyc26CVRnYf47+6Kz4FQ07Vcnz265
PvWWsFZF4xPvfW5ggZsJ/HNwOjLFhKD9OGr1alcJ1ymiWbG18US0ZpjPHekdZIQWf6mjpz62Q4eL
0bCevtFk6KLvCUPnm1gNb7+jysvK9A0LDZkLOJ6ppooIf7LsZPBXF/ZgvA2tV4knxWw2TpiAdp3C
CO7aVsL6q7ocy6lRg79n8kuxDrWFYLXTUoTyf1Vbw+iYnyEadp+knXn8FjGpTdyWd2deL5JIhRcZ
+MuJUADvHlzACsBNzoYvfmQy9zzlaQJwuvVkLv4Bg4Nu8H+8eD7QWvPNRYoLSWJ6NwuYFw5EQ+Oc
mDUllfzxp/TeY8iy4OEsZPyr6Qdvc/R4TUvKQlnjeUQMlAvk7m2V4a8PaBWmk1sBMppTqJNHD9In
1BKOCCxziA01S4lwubF4j7ZxM8xaCpduSMdGd9Tec8ulN51r8SoUhjSgfe++b8nsNwLAAQUysrJ1
NWccD0H22yg0f5m0TNtcC9spownGqap8ddugimLCsJok1Mfn4rt5/Igh4yqANzYpbb0liM3OetfK
r4TydnOIgRf149KKeBReuQhphct6YjylaHO1taOR11KWTm8RvL8zf/Gr3E23WwOBfF+2aZBdHSzf
hWQgw9aA/nklF9krs0AONnKurkErikMwaaj9+H97ZmEgnUA9K5deiHfnd5oBky2Pr1NNwBXMGLuZ
kr6SXt3z7aB3aKVLKyTqNGiCXV4JLK8J0ygfAXFUqVd85gJSxqo4pD3kx9dl7DdAVxrOpRQbBmwI
06281RPnHznv7NKZA+bfov+T3uT1Hk4q8QJ0il6w0YqxMW1MC0WYfrm45GggkTMxINJtY5sgmvcW
Jd+LSP8pxE9Ojb8QkcJOmoC+6rINXeKhg5y5OYB3g5nTnH/HQKMsih00w6HfEVzHPMXeXe0GZGWW
q7pNib6SuIzIpcMFLf/RdvnavUN70ZKz+YFctDfBOCLg438/yMo9jdBUH8ZtoBgesLSuDd0l2k46
mWr4rIVXTHmLh2NT+MqIeGTI4+cTRshYwGrej8VpYGE1aZzvz4/udiKDJmu+Iz/piN5XzeeetnGP
5QfbsoCURm4yOaRpMlZCJBoXRxHujzXZqN8wHbOgidcOjbUJBaKFlBDau34HEFOPoE942phNI/B5
yMAlQbkl1cqZZjMND2eD1t30lLF1tmV6AXm1lK9cTSN57jgtXnrniiAqV5dAhul45aNBJRvJaEKx
aUp5dSI9G0SzZfffXsYQKQJjt8bVFiDuJkQU6uApJA9HFVyyuwOhgMm+f4Pb+5+NU+bkUUHZB6AL
jG93tLCTuquamxHdkYEatMdAoS/vsNs3mqB7f2EEV3mcRFSiNUQT8T/7Rnb8pUtjTLUc7uSTrUjT
UTx2QwGm4h7tGkUloJF1Wu8mqXHLpt76f110Z+ANRECK+TrjcYtFCVch6Qeo4SVMFSLC1m7X2xoN
8QDxFxdG4pei6N3xvLJy4/hW/ej42sQSOtwaaGxameSYbizdL6VOnoyfNtMy5KHnk9O5b9BYiSmc
YohXiaXhj3xDTY4b3ujROLyls62POUbmqqvr+hfWdScm6js+zp7K0QnAGFMJj5zCoSSkoleYV1Uh
exrfXgEVBSkEck2hRz1LL5Nap392zVIodU5W2Z7xnatLTHJikvuUxLhyY3nw4WtaQmy4O/Q4MQ/6
jHvzJQAmmvDv+VO2OzpnX/FeXl3sAqNEV4lHj+GHzQT60rWafpBxnv/AWnX0SxlM1cyRQHma/aWs
I3N8QgK2fsxEBaWMtveAPGH5gmpMr6mk7FGtH4LrIV25rSK6bVOskNaNHxj5aldHEtrJ/dV9CJSM
lrBAQ3WgPs3wyGXt0J58VlXjFKI4famTlKZZ7ZdSDIC5re7enUsQ410SSiErNrdCLAGIVeMlZt5c
AI5wJ8gFJnj0A08rF5715ydQIRf+/9A2DwM3e+SxKFCkY1IExxRCEyI3GfX5PfrwRSXttxLzfHOo
h28Iwm9SMw85guOpFPEhigyoa4MXhhOFy0h+5F8ssFfYUJXzgm66mN20n99txgH722OG8TYEERal
H3V6KOlIziRNlVU95Od+OSMv4fwx477rm0T8LM4sS/zTjDJmyy9jIT49emFnq7/zx/WCzUK2GpZe
HJ9V+c4ysuiwEcjpVN7ppfnyqPHewNa+P4Kp1O9R/2M1sXxQJUWloYldq1rqB4nD+xqP8ICCYJ6y
HnvS7Xn58pECJEv7Eti6/bGBTMDfRapu0tEL5jPoQg6hK/liH0xtRckky/y/N1zyllNY3b+5HRFp
48ZPWV1DjIq3DcVR03I4Q3XuXyf2gdLTlCLQnIGbRS4myu9ZH6aHt0yaduObCSsdFW6lsZLW0IVH
EvD9dqa+KCJs1XgWXaldLzp5XrGqUApJ6FzPgshgQS6uyJjbN3kRC6Sm7CgwJAaWrdfb3fZKXWz9
WI/PjFZJCmqebwOZQ937zASKzQJbaGlwlIQHPWdQ30qgT7aXVjUTrGx/UVFRx1BCSfmEIWB5eWlm
EqL9JLEOBm8Fq1NzX9UfSfb806pXdp5GnEyCdrp8DfYdnJ1aBccXgnWQHNt4mohIZkQMVZorTwq6
ix5KxnXHRaBtiJ4hh2iaTz7SOMpeKHc/ACA8DNOJurXlWG8sIkw/UPxZ4wVjSiWtS8kh8nJ0qCk5
9xnbxi9tw9Smvs8psdD99+WfV3bl+F/6FCx/yDmf0OPq3Z5rnTloupdr2YnK7d+uDWAW5c00qpek
HDflmsbpDJ5pCqhzv3YiZz30Lwsk/wsSi+TfXapYE35aONlvCFoy4QWDSFQ0lPdZGm4hKkQyvkWy
OFGwTk2GrjbZEfjPm008m+vByRdES5BLHKBxAqezpQk95GZAe40g5jWsUxi+cdAYe9pvI971Z9Ol
Bm2qHyKpY2FliFQ2tFsHQ4fxb0xGxQEpIK2T6LAMbD1Jsma2JdKOoiHEbTqXc1E6vwgUMhjkRnND
1R6tiO5/w6Q4G4E/pCf01a6yE75bVlKuVhsMtvPCg5Ss1CGFt0tUyjTHP9IRaZBehiuUPzW1O9Y/
CUse6uwfWIiJPk7Fgeo2ddotndxvc0G7bRQI1FFsC3tUaKADtSZhBxdNk2bMAFbKwkge6p7O90Ei
YMDsZd/+eveplmM/Yu9h5y+PLvixOlU1iFVaThVU3wWeN3/4SvbB8+iZWyU5zuL7qBQz8gLPMuw4
S2tn9mfb2LAFiEVzrko7cDybJ+5l+D+xJehrRjjzAW710PJbtHoKDUIwXxFE8ih/NQQoYBWtJLI/
KYUJQFi0rul/beTDi3YCMcL9RUgGlRExu3CvYp6e1E6QqGu6i+Adrd64d3UqB1wHg6zT4oVosZi/
CvLk+bKfpO+hwGBCaNw8SwL1XAahZTBhDChIQA4kQnkJJ4AR7IKrpPyItr8GgT7e2RsVE6WFDE+U
xM3Vgjk+QRxKwYb3i3KYYG+oVbd6DrJVgG/EM8Cyx/Mnt6+XiR+rsZKEIpa3vqrsKV7gtseUxBuJ
iWbvuTw8EUbIfZ4it7r5S9u30ww4k6kOgR7P4a2CKWH8BpWEUoolxoJrVKbRumgKilJnOffV6dJF
hN859Qr8v/jtrewKxc4sxKkzICJNxxtXwpTb+jy7+Z6ZNt+F2G4FebLFXi++1U8x7ajQYfPWcZhK
OMEGDwIADoa7LozkKz5ywBbyKFA6GavwdvHTNuCMpAP3imE0P77jCG3/crDj3wxl0Mb5s1/QkMi+
M8ILCZssQQbnuig5vq4H1KCFzYfFQ6Dypoh2mIisN065+OnQEDQwMF2hVXRPXmN9DIpJNcmUJRNZ
7CBMJ6dR9+/q+7s8FOtKUlsfasqxpoohzkcxsZXS48zTMy/0r7bz9uGAXMfypeQYXXqXHxJ3yV9X
uYxWIAm30GWUq7KZVfxyYVssNvoZsAHmy6MsBGdiN8mDlxtvJ6QpnvXRcvU68wm1Y8u2jWZBeKsa
xDkSVYd0VKFlmxk7lhG15Mnhkczk5ZrGzk0aO/VmVTKhaPg6UPplwIP1B7Vy+iBd6qZe2n93c9lB
C3t/3JbHKjsPaL4wNnBWxPmYfnn/BcM1tPX3DYhbE1Vcaq/o6t0TjKLseMic60VMSeRWdpXwkXnb
AkptvHvi1wQV02WLsq9edHaDJj/uwE1GwgDLjP1i/95rX25xgX/v1fQlSptsfXXD50MrGpvdBBGD
a0cSjOfe+7qk4wj7x6Pd+ZnGo2PpD4Dc5gCzxZzCbKowF4C/R4oyQZUu/dQJd7AqcWJHE7nLfteb
bJcqUkJWm0ZPXNPpM0J7TCWLKf9LIb+dBcdv1GVpzWd+TpEbKHGHYWmW316eLXhOEHpn9s06qfp4
qXyLdakM89zoD2Xx896Xs+fEuT+dxgHREhc4OH6UNi38nfSd1c4S//ffIN0+Be0LPdkiGgKA3Dsd
1JCJgvKcPnpZZgZiTdvSYo09UmhMva7iAZBLl6BlRjNAuICPX5IRwlwi3GeIAqj+zZNGw1fGlPaH
GfCO10m1ja/rWqt2rpQ6EbOn9mmUeYvcdaY8+xLZEMM9u3FOfoKPOOcFnu1SAnf9UxqZIxcQVLF2
+9tHEp4Hx238flNVQxPNzpAeUNIU8rub8ITAtkye3aC65TdI6nDMe1Z7xFhFfoYZ1I0jAdcFGum+
Ol0dtkvJ2wq/iHNXzYkHSov8XuOq4GzcjzKesEYm+gtkf4AQo2TdGrXxAnEh9tl1sGvXBymL0EyS
vOlBrxyn2mO9l2NzvpaYsNxlxwwmiawT6t7SS3sAhGETfIqFi/jp13MTdkwB/2jpmjsqA+1AAdgN
sotWj9qVbFSkkruyaB0ZZNNSVO5qceRnFod/L0jT4iyBQEYBk2U34GT02xv6kJ33y6tdbqL4Tueo
EZ7OgYWZXIZitsSu7ZJjPgNjv8GH8tjVWeVFAE2K+aVFSd5NZk17lBMtsjgkt3PRAL4axjtB/X7q
xMr5Z8HlCWZkrv5rbisokYDbKZX3aoXTTpf0M5e+z2wqbRewiRWWIKtUiN0aD31P/CtCHsC/8UD9
N1zDN1fdHCRcYuJKqKytbHjN0CJmhR4DFbiUiTXE09Exb3+2Q4FcrDDkQgumeGJ8brKzN7Tv7Ld1
pVVfJwUPnRMWsG/TBizU7F26I14Tn59e5DtXfrrQ4Aeo/nXzQDxPPZ3vgYyPeS2DeT8ICfF/IL32
yFsNo7dD/1YkDs8XQQr/KqcwQqfLKDmylIg6XxipYylpMkxenmFwI2kjPU1ly9OWoi0Ur6p9h5fo
LcKVt5QO2dYqpfIY3Cuo59Lf6MoMVHXXqZcHbETFWJ0Hcu3sueO3uKFTIityzXWn+AFrJmFin1w5
QR1toT6VjeSufnzoKgY+hXkT8veJVoOuYBxuwxurdgK5FCFEhI9DitLuf6qKY3hvwB/gUZNFE9zg
t2rIKzt0fsIzXZhyRrBJy/dnAj7gBf3Og7M7K9cGfBt0jN8i2Aj5sGqNrcpRxqmaNhCnBOUN+i1n
x3Xtt2cDTvidEJj/VbELkVgzRg58g83ZTZDs3ypdE5yPdzSztOkH1gKCArxVgaUdUgp677u/K/IW
n3VtmP21dy+ax1X8x0VmGi/FVcNCeG6KqLwyOxWhp+1FFjBAoY3NM9KzK2y15dQ1wqHlp5NtV4G9
MglbjABMgRn9X661bQ9EyStEiMQCgym2c7Jsk0xiFB3eoWVJY9CIE1J3kYN7I6boDhvnQB4hN7Ae
2bjqHab5buiqxnInb+PYxgqK3QotV6XqZGoT/TEHw9wOZm1ltIfsS+Rq8GT7YPo/WlCr0HYqrnhq
fLPTkQ0DS7tOvv68XhyJQba30tkkeUtTdRMnV9rwG8mZqQ0DvkNw/tlQYd5bc1ORKPK2mcT6IJve
oinW2ZJKJPTmaZmVsT37VnbZjs/g738EURkZ260sQXt1YOr6Q+S64qr15BYYzYXFuz7Po7hWvSpT
/Tm4EAWjQWJoLz0QpYdFn8HSS16lP3dtIaKMIEuiT6TW/Nq1gI8xwQy1VWgd4r64DdwwP/zrl1Wl
w4LnUSxoCsbRlMtBI/pMyzBK7Th7G1aXgpELctPsStUYxDTww7WR4/1QGA7QtoLqDV0q3Rz87c/5
i0GMfwRdrd7qe28r5tINVQs8OtLqHMa5z85E6C/W5v1Ze1FMvN+M6NYhbf5OdsfFeSYmKwjNBjAT
9mV3I9DTsHFOQSmJU27qu7Alb4xVkPg+Ht4nGo6oE3h3ZWHeDOkSe5D+rZ7pW2HwobMpcvimf+oM
lq1px0DecTWAHoh70RIKJiUYmW5Xa+Z2Fyf6GaXwTd6tEm14NLOKth8je5jGABwC1U5UT0XSav70
PEN+2PYWoezrp2McY6qIMAipMOxky+zSBWUQDJ13IdYE1k8GAgX3aGQ3z5OmpABR//nodRirezRx
i/J2vI7FCJ4gNSZBTjvqmLPYd6l5fVaSV9AcuKj9VF/2aPPmZkYeb9S1XHDq8MMekzVxgJ+ymJRg
mHukf6TrpSPLDf/iuk01SSGUl93JxA29AnL3+EvvhUCRuTu4YQWGCGG9UOa6psSsouEWfxCHNsQb
2Duc/lDAzuCWDXUAhAvdlSI7v1jdA8n7Tn7qDGEdtqJW18LfpkgB8E0Ud3NZYhJVdFJU7uwMtIOY
fU4WPhxhc/NdluMZqUfOsplbaKpF1RswF4x5D7wo8zcPDwIGLWnCPermF9YHGTwQammrk1D7mnVB
IspyqElo01H/ImGr16r0BSlsi+zvbomhKMJa/FQQ09LXbAmwOvvQn7OpLg0pOFPIg6x2XIgklU9f
npYXJFsO7ibhHb+3D0hGTteaJpXLAO5cpSgnrS+rnGicUUD2NtfUX7jEqd0MoJ7FaMcCfdStkwtN
2j46aQdbw7yTkt5ZXzEZPzdDD5+nc7mTw/SMWu3fXZ2ynAQDYs3oA6j4ulHzBxhXlmchskTRPVgs
thfrDDHZzkh82n9Cf9yxmtO8LJ9uJgUT3DjHgcjBjivUw79ZK4xNS2pGFdx39TBB8ImnwBNHqY1h
mPvWuktSEmdi+vr1Y6g8CtjE0KS9BKgdQ3rgAxZZ3xjguU1kLi+GzToNe0ZzTP9eGoUsohtmlW0z
YBwBPodMA2JARRdTBzLekqDXrSu8MlYw/0tX3YzCOlO99DxN8l0/LQFDzEaryk1udFU2dJVevNGV
9rF1SS2Iqt8cZc1nrLAfXkXnEWDSp4+q7zH2RO6dUxe3qcynYSdvOuFcddoawU7ujlhETM+Iaiy0
vsIGL2/kH2KGMZu0wUYkFZEKneHGRTNtFrtqhHYi1nI0/66iyUzM46bBXsAQJV3Bl8F49r2wb2S2
xo6pR47E0hbaCOoSqpG1DFV8tmIsIeWcMLN5bh1hf+iX3ckyPiNBFyPqu9olNo2VfDoCLTOtbLon
UEEN8GB3F1Rr4ELS8Mc6v8IDtEuBbPmFapxQxwSjP3nXoFZ68labzvla+mro+otnwSNGEVKhJIdT
PbMyDfrx39SBWjlweHb48Mm1IhW05qTFbi39uXaPxSPdc+WuPlEyasEUdxM2s2yBgj1B30I4iIQ1
rggKbS6gPaM5H1nT/nsoKR6wpsScHmM/fcnuQn65KG3K6MQt9Z4UdzsRoft80f584VbpyKvBi3hN
Rz+V8RWKVKF52YCZj3BACgnFKCAKsyIKeKW1CMLLqkiJkeI72sVJ4RsRi0shAiX22/kJkQxMGMtD
fTfi0RMyu5cmtBfI87aFjHUXDc5QS+/F1/2MZhd9reBtfXz9FTgOcHgCgkZW2/wf1ISMQBOMJXLV
mxyUsULh0fNrfEAILr0oell5fEaF394Js0CfzOpHXEFzHQidzgtH6vG8pay6Lt68EJ/Kknp7YPaR
kjYy7STSteoTzJi9iRWDL9/Z6qtcQPWl3mgARICz/6NQAwd+dNpimLk5UKZlPVBH0giCfcjjQnrl
iNmB4Tec8o/L2BxAERLeTWNihP8iy4awHZLM4ceP2ccXBa5z2RgJ6LhrxAMOuF2bwGibJEqzxfIc
fN7U3PBBqdLoAyZAu+WML7TfexdLaFle0gDkffs5nq4OBQkWdBgkHuHxA9dquhVevCd6SVszPs4r
BgNO+LUZQGuTzcwXC2hTOYgTwVxVLXRZbN3zqDgJ5eg2ItBcTkoxH94cq6JAFm4zgCCux0UaBC7g
WlbZuMiuRBUS62+ZIcMgraG7X7KSdY2DBOHlfG6l1awUH4PX2z4DTY13tOWoBNCFtXB8pMZZNaeF
5O2ChdCZWbj0ea4WJlX0XzGwpQTotL9POPvucFTVsb6Yu42MzPLHKoF1DnEdL2BnmhSqE2WBupgu
ekCD7iTSN/X3AL1aeXrqBas3bEZbV2Vmubr+LxR9clq8pkRsvemk4YygdGKq8YBGzz6ZKugvUY9a
+0AIPJ3NNZCOW/7HMhpdb+8whznnBEMXvZwRVnE8l4kYWS2hd9EfMqj7QXx5WxSyiUTs3ldH2j4M
r5zMqmtEVfYlXqs7dbQCr67F3TG7yG47/R/E7C/HeLM5SdL6Ri3iFG10xgbuUTrTPhuw1iTDmYSr
5ND+04Y/pUY2rovleopYF3BvrFmS7wW9MekQleN06xC9ysKTmAgDX14D3Q2YiMKPB0JOB7JlzOpz
V6bR6hEc7mW1Y/qpmXi8wIYksUqWnziEMtHq+eXYDh6I4reS0zGD4TNgFWtaYN5Mi3C2XSTOHEix
00afVNSlbYxDOPrZ5lMu4uu9FAehXgsBR+dKxYvXfUxuh+cb5+rNhFroetuMhqQPmZrHGUehLZqM
YK5vRCBHLXwB4izbdpluUIgGMbEGrbql6LgjlpyP/pD0gN3VsRQZHMMtdtbRGy+jWQY16Ef3F4Ur
vKZXlV8jPtyaa8cK3DoXfMWqprirv90rxJ9bLZIzHtsfKgfU9XpiU+sGTTaCQ30j51JF9cwDDcUb
Gfna70s57OFVYL2lwehHOb3/n9A/2Chj8atdKsq3at0erC9HRcU3PqSzfsr/3Au0uNY0MHbqW5aS
V8x53913wDQiOWzfHFrtq3c8OH9cP14kdBKGQ9nSr9V3qQeoXrym2NjERypzox59hXdCQMI0MBWg
sZrFuMgrcxCxldRVUC9bPBTyS0jgnuLtS8qMDHTCSFULb/6hOx9WgRYoBglADjFRPK1yPHUwBX2Y
HgmEruDHRgxzPQK8j8LrARanGKnDRrbf/vRq5epKcHtySND6fwm9daneA9ZhkQRz+DSOFyAYGPMn
GCt/d2OHTIJxbQm964rnZOJxVwrTn2bG+N4NuYBF7qcX7JWiEGseCqgClWK7v57KXf+x/RVUOQie
Ik6+eU4nbK9zQ4ezl60LWxuEukXOllVbuSpwQNam0AUNuTc/SfpNuuQiY5oieF0NdF8kTzHp9Py/
/oZsyYCmOAgtArkDR8l3fEZkw/tBZhS8zCezdRKiqqiI+f9NEIoEkFjKvHmJPpxHKtxh4Yq80Be5
SNqqZWnU6K4sfo/mPjIAxfyAwoupFUVAn93cZ6oB6618vsenFDl81JnIhWmDyK7p78Hx77Vuppg9
HNOwrb3CnRxz5TW2WDw9Rp9HudEIp2rH0m5zXVFXb50lAtykmKC7ofdvBZFBQVU2O2ZgsVM5+4Is
t3uYFp6nnCjPWccAfZy4fPNwlEAhjGIxPqR1UlcyT5Dq13L1JYPty/iqm4fHqu5RFvDwH7cMyvjP
Snu4JEBQZWCjAlN1G7mbutuO62kNa9llpxTDrzfMmVCbYT2Z7Ik1muJTs1jeqmuNql0klO0ABVsU
coUM3B0ui5LQq8HFXp1sF9jg2YCeD4fwTAHsKtUJCCS35spafvK+Ro0/0rcNh3BxMrBOSE6Vx1/e
7DRu1GK/fK8g1X7NeYKApb1kVm4oP9VtgBSi9fJ8gI1EXJ6RO55oOukdUzvovINolX4bbvZhMdMX
Axhwz0Z2rwNkSTKCFRskBC8hUn5tPEH5sFD4i9FUU8sILeC21vSfnqhlLKbR6w6GbZC7fdhDcDz4
+AkL+ZPnPvr8prHrOExjjckvDahrxj+/IJOaKoZ/yiEheXd3mDJaKeVDpgmvxQpzQXF2Jt3TrrCf
exEfcjT0HBMju+jDo4ZUgsAnF1guGa1tgeIgIOwltp37wO37BDIhJkF6YMh1GFYYrIp2Kef5qF8b
iQ/NfibExhUo1OnngGxAvkaPhREe8U0O2mJHCtNfL1oikzy7hbotQOa2bKXdynmSoh2ZMi3YKUSu
QT8aQjQQMcw8oboZG/+MXAomfVdICITanEyG2Mh5TyvXDY1Xfbk8AcA88MVdoamDvV/kAOHVpQO7
r8d/+3yQYG9V4MgBcwBzqKU2oZdbx9pGa1CvLMTgvZgDXtAPdtvmrKJzej8TUDx6w+vaYvLdhlfU
tOZ2J15msYCRrWN4VMZvJBkG4bOPEYmiscHtTyuBIcN178BGePfhZYqSC2cTUC1JUgn+TONIXcFS
tcb+pvk6IQ4GCKGfhnW2uoFMVJ7cAgwslvOit1ep8ko191nZql8PwhKjHjxs66NmdBtjqkS2SB9p
aDnC4NH80t38W+VHIyudIu8AsNhm5PpReu8CdotAHY8PeBscBrnUugBnSBeiDZXXFDhx9I8tSSg1
s9PJ2Q8sXYw9Ix3xb/t+GVIN1fwoiF+Jy175BeDcBomzbtMBl3FnN4DhCGbeJfmsiYw+3GcRj9UX
TBOARy/Kcppd19sAV8uI8WVnB7HRYfRloNrtlXjJyAgGnxbSaji54TVT5l1lAetgzp5szUgEaqXM
fExQzJl0pDncKdgtcvmfrUHb/mVCcV2JgzATlc362F3PxGULFwnNgPJLx5nFJ1MCCGwx2EirWTvB
OXb2JT9M706yMZDjAdOld7fIR/YP78Xzucqk8pmqmW4XltGTn9QFc3U5gGEC9aNmwqJ9OewlSB30
POKQ4galbynXH9eTVccmn7EzWTFnjNE2OpEWiTini7/4KIHBX2Y1UgbzeH5eHH2ttZQkOuKRVsyL
jVRfDk1kDew8pTGuSbb/qiHoaz+NdjOhajBpC1t07HTkm3NCbdDJOPdHjq9/OvKpzVz/8goo+8iA
RubWB3VR0qkyUSKPSgxR/pfeFURTgD1Epz3kGWFTT9+Nyj/TC9le84RtTaQopmuM3BTtBKTo8X4y
2NWmPdm+hTNFYePCYK/R3ma1PB27r4kpxWzXwS5B5iX9ZDHTkxpNG6VshdWoXNdmlbFHGxMJ0BLv
mG+Beb9WWpvR6cbP1M8bWkPw0CTeA5B3goIr30Qy3XGPa3bWf13uovU45jWvpJU0eLi5BIoQNp0V
6w9AHR4DQ496qHGfw0OVnXzfEkh2c5ak7PDgqwiKm9C//h+0TQohr7usY7gIQY070n4mLRS8bn43
91NXWCJr15HG6DYNgVvXYK8PRnkiDY0TvjH4GhZKtSuU2OtgZNLxMxBlVC3vxzewNkkHI2alXS1a
EMgQweWpJf80MwfUeNsyiwoDdbe2Y2SdjXjlB+vEnKmBkHo/OcnpjHFtpyIvnTHL9q6eQqnXxzAV
0SZv8f5vSwzHenCcRz/1C5tJv1ucy+87gskPzWucY7cmp58ZuOzls8/wwR5Lwid3fn+BbLpIKVVL
BCCSQfGKrpSZOl629+vrhFdoMEN4z9LUblIF7fWvNNeKCzhKS57kNymdDunCUSBGjqU2uNOWw0p3
RYIk+fFWb78g6FeSSOIacCdes3S0UwjnIZlJXECpw/3YWDyObQFTjYlSIe/EvnLRGlK3gvmqlQrW
SePdIHFRkmlK+CHeWIqnc65hcNInqkoBn6g7JhUx8YnVynZULIyCP1qyDr7/uDjNge55blx/2qGj
agbn0vwfb6tLzE/00l8nJ2l7ct4RTOBFQEnGtYSLYmqoL6hz2bPy4Ux+PZXL7buAUR8WI51ikKHz
nmmzdr4dV90nCOsZ8xKwOBH8NKaAL+SOqRa4vRmAur+mzn0N4q9KkTdqAxqfxJ6kz+G4pQ5yYzBy
v7V3q0j1DFW3Qq1DoDUER71dBkvGFiweRDC0yybXr++4jWo5VReynaFn+lN06zWFtGcO/2b+VFuR
3rndY5WS2UfHtvoVp2zHxvLNzwycmmLdxMauH41n7aNcIovR8mWdiTcMAikVSvzHkO+L1QHbnB6Y
SKVvSQ6Z/7REZ8nXVKhazqdR8nDng4j2H8UFPHaMjWPeaazPymBaAo3fsNG8qdKZFt6uhuL1cAtF
MByL0vDkLgwG1+5wwDzvdre7iDUcBPjCHtrvGyj8D22uWpMfYtuHEpIBe9jFaavZ6kegdRC03hoX
2ztXdDBNRJYhyogZrxPAQV9KO0Gy50Htm5/bnNGGtD6eFnZKF2p+E3n1cW5Nbgl7WZmk0Vh+Oo2J
RWYVrgby0qg9taSczqwpE5aMT1M8iZVB49XcyqHAn4FX+INu3P5w+7ERfGSx5oa6RKTdbGpPNr1g
YN2VfUfE5YSWhPVNSFcAmPJeP1qwXpMlubwGp6gQCx6EjrOEq4z183lhOPo3H5jG8G1PxdYfpPeH
00B6EshPUJRtoHj7HVacurYtTXWPWNWk4+nFDh87NmHpiLa3o02cy7P4nyitcDxNQR6UefOyDWMW
tuuJ5pFM0kmE5WPYsLpmhrmPEzLuQ1weMKXgoaHdluBMYF0JDPZFCCuxEEir/q1HkbNwyPkEWdtC
Nj3uDpLZ/LDr24qIcI+7gGgWhgarmeJgzrPoYamdOPLCUeF8OaOzq7XMiG9PdfFR6y2hE3HSzTx6
RcyRtD/JqReJzy0dU3aembZqUmkOPo3YUM7knRn0/mlMS9uAzkemz4Qs4ZN8Qe4lzivRk+IRbenY
ny+9dGlE53yD6Uz9nFB7C+dc8rf4vZw0g2m2FyD5UgxOpIIkqb1+KZxTmIGnXWdthnfb9r94NfpT
4/gNy0vZQ2GQx5EGSjhHmEvb8CNgiETUtjpe2rG1Ezs92KlTG/1NkaOk8Np2htbqnlA1WaBKUkH1
6ou+uVcxlunY8exa5xOKuBCsKXzkJ2qeyQfXMcGAGIbORGnAyUdUys32gj/JLnNIxaR77+ZBmju+
WAEWnKWPosXikwLfCKSS3n807UoikXczUOPNkfRgxFxlfyU3Lev3G9eWac3pdQHBNQyVJ0v4Gw+a
20J7BG+NPrqGJFtr2maWvY/siyxwUiGQAOSTrkxh/0My2uulGSGvD1GOp2IRlUT36YG5j0y7Am7O
usMLZjQlRjpLQszDkBl9TTAUC2JNQApKjh1aW9MOClZJQcGwX1tY3bJNfEI6+LZy9E6OS13HzmXR
b8KT4W020Jc1FwYbTzCwOXKKXhlXnBKNiK7HtXI+E4lY9aPUGiCk5dzMBqet37YQ+C8odjABulLz
osOjk2PGu4NV1qWY6RwIziCFzwW8jAciDz0wdwS/cbpEFuh9ssKdYSnpwtbnlgjyk6dWhFdGzZZi
1IHqQZc0fhdMRMYonnEGrcPWPCqah29NrDCGtmzqXHdycNcF8m6cLne0/VI53BWg9wDR6VzSYjeC
QvH54oFaH2AI+Rzwjcjp6XmspotKvO10U4Oiuywgu+ZgrPPM27zr0Oq9bpgTaEy0tPNbnVyC+EjJ
NhgqFsGSL2VtCvzDlFQUCOcTN0HNkanZO3uj3Tw37FBM8s4bNuBH2CKNBEc19zyCj82Ki3NOYpAt
zCz6v6uUds4wysMG90pdKFfv9lpinWcnsjHRKDzL3V61yuKoexRaa+vwpwuxR3lgYF6V4TK8Px1F
sHenWfnC/drQEgWGcoc9xGWc4u1K22agY2m+d942q9Kr3KZTVxeAGMrBy4P+uMv6DwI9qpNMpt1F
MunAxyW3AS6OIPaOkMd016+p55Gv6TBT5qk3Gx47osffYKWH/HZMOTMvz6vNiYAGLgM+fDvHhwHl
DJAtzUFsZd1Qb2MS9xUx0MB6hDZn+4TDYlLMwfU98UYaOyqSURNQ8fJ8JJu/7zSGIonziqOrONix
CK0r4NpuoQ7yujVSVyzKXDtbAVGZtxmG2qB1OJ4fsh7r7G1FgkmJYHR1DYXBfCx5RXZrQ4LmW+qW
aICRClZ25STE3B+sfM9W+pExSBAWaAiWPvDXwUq2lUymH4lFt63VfUHBtu7xCJtB+n5HxZ5oBO+d
dZxlIDe6kL1tHVgqnEp3W7bKZZccFKzS3HhVQpnqKwA3cLj2YlfeATocnWn2+HgXh7q0wlDVLCw4
rFZJb3SlpocXyfAyv5mLCZaYAbC3xUoz3rnFSXnA1zORsKweGvTbCc63NszbaptLoEHdkMMO8NPC
xT/1ZLg6XfdXuXpzzmBdJee0Pw+U4TtNrTvqIMsaxCSoArLRHK1168xjMYYVSqKGk4GSfXorlZe1
gkHKfs3btiL+7fcxBtEbThIMGHHnm0XCgqYp0Vhz4dCesZtNdwHw0k+CPoG8FvQJNim83TsudQHS
QVWMxVYmugPoooxFgQoebTibCZhHMs7ww+TlLmgB+p7gux4U8ItnncY6s6ed6PoLoy5HLtsz6nuQ
oiGNfsG+y8MI2J1E1ZBjKsJUcbhGnuIYw/GAuCyYyXvL3A2qluI4TbGO1w9ict3RLrSkYOtD00GV
AkhFZ0xHyn3K/FmZv4O3VN54219CH+rs4guQLIb+/iJTOOMdvKSZBh3reyM7x9N2BFgsVJl1+ndr
oQqNybkvpFq/rettX5VQ4FVudG3wN9Sol0g+k5q3YM5XS+TzfEZAhzFtBUwwn+Sl020lkOsBtUhO
bg9uJc4tnqoc5N033ifupPScICiQW3TBYVqGc3Wkrhveo7fpYxYY++LCmdH7tMW8ZSWGr54fj4cs
/C5pQ1EWzXeAcKWNI4SOo6ekVU8m3xsDRbgZc/Voy+I24X96u6ugQEZfexMcn5f+Y0G2HKRKbOMk
RNL5JNHCqIXQt3Jwiov7u0C0WuAFtJYEwFx5aLCtlofF/JDNeF2EOw1PQcIzsU/PFRiRonapdjMh
RzG0gT+VdV77CxOLYUQEy67h1zbSW1WZry6XadziG5O18Sev8eU7ffooxKed78N3uNKQ3QCWVe6L
3JMRi0pDKXEO18mKYIcpejaVK6r+mYz2Nde9VF9u+oGWaUGHKJ5eKElQEV5SO+adBkNZJjsoUaSH
/RBS4knmvZYiDDIQ3IDJY7dn8tIRXnGcnM7oLp6KSGXDnwwBiEhEncIMCjQr8tzefsTHx9RLUoFN
U6yIXVvA0nJ3gDzKlSJ2YVna9QNfG0Ij6Tuu0qa8CDv2NKfx6Ug8cEpFIRi+4Z9BJsRIDCHosPsJ
gOgLaV17kng/XQeolpqOTdLmHtKcT7nOKyvlCaHUABR9t7VkjkH1oIk8Wyete6GJVcm8MyT2zgJK
f3LK1bBsNaSdiINFBYPH+hhGSxqgff7eBCdFIFenTGfREDxGVyw8tipLDAeZQ97tIFxqYnbzzX87
ZP1ayin1s+9hIud6ONXw2LiESUuzmSELACiez1VVxkUu9kj5DWwbcGNRBUN4gt7kWSGrEsZLunWJ
ZojmQ1yZC+VlYW7F1zJ6ORMa8GMvGn9FGCTG70YvrczM4x/A4tklUlfdR0R8VAkpRu1asCipPBIB
p/+l2zy6FMiiOxI17nIlWS9VU9ugr41Nzjyix8eitugWsyRomSLN3GJYylKvu0CfDM7GRB9+ojhZ
Wcbqm0QNdJT1bFNzIh/NcGdM7/4/rxNOMtKGBsj6K2yhwoFxc+8AfOzTS6IYqlDMDPqSfpC8OMrj
TWvSNP02P/Fi7LUJBOj8nRH2N6SFcFiLe85x+jwCtAEItMfEatRaKoQKaVtOVnd3qzvnFDUa7wUQ
R8InycYd/SXYqsDxWKJS9fsVxX7GPV+ACVn0gsAusZuTBw3DwB8phNaOtdVGbV0p0Kr44roanjlB
kLQqMAGUMQktDwaMNPX7/DPezobltn+U2VM9MglkJgT0GK+kwjRus2FkqjxUGq158c8bBmyLCbmm
WxErZsjGXzVox4lZUjQMwfELLKATjsZ6o44zKe9l+sjtsZVJDBJLWLA+ocY5H7fSeTlBiIe5llLK
RKfRrHE6nOeWz6TfuWdjZjClSaQwEox4kg1H7qVb+2jc7JUM0B7ZWBmagBl8Uhpj3102mJ+7v0IM
s9Hupr5nSvXWI5XklYfyf1ZBdLu9ZtKNV9zzMB2Dc+uxp7XIghuY25uN0WKOL+0/EuAWWkPMWt1l
/pKaeTd7WD1lovgFQpiakmZLUu7gmBHUlpLPodwq7yEZS7XIDYWpy76BvWVxqtTVliHM4iTL2V6f
EnvWkJCNGIoejcbkELhkHdctQ6whS5I333ecXnYYErmIx4SacODW14BFSp1stLu/J2W+OHgkk+Ly
28rboyEz1ZsR+YZXOPz6WswIE8Licjzdx6SO27msYtPu88KZDBmQ1x0HDKV7QQjw4FOpI2hbrJD6
vIfyR3h9u1ss8QFYXTaqLbbi7a+cGIAQI52Y/oE1qVcxrk3dAOsMCio+0O9H6Aw0ok1Uzq5GohX7
T9RLLhNHDl67rzVBIiOI5wV+v0jSEFV0DfBQVS2Qrx43BZJho2IKjVRWyirG0MTguPjIrpzOItR/
VKSCjdPgGV70g2YSKBUSMlP81Wr9V8bKX9QLyaKwTKHOYYzw69JFYH5T05rSOc5E/j9vE/UQoxWW
Xv8+dbW3x3bWSO53cURxrVvmShq8e/st3nPccTKiUUgREVVSiJbXOfY6pbGzQcRF/xerYQD9hkyH
zW55gOcKdjmr39mVkB5FkTGZIyBYryyoeZjzGSe6TJQWqetjBEH51KVi7C2BXZ5PY4+0k5aSsqsT
bbCGFmKPRPaapcdXthbCJQuwefZnY0z1TQ6L9Nmy5DdA4mD6ew7hQ6Icr3B3xpFqLIE2g1wXULKk
jSiHoqs6LibdvLvbGEziMRGwu+HNlqdai1sOCGZ0aC0PCP5HNhxoy3HfYayLA+He8y01KgeJItLc
h6YOfqjh/whLzCml69kd5V5oG1hGYzeANcJXzYGZ9V1Km0BRheBgR0ojoYvHby64wK0AManl2+0q
LZB041h+7ptp0MaISObx4rx+Md0bJyTBC4dqoKZhdCW7XtkLxcrSVeb4kGdVUvdzfmlCKMkn0aJ7
p9oom31FXd+SSbs6gfIWwwz3X7yCjxWxX3aLgzmFJ9YbGhUB3v4c6lrKPaA2S6yPe7b9nCwjyGeA
SU9MlcfUoV0I8MpC2RiMUFkrvf0Vtfx8gxUDlMgmGLQ7NKBjJUiooHIY6vP7oob8B3mjLRNLEkNa
SQwZB8Hfws8KTUD2KvDKw4GKTZ0OJZ+sa4Ua28gvXEfT8giJPiloZef25hZZt6hgHsPCJy+zURxT
ZJZ3W+V6RWxSn7O2zvjLZZlSih14JEC3DUdtBv7I4cMWbbe4ACAYb2segh3psVuxJHGtIrRw36nq
IK3UG+2diR0AR6MozdaYUZCQlPGV2LvRxvfM6ENBjza+uHoqiKT3FglS9YrZdtUDj8axoT6Y+eAo
qIFd6jMXOEIKhdY1QRkhout7s3GCsIqLuIqmxlDsr5DxVHHEBOFEM1bemXrphQQMeTqIAT3ykWqg
57du+11C4bTzffYN7h/cK/HQaFsZ3RhjPOoS/hQXDeMYKHu/G3371DB9+g/ZHXh3Us5sCthMn+sK
DQJEJesbVbnM7mYlD98CD0HVpGJYSwceZ4HXTMLfsG8H4e32LRIZ5bXDbiEEjxlIVEwAbQwSnfyb
Eu2SrGp1nsb4aodg4nFazAcO0GFJiZM336j3zV83RHmJt2Sb10M5NyaolaoS2ZNcRPTJI0PRptck
Pkjeb2J6AYvp5yjr687jLxyf+YTKcTE5Dzv0eSDFGTe+bftLYo9JFZjsIPzsLUAYZpyBFh2bBo8t
GqK0EulKYJFmSKpnzp5+nizH0+6eQugOKBw8SEY+0+ScXEtJ7TjWfAD3wy2XZbMcdHFqBQVT4HtK
Ms9oXamUt2zWU6BEb3jQMW+TVps2v04tYhcl3H5PAaXQuu53RbUmjNkCTrMdjsUd/bRgoIiDcfp0
axyHmAoMh2WdDgl0lSHoHc80COjRG7VDBqMv7EvHbR2646VHWPRPajmoAWbMq2S+QfFcePfrC95j
QCCBwiCQKBa9ilT/NqsExwZTj42BsQUaV6hUa+0EnmJsLF77vsL3xLTDIzD5IRQZlYoLGuN9szz4
en8pTdiRyqGTLlTDlr/gtF8XXwwIHE6/64Le8QPp3LkpWHQYsHzZDz/lbBJsoIoU4gIZf8EAN38T
JGi6F0gby+/YMMZyJyfLcnzEUMlt4zbeQ0CGhOsPxiNmdi1fEGkdceY5zN/75pCrmgCqOgbwDiVx
2JnuL9I1oCwST+mXPCpJBUcE6lv+XmaCu31wg4oQaWr+5ZS68yl/VcT2hKIfK9y8LNGWCqGq05ET
YJJaAt07Bvhl2CQaLJWbByQs5iY30vcYvcWl7xy9urP+SNlqagnP8JoA9DKj9wh9t9Kdxak7DO5T
JaKw+/WKIVVdz9XKszbfIR728FhNupbdYFHraYxf8T1NbYvsN7Il6dCz+hbe/igO2h53Ivhl5QrT
iN1+VXY8zMMCMDZyqI+3P0oiP5kIKPE9RFpwq0hlMJlG/4dVKASYIXWrye2IidzAyOfAwOlg7k9U
tIaWBRTCul1mLZ2aMcSNGcBU5c25XFDVCMhpHMwM6QE0u0uTYBj7Wy31Q0NLoAyFB8Bb5kS/Hiw3
BTUaEq0PERPQnllVeXmGNrq+El08WQ+jy6XBguTI0lFPCHNUGDxL8MQdmcEg21qxT49FR0dFQJhI
kRtjYAssND2sbZTbLc5OsVnr48jVUwQ3V7LKsuN30XXVSB6qc/8Xq8nEsXWkgm6ZKJdHL0+EnsXS
DwzV9KKhpALlYV2PNGsGBZXXTqol9WxiR5fG/7RP++ovwcKkygvc6g7WTNqZG4TWPLBVYChtVxQZ
l9eoYtAlh34dswLSPtN0Elcz13QxNeFqXcH303m5JVQa7KiBJe6R07o5ui5LXTH/EGxQgDL8w7Yc
xtnP70dcf6PySp430i/xiZgVP+iTLW0yytSzaRqfIN7+n9NYnbzT7qjz4uqYVIQYjbdGL6+f9LGp
c3k/YGBreDyg3sjoqVDHZMnrtRer21HvHyGBwgCF3CJbD8UhkiF0kNuFWXZm4Mb+orZB4LtvftCB
0warhyxbCX7iXWYlf2R5KMKu0QmK1kFeg+LwGRew6lJxnHg/RBbi/yXlYz75NSvtZcoZQgCWcN3J
raUHKxpULsl48Jg8x3heY93Y7au0PbId3micZQXL3uCVa1uQ0fwb0/PUx55lLF5mOKL2b00AMH2P
LR32VFpD/37+cIECLVrkxP7MS3qUlv6JZPKdzBNfYVkKmj25gFiRYvItw9OC+Y3d9cqd8VqlMxB6
BPNUUS0XUaGT3HzYnFI4ZOXYXOczlrKZ1u3gNn4vY6xuUZYtIRC7lHAgCmwBaFA6cN7BMo+12VPs
K/ftZWjtK4YaXVgKnhi9T8HaOLH5zLfBqSjO4aOR+9YKdMkXL8vPoi220UBFpjZWADJs3sAbXDIA
HIKv74on3nBPvLoIZA41KDKHYWwDxvnfR7LGaA6cTAc8QJPLjXZAt/K5ZNk8sPZl4DbXRdkXFriC
52CCqqX16h1KEcLVX54NL1VOtODvu59ds4BJSS+BZ90bdd5VVADMujliFRA83HS612pAIj5M79i7
Wn6I3kQAQTPCTe7i6quqlEWKIhprC3rnm1cSw1gVxxIvoqgfVovkRPfVhvpTlVHQDQjRGisCMStS
0Ug96EhhEuFKWDjwMZ0YpBSTlRC/BXIrZOLk7TajK/suSp7/RrNmZpm90CzVmEsb8kkT7V683+JV
BpOGxwXy1YCfuCda9HmjjwQXp2ZQUSbKqaeKOW8iPZkgLS30pkDlURomHQ8Q1tj6yYApcD8c8eMP
3avFELzQrdQlS15cs8FlgPulggqWogzSnhM1G1Me6RgWIUryAAyZd2Hkjlr4hXw/4w90xMiLQ66R
mzHOy78oUcfNSpeXzjar5UbxEX2rcWXCRLmj8Q7mRrNixEA2D6m+rWTSFyrja2+5ySwyXTv3sicX
SgBxWfMPQQtfnzT4Ffk4hVHAyAypdntLTGPRxfqsHrqDsHX1LgElk1/emMOMtQvW3Y9oxiq+nsy2
h98UR33fZ/91qjyxf0hN68Nt3m97k8HxFmZXKMJkXnc4z6+ZbVl9kq1RkoJ4NtCEbMfUwLI+igNP
MG3tu3JlscMMAXZzJvThJA4ZzJEBn4c/kI+eH8rD4idrAVGMyGNJUzElvNaZz4A5T2eDAYrmYvsk
Pv1M83n9w1WBVGMjKEjYWiIRHcC02MZG27fH95ve8Dv91WZdM6FjgXV0N2Y8+qediirqR6A0ukrn
IA78VQoJ3qUbFTvdCUo9peGMcWY61Gf5ZQ9y+q3Z13lSjO5slNqVnMKZ2gBkdhZIFNZyjg8Fe98C
uHwcFSJtFJnkWnzpjdPYSLs2Hw7as8ltXCJjvTu9mCq0FyS2x3Ky3ui6jiFNPTRtPY+hn9iETTzE
ZwyTL2F7P1ZMAEgjU8zHEu2GSj5VZNlkU6x7FY8dj8FOut9mYkrZqqwzJHYf70uVUGMGAv/sgQ08
45l5/lNnz+GMvrdKIGuWK19ZtH1oUELAtXnUDqBmV6l4LxGmCa0E4P8jC0k+Mp96/xKIwzNn2YSt
RrTWBqfRSfEkQ7xdBC747ISKpxvddyv+9HbwLOxlITbigezTae48WcKL25BEsB3lHmbX05tPwHbp
jdOsN84QD4SGs6lQEwZMhK7mttDg5oy0kQeSyi77OBucAlOtEZqTbM8mmb1XaFhM8C+iCe/9C/Io
aQ1+ivrQtpvsZqdlcQvLn2Yw08qUOqFuiz0OdvDEoi6qcWiBdZi950hT4O4l2+SpOK5p5+Ze5Mdt
PdEapvvJEHt7Eg4LfT4DXJeAd8JCBc6YylS2p/XlNhB9fHAlfC47w0oyyfvlV0MYma7ZflLjcHg3
l12d9+bplUjfB+HednD+lQ8KyLH33v4LdXHMtKN5mco5bN5OpcaFLwXFUFcIBO1OSatogMe37j4i
FYpEgRivim3Hsmwqy6ndEhhHhMha1FWo3vhli/7yyjrgyqhSBPB/GcMb8ZrKURR3igOFAUTJTB3Q
IZsk29sGPqNyVuE/BEZN1jmqucNtgbX2chjNXQ2hIqISmqsnHl+dsSHW+AGHs3itRxmN1buii+Ia
kDlWLQnkfhlrnxeE7XZEEB6Y+iKvXp+nv4a+JhPes94Ket+66K+B+9W7f06jblM8Hrar+owDKTkE
jNUQzgRCjUrk2RIdSiGSWVjvaFIzhFPkGm8gK2LwVqQLWE4zOtJiZI/MQ3yGDte88B55vnM85UoM
f+GtJx++SmfLSli/tr4AI5T1xGTH+VHDlxL0jbxjfLsOPUI29pEwK9roYvLqiMV/QpxxJRNXRrLI
+RAgA3vXSbc8oTJGnDN4qvJRYPzO5WEtIKLUGgksA7yCc6zuvb9JoZBGUEBqD55fkaeqd79OeAJt
oiGmBY6TykPAkjpgpAaCotYdipKpni0uk62F0LYs+iaOYLhtaQMoZEWqQDXAh915XXsb999YLjKT
iNc0nCeqRXR965G2djsEVUIZpGMxxYo+82dIxjel9uvQMxjKmoOGHX2a+TgN34lzMb0rLlS8W4tx
Q4/NjdZtwQMUeUUfzlZ8DgBMKpCO00VrUGUjvHes7s9dVXpo15paYhW3Sidlv+khRXW/tJA9uVlU
lTCPRszF8mv3kKSDl6/+hDrSFj3NlNT9tnpIrhY0D1sZNHxHL6wF4jrH0Erx5grdY71e1FobehYu
G8EYGjwMKc1BTAVhaZEyt72lq28KKRHdcAx2MtYBJbOPBASYwsk69FQvX/LYnMpp/Vr+GZDRbiBp
O9rtdyoABrdU3o8VAbyF71XuvUjYwsPbIqqvBLAzMDtQdRRxtvfBd+tUfkRx9FYkYEKjjQDdblWp
Z0ublhs0Ycnx1t8SWGf02U8EasHIO60DkFLB/cilmwBPbVnivUTiyR7Ssmz+zj5rVhyWLpOkTqre
j0xN7SMf1aLDam6c//hnCPjcw6weybx8yluwSh/AqKlVS66tSLaMMy0UIBiDehmV5nokyF93ho7D
XYzjcLUNvE9pNdO7bHhOsbb5oRvgubvrq7HfiFzp1DEn029U1d03aGEi8smDvmK3giZChs78UshN
Na502evA2wGaxJVqKmUj+OjbbQOo8qT2T5R+AXEeIjlxj7X+MJd/v9sy8LIDLiz11UJhY9lJ94GB
cAYIX3sptda95xX6/Cq+6EnbK3m8CRKXnR1lUbd5HTdeywS/0AMrjWcKWEo4AXnefj1H4wK2F5Qk
as0R8wdd1uApXV54kke7YGkUwHKbQKjQEkfinVoiGU2v1jWUwghp3+VQwRW5xYqnDgjlHmqdrHhF
hpuyVd2UjHobRVlseLffMiQoylfJCfQzln5fvh6MgxWLM25IuAP8S5rQIjHrC2J8jJpNjy9vyOAH
Ipm3c9JPv1vh89Odz/0UGZFKjXc3hnhkLbzAJ5WlLcCpwVTge0spLdwJJOoCMyJkNdfjAKqXuamA
A7odKW46e0OkUQda3iECA0W0eTkVRSUCpxS80JCB6AJLMzY5dHeGoEkoBBaQcpC4lJ1xaEMLMbcj
yKpyF8UuXT7PlthKN2xZTFLhJYtb/WV5ZeXNMkvwOHx97lzIIVG9wz+FCjc2/DiSPihJX+f6577u
vAD61c5mnJQ5rzLj4bmdmyT20GrlCSG7elbNQu+HbbFQ5G3QDNGginXMX69vZq4aVHQ02KX5ReGA
uEY/TjIpWABy3r/1SxeLoqj1yYGjeEXE/lUDl2kUZ+vbtTuHDLIYvwNTXfJEyH4Mj3Zlms03LqTb
`protect end_protected
