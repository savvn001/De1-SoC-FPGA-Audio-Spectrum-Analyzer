-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CYt5Iu0Q+AQ+IkMRXfC4jUNkkXvQp8441lMsiDek172jppBTYcO5j05LhR92wuZGKeB0wW+Kf4kl
NwCvC0mtoBEDnh4Ut+YX4DOd3LbaAtTcG6QwBldfC0q/LEn18xyY+hiwQEJMdGs4OFLIoZGtXgn2
p8+IERlylWS7VEbKn8HMRHHZaug2vkRWStgZLwxFqCuKL30b59cBAftsgwLaw3Iyzlht7rCcNgIp
trxn2unVB6d1hzy+A4gEuN6DaGP7FSSapUEY7ddkzV9meu2Hi1YG7cu07vjSmm9dr3VuupG7GwlU
7mBjWRZJ5NmfgSqDWnjzf+0NfCUBeh/Sash0DQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5808)
`protect data_block
qNjfnYjCTIbW4I9WAfY6VcsfkWLN5riwf4qqjl9Enbg3+wAF72efWPubsE4qpdN1nGQZ2qeuQ9rA
wpWmnH+55MZBiqzEhOUCIukyOJrrkKv5/Xry59eqDK9y7gQjLcnik3lBNh3LkWLvuJvtHcUjIZoE
/2acOXN83C8S/R+F+UvOktWumuktbQfwGjE0n4zdniqfETDDMCGcXhzojTJCoukLbzMvrMJJxYMp
+R6tL8tWEEc67FmBWFvmh71NQ3zxCLsM4NPeJC+akqI9i3ZhryxGx/yfcm5owA4CSn4Z/FbwUU7P
OMW5Oe09v0iEGF/5gETV6VCP2HzIThd8CRj3oCpE6H/cQZCGyxAHrGrmYCBEDzZ2UqqListrJXNB
xk3lhz0nSvWbPsYHKoGHrv+TWNrcKM9hs3nW5/0GvkLX/uPapGc1UqCEJwH9KdvDhXawuLbifAE6
68lVNXjknSW7IArNxhrvF3KU4tBu28uSuKGU0bxqvKfiVliYcdN3J27QqBWyOvblRS1AtqJ569d6
E11KBauBDsxK/7KL4rUh65XdnhCBSRywbvs3sU5I923gMMT3FSTphbnZcQsLm5a2lmHlZPzRdaNl
CQtAp9v0rHXde8O1aXge06j/88XFqMuS4xHHKn/cXJB2qgotIu+p33ktALcMx1sTQ6QGzK1luhgM
Lf1ozyFrQ5EVbceVQFkbWYTm0rhTd5+phQqIfbqy8eWWTlN2qS7afXX5WwQ/jydo0CbrLBKBqk6+
iZqKFPvQutjWs9rOyPzWRSUOGjYyKpBiINcQyejsXlWKgt9drP1Amy9ILpFKIMiHWs9WMxD5JhCS
DACDRdUkYx5HAhGkva7lfSEpJvdFKeoFDCF059OtvQvdSSvKnW3af98IKp0+PXJac903D69pTjuX
8OON9lkcrLH1gKxTu6e2J1rxQk2pdzvdIt1x2FcC+RQ5a/wr8gq79DYmneQXuvYiki09x4v87xqf
e0cIHWVfGvhaxCKm2bgM5GheOFkw+qSuS+Ecx1NO75UD5SsvcjAfuNYzO/XGsnMuMHS4RTCJMK7J
PsNA21UKE0nkh3gJfpp1mMqyts06VmR24P4kqGOb9BJ6NK1IM7cdXGLSFNiNw4UVW1H6XfLSsbA3
E1D/VkT4lJY8jwR4ijCUXTDt9F/+6aBHLezw2cR1Aw9WUqcr74XXUScZhkjANBr20oj2O7N3uAKb
xRygWp8Ujz90nAb0gLPBsM50y6eS93rlLQhnGJEwvcM8papuQqOAQQQa7FrU6SqOi15TPpI+BQnH
yVpNXXj/InCTeaTGiaU0V84FNOyMLAfw1EXh4oWXG1xU7IFxJ8Acwfrq0GBuftXfg3thBM2F7ikm
jtgFuosgbxyIe795SORjmxMz+gMGMsWjmAfcyWUjnOXZjO0WQVY9R83tMstSGa4JvYViw4rL4U2s
FxMTBbevaxQMalW0GomCTp1NDekfrH1iFk5s6FXWaVSSVQYm2nXpwPdoc0BI4dyazkJ2c/KZ/khr
iy4N8cwX/ebkXjTXwCUJ59OO4meTh7+i3Hi+AGbr5UBx/FH7ZwoInsT9dubOdDl6sm5j89iTWiQA
ZSBvltytBCGcAYrSzb1jG75u6mbYHeTMyvjwx9oYC8O+ct/o4WpkVMDCIop9fFYx8AtDKWADDizM
CtRsk119JSk2/RhTthCND+RrQy+IUp5B9qiZaaBuh2tMuhy8ImvVRzXhsp2qJ3vIXBrKzt+eX67Y
vVIxkAB5pGa+wtmJYqaEPMjEmtEwbFJUAi9cOVVAz9m7yWVrMbFAd7FK6Pi/XKPrPk4xRYziV5HK
mTtfOQoZxMw0ab+HhzpoUml6Da+GOL9GVsSsnbT7XG0ABeG32NIkmc8VQMljuglYJqC2IociM1ck
jqKLSK+PNYYIuoHcOpPPKX8RGMTngutS2DRCnTfuEXaTMseVRQNzj3UdIAgStDwRzO10iZXSWYZy
oI0x5OGbxP4Z+DWYFgD1bD/TV6BYmTDKKXgc5ctPa+s+mcEwHdWcp+uWmcry0ZSZcZV1UoH0GGkM
MVJHbvUJeEsSWlCYVlspirdWrge7A9Ad5fS/L7JDscX+55csGpvSXdcFoxx2iyXdDkxY1n7iAbQO
ONrEy1p0dFmquFMYESrxD247gRogVS/+zVIsSafTuUVdGu7ZGwYclEYwW6bV2XBg/j9biIq9+yIR
k7LcCN0AlZXkefReEUh1uTHMxdPlEdwYlIDIbDxwaNA7Kofuqu4IEu3cGPRrHKgpSLrV3w0Vjpfs
Vy6ryYYm4erIaf69n0yUUYCW6ej2HRLZvw8SGwdF8l0M+9MAFJrPx0xGyEKNk9PEbMqJMP9jw7U8
N9bNg7LCpQRBqEEw0EDSFZESwChL2JBNttc5qdm8+ukdEtfcBbPPN4e1IzsCi+pSHDAt2cpBVjH1
KvIAnz6r08OWyWPH3HHEvpQMy9OHGG857oQJFp8kwxGQeKTIJUscjkxmj39vM5xVbyIEOYCewCs1
D5x2ARy0j8B/mJxfGiU5K6mogHlZRfoJ50dK42H67jY0oDkoCzR5R3CTEqghZHn1Tfv5vdZPOjG5
HvDRBzaIa6Xj0OnbB+wQRPnCmtlmRb0N8b9pdVyVFTaTDJnK6ccyYrvTgXhwMVPSQKdQ7mTPm8Ac
E/L55j2MX1IqiIQ0AcvZyFr7cSU6j1ty58vNfvfp3egMo/qdeayT7jMsVZSMRqkg0zcrclfHCTq9
knB4O7/YIFTyrdDIv4QW/8upM0XNAt8G7gvJWLGnPxOXMxfvufrigtxcMA4SqxcnRJRhwbAu8mkP
vyvuW7mLos3LpWax4UkHJPsjJo/yw1F2CJIEqU5H+DjvEwGnHKf0QRrO9orT1beRtDV4fpMpmILS
f2u23RhKvFAR265KQZsgvqRcnAbv2jdH6IEGiHxWUEDTGpJiulLL/bZIKSwrr6HqqxBxnUvpHG1K
xJ2kWmjJrxwxk4YT9t6/Dmwxm3nuXuAFDEKe17ABANTfIqD2zbqIaeNSrCsO5nLKvJzyOVUgofWY
dOAKa5fm9T7nFPoOgtUetvtIzr4L9+eVfIfE1GgBkGwJVTlTRMlpZjPo5Lh8UAJqI/941p2CTLFV
W1gW78mIWUBRi0GIctzv+DsbtbdEpItsE/OABy3Dv3bcADI61IGkunT5GH8CTy30Bt6RZfP8pyTU
uCYwGGBJ7myjuZXDEI73qBBFWmiTVpqE7qG2OU/zbj1/SQS27xAMYi0y2zyyEmp2gntoo1LFGgZq
IL06So57MUPOheB3V3+wTmUjIGbJU2FuORQroBSh4iX9IQUq+5BKQtD+1rNahmOmSmrnI7w2w4n4
vsv/+tkI6WN2QPYyHuwylcZDEqHUTaJXO0dugVqlZ9iXnYTtbIscTfT5yz3TzqatXIQIokZ0Qiee
Yb8EDlwEwwOw5lyqLNjmoteBJv60I5pHyHUCmCa4m474SxmChaqJmNOAW26fKJ0PioIvLtNiax2e
5W8ca+NSajRPUurP4BXqNDUQggO9p6mlAF/ZazY5HVg1FPqcSqkqO1Sxf7DfnnKHCe/5BkZ0uRlB
uXy8q2wOz7H47XudBM0Uz8iFoZM+bO6tIQkC8LHvr7Kj/pLjgSLMjCLIrGqMchMsy0FrFxujt6Oo
KpKYdlzYMwX7tMlBu9mlILMe8jPI9aA4bVa618YS7gt1+qJPN+bIVrc8aAHjyr11mZOv0H3sgWnZ
mMfM+VP27c2TTCRKCue5RGP0QYzc9YIeBS6dJdrGsKRK4yIe1av7baA8XfK279iRG1et+3j6PSTz
+Z9K4ylDN6RtLLLoTSDXKvVnHaMtLd+X41IoHIF6JkWAgp3IDnsuU78AEZOKpewl9PvlOFLm/8xM
QnPL+oT1BNpmAqEJF178JH65ii32/eOzULZGTS9wSXvi78Zaca8mJyWz/fA4T1KQGDvPq62fvbKt
qrhQx4JGYQPci6+jFbN7toPUzh9froNkoXtKDD/7zCbgRVwEujJuMnDbxoOQBnIpM4cfrlHZqOfr
u0BDi8BxVgNETRPgiSoUm4L9FTqT15UpMKvmrOHoooiYSHOF023xE4OY2iAQSBa/CCjqKi1nKqsU
vFsXNTOkQO8DhSEdWf5S/TwRPwuEqB7u8/4TecIwS4+jl/ZA6pb1m2xSjYQ+07ivCCWW8U5ONb6t
Hac7WoFWB+dYiIKD8tkzn0j0KNDUv/KITzcweoTCTUkSji6RLT1LaMqYyyWr9boZ6/eGX+LDfTjO
9d4/snlw48WZnrEAdYjYQzw2EEYx14ZB5qgbWXRY9NmsDheXLouyj3piyjzbrmiVZz3i6H40wvZb
EezzJEnd/VshE3Xz829qFeGAExWvA+fkW9O7l4JgfhO+BorKY3Y4BmIy9C1xKFtYOKQMhcf9/H3e
W0uC+/IAb5SMormXwWqOnxUjmwqN+meykOnyZQBhhp0wjiymqCaapZjiJ4nfnZqcKHyGWJAcFUjp
HTHnZPCiA2MfTaxHUhN+lXR5Tfcw8d0Bm3RC1LSEIq5hLLRO4xc/SFGdcqq67O/ohjMjW3AyF3v+
8kRMzFHk1ZInXjMcCIMAMVfbCe52WROCK8O8JGiOmKEvpTljcwmflNKfLky/jKazf6EBf6R3sX4w
Ev4zJYwVSzP1m4sxahZUuYKFykm/zCPhA154brioOYqkGrvRW3DeZ8V+02lvCJLX7xcVPS+jBCCT
v3+TEShZ+HmQPb+gO/2Ss4XbT7C69esSubahIkEMBazPociJbKU9yFnGqpB9N06mNaEI9Gbk9dUx
6IJNX2DFRh8OkSLocvAEVnyc6iza11zYU01+D/pyF4yCn5yIW+xhzl03ICx0N6WOgTv465Rj1bCz
yp0aS4XnQnPE1X78zgT5qXZjT4g6vCXTYoIEuiX6MVlZaBKbQH0Ul7W2KtFn/NxtXh3M89e9gvwP
hWkwRA49gGW4fLZN35WC/Bu8GgEjiabg3eR2cyPX3RkCuq2a1jgj7rmSTTnasN0XLutpAVxPDBHn
O1meAysACPnkEb0+9PRmsefIL355+FZWZOtVJ1YBU/YJh/Ch300Fn1Un6HZowmAJXUzgyKaVkFpg
zDSSMV2DyReFkClZeHNCzg4qwChYdXnR4jh+lxEdo7f5C4ee95+CXWZTSBD6xHPq4oX3bxMzz66A
8FPkZxaabgdyhVeVy9pkaOqSQSi8QMdJvyo46IW9KYOVf91L66YPmBbWcQu5guHIg4oy0jDT4kc6
Vkbu6cOuxa8CMrfvvMPz76ori38TC38EQYbh30thsHAqHgiHYE877bKDjvEYM7b1pjzu7IJUe0np
czGb0rn05aumY5CV3wJRUFMmuS4/AdTvCJnrxYu0Em6ZfaDBfGouD3h7CejJK07+eifQ9iDtEPlN
9TL4yLNvp7fcOX4YmsOg8kJryljHcAuNjW2N1DsxcIEg0cVlrsY14Suhue26fcfGrhPJ8ok1k3NC
mP74XnVqFqAn5FCoop8RD61E93B6cMS8tliPY7oZPM5iZitPNFmeCglM4F5y1baz6d59qVO45+It
A7dfYma4GyJxUi9wWU9M6jolujxfRQUngHRQCprYb8KYEWoXzKEiRRDUq6oG3+nrVe3A0dIjd6Ot
dtgWXKMmzELCzLDDWcFTRx1sN58lIsRyyd0N4qWtmLKffpFNKIkruG0jQAaeEobTwD4VfyQZz0TN
G/u45s7bw31ArR10+HwX4mgyv1o7hlXPX/l2idFf76xA5jOIX/1NY4TDw13EUARl33Z9IvOq0357
5Ts4gvL4YHFp7tKOs/S7OcXIHIpP5LW0+7twbqW7a8YYrtbTrdnP2SjUCjqR7G7iZSRPNgCYbbb3
Yr5GNey4KRirZsVuBnIB9Vq0MkklE6O3UFXSBhkDGp7TPB2AIpGspt4oTMZBRDJwYDZ/ajOANF5N
PVL1y3HohKxkklk+XpiP7BJBsdVq2fLzg7en0K6yCq2/RUQu9vCoZrJ1czzkdW0FU80NtKkFNaFr
ziMeyC26efXRV4HC4zKZUIpX6Xiyhl1Jq+Bqc1Q7T4E+6Z1Ulh5tWzZX1p14qUxV0hzFoEq+RWIg
kxb5whxO2a3wK8BbEW/mIQ2n1QEQOoc/Z3Bmw2NYJQksCYZLhvUgiQsTKaBNZYru7a2dfe9gLYJY
1jR6DN6qUBPWKCl79KuTaJZqGdnviBibVJAatD656YUzjenths2q3t1e/Gv9O0HdR1wCDzc07yaj
rBxxcFTPVqogU+n8B4G8lLrMwq+nHmCNQN4v8WDFEMOFhx1rhmwCXSztma9TipAF3+oX+UCxxcw2
chz6YoqBMyxbAfuNOa+yAw7iavqjxyZbjxsTQ0GXscGyxq1xX/o6usdkDOw6VwLCxvkd2V+K65Po
+1Ir2W445aCzkmtp17gre9qMBNFtGoOonVGdnK93roOmKmZv+ZeVYlmbL1wNh+KAQMZd7eG623/F
vEAQOl200YUyW7YvT7WSev8H40boQ8yQ+pm5HUMT4WJrs3K6lZqR3MtrdIYF2gFfFX1XZHHp1pnD
yH6r6jxlo3qYDRWI4RRHiAvzbBeJIbEJV4nfnZ5Og7Go4BYKLyOeyEoFwFFbd1N52IL7qf+RMKnV
HH+KH0vqU1ut5oTxA/JJLHKN2Khc/BkwX+uab2xIiWrJ4qzKrwIHKCKmaySvmTHC9iQ4vpaSWzDX
9+QlFme4s64wEmCso5TZhc9/nPBDpnWvVb1MhZkmNcKUR/H0StnCCjNyxr1g3UnjqwiX4iDPN3ic
/LGMT2EiI//HsprntHBD2RvqoyBG3SS5a81gO6Kq9+6jvy97wfT8+jS8ZinMptwsYm1ZFzc7cjTh
3zkfQKoHF9wCIZYdqm5ieG4cxFIV+BAo81f50kyvCB1TLDL8bVZa06qVCWwrBJ1pX80Xe/f7onGL
93OZXze/je6R7n22yog6QrHf+zinWqwcN04NuTwmo5dScAWNlPQpvpNd4y+blrbdLeZL8P8DGt+h
1ubS3PGXzmjbXDj7w/gtWeFW93BIB/jZsjNJN37MqdeBeeaCInWIxFFt/+1YboownMGPkBPIlPJ9
E3Gba+PpMZFcHWmstxdZicMbiUrwt3/5ezNG3pvHidQogH6b5xJ0DzzcuLLK/LAej5yXdytsYFjV
2r3aLdt4sTstRpbMhfUWC4etZSjb6hyk5326vaHMZ0dVBsG7fYfg7sY8/cxEYXPbgSAM1yiBciBy
hmMFTomynAPiljbwEgjr842W7bdWmgEDoQkf6JE59OTNQRp48FR/lvESClPZL0BNPD6z7eYdMx5A
Vry39EtHSk2XfRzUbBpTC1kFqzbOt0BNPiawqzRww6GU0hk4XwV30m9Ryz9BBVdNuO/gMYaCKXHn
CHFw2bn8tgOUUZ8rQrhZRYjKOQDN/ZFQBYIgmvQSTn0jOW4obTvPwAYUd4h7U7/xRXnr0Tt8Gg7k
SNQEMux/ral+8gr51LrlPNGLSKsse7+14FXnAxB8vs7no/Wn9PLESAEyafHoTIhM+VW9uH3UZ5ss
QtRCfrOOagM8SIcVfhvrD3RHy2z8NC0xTXCw0Ptw3b8nunOziOkUcDJpN/Z/5XMZ2JBpCw95l8/O
/djU9DNzkEpnLPQyReHT75dNpbVjsZp1I25EP78Qd5hq0plWI+7KQHxltMAopD7wGYYGtKFXdXYP
hwosRb6UVH6lWcBbEcakiCtbG6ZWy8bGeXdOG90/g1RTdQaUD34cczafENXAd5ZMIEqZ
`protect end_protected
