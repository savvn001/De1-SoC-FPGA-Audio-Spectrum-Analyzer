��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl�"u�6|F�jJ%
Aڣw��};�9�D��[��yKה�2O u�s��4/S��)�r�R���Tkgo�R۩~����j��l� D��5���+�HR�?/��.Fn4R�l��3��8e@��S��� %2�|(�Sʠ���|5�~��@�9��`��Zq���:ٍ_�_[e�kh�pDN��<(�������
���![��}���>�`P��{7��x}n!���c��������p��v��+Q��0��}�a7,a�TJ�w*D�;yvX��b|Yw�n�0�!��ӣ�L�_�_�<�j,W��1�P��"�"��~43�������0����������&W�{�E��Om�烲2�Q>m~��� h�m�5Ov�&L\����Wv!��=eenق�C��`��~Ӵ}?�����f(����-��g䒒�	�F��+OR�t�O�'f����S�BDi�,H�e�NY�-j��W�����+�e�s�)> :'IT$������1Z�-�F!ETZ����^��,�V9���S|����r
��H���K5�ե��&��}��C\�:��LN����e�;�ӛ��{�9�&�pJ>jpJ��Ěw��u/�g?�.�hIg
������bڗ��B@|��[�$/�݌��n8R60BS��I���o];�G��;
V�)� T�J'���g�MV��%U~��30��X
�}���<��'Z � �i�B�!>4�^j�ٕ��-W?�Wx�ǻ�%>�z�S>���X?���F�'�0+��k^Icַ��-�6�	z�A��e?&$��ó������I!�I�ri�E��3b�<�Tk�\�\:'�-XZc��:��xLR���P���`wa�f)�_� ?��יj�� �*4�?���r���y�.* ���Uf�-����h+쒦�i"��NG�i,Od��h��4eИ�U�{Ph_,�z��k����p�33����&���x���Rr�������Ch���k-�"���R3�$��ۼ�];QÏ. S�~m�08���1�4M ��k۰�6>�ÕT4��y�D"]���3����tꤔ�!���7M�}o���^��� ����	2���\��rԹwqhަx{��鍔��}��vPD���
}p�gI����}��ƣ�#{��CfT͚\�[A�*��nD��q��ѲRb��Q��6�ۚ�^�Ytj����J;--/�?�ğN*�JQ2��q1�_\8pytD����薉^�4�b��$��dl������O�<�]�S�����#x�F#q�N�z�Md�����>���~4�Q���[�:Q������q��z8�ތ�95m���B���W��@:U�R#����$�ػ/Ť��+�ٺ�a�pڻ�Z�K�h1j��;�#G�gwOƠ���Z<C��-���e����qT���K��g_E/S���a�=F��H�s��6�;���ٗ攍��U�i�a��0�����:C'�f������l����({s����~n�n�.�{����u%�p�I�t�/q��,���rQkBڻ��?|��V��V6ho��J'r4�M��?��so��wbްq��傷�y��/|�R�@��,�b���1�a�����;:E��M^~#�Z|�2ߓ��C؉�/L�߹�]a=�SR"{2Y�{A��V��my-B�l�
������P1q�:mHށ��?�Y�z]�-)�u?=��p��n�����+��z	��]�����	����=������L��!\�І�n�.)<ұ�P��n�'�씃O���fT�w�s�?	�oE�=>�"s=ʳ�S �v�:���U�su����ܱ�1��A-Yne�N ��+	�����	!��f��(`ܻ;�r��՟~8e�<��T����E	��Y"|�e�Y�;������	�&Qj�tc#���Q��k^�N>�#��$|�����=�@���}�Y��º�MGƠ�J��(����=���YsAw��''��g��%y��Z�36Q[�>�U�)��P��1��1���q���ƽ7r/A��Y��w�7�E�ٚ������ޭx�Z����ٙ�ay�����}jHb���G�l�ˑ��hG��M�M�����N�2�#`�	֬��n$a|s�x����ه�8$�̫
!�Sl�':�s|JZ]C��4U�g�/b��9�W�(�����&�TCp哏�9�B�u��ʖ��#��%�q$�����p�΍
��?5:Չm���-���mX�=W���YM߱�F�h��E���j���{�e�ذܠ�Y�QTy��
l̶��T��֥���t�D	2��pDH�f���j��6�xWڕ���6[��̂�L}�O�"&���H����.��7"��MI��g~^P�{z�zx���,�UGM|v��:�zouh���2��	�+ac�h�v��a����R5�h��">K߆�X=@�wT���hi�c����$�c���g5����2D���x����33�k�1N�`�m�u�}ϟ㍥)��b�=>�1��Lܧ�&�Ɔ��rs�o�@9�.53�(4���8n�;nAc�5��
�τvȏ�y�ȭ�r-��)�e���pkC���WB���
����V����6�|�ԱV�YpT��G��V3�?���M�V�Y *��Z�9>5�����
�yL��5�eS�������:'ތ�LH�����mm��@.P�ioYa�J��C|��f &pM����lH�K�_�!H7�?2���pC��|�<"��?k�2�j=R�e�O!�`����z���r��̬��7𱽹��`2 �8$~A-/�(v��1ü���(�����n�N2����/���������L�;�7P��5���q��%d��=���w1O0���Y�A�6�)��2�oc	�9;�le�� uPR��E�ѧ��a�_�g�����;�g1�k߃P��2i*�u���Q���0���u�]#В��1��a\�Fd3w�gT?�Rp�"d����3��(�-`��6h[?7�+��L�
ۿp���'թ_�nII�cx���<O�ch�W��R5�yN��K���B:�M����	oR��2�=��Kf�B,�@E,���EV����і��k�����3b�ٹ<K�D�3���_�xI	V� 5��X{��N��]]	�X���Î��#=��a�̷�}�+L(�G=X>���*�u���8;�7Z��'(ʭ����y�� B��HӾ[��^U�wm����UO@�Hj����o����D�f@>�E/Yz�4�x�׏��������@ ��2�{)We*ɖK���59�i�G=d�9+��Ke��H9�;k�o��@;�'Pf��X���;�V�(&�UFL� -�(!����5������8M!���pۂ9+��GP���O\��@��}iX��Q�[;%Uy{#.��߿�N*���e���	������Σ	�%Y�*�!���؄�$�E�)�ҁ�	F�?���q�"��$=}p���Y�����D���\g��B.�:Y1V�U���8�Q���N��i>x֨t?v�/�eB]�[�Ga�X�O��	�8pJP_J�&��˅�H{�,C=se��03�^_�V���J���m#��5�?'YR)���n��:�S����l��x$�+b5݃{)��|Ml���w�-��bwQ~.���?�}���_����`��O+:}�z��G��By	��3���,8��B�F���cz�$ngη�%���*���`ʩ���D����/[�$'b��ˤ�1��Chl{�v�Ǫ��p�0>X"�2��C����TA��;�t�7��&��uDa޳�^�����F�wz}k�"2�Sn�VfFJr�����SfL�ةP>"��n����t}O�d��Oj��)Ꜽ���ُ0f�mۺio�U;�aX����lπ�B�ƣ�w�x�m�0������W
�HD�r}9�,���b~,�$	~��7�;h�T���L:�N���WY����f�Z�f+��-�(W��Jn��/Vz�V2���D8�����P_`�\b��V��;~�ՉG���� ���_�,5)�Ruuķ�~��Dz��q9Sc�u�*�2���>YH@d&u�E���9?�7Z�yO�n�A1��X�fb�E�R�T��T�E��nD	S$�'���o��ńaH��Y��Qr��X��*��+�"Z�xw�L�݌8$gn�eŦ�[��F%f��h���el��b�LyͲ�2joH9�
T�ƿA����Ia��+=�CF�L�{И�PY�*ov*D�ƈ�)xԪ���a�H��eZ�g�a{�����t��.�尿M�)U+�n��Dc'��z�������屑���i�v��:jn/N��p9�yn�5'�wc�d6}Ns��:�ke�ǲ�H����NU���Dg$��B��	�,/���2,��6�X^=��WO�Q��d�&>���n�#��{��cs����we�ݢ�5�*]To#O������6L&��v�n1�O�XGֲ~z�h*�����L�u�r����nd�3[��� IF�9��FN��^Y�DE�O5�`��FN���a�fN0�xL�c�[�	��\��^���(�r��k\�9V��آ��1���x�MJ�>y؉�E+�q��e�"E���j���U�m�ݛD�:s*������5[���� ��N����o+�Y�����w���ɉe<\j!�zaxd��Ht�o�c��j2������8��#p�:w�G)��K�JNB�xd㬍���S�}D&�C��@\�� �kXh���S'U	΀1��)���MF� j�w���.ּ���P��9���*��=�[t���^���E��Kބؿ/t�^�<"�Z>�weV|N܄��B���`�^�2��2�uz8E����_A�ϭ��7��d�t���(Y׮�J]�:�IHY��-�䄖��n��֐7��g�r�g+�է$E($���~�~�>���$��-��=���N��H�8I֚'������'�HSv@���e�u�A��޳E����y���r�xO�"D����������U��)���׋�>�J���u�Y
���)����3�,5z��^&Q.?*��:%wz���{h����It�g9�B�ˇ|�^��?l�qGX+����C g���~ 4������ō
��Q�e�~�4����1w��c��dJֲ�1U*=:6h.���և�v��Y`X~�=+�78yK��޳�:�ɤ<[��5���Z��=��7�Ȯ���y7�Ղ�:��8p���U-ད�K	����#��X�Z�9���O}S� g�-3>��@��z�E��{��yT[s2.\�nųZ��5!���Z�YV�$�B�U�{v�s�)���nrUH[q�3������ύ�=^³P�^e��&X<J��E 3A�f%)�,tN�B�p��2ܩ��Ĩ)XDr�;!�qɏ_�T�kU���E��󧹤A�Y���h�J�p��o�$��R��1��K]�o��m��NIW9��2����A�Ǐ8��)�zF���8̃� Z%��)/)�q�O{�'�d��sd	$���EJ-���q�ɴ� n��d���$�9{�x����T��7^H�pO	x��h� i}횬�0R����TeE]�ީ�.�����WNj�I}����{#�3�1.`l�]3�ߓaEc����6tm�;���C8ؽ-������dt���K��YYG�1����%�Dc�����z���oz\��8�K��q�}�T�Bˆ�W�����2�x�#6�X���Pf�\gt�R���8aMGhW��*��Wp���|,�Y��
Q�f��T�������\P���h32�nY��'�&i8�y>lV�����oߜ-J4ds�f�J�E:'����y�rC�e��SΎkT�����-���U4�Q?��h$<�I�"�w��e��7��C5.T�D!������)]}S������.5{rL^['VL����y��.D'���':/9����v����a�[���{"�LY�:E�E&�X��Y���8=FҬ謹��ݕ�_���+������~X�-G8FF7�s��������C%�����d�}"�ĭ�Y1��|6�B�|�aq�o{j�k�`6'{^Nwʞ�\-O-9����4������"IC5�t���=�F���t����{�X1���~�d��b��5��ݯ���p���XY�q��Z�.��@��'6^�FYv|�E���d�|������D˅2���/�bE��ٷ�9��My[�{ݽ� .� ���#s 5I����q�u�'ց��r�o��/��?8Q�bO,��Z�.4f�m������Ll\�~d���d=0[�5�����5�,0���4�d`�>ƪ�
�	��/P��f�>�:��-��q(c�����NaY	���^��Y�f"�gN��@���+Z��?��,0&���ZU_tz�Hr�4�rn�[�*�~g7:����#}*7ݩ-�ĞZM$L�*c�98��6�g`h�W徔���!�����bo~�t6����()�&;�S�Ȝ sG
��#EПSs�t5��!v������DWt�^��ʯ�i�=�$�e��Tv �j<��P�S�!7v�.*S�G�pZ{�v��΃����f+Xs�������t6"�B{�k���:�<WH�e��4��=т1��#�g�:���ۂ�H�r�[!��<�VS���s;r�/hLuŚ���2à�l�I[��u߸�$w��{	D3Y�ذW���*��O�j�Ѕ#�fp������'�j/�%��z������=��#�GR�AR Vx�uR�n.la�nO��}P�z]�,b�>Z��b�Z�D�ݝ0=n��`�>4��@���`}�`[6�-CB��~~�?����s��۸��ZJ-�8��ΰ�iݢ�Vwe�)����bgt��Et�q@�-h��V%u��=����>жE�е�L�e��|�A�j�s=���R�V��`L��=vr�ZR�Xǝ�~������n�F�g̵�je�FܹcGޗ: y����̂�jx���TY�|��1�Y/�!|� e�(3���Ps
�4��OQ.-�l��@7�q��Fa�S�=��rQ&��A����ҍ��y�`��[�Ÿ�o�02#����i)�gsO�4I�Hï2^��je�ɂ�~q�i��lBd5�:DT,ݮH�ߒxt`+�W�	�%VMך	$[=�ٵYj���|^�~�"�L�P��������9t"�$[rR�EU����́��m����!����������QE.����;�b�cᖬ��c� �	sx�$:A'�����~�����@B���8��k��e�3���V�y����*����V?e҅��fD�����f؀Zwoh�L�c���s�P�{�'g�./���Sa�a��P�,ޘO�ႂ�\���A�jg�NK�B-��5��~gI�F�������+�ȇ�&�6�o�8�~}�S�@�����SaF@*dK�q��\���5�GĎ�����\ޫ�����L��~������H   �惲�}!|���^0ý�1yE1��K�j	a�w*��#��!͋����a����0e�iIb�4l�v���Q-Р�9�͔!wi��_0v�p���4f�ɺ�X]�Շ؍3���2! �����,'�&�H� [�|rWВ��y�����HG���L�'\�xIf�S�⫲C��Y��O.�z#rL�I8��w���RX���1���JE�!�=J�C87Nn�T�%Q�b�H��Q�����l�(7���X�~8��`�)ˢrNl�nj���$M=��3��LI|.��#;���W�����f��缲��Q]_�"T�N��y�V��s�zY����5Ӹ�9�?$_�H;����4;�HV������7��&\��qM�×&Ƥ㟤��{����qoL����R���U@��w<|�EKz�=�	�*�%�3�Z���#�
f��{��7W�;Z�����Cҝ�$xO@�2���֞���4zB�I��v�#�ǺH�� ����u �z[�#��]'���WF;����K3����,�}`t��0�YV�C���N��SrLbv�2�RUلYŶ��2�poF�$�̚	�^�1�6M��q��(,U����CI"���h�0z�h���d<��֥?��������cr�'C��K�e�v�~F�{��F++ͼto']ɓl��Z��@�����f��˶3�,u@Ԃ��E��������Xl}%eR�{��R	$��kGaED��:CO�Za���MV��I���Z/��4�*���B�r5fa���C��YB�˓��zڛ�JM�ä_�"����^Z����5F�w_�Hsl9C�i� ��q]E��s�Z��j��P�Wp��.��͌�/����{���T/�؀�$L)lG�������
F�+&xe�+�%���h��p��'fw ��l8�\P� ��e7s��L{k�;�Z�\ �������C��5{fA��<Jg+��]�y�Y�UV���|��������"��0�?��!������W}�Z�~���{ܒh��	���=u��S��ɭI����\6�q`� ��V[�=@��}�������&F�W�t�\���~as(0C���9�u%�-R��y����È���42���=7v�[���]�
^��Jj�p!N}��Q�fyi�8
Q��~�jꈻ��NS!�saq�%���&i�K���Q�K�F`�nU�D��W��(�$�a�*ndMf����)�	Eɥ�pY3h�<M�СW�A͊���f?�{�����`H��S��}^�J�Z�2}w#o����L�r	�oO��j@,�=�S����7e�/�+�ʹW���
��2�N�����1+�d��� ��U^�Vh�a߲�����fk+j5�&�$�E�D%;!K����x��bgKм��	�,��51�]��t>�ԚLd�����J��4o�H�O���#����.�3Ņs25w��=z�ެ}�!O�j1��dQB���35;d_�Ν�9N�v�\��Ŝڨ?�3����5jb�����'�WR4.qg��OӋ�A�� �m�hg�[fV���
�z(����F�B�}z�/���A<�<mӱ�Nb_�N��|e��j��JQ��ѳ�T���E;��_5�!۠���iX����Q�Ҋ��ݯ��A�ĝ���Kx��!��#\,=�?Jdl ��jn&�k�����@[l��[��P�V��~�B�W2��A��DS�an[`,q�$��ۼh嵿]3�?ƌߖ+�D�������8��3���Yݤ��vQ�/�\������o�)C���1�i���2'�����BÙ�:'K:D]�(��O�v��.�^F�d��S�B�h귪U@5�/��D	x�©���ׅY�~]���̦;���O�j|k�����gQ6�jv�W���hlkh�U��Ѭ#^G�c��*$~Fh�#��9F�O[� �7�:]2�Z���"uBlȿ��{�~;��;��θ��K	���q�ߍ
U�
,Jn��� 	�UP0P�h�G��`�SH��#<���4fi��o!4�D�O;Ҋ����zv��e6�<���MaYL�43:g3v\������;�����tWm�B%V�5��9��d�=�|�c�2�?�i`�R��E��z�\��tɟ�pq�Q_3��x�)I[ɒc�Q�t����R���E��b�纭����B�(ʹ��ppS���_bĆ�^�G������Tyu� �d�E
eQ3,t�э�գ���*���Ѓ�~��9��g�$:�8��^́���6�A��T�;�{"e*�0��VĀ��q��a�T�SDO��&�(w��>�ٝ�\�����5�GN��l&_~�܊ٳ��|R��z2��bZib�㫝���ʠ;+�;\/��n�Ղ2��q������'sy� �o#7�ݫ,��Ms�t�;8�ˡh���~�*A��\*B�C�Cg��;�fR9�?b�U�	��N�F�`nۍ�^���PA��$�H�Cz��i]�M����oP��gS8����f�#D�����Co�NnS�m��5�t.��p���)�i���N4�|�Z�⧄vѡQ!�"d�p<i�Q����%����A]�g���z>���=j	����F�B��/`3sq��[^��Lֽ+=)���w;�Kż;�l/����k7��0Zx���.�8��t'�O�[�^@FyP�0�����B����K�@P�LwՎ����G����t�,�r��z�<s}�^��XP�i��'Ě�7���q"�����R�M�)�_Pt�,��n6E��=\"�z%3E#<eP7Iqq�y��7G,/Sq*�t�Q�s}����[K-��T��=�*~�C��U���W���+h� ��Y�8��%�/�ъ�a�{���m�	Q*1�N��6q;��_�$(RW&��Fɿ���:C~+Lոs,��c���� �T�H�?�v�{O&?	��.y��ɠ�.�{�<<�k����j���k�T#��ܾ�Q�8�=_%�j���!���܉k����)���&>5bQp�Y�]p���2�_X5�R
�d�a膮����>Χc	�f�z��	݅��l��-��O8�.X�h�{;����O�����	�*���E��<��W��X$KaƷ�CE���A`�ʹs����W�Z/C�G=m�?�Y�!Hz��FjrÑ�&i:o��hK"\���3}̙�ZZ|����w1Ű}��6U��rj�e��W�a���N�(��lRl���*�E����������#)�I8��/���2������v�O
�����+\��?{Q'&-3��{�W����^lD����\1�C�D�a�Q�J�ZZ����HY� �^?K�2�a��[%�0��p�C�^M�U{oQ��8A��b���a<���؝�+9F1K�e�|�!�����d���x#�B�LСy]M�WCN� ���;o�p��5��e�.�q���<N�f
m�T
"rx�m��,u�^�D�3s�B����R����^��cy��`7�`����X��b֞�DP���~��")p�F�![�W�ruw�rjc-��8��N5=�>�PYd��-�a5!s�gZ�/�dn�|�ϗ�#�'sW=�.� 6�4:s9:]I�ٝa�#��u��l�(6#se5�f�R&���C��]����*�n8����]t J|��eEQm2��"�R����ًCbbqr�G`8(w˴�k���0���C�
8/ȗ��
a��FmC��&ӯD9����Dt3�H4?�xy���[�{�����ᴠ(�K�s� J���T��'(-�F5`�x��M����H=Gh?�Ϡ\�Mt�z�3��/o��J�T��K�<)I�X,;�}[�����T�r��8��S�r��v��`Mxt��Ձ�Jk�O@��D��s�9�6^��j\��n��ɍ���Xү�֋5)�q�9���EHN��#����lF�
C����/����c�!�G��M�92cb��&� C�	��Q�����c�vXɃ�2N�]������4pj�����+�H�X����P�+ZhF�h���]���4|4�X���H�;n�ZB�Ŵ�DFE��Peܗ���T;m��j�����X�P�y�^w��ap]t�?�	1��qp�8fB5��[���|ӥ�n�"s\N�� (���}/���d��`F�L��/
��z�/����1 M%�]�(�K�4�^�L�e�-g&����u����^��D&l��T=�۬��S]�� �h���Z��< ��D��&�J�����$"�
��,��u�ZV �YO���f�&��|��/y�$���Ρ4�D���#TQ�� *�/��w�љ��d4�7��|7���o�0�Z���4�t�(|t1��&�(k�VI���M9���"�����8tk�̀y������l��Z���m-O��R���։q�km	Q�O�E�Q%�E����(�C4�[�?�[$sWKD-7��~��0va���,����{L����bw��{��`��T���l���iE���C��I��a�e�lN�*fN/п^��!)��̏�۞�#MIse�����t�+�`��st���JM�a����35��N&E���Ӱ�s�!��*�#x����
i�
o4��id�/8qg���+
��TT<_Ȝ�G�>j~7��e����!�[9O�T�ʄ�el�P	,u�m~v�rb��XBw���y\;���ٌ}-9~�J��(�P	Θ�7J�;�}}b��s�9��7!�Ք����,�s2���k[o2~��kL�Y*��/BG��a�1��s���l"Җ����EZ:�����4ߌ�U�aa�>4�F���i6[[�αt�h��Y�)C�7	42/y-)/;6y������,i���=��ZmDΝ�z���YF��Z�"m'LD��������V��1�A�^�:f�#����2���q��ٲ�@���,�7W;���M	0�p1�'�;ӡt�a��D����8g�� �`q��{@|��A��AZ�Qm:?0o �uo�]v�*]� �#3;���X�y{�ڝ�衯�,�����S�4|2O��|͆�
-s�����C��g&B�3���Y�+o	qF�͡K�r�_X5Wnӥ�n�CÓ�Au�ٌ3��f��H�X1�]z�	�?TP��
F��[p���>��(p�|9HX������"g݆�`)�����,uxf�s�o������/��C�j�
�g@y6j$�"(��&�y���qI��	va�	h�s[�R�3ԇg��)i�I(� /��!�sAt��PJJ���>}Tqt(��N�5zO7j�j�)��F����hS��Y�W��q呞+��I���o�Dw�mV<gl���6�WO�أj��^��;�.T/�K{�#÷�!4�7�-�a�B'�V� 7� ��o�h��,�����vj�����m�!GF�������Y`ۙ6U����Vn�X����)��σH/�E
g���t��+��b�+]��*0=��y�Z}���d
����)��~!���>�x�?���@yC(\��d�E���NM�ۣ� C��h� <'p�97�������d�[oʡ:・�Ƒ<5ލF�e�?&��i��`�S]#�/�v��)C @�����m���u�λ�?�2�n
�sa}�YW��k���"�3H0C̈́�`0�$|���T��|=1'�l/���;��@��t���ʹ��@X���b^>�G�R�`re<���XA"��;�i�^i�HU��;\/�%J��T]Ls�<��a�"�B?:ʚ�lx���4q�҅~�����%��Fg���nM��.�r7����c�g������E \ ���
Y� )8�'z�r�Px���O��&h����:7,��eC��l��[)�:�z�9�غ+��o&�=Ʒ��S�Շ���[k���SO�3-t�!К��N�Q%'�%RǸ*�?&$.`A�P< �"�K��p�cp�_)"+�4D��N��,���������0��m �S0�A�k��M������Q��YFI�&&���_�>��t ��۱���Bm����=,��K�Y��-'{O�>��3�Vt#�R!�%�I�!�T��ndtHu���9�Feh���]oV�e"�
�-����+<Hb���l��(�N�c�x�?�dh�fJO�J��Nĩ�%��u��1u����4��g��
�5��Ty��@�k��J��ʼ�D]��'I.:�V\b\WwH*O���.��΁���X��a�ţ�@��d>�J���@(�?�����f��S�w�ri	o��xMe�51|\t��� u%o.[3��|o��r3������D����'��*�%d��{� ��@����U�����q�m��e4��ޢO��S��mq�����]�爂�@��A��
���[������}rp��bǑZktJ�r�~�K_�.c�xw�˚�J#B�MH�
��֓I����>X�c�����r��w��:,VH�F����c���PiM�s���o�{�i��A����[k��F!:�$JYHOj(��An��� ��{!����M��y��p��E
+��-�Ǝ�t�&��p*Vl��cO�Gp�K>�d�,��n���s1��O���$�ӿ�a���	{�R����t5v���Б��]d�y����o�P�����Yb���	E���Z;�ʐc���X�ڨ'2 �oM�1�4
Ɓ�F��zH-�u�kn�HJ�@��
������`�|$ �\ք4f������#�9���+��'���j����<���V6�V�_.A[��oI��۷�#G�[;	�N�Q�H���Jv��eT�!x����1+�����8�k2VO���h�y���rn�L�A ܲ�1�p��;W�(^���q��:I�fc��-	-����Q��8�e\rlm�1jq��`f=���I��߃feo���s���&�S�����PA^��̱�~��o%qD�#CuD:w�9	�����H"�1��T����ʄW��l/�Ƀ�S�0��	A�ѵ���^�H@=��9:�gA��V)��_�ĉ_R�8=ü�?�O^S��!��� {[������I���e��W�*�x�aQڢ���#`45/�����k��)v6?��z'n��:�^a]`Z�>6���=Jј(%�B��Wqr�!�y5�p��v�ƺE7���cO��%iB�R p�����M��4��6e��|)<=ב�[� TL�#"��9q_$l�m�5'�.���.��-4᳗e�W��^rl��-=�c�<%}�������̐x{�<�A.s*��/)a��,�g�s7W��qע���ʼ1#ynSNS��D��&�D�$xB22�Dx�m�Kuuꡟ���]�XL���Pښ˩���xu_��EDx���y:<f0k��.]aa��,̷L�9�J�Z�ɀ�m6�
�ܻ&��x<��G�K0���f�B��E�<��,`��ɡ�fV���w	zu4��X�c.�������Y<n��5O�sl~�s��S�(;��,�����=.���7[h��#'}��Q���>�t�?�Ƶ���/ߦ���wv�Hi��b���L��Ń����1]Gr�y����:"]{ŁU�l*/�m��_#+H4����� ����ap�&pm��<zd�j-��Ƭ��(�F�ԋH�~X{��4�{��4�H�Q\���p.Sm3v��ڏ/1�ߊ��t����7��d�������U�
ɕN%
���s�ľ���8Y%F��c�̸Jr�aE�}�����<|��k��(?���
�@���'�N�y9��/w��n"ڻ��${�z�>���P�	6O�ז\v8@Fݧ�IJom7���%�V���������m+�g�1��]��aÎ7�(��%0�g�[ V8�`s���e�c�ޘʡ��]f9�6hʍ�2]���R��2D��{���M��r��N����<�EG�W �$*`}Kf-�P>��8�q�)HԢ6�����1�,ߕW=Gz@̣NJ�f^� ������8��Ѕoa�0Go��$'��#��m��U87�q���V�P}7-�ӑ�A
�|�a����b�"��<���z�zxk��-�|��\ŏK�"�W�h ;usTY�_���t�^Шw~Y�����?W ��ʵ:�[���_��t�+��c��Jk����7���0��~q�;��/5�x~c�Zi\�*�#gF͇��z�$��7"�XF����B��j�r}'�M� W<ؚ�Yt��E)��M�J�bQ�2�qq�I��=��p��L��=i;���%�v�vH��'��Y&��O�s|Q��V��{NI"�*��	���Z�Y��Y��
|Q�զ:eW�0�Cv4{�r�֣��OŬ�D���m�m@���J}Ș<����KYz�'$�U�f����`���>��U�z���|�T�9��O�5�z��k,�Me��PF�>��
����R`H]���Bݭ��丑�!{���X����D���W��Oi��A�g�p����ŀ����E�=�Ԫ��S�����ط�y���x��ɤ0n2A�=[�;���LX�e�[�^�$?p-�Zȕ�	ƿ��c�����-�h6�f�碜.���V�Rb����^[9��k�xlz4���ܯ�?��x�>��M<m2���D��P�un.�V���M��k�d���?�cwsH}�H��0�X������ƴB<�p���A%�[�������T���'����	�������o!��#e����j���.M����@9T�G��<�V	����=�<Sf��z_��8k���?�^�����2&� @[����۾�㎖T9l��NE{��ڒ.Ej�噂�^1�5��	���,i:������!C�����Z�abX�I�e&���.����?�$�>hn��_�z�o�T��ْܻ�،�����*�I�� �K�YSj<�n�K�����nU�~W_,0�ÕR�m+���xcz�/_��Mz3q��N��T�;533�[8ј���`�A�UQ6�,@M�]gc�Ց��X?}�폤�6��2f4�*>7�-����vk0_�o.j�\��y
RS����W��!?��aBּ�!8�����n?("̶�%h@V��HB��wwL���7�!�|�Vo�5q��(g� ������/�b�x�Z�.�IՂ���%��)MJ�K#��/�V&~�Ng��8�~�#w��w���*a=7-�Q��طj��b6�61r�㎳����ۉ	"�Z�˥�z��Ʀ�gI;�A�ʓO'.��dl|
%�H �P2�|�H>�?!N�0yU��lO����7��بg���k��=�(9���.]A8H�5�62N�4�u~��W�5����狮3��3�+y�e���h�=$�zɳ���Y�^_Z)�m�|hk�[:��K�Qw4d�|Cu��z��=5�<ނ��5>�1��._������4�l�4��#Ul��g���A3�	V:(dk��q�WZ�ή��ڔ^+�@�u.؉�&�Ū�E���>���Tƞ����۠�\t���U�SP�U�N"ll�"��;3�Ȉ	gL3/A�f��C��Ni*�`*�i����*Y�Y���6�g�/3T�+����[�S��Gb�6�p���x]���`�%�� ���W�0�P��X�%cl���WMkی�����9�a�>���T��#d�*�掺4" �H3���|&��~�d[/�l]g�'��Z�k��-	��"��S�j��}	sNq���M�������!h��S�!�1b:N|c�vLQz�8�O'�7����s�R^�$�dDL�d&��ʕ�~�Q�P�|<�1��!"�RM�Dl�e��^'�Y�E�߄	�*k��V(}��@�x�!xK�������J$i� �We���pns� E(9-�5��t1f~�
��˓�k#Y!���[AyV�S�'&ߋ9�l�<ϰ�ß<��������p<����M48��`��.i�O:V`y�~޵��z���g�L�	o��|D!1�@�E�(~�bF��VV��E����l!x�6�fͽ����vM�Pd�f�!Vn&�a��f�| ;V�'%���C9�'L ��M����qQV��+oe�I����-���|�������T�o��>�*s?5Xh�ي�x-ȗ1������Q΁�|ZCJE�MZ��l[Hl��\��P��ՊNb	�&�,K�(T��`&�pP��}���v�B�j��-�^�P�"}P�S5d���[\�|�1�q�4����IT���zf@,aR����R!hG;3��F:k��!)ut�6�"��t�L��7��bt^���U
C��r�/��y�d�v{�֬���n�����c3)5;�x�K���a�`)�1	��Ү��o�����,��/2�A]h���J�'�1���M#����$���R)Ɣڸ���]�o���"g"2�A5c�JSQ-A!y��-pk��b�w�ms���~�����i�.j���.P�qk�Ք�4��J�ۄƧT���0�M;3����H�W #T�a����[$Л�`��:�8B��*���G���ڿQN�z�[��|���tS����N�@�QY�D�eJSLr����T3:�<M^��o�a�nu�_b���IP��ʗ��WxU��Af���A�d�)Dj�\��[�^(��S�������h���K{+����U���(���݃����m������Ɖ�t��Y�~Ћ;�}�����I�o߽b�;��O{���Ba���t&!d�hc��(㒑���Jr�NҲD	�Z�E$� �wɷA��5���y�}���2�Z�!_��ҡ .�0W!�^���$�	SX����עj�tw�����'#x"M*5���&�#N<��쑜<��?W��դ>�r@_M����$�Yr��b��}gt&'�_ԒQd3�A�'��[�:���?='���>�)@�8���X��N�}p�ݫnJ�-ү?�V8{��ՠ��S��g�FP]P�ϰr��ؔ���06���E6�\��wᕜ�B��;A�][6$�����<�0�th��a� ��r�/�.-f�4��p��RS 5#aS[�f�2g17�c��2�E���$ɸw��l�o\�`�'/_�pw�C������pCüњyH?�[�y���������F�����Ȃ��P�5s�Cʨ�ms�dN��wx��%���"�5�q	��VԘLƨ��K��[Vܦ�l��s�z�;-�	pb��k8&�r�cQAt6�wJ���v����is���B{�ܡ�}bA��zKiǫ�t���Syd2�n\��1��႙�)W$�d�6K6�=�l��z�V� ���ƪD^6���n��_���vݾ6���*��� �fI.������ר?����R�(1e�#'^b$�I�ZS�c,
Զ<&�#�ބ�^5 4I��l)�g�mc�@�<��2d������������E�%�/���?W�;��3W�FX���]��.�)��xV��I@�y͑ʺ2��Q5|��7��}&=�8K�e��?��ĶC�[e��֍�֕i�5�{
K:�����z��1B�ʒ�JL�jj.��h��}��q��2����,���j;�@S�z�����R$:o�R��7����`�rt��s�!�4&�
o���)U��@�l��￣��h�����B#+>6J&s�ΩO�A S���bz�be������O,�!.#��ĎGj���C�'����/���A΃�]����-9#�1.A%���� 	��n��}D.����`��I:�@�A������A4�#��ͪB���&{����D`�ogž�����-Q�}��|P[ͦE.bI@������r97���� ��c���<FBL�1�K���t|�2�����!������6Ǔ�n��t?\	W���ŉ�q�v�M-����v0�
�̦U��!c�Tx���c�t}�t�2S�o#k%�2�l��:�z���,Ƣ�n�Z�w��j� ��;�=�� ���� Ey����5�vV!��r6<�ů��+�[��%x�w�2����
&�Ո��%?��.]�ۊQ�
���٩<���W�?����Aa�̎���ijaB�(*7�_��c��mi�� �������wVI��ȖEOӢ����`�.�l��D�iMD?��؄�����o�ɨ8�;ZI�,�N�ġE9�����7�י�X�Rv��NR���D�>S)�|<ܑ4Q�x��2��t�%�ê��҄��v�P��Q�{{Mn|L8� ���`Ռ�d|N,��p�Ũ,���g������vKU�#wZo���Q.,.����m�����~ڻ�G]�6�M�\�$��������j�>�q~ɧ���;?�������`�M�b�<�-�I�I�i�8�**��F��R��	��?�Z|��C���"	b��c]��p�[�sF�6���t�l���׎ͧz�cq�VL������wN����g5�&8J��M0�/��A{�	Th���
r$Џ����hl�Z*%����cJ�w!K��D�ǚ��_ѐ���}.�e#HEs��Z�'��oy,}:�}�:M��q�p�QY����u7.M�^��S�o �>2����
�u���&�a��֓�5n��/���X�~�7�ZJ�Bc���Tp�f�x�Krn��0�g��������mm�vH���UmG�
N��ڑ�dd��j����rN�+(�u�](�͑����ϞU��tM�J�
~�(�(xa���Ӧ�P�O��7+�2�������1mW��s��X�kJ�9�,ljG��ᡒ1��3�$4Ma\�w��ړ̽
B�ra��Q�n3�I�vˢp�s�ѸI�c`�c��M���q=��0$��Ոh����]�O���w;@��9�Bp��녑�E\��xq�O[O�Ҧ�\���C�X�+ݳCGĹ��ϕ7k�1*V̾尶�+���_��I�OhтT	��	�KU�gk�dg��x陈Jo
Ő��T�g�9]>�HN��8�Ҽ^�\�a�!wo�������� ��Ә�m��5Z#���z-v�I��U�����]�|���\�Gu$��G�!/����*�8�p��/fh?CS+�ٜ��[�4B���4� ���/��F�D$Tإ��d��A�z������G�ڱ�-� �5s[���7!G�$��}`�+�*!���Z^iz�nY��hy	1���\s�2	H8+�84�}^IB���8>�oxd*-�p��������5j&�v��!�ne��+�M�2NCѪ�=��2oF/����c��Dj�ȥ
wY%��S�SC�3y벗���E�)o7y��S�_$�| �µ�x޹8�<YFv�6f��4�%��D�����J嶶����Z�&#2P���`�=O����/�ǳ�Ƅ"=:t��`x�`�`���;�|c/��Au},�f����}Y\�&��^Z^�t�p�K/J�̒��������:�����l��+U~�
<e3���+������̈́�r�xM"��V���"^B��c=�l:5cd�@"�~a���
ٳj�"��[_���Jdڞq�����6%*}��ӳ�P����+�ٝg�k:�FmRv�[�Xl
��	�<�J��L���u}d�[@O���2��(3����K:q�.�&6F�~���7��>,�b���E�?�C��t�*�	�.�:*�,g�Qk�l63{�c����f�����(qZ��.$�Tt����}� 1�ި�����6X� ��l!#Ú}��)���"!}��F�B�j*� �F��F���4�W�دN+�$����lب�JK1rz�i{�p!�y_tI+�-���m~n�I�\zM�G�o�ok�1O���e2c~
��(���k�>��}@k��&���f��j��_�1`�T���Ru�F�Q2ٿ+��/��^k��eY}f'ǳ��Ď��i�ʕ��Ѿ��>��a�L&U�tJ���b�d��lf#aq���.��XjDr���סK���b:hbm�T��$��h�(b�1�� Y�����^�PO�&=d�6�Jy_J��+��C0�I*����QQjy��Vi����e�L쾬�x�ѧѠ���z]A&��=N=�q-_M�����b�����Tٶ	fǔ�,}���nFW�}��1~����L�V%4V��lǅ���W.~E���P�U��u��!�4:�D�@��e�M��vD��*K��p�م�<������^:L9��˿��_�3�p���d��97G~�E!Sܣ���xı���~MU�#Ӄqp�&I&u��45i妟w�-�TBήv�� ���=�oG�a ˋ�һ$�{���`�K�w<|���bʆ.�()rs�V��p,�k�se�� ��8P9~!?&t� ��<c_ʶI#������z$�SG������0oX��K	�v7���D}�Lhp�Hq��ʚ�����D�vބ�:,�J����2����^���ƭ=��cʚ�����9<i��i�!��~�M>L�����Ws?N,Z1����]4E��&�En�~�LmE��.O_R�щ՘����k"���A�
���1d���VeO��ÅW�#�D�l��D���O%�>�,p�Ob�aP�RLsx��s��+m{�}�}��L?��_i��C�K()��jM�_����޷-l!�0n?juE|>�cO0�$z�q�Ec����<W\τ����E�ʄa���x���z|���(Uݦ�C�O����8�E�����Js��NN�vڷ>�d�<����v˫)�u1X���|��t��f;eo�G�~�>�e�x�
Ȥs�B