-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fxgL/hOEFhOMhfWiYeUgKYXHtyPKAzinK+VbiZuucx6l/TFvlTjw6/k0cPlSjqaJg98zWt8ZFNzO
AHW+XA04UsC+HaDJ/PAHxiPKEtN9+TTwtuMxvcvZZqboIA85sjY6GVNWZbP7w5INVZBDMQiXOWUZ
v6d10NIS7b5ZcKTniI31TsmTSqnwnmCcmzsZyYf/rdq+J8cYuwQNdX15TxGEVSQ/5zzt+aD/gP9D
tMQiqfScwXJ/0YUWwICVW0hgneB58njod9T2rifirR2znXAcTcNxYUiXMfldAUue7UG5PUupc7M9
FqEJCC0lxBFnqesGwizTSYNVaoHpSEMJZpQrUg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
7SVfStuLvZly79TeG4rGVwcO/oyGmVgE8VYV4EvkY8PpTkF4EcYZrgzUd0FjrdvFvZEGeGjJ4v9n
xW2qcPxhR4IvKFhxQRCROEe+tKWgXrw01ntrYbZ/oP0upZed64sfVJ4DMOM8LcnT8uORF/sjwfk9
oHPR/3AJAZXjJufLhRLfEt0Q0MV0Ez1iiUDJpLNqQdQCM8M7RFKOYrzCK0tSFpGxBaaL/02eldi4
3tXpW1LYGf3v71qRufrcvyEJnArSAG6/6aFjiPIeRyuRCadIXqY1pmf9I0pOWjKaqrc3jSd0ktqp
FGF2BS9HFVmi6ULMYxPXP8G1ssB6CCGkkdn7762xtt3fHcnZw3sKTMf8d6/8nTRsKcIwPgMaPDIf
bewOX5of9WllXe5RUxzvQ/YIRcbYRtsNQA4in5uOTmtLEkeXDj4VsSan0nS2tcSeJaeEV6x3bZy5
Vk1VEx/Y73KOKpvoELvsL72RnMYu9Ls08ivPJm3ZY9H51HCXp0twXxwO1uB3wYPlgYHVzZ1bbAQG
6qvnLRpiWxLMfKa2S6eyFSHenagnwLsDWTXkPOpLzJyW+sUGnwOdN5+MAIpd2vSDHpIvixFYs9dP
e8G48cIzK9g6l2eZNA9lRx/XvTIPKTZLRc3Q5tkG79Ee3X9ZtaHjf4HpVsppai3pyt9TWhLhmgLR
V/6PbOBBHPBy7DBwV5XOMxTHU7bXKnole2xvGpbH04IeIDnJ5uqLtDgWHQe8m1yECUWwMc3IzHLu
sHoSdBIvGkldSnvnoaPNK3ca2gF4mMfdoY2AH21O42kbNRjJxSjvExcOxjWrxDhUsVwc49J9ETqW
MmI7CNieKHbaF2vb2PjmXopkw6cdywLmmT9HBQjVkJUd/gBRk93iNhQc5hI94tabbEsTaJNOGSYi
5FsLtB5eHjb3AwHk2qvnXA6MCKAKqBjtq5kvuhI2JvqcfHul8SlRt8OcWrO/AvyGeFN3R3NvEgDA
cmuXyhAVttd2sySSXYxrIKSz7lLHw8lXgSFMBZVoUbGp5rAMU6rykNAJf7cUXlE9ZyQwOF6CxlZY
56b8tbbe6jfidjJZF50Y53BPva8DpS0Xieuxj1eYY2WdXYTOAxAcyYald1sbjDWTt9KN42OJRalt
1D/0VnXyazT602bJCGZTZvbONh6g+fv0Pv/0612bh3IfrsFdoppsc0ifT/umUq9f862sQHYls+PR
xDnAXpA4d8qdFSWE2BvIcktwgEQecYjQfUGdLDZMFnGjaADjzJZkR5wbn/0XKPj51Dv+rSGkja4c
DB4Uiopnu9h0/OD0o99UP+7FeewIGz5TDHrlOWTZ91i6fK3Q8rNzIPuLVdgVna3bCCpazuvQM9qX
YKehfLLgE7jFn5O3Fxd6KdfWSQTuZN8HHeFrdbynkmwedhP/aY+HV8nJDreI5ASJLm7f3w6uYHIB
+iLCvrmj7Uo1UdhIpwJX25Nr/I7bLhMFVuLO83DYTS87WzNWOYlU93GnQweQ8RhmNmmlnBFXAt49
HYIJiC2RjUR/ysqAtwemTbdQg/hh/hPWuNdkCa58smOAtoeHxzOsyE8U422AR+bFA5I0/8x9UzPv
at0KZ2M7Rl+Gpyrw/ljEsysyeQLgaLiB6FQaH6F2WyhA6iQ6bvDhCobokHUBen0YtVBotJcX3JJK
rw+DtAnGhrTJMyq3+Lxa+e4DbWnUdDXejv23kxaN8kn46KyOtJyrMPJL3gv1wwOhHjNj/1QekKww
9r+tQ3870h3SgJmuy3iHdaovg5mqNd+V6iv2mBTHHgnz2V+0kX2W+yFCQUlGENvjGMm1uIDz5VIv
VQp4zOafcWfj3UoO1ryRZLt50rLXFusGJH+zTn+sT72AK3xdDQwc/YlEbdKGI4WFDKmZUqAeiFbi
mPnXsp3FvtnDEeXnCl/jgQY9vqAz0cVjfXQkpqL6jCARIWrLOZ/Pn8y15oUkD3kCsP31VDzVv//z
FzbasvvIPA8D1/1b9c0xOfJazpgtcwUzD24te8db5yMcrWZfJF81umgIa+ly5OtdBMdeZxWLr+G2
zuxMfEVtBKfI3JgcWbIrI53j3VKPCGBvFLCfBtH7baqnKeCLG0SDriBdC5vU9NkmjVstUWJR/PdH
X5C5EQFXgOjWxjoCS6rZ+wpWCY5bN4LZOWIhNSonBkX/QJ6zKCkZ7mQR4bJFfz5iy6oj2fcKxafR
IcMjjPoqpbpjSNqBzKdvzTdfu8DfVJ92uRu24v48X2h/p3j/BZhFH72NPT3+VPSkPvbiPWYjBtqw
pZfeM+YnwsoeSXX9eZE1j3kycQDSb9mbKPUeqMkV1pv2Q5fFtLesfh7C9vffikssU3LzkCp6nTcJ
cZFlGkDqzHuvZFsLqjUXJSGXqZMxrpdh+iKQYwzY5k/SAikyWjWOqe2qK4cFlBxXP8b0X31ZUAPP
z5I+S7qtmtcL8j2Ll6GfCujjFBvxPFca5PpeR2KlTfGMjrJKMVwD/qkSUw3myPzeuMEgQjTdfuZP
VZzSbYMYZSFWsD0LdSqemcw7r5rvgi6Y9tA0mB1lzNMq7Fi5+tJPwOyDN4pJDR0oCdn5lCGG3aQU
jX2hElC+m5kFFVI0Nu+ftYSHMtaEkgklT+EDb5RRR+ZRTmIlhBnIPdOBnS8KMbfcejYujVKlFTi3
govmljSceQvLY1Jl0IXVff6awcv2/+zZwvGol9ofW1Ij9Q855Cuu/Yl1NivyttQuuMgqKHdrXOuq
bU2+mVYp7GeeimY31O4UO3TI+qJZaCbr46+SzzLsYoHFiIiZbuV3BHKVpVsaFW1m/ZGvMpfYzDBl
gtzAzE7u+WyV6nhFxB8+bUMVa7QkptKVAgGNDlQ8NVtOiCV1IWx4U6w8irp+WL6j+UAsQlLHSsaG
mY49GbeY1ePcBzhBazCocnPG8SO7KVEHbSnNehRGYiM2wDisejqXScrTDlE+goBoBq1RGtSPRPXT
kVk2shwVi0C4EX3NakahCzWfmKtTRbZddWFTuM5BWG6xOJimO8MQbBp5jekLCMPotv7Gjt55VsZK
bOjDR3tSqF3al4yWZBMNxc1b/up7+CgciEHpcjMOYpoCPXbs7jwbe5pSmIyAfa8RO9iMfFPpXVFZ
FPMJ0Hpu0s9wJ6rlh2wwgBOHKmPy2YDLA/3LSAvpqxNs2VVTuiTZBWjqf/UwLY3dtOHYkqZ5TvZ9
wih4a9TTifRITXTudahjZw1dyC9BBdFLGdKnHCkhpPIlRvSVb5Uw4+Y2qKiL4W7RjEM1NwpAc4Un
qksTeMHSqUJMm/bEDfZos4aCVBph0Bsltd1s6hOhSE7WiLXKdI7zT43ru44670pOXNsCLKHq1I0M
DLKd72W+ZqIRaYt6XoiBdNJS/V6drwMEUTW4FLPqdTU8S3ZQOnBRpUZ+rklSr7A/tsQ2JrSlJxLa
qc8Oa3EVKfLYkUzJnJteHL+tOyHxMWe7OuyJ2uFC1vsGAyEQ6SA6d1PPkWr/Q67dONVxywjA9EO5
z1q/adm+xkFoKj/5WAVDzv85Jwc2ZbC35FIdysyX9LW2WtxYiARWI55b2tHMhzGgJZVHmen58zH8
8JaunSbiUDg1ojiVe2Mpvtdghfg0W5gZunpv0/NBpftwSjWh2zoEoThWXDCIKkIeRfJiN8gnuV+K
Kq/S9rx29p9J/Dff/h3CymmR9GngDd2JtlK4gppVwN0gcfeaQ1Z7H99TDN///h+ghyX0imxvd0vG
lfctnaPIF+8CwFhKm72b3PwPVThQQpngM0rpRG3s7vGQpYtTkMjOwk8IsxDU3eyxIV4hBHsGKa6Z
JWqDLJggMes+1C6BQdwEaKewsRB/VQvDjWxr/LJStubfBYdzSI0kXrKznbjCLGQOs221OTGJJfZB
yLnyQFwCDX1zca1emWDa1VBwgw9RJoCHpIRKT6U1wxUYcI5QwDlCGdcvIR2q0etlkZvLGGUzvOGI
ZEWLZHUJ/ufISVc10q3R4czEgN0MJDACDUPYRt/2gHoA+1sgcZKSxdwej8QmiyId5ClwZwiGkAU0
gSss3oNiI9QIpyvX0NuN0qB3wSH8DDI3Wcs5tM1YAZujzVS18pQ0MgVLINkvK864ZkRLffhGuFZa
xHl2UrmmP3ctM7P9Jq5o+q464osQQywQneiamIBGj2HHuhoya5pBJvVLNBg+DFeCYLL1U0Hw9xeo
2LwKs8Xt0Z2R4lMQQY+jK0R6pLQ+FNGUMqwEOINokKhVNPLs4T5atm7fXa2dwEf/UzQnob2GswXl
kdNf8oxgDNLU2s97yNb4gFm9TNr+UtPqKHJPzYMDW49Fz/in8Q33OjpGCKo8OyPWz40NFNG0aKfd
6Ynd2siKKwcl3RKX/+Sb4rgnmrwLLfQeGs/DpmvGl8ed99SsfoX7gGau6xFDKkFAqR55RnkRx3Uf
kCLvJFpuuoWu8RmB0Tg88urZtQRhbi05tfcD0EZ9OPoDUTLIOTBmQ7WpxNEYtrcCV9b+f9Q7xSMk
u2EJj8NuhYdTx8yAx6sUxugMblSSV3Ft7VK19zEkbCs2PONUm6qbas46fsM8B4frN1p5xzj3t6Rw
ghhBgNCbU6HR19oHNmErOf7utZmEbobk3VDqrZg9by3QI1OyMZqIwQHEsYPPrdLnKqMBm+8reWqe
SphEfAx0wHgLry/8vUKCchxg+9tt/0iI9ikU4ezwbpBigzlUp3BZ1pQJtjAdY3lxcdzJ7gc2HeVh
fZ49cum5lSjMuKYK0J0TY9c2xU0Gq9bxeIpzsiAlq9m2cMl9SvKNBcg/EfZtcqDLzIawKjEsn6+i
Uub7VF54YkKQxFQ84Rp+nkBQ+VL85v2jNYXu0aQNmo/TdrrKFcaG1Zu2qpq9Dwlc+AhtDoQQFO3u
d5M3dnxvW8YWbuMpMushBQa4iKOd7PQvTrezUJQKWaOdfnPlvBcrc91BEajdxH0YrRZRe5N/nuAb
kXrk0SsbT91+YOW2SsRM1DFOdXmMDcCsDEShdhWzoQ8cvD/RWLMn8KTryj/76Aa/6mi8Ww3pCRo5
trRuOLiCTFiK0NThRs4L4s2XKOkIyVIDohOD5ojCore6PFSPdZOWHhJDhF5BSwgbcVlL59tHBTnl
wKLOc3SbFKunBK0ylKu/Xj4i4ITz1wx+dJ4j07rwCQqiUcXEvtCkW3shbJhVdmdJHj8uHOCbDQDC
yHLk/ExII6YYJ6sTVbAArevI/g1h9dc4CjEXI/Yev4PM2uMwh9HRN4ukwuuuhT2/SifkP9JUvAlx
UejTc3B2JjB8QIBRM4K5qcKguJaVB/ed+8Gyaq60yKkEZRmjHARn6FxbRxNJgsBNeWpADZOJo9Xj
0YyiVijBUfbe9qCvWAcvzGwFZk4uNVvQlBdI2saC+73uHSy7aKbR633odra2c0mJlf5/zL5xya7L
zLB/1IKiFy9H6wM7Jwi4PVrZguj5s94gNr88alIxW4muufg/kqbQWAKTNdUZt+VizkKTggGkewz1
QO/iiVHsbP2j4RYf1kQybYuaSMI4ZbBvBbNRtuNvn+8XJHpkqjJ8WgXLaIfkSZ9Fa9iJLcOsUqeX
t/M7Vk7sV0u6InL9dU5GW/1mX1YuGz3jIP6JQv4GHvyCA4uTnKLb5E0Tn3AoVBfcT3lZLYfJNPAL
MJfe6D1I1eHx9LyQCLAq4iYxOwtoAEjuBLiUvWw/Whvidq9ExQm20hjFGwKFCz1RWkbZF8Aj0CCO
cJA64XU7oA/OLoyxEyl3mbyD+KoFxy1/jVlfF5+v5DbsxKDJ9nlWfDle43QJbBwJHqy292Oe/6/a
kWD3CX2sRLhzq8brdIL40kHe6K8dzpLJgBlWh6eYz7o+HMvC1AQV5aO1XPwYrLRl6vb/mPkGdaKy
U/jZMBDn87GZtA3Nb1AHtn0sIjE32ajHpF/CFzW2wSes4FfyOzQBfi5ZF7ZPVMBBYXkNrbkP0EB+
Brvb/JeSXgb4lG8GkBE5eMMPf/wXu8TwMzKJqzYfS7q4fHYS+yRSWMyiS8rDvrLPVjY9JPuRjE6v
MQ0V6vnK8uDicEJePlSjjUXtbqWZu1BjdSyluhsX0wbXkZ6sYfTA2Z0bIsU4oC5WODoQSROxbZ0x
oPhWbK9w/JABIvTzpFEY3ibvzAfoFRUG6rKP9BjxfeoMXUayDiEeHCbovjR3aU8gvgOGPV5hcH+/
05wNy30lLFhp/qtkoldvGq4TE4HqxZAWKeyYqKDI5mb6D4fdUWQfJgpYitGLhUhqLPNqWY/ZYMnc
J+SKxoOxXxewv5G252HXhELiIaQQifpS4P8tflM68lXDBOEOGjU6G9utzt9DKwr4eNgzBh4kFEp0
Shb9M1KAlb+D0YjiFQ92s49N0hiehRZLeik6TwVIReVR5BgnkLlahQ8Ex425sg+ZFOZ8fhH0GTYP
SieIGCZ2QYBTbTYlLuYMzAmAbEkcgRCvBRsupINwqlNXwIqkVgcdz3TGnW0zasMUQJV9F8maDhYM
+OVblGbliNnACv78Vv7O3fr0SdbyxbWcaTG9q21pb0Bh4EtrTb+aGJniv8uK5oSz4Hjpkk/W9tfW
q5jR7d3VchEBMThYY3kkSJAxc3nNX8KP1VCOG3F9dLIAA2eB6Es4mC0uFXe7ER7GH4AeM+5A0fp9
nW2KOqyf3X7P/v4uZtzUrXs4UUuqVm7vXEKeOV7w9jh3zzT90KKIxUqEiESi27Nr3SQkgroizK2l
Gh1pxfZlIrwdwO63pUje5IyyYNGialzYq8LFVfiBkOv8BNQVsxG6AOR7wGV92JCgccTC1MTAvpxp
+/6a6IDnqA24q7L66IVcQzk8rs9ZLeqfJ5RREV/9kgilG0r/EtU8gxZfflfOD6O3pTTBNxXk3gos
/jtiGnsaDHewaVDnp3iW/LR2pVuQcs862F2lpy+XOtmJY6AMTfCZn/NkImxnsy2d7cblhsLad9OX
/0gG1SakqpEH0rAdlgZ4tFPHpzz7f2y5oHAi3uQsCPv0aKqn7ZmwjZrwU7PRRZQw3QP8VAnDCdoB
YWms+5KwbxuIEoW81SrAYmz9SM6NualKTJD+1y9EmCHdLcN4OMzK5uIGetj5Rec+4SsO2WewGMH4
jGxklJZfizNh+6QWqOwYvkDyxcCvxJ8z6Q2BIVZeGXE0yPl3eCBWnivKiSgd+bg5YfLN8L7HZEsU
kuLylkwYlaqrut/0+gMaCYW37kc+3FZ7gIVvztVAuJJQZxKTpYmA2qB4rs9PChRn9AeDycxKnsnE
3ztWWI8g5dGehQAoMBcPd1UkzNjkxe9q5TlT5PolcvfKsKXddiKfSY54lROWuDTzsn/XEOrqTMel
hJwoqj5k/f8MQthYS1u5CDwmNS/j9VnMFOXeUMGlx4fTnC/c1a4j5g2d7/rYBVWXPkXjin4bURxm
xeWlJDq3e7vUX0E47DOmzEZ2Utp0vEYX/mGHSl4Sdo1KD9AESJoO2iImTzfFkCs4XtcHZHzXDFMY
RmRha1phXERQwF3d35caun8S94WwDegjhmU3yTh0pKZDlWfMvE9KrOKhvwmZzs0nWIx7CCqpyPSf
C8bcRgdSEohkuvN2xqovaOk329ej8LlILSV4qTqideqYt4ncGQk0TDtkap1H0JqKMP3V7oWpqswE
CHdDXdy95/nJKXh8yQjqEDzm2+6zkqkCKf9Nase491aa/72l5xARZNrFIK6nhu9OEwu274IFMokF
II8vGKiuR44WUsiyilXMk+OVPrNg+cXa7Q4vCzzy/NZ55F0qHSrD85FVZNfhW5VZpGxtJ9wjM+Gj
vSrhg4Sbbz12YQH32qtDRaprLeDAqt9Pd1qu8aKbbq8xXLGLlibvudj+SGjV87pWrCTCF0oM4hMk
DLi7vYB40p6OCDMdlOSlTL2G3YKVP6yZgturf6pCc31hBqWBivEwz/47MjDiTsfDGGUK1wH9FoN2
D1QEJePnub6zPp9Jfxr0PNOQOLTX6nLzRplaCDAMf2DfiRsrHGjGk/ULjMJKWMcxooHVGCYBPsnR
3iOvf64lGTk/nYWxupcMOrtFJ3EV83GdBPiZHtLYPz6UjXegl2pgsHRBu3Zfzt404gAN5U5VrKhM
59E0TcM21fpuN0GCRLTf/57cA5nQMoYPVmT6/L4u540SFRMvYyR8ZX/V+d6H7JPp7LpNpGGKwMLW
POIr+u97CKKVcbMDvbvRUIN5u91TJOIVQuzC15QVFHdqq/5neWwulwpR5NFOiGvXbUhnejYilfDR
p9gYoOc2XnE4WVkR/rnLYi0lYh4+O8Zg2Gwp+dxqkMR12Y2Q3r+IFwuYWwgA1EWjs76dmO99yaKs
d41aTSXJa75HjJbrQO6u+20SeihCD+Cm54ukXjR7uOpBniSZ9EAeCWUBYhOS9xdJoMgzYKmUQl9X
IAozj5/sPZy0SFDDyRhjwstcxBmOwLDfXHZrAyo+GIs2tIRSIKOgIhzrvOTV3wQr0qmpcevD2csW
qkqosEMeLHvl8Y+ToFDdohS9v8EPp6Vp8O3NW7l0JwXfjzRy60A++g17Yedld+OPd+H7cg/VujqJ
jN0QyIpL2JMhbCIpr6Fc23gNIluNbUZN2d/TNtIZevX0Ro/lgP4yYCMkYF73F6CpX35zJGkqBiZc
esiISC+b9d7KjJ1mW7Qv14ZRAgzqyu6BCV/qWWj6ra67WBVI5iNFMN0ap1LKfQOgl4Ajg/WfXHl6
VJgR35q7krtcrjM98WLN5X+cdzI9juw8bAJ1XmBDFxFfOeeJS+IfuKkNiiT2HqAxBxPjvysMzAiC
P8vkNh1fz2/gDnn63+6wnkIBJb2h3KVLxcCB6KoSoqDZgUk0sXPLtYqe2gPr89CF8B3cQOxVsIAh
+1mpH3l5gX2VN6TlQYVYaYes/1jY8G3k/3mYyzLOZXbqABfFMsAWbhRQ1VJpwl0k6w+tqoAvGNw3
YqsgcORBgyxAkNdPFif+NkXSh4PJZfTk0BY9cMeShDTG+hHBHzbyGPE3iwmey9dGKaPBbwCvxaP5
2Ddgq8z3jSTJUG3WMIbXS1nUO+4Xkck86+7mq19cGMCSkQqJ7bAk3FgIxBDifV5LLCJ9nbj6oPlI
xe9RMe63l45XZ5ycj8YwKkiKsPRgSa2xneNx4QBrh+bx4OWn1T8lVLdn7OwexTb0640/eNK8SJJX
K6+XOhvoc66wvCrNpBB1a57utqfed9alxvQgnDwOGxTNhNlmV/P5G/OFJuuTlfgHFnBV0HMt+znE
gQ9XDavKJ52goKpf3xP6vxZrijM9BRZI16Kh+cZC4k+p+yNRhGLqjuTk44rk9iHB1gmUQq+nzeyz
ig1WqkbucFSmewBLRIxV9V/iQd/tiVNvQrRFnGktam5bm6Fc3SMSvRZUgldpSuEZRzx68Ecs/7SC
BPWSimjxShaxBN3BWbinwJ1peeToJA+lPC/KSmD7SIGbhwA+6B3ZYFkFIw7tiDivkcuSzkmtpLaW
U0GzqFfeGgWmEIyi0/eqn4S+fDhW97x7qwhCHgxZf1s4g21x7m3mYi5cKoa4Bn6DOgaXxa8sGwa1
EycpY7ksOLWNcOC6kvLdhRgQLtCprgFmin/O5dnRTv1gFTHGfLCjlM5GJ3+Ll6RO2bfc/15MuQpV
DkJdCw2+bbfG7PG0EE3KKegirrF9IIPKaykcHUAKQWtmw/mrS4AeSd9LDM+0NvUxLIfsxx4QU6Cm
PTY93ZrjnNhNGpO/iIAIJ7t5TGZuzcnd3cs+FXPxarnxtwCzNBx7TthvqwdNUepG4VGGTSvF+ZXO
fxjuMNULPERojee0z5Hr7mem7kLqcL3u7XJrf258uGOwVlsy0Yh4Q/2FLlC0r9Tw63/NTat4hGHF
rlF3irpU6c2OHEo9dM73rFsgdSk2rGB3JzEER87rhnFQmgGbW+gPwMMrGrNwjtYE4NW0R8dWFcfC
MCzJDzSy3N19uAbrPvxhpuF+h/q5NPFIAd6n3TxJ+D4Ke3KvujNErhv4R9JSwpaX+lLhKAEL++Ki
Lch6cYWmN7zgOseqBMwTTL2DsOIzzXJhXpLrDqPApLtINJG2PBKemRVa11zAfmCjsfUlpMI=
`protect end_protected
