��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}��,d�)q�n'a�s�0~��N��C{�OƪR�)��K����Ņ������6+��˗5���#
��	�Wl�x��LZ���=K�r�bH�����[r�u���b������9׋8� �$&W�JU�+~ T�~���M6(���W*��FC�:�6Ɇ��]\7����,x�&w�gx�}�&��&֎Ղ�6���L��t�pA�4z؇�}��T�ny����M���;��$�ͤ���Z03T@��@n�=a�C��B<"����-S�uI&�>�z� \��T�'�xO��?+R���i��n�T��� �xLV���f'�&��h?� �8sഽZ17�i�����	��8��)K���B�w��Z�#V���z�Mt���<���^,Wś���ϴLJ�)��e����((���L46�N~��h�g���F�x��"%_:A(�vHR�r�q?�IX��SsM�D�իHcL.}�Q�%obOF %G�X#y��]h_.��@Ųp���a�Jo��qC�-c:���AJǐ��#��ǩ��w��6��;�B�g$z40Δ&����"�o�,�t��D���<��4%
�Y����H0V1k<���R��q< �S� �+�+T�s�i����/������務� ����� �NA���I9l����52u�5S�>U	i�K-���F59\>�����H�%��#d�i��*�2L�t�FStH�D�w�x��M�����-�
2�t&��@.˕��D�z1M ��U��V���KVR��ٖy(��9A#��E
���4��<:���11,2��&X�ǅ?�SuV�]HԵ~�D��K �F����*�]��(�lbO:�ܾb��
O�7z�P�b��p/���i��� U>�="�LB~c�86���.�GT�Y��K����]��?�W<\[�:��9����'��&�Bi*O�����v]/r]l�V�G���s=��r���Ư��ڝ\�4t�x"�T#7��7�/����vL7�p�%�&��NE�4șډ�*S� Ǜ�o xfP����q��c_9�A�H{�]�C�Ek��yW5�V���Ԫ~�>:�œh�n��V��*��N���U�Zߜwzl�#����/O:0��g_����W}�H��J'9�n���<G�%�ܞ�sL!?�鮒 �=|��b���aeiyb�/{<��a��Y�[r��2�e�צ�Ơ���Pd��c���-dN5i?Lq�HmZu-�L5�o�k"�$����׾���4��I���N���9I�ɽY'TF����D;�98a4Z�)t(=�e�/h��wQ�v��8Z$�>Ȇm �*[�a�� ��-z�0��@�Ɓ�Y����GB�1��jt��,(-J�Tѥ9ƀ�wA�m��BI�S]n��a���(OE�Q��|gdz �?c��T4�_���{��F	�A�vѰ���%��{I��.mK���;2�s���5C�%D����\Ą����Ւ�K��\��t�aSl�B��R�wDa���E�c���1��I#�(�%��V�b9�]n���cR[�9㇆�B�6Uk���ݍ������H��V$��a�����t8:���w`�nl�s�|'���5���iDf�.���o�Hv�&�Kk"�'����VA�����7��q�-���Z�@�f�k�`G�QG�*�N"���3"l4�3�{�[_�ƌ��Z��$&��_2pn��F�����2��΍������>p=Ա��%:]Dh,��'���c���v�`� ���c���V���&�c J1��F�u��K(b����7��7��z�;�K��F�	&4|˚T��t�3k���e�a�%�р�_��O�2��NY\^ܵ5l3!=���!�o 3#�X�/Ta1�Ă�{�#9�s'(Y�v9Xn�������T
�M+��¯�z�%���r�W3��{��Y#6�"�s�,m�1/R|LAX�O�Z�P����`C�P��������?�j ����]t����%q���0�'v�Ln��c3"�V��/�����۳�UX��nu�,�2�a�h������������\��[��RW��<��HY3s}ԑL�A�!�^�wԞ�vԯӧ�R�U��/���-�i��H����S&�����W���	*>�fZMdBhҨv�FtJ�8��!Hjk�N���'�mڡT
� A��������oz�wb婂�P��j%���S�_0օ.e^��T�sT'$��ֱ)�`T�E�!I��uU~�2���[%����.�k��s�ؚuR�k��|�q���G�����!�4�����	�*!Qm�$k|�V�M��
�X���!k��iT�KW*g��p�w���TO�"��r^h�P����*��S�>N�vc���դ��m"�)���=o�2���j,�|"UH�x�5nFj!�ȡ��V"p��Dk5����8�t�7����] t+F����~	�	�ݖ텘l;0�Y^"��
~��s���..��`���iͥ'EZ. йӳ��W�)�y�b'��ٸ�WhJe`�-���L�I�ku�ͻ��yCao�ȅ[��'�	B0��Y�Q�\�zB��.F�n`�ZfNŧ��3��$F�/�>�>��CF5�<QȔB5;�vf�t�����x�+M�(��o/%3j �7����Ea+�����%��Ƭ}ʸ(J߼6(��H�b�Ďr|/6���ˌ�d�%\��K��Ѡ���b�4)�����@YĩX���	��xc�=�a%:q�t��`��Q�T��R���}��L�F�2�z�C���:�ObG� �=��Sjw2�g�1Q^�5bj��R�B�Ñ/)G������\��/óa�5�����0a	|	>����Yp���Y�ɜɃ��u�����e&d�O�YZG��7�Za����Of�;1�T1nH��z���t��((�p�Y�1H�0����w��Y�#��أ���ڼۭf�݂(��+x{I��೩o�{_���H���P��f�i�,KGax�1�+�M���pϒ:��u�Am`+XF��H਄;��^a��R�5�m��gӜ%�U֨T�.�V���^�l�8zM��˞`]m�V��49��Pd�`m���0�)�F�(:X�*��^ ����Jb���PJ솀�5�.+88z'yG���j���1��eu�;��x���U@�J�;��Ѧ�g��b��Դ������k?#����tL[U�t��=B����s�(�:גQ���6H���3����VҞE�`���P�E��G�Y.!z��"$������4��:����b*{�����/�H-QO���� ����j����8�� ����Pm&K[�I�Ou�*���U)�3��gY{X��K�T�	�f3>�o*����)-�T���gӿ�d��q௑&�:�#Tn�S�����Ā��I~]cx�`%�����_���x�����l���w-�gMU&�N3?7��\T�����j&`��xwF�K7j��A�n�������\�9ƞ�3�o����c��?�zcܦ�7����/7��'���+�8u|���?+`XI۹6;��%��s��B:T�P7�i��094���WyGl?�"ə�#J��
Pm�n!k��x��t9��>ǟ�����Y�6&�C�g[)8�������-AK�~:
TBj�	vA�2F�'���'�/��!�����s%Wo�]_��\
��Y�4/�Ǭ4hb�m6����iX��BgRUx��mV���|���$ŎlXA��Iz�3h�4s����t��W�R����r�$�s=�,����X�i\�J��,�
��$*r m�u{"T�l�t�Ԣ��VTr�VW�e�F�K�gc��B\� O�����V�D��=�������ّ��g�\m �����Q�맠2�M����ؑY��x�?�� M=	^�������O"��FKنq��2l��u��4w�uz$	�6Z�1Բneh5�帢��ɦ2�ʽ=�J(>WM���pH?ZxW���_3�H�ٗ�I�F�MDˉ �l�;)'�$Ð���j�t�z}����<$Z�$ȉwC�	%��M9u�f����+��S�C����"+i9�I�2_%"�:�z�C�P���X<b��p�I-��VQ�Pչ ��Yw�''�1WGV��j|Pn/�`(��A2w�tM>䞛n��3��7���@��\���Iw�����W ���.��dg�����
K��JPj (w1 ���4%�5xĐB��6�*����C�`��h�P��iS�JlY5�huE���^f�;�Mh۴��R�dɶu�� �k��\�5D�Ր)F5Гa�.;�g���NN��N��-�U;�e���;�J;�3�W �=���?�u8���K�Vpr����qF��y^�������4V��-]cI��_IY��.�&�*&i3��ʭ��
���XhH�f��[j*���4`Dx�ǣ��,�7Q9Z�p4ɨ>o�J0쮃��dyjF�a�5�5��M��h���Qx�2�Uxϋ�;�La�rqie%q�|��)���7���2�*��>�B^Q�nz��߸M���ue[�/�tk��n�k�;�6�&l�n�`Z�Tx��T��-��勵)ta!��>����ó��JD~(te��$6�G���R�*,��&���䲁�N���Ks�Z�R���0}�A�H���v��6��}{���7
Ɂ�������>8��T�H�i-�!�	S2�>N���i%�1v���U["-����ȝ, �I�d���\\�G� X9�<�D]�W��;����$οL�P�,�K"�$>�K����.�̼�����G+~p�B޼7�J4I������HI���W�:0!˓��4f���_�d�%���`��a26J�̬{z��!J�ΰ����� ��p$�/3�c,<��}"�E�?O�ƞ4�V��C�qՍ���`PA���R�g�#Xւ��3�^s�?�h`}6:����d���|��Jר�$)���t�:���@�_n�Cɀ�O���R��Ӳ�a�7A� �
/�9ٖIlns�xJ'��'�~�Vt� ��o-�A�*���י��Yn��l�Ý�ǔ/U�Ί�~����P5��f�4�n�R�#�� u] ,PְbfY�,�PZ:���i���C�f<������:����Eu2�a0ID��I���ԙeT�v�^쯲)���RX
�S44wT��B]%p�!���`�Oԧ�O�?�H4�N���1X�����,m�f-����������	�fu�'���E����O��Ԛ��35G�}�܊�۪�=�uȨd��8h�s��]���v����0H��,�I�3�[,hF�do=|�_�[M�`A	R��
@�<-փ�[�p&�?`􇘁�p�\1����as����Y�cČ����u���dد��<��#?5μD,N�ȗ'I�"MY���"0*��=瞗 L2\
$ ϝ�^��5�r����qk�0����<��*b}�'�"#��"h[��U.�!i�rx)U��-D�|�E'Ý����\u�+�Y�{O��~�g�y�jM�bJ�]AhVbݼ<��ޱtg�H�p�r�>q�쫪��B�	
��<�$�C����>�#]�M_��c[�Ճ�B��3j��DVK�e]�~��/xp� ;�WD Vw�������Y�+ߊ��9U�w:&�ulO��]^�A��JhZJj>��1a���;�屲M�b�g�9֢�ЧMP��"�
D�1j�1ih��j�"�"& e�U�~Ӡ�yibفسm��?�����	�F `|����/gU��6\�rZB��q����� X�o%��ZRB�/�<�vE>+	Bi�J�sh��?�XX�hͮ�@��%@_�~��ܖ$Q+�ݲ��ܿ���n�~��r-���?��b�q꺼?gM��=S�>t���t����X�>q{��~�s����%���&⊓d����SУ�ڰՐH�Z�ZʩH���zEB�;Q��������O���'X�0	����{1��[�[��'w�1�"^"H\`쳏�z���ڥ�q\`Yl?�EvNb��Lp6�!2h=4�_��O�_�rTS:?�&�mv("��V�CT�%�o}"�7/����b�{?)���ɞņ0�s���k�`�,!�����y%��N��9��x�(w��u��'@�7cj�;7�6���PD�[�B=0�e��d9��3��",q��=�k��׆�ǫ�L/+����Vl�%wZp�� k��<����{_�VJ+���]4M2��h�N�N�#� #6��́�*'k0r4to� X '�g-�<OY��H�p�[p�ۧYO0s�����`=M��|.���N(@�6��o����y�g�;G�}��/��1K��qN�"�֦��͏�.	�{���L[��D5ֹ�:��3Uߎ�wߩ��H�8�5ȞFqsO�����/�"��8)c�>;��S-K�����ه���ܥn#�j�G���Q6�J��O<�x�$�a�*�-u���9�"a-�v7?��œafǸ�2&�� �%���mbH�����49ۏ�C�c"m���:�����7fp�I7��oLBn�_��5f�Z��k��~N!��j�*^�\r����]��������a�v�..f	��"}�2��}B���@�.jN8s!]�Ho��(�yPm�HZ��#�R�04"�u��5iޞ��#�O�t���F)�g��sV��S�4>M�bf��޾�q�& ��\�8�'6"�7�'���~��)�~j.��2)�!��K3�P{@K�S�<b��>KoU�Ulsy�� {�>P��v����ܛ���[-��� x������}o����!��؆�]$���"����.$�JG@7���V��$�y��o9�� ���g6p�!*"=y5ch�C)�;���@�l��g4/+M�"}���v��%,")���"b��������ۤ�ɗ�"��q���%����U߯g�]�.eF�/yA i�g�M>\������3W��;�k�����bx>�luP�qן�@���'��]�<�*�[R��Z	��v3��5@�E�m����D�2չ�ȹLU�u$�['���)���;� �^���/�No�|�5>&.WUO<�dE�8�3 ��'��%1۽^1N�u���Lu��Y�a1Q���T��N�ny���T�ft��J�q�C��_sLL��Y��aF f�l�>"��|�l%%�5��aKx!0QHhO�ibOt�V�g�Jf����Э������J��z�էq��EASY$�*�\�c3zMf�@F�$�C�fC{g��Eh]?��~Q
NF�Cv#0f���}�����kn��A\����|��~�<?�EH��P�xg�6C�Y띕	_�/-�F`��6����3����)�+����Z�H��6�"Ĭ��X�+W���Mp-�%�=�������1�CFƏ��W[U-�b��{u�G��deW�*P�%��J8,���9P_h�{_�}���I��3�*4�ȫ������xU_�Ak�� ;����,�;�^�Sk� �v�R�B���%$�ȣ�@B�O�񛖱��ԧj�9o'*q#�� ,wގC��o�a���C�L����_T��w��a����Vx�ܒX���bȔc5�{�6���	ǝ�e��j��o=J�:����)�T&h�j}p�X�z�-��eңy$`����'���n����g��os��Ũ��1%��)b�x����%��9�d�RF䊥��:���g���_uf�<-�9��\�B��?�e����,�=c��������,Ф'������i���BT�2#p��˾��5�^z#K���wS���/��s�6��7)4�e�c+5Dn�S�3W+K�J�Q�����H7���0�k������h�����x���,��FS,0��QŻ��"e��i!��F�\8��im���`r�H;b�MW��jG��n�21�/��B�y�*䓞	�j`/�Z�,~��:��X���˲���M�Ӄs���_��./9��f�r�mV2�jXDqƽ��ts�n�kBX���iX�9U��H. ?v��Z��ɗf)3⧅�V����q��WG�d"�ZD�4D��.���ܛ�x���<$+��1a�"oσ[Q[��uC�q�2=��.`��"��e���?��s���=����%�cg�QfB#1!�a~W�"�6�c�`k(S�v��	1�	0ueL[������3����F���Vō&�S�&Ia�^�7��0<�5Zi��v�H����fC��6__/J��K�'��9�e�A�*�#h7Hsa:��zI� ˈ����^pV��)^	��!Sn�~�?K@��ʯmē�=���mȢ�Xu��Ԑ2<�����<H�;/��^�����Y��D��O�%f��?�R��wo�Cd�SA����&ƀ�j�M�<;��k���w��X	P�	 �ݫ�������d���a#<�Ȇ�ک��a3�R�J[1�ύ�Δ��\��6��W��,��bXE8��|HN[@`�_i��n�`�.�-" �;������]o0oΖ/��K��I�A�Ie�Хa�h��|�#_�aG����@b���JBg�r�����W���+�\pW<�q,�7^��x��^�o�o-�7�D@N6���1�p�c7��qeY_S.c�::���"�O#���R�Æ�i���rM��9)���.59ni�%�oF��h\�b�O�'���$<>��dD��f�P�č��ă�)���n���Ah?>���v��o��D�&��G��_Nk���S0�ܢ�9h(��[5$hמ;�l s|R� ���	����~b��a����#+�d=�}p
�k����ߛ"��31@��i;�x[J���Qʆsi�����h8�i8�o"��P� u�3��UWFھ�8�B�d�!�@��&�ٱr�BN�nM��1�����)�*���{0�X8~�-5���7�9��Kǘ뮋c���b�#�Lf� �6�+_�!�/_���r�z�^'cF��"�>��u�F���ӝ�UM~A!��S�%���8�����}�Q�pթ��BN��d+�Tn�2:�J��_pN�n��4@lQ9P,$�\�6K!�&M/���=A+w�p�:xd]7w��p�I�����6�􋖭P�����D2�KΖ@<�~�7)}��#��i�/0[&��(s1�-�*���1wF�]+�T��i��~��\v�4eKߨN8�J��aq�]B��|���`�k��izx��a�n:��߼D�kj+q��9�_��i��I:x�E��C����qz)7]9~�a��uE
�1
"]7H�=	+�.��.t�ϔ�ٚ17�<Dɗ�)*#q��a�"���9k� XY�ڵ�e����A��Kq����tR��ɱ�A��17䵽|y��a�]�̷�k~|�`e��%�#�T�J��{Q���@ +N9��g.9�Œ��� {�?0_]V�:/5$	��Ŧsor�3������U��M���G~��ɧB�=��qdZ�hq�U�� ����Ő�{�TԼ�5ذ\ί�Q��
�<��UK�������{g�d���ވI��H�B�aO�2F�5,!.�: �<HGe��_�(qT��`��c$UT��OqQ�������Z�b?V��V�ߏi@�'>O�sm}�/�b,|�!?h1�m;��q������̐æ=TW�y����]K[ĥ]�p�����.ۮ�Lߺ}��y��p+Z���#�]��c�u���3a]���|P����f��Z��%0�vʡee�hl6��zmY쐿E �I����U�#)�55��yX^i8E��Ȩ)]���EAF�_�w�/k� �^�����1�~��������V��8$"�ӟV��VN(�1d��NgC�����}h2��1ƶsn0OOCÖG�*��*;��}���V��{�Z-�CL��H��ɿ��G�gxV|��ghYd�L�ո)`F.�q�G��V�"� �nǊ\�E�����G�~%����ar�O�ZU�#�F&[��O���f߭�'�?q�'��D#�A��	�b��]4E؟��:ӐXC-���r}�U�z(�Q�h_���
�ʌ]>yKӂ�ʿ]��jKM9�81C"�/j�D�-��N��YT�su�؝dL�(∻��jLj�9��XUh��lMX�!�_V�eM~����Q�R���Ő���l����(��&鿂%�}N��fC@V�|�*��'D�{��9�w������c�^�*.��17�a�,���7X���+��]�b˯�l����mzݰZ�e�^�TC��D|�#\<�R�"d�¸*
1�}^V���>����5��g\������1
��?���k���%�&N[�y �x�A�W'�[m��$�
Q+�z����͆-�f����v(\*^��O�=j�Ҷ:���{��V4Q�-G�#��ٻ�����܋��ၫ.�=�Z��G� d� ��ûJkO����K��Gx�'p]n�zt�m��'�o����|�k{�d�s�5tbE��Y�%�K9�J�`�21�[,�p��ɖ33��9��!Àa��,U"� _�(�F��q�)2oߺ$���)�R� (*�hʺͺ0��}�&����5���:[�(P�ft }���t��ʞ���q��l��8{k�ԫI��m[�c�l8���e��2^�����v�T��& e[\Π�iB��R96d<��#cmX�!�	��DՁ�����:��VS�z��id�.��ߏ<=��x�ĩ��5%��W�)0*Ğ�0,�������?��W��I��*�s3���0�����J���Ƹ��O:��	�u�Q��In����ǇP{	)8V/���,0z|T��qz���V��N;�L�s�?�P%_���6d��F�(�� ����/�ý1tWŖ<�]��E�3�lbM;�6�^�37���5���"fŜ3#5��HN�Z��w�'v���^{W|h(��*���R�͹�^4/�6�	K�|�4'�eɥ�:T�����o�:�sw���4�rK#�K���\�7��[�4�K�Zhz����6��]�䫜�I0����������)�jɻMˎ&���B̟���CQ���mY�������LA�Ф�J��x1t��n~��3ꖺ뷌�y.�+C�ѡ��v� ��.�1������#��b�j�=EͰ�b@��	MX��K��n��M���H!׺�h�3C�n}˽�Y�����d`d!�p���>�L
	�"9�BVF#@.�v��r�ҍ|�涒�E��GP1Mc���{&�$��$>9z�`�����OkZWY}D�R�ﭕ�S]y�c�y��O���<j�������Ë�|�W|�.�{���24�Z#y*�RmR����n�\r8��`嚼�y��C��p��P�u���L6���E�]�cm�Y4{s@�B�a�s*~Sax���<ۨ@���[kp)���kgxvVn&��CΘx��G���Q|�l{�7�@��]�E��˒��$1�D���z8�Œ���xrlN��n�ɵ�U>/����B�e�-�!��ڐ8S��0���X��@�f*Y���(�]}2�0+���I�G�.Qt080nQ��ރ+�����f�� �� ˤ��d�1�g��m3�*c9o
��p��B^����ds�q<���()�0"�Y��kT���U˨�B>Y���E�ȼ�6ݯ&��͖B����~p��)�(���lx���D]�+�����թ�l
ؚ�nZg�P���jƮ|��t�Y���k<*�F��4X�F��¯�;x���Ka,���J�B��������L�\����ư���������s`0|�H���C��S8�cs�O �M3�j$������@��!_�J;V�/_��Q�����}�*!����#�6���c&�b�M��vB�	���wL��v]�V��Ng����ͤ�P��N+����X[��'��5DO��]�"E.��I����,xOj�z	���a�h�uk$s3���j�q��Ȓ	.t�u��M�	
��a��-%,�qل��
y"��QbD*�4]�Fϓv)�>���9T��������/��'XH80��-�I�}7Ίt��)����p���\o�m�JI*�A��&kY ��N�咤�|D���)h)
�e8}�*=��X4ERh�Z0l�_5����X��Wr��.7o����=t��f�#��Mw:�6�1j\��Tn����>u�^l��
�ݫb�ppA�5V���[G��q�RY#����c���?)�q�aiV,�������"9��[ª��)�-��*pWK}�XHx��ǹ�J � �0������\[ ���s+"u���yh7f�.t��W���~G�@�8m�%PPg���xR�pz�5vh�\���۫���}>�?PgX.������������b횊k��A9bQ�CDz����e ��pY�ĥFk�1;m� u*=+x�#;��s^)q��DaZe藊�r�Љ|��.��j#Df���q:�
�q�x�ј��c^����T� Ař�%9�30Mb(����e�Vb��Z&o��W,2�}�D ���;��-�`26s����Z<8�ś)����(J�=�ѻiX���_ϕu�N�f�U��a����rp��!��LN6��O�5wedŴ�[bL�$��M�%��V�;��}��l\{�60��"a��/��&��<�8@Uy�����d�bW8�V��Ix�k ~~e3��4�9�L������i�Τ�ń��Ms-%6���BX�O˫����=rjk��.�b<�����S�P��L^�Y�Fq��ɳ�*g���\�3�̸M������ĸ]�F+G�h�H��t�)�m-�^/Ǜ@�ؒ@{���8Y8��1pG%��O29^�)�G"�A*s3�� 'y��1�n�,���Uͥm:nF�pωE_�������E�buu��_���y�Sy�W�g��$�F��9�;�^���N�S��$oW	"�w�gZ�����Ӂ伏7�t��Ġ�\�R�Ct����Fc� ��z����Im	)� ��zn�҄$Ԫ�~ۙ��c^�r�Aq�[��2MM�!OB�-g�������0�w_f��.u7նK3=l#�lH�	�@�! o�[;n�劔��wT��d$�'�����+^1lm�6<�)Y����p?O�g�]�I��L�u�4F�#�m�A�<���_���TqR���]d���CVѩeD4��Ul�<�W[�%w���0>�TcGy�<� �(5�X#�w�L��Ot�jCzK�f����ro<���3�&�M� c"�|i����[oZmY�}�0��8����C�+�� @��N�Li����fٰi#��_8g��)�R��
<��?�`,Y��g��Gs�����0�M�I���E�(�w�Oȶ����������,}���=�'X�t]�F�7��a/�#3>��%����7-T�w��`��Z�����mR<�j��������reK,u�M�G�V�~���]�9��zj� �B@ܭ���{Tޗ�`B�r�i��n�M����t�j<9k����ֵ����9�/)���$ܚ:].�3N��z�;�^�X�������O��[o�m<B4��c���1�����|"�뺉7�Q��@ּJ&�{�r��U�շ�f�?e�e�Mpx)Z)�=72���#n���i.�V�^i4D�;���l��٠�A:L����I4�v#���\k{h�y�y���}�T����	e���)O�����1�s<WM����T�)N�?ևƉ}�[����kT��%՗�aB1DIWPk�C!�0͟��ܗ{�Vq����4����2�G�ay��W��Z՟�$���4[H�=����P4�z��H;�0����V뷿.t��v��Ip6��V���򿎣A .0��=���]� K�F��pi��o"�*W�Yad�͖!�T�Qɾ��կB;G�k�S�c=KS���O=�cN/X���{���sE��#3�Kg�vĴW��N<=a���)j[��75ↄ,��/W7���M�;B3cXY�՜��W��#�2� -xXQ��D�������+���y4�����:��Y�/�s��q�0�Ń�[Lv�֕��i�M� ��$��D�=�n#I*<ML�M��w�\8���/_�ku�@5B��/heg rʃl���$(��$:�ذ�����^�F�\s�2�oq�j��兄�b���<ǇD\��t|u���zlHP�W��|`�i ΧX�m�rj��`��u\���N��+p:�uP��І�^�=����ec��k��\i�1� -����D�7���D��ek%��9�SV�J����iLX��q mR��
O�I��·s\�22@���J��;�p���k�Dr&
��)� ��sf/
&i��(��d#z$��-�6o}5�o`lc"����*O���+��:�Lu�'��d��t��pg#�"�-�b�^n* ��%@����H����6�cޫ6N/��Ѳ��\hj�Qg�Sb���t�*se�g孂����������k��H\���6�ۿ��p/-����y,/%}�%�L�G�����O���a���ػ�����tu�E�{��0:HT3W���[��{�C�RХ���F�z�e����BP��Ch�Pg�pu��;�	;,I�Q���P�+���sX;�yx���2��1vI1<�%{����fx����D���{T٧;K��t��a��.Ҭ0��Ɔ�8�������<Sm���N���)���W���;�+L"]M�Ơ$�ln"N��@�xE��mዧ����_�^^�.�e���EE���<��iT�9�g���FH�^��5��$C��z����ʴ���ē��+�6������-�4����)� �/쫎�,���)="n)��}�JdM@o���o1���Rq�Z��'Ş��ˉ���E�B
��Qn���Pd����*U����UI: u�
0W)>u8�����j��8)��� Rr�F����8$���I�~<�!�I�\��m��j�|��L�*�]���"�o��T�L>{��){)�;�BL� ���9I��"<�a�UH��w
�IX�ix�+7A���K4@D�_Ã~���0���*�x��R?C����O���%�9=�T�TӦ5˞��>��,rd�{g^�K��`�|�Ӣ�s-�r��P���$a��h�_y��m/�Vm>$�?�Ǻ�����|���1�S�S����F*�1��߬h���*\�B�j�P�B�I�EّoU�D��9����.֓�f���o��M���%�F����>L1N�\w�M|���yi�!��<�x-�G�Dr��|�O�}���G6w��,0���|_B�MQR
�c"�n�	.	c�اy̴�Ua�?�RՌe-�V��G��w9_X�fKV)viS������U��`@�6gc�]�i'I����^,��7���'S	�j�R�L�[ʡ�L�w��X�}`6r��� �yIP���k
��3�3q�d���
�""����2�j���/T��j�@vqv��4P�7Lό�B[�>&Q�K_d��G�"w���G�GO~�L���8�&��x��4�LuS��oX��l����	���Y�vיƣp��h�����o$����j��^�����VW��f��{V�gS�ESqr�V2�I�~~y-�����U�y۔��C`Ouc܇��d�J�ޣ������,��ju�[��z�2��%3�_�~���)�fe�3�r�����M� ��O7�tWu_h��[��L~ |y��I��Ɔc�0���Qqj(��U�fbߤ��xq�Ư�=^�������k�r�n�2�r�#�Wl�4|�Sab_K,#�2)�C���X5�_zt�������]V5E��h����*��͍)"���
�)=j�����������*�g��q)	����<柒n��t���;<GJ]M���Ѝ���K�7+z��98��<�G���6q��	�^���C�l*Q�#*Zq�����HZм@�D�� �D��e���u$b<"�k��i� �O�7㡰/�TJ�p�R�E�z���1��Q�*a���k��l�@k�DRN�G2 ���s��c`;'�0�Z/����V !�����ݼ2ͧ1Ӟ�z�x؊��`}5��Z�A�)���u&t*!|��	1@c˄G�,iN>�4��M��Ǿ�N��X�\�^�ZusR�Β7%`�`G���Y��H��j���:��&���q�5f�-�>#0�&o�<��{�5�$-���
S�C�1�����'k�2�,�����E��N{I
}��)zUU��_S�Q�:�K����;zi���p�tv�'2��1@��,I�nj�/{��mISo�6��K+N��6���OL]��ܸ�����AÉۀ+�GϧG�{a�F�"��/��Y�1�������up�H)����&r�������&�S��Ztꦨwgg��L���=�R�}��qm����,2.*��}��?|�T�O�-w�W۸�Gs��uD���?��%)�E@��.M實b7����2�28�r4���I��$��O��� ������^�3f�L ��Up�����?��9[�(�k�D'A��&�Ṳ��Q�'�.����Q�Q=}����#*v4'8* p7G��<���b�3�w'�\���E޸��G��4Dw|n����л2��T&ia/'p��-5�d���L���Y�Tٛ�*���F�Re8#Wy�+��W��#�n�?�����#C&���}_�~�|j?�Z/�¾ӿ�7ѫ��~����1�#�%�%Z]�$��b�	�q���nh�5���<$�P{ ڭ�j�Y0s*m�����2�	ھ�L7<���[H��Ճ����8Ral˿��{G���
MG��ʢœ�4��gM���9�iN��i�t�������A[����85)+�%�kL?�0�~���p�6�;r�(�s  SY���A~�Q[g��b�|��~4;+y�GsW��o��z2��M�o�0�"番��9�ޜ�l���l/Vz�|2��l�;���V�*h�O4��$���z0
nB�kqؘ</]ti@���l�����'��;�̾si	�\Y#�~�*�5j+`
bX{m�x鬳tH����k����8��8���Ikkѡ�L���]k�}��[0��z��n���8�U�@�q�8+ͷ�g�O~-��PJ��J���1:�*�N������ �f�S�T;
��~Mi�sV��5�k�� ���ǢHA�]2����5�wQ��:�]`��!f�SJ{2�s�b�8��k+����z��hY|��������N&B�r�<~����M�yB�?�l�U�׭Û%����~f�e�ƾ죇x�o�+ɉ*X�Sem���d\4�C�qʠW���*t��ZZ���lҤ7����pB�1���8]�{�r���A;w�y��-/ g<��%�!R>&$_��LPb��N'���N��<��,$NÝ��=1A��K�~d���7)�bO-zD�"\0�fd:SHP01���w��t��vT��Q����N��F#�6){[��UI�:�kDV�� .�1/�|c��G��b�R��;i{���$܇�FŁѝ�2�v$q��,�r�@Var3��?uU����lHTN�����JW��J&񛧧08YE����_�-��=�mk��*!N宮��G���m1d�؁\��Dx�a��B��Q'k�x�w���9`@� K9��M����!:Uۃ=��D��F�y����Z�	�7��Z�f#I ���]�-ss����
4�:"�4�ʝ��M(�,�2��n��$ �00$��/��n$��8�8i�ɺ�����{��eb����%>_oI����yJ9K���lyՓz�GBp;�ʑ��'� �&��F^[���w��L�b�~�	����Sa���l=�����N������pƔ�]Wl2�����!%����\�'ۢ�b����e ��|@N2g�(LB,D ���8��C�h������NТ�7ȵT�d�0�F���w�î�Fl�3��\�#L��v��Ld2�|��T <�I�ل�f&� a�S�Di���5���- �?��*	��P?��ti�u���rgQ��A2��е�	�W�� �g�z���G��(���<ե��;��{���J���jV��8��mc|��҉$qI�%���/���Gg�c��߹�'��W�ֵF�B��x��w����m!W�#`�̕�L�.�t���$���8M�3ʦ���7xd�ӂ���*;�u������KG	�e��>�#��f啧�B��9 H���	��q�YD_$���!�e`���-N���`0*=�=��b���LZ��PhB�cj�h����ȹ�H��J�O������d�Y�\:b��-/�� O��1�F0�}�Cnz��*���e ?�b/�'/ u�*w�el���D��V��R6�������ӳ(1q0������&��/� x�չ�"/UnZ)8�,�7N��:�~C�k#�����{ϓ��3�&\�˿E��p2\㸊l�3��O�ؿ�`�#�l� ���	��7�c X���ۮب�0����3<Tѣ��p��DטT��B�|F?�>&�(u����'�Ї�4#��<����m�y�kk���M.�V�J���)����}&�	�&d�@ϯ[ɝV�� �M��~䧅~@��O�=0ަ�i���&@��]��\�_9�ΰ���K;ރ�'��X�S�
s�{~�N!ڹ�w��*R�R�b�Yڥ���T��~N �k;�M�F�9�����+�0��2֏��*�,δCE�{�̔UeP���w�0z���#�y�r��a�����E*��-P0��y�e~��s�Y*���w�y�;�V����휰l�\���m!�O�No��!o�l����%�3�����ϸ��l��"�n�&�]�s�WZc��n��5��?�/ErZ���,��R����\���J�D�W�����+���4����0��������
�xj~�7!G�m�A��𧥯d��"_�ح�/� �?����N�A�!��r1�p�����,���F���a'��aI�b�ml��*�q����i��A�&�7E�?U�ϯ'��38,7�*h���tz}�7�*A|BR�/�W��N$�XeS꒠D9}�7�@~����.㋪���-��D��h����$L�����P�>�]�8�8�W!�N��,��l'�����/	C�@���T��|)h���x/9yCU�NCu��cF�(�b���i5�eGl��'l�kd'W&�б�%<s���4}��B�ǣgF�ɍ�0��G���xP��$����1��DB�Q_A��X���%_�m����t��1���Su���ˍ��((�A��z;���Zl�����z����e������eaj�裀�q�?��y�u  ArBG���5k ���Ly�w��A4Q���m�7դ�������� �Ve�OS"I���=D�J�����K%V3+�����L%�o�*)F�9 �'��rm������-�b����bS���4ԙy���,Sʋk�M�X\뉏��Tb-�Z�K�K��N0��~5����aed5b��8�P�y���k�)��nC�ɲg�D(�Px3�pXlW�]n0��aէi��[��P�9�<��v#�-u�������ot�R���a��w��s��qI>�zu�U�5���=A����-�!��t���CO�񛴜�x�wL�q."CZ��sw�΀���d�d��.�!��ID��چb�����6���-#���a;�<�P�G��	��Dsc �͚!������̽�1�m��*gi�2FT�V��Y}�1JN�v��Hh�5;"ѹ���lq]&�/�̺���Ce�`��m������H8��(F�P�ZaG���D}�iy�K�×l&'~�KV1����O�]M�;I�]I�;���d7��#�wj:�6`2O�;h�^(�W�$ckx3%S��<�1R��*��q����:?�	�L�.qm���\������jy���p�,l�jT*��b�c��1�6�@�S!,��}��8���|��~V?�5y���p#�`� ��y!�Ɛ�C���ߒ
\͔YO�v�w��6T�u=����� �����AK��8�`�����I��$x٭D{��ꣻ�4�\�J!�>(P��������+�u�Z]$�,rG��~l�(ب�Ig'����B� "�q՘�]p�)'������na�q ��Ո��ѿ#��y��L�,!��υ*��`&������$
I
�*"��"���q{�t��
.���W��0��6j�\}5����֖s�B|�t��BL0m����X�L*�|9�����烅�rY�֞�!��F��n}�7>�%;�}�C]�!���l��;.~���q�@���v�w�_����-/|���gJm��@-�Q�Y�gf���dF�|K�/�ۼy;�g�(ЪO��=fe���4P~���}I6�~e"���n�%���LF�/5�,a&Y�
��g��3sL=�>v���s�Ń��0.��{j>u�wFM�l] O}�T�(���&i��# ���go��X?�j=��x���C�gה
�H�ه6,��*��!E{�.UD7����(�|��M˟!F���7��)�D����d�=���*���t�VM�m����O�#����3;��'1�4��z3��E�f��~A�H��/9��-P�*�6k�]�%?Q��X��!�e�m~p�,�|@�v�#��#:�պ�ڔ���u[��8��T���tG���Zì=��	�ݐr�	���dy�=.J����d�C�F�ekPmo�M%1�5�ؖ�Iu8�e#c�3���o�?�d/��A7!�5[P�|�ZK>'�`��I<�A���D	��Z�UQ[��A� ,�	�@�,��������j@��"8@�M����s�4��`qJ����\f҂���Q�{(�¸���[-�� ����S��q,Ȧ�_�% �����Ep3���6��δ�Y����os� 	1M�{�������9�?��y�_�7��B�����s/*�Wf����"�������y�fi����,�F��ٜ�~9�7�A
��+t\�
.3���5H}����OvIr̆���a>T��ԣ	�ќw�����)�W��'4.ӮI>���/Z�f��`1e�m���f֏�A܅�HNP�@��ڭ����]Y��$�h�%�ю4J>�!�E8�E�@/�_j
T�#v�/�{O�UQ{Z_�)�[x��={Զ�*k��ku�H�ݴk��B��64<\��0�o�V��S�[� ������Ln��,�	f=�k�V�5�dI��J�=�qg�$��e��u�*��x�C�q���l��r��K~�w̷S������f��A���Řrת�����E��tZ2��؂D�]��l�H��BP���Q��+���v�¨��=6>R�,�m[^�V4\T�N(`�Xz�ڂ��������F�V2�����AB��1]|	ִmۂ28>�+"j��\���0�DL,p�;���yߦ��l����ٮ J�n2J��m�w����
��b�Uw/e9)^L&05�_l�au�8�#��^�|~@8o�5�:=�/h�p�J�Q<'od����,"����+����{џ�~h��e
r�3"ӫֱF0;r��%���� ���v�r��կ�{ (b��U���w֡D�|�,S�/L����%l���E|/�1�]Š��Ry|S��)�q�
�%�6Aukf&.5O5�_��S�Js!S�@�2碃Ds6޽��9�z��tF�z{�̎,����xqH5���1���L�qF�q�N`��Cݔ����6h24�r��;��F�CR�T��7PK�H�:�t�o���-�v�sg>��E���A�����K�;	��L�2�ӑ3��Oƞǒ��:�)NsB1w+�Q ��&n ��_��3|7�b��!/h�\���89'�('�P���urB�j��z!.��#�ݙ��}GU�6���Zbx��ym
�@�Z8I���O��4E
��Ǩ�+7[%z.�U[R`�Z�A BnY&V�����]�g�MN�ʔ��[S%�n[�1�|h��%��I�/�7JQ�K��m�?js���,0+�Ja�%�|5�CI� 0ǆ#��`�C�qe���9��=��p[��ao�@��!���
��%��"� >{L�ª�!_���	�j���5�k{�Ne���� �o�o4]�p��(.&�����H�`�m�e��/8$����:���	�T5m��7t�l�o\8YO�G��ѡ  ����ۺSW}�%�����	V&Q2LQm/q���{MW��ء�[@� jU�q����D�H�R�WVw(���T��� !hE8�s*�Op��K��G7�胗�o�LK��؊/�#V��vE��y��o�/	����`%;*�dc)jI�U���I��ޗJ�۸��<��&��C�4��	�̀n�u������X����0�����i�+��{e����i��=V;�~
{��
�޷����ʔ ����@6Z٢������9��Ł���C%(�FX��JwѤ�ų�8�̓v|��GV*��8�I��|��k�L	$;��7�i9G���������x��K���tc�]6��:���9m_�Ĉ�.q �0����d��H��<I	��%$�k����|��&7UN� �չ4H�>uu�r���)+���W6>��2X�w�D��!��m�,2:��xZ���kS	��3k�b��W�։�:�LTD�m4Ӎ�봷����ɟ/U�iZ�{qW�
/�)܂ɪ��*�v/qqKB���-���Vԝ����Q�wpf����/N��4�S��x�9�����/�~�
�d�_�1O�Q(r,MA����b��RP�%�Q�v-�%��U`�kF��VHuMum��wn����?��MD�c�C���¿j��e�z���?*�ͬB���EY(,-C@4L�[��`����c���?!��Gl�R�Hr�u=]��,�U#���F�+E&o���Z�B�q!ŸD7_݄����:X7�ua��g�U&^񬧳���洳4*��l=eb�v�O�=>Ɖ9J&ĸU�m�� s^�A�d��Ac�*xp0�w�V@p�� ��ru��5��*.�N�̅��hl�=��k$�p��G�˴���Y������_6����.��,�nL����)!���������z5ӂ/�I*�W��;}52�"?�d�F���<�E���tÑ���ѽjb�N#	;�Pg��b���?���k���[xQ1ۍ)顜`��>�"�]��;��̖c���Ӥ�Gرf�;���M��gٶ���eg�n�}�`Ŭ7�+j3�&!E-���Ͻΐ:��_-؇��)05L�t�S�C�^2��KT��n��$
RYo���꘢%������<�%��Ьĳ��S|"��^A�Y7
�.I������V�S+�0|���ȣ��_���MCQZ��"�|��1���t�2b��Z$H;���9���Um�B���T��Fb�<7�N1��Xz�ۓ�x@I^���7K��-VNϾ��6DPR�9~�r���
���Ԋ�Ek�����-=�l��U<�E��Pl]1qO��c,H%�"���:<٫�M2�d��zar��r�0�FR�qE6<n�����+�	��Ug���������1�PO���ƃ:<���+/v�F���x+g��IK�>�Fx�DD�v2�ϖ�ܖQI+�^K���8��l��޸��ސ�`���_1�A$-.&Q�W�~X?n|V�仓����%���5��q3�J�����3,��r���V6j���O���|����ķ��q\�L���������9U��7�h����)�x-�ɑ�o����jQ���@`����!�R�S�{^B�A}:��d�5q� �1z|I/m�x�������\�b�0{8���@Yʬ��^6�8oy�� z��1�m�E�ˊ���;巀PK�yJ�������(ͤ��HT�:�{S�	Ғx��l�f���7:
'/�
�ĺ_[I+����pf��{���4FP��!�m�qưԞ�䶕)�s�UG�G�����8lJςY��{�E�� jo_ߍ�|��E�ã��"�[��y�� ��ɱ��:|�)\)j<���\�d��X�����,�hɑK^��`$�Q��� �.�A���=HU����<b��&Ձń�z�@��pVw�q�i�I �7L���#��j� �C`V��*M�D2�*! oA~��{������,P�t���_:�o73�4��{��{�|=�[�0ۨ�reu C�s��I{թ8�����Ƅ쮚cH.��q�������^��ď�F[|%={6�`���G�Gیx�ƾ`"��@�~_K礝�R�{��2LrJZ3N;��.��+.CNc�e�Ծ	:%��8���,�/YY�i�.C���e8+l$L9Yʹi$@,�a��^w���.΅��>,���.�k98�;?�f��\�g���]�O�����=��h:-'s��xDi�cn��U�<%�'Q8$/ ���1�d_�^$�I�Àj쏰+H�I���4��[s�#l2.o�0|fQ�f3
�z�Y�7]�}Bv���8�Ջ/���!j�3���F����n�z��b���f���U�@�=ўf�z�J��0��R�YH�ވ�wA6��*о����gc�@��p��r7��R���Z�xH-x�,+6*�1<iha�J��h�l��3̭�+��;Sv��X��D�^wU�|t���ϭ���*��3黍�W+�E�ɓ��q���p1�z8wz.>B[Pis�s9yW4��N�r9���$Ĩqx�_I�f�xF�N2u7�t�B��K#	����G��E�(����RkG�*E��T�v�P��;��� ��ۤ/��U��K�	�9������f d
���F�1�䉵����*	l���i������԰����J���f۞��!qbc�U/�NrI�?L��fD����3�:�����Iu��=,9�]��A�ֽb�$��׏nb�(�~���4�L��e9D�C	h�Ko��]-�l9��e�sAp3�g���D���9�AmE&�o�]ڨCF�)ކ	��[5q�aR}��&8Lϥxgr� �BG�\��j��؏�D�����-��Ո���V�H4]���HLߏ��Ka��@�%�'�/R��'���;�ͨ1L֓�Sf���ư�`.�����`9q�[ɹ���$�E�;��� 伊G��>�(�^�ٟ��X 3rɎ�U�Y�9���.�(>�L��]���V����kpJ�����.(]�,��z`�4b���_oʚ���!r�[��g�ڳ>;v�ΰ�p}��I�3����*�*i���^4���Sg�Cy����C���i݆�=/Q'x�4<(s���=@���0D�yy?`��# �и���j�nt��7��Ѫ)�u#����N�+�Qr�2�<�oRbp#������|�7��`�yHb��m멺�c��ex�]�]J�����Xo�7O鑺P��{%��+�Wv.��e$a�Z�_�4ߡS��C�	'���V��ld�ЛK�u^�n��?^bs`5���=��d�{�"0�pFm���_���3q��7u�k؋����R2P��=����J��C����E�@��u_���Ib���������r۱:���Eo�5����og���{	��O)�]��}�FQ������3C�p�ǽ`J,�ap�5y2����+*�hҙ��vw �]J|�7�`��(�����^���:��G�.t�nL�̐��7���\��ҍ��1�~�Ya/΀���
?���)��xMD����=��2k�uh.c���sF!��(Ҭ���%Ϻ�x��B�|:��"ߋk
�@�˥H;�s]YYyLF��a�j�c��k��c���X7+����0���~/!��iF3ˠ�u[��̵����(SL��آڬSݟȜ̴�	�,f%���M���x���K�70eW��GJ
��k��'hf`��I-3�X9������ֺ}�A��"�f9FcT!)�����ʘby���	e��|];�^�Zx�e�Q5='�7�8����M��b:��'�(����U���y�2�;���M�A�j��M��()h��Ʋ��H�J�T]��8��4pǐ�iL��Z֡�~��"�Qgz��U��@��p�]�/QT�>T>���{�gb��9�����njt��ب/�kG�ɍ��N{?3��x[
����V�ȅ�ѪG�YA���o����ӽʍ�Ț����-F�|��w-���)ә��GϷc �w9��"���.�vQ)H�(5e�y$9��첱֜�$���6Ɣ�,���o}�0y^��m-��u<�}���m��Ğ�ᆹH��=sMn�����Mh�����Fk�RT��XGl]��*��-�}D�C>�B�c�O_?��A�^<�!���lLNΑ/e9)yv�"ו��"T���X�b������t�1�>�֯��6�1MCԳF�k���DT��쪷�p9��:�yA��NU�%�h��$;�E(x���.����)�8oR �V�!��&mC�'?�?	ԧ@�N6�5ًP��+4���j�bG`�ʎ`�Hۊ}v�1s��Sa�1�.z�Ф��,uQ��3�_g�ӭʛк�͛R��u�
m{A���B��:������K�Ǔ�/�Q�����(��-��3=y{�������n�~2���7[ce���
�z6�Sa�aIOv�ځk���+u���X���&c6��B�B����Pha�<����i�F�{6�5�?���q�D�[�F2$7b�kH�B-�uH6��,��澀e.l��;Iov�je�s��W�2�R�ķ#�����Λ�G`��hr�t���\��$p�	�φX�`�c��h�C�����P��E,
 t&��-T�����$�����ĽB̶$p�����Bd�>����-m�(3����3��ꐶ"��qߡU�XJ80���쪑�9�5���ӷ3֤犕ҋ�76�}�{f�hs�]�a%���lε�i�T�x5�η*��fc�D���A�Ԃ`��43��
�#����g<�v��@\T<�"���N�B:<�5͏,W�>���Ӑ��?���!~���]D1Ky�a1��f�.���B��Q��t�twpu����֖M�{?9��{����󉰺*kZk�x�&?i;��%�,�+�翢`9�#wd��A��`y���+Lmo%a"r�vܥq4U*i��	YK�p�E�5
�A&�!�3�U�Jx�
���mp*A��ݗ��a&f5�5k����{l���&�x�H�mm���^�-�f2��P�P,����X��P�_��Rwt}��KSfˤ��M������_��^bg���/'�
>������X����~�	N9C9��5������Tg��nLk���}9/I�T��=]�z��M
$�����0�f�ԑ=fZ[�b�����i(��r�b㎳WB��t������r�Z�o�'�]��K�sbhyj�
xF� @�6&Ǩ�$&��S}Z���@����)7�_�.rur65�Z�P5���5��a"V���j�.�/��ؠ0����Nj�|6�V�E�20(��#������[.���{�+g��aO$�q%O��������1�h'ą�[��F���	?��54E(|>�,G����h�wNaI�/\[��8/)
Yk�������>�zt�A�\�^�Ed�k��.��l��(0Y�J�P[�����p��p>��P����?���?��A�+��B����q�U]��i�E�T?s���k7
���H0 ��I{*L���v��9��?�MmcK(�{]/JU�1>�8�s��35����j���y�/�D�->:�h���H��L������`��>�5�"g
���Eg�myc���)���$��دu��{�p2a�(�ݭ���^�v�^=~5�j\(G�+6U@�mp����PXR��)^��M����x� i�0?	��:��z�l��[�1*�T�Hs�5Y��3�צk�o*�%a�q�{^w�u��>L\_��]�-aUP�y� �d��ce�'���G�?��2^1�=��S�z��j�P#@ޅ9�y��o���ɚg:�*ye=���3&�>�HlR�I_��i�s� ��6��M�����SҍAʪ*������ǆ�X����ZI�b�q7<��q b�"�f]���Y�?u��Դ߂j���p"��-.��uRg�0+Y���BoiC���#S�i����q�-O  	�0��L�C��X�l}V�Ҡ�;p�ڸ�v�)�|��oJ�Pru�G�%L�&*|���gT0�JQ�����I]mw$�"5u���.���c�7����.]Ô�����N"L�yWC.W��Ԣ[!��V�G2#Aɥq�����t�"x�G�Ҡ)�7Z����/f��9N)n7qSN��8�u�?R54/�����Q
�TqN<g<��q��j�9���P���>���G�W ρڬ��g��`Q $&f�xYj����W:�l��w��L�$e�����T�m"?9:`B��y�HJ$��s���;>�������s�n�!ͬ�,�	0���I0>�Ee���*�]C
=ފ[ /�q]f0k�}�G^��1^�}�.�M�57n�D�"V�Z�&�"�5��؇M�&`I���2Q�ym� �ݡ��w��=оȥ)D��,D۞����l�p��DA���Z��nk�d�_4�<�xc���]W��m4!ٻ�ECl6��)�-t �%�Pofy�R~J��?��U�ǅ��;%��	���ƅ���jA0�_(A�ZOs���"V�j�'+'Z����p*7����ƝV��:`��1%���������M_� X�Q���xl��&��tw1�ed��������$p�}��V��J韰���EdĀ
��+<^k ��lC9�֢�����C}M
G3_+��& ��|�1�����ˋ-啗QCͲΕ|3�EՓ>�l�D�Qj��u�J��
n��Tfd� ��)��t�2��:�@��2�=�/���O=hI�:&ߩ��P���O��,��4���_.�~}cʍ�Ԩ~��0���>K*�>	F�/�� ڇ*�Hj�}��N_ۊ����}��4rg=�4(��vMga�2h�k�x� �'��{�>����ż�o�*g�ڮm�%9����J�m �aO��']���bb��W���Zi�us7_T�#�V��I��,�^����l��iD�ٳ剬(򴣡u�͖��B�$m!p隰��8 ���W)(�����֏g�8���]��]�[�Dֵͱ\�]�M ��B�R��6*��	!��9��e�꛴�}Ē�E���׶��.���2�۾�q�H-�LX|B�8W�������_K�W��2��ɂ��&�@VWw8Δv�|'A�@��2t�h4���,��#�#MJ2Kц�����$��Q��������I[���W�>ÖJ��o��[�
�Ф%ا�6�w���Xe_Iϯ��'��č�ә�%���HH*�i|HNBR�̀71��N���2�>�P���?5x9��U�6�k��2Q:���(��G\B#8~�YNr����vJ�e;�3�I�9\�W�U��0�����L�F�}�BJx�[|]3�z��O�ʐ@��V,��x/]D%J>>�dթQJ�9�$�;*Hw��α�ةOP犯cIm堿ص���)��ēҞ`>��"4�᩵:�#�=��Ag��H�4������"�)�D�F�n�D0�+�.���΅E�������E����Aǐ�-؋L��T�V��V7�x�'(�l�5͋���W�w��)�:��[eʂ�~&0��"��ҲU�5��9��\ZNr����z������O�En���b��D{���a��J!'�4Ѣ(QB����qD����Qu�J�ꉎ���ד���أ���I;dI,�3�ʎ�H?�$:�I'ݭ:�	���vZ)��c���壙.̤���¿����5��W-mU��`�Ǩj)�}Qm텣#$�/UX5fﬤ������z�Kh�-���=��s{ ��0s�������R���ǫ�C ?���� *X��Lh�Y<���K�����׃�n����Tڌ©ub�7�}*��&�t����c��>�a2�;��x��ڶ�e��^:�}��W���'~�r ]�W�����/Y������d�¸�n����dOC��<��B�n��:vM�fuE��iAUH��Խ�~�B������V0�r<x��������Na�Q�4�_�<N��@>��`J��[�Gi�����@1�8���6��[ �����8El*����	��ٱ��3�E��7��|�/d��Ky������?���1���+V����*˴(Y1e^��lx3�9{~�17g�~�E/)�8,�+\pY4L���%�-��$u�zh�g�T�H���Uğ���<�>��Q/&߹�p+��>y�q�*��P��F����i�Q�R��-����ق���`��B0�!���/���7JU3IZQc�6&�|��g@r�zS�=.�����p.��z�;�I���(įs��d��.��7��4q�sۈ
�Z�]������@<i�g������D��*"�N��Z�';Ss���H���̟Ô\�vLW����!'�nݤ�� �n6�1@9^�>E_H�k;GXOj����Z4�Cb��z�1�s�O�.H��b���5f9~���mE���x�c����qb=��fA�EO�)�CES��7�O���<IG�O�9��)soꧻ�H�_J�t��xي���y����e��2k�Qaq�1�T4��O��Yi舚�/WCW�J/�»�j����f�/�����4z=��m:�b��ԾU�$T�*�im��N��e;��aqK�o��v/Q���A�1�;��\U��5��`P�\�Q�?ۣg=��ۗ�����M�3��*�[���;~?�\�������n�$Fx_�?�0�E ^�o��%�n��~<��A׍�J�F���[��DY�34l.��>��Z�P�=���j�ln)�$K��UǮU�_e��%hs�Tn�q<�#B��@\:��hh��jY�v��"i��ώ�L�lj��],�u: �k9�rF!7��ѻ&����RN��!Y��'޺lV�9����O�	.��٠&(�Y���ԏ��8��K��$TM���t���MA:j�G��V�(�Vj��P��Om�?Z��h#��@r��_��^tP�E#��U 3�]�q��
p�K��'r�@���X'I<6�q,w>��C|�����¾��s�V���3�'���<_w�غdA��M&_��xT�{{t��B���!NZCsB�R�3;à�&�S���>d�u�A���.k6����i�v	��pK^~
�#=y"�G���+�
�����#��&�W����(n��G����!�
X���T�[U�����IS歆�Vf��Z�G��a��� ����yi"`�`�Tb=�Im�С�]�d�oH�'���5p��!M�_�M�ẋ^�y(����õ��1�I;����_v`�x�����wr���*K��]����<�U�t\�>P��/ЯB�d�R)UUY�l�d	��'�j��J^O!�s�tE6\�$��^��3&Ls��u�-���Lf�w?�/�)�2��zԌ�+�&�QD��=l�`y����F|����Z�p�NV?�&��E�j&��]��Cb�D-������8!7e�كݴص�j]�������!��E@�7B�i��W�c�#,b��@t>C]`o�ϝ�ا߈���ev��㣔���`��P����G��GA�q�k�K�a�4�!m��z,!������f	�V3pUd��f�IMT2+j�P�f�SO&\��Z��{r����!x�F)f�����Kf�r1M�W�\�~�/��<i:���o�_���i�uB�zD�.���`�zx!��]ﳥ|�=�����k�2n��[o(��PP�C��z0CA3G�6B5M%��dHBRZ˪0(�o�T�9m�KV�k��W�<폷mM�q�O�MivgfE�&�~�K�������;LRH���Q�M���q�$�v\��S��5,uo%5]@�7>�wWC�qfh�א�Kֈ�IpU�Iڔ�N�@�����(�����zX��1F�2^8�l���9ѱ!I�0E�B���E+UR��L�Th���u=�pu�R��0�]��z,��}�#��N����N)}�ۊDD���w��б��T���׻[-��CbP1���������L�[�Jq|�x:"��q@v^GzS���*�-E�Y��a��m�V����}��b_}��a*��R~Z#��!Hԁ�b��ڲA��J:�3B6J]fa,�]�����x`4x��t�p��P����~Zg_5�[Xss������_)�|����vH�%��@��hd���_��-���͎$8�V�5�l��T��[24��h��1M�%Ba71e�����8G��!cq�y����5T��x�%w=	�!�&�����$8B���,�Cj:<߀������傱9�7��Nk	�f�]��xq���-џ�$"�]g*�����\��{�22�����Y5��vo����֟��B����#Q�C�z�zA���`O��t�m;�#�8A�\M#p	�8���V�ǆZ[��l		5�|��Q!3�=�$���	,�i�Dp��X��1=�K�LB|8�xJ���Ğ�����Ci�κ���I�P������?��׸�գ�Ug��<��Ϭ!�	�)L� gu��0�Î�5灠i;/i�h�92][�OWiK�11�T9gx8[ǹ��|��pi���<���y�g���c� o����_�5�Z�T*�.y�����9S�����v�v��o���=C�s
1󫁖�ԝ4��q���ׅ)�9���O�B�N�8 �Jw��R��hP��d�j�AcRh����-�}r���10����ܠpgc�l��8�П
dP}��>P�L)g,�"�L�ǥ@��[��.��٥�aa�3�\c�i�mg��<M�-�*���Gd��G����LS��)0!�u��.)��Q�/��$�O&6��?���"��"]�*�+	=}%*{lJ���%���P��1_fL�����8��M[ݦ/~�f��`o��cmî�<l,���F�F`Y d�^�yg�s!P��O�8��<�{O�_B��ji�]7���J�_��D��%V�Ռ���s�xis>��r��ɽ��/�t.��kLI�������9��G�k�O���A���+ ��2�۩��L$1�r��+>�|�����/_xs�oӔ�B��1x��G����G,!��n��ǡ�K˰(�Ƴ�RH_�x�גn����c��u���#� U�{@{�e��oћ���(�IۀL�\�׿��Szj:V�����C�R�K�%��<u�q�Pu=V��N��j�����^�U�`�`�?�3��FE�FBU���d@�NC�k̑�s�>[~�s��UI>P��R�}��������D^"	7���;8�~S7��s�a3���(��{�3�t�Y6$����P�yM�/�V� n�+t�ہ�j��Z��>��Э��~��Ť1���p�MU?D�_���Ȑmwcެ=s�M�3���g܍���fkr�&v6�.�c��rK���F�=a�y:ȏ$(xo5V�+�B���w�O������^�r_�spb<]�>��0�?۔q�"�][�������(?��9|9�up�g��î��9�Ĺp��,{��z3��`��?�:%����R]a.��Ŀ��4S>7��<0���U�Q�t;��7~�1�nU?�Ap�ǂ��q�Z:ꮟ߳�*������*��83�c����G��Y|�eZ��#���cM{bdK~bSfsæ'z��xy^�2�#Z����(]Q7@��� �����N@�u�:Sƕ�]KJ���3�o��p~zBe�n'�Y�2�Ԏ�/��@Q�h��k�?N�Y��Ka�
���mg�"������$�]$����+)]�����C�|c�6���F�p^6��Em�n�2n^N�K�dE{�D�w<E�5Ϸ��M�`�e��B
t̰Ԥ�D4����p36t����R�'p�r٦_��v�B��T~��?�15��Z��T�ZO���ZP�C`�H#:��M��?����ݰ��b�Mm�o�P
#-�����T�UQ���TKu�p/�h��i�;�����y)ޢh畯��[V��Φ?{�En�� �g����墎�2�]E+z�	_�R�������&���US�L�pWW�^"�r�h��i'h��9XR�7���,��ٲ}㖀L������܈�e1��혳��f��B_���PH:�&���g�՗˝�䛫&�s$�f$v�8}i�!�*�!.��M���B)�$G9r-�*���Ved�㡌���M:�qeBev�&�0t������S�]����zg�䯎�ú6�����n��3�f$�����8K�m�T?��o�;�]E<H�$"4`���G>d�h@�3�6��� ���q�����g�Ԥ�� �椂�j��|Q���]As���M�\�������F �h�b�;Ǹ��/��g� F��=�e0V�Y �1��ڷx�a��Jd�m�כ�6P|�N~��|������K�p3�Vge�����1���>�F��T����[�Q�c/g=�K�Q��`���ɣ��
@�Y�q�hUX�d@�ц��T���~I}�Fh�~~��mn��A� ��T,X*ihuU�E9�g��.L���%�Nr�����"5َ;�@�?�%E���m�9#��9a���N�w%"�p�'l�\�R���x��!y���n�f�
�Ԑ��.#%�K�v9��!������gՙ��E Rl�56-"�>��bm&!ܖ0�^���)��o3�;�4��k�����`�������
�"=�)��%�χ~�����Q����E��4v��1ѹTk��|yr���Hy������̹[��R�
�on��"͗�xi����J�"�>^0'*��M�֎q@��fۢ�)$�ly�qRN�}�@ޮ_�]� �U�/���ޥ�����!���bC�ͩ�.�ab�X)� ~���}R�y^��I%�HyNN�>/�O�KvҖ.:iѴ}�*�
y)%�	��P���#0Gp��������:+O��C��*�����Kr�\w����<3�a��l����U�b(s�����^K`�ڸ?�y$"!z�AHj���c>t�T#�l�h�(	�/�x��Zf��=D�ɫH'ɐ\ϡY��ppj~J+\�XpTZ�}e�^!�������jb�gXk�g���)R��AU���4��N;�7�wiz;�,��\K�����YPs��l�ՠ �7&��K�{�]2�
@ �;&?w�I`E-�v�������,o�<f����!���� ��; =R��d��4U�J��i��ԡN����� �#��������x��	����Q�$�uڏ�����`��:�|ae���F>ZB�����gy��F�@iKl5yZ:��\i�K���N�ua���B���{?>,m�)w[�c��U�����xB���(湵�2��)W�t��+~��̑�{)�V�Q�[���8�����DW��H�w�.Fe��Z��f�N���OGD\���ı�V,׹�4H|��y�d�&4>��5'��h�=�̼�%�4��َ�EXF_⟡�vep�un' �7>RB9l~R�E#zE��'OG:l�������r�p`E2��r�s��k����?����1�ⵛV��`_7?.`ӯ���I�֝�C��`^0���Q��^���F�Y��6x=�~"��=��Q`h����S74'�.�۾o�<�)��8y_�Rl]���v�<�F��`xN=0iV���y����eC�߃~f�wWgG�h#�^����� G;e �[Ln���h�����s�h��;&���3��g_ �#�qp�)ml��붑MY� }��[������Qx�=˼2��������O���Ty�k���T���^|���rgO,��芔��"��l��_RJy�ح��v�$��zףY]Q�*n�ϓB�FgB-�J+JYz�y���tF�������0�T�'t�eu9r8�)(U�p�
>�엃�Rhc\��BV���9Szr���j�~�2D؞p�x��W�8�e��������u��?�5:���H�C�B�y���-�A��-e����Ičx��ʻ����a��r�>K�c�Q0'�>U�I�.�_�9�.��f8�cpc"���O�S�Kn7����� &3�:l��*ShV���&����'x;̬H����o� ��<L��;M�}�f��wU�m�7]c8��4h��f>��C�5{�Xk��a'�d�l�~>^�I�$ϟ�c@aʺ���WmwP�&��RU�N}�E�n�T�6.P�����:�d�y�{��3�"�~����N��^����I.�P��ş��^���?�'E��:����#dH��ƌ��]���~��'����j}���vU�d苝|���dN{6�&�)9r�W�����$�I8*�A��U�����pAQ�;�c�V\���ϊ6iu��AD�WI�T�ў�����E�=.Y"�Y��Nh�[�{�>��D	z�Ƽ|d�a[5�ǒ��,,_e���S\:�Sn�ir�Jf�x���.�*�1�[�[��ϭ���U@`�=|<)e�-X�w��$�֖03$�z4�k��(�!� �@�JM�e)'kݺ]KU-���6�44�R�O�������z'.����A< ��a�w��&�}=o8;���{��/9�Ƣ�_iR��sy�<��D���k!co6��A*����G}T�p$#v�Oפ�0浈�򧞎cN���8Y�z��1)�Z�?T�ü��q�h�V0�LK+�`�VSrI�EE!�8����m�*�\�|�nԦBO22Թ��Z�SfbK¿��oC�c��RLk�Ce73C��[|���)H��T֢Jy�6A	�[���X�c�Q�GMj�(�K��}�Xn,h�̚Ic�<!䘽�O	?��z[�/����_�G�����~�,�[�Ch�<��2�(YF��ճ�α<w�}�h�U�]��P�N2�E��Kz;���
)�~�ېђ��s��h�\LE|��q�л&*����Z1F��0k���r���)�r�('Rǉ�.�ə 6�Q}We��� E�~ ;��x��6���[?"�,[�¯f�r� =�S])�Y��� ��&Ì�ñ����7�v ��IQe�>�� zlH���{b ���'s���G��C���=�"X�A3��������)l�3X*5����n9����*Lfэ���ɻ�0�{_E�:�e�q�&XD�����r:W�����_���t�S����R,�&>��`��sO�7�J���[
��Vy�	4wo�ݮ��w�����q��	�ɓ�>LfH��O���X�#�M�[�v �gV�l��K��f��8���M«�?�*�_a��k"c]
���k���Tm@�w���B�HC�ДY�W]�|5��מ�0�Ɔ�k�&�^>��,&SzG�W�ȧ!��z5D�:��N���>X�
�1�7��|���JYXR	/j:���~� ��XX&��*��N.Pɞ�ڵ��]�1B�W-����e0�W�=��>8��{t��[�>Q�������bk��{3&Hq�ef�r��/�>V�(I���(�Yk1��ph�{�drz#�W!��c��E�S�~ȡ�,��.�S-�i`������6y��%�QO��7vw�A��j�A�t��S��_��ܾF��i�ɬ�E���l�=)���̐��V��3�^���_<x?��/x(��Y��g-WL
7<��.ҡ.�nb�S`�o�h�`_�j%OPV�D� �U�Lt�������_�(%� 
1���i�cn'@:�fo�lo����O}����'�Ŝ����7��U"��b���S�6�s���4�L�#T�t���Δq''����٣�	�(M����;�>fh8i��j��М��^_ל���v�3T���(�Aj�3|��� �x�C}E:�9�l��"fK�7��O��)}�n�Pb숢�$��:㲅�qC"���䯨��/�3S�H,��,�[�'��.1�W�Jѣ�G��F�3����^���`+=��+��xjKu��		�����
n���_?8P%7n���8c
��c;� ��u�I8fj�J�z����qv�rz,5�� SqV/���iNIq��#��h�y�.ͦ,n�c��E�6�éҤ!�2as��j��ܚ��'*0!�K`�}�Xn�,��9��C�y��4Z��8mX8��d7�ڏ%��ň 1l���v���J���9nS�W�5�w	,���3�d�j�T��%��.�'������`�@>/>�tM�)$���<��? ����_�`��^V�oV�ٯ]���ƃ����oX��Y?[�^Ed��&��d�]B?Nh�0����AZ(�㜺�	/��v;4�2+5�YT�2�g͋�����\�D�A� ��z0H��z�s��o?���7�[b�&��.C֩s��|+��Q:�~d��[�m�s.��07����c����9��;��G�&CC��f^�
���BE������/���ӳ�E�U�Dﰣ�xn�aUL=�@�����t�p:k�Xh�a\`�K���ٰ����b��e�Ă@���*�T���,;����t�T,���I�@��Le�2"���C�nݝ.�04��i+uI��؝���e�m�4yb���&�,�ʬM�
���ʤ�O�c��� ��� �S0���� �Ղ�M�~2�5�*�2�K_��+�GW�:����C�z���hܺ6��$)孧����g~f~7_�_V�U��5_O�*�wMB6Ĝ9S�:��q�G�6�#T���Z��3�� %Z�PJ��}����Z�Xi��	}�D��s��5���� �C�5=t���U�p�˺6`�+8\9����X�K��v1��T����왫;�\]��V�??P1��2���lt���/��)BAd3�_�;���3���;5T�}Jz�n��["3���b��A��(��x���'���̾\�=~�=y�.,d�8[�h;��1!9GP�\�-�"'l��k��0|�E���9�KA�U�V~���"s~cf���c�u�&ӡu�ib7���X8��z��sxv�
C��(�V���4��pƣ���_�`�i�V�l�� ���K(�`�L>�M�swR��[�=xXZ�$��/�HGcD*i��B��bƏ0���1�HM���[	���,h�nj�i��5�� ;�Ԧ_��>Y��:3.�7�	5����G�����W�8��RѩA�ء۫]�׮��w��dW �$�B���>���e�.w�j�g)��j��>�pA�ͬ��XB��
���E����w�Ʋ$Q��xI\���K� f˜XJ��\�������"���8�tA�1ۮLg6�E��f^�{m4ŏN� �Ώr�	蜱�%�O8�=����E��|B�ӎr5:,;;ʏ	��]�~�iJë�M�jtE�c��9���j}�A2-�0tGj����_�v�	=���l�VIn���){ZVV��'_�ǧ�ٻc������8��G������,�X�����+�<
7��>ҐTYw��<�U�"�C��f\0��m����`n�͓�N�l_�ɦ��$���Ԏ������+4�<�C��q��/�;��㏉���X����'[��п�.�:$�a�w��i9��Ԟ�4L�t��F�O������K��{L�����NN�q�Σ���b����m?�y1�ykRR��a6�46-�^��8j/{�oe�.��Dod�.b����N�uҬ��B�?عgd#����5�YF���������]����KjM��?'mZg�Y�� ��$�)�K�pW2Po_'T�gߤ8%�jn	�����ԭqJnޡ�æǢ_��D���l�������9��5�ߢ4����F`�O�:���}e`�{���#���+:�*1x4�aL�꣤�Ò���K�C��Ut/f����������Hm��5/|௬��]��{,�(vz_m�쪱Zy�a�+��7Xrt���p�7Ҩ��au�-�(�W-˞�YzXj�5�^�$|�p4�����{��grNj�ϞW�)�&'��2�%���?y�	]2w�z�ݳI�6m�C�44���p�g��k������>�(zd01�=AuC���.)S���iI!n�+k�W�(vq�Z�		᷐eraf����s�54�Ĥ�$���?DڸO�ޖs�VF:%���⥭8���N�pԆ\���u�v��7R���8���Л�	�P��G����|1���
�W�%��2g��N��P^��ߏ��ʉ�M������{�l�3�q�$|���LYw`�sF$�e���Q͡}��$��Mҹ��/tf��h?*X�D �\;o����%�ڋ����P������L5�9�4X&'^����5�Ǔ@?+e�
�;��n�L���Ag��s�*�[��4"	=bQ>�?A�cI������Ќ)�9L�Enp��O+P�p��);�!�l�R`8�c	�×>5*���1�����g(@Qk�$�7�̝.b�U�ʠm�4t�4L��b�N�c��A��9� *P:-ܝxzI[��-S?�/_�=�iT �����+�OM�)7�)�������&*�u �T u�\�����|��K���$�moW ����ΕJG�+�A��B����3���E��?�4
�z��&;�q~��1�y�ӣ�0.`�cg�u#��0V��Gf�ߨ�]�H�SO�a88NW�}�]�=���D�����t��D�U�>�=����G�d���*�ߙ2WB0�J�6�M	g��*F�ثS��^����k�?����0�L�p��֟9�|J����*��I����C��� 7�Yl?R�2�Q�����׳����[�0��������-��D(�~�x����^\^Z���b��D��R>�d�@>�F������rbqP�8����k��zQ8o�9�lp�Yh-D_1�G�,�F�X�Y
�1
�7ߙ����h�+:Y �@��K���~ Gt��Rv#:����(�Y��(�Bu�vgle3sI���W�ώ�3���q<�Vj�2DZ���
����ֵ���յ9U�����%|Ĩ���rMd9d��nx���������� re���ㄵ&p�R�Y�	!O���m)�415�O������WW<��wR�.���qJ�}?q�b��b�tK{r���V�p@U-!8}@��w}us\��	����@|5Ğ�
w�/�=\��0���m}�BPGI����B��`���6�!�u[���a7gOAz��e�xu�r�D�y�пI�)� (��=Z�%y����[�cJd���ԧr3 1��ԥ� ��(�ք�bX�ܺ�T�"U����J02z.Mp���cc�E` �pD��|]�q	I��,jW��B�n"�ǘ�H�+��S/e=�ކ0-<gP�v�W�aW���A�E��צO��s9���O���n���t�7������h�Ϸ��ml��|�B�t�:f����A�����.
#�,�
��a��_8��1��{�N3*��[��r-&�hZ&DT=|^!��^��/���Qc ʊ�����(��y;��������h�)�V �d�B�����p��;��6sr��c�����KH~𬰽R�!�3�e��3|���jw7��
�>L���YNwx�*=8t
8Wj}[�u*���_i|a4a��z���[�o�4�G����?[1^#����~+=o�f�A���[��P>քOX!��]�Z�>;�9+L)��#$Y׬�TÖ�����ꋜTX�8K
l:��=O&E���x�m��KOr/�r������ �"�U���k§U$�ڥ�kⰿ�OJ��_Zx�[�A~2�
K�������(�-�<��K~�`�I��.�i� ���>�$��P+��9���OwC�Ԉ�����Lm�/�WAD�lOF�Z�&��������˼��Л�&�=e��@v.�<I�O�s�4!ԝ��/�2Qb��<ᮀ��p�(A ��a�+�BX�e�\�J���x�#m�=~~���[-u��8-�)v�ƙ�x��p��e+�ݞG�+m�j��L��O!�k�G+0[�����ٺ��� �EhiNf/�S�}���)�Ȱ�D�/��B~�u���z���P��qt�\
�-Qor��- a>B1+���Eho���ʐ���N0%��,��>ŞFF)�&Q4itH3���"DTS�D���lg;��<�c��_H6v@M��o��i���$���V��|R(;<�a|}̤{��@�a�i�м�|��e�Y�ݨ8zw�aY���|�<��c[5��uU;�q{M��)P���/S��_D���������V	'L{����`�AwZ{UVB+v�����Ht���\��������b�VV��B0[3r��� FƪH區�[i�%r�&�s���chZ��U!�D�s`_�@�a�b_>#�z��_>Z��Дr@�t�&{g�Z�Y phꨉ��������P)vn����{���$8oрXI��������:A�Hs�͍���p�D��������+��k�;��;5e��[���]
�3�;\b�C��ًϑqG�u���EU�L$z��9��z<�(6>�0�U��fo{#{":����B�y���Q�|����ιY_:�Z�{" G^�,��@����3N��tS
��C��V=*�	��׻��k�6�t������� ���W ��
]��x���ǀ��^�˒�ci#�1Xޅ	�Z�4�}�5�/ǃ���S�yb�W�M+y�	���<�e��	9��I�_�'��|k`�t��=~q�}C3�����J-qߒI��m	$`��l��ӥ`
J/���r�ǉi��ؾ�"ݞژ@��oڈ�A�7�{Y{�D<̷H�@P 1W��d�����'���;Oi߯O��!dƑ���?��C���?���m ��&���[�+E1qsp�I�p.�}�����R���$�8 ����6�ݽ�vL�9t��$͒w�D�vy�4�������!0��JQұq� Wg:���s�"U��{M`�(�z��`�[���F����7�ny{P�3�6DJδЇ�L�T^��a^���P*���Z_��y��w�nC��{���O��#��J�:�*h`�1���k��Ve:�t�
_W��lQb�t�������C9S��0�ăD�Vsk�BF�+0�ʯ+��u�m}۩�l�,�fYTG��< ��l>�U�^�ZD�����@sL��<���bs���`�Ή�ДT��@����v�5���<m>oE�z�ݧjM�c� �M���6�:�]�$������z*�6kbOq�n���³.^�P�E��-a
s�$3���#��*z�� }8�V���r��)���`��ͳ�qE^��xo;��k��h��F׏?�����3�?W�*\��aMq�p��Y1�L�(4��U��ӊ�m���Lgp�0��Z��z�rr)�"#7Ln��
�^5��iR��n� ��
�N���B�z-;>La��{p�3� ��I�я�)�iܙq��A�_e��A������^	�jWhCڞ�'��D2�Ρր��?��"����Ҧ�����&��gN��.�sb9�'_P�{�=���iQK8?�sA1��f�.	 QN(q�8�|���n@��7޺�c7�����C�k>��x	�7�ٝ�<�q� B������ו�C6dK���h���`�	Ҏ�&܅�l(g\��z�
��H+�J++��!�S��Q9�,�a��*�[fz�������{�7G��?WZ�|���]Ew�������'>������f�Rp��젠o����9�/�|�~ݫ�;�=Q���#��K�W�6ͧi7'�3��n��F9:0bv�AX�&��ˍz!KUN�v�K��4�?@�s�l�_>���B���LT�<C��h4_���4)������w_@B�BWc�Ӌ�[��4�t�m)vV����kY4I�T�~�f��P�Q�\���l
l.o��?D��:��1���⏳��j�֊ʼ` �ޤ��x�vq=4����9�$
h��<I�32=���zl���� ���!o˚(�1C��ٵ�|;��b`�Ěi�>�������HF����n��)�L��&�8��g��1�ϐXq! &����c���򗏸��e��^JX����G��2� �B����Ty��^�V(���;�p��p5S��&mry��
j��<��(V4���V8SR 	�r�� �W@P��=�s�sgZ��6;�t	�e(��F�e���J�Pr�^Y-�����х����u��*�{"Y�����&�,��?��䘔K�=�>�������`H��1�(Ƣ]�0Abї���|}R��`CE��堘������="LQVMVC.�v%�'A7��J(v[q�)H�ݪT;v�%�����x��v�,���˜"鉰B9g�tq闙$Q�Xo�򗐙�R��6Heo�]����3٧:M�j1�ؒpo*S�����}�����|�fѡ �8R�\%_�E�髪N6#�)<%��('u�{�z�c.�f�_��>����>�G_� �����w���*�r������д� L��t�oH㫖��ř�b[Nq��k˦�!b��`���
�K��lp���;�!h���R�w�IaU���t�6�I�}�%�q�n8$Yio�`06�',�]�ƏN�d��K�ɠ����m�<���Ԫ���)ʥ�ӈB��E��#�����L �ݩ�Y�q3��@��j����q(@����$9`�3���q�qy�{0|ܰ���,C�kI	P NK�Iё�N�M���V���A�t�P�*�v~%+nOt.�Fz����<��?M�Ґ�s{���������K��"�Yw.�Û˕R����������S:�����x�\�^Ow�#�^��_\���AY���[�^�#��l��#�d���z�n�����QF6{k,'��{�����N�ji�೤�n�>^_u�C �ܝ}��9g&��4q���ҍ��%}jF(Y��+&(���=����Ϭ����u��ܹ.�����~\���A��h�7���\ո\vW�)g.*���5�(	�T�Ǆ�UH�&)�y���[)Y!���a�vV5x`p<����V΍���^����F3��$�RL��uJ�"�v�QtKkk��H�C�V�}��_�V���v�s��PwsQz��.���E(��nIF�c����Ku����N��VEi~!l�����}�KFV��4�Ÿ	�f�30e��'~\D����*�ç����P��%_�y���ߝ��jv��њp�o3�	,���E���R�%v�6�����5 )�?zk�&��]\���<���M� ��
m[6�ɝ���q���l*�gZ�FR�@dm���x��i}���Cbw�Gs�;u�5,J=ֈ,6�U�ܣ}����%L���W���]�Gq��������R过���4v�[3��vҫ���aD��'Z���%=d2�#NU��3�<��({ʋ�I��HT)?bNQ�_
c��>���,�fY�)���Bp�
����=:�l�G�N0J|�&�b3ʞI>��Y��Ё+�MN.��ay�C�?�V�,�����ʔ���K����4�Jÿ@(g;I������Y_:ц�� 
���MI��/s-O6=��C)�(A}Ee��[ {���09vȈ��]�e�����)�r�v�3\��(�<p��Pj��y�G�
/��?��=>�N�I���.H��3�sw�_�$�z8M8 ��G	����j�����5�ʥ��x=��j��؛���*���+m�?c����<ÿ	��Jg"��XW�y]���1�r�b
׹�/��	��Na�K�Jʄ�Ū\����&mTӂ�k��?ԅ%��>����+q4Z3B�pMLL��<��3�ğ0J���
���n����h�V3P�i+����:�kA��ٯ�i*fg�Ng������n#�l����lè���0���립�˯�J��V�7�x��]�.%p���Nyg�{��ti�r,��=d���t����/������t���$��fHzZT2;�+ԹU��hG��-T�jL5m��[�@ae��Rp���l%^
�	�L�����bFP^Te�����q2��B` ���U��7t��.aO?�1�jNz��d�� �F�i �2- 1����RS�ܾz�����p,W3;y�3g�Ҝ�H
߷��_��V��S\Xp������CLA���1�B�Ϧ
�����N*��'����-f��L�� V�5Zc����������6��8hF�T��[�4�|E��㶥��u��LMǪ

�]6�4°�&7��h#��*�[��R��T�}��u�I��L.���RR�ΐ����D�ћDW�O�u}Y��P��@sz����!�����N�!I�/Kv�7c�Zs�������`���`�U6B��f��|�ܒ�.�ӕ����F���X�j1�Y�`�Q�A�����GZ��"G�r�!q����&_����'��:��/8�0 >y�4�I�2�������(���켖����}�~f��g�I��A�EŻ'pY��
�f+��ײ�х䁖ό���l��D��\��Cٓ��o'-�XB�q��k!��2���7���\F��L�����-�����Ɵ��}͹��u��Q���hs�j��
�J�IW�~y��m2:��B��gl!����ؓ��E_����3gx�pĚ�y�C�v���qA�{7�5t�n�,����2��w1n��3�UY-L�Q]�E:�db�C~��2����4�&Mh1C$�&�T@9#4�Ȑ�~��o�����ѐ �b|%������+
a7����V,��RUM1JC"��%O5Oh�JN�D�/8#V��.g�3Y�3�>��W<`�:o:Rը)9�OSLhB��H+�,���[<�Y����z蝒���)��K.�2�Ћc�1�l��$eC�3=kT�@$��9V	��2�5�{��x��M��j��0��@(��rilҥ�힁K�%�F�.;	G�}PP|�^"o���>dMˋ!�}x�58u��.PV�%$Ͻ�H;}		�<cch)�e�8�0�1����z�Υ�o�w����19�I�N;�#�3̺�Yڐ�uL��֯������:ས	ֆk{��W����8k���抅S��#�r�Xkx���0��.|J[a�V�&(���������7�h4�����T䌌�r?*��V�3'1M
vse훨�DdSۀ�~~����J�p�Z�[څ2���W|bp`vװ����9to�9ɽ�<�jQWT$�`k?���Fp��NStt��rS� ��Oe��d�T^�5�֦~���R���%)� ��bF��7�eMI~�(� �R��s��10:v��9���*�E�Uc�]�@��I��1BS�ހ������h5���F�=q@��v�L�d-8b�a�{怩r
j�\I6�يO´�p��Ƨ1qN�uw~,m����!Qr �Vh5���Wm�<P�r>qN��y� �U�	�
�7޺F~�Ei�Y���q}�E��}�*�*Aܐh�2�)����!ZU�Uץ�]b�K��s�WU'rX��<p������v����в��:pD�<,rH��̄�ϗ;O�R�k���;Y۠(�+ddX<[��"Wa5!(�EK�vr1>����x���v�����|7�0	*��F� �F�LŇ��o�g�6��O�.�j����<� .̰��q�v��Q�J P�7!H�Z��
��[�J��ZTߊ�q����3:^�ʭ0:�W��wh:P��;����de��L���-�\$����E�j��k$���R�?�d��TzB[�f��trb/�5�z_���)��f�
�d���c5d9I+j3O�.>�-��x/R�����R�N���[�n�6�7��,��&��y�/�k�d�z���@��D�m:u�3�}N����,���S����ӺG-s�u[�99	n+]�	&�T�~���6���ݙ�?ȍ��T4bwl�M����T���R(�l튻�Hi)�x�q�a��@pc淽\b���5QEjF��Ԡ&��ہ�@��� JY�*����`�ބ ����W|�r0xN4���،/TWo��c�#_�v��w���p.dw�E�Qa�(�#���E���m j���>7	��a��>���ٲ�a�_׸QH
`DC�$����eC�;�ぽ��	1�M¥�k�R�B� �TA�� �ƹ�$)������|;�� ��53���x�!C3؁E8�>�+��;ͻ�.����
�zk_�>iT!�"xjq%=��[�S�/ ���`׼�2$Zޜ6��p���w�a�d�oٲ�T�_o�KHR��FU�>��%�,Q~�R�S�Zڊ%N!N���<(M���5v��������gN��6���M y^�P�	AQ���z�|����W�_@_�v[�$��z���SX��$GSs;��B8y������w�h�P �xy��j�?�.^�lBg���o����Jwl��� 3]E��F�	�w�2�׏7U�&�<C�/09"�Ù��`/q��~Y0:8�b<��88�n�+9�F�n�&�"3��Si_B��Q���{1��p�N��4?4}J�f5����f4[Ǭn�o��#+��#XJ^r��7&�6�4x�������X#�f��k���\���ȅș��7�Y�g��ٵv��ތ�G������f^��y�Am?���~��9MM����MF��ȝ*��:]�P"��M&�䳯��������v�!�a�W�b��ge^���	�"&P?�sZ0N��w���n�	o����/�R��O�N��Ws��U��~40�I�Ņ��)���s��j�ev�������\�:���&Ƥ�\y�`���y[�0T��EWDر�l�5��#y���3�ږpmr��^2r����|�ׯ�8��#��ㇷ&_N��������naTe �wpnũ+a�<���ǉ�#q��}����Ax����iQq���.��zg�ǣ'�Z��ΘW��#�N`�Ԇ �v !��/�"PcǾ	xi��s�e�<[
�Z~��a�}��2?W��3{b�
'Ʉ��]J�0PB����w�)W>�t��V�4�Cî�B��.�-Ǌ�(IN��Z �Cb�����W�5�].���&X�[�@!��	��ݬ�+�w@a	t���Q@��n�hn�X�o8��ҽ�S����Wt.�,P�Ut5Qm�2��층�Î�]��2P����Ho�q=���u4>L@�`�tV�А��.��-����� ��{�Nz,��x�{�.���-����N+��hB�6N�1 j�ּ��ck�et��*�Pe��1�Je4^�,A���DXA��o����}�5�>���������v{X橏*�.��$J9���𑒬���B�l�x�G�L*�6�X����Kvi���.���5o�*%��� ����_8��i#�dQ�iTA��Ա���y�� ��Q0����ګROQd%kd8_��32(�׈S-��x+p�7aM�������iQ(rՄ�� �����抚ٿ�\�^9��c|�>�g/�Iy	z!��͸�F�{^���U�rS�d�/��y���]*���� L�$��A_ݿNp:��t�RJ���D�M�1T�>��7I�b�ET����j��	��R��-�T\o 6�e=��v�U��