��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�4V��yjHOS�;��3�4�y	A䛔��~�ٶ2V2� ��i�9e��O�|B ��莫��Ɗ߇�o��
��T�J���̃Z��*=��1 �f���-\��H�5g�\
�b����'���x���|��l�����Sd�0�q�G�&�;��.��0��c��{�V\#����/���9��Jݺ�Y5�U{BP��?_)
��I?�^t�b�F�"rW��h���U��$�*a��O��zX�;'L�t��ɂf�W)ׄ���t��n��6R	t�E�A�M Euٲy�d(ӈ�I�&�b�.I��2��$�����EG�0�50S1ٖ�I���6+��w�݆1��s��>�|c<�#+��fn�0!4�J���s�m������n��Yl���nb(�N\S���p
!#�.�|]RC�q�j�L���1ا�v,����P���[*&����^O��"z���9���ć�ť�^�FJ�AXh��Sy�(f�W��;o
���ā�R�ch��sƠ:��lg䝎��g��C�B^������Z�,ª>{�&��D�[g��1���"���o�PYF+
W�]�G�.�0[.��xǽ����!��g��d��X:���@���js3fX� �
}��h���!�F5s���d6 noX����� ��$9j���O��xW���5����I���b�z���d���y.��gײ�Ҿ�
ј�fN�mE��;)�#�7ؑc7����a����>y���"�D��7��J��z"ts���8T�{���'o�.t����  ��W���l���� �������!4�j�z�����H����6�^8D��	�d����;�_�K�4��گ��C�g8Лu΋���}���(ͻ�bJ��@��Pݍ-T#�1˦,�h*����Gq����=o/��2�q�{�,�L~ +J@`��;��)��g���ڷ����z���Z�LT����#F�Wz�e�IC�7\Oe�u&��R�&sb�ܞ�����&`��<�O=q�:1���:���R���yoĉw��ժ�a�	�ܚ��"�W�hk>)Oδ�(��s�p�ZxPc����{ ���N$�Uʮ�c�#j�-��4nqxj�b'��1�Z�j�$�xD����G��z�w�x˕��g��V�F���^�%WoP���O�Ć��k 0ѿ3ٱ�fW�7��Y�=�S(V-�U,�kF�Jq�V2Ҏ%�#w�;��z�d���<�2w���\PH���'p�u��}O��dY���#9�o�Y �T�.�7�*JûYB��΀��������X����d��X�ql^���82ߝ�"`�:K��I�SIaR�X�i�i6C��Ȱ�P�'����K���28����O�w�̄H�)D����j��H Aw�OɌ���v%�������W���ď��k'a�F���ƪv��t����q�eٹr�e�b\�wj| �k1u� �LV��'�-E��~3�kο��b��Wh�PkZ�&a��P���`GU~�j�$3t��n�/Z�?H�����;9�6.�lJ)BbP��v$l�����۷��r`���p>
o` ˆYƋ�a����{a���"��{l����iG_a�P�v<�9鮂����~/��Kݨ���t�Eleo}�+I6��[C�W�`6�BC��E!�ƒ�JCNddR�+�r|'NBB��-�e�g���!Y�گ���A=��[?NA�| ���*S�f>�P��{cc�~���f a�3�?{��6��j���H�%j�a^i��B�=����c<ʸ��:��F�g\��<�˗�H���fZ0�g��U�A7�#2W�`�[j�3i�VƂ������x�̗��'eb{�m�)�jS������n�<��.�j�g��w}��^��>�D.��3�K�&���O�ɋ��$5��?�p���{^�e7����P�r]@��*���v��[��W��b4W�	��J�.Ev��v��/ork��Pm��^ ���Z{���G>!鮙�Lؔ�P���s�1��.�TD��b�iTI�o���1BB��K00k**�a�ߌ�e��-����-j�v�� ���k�J�&3�W:#��@h8B����X'�t��k� ��:Vx�����K�e7��.T���$����t&����B�cP��������� c-�V<"�I�X���#`�X��l�f_T��#�P�i�}��A	2��xV�K�	����9�=qJ[�r, #���[��v ƀy�]Y=��L��ۀ���2��P-�<�jSA���78y"��\�Ra���p����؜c�ܬU���M�j�߾�O�5����I�U5A�7><�^�5��C9y�kM�O��iE������p�)�VN��̩���%c\��V��by���čԺsLO�6P�����H�3=�L��Z���C�|�z�t�8JP��·��`z�O��.�0t/T�4�YTQ&Bo���
�-E�:?��{�`�b�@�qܱRz BG]�n�u�D���%���`���?�p�T�t��8&� jiڪ4���y�9�~�}2¹/7-C`����)
���eT����/���,{9�H�J����ZY�ߚ:�H���4y7� V���zG�N#�E�	����#6�4����G�E����և��P����'��Y���m�T���xs��k�j0^&#H:BT5�+���8�]����D�6���-7qE�.�/FWZ��̽����L"�ŀOg)�v�R�����UP����@����$�Ɵ
A|��_��[$����)��	�q�����"rڂZ��d�3������KyOq�5�����9�{((w�� 	p��[�R�8ʾGS;�1����(�y��сib	�A�:|	U��F2�>�CՐۖ��������h� ]���UV�$t�p�2No�D��f���g�K��4��� Q��	阩}m$"��j�$�x]$��<��3q�#׷S#�%f����Dm^ql�����k(�^���B���j�ovg@�w��B�V=-T�v
c�Q�M���V�y�(T9�����(,רd𤎤����>�ǁ�H��"�I3q;���{HH�ٹ�J@�Sd����4���~��ܷ�. �4�A3<�������K�=P26';S�$�a&B��G�u��ՍH�Z�6Vq`��3�f�2�W赞���(���?���IO^ �g�!�s�e��q�+{���K0þ]�E$V���5�o���MYp�'v&qj�)Ԡ�𬧉l<F�i�N��L?(������TY�ʔނ���x��O	��vd�*P�4l�jӰכ7�B26��nT�S��/a�L������t1&2&�W�bsY�dR��������Ro������~{~�q��@9��<	��$�r�n�����u�uI�NK��B�'�V�G%�Z�*��!֗1�Bc0mلϼ�A+,�B�e�RZ���mc�������r#��	+K)��r<BVhm[��:�Ӎ ܝ��$Ғk�"+��)6|�d*���J�S�|���{	*�a��>��UHL����Lp7�V�r06�r����kM6qw[�Pޒ��g"o������t?��"Ca�P��T�V�B	��
�LѦ������:��V{����E<�߷�EI�z�Uqv�~�w��K��ŵ���������N�:�~�c��<o�+��C=T���-����:F=w��Jׄ�/�xQ��Z��և�Y��I]k��{ �4��v*RKnB%,�'�d�=�Wm&����B�288nv��͜-.��)qF�ޚ��T/ R����	�$�`=�6"� 詮Ѱ���с�T �њ2J�-c��p�A	H2��?�K9�;��T��Yf,w�T�z���sY�[9������T1{9���l��8�G_ֿԨ7�PJ<|���}a�]��g�.���M�������'�s�9����Ї[h�
�v7mz�S����Ђ	��/�>��k%�E4栙��\]��lP���["Ï?�,�Wʟ�||��⚄8��,$�M��@��N���উm��M܈��x���Qjˋӂe��@ G\����&>R,��b4��F��ʇ�K��cE�@dn<���&��4l��Y�a4�7���r1%�og੡��q5�������Wv�:�X�5Z��FA�����pY�Bf��ђMU用WT��"��2�����ɪ�{֨M�!�	Ě^.D�?}@�����6��%��r�aZ����b)�"`�TY��Pr};�H�~�������S�U�7���t��˖�E�۱U{����� !�u��AӜ���	��y=B]<ƈ�\_a�)�U=VA9=9B�����`�LTk�U�:�������Xp�
3���e>A�)zz��B���)-���.�RR�S�q���v�I����kT����sMȘE9����>t�]��m��y����r�D7ۃ�-��i��lc,��S9�������V��C�S)��l�un����}8v����S�q�0��ʉ.�5�It��Y�8�U��b��!Q��n'I�N�X�Ebb��{{�W/�y���i�g���A0g����(I��]��~���#s;T��bBؖ ީ�J�O��u>�;
ri���2q���&�ߓo�&g�;ۇW��2�RQ ���y_��	$6���mq��o���t��N�S�G;@��ϐ����,*�&U_��4?���%���d5S$֘:�+z0_p6QG�' ��Rs�`��SH����2�UR��!z�4��Km�@���D�9b!��p�i�*��A`Ɇ�<��_84��R#Nb�9�o/�j����]�U�5��7�Q�ҕ�����G�|7H8a��l-��0b*"����	�����럦���yD7�-4�2|�<S�7��r'���� '~}�A�bzP��<�?�^�L�&�$ :���.e�{Ђ�_��u�}�+=�(jn�ϑ��ڲ�AN۩�Ҥ�����M�A���,�4T_U���t��}��'�h��]FD�?�	�D�DXiYL9�E��.�d)&��ښ�����l��UQ�����|��9�*-Љ�L2.��$P�6c�?�[ 2׃�b�㱄�����6�y٤tpco�:Dh���$��-��[ڸ<j?do�@�/TT%��\�m�����K���j����_Tt���FAw�N��L�G�@�?zi;��M�v ��1(�ҥHQj�X�F��^t�,��+-�I��^v���믁�/��L�>��u�DqUn߻g�Pd*���g������ݻ�
�RD{���/�8���p�<�T�2�댈l�0lE�ďWҩ�5�-(aX/��2B��y�����Nʛ9Iv?<\�??/W�$hT�� ���6���]sp�e|�i�g:�;HF���h�C̔�Ba��iz�'���HJ�x�|����*�@~�H˖�~�C�1s+V~�c"�5V�$#�~�RN��d��T�O�VF�Hn%{�$�/Q��	�ɫ��y�iF��;��+Oe��-B�������7��"�az�6be���M�n���a����i�����������^"�`��V���8��֚W>���9�

���j{G�JN��\�I#1o��}F����%����k����ـmG�)�L��A��ڴ3�,|O��'�����V?�i縱��-?瘭��4ȭ����P�c�F3I���� 8k�<�A��1�7�+�n���)m���T��S�.$���M�9t��N?�y�yo\K�u�<2R,�N��Q��F���k��9��3<'}}/��)����&ޣ�R�d� �
<�E���,�����qN��KL�����ю���"W�d";�I�:-�H�[��j�h�w���=�5 �Ϩ<�	�J��'����~jx9ӻ���CՁ̧@��o��9Ȗ�ﷷ��!i30W�C�0��vĺ��B{��I��)�x}�]���������J'�d:,�e�`���P��1�*}No��aDl^��L)�l+��a��_�*�q���xN2I�텿1)޻�i���'X.�_W��v7]=�6��Hygեd䫑�S��03hg�rbL9Q���@�1w��g��7N����]JW�`�Ƒ��!20:9Gi�*U58��\Iջt��q1)ֻ�>#]������ܡ�HlB�SS�_&6���C7�Yp�o�s�V���4��J
��MX�8O戦��!�}�&�?�.��	�_���0bx�<���f8��kY�/L��0���p�_���E�<B�m��F���{�-�Й��/�f��!5z��Eo��R�cպ���$Px\O-dm����|?{�����h^�~|�w�Ǔ� ՙ&�_9��Z�gxj�d��+���*�� uĴ�pk&��Oޙ3�w�U���s�2~�?�%h��)�`<.pil+X}�W�
-ϸ�ii_�=�^�%r�	T,�;�r�j�Vk����4_3��~�^O�px��xa�#����,у���q��4WG�KV3i�j������� �W��MR���xί>��:��/�w�t���	C��R'�03�(�����H�e@�иC�:�!;Mܡ�w��/ѱa��C�e��@Zk!��J�,�hg�<䶦�vp�8i$<<iH����P�;V��h�g��.�iꊟpz�_�^���s,�_�
�؝�+K���������Ķh�;p~﫮�Q����:M���i;$V,�6�?��[�l��o������M��䯢�4��i��Ӥ|:ЩΔ�?jk�A��::�xklm�}y����8�H6��h��j�<4(Z���fh�7b�{�xN�k4�m�#iƐDYZ�=�d(��Z�mKq~�O�-iTELF�<3m
�ӹ&��ĂQ�5��z~�O��+DP�+ўX�U��[��Ε�?(DS��
��_ ���O��u��N�˹�Ы���ӹ���8�M)G�`����2�Il���5.��+��gW@�NИW?0B4
�TkWI(��q�&S�i������[��d���C����[rR��"�nο���PN��@�����t/~��Hs<%o+ӅW�Yk�-���:J��O8�v��9�r�ƭ�Pz1B�'�<��]�8���Z���� \/	�z�>j��\r-,\�>�RHv�����xm�3p���I��LFPFߧI8�T��d,������4��Y��5"����{nA���C�j�]�Bt	|ȳJx�J@A��p�C��n�2����^*}ў|�Ҳ��k����vןh��mz�j^�ß%B�h	�e�l�����5>��!�[y خG\!5�Dm��"�қra��̝���k�ĉ�w���E=�8X��g.de�Z�>�S�1Ñ ��xB�HT�4WKe`SȧI�$=�q��Uq� ��i����ܠIs���Dw�.�W�N�lW͞�<�3�v&����C�/JvP>��EՂ�P>V��ԣ_�2����2�4��L��@�^����i���^���>�;���f�����j\��Ă��
7ߩ	y��FjK�K"����v����e�_��v��������>^YY�� f���'��ݚ�[(���(%G����Ȕ���p��S��ܱ�ٶ,X��CV������DO�_#ǺĚ-�r���ŋ_8l�3�Gl�&x�!(������V��&�~M�O������s�n�����r	`�%nSY~�.V�$(����v$7ԑ���k1���J���f��n��N�܆��<���f�ş���'4��H��$S���q�O��3F�v�d�������M�u�sd�g�UPt���{�Iɡ뫂��c���ʘ�:C
9��X�)�*�.�	�eO����I9�Z#�AWԼ�K^��B&�a�����M���!gq����ݫ����!���!t��j�x
���YA�!Wj�2���Ftv���_��k=�hvRm�d�\&���ٖ���5���0a�}hV�3W���S,u~�E�)Nj(H=$��	e�ȷ��GjuS�2kP!:�}����`�VE�]�6�A�֛�N��yk���eù=_C
�Ka����c�1�����Rh�ks�����ȉ��ЫeC���9���	In�NNq�ΐ/H_�n��h0�	*q��*�?�KX�YV����A��4�ޑ��4��A��S�^f���9� ����Ϡ�֟j_�Ko!��厄ȉ���k]���	L�[G{����qƔҋ̛��D�JG��x�Ad��4�!~��!�T�jTF�"Fi�h|9��&2��rO��Z;I �Ē�^�Y�P!��p��� �X�.5�n���t X�0���81>�֍�3�i&������eF���@�MNpz��2�u�U�`mM�u���~KH;�IND��]�Z |�Q�N���>=���9l�t�#����b�m�'���g#��B�ɍ�PH�<�@>DHp��������2�ÈtN���YK���>䐻h��Ͽ�M��h��CC�9("P9�`<z%�_�)�e-0�i�RԄ����[=��g<E���rn���*����}h9r�ڐN��!�� KV�Yp�:�WS��Sd�<ib2L�r�D�� Kz�S5b;/!�I�׽�E���潇��9��g(�m;NVΗ�B&W8k�Ro헇r��Jg�z�Q�kp������������h"ӼJ}�bk���%e8gYlD��W�~�$xZ.���5\���dN��۾N�,��)c�{�.5�#���A�Z!@��E�Z�?��Ց9�
;%�z�7��4��Nb�l�� ��2��h���E��ԧ_�'��q�*��.v��!�p�Wfw���;�p�m",�"�*$n��{ �-�S�j����_e���C»�����(X#t��d�ƈ@ض/?⺠��6!
u�J�Ĥ��{A�G�C�H����jjx��X�O<��W6V����!@�z�Ik�M#��*gN�ZIx���	q{�)�,�&��m��3���sOJ&�텦��4���4=�ףt}�e�[?�5���*F8E��m���_ѢZ�kUx`�C�J`�p �vj2���u,��
�����Vi/�H��[��4JL�gC�v'fP�j� �2q���WYŇQ�sMɳ���X�+�z^`�R|�C���������@Zyp䑆YZ�Y���u��Mvzҹ8�X��o��i]��j'(*��!��q��~&�cG:�?���1f�t�/�2 ���� ��q���FRh�}^�C	_�ha
��i��-�
����VWds��r@�j�x9���n�-�u�&�1�� 4t*3�Zp�����3=Q�����s�eq+����Qe���K̤����B��r;�]�����|4zj����3��^���j��!FnppH	8��Ζ��:4�w|xv���O�C[�IY[�Cs�"��$�qa��{��[0$!�B%1�O�&`���H܂��hܧ��<&�8e�����EA�҇[�`�E�]� Q����c|6/5{ �q��&��qc`���A�@R6�?����Z���ҙ�[���L%���"��-��	��iǮ>.�g�1p���WB̨y�;d[�=Yӎ��^���"+Ґپ}�K�ֹz2�f��z��^3�S�){ kfD6䓣�qf��/}�+�p����v����Μ�%�U�֞xeN>�Yw~�6Sd{H�@�k42J��I3�L�������	��{�"��Tۭ�nʵѩ&F������f	As��
G��3@�,FI�.����Y(^:�$*�b�]���D�I$!N��@<��Hp#�t��A�`wۋ���n���w�>�"`8ojp�Ğ*^�L�n[;�Df�`aN�r�X��M����'!��LB^YK�|F���W�RL�Q�I单K�����$��㊟��?��a����J�D=z��難��'�8>�X������B����q;ʾ����]�_���q?��	�3�D5�_�$�x�}ZO��>�r�i�g5u��:(<� �T.u�E���䜕����q�~��6���o&+E{���������)��b�o}tA����2`sZ+�+�b�n��7�G<\�^k���k��R	�		ׇ�53R������wRE�(Bه��O�%K���<@j$[	#���{J�&H��~��1�g3��#�PV���9J:�?ǩ��������R�[U;��Tn�>m9���|x��Z�D�8y��#�$aS%�^}�8�єZP)3��1��E�*bI�#�\�B�#�G@8�����A��lOv��}ͳ�� �q�1�L�X��������|���g*�c�o��4,�m~�:�T����l�x1�q`�(�s�;�L��q^3�B�&$�o�^v�ۓ7��#I�z}|�U�x�YN�szk�z�e�t-S�K���Nϯ*��M0:M�����И���[�{7 �#��;4f���qk���ys�mti�+F������+A�[T��;^�RY���é�ȯ����U���_�c�D���<�c=8�mӣހ�g�J����IX�50e�
�_�I��g��c�s~� dYV�g/�X�IzC���y]>Y0�a��%;\��E�,r��8���c�^�f`�� �`�+�>/���(�����d���PA���-���_�00î�e7!�X�e����`����u�+�J�!�ii�tR�=�x�Ed7H��J��BgP(���w�I���j7LYػe�˨����ĝ�a�y�!�/ףJܩO��l/��)rWǗ+v©u���f�c��Ƕ����_U}�9�<`�݂׻��;��n� ��H\��.#�~D3^�w�*Z��<b+E�Hb�w�g�bp���s1{���t`�	����M�7��	�_Lɟ�ﭠ����P~��4V���o��Jٰ{�ʃ^� 16��4�9KP����	�_�D��2M2�B֏QZ�+3�����W6�>W�ķ�T�2J|Q"}b4�`_�jh{���q��x���!�wvj'p��좰�ŲL����%)�9������5�0���Vf|wɯ9��[�����Vw�4��� �ȃuu�k���
QG3�:kxh�W�ۢc��6�[ۅ~��/Zه���C�
�(�K�����\c�p�?�76~OЧ�i�(h�ޕL?z'R]}�_p�ѝ��1� b�̽a������=�!��R��Y؈�m݆=o��7�����};�MrA��Y�$:��F��չx��I�`��\���|P���6Lѕ�0�a�C�A�g6�j4�_Dԍ��ϥ	>�	��Ԡ��b�O�(!�z-ÛZ&�||Ep�9U�L��|�t\�S9y��	�-���V�9�w�wi#L��Y�w`��ˉ�M8�y�*��x_#{�AI���W��S���P`3�Ķem �o���bn����b��Bi��ބ���+?u�YS!g� �:�F*�$�n=��!�Ce��%h��\�w�Ɉ���+I�;�"��
gd��c�.���Hc�;ӆ'q�$^���i�Cs8��p�*s<[�(�eTԤ
S4`�{�似��`��.��)~2�f�ɇ%��AqV�?��d��Z�|�%�UXGX=_���6�"��*7�[�x*&�m]�҇e�lB����@:#���"��w��wq\=$V$iA�%�e��ݭ��ɾ���&�tޑLu����݇:N�WC��Ջ�W��f�[cW�
�4��.<6���3h�"��;h�ɠ���4#�8vu������UK����9ߚ���Rd��sԄӎVX�+���5E#����|��)F��:�$�2P��g��y��<CT���>�\	��s���Иߞ�I�a���,�N��m��؄fY�4�W�s���?ǁC|uUEk�˰��Zk9mX��1���Yy0���"���F¬	��?�u7�	�ǀk<\K�	��P{� ��'kb������۲�����o�P�4�X���J
�󔂐^8.����m��-���Y������qA
�g\�b��;7�
����+�g:n�)�rYց�
^��T�L@,��b;B�~>��}���l��[�YN�w�/������JT�b|�.����$w��#��.��_98��u�CZ�ݻ������y���"���m�����׃ 0�G��u{;��r���3f��5���y:c�컬
��}'�3S���J�k�Q���Vs���#��GRe��}(�UV�0�>�&�pBI�!J
�T��[󵦆G��EN(��䀓t�.;|;ߏ��^z9U~����9�Z'��@Y��E����v�6|�� ���|��)���%g�J�V��ܯ� �B:�*o�����D��MQZ��{�U-��nm|4�6� ����/Tfu��/�?����~�w!],�ɿ!ő��r��C�D(-�Y�]��	"��8�~�G��u� &�lNCc(���ڔ�T]4��Y\�Φ	\��?F�[�4*`f�8�lX�c�q���dD3�]}�mu�"����ɆY2 ���ʠ���En\�01��^�y����|f�Y�!�\1���A7gc��9���5\�v*�Δ�j���ϻ�e\_���u�+�ʢ�lY���P?��	ot��G��;�gqV�-{��M��>����nyO*X��u����'�!�T�=����g���+�/�q��z����^S���L�*,o��Ʒ.KX�R+��?�
�,D���9O��S� �U�еe��Z>��=x�8�Mt����	�����A
=�AA�7�yd�X[6����!��,!��B�F�Y�7�X(r�KJz�[��2hxzDc�ǈ�Η[?��~W�F#���������ʨ.h�o�1ցv�d����k�0:�Rl�Z%·�y����;��unm���ܸ�_�P����m�G(��V�ސ�5��iֱ�
)3�������$�āt�|�)�F+o�!��a�My�49�W��E�wE��1�]j2�
(�MkG�=. ��V�v�{�_w���ND ���yP��y���A�l�����d��g���z7���1"�4�2��'��Xb��b?Z�����J����@%L��c���,�\Y`��	�C��9<'��P��ؐ�ʵ<Y�M]��n�^�U������N���Đ�?(Ww�v�+�֐�'�mF�ˆ����#®����h�{�)�3���	�y�BD��-�Jb�i�;�㄁��L�ߌ��˔7Tw[�6�Ԝ��@m
�0�L��!V���U&���!�升�`Ӿ �P�O,0>��q.T2�lqW.񵮄���~c"�#�c�5�x��偘�|w0�2v18��#��z��"�Jf�?n��_�j<Y���>=�{{����_�΄9܆U35>�0�dj�,S��%��Da:���H��t|�_�}���.����JC��P�8^���n"I�����t��5l� ����#��好��+B�k3Gϣ�rb�h��C��}�]ґ��q�=��$������ň��r�r
P�h�D�#��\e{� �v�
�C���K(���k�y��~M_�Is���.zW���!J)]���y� i�ƍZ/%mU���.��]IygI�]��0��G}�z�6�uWYҍ�3�m�V\�OFMcM�����[w�9"�Xc�Cjs^v��󌒍�)�-��(�ِ�]���o�B{,��R�6�t�x����!_S;s�Q���L��j��1%���D���lC�(���� ��;�E�3"�P��L��։J\KTD]+����'���e^����� ����Q�����V�Yl���
ӱ�<a�b4�p��f�ֳ�<T�?rϛ�6Z'�rQ�YT��˟�v'Vb�V�%Y
�+�z��Ok��]���� ;,���'P�4!�֮u�qe���3ny�I���Qj6+�t&<���<����zX�4	��$L�s�Ws�}X�ax"�h�O�]p�JY侪4n`�>aAk�	/��*�+����J2s�P���bE�ϑQٖsg998�Be��Bi���X爥�j��R��o�q `�	��_�X���Iڂ'��Z���e������`�7b��9
���U�6��X��<N�&��}���&y�\��ѲB��~��]rr�˸�)l8q���0Q�9�浗͂ug��@�e/d�\�wt̝�x����)����w�	HR��X6B�g]`ë�!�� �ZS�R���.��N�H�,���8Z�Mq@;��EF`�b�im���ٽ���CH'4�z1�S�O�VV��b"�̃;{����8q��ͪHL�[��D���NՖy�NO����q�s�[|�[���Tc��%Q�Sކ�  ��n��:y8TT}��L$�G";������i ���/�U.� F��Bg���JP��)� T�y1h60�F5(��X�����YU>3��m�-���8�6u��uǋ�<F�m:�F]�ݫ���Nj2� E�s5B9Eq��d��w؆�_C�R�2�A�X8�ʂ�@,�g^��ʧA�0Gt�k��g#I!�U��r��ᔡ���Ҁ��lp)�	� �'�����,�'bHZ\����V���?���g�T�j��5pS���"�%=�X��/S��9�ݷ�5m���|0T�y
�F"�FK8a܏���"w��[�u�����K���1�6W�&0?|��p\�$�bJ@�d`��c4/���v&�pa��:�\<+���|Ǚ�V��9��U׵}"���@.[_�mMՂ �{�7�FU�~˕��}����ځ��~����t�r(Y�������� ����]D4��l���ǀI��h�IV�)s UH��N	2u ����66V#8�P��������>�xA��Y�uP�ȝ��2����/�	�j�"Y��W�$���k'��ѭA��wڲG��m����-������v�ǤU�K������G����������_� �u�>������#I�`{� ��[�WL��<U&���! d���(n�*]8#�_���.ju�}��@�;��vQj���P*o�V+��;WA]@�+�w**GzQRT�X�Y;c�a	s��D5�BYⱾAD-�Km>)"Oc��v�٘_�l*����D�k)�9�����d�Ca-����#p�~��'��n`�ˮ�zJ���7]��A+'��o��i�0Xt�d<�(��=z�1߷;�=���m��tLbM),aUT��#ȫb�*r��'	J�R7ZX��-��dg'$�=j5���_�q�Rd?�Nf�q�i�t���l���^��v�7x�BƠ�M�:�5Fy�I�T~d� ބd���d#�]��X�2c��=��^V��~HE�"��iq�f%J�*�	�?��l�ɣ�PXBg1�P�_�3�Й�#: 1T_pM��@����T�=h�Q�<(\B��Q6_5S��7N[#��x#1�V��Mբa*S1eYm1�ŽK�~�Mv�?�l���]�i�IG��w*���jm�_�����,��'�?i����۶�L1�#��$��ya�E�<o)�|v�+D����]C��2&Q�2�y�YJ��z�9,h�^ �����J�[d��S�������S��#���|ȱx�J�~V��RM���M.l��/W�0�-����ݔ���c�vE����-}E�X�.�F�E��N�n,GO}A9��'dQ·��i��qli*�4	��>��娅����hR��]b;��f�vTF������GYc��z��3�b�4RԮg.rX��,����o�3V� ��	ʡ,�p�_6�]���]�U�r}Ţ��>^z>+V._�&�y�_M���YV�g.�TiY*G|e�o�
�� fd��m�C�L�͵������=��rD��9�G�=௞�ǎ�W�y���_��jW�ΐ��̐��`��r���8���aĘ�x�
<��֩-������<T��6��}��nU'�����x�aF5��m'L�Y�F=j�}�M�I\���us����'N�B*��x\���M#,��v��N�K����a:L_]��0)��n% �w�g�IC;O �b'�	�����-'ls�q)�2J�Q}��`
>�BgIw���2�=/�\_���&�-#��Z��(݊p;:���.O�7z+�P}8�z�Z���?v��a ܺ���5�ܧ0��>���j�R&gbؤi�Q�����ҢΤ(���o��v���쓍���zJ�`����y�c��:��&)n�k�QH@�������Y#�u��"e(������9Ԟ�Oƶ�ު����O0�wlsbb�Si2�癬3�������E�%��!̲K�et��/*V1�D%��#��ⳏ$�x'd�j%?U飯e����1�A����)]a�<�GH�h�#㔝�F�L;��϶%��Cx�њ�:����\6O���y�֚3��N����)�������I,����?�ZM��1�)C�w�&�E�K̵[�Jd���@c�������+�������6<���w�l�����,����1]�56q#zj���#��1�T�nl]h�ƻV��Ţ("b�9����_��u�?]"�"�0���mz�W\ɻC]��O�ej���	1<u�#�#�`E�31�+v��x:�R�$�[4��3��b?]�՛p��L*�z�h��C30Uci�(c�[إ�{7�޿0��E�.��;`�'�jo~�V�\�*�#���5�ȫs�D �TO��Cn�����T��Aԛ�5-2�3Jc��3¸��@��M�8lU�eSv �Q4�l��:|�V�i��R
�:m�,E	�4����$XcR��.�oV��>����ձ��N@��8<�L ���SH�����I�!� ��iG�F�P��g�Qa�*��{e�Q�Q��������� ;����5�j0��T�AL��4X0���Iy���E��HL�AZ�<�N�f?t`���4lp|����JN/���#�����x#,L��=������Ż�g�OJ]�a���>��犿1��8��q��H�,lie_��Qz�y; 2~���tb)>�1g1� Ō����.Կ�����R�z��/sb'�,!/t�y
,8�&����)�!�ףk��� ���Rb�#�S������+V��KjLZ�� 	�juG����
��4�J�'��X��B�kGB�`�1&̏?U�R#����+%�9������� �����Z��c}ܐ����流�
e�+�=*n���D�ٝ��r"'�$�	�Qm��]9 tT��[w҉w��'�P�tr]m�D��M4[�@	]j���j�������Y8���:�ו�$���A�6�H��
N7'lb�ynx�G?��9(깊W��5�?��mj��uy?V��==�O#��+���Z�=�k�H�f�l���+f.2��ܤ���!t����r08����h�/�؋>����{��L�";?�U�&�.)vP�Iw��κ�N��&n(�e�&��Y7
'���G}&��*;<�)w�@L%YmK.�t��t���Ws�?��]�1�x��8x]�hĎ(��@�ҌO��J@:b��9&9���c��W�����\nޕ�����&�����#(��#����Y�$v+h�-�k��~x<�)�l*"b%SXT����嗘��e�˰����+o���./�.�8�l�ktN����~9��%�y��'�:��k��j�ĸ�
�&惶���Y�?�������}�I:2�fm�\3ofsxfoWE<I����x6Z�5��(�ő���>\�pD�����̝0�]w�!�_��I�q>6��ǟ^������Fݯ��&��IZӵ0wZ���N����v�Nd��A����\��8��vf�DIu�GeN� ٚYi��6�mc"1���k	󲷾�l�6�劫���o��.�{�`CT@�zݺ9�Щ$w��V��,9<��*?x-��:0６:�A��ٴc_�5Y�;���t7�����OtZF��td��[��H�֐Y��0@"�Cw%M;i�Gb�U{HI~���t�*+�s��Y��Ů�!O�@{�ȧ��� r��r����{�,G����(<�l��5�K	BY�|�O�Y6���i�Vu���W��̩E�T������!�n�iڛp�8�=2�}�*�pV*,@�,�Ӥ8<�>�dR���%�A��9�ы����u�β�c<�r�!�A�ݑ��,��͑U���O>�I��'�V���2�67�T�8`���pE=P�m��eh��G��ߌ��L�U�ӱ17��AFA䓥v����7]9�q%���aE6EL�ӵz��\ck�d�b�=l#�.��Mߝ#K�m�Ҝ��6�UF���� t�MR2��D ��"f`>���'��ʦ ��G�$%H�L]��Z<����G�-��V�_K}�&m�ꔞ�py=¥�à볯ꁭ5�Ҫ~��-���x�:JR���|,2.K/���u��������=�w�����b���]��Ĥ0Wu������ 4$���*{���M��<6�ְ�a_MaA��_*�:�߿HW�-�`�RS�1�T�|w~����h<ϵ����;@��~�B�S��*!J�	�:2��u� yQ[ A�@+P�P�����/}�25�?(H�}�w�)�����8�A�ztո�:��D\c���ӆ�냄�Oh��	��\۫�.�VH�&a��t�ւ�7�^��
��%$u5�����c���yL��+��{��ȡ,Vp
E:,}�j����X�&�8��h��ESU�� 0�7�;f:+JqÃc5�8�̫�R	^�#�q�$���u�]�3��R:%�����|-���j�J��s�ڑ��/O�$�/�GX�V
=�ne�\B��g
�^{ܦ��.�F�ؾnS��g zC��Zb��G��K�<q.򁋲����1��ػ7FwqvN.eDDFo{=m$��	����ђ>">WbE�B���Rf
q�O2�G����2���e��RO2Z�x���وUH��r>�8-��ȼ�@ιX���h#6@ހc�ژ��2+�ci���څO���9� 6������7u�p����吩�0r�I�$�{{�ۅ��c�1Y>i`䠅5 r��t(&Nj��5]��y��\ �'�����-&�N���fߚL�O|n��>����mq33-�M��I�8�H'f�ϫ�Y�%6M"1!�8� �.�G�Oa\G�B����r�Z��/4�n���s� �,J�3�D�@ (#/I����m�glbx7!-����r�KZ<캃���O�g=�5A� @�	��e&ƾ���L1��
& �sm���ނ�-��E���8[�NU�2�qhTs����G��C(7�b�u��oFB7���sUE���QY����z���^7r��#���Gp���n"5�;���U�v~0VZ�M�S�l^3�Ԍ���j��k�d:��P�ж�����r�+�8G缓�!�q�I�V:�)+$�ja���;���a�O�G9���JYC����׻�h4�,n9n�Y�7Xc˟�xQJsw��<xy�B��;7�+�"�d�E��/,$��uKj)i��|��;�[�q��i���?�I��w�q���U}����^�d:�����t�ߗ�o��b��i��ைfP;��j�!(%�2�$%������ٕ&[%#�I��K4i9#�g��tjm����9|��i*�j:8���bj;n�	)M��
u]1WL�J�"Z_��5 M%ʫ��M�"��5@6��Z �tC�����9���<���O�_�J_[0ui-�.?Ʉ��/�FD,<MIi���d�ۂf�����k�~��ϥ�,�cyjRk�r�Ӷ4���%�k{�����W{]�jMw��>���D�w��@���̣��(j�e��KA���H��O�2�z�l�����z~�3%��m�$���������E�v0n�:E�r���a�:��l������"��!�z�ān�e����ʎ8�vw[��{I��Aۯ������1����౽7���'�{�;��"<��!G���W[?q���������}V<#<S�ҹ��P��0k���ʥ,�[>yMz�[� �9)�F�����|��0SdX���Y899�%A�t��[���۽_��f%8�g>����u1�]��q2�V|6rA�DP�K����ܴo��}�����ډ�����\��V�{��
�;��DF�|cG1�b�W�UG ��gBq؊)%^�ѥ�nA+�����,�U��ƹ8
L�R��BD>!J�3�2��ZN��E?�R��~- ���/��s��k��&�k�m�>e.d��$B��M[��d��9��د�8��O���(DKv1C��Uw~g���;�Ǯ�lCy�j�H�_���Q�hK���E�JRfM�T�a"�Ǉ�k�_0f~ߤfe6��4�I�BJ+��l����^{��s������R��#)�����*'��Tf��ܔ7_��l���{��L��yn�����r�M)�?+����g*s��5�兢P�����"�R��}�7E(�C��/|����\5�zZgU#Ԙ�ÒG����,�Փ`5D���	�P��4~L�R�`C),\9I|T�IM�$�z\����l# �Iɱy!��^��s<�w�����b�3���f���u奁���5��g�%�F�(׀����I鱙��ZO=9�MG���JZ�Dvp	�t}��
�1V	O1� ����+��;����@�.�r �ͷ}�T�����a�{�u��|`(o_f��1���S�A���������u���n�5����Nk�G��f�+�ыFOQ���3��xƮYÍ�Qe\(Cv~���v'8�y�|$�=�1ΉI�W���S9��KJ�#�c���N�?�1�&<���Ȉ�S��Շ	����?*G�I���1�w=�2�����G~�I�������14�b�I@�yN	r<Z���AyA�IډlAڏ��< !��c���n�)M��l�8�A;�iF�"��Yؗ��)�H�c7Cڍq0���4*Z�>��t]h��@R�ͻ�{��iO1;�r�$#D��يo7	I�u�㧂�!'�����&"ɫ�O�7#�^(��\���t�-bۗ�C���J�x����т���g;��b��e;��q� �e���f"g݉�w*{k9W�?",��2��h.��3k��G��z���k��}kf,�ҡ�/���A��hg9D��U�ΪOH�l�00�|
`����(��&����2�>㔢�YT�V*dt�gc�#~�YV ���Q+Gx�SW��j������� ����#m�ĝH��������[@�@��!J$�����U��S ��++�UT`�T�|m E�(��Pr2vp�dJ���?>��.E�M�͒�&K�Ua�TN�^����]��!��Y�Aֿmo^�Ti�$�z���gzx�+&�t�$t�%�1Nk�4���R��Ω�������.݀зB��j |����ɖJ��ܑED�-3f�$�R���ނ��tKi���q�Ft�����0�Di���軹����u�tM����c)n����w�/��_�,We ����`hI#���T�. 8'�H�y[F����҈k_�޾��K�  wW���Ġ��^5#A�T��e��V�8ϖ�3S�czHw@9�~UW�917C��^Y�.r�[�ʐ,�^�� ��3ߝ���3��M�<�lg[�j�B̋���a�-r����H����%�6�n����EP��̲�+��}U�28�e�^;�k�������q洐�P�q�����\eKs7�B���vE��ޡP|���x��ѩ��� [�n����c �[s�ד��
����nb9�W�#�`��'�����_�����E�f[�4W�,`cD�9O�9��,z��\�͂')�cT� b�������3��M��Ayf,���Ia)9M8�	���G|��j��}�J���Z�3��� MT�ds�OJ� ����沮�<[�r�!��NH��������,W�l�w��V�.�Q#��;*pܯ�!v��B���0GdS=�b��6��1ɗ�c�6`�K���Zi�-{d�] P����p-8
���C������'߶5���HؿlEf�ێD[��>��A�N�廦0����B���߫e1�$ϔ��"V��t�L5*fG�Jd���p϶���M3I��)]����dhws��w4E_�3���f��c�`6�W��ӟ$�H��Ვ��T��}i�%��Ɋ�~=2��H{��9�u�h	|O,� %L���|�0Te�W0]�#��V粐�8��p��>�� �^!b��}I ��Һ�������$�<���̜��3}�qo<���IԶ�	��J �������C���-8�T4�����]�#��������<��ZE����p�r�]��#�[��; ���hG@oB	-?��JB]ςe�s�W�MqԌC5��/:,�P�n�=���ƭ��I�oP�Y��SH-ke��0]u�_�a4���n���"���ˊQ��q�,���D�^�V0����n�,�x�I
����D|e}�ڌ�O�E���o��"	����`�J����n(��x���П^�M����P�ȋU |�Ƨ@B�<7�Ư4P@� ��Ȯ��N�� /�V#�_��w�Ǒ��T��C X��k �4���7Acoyy�����r23FQ;�~�-�gE.���}6��]������$��'9�3�Ƴ����L���ik^cd'8��t�Y<M)�T���C�S�@�;}�� �8���m�{�[�jo��Ð����{�K�,�!�����y�J�A=�e���/<H�ٽY`z��X���p���m�ꙑ�'N�ꖱd���*�|�-&�#�p�<kj-��3��rfP��S��ʨj`填�1�6���q5����w���8ߓ�`Wـ��m�ÿ8v�{:1n�&��� ��B/g����0'_�D��)��QX�LO8��t.�s9-��ڊ��Y"�+��W_Ţ��P��Ԑ���P�x�iM� ׃8��>����U�P���Jh�W����a�P����#m�����MLa=u���_�=4����ѐ�T�/��-�j��C��K˟&)�͸��tU�I2r1���n�c�#[R`?������H����_�3b����������CSW��9:<V��ͱH�U�X8�[�mԩf���9Py�N?�\���.��l�PVw��?�m���R͑j�q�1�+���Y ӎ!�E?V);�t��A�5� �{=�A�$8����oI�d`��5��'}|I��g16�Ԕ�1��o߯�g���F4t���8�O!O���5�!vPu�z�}S�Jܾ�`R��'��.w�+!Vxژ4@�I�oE��/Ɵ�.�G����~𜛷��ؐᘤ�a����<�)[�'�2cX�=�h�ڛ�B�j�\�Yrn�W$q�����moG�%W�lu��g�U����*8l�̡4����:i^�O�p쪲;[�T��\�H�]��B�t��2���f଴8~��VNN)���iB*-�Q��5�3�~�)R�KX	�9H>�Rh��D*^�DcxXmL���VplK *'�2P���ܹϬ2�9`O��%\��7p<���q�m����|� W������@����������t1)�\���1v�!�tշ�9qI�~��8��zQ�]<�Z=R�7<|���	p�|�R,-0�������$&w��T |���)woؽ�T�7����1��0��۱�&eT^�Q%�y3%�2�]��&T�u5�֌|���4�e�Z?z��Y?��UЁ��d���򑊚{��d`��5��d�(�Y�����ڄ�W�$�Hoo�\3����J�>Ӏ>}զ���JK�4�����RhVT�w�vAqEv�FuV��v���	m�;���St��P��2���3r[]-�=?_D	���Ʊ��;>whc?�bG���}�	J-'����?&W��$���`��d�aiH��;B�fWC!1����q�D����Bӥ�|�=g��ܣ�Z�$���v�m��]��^���D�2�u�OV�.hp���<?\s j�`:���O���/���=�Tmg��G�ם��y:3�\x�b����=
��&�����C'�S�nz�d �I�A�������mz;�8�e}yggxYPz���s:�,�--���:ʧ:��9رx��צ�N�o�5��I��k����$Z8^SO��}��`��m~�#3&��^�e�o:�~ �/�Ud���`#��P�"_q�bx�����e:�K��e�y%�x�� �vÔ��[��R���m�}R�
�' 5vĘ�`���w CT�Ԃ��"�q�n>��`=���|�IG�ז�P��I�������߀(e�2��eSw� �J3g�"�
<C��YjHǎH
�fz𙗺(��9�GV1?��5���μL'��OoC���
�ג���3�]�;�r�&��	]������f4��
�[���D�h�	N.��q#������6_��A��Ot'����bvD^Ʊ�5�Uf��Lٟ�� �����{/Yen��Kn{-��l
Zҥ��U�̠�.O��.kl��W�t3is��Z�՗f�w��'fB3�J�[t��9g�;!���y�z�1�f='��l%5�i���G��C�����&x8G*�s�̌X��b�
���'y�����&��9��_��E�.�ϰ��,��&��/�
��dS��`��u;���p%>�Y�=�_�y�@�hU�i���N
|ar�I�dF�j����+���k}�|��1�7�(+�`�ɞ��g�8#7,t���2���!%8��^( �@��ri@w�VS�2�[���DM�u�������t�y;��H}�З�4]$�7~$��^������@\�M&ש�ΰU��&��s�!V�!4�V�gY�c�o��tn���+��. ��uh�<%��d��#1��Ǆ���ي-��H�X\;6_W�H�u�+a��MU|7���j��t�)X�edQc�3��^ �<�,�<%/�QN'���@�GY(R��W��W�g�nT�m����n�?�~*3
�io�x;<�3�������р'_6�&��l/��ޮ��w����)����u��:�iS	F��e�$6��!��My'�e'��#
��G�HxFI9�([,�،�0�hʻ�)<�[�k4������f���UǮr����Al)��E�e��L������#>R�K�L�cj����3�qMd4�h���V����6��O��f�ꩰ��m��g,16���i�S���gHôMGTZ��"j�����@_�����-ݹ�*���pO��U�!�2H"���J�l�^\X���d�a�c !��8�7��s�㫔7��x�;��Whk��+�e�1<)~%��Y��tf���g[v�G�z���ki��Ƿ��zz�+������d7��FS���,
Ёڨ* �
1QwKծ�l�>)��pI�*V2Gz/QX>g���:�GV���������s��ʍB�~���R|��\��V��u �L��|�]��R,W{�"����3_�Z�����a�%�5�+Cn��H���6Z	{D�:�#���Z`B}�"Y����2)�H�0��2�F����F{b	h�ץ��@@��F\fj�k��F��Q�n�����W�����Ε���e�}VT�
��s� ���Pb.�,g��n�3#���]����Hձ�\����.�B�`���J�h2�I���n�#�ȝ��:D�������3Ɔ2��j�xG[cQ_dڲ7���pu��Jo���4�O�����;���_e��*P��y���*ٖ���r_C��Ҟ��]��C!(O!E������t�L��:�D��*�Z����K@��$��]��*���u�w�\Hۉ��]�:����cۃd1q**(��Po�ߗ�@o�$Sd6��ژ8 �:v45D�h+j�����hGbW���U��p���m��x�Fj��� �|�wN�S�b�|�~ �~~�~ϼ�����	I�w���i��x��: ���O���^eREܡ5��D2����s�)�QoF��h�]��%ta0���O�{�����`�֪+7$/m�pЃ+o����(����6��u9�j��R]*B��s����{� B2��qy�~�ߗ�D��b㌞�Aa�M���S���~i��t��߇(Ͼi�rҘ!hP-]c�ꬆ]|J��[ �|�]gm/:��R+�B>����7Y?�v>�� Ƞ��X4�xF���N�|˘?(��1����ԟ��)��F�L�sP�ޑ�� =����.�L���3�<�~��KR!��W��O15�еaK��0B�y�'�N WH �V��e��O�Tx	' ����ĩ"���пVxbY��Z�ώ��.	xq����o�ZC"[Lr�=��ߜHYeB䆣G�x��_�=ZC<�j$� �i_Dv!�M���x�b��.f$�SK�7>0s��
���� �p9Z�2cJ�:�$E���w68���γw����aH��ML�Cvr&�AV=o��Ld;2��
XH��c?�fc��}�����(d�V�����<{:~����Җ;���/�+VA��h�,��K����ZrxxFH�:�C��Y5l����/��<k��:#�+��.lX�@�S�6���tՄ���L�]�]�q'3��39�k#Zv[����wP�����m��DBʭ؉�B�l�D9ͫ��=Ц^����V�0� �f����E`
�\�-�I�����W�,�A��������8�/Ҵ�6vW}{Ie�#yFi�$u�R��$��>�e~�6���rU0�N��� _6�
��tu7���l��!����`x"̴;�����e]ē�#�s�V��p&��`�A2�m/J%�������¸䄒
a�^9�W�7��)���I�S�w���V5DTOw��"�����p@��z���|W����$xx4���23o/!���_vw�<6^�p>8W�4�A#�M�A�rRc�BZ*�m��#�d-p�/���栠/~�+�@���Q=,9AW�]����z�E��}��b�H϶�~G%w���%�Y?S��`�V1�d|�h�j©��z��o�ߍCԵ��K^%aZ���y�@���������c��hcv����XAd��s��sn����@��U�QIB,t�@�He�*�´�}��䣸�y�pׄI#wD {�*�e댩{��m?<B�)څ��uQki���-��!P9c���Oq}L�bwv�~�\�b�e!�;���P{D�*𻷎L|8�����7V\z���PE���oV�2$K��w�P����%nC��4�U旡��肅e(�����Ap�Jܨ��XG�r��xșXڐ�*������80�K1�@8�XʘᬠT�ί_;`fa�ۑ���!~t^�Nb�	�W���8��)'���'��:�x�Ih�9��q2�ᄞ��ĨLY���T�noN-��7oi�l�wIKY��y
�k�5f���������JS	m������K����Z@.�`({��dLU��F����H-;����uU\%������=���*�1�]Fe��7jxT���.NW��J��>˪8����֙�Up��*��<#p��#k���qj0`�h?l�*P5 _����ʸ� :����JJ���q��nˤU��c������6����㨲8�'рY5�c^�� �I1I&M`h�Ǭ{O��ۇ�@S}z��qm��%�,��S/�5�za��L��'A+���a��J�@��N�I	�����NӼ���^��tp;�Ј�*l�J7�}wl�6�����G�+v��2�,��=���v`twF��VrguS¿|��^�+��y�U����u'�#��	rCa�>L ��
�J�����yqF��I"=(�w�(�>��͝��i�o�2s-���=J=�]�gx{�T��|�T����!�:��`3Qg���G�����Z���x��{���������}ߨ>����E1u]����������ř%�� <�5��m}�W���~�d�?�=���U�����,@�̱��D@��^c�aRJ��*0���au���dY�Pӳ��`�\X��u�h��]jmK2tY	lo�Ƨ%�O�D<�a-��Bf	v����~���}9
�率�e���g{��x�<��[3�\����cS�8Y\��K�%���3��V�Pv�^��e�����_|���Ulb�X �$�@H��-7)S(���B�2�X�B�v���	���>b������H����"���@1�|6��rʔ�Ȉ�&�b��.-�k�{_^��Q�/ 5�zR�Y��A(�g$R��P7�Hj")?ar�jf ��M������Vk��`9ŭ�F��-+�G|J�0���|v6��mT�#�kuK�2E�{�aJ�p���'�O^,(K���$?m#�}��f.6��?�6מ�!�t (�Zz)�%Aq6���'Rɵ8t����i|V1^�~�2� 沚��^\�A#TA�|윱#�����v���K�V��:����	�1S!fH�^���UM۲҄(�:��N
Rh�@�V9�b��0��p�G4y:��N���`�l (�f��/��.��x���o2I
���b-�AnrT5�<<PfA*��O��hPN���G��E�$����c�4�9$��
��(��g�&�<�[�PO�X��������S=�K�^ñxb2^G����ɉ����|��Uf�̟*Cd��Y[���v0�lw|�&|9B�`vW��a{<��TO�4[ '����=�އ�Fh����\�M�����.�}�h�Ӹ�0P�c��2�"Dg�4B_�:���Ʋ�b�*C��M�5k�)�1:�[��u���yq$I�4�M�����y��\��˨���	(���ӥ��(��p��3��i��˭@2"*<�Z�᩠K+Ӓ��,�42��:\\��s�A �Ht�a����sP�I�F� �;4x�*�:�����c�D؀Fs�}�����k�����P֛꾡)���Ǹ�̢Q�����T�IPT����fR�s,��>�MЏp;�%.' �K�XH2T7{�D�p*��i�%�̇��5��� ��5�����!뤟z���87��}�άg�p3����3j�{x��ķ���W�~� �	s�vӒ\P36�i>̞,8J{��I�o�i.�F��J�	͠H1XVFϲ��g�.�'���S��TX�2���OM��n�j�{Io��Ə�:�%��O׳	�ij�V���:\�_��2@>bk�L2���A�TO�1~�	���i�Pч١����gc��f|�%����ռ�e��� ��Ujk湚
�<�3����_ܔ�JxS��/>����7͡+e��\��+[-P�����}�[5�攓R�9�j��w8�;��⡬��L�1��4��ҏ���;R�a3�R����,�/
����!͑��?��W�%�-���:gl!�ب ���j%�n����Ξ"]�e �3�.�_ءo�dW�գ1��՝���oPyX��y�������s�O-���_�l�������M��m)b���L�����{;4s�����d���Ź;&��"q�l� ��P����A�]�~�Ɂ���[J2�ަ.��ns{%5��V���)�č��0
�$O-*f���/�����H��
���Jl��ؖ�T4�������BD�ǌ�*}}���DU�(�U��!�Y6�i�kb�el��|�ٌ����a�%Jl�>鱣݄��.p����"1M!>�};� DqLC�	��a�`b��X�1���"z�ČJK�:oz0�0�pCK���1z8��ߛ]�oSЁ�;����Q;��� S���h��j[�>��!5����`��%�-�e(a&*���Mq���.�F�!ʹf)o�_���Zs$�g��bD9�X�Wq��3�O�0�4�n]��o���+4�e<��W10��V����RJTp�HL�R���%y3�רg���Y�ٽ��cdw��嘴��Q�����6��?��H��(AP��7hhQ�(�L�

"���� W���(�t{�VI��_J*c _���Na
����^b�3�5��ǒ��p{��vp�� �EO�)�����A�y�*1V�����/b��+��Z��8�
����s�[���|d8!Wn)n��r�����(('��c8`}�v�O{�sh�]�g�V�,�7�J�eٌ(�A���6�w�%����J�d*Z����&�)_�r�`�0V�͘c�vȁ��6�V1�4q"ߢ�0�!D�`�f{��1�&�	�QO�#n��'<�6R�O�vUz��Q�*�GP0��ЋD� /�C��)��i:c5�`|���Q�Tڗ��%)���E��p��|���2�a	V��1Y"*�J�\nB���,�>�m�&��r�r	yj�k�ڕ�:z����L|�}�}X�����6kd����a�#�(�+*��n�n(F�-[I/�S
`1D��ѧ{RX�]]]ٗ���{D��2�#8µ����Wz�lz순Q�a!�W�g9n"�~<����3�9���Ix  qXM �(������q1�����v�Y�+/m�̫hGa��`4�
/Z�S.Tpp�Q�:��^��n��.bb��.��1�L �.i����X�!�,�$#��!)/�໩
pJ�Y�K�j`y�w�� �2��0�*� T�j	T�q��Wj
��c[�N���=j�dݸj�Ix"�r'�������ͷ��ӣؖyب���@�؎
���l�6��/xb;}�F���R	J�8��g�kH�}|���o��$�ʾ,�+���2:�e1:�e5؅���^S>��L˵V�m�H�H��K����:� �f?�h�}��x��6�8/� H�dqڴ�g���T���N��@I�2f��Y�`"�'-Eu��dI#.i�4p��{Dx;'�Lv��H]BR�|�ɳ�!Ɨ*�HHݭ�[���$�}�`��- Mѥ[|�#�ȍ0�����T�V7?s&�s���ΠL8�y��p�Ŗe7�r�DD�V����,��|�����^���j�m���3	���V&&L����&����Q��!lM�%{����.Q0Gm`(�ǳ�+�36񼴃�
�7-d��ɻ�����1�m���Ԩ�ʨ��*&�����#5;�:��B�)�F ��f}��7�a�o�aeGKpD+h��9`๦�	2�L�ـ-TL�<T.��?m�*�wL����^�juB�w��9�lE��wϺ�𦃟p�X�iv��.�<�qO[�r�Z�y&ǌv���w���B>g�<P`6B|�Dtm�"�SiT��
�����`�mq�g�Cd����1��4�<Fby�`�X�r�G��,�>}�C0��Z������)c}Z�#�9�Q����<�#s;���	�eT�R��a�Qq��T5��'�.?	�a+�ь�������^�:���Ǔ����K���zR��cD�V�V�ec]���Yr�'�7��@9�W.�Y� �7���(e�f�5���<#	Њ����ȗs��CT��u��`�������֪�~�N����(�B��b����:�d��d؇[�r�ͫ��Dϗ�#��8��ӌ�@v��`��x+8`%��(7%�D����}��:\�fwʒe�*�|e�ؔ8¬�����U
�h����#����D*o�V���21`λ�m�Å�������9ѼbvL��:����]��P �˂�:�9�!��ǽ�`�<:l.�+<!М����!ɪ�\�@���8����M#���JR{�۴��?�ǿm�x�"��kM�����v)z^d�d�n6��+�޸���KOV�%m;�Q��o�8��A%j�3�@��[Z�`%ٔ<NfD�Ɇ�l��9,�����{�8<]ׁ�c
�����ݘy����lKnB�{� �3����FMDr�5j�t�����
\��;+���;i���D$�ፃ�����y3���8��{�?���R�U>�]7�ge�Gx�����1¬��O^�$�Z���?c!���:sE�I��N]&&!CJ-
��k�}���a9�t�S�Z��K$4�C�L4�[|c�b�t"����XZ�ُ֨;�ϟ�\���G��IP>B_8.�fw�6o	��`;�aT�U�'8P#���(�44�V��/��W��vxC�_�v]6T��_��7��r͌ 6T�v9��5k�u�Aq�0��P(褌�pY�c�>� �7�A~��e��A��O�#�i�<��s�:,��H�a��;�w���ME����WQ-���c��;.���K�d���mkFF�F �
5���C�.����u��U�qם�u��V��}o����-�]-0�}������Y�@�~Y�B�k��Rw�����Q�!�,8�ɶ7�@�"�*����+�ԁ��6�>�$�s�Mп���Z�)S��zp�mI��m�����A2#I�4�2�R���J���:�e��͂xQ�Ϻ(���\\�\�fjs�f`s_�vx{������m���#ì
����D6ޠ�[;��+�J��>Ԟ󔾬?�hX�Zlɠ�enc�I��O�"Lǋ��1+��\(E|����ɵk��e���>�� n�G}؜�6��?��?��b�֪��0k�❢@�2�iq;�q����+ի!���Ӳ�L�1����ʝ�S�p	