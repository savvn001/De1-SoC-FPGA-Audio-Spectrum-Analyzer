-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TZF3jEaLQzq8sQZBqQzdZnmldHmTilI+pCOVTZQFOCljHSSJlNkY458vDgMUDyYXxtYA8UeARAo1
aYqf++h5REDH9zQcnHo/BVfsth4dpMK5rIw58YbKZ18q1ZrJ13GX3M7SS/OK+ppdqmpkIGwSV4GC
QnppVQMEu9CeV13Tci6s7I8l3zQg1aMd+gFE9embVbgz1QIBTI+Mc+6fM/djDCIc+QBf4t5nwOMz
3/nmO1AvRdP8aQtAW98US27l7Y3dMAm9EPCldFAZ2/V/gznmbb8SyxJ5/FOlFzMRVRIwbweYHn7x
jQxxcO2iBxXIg2xaWhnN/ZkGfswaunEik1qGXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
IVOC2EtiYM1oie8LKg2Gipdye2asWblf9Szq9ubN60jYxZwlrr6yoGxWZW6ptBSa9BO8QTAEyKe5
+ZPpsvoCOe+ob7ugq6SV8MX75jPd8Gro60gkUfBX+KU0BJ7jQZrj+025x6v0s2ho56NKNUrUT9Al
VwZdW1KAJCRQ9/Nfphpc9yP5NWoj7ria9wRS6j7K9R1LnfGmZr0OF+7NKoOfsevRBD8HWGyXPjeI
Y8FWDXVXtVPSxfyzpwqOeLVMXXvXqPSGNp/Sj35rFCVYidESKhk9LwaEHV1z2Vu/5zjpnQFM3uY6
3YwgaSbWZ9KXlZ7MTVUPH03Vnd7+Fzzu5MqZ638Tk5Z0mlgsvMoO7x+9R48vS76+2QGTbLEGG5VB
liKsDSdziY/FplC5030axWsiyteWZLNoh2mRYzw9suYzPRfM8XSGxfOGjetCn3srbZE1EagoSqtN
AzMoYVEsupz0uDewsNUtFFTve/fkic9D3ZBJXmE2jXcB8VkNbcTjgg2VWoFowuqaXGPJyxhRpFCi
UzbFHFtD4F5OaHedLCesUeub+aJMiFq4LiUt+/z7FTpPMcO0L5fE7hWH4uRbNcLOhnGBnu/ol76d
aHx6SFWUBc/WuaH3S1wbLL3Nwwq1Vrr/HEdygdwRi+HnHtXzCWERKJbbDHHLPhfezMq29eHaxlz3
a2IQyUkvlRauHIpJ2i6m/z97FPK0LjiQDVxxvCdtg4DTsIcF1c4Mcnm2ES1iQX6QmshykZCkBfVU
rl1bKqnfS+/iH9ApW2XlqpFpOamOtFz9wqo7Y1/h7HPkVwNSd6eiyusGMcUNK6KVCQU+fnsL1FZQ
gjAOV6fab5Pjkokuf2LkjfA+BhMC2Hq8OKZ9oct8Gofbo4pIXIj42WHYI6t8IEvxNUej6ImdUdA8
Ud+3c+anGaW0qtUWWV5pzWMHm5YhGUQ/uYdVuf4kD/nYAgjhRBTk2cwK35I2Qz1mb9W6jHtXLKqV
i6VXOa7HloGOIP4GzATeFehYFC08t16gGHarxZjH3tJbhjJKqmwXcWho0Z3GCo6IzsYPowVJ9rBW
wtsxMu1kySeqTdj8ErE5+5VG4TIuz3Q8mauX0Q3tH2pnPwFJx1L4vMS2oYxaeIETgWkvbGo/xxk2
97P02T+tEW7t8pMZkXgbAER5p7aqmVKe6WLiGUfGLdTWciWrvUHQko0HxAbN+JYkwJKtkIWbYH/2
JIxBNnkwncJjFNW5j362rWj/BlxXjak9+KkVpZowM0Uk3mZAHL8TJjFxM6U2XgUpcTAh70t18MRM
k5gjzIQSIWqAI4Bg/rfRiGpfYRdc2yA3J69oYwsNx64dXhgKBF/IyuKCw5KluSggTPelwQdQnMsR
rx/fEylQ2SvSnDe/uTGA6qmR7ZjslAtq3sgM2lXJyO1A30Ct/KGntDscaQXqPV8xlLjsTeEB58zs
3Tya6s2X/Kz6m0FYWEURZxGBuD7Rbgfs1en4OxtDgTUCktDthLwU966Bp2VoUp7hLZMIMBb7Tqcd
LDvTwML0Gj6Kx+hlB4Ze/0S+A4PXPp+RCQJUIBrOkoOJd4BPtUUCphplW5tw8FtoLrvlM7hr4oYk
Q/ytVVy43aeNCIXN6cZBlFuFn06tLIbXJLvWfnnxzpLOY9wAZxSL2CkK5JYI8gIMnb9vJuPZLepG
z50WukRe9vXusgCudjRA5/PoCXd4ZIm6uzaQWzStjMh/80PPWDdLDvaPNboNbvX6buikYlo4fj3H
bzmSLfpK0sEcWsGhkE0TGQOhhlJeXbEt2jrax5nK6FuShxxlqIm1tQip0yfTCeFeZ1lSv0AGKdOh
fKSXpKBYJzDVNFmT0UK/Ldhx8FUk3rfiaAvu8w2qn2yjbJiCE+bk/8JKDSWQfbKz0bVrsr83/V1b
2DzqrhlWrgumWj8NuHgiuuifD1V1gI/iz0J16TaglapTf6p+jdmW1bMLco4zp6K/X81yltAud/r0
UnJ8ROQO5JwVtiMY1o1csllGVFzuT3Lady65+8gN+9ZrmOt477UhQK6PeABzwm5lzAASaSQ9+jmV
Z5ihgFGRXYzLEjj/7AAkKOrSFetcx5XmioPBSAd9nqTUu3yXNou1POU5P3TOEuDwbwwkoQXlfvrg
6LOyJ4xmw6Xbv5EqwmNQekSpsP/kIOxsDI+uB9c/d8/athbKQOOABCkaR5ugFmqJyTewdsgTJJoH
5TSbMBub/UWz3UxARn3lPdGduz4laWmLrh6YvI+dynmS8DJaEAHCaAqk27rsdbBk87nil5NurQmH
/9gDIPM0Yapi2lXmlgiX+6BgxYcPLpj6G30IBF8jRdqK18zBswJPgBXkIBZa/aWQoJWB4yWpdBpW
UeGeYYsl5jfJLSsjfo54HewBdYzQptsyxzUNmd1buBhI1b6JbFo3S7LRY09oopnbePtPR1q749Gb
gZ83Y8/GRf06PZSljwXF38W5CfZVZxKmiV3EFvaCixD1n/nVxEYwBSVmOeWHbxyEk1JJQMyY3o1x
hUa5KZmOx6y8Gmey8GZ2wAZwamfaetHx5gtn0P0RF3FTLS9lKb7TjbLhNcFNsw9No6UxXRVePHBZ
8fV97Oc5tuCZDcfgo9CdE9V1FBSbA0b+3iVLYqpQwsjtdOEfvgteZB2/THkmiJjFEhA4XdTM7Bnt
+2jK7jlB7aMzUunNUbLb9nfhzn++UzgsPzxjAehXM8ZxPSMIbtugO1i5KcXOcM5GFOzj5Q2HFc/F
CmO4NgiUSoDarz+Tf863xYy/ggpboLzq4/c5C1vHH8Z0m6HcktEF8FA8PecemQe4AvhTnV5lWeQC
9GQ1CYHXvlBLhhfpJCBW44CHN0gV4oe/VRI/HuuOuus7mkr0Wf7AIVeHN3je9TW3Y/L1unu0C5z7
SDGtnPym4PQx8yCLhugVGtybuGXVMT+EJ5sbDfm6rZegctL3bsPVl0lkuLZBGBDXbRMe6pDgVuRx
DKvDVzEtrZRyECHONw4g3x7xsHxNFlR0KZAP0EO6Q5og3eOl31xTDejOQ45MDD65fqKreXVO3+MI
hHufkmfM8OTisCDmyXjOUCLjcQgHR9Ni52GhsMFbJyE/g38k/QysbtNn7xiQe7rnD++EEM4fKrsi
E3cHhxNECtuMc2eDcLGWYFRyDVupuWmV0REXedwBy2ZSUF9GJU5BPea3YpKHdR+yoAu859bm4iyn
LKWf+G2fa8bq+ZXPmR2AJIJw4UTMC0yaj/zbWj+Jm52H85aQm4dYwrmln/2oeOsD2HwUM/zj4yhu
c0Fcr6rzzXUtwFEZUJcKxqqir6R8ZTi4znQ82GL1VuYIzilirDcYcaNNd3vmsQWnDyVHnOGRnJFh
EwRCHU2MwqXx7s0g/qHKXDBdvMzVTrtHGPeeJ5O+gPRQMqmRuFTkVqOwBYl2OQdyaC7eQ04H+PaY
H+Yz1UDfHgY6AnLRvGibaUod6YtcpVDuNLu0JqzG8mQCD/M3Hp54Y6ysThpfnclvp/1neczuq0gX
0bsRg7O4VvZQ/Ha+hqCQ8djfeZq52V8qAQy4qs1RJmsrgAhEeRiFae7UmqauPvQJOMkQBEYIdyN+
PA+eO0/9PLaNWjLUgh7hebecVnpDRgL3zR6bh/JNzz9DSPR2cNKXiF7hrU9hX+WGLppC+R6cISF0
JgN77xdnPWT+bBB22e7jLBADV+NB+ZOcMC5p00KFs+ROJgrtYsxcyB/JMKQd5c8Lx2ZYmo3Wv0tV
FeryyhG6AU4IKLHIRl4kVsTbkadF4mu8sFE30eK6b8OoH9i1yFUQusuGosY0zBuF5A7/89Mdo4d3
dwSmOdDZZQTvEhKXKNNLXK9fhOw2hZaHvvlyIrTYVcJx1IP7SZDl5PIEp70oCWCdRaDR7khz3GlJ
u0+bE2ctjmqhHJn/NQtjvUunrei+F6OzaDjo2RD3Hj9fD5V7UBBmwwmllsPcVUsLMHF9XLfa0mEC
adsY285sHJxUFAnZBQAgSeKpxAxKX3tIwt8aZkpJ0X+4tE/6c8m7ixTLMJHAZf2ieNr6QTTSGfvT
L/s9FlnkFmTgsvTzCV8VY+Yn3nMbYwIzR7OKNPHBp3V0pqR67qF2lAmqReDcQa5lFv6eNIMihqta
suGr4AnO9tWKjVcfBlofvN3AzL2Gn5Ad8kjna+v7lVP6+RFDudJXWJA+q1MhoihGBs2aPvg/lokb
hIA/g83hJoVlRIA9oPGTUe9egZLfrXZVJEC/k1Bkaxvfp86iZk1uW5wd+lEyxo6XhJ7wXW3QkH3Q
/Rpx2KX6ahzXpyZaDSOJmUKc46IE9hqe/p/vzHLkAiFLJOCSDocGMWYRwhheiX6xoWfR/m0LirjL
xmkD6Mhl/wyu1nGGyy/6pbai2UtKY6Oxhg8zDvrxJz6Sd1ZN44x9Ggfr3RY426klvPqMRNCKn8J2
41vG7WhVgyexNQAVEnq6UQbLrEBL1HuWkGNweHEo3aatJTilcA9R1r2+C5U+jtG1WsEYKdJrZ8K4
LY7kdoWGJP0AIjM5Psbx+nZfkLEJgXK25n2AsowsJmRPSET+gvqTnsOLkr++v+Ev6pxsctl4Q5wO
t0NGwpvN1uAy4jwg1n19hvFOGlm/hhM9tVpu7PCDZqNF38XWoi7XWs/pwTKLsKP23QIOJ1k32/KN
AJX+z2YH9IxmU2hpr5c+aol2ZKkdClVgDdqk/DuJkpZmM5QtvYxYgHwmME6rwsvIfWEDMAWAcoW/
11T8qDTfCVZh8a0hF/AHxsCDlJln361fzKANa670haF8UUmOop1zHxT28s5Y0H3LHnsVEi8bFZkq
ijHaj1fpbbqFMhufP8BWmhj2rEh/h697jrwbFOx4jpBpVMskRBZUKslHwaP9syUTaYewtOV49acx
+0t4mX8xNoVU7U7G4tSzzFn20jM1X/B5AOLaWXmvPkxTXa/WMdDYbIf18TDkoNkmk7w22DJx3DuH
ZWfTRTbrlTkXIvy8rO3nz0ogZy++/KxOsI5EffOKC4CrsrrxN2jOP4G9vP5+w2yWP/+mX4aImmzm
4By+GYWRcqeHM4MbfhxgmPYsymPlQ+1JNzazoI4TMx1G6QYaC6Gfln3JGEEFtRiMg2e8W7KNR6RS
b/bQ8JM4yjc4e6PHCzRMB0tzwc1xTK1y6YlkThhO/gHQwSTYkNq8WRlYW46Qe1TPTOSMcwPlpanH
21acffwJlas31gmWjT1obJS0XrdGSB+ERj9JCpSEQtmDdZUHKkA7qU9qnx3v/ZftmEBTec+F5Bh8
WZpWMckBBeh5K53N6RLKV4ecBiBsTYmhJA/frurRrPy2OVlMEhPlwmne5VmzaQhe2w1V6RpMAenQ
rsMKwtZvZDY+nTpduyzQhzN5qnV2PLTEPeLkWEvSQpIEovIixFuj5Pw6GGHc/U+x358xspsvM7R+
5nT2jN0GYebuRquz6SpY8SM3S8B3Zlz4EMaP+x4ODO5tuHt2SAamYg/+M/DFSGN69xasUD6P3/XH
ncVnaXv7adUdV1K6hx2NcACK8FrrOpj7G9NVnu2kHVWt/vBmpizihApC+1CwVyzlDC6Wy0x37GMn
u/+Wvp1CpO2CUpzYa9n03oqAQhqiolT3E/h+5U8KFg+yNOY+DtOryVZh0wSNc98yxfn2z6a53qt4
XnT+LT/ymFqwGoY3hJ3s6aZisu/JXb6aJS5hZvsvyHtXqyPq5Qb9ZNamg0/L3M/lB0iYj9j9FlX9
GGmubOuGmo2ENuE1bE4YGTkpo14o+SlXbhXoS2JYo0W+m4l940g/GP3xaLUEcOhxBjTcxaSEXeFn
kCRnz9CHmFqiyEJAhnGWkJVvzBC2iH8I78X8e1pB6bpRmVirM0BL778oTJKZE2lz0Tam6nh0X33c
3QgMGVkMdoC/6WM4HmOcLVpBVu8J9icxToOImrT/kJN15uxK9urs792bcvCo0giYc7kl7z3nYTaj
D7s39kZPZ6twJrB4B3kUMqlT6W8xJLyhZfDKtNmVJrDQaXGpiBFQZUc6T55Lvck1IW4boqm4vxEL
81lCHdaq1XoQQc9tahHTjnYvj0/OyC9Yw3h5ZA2UZ+5/QYUrUxjD6u4GWIwa+/fBX4LBVRx+jKMJ
7CVFa7uLMsERzataH7yetSXq1hxXrcroC1gpNMoAddZMwG7reswoSTSpTNokvw2zNA0T2pqVkGx1
ftE04VyFM9bbVTbAkUKOP//mT7ARkwys2HXbCSySGGA+DUGLPdjvN+cLEK+ahlwd2vMHtB0zcFHU
yIOnzD6iOtwSfdMsC7u/tPyJfsmZKrRTOBVRbWm6UJG0xQsk2wi625eoJ+ZSgZcj5V4ZTjxyBXKV
UVgEkQHfHArTo4FJ9jivC1+ttoy4L6p7j1VyKp/R+32e6TcBo/j9F4DfE0PIxsNS/8ufLC/A2Ga9
6TkydTZvgi9NaxnYkY6oXKh5D0/92rnzGtU22WAtfukGJxZ926b2S9iPUUqhmUAd+whnI6KpYTBb
RaKXjkscd4Q7ZqWKAij0I85Xy3t8kSL4LRv8QLQYydkKOXWHQP8vy2ah9NyJCJCSNDdqMYidDU8C
lslaLHHiABSHbJGRWZ7tjDdk+O245lZq7ByQ4V9P5k/9GmxOdTvAt+XQCyT6g2dqsY7+IgYTq+8Z
kgB6RhVsGpWCk323lrN6OR1CrXWtnaXRfAARg/pvpNLP+gweEyuzsN1JWefK/MrYtyPvVYUMI16P
MkVv/nymbjTowsC0j8ZDKe4d7HLIQE16QAX1M/GHaYErqkKdrCuyCzQegkc2yrOoF6T/YLrEmNIu
sylLAp1wtXUbweE0q2RSySQbfyDT9UyJ+6X66pP/67DxvTX5YZckqiYRibvwwIE1jCpxyJOsCccA
2WTV5prwHWRRzQ4LP0BeeMBIPbwkNYh2pnq6ai6IpCGzfJzEXtqW09Armo79J0Frc+G8wijk3cXg
MI4uK5+FKj6f0RN5h7CaFNCZ+sZeaFZMGZEuEy/rSezD3jrGa+Wc1p2k8ZbnamghB6iHRr0laJZZ
FUSaJJXlZMnY29z2EY05bk9qEBd1EoOeJSK+zV882+q7hCPjR4toFEpIK8tUyIZ0rsoye89r/X7O
J0Yk9UuLlS7QgBksYIN+Qtybtd4h8sBcoL1OEixzxdq4OMB4t4zqpD8n+98C938n3NH+vL+SDs8Y
Nllko8b7J9HC6g+Zm/cuhUpVQCD1N+iQJgalZICtVHpiI/zPaZCtt7wIOnZndQWgbHySaNsZ6r1o
Jm3UNdgpW/A6d+ducHip+k+FQJPACmS9u0iPX6HaH9SiaxlZZVB3HAD/1YVerDe1ZabNwlUwpAum
1DtCXSST9JYWz+9iQrL8fxkVNHypz6BC9qfiCiQ3kndF3n+cQtYMxG3khnWfyoRaWgWsq8QnxfiT
FSv5x4BVcX5q8Yc5VAEdqnIP6lg+a8gQSlFfq4emCcZxHAJQb/EnGUpiwEzAdBBEHLgDAunROTC9
GHZfmwCyTo7I8vVWgxBAaHdOW24jY2BIwkxRBSllKvBB6S9R/o7qF5OelMt6y2Qzqpi+WKygr9Bb
SUYTtZJ8A9kBuPGJWEh+vMqCouj8sgGZB6p5SQ7nF5mzodn7tMwejZy+8TBoJYcbdeqJyv9JQBE6
E2clgbJ7bmvyin/zPEn/LThthn5jpkT49DVq4rUEWzdWro6ZNf3OFUr1uXBNUeoTXMG6RMNA0rE2
3gJQ1e611xFaut4cbSIlPF92VoTweIb7AREvA1nx5sNN/fUpPYggnAYSEPMQTycSEhpXSj0bLQN3
ctGmZNMat3XLhhNogP843vQ7X/Mkcj2othFvMp2L/+lOB4MQ8L6X5NCDdGCfR0hnJcd6Ac8uBJYH
dV5VqFWrp1+Dmr5McvWiId4CD5/u1FUzHYzPbM0PkxTuk54wzZ+DrAW9m57PnTiNcx0ARKUojLrz
7dlYmE4V4wqOfvY2/AE4WBUHQTA+aGq7QoZG1vL3U7qBpXjpSQXGfA3qTkFIdH+lbF/8+MWtRaX7
k1GC3m0B90ZmgnS+DS3idcWmAZ3I2vxnefKiMYc6jpUvDt3XUzGa9/+V1fPMHFJlZ3E5ZgFG+lJx
jgjN0D0Qwsnk4EM5x3e1kU6TkTfVYz7Kvc+0hXR+x45gtINIKAcm6ITtoybhvaGVfNYZaQhEth7C
Hc7WePFagXmI9q9uR3HoAKk3ykmah8Mo9dqJ+9tNSWcELbTF7kN4yyOb5UzR7Qt+y4jXacILVeA2
8l+93Urzrq2Y19dHBMMzL2deVljY0Ys963BMYJziBKD2q2ZJ51TEXWBODRVUVcEfEEnuYueCjv9x
6+rLImNc/pN2FEgveZ6XCbBf5T1GLBTSVRDMwnzG/wfCPNWcp2ukVoCIwLQakkv7MJvfmF67Tms3
Rw8tUbBsQQUbd84kfX0mHjTRD+huo4HlXelrvAOApcfo79bjgZPRSxiA8wScCtnxEUriaNVvF0WV
rCM2N5Y+359hEEH51tA501/+hDUCvF/3ht2I0+Edvj76WLuoJ+TVdPshEcRd6pcMZrhxqcjkOHNi
Eaz6Hf0BB0N7o65YzqwmqZ/xvMMliTHvD57GQtXB88f2CBXdSMJ/Nh83roerRWeNWrFGrKGvPg/l
BVXS6SvgwMfONfvWmpACB0RJ9urwfMXhec5vFGfno10RWjimbItN3wPFKjndI5VToKnK2ywKg4RH
EFDBzR/Ri+JIsDE/4oU+YOS/bGOtlhNOTUPQ9LOGc1Q4wudQ48oHh4XYSBzW5JrRJYdG3XkADxak
8MJKAQT909pvqBg0CSlSRWecp1/Xv7iQRN5lZpORbGDtJ3nU89Tj1C0vH6SU1D2tkIWBW2yUathS
4wF87mBEnv13BZ1626TqZ29WZp3MEsydJqX3Ng77vyslHH/nQqKFkMDSGrUctcMwMa8sGlG1L+lr
/ZBwss6dx8h3PRdgbbmNLeTMNYazRJ/k5R8Y67K41sCPexBxMAFNsKxxFgqLfVGCsn9UP+MAFmIf
y0q3HE6q4dkALlJ/UvW8fgGOr6akmiIeVsyD5FUOAwS+1hbo/g+OkCAY++M6cXgHcd4vlG2AW2NE
PwgO+zDi19L1SsnibhqPXYzyi1mvyw9x1eqPFURKov3Ojx8B523MXNoJKKDwzEgqBesy6ByDMs0S
Lej0I+oLpO1psh6SEH5cI3GLfaKv7e7VrY/kiNSVvQ9dxp8qNjG+mR4sxS7NbVR9ySZZ9yIB+Ri7
2B8oe4UaBIbHzRnSuGIELW+rC/oWdcTLsQOQm8PLhy7smZFRNCbLU86QYeA6JFAn/Ry9zL6dSSo6
hC+z1t9S5l1nm0KxaUeOmUgerQFCYEXMkbEiuWQJ+tSVZ0PXPobmTWEwGOGLBIGZzGfmUNUkFnLQ
ejISYNdd2odBY+ZddREj/r+7ItwyRdelnvAsu9VMhFbcqfVWlYNNAnRh5B9zUPRrPBoDvxGrvI46
CnXIcWx04BpdeRAilRK1X96d2ioafZEEpBQ8WKq3g6J4rphYnARnjB86V3ZpJnyt1WHW1AS0ZOxs
CTZncLgYDa67EfdWFRFw0SNzTAHXEbW9/Vk0emwfoade+Frwu+rUadnXCZTpedOzSWkKxnpLpfFX
+K5uMxNmf7u+MaU8EPJ4n8hIfd+oypLtJsBGkMB3u7gLBK9zAnoC/Mmk5q8AYuAzLbTWx0Ro9U9Q
MadgHN1zuK+qaVZabvRvLbwXOh6DpqhGkT0OT+/WBF7oYsP3Qj/trDJ8P9r7pUnfsm5T+C3wOI1a
eDy3pIwKUN5PvH0XX5jHnghSPMDs5zVwlOKHy3AFf/BaBSEY3ZabIbW2+s85FC9tOxU7xFwqcQsl
dZ8kbHNGkSr4d6DaXZGB+9i3xvvREV7H8bLAI532bcbY8GYsK+3A/FkD7L1BiucAUGqLtLDVaNJY
8lItz9GYFW2ztThS9D7oWEJWLdQuk2SGDQdapXV4j5jeMzyB1BFcgKItoXf2Xll6cT1iPmngC4Bk
mRKZOQsiTubrNwlro2fXQWsNWJqHLdCI4g9/n33QKI4ZPG7zpk5DSvV+ut7JsiaRk51baYcJcu/m
RQ+ku7ERGiGDWHZyWvzgyZlluplZMPl57w+wueqge+pgLW0n2HeK9a4++Hf5ZShY7rlUCVoz+tff
vh8AS/2NqFNmBXO6odxh4TBEJXgxvGK2XRPhRie5pp+buJg4IEut0oyA5OPIlHsBB82TdvLx1E5c
tYdrX6js2HPwFCxDwuWuNNzYSjm8yYgq+KLjX/ynyMkt+dVKGcZ40YabqJo4ILcNnPg2TYTanyk2
O4QuwRyv10gUg8+sJcsuWg44+j0rPhPI9qdwmMzAbfRyx/KkB8ILa3thFVq6YKSynVDY9U5TRnBm
ZCoAzlmcM1aHqUwWdUVT0Crri17Kc4sJijZeQEcrc/wA7Bdg1BNAreZBpnkBv2RQ+wvrBH9wSbQ6
SION6La4UQCLN7rJsOzqRmdkdbZV0NqccLYJiE9v+EZwypBfMJKa37xzyQSS3u16PUqajUNN7ERM
aGkUNTOWhEYYGI8zXoRsnfVRZY8X3Ox//2iL1IIj8H2VXasFlkIRHL0LmbTZFq4/v3L/29ofxEe+
OOuCqev+cpOexfXtlHXol3g1tIukdLzPtaFcGqPUWGPLvs+WzR6+w7BeM8hRVVSnp7z9ONdORnGb
H+CVQJkzxEx4p1i9D9nw8af5ORq0yaEXp+OnyNCnkc9YpUBOzkmVHsQ6MtzC5ldmdUgUjQqIbHs3
+MC1rXU8h0cU9LOh//VVdNvT8gzVg3x2kSRL8O4EQ0Vq4SibzeVSf35Vz8Iu0fhzpSXXCIdr/Od9
mi7TzTw+Quq8CYh2VyZg+ya20bYub66WT9P/zUB6Ve53jzHz5ML+qFOYLDkGJVKYDmpco/sHf+gw
kSp4nY+dLKlrWcXod3gEuFTEnrplpfqWitdkwDvbJKvZxiURfPf7i4AUHrk6OEAYzEqqZJysmwWa
sKjvzoSLyBFsXQIXAC6GGMJrjfYeN5HeBhRXMEDX/gxbLAMMxSC11jf2GF5sWkWDq8u8FF2yCwpX
EvV3pc+kd07bbe0Nr446ueqtVGxEn5NbHz5JBICiZsO1Ipn682Rs+gVEuqclJM/ClVlsd1uVRIE/
ZOUZllAM0PFn8uKAYsui/4OyfAbbxcLjkb1EUy1dcxfog6+XcuXTctOqbp6TsHujRmuU+Ud6IHrh
EqKqS37RaJ22cgj22KC2NNvNT0rNeAyguU52pLFJ8ahxSB9GrENvnYGMH7jU7y/VUaQakf2C8qmX
nry7eXaEbgKLK0nGgVha2H5/4gDcD9Ewp2wF1SDnMU8jQcsxtnStA1cg0esiD9B1cc5Bb6MhtMQd
60taNQT5QqJ0Ako/Y//tUiBX47izsaIk3+MnZzi4drqC2FPbOW32nthWdz7zyZHVjLAm1drOwBHk
nigi3C3NKaqgABaFjSLBbSF1WBtNXBHfp5Hyr5PNgfNCOOT6FAvlfl2gIXqKai/PoBbfrzG+Wkg3
/lr9A05HytlmgtKR5iWn13vvDGraogtDv8OE4ckYm9rsJ+iwCRhYaYWSSmg9uWvaVHJeqAeYDQxO
yQVXHEn0GgDg0oyRTTv+hoZMuKEv0F0FmmQTFJ05WixdcY8CDDAp5evmsV9VXvYlhGIPkEwJxyda
udul5qw7D5KGQdm7hrBpCECU4sKY18hF3QbKpdXrK3KQxbnCQeM1P2wuVleybKLTBmtuClwHSuXX
jd7a/La3H8E7cl5UG4cDHZdidGGG7YROjfeiz5pmUMRl1U2Lwejc1DbrdAWVXiCFNmWKIgyrRSPp
Hpq8dpXpZT0TxDpMKg==
`protect end_protected
