-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SpXWlgx/iv5qVqGwGHS3nfZd54Eiz+2MtPJFJSU9/V4yMBu0S9eN0gK7pCS42ypWz9yjv+5qkcb2
Bn7J0LbqI7q3rx7HsxeneIYV5Ft0q7z3Gd4D7z5jRg/iQC3Kyh+bjT/W7EoGX6oAM32Zbot74dBB
Fl/QOqUXoayp7t6F507rRch+y584l4EkifKW/CKW1XVdlvMdCjWFi4tsdi+eDrpk0IJNQasPKCDL
7tb+qGmyAXOx4wAhViHv5lnKISxLxDNWWJL/IAKusm7R78agl0D9DY9dh/D7etCwwM2IYufdr14k
FcO3185g5Nuyz19E3sXxKqXWqrGGUdtfSio+5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
h+8I613LPiI/j7Pz4joGRLj23LnbrW//x22TpRcKUlwDT0rJnLrWA+zOrGP9Pc/ESjTPksUGHpAZ
eLSZyCe/Gfj5P90JPBAETvmXIED3Ewa3V75Yk9FxdKKatAGuOJk/VXn+GCHEFJERzlqrrH5kHQ1o
3TdOYW5hQjaGiWAmCnt5G4UYXYY55qNeM8Kl+r6uRhSqNohMRUZ60KmFkrit9Z6uTV7PEw7Yyuf6
inK2c9RNW2hIOirpKrnrjx3+OtGrQ3traPsQm/3ZEY+uz5XgLP163+xSjFVPP9Yt5nm3CNU86FZ2
cBvSgD+/sNOUkTPAeXuwBNNB1//5jlZK1Ao4ctkTvbnn5zSSsPGcPkbb/zXIOaCOmuZLJyEzqQR/
lCdvBBDFgyxp45KjjlAvYkkZayli52TBc/j+Ge0iK5CNZ0OkP4BH0eLlB4JL5I8FUQrWdy3deuCW
lym3d/2+B/qZLL9OalHxYiC8H5QUU0Cr+rjO/JxFJFVbvRNN8/WyFRjMGzgKmrIUw1C6TLehX5tY
pytDU3G0Q5jBja79e3ilAaLiefJ/zboX3OM+t1xQd/nzINWfGy43CzSq8DcmKY4vLx+n4nRU3B+l
4Zq2dDt0yd9U/s/ScPIgU+M3k3b6UsW0lY2eQm5ZnL5sm4mSZLTPK25XSnul85gqrLpoWDr17RZH
mKb9K/DyrLWSMrW7kb/GLidZ5WYcxkvSC9e3tpndNAq9nOHiJHgnxax6U/2vlJ2PFR0w7h1BoDqW
Th8tUzZOK/k1SHc33DxZAOySppN6WFNb8XaF6q6ZW3eJR6fAz6rbfu6Vi/doyyr9FPIqFyonCHvV
axZvxBbOfhUoazX6XnHG643Vbjqx5MBq3GuNBCqXxx/cgyyV1eFYViSfziFu/Ax0G+oplchpeMuo
zmXnrlgzY8kwPpoDOfVoD6QUaRHQS77vzjLQRvINkVzIXTcIRI0n79cqsbn+tndJVjFi5cmtbHnS
Qy0AsbjwFe2zOYmgHIkWh+b/niujUicqPRHKAct2WM+nuRdoMroXKbLD1cE5uDl3yZ8avP5TYhEh
CVDYbYjoaSYq9jwMuLBMv717Wz1W25I821QaGdCccghikAOhEqDk4KZgF2oW/hnslp9fZ0NOsba6
vqM8mKYBDbLBXt2OKBleFqVtPJh5VA0IbmHMVpVlRsjf7gkid6VLs1hMEcMfgqJSPHn3RNGG9jil
HHxvFfYpEXsaboHP5fK6fkOtDCVb83ELS6E9W3WeajUbFYP3n3RGXvI6U6C+RuY1J5LMQgoKT9i6
5eZTQJsJqdnPp3O0pn7oOt6FW8MtcjiOhI8H2svBqjsWnmM1pXHr7Tb8JkXDAE/0QzyILRIYV9dY
zDUemZHfy9AzIaOmVx4X1YzgMm1y/ftt/9c4T6sHpMpgWUDsNINjX8D2PguLVhcOaAyXwEk7WNdr
jBl7b2hPq+S5bj/GA/WicNAgwVjRG/iUqWeCp2t7tXIeX+pWcyPqKZwLv2nuzM6TtfMKmRn3YKhG
2zHXGtQ8WOObq4HqwsJwGoHwFGu/2iHZuHKcELEml8B9w8tbEtdzvZpbOzC1NFPIHVWw+h9Z4wuY
1Zg/Sxatp8l0YKsZDv2SMXW9vLHZLoVD87PlhLvSbG9+epzpVKrBA+C0E+OtRh9YtXv0y6LAgoh+
/xkcukzGraqRi2zbVn+W5x392coROP873J7chnanJ/jCrPLT8LSU13bGFSl8zaxG7vGaTFv0T2L6
L7InvdCAuUYZ/A4MhKZFgYf2/hlQAcRvnnF+lKd2c6AIliHHgqWmAF1oBGHgbXqPfkPwMRcIhLvd
PNODDjJyV62P4XDJr4oEVWF7hrpW0CW8u9eaRTtRUN1Vb+s/eupsrzhp4qeSVEQw/zXm6r26WpbR
9LJBHBCskjtNsmPxHXYY3oJ1haGxZEHq4MeyrlMcay/aSikzXJ5gtq+6MlRKnL19g5fJd1P4oM0m
EVcGiKACBCc2KsF8QvkjhybVkyu+To8G/pqBx0RyMLHIMBOzNNVAgdS1X+ORyIS/hZv/5LlEUWXG
xXtwkq8mAb4qcFcW3CbWaVibZr5z759QQh7U+6ehiOg6oAbOD8P5/l4/KcHM/SioO86WUxXlUAru
tskmHiMsNIx2nN3073/HGhIlnzcdzIet2YSVZq9NJrJJYlAeWWYCOU63qk+wm64T7TiqMHhXfcCh
vwsm5F3FCgfsMNMgF0eSdO7EkTwtA3mnwL1bY0JnTsYiua3pYTbOOv2HJwHEOeCGQkdFp03OVUbw
BbShlixMFBFJ+lzsrFJtcz0Tj2LTovlJL3Q7F3VPhXwUqGVi4FsnM2Wcd+1FQ7xvTl+l+uBPYCLL
InYpMQ+yCjMi9RoJS7xYY82qQZ2dozHqi7ADQNvIFZ0vue7J8AMdSrTIwc+hW8ih7iGfKCSVh/i3
5ZhOc/IzTmJJjMEZP6/Vq+XCzwn5alxVF/mZ01l1AiwiV9Q9RmbaiWX+ho2Y8/XXrbzOM9VfsVzo
cM6cgueIagO6EPtaLRXcTSiqhLcG3I3ZwlX7xYMxRipWP6nm4kJctWy99TsoTtWDNwigjOYFjImb
H3O7cyjfwDfvyZ1NXU3EDFrlu7G5mGf0mVvjJ9xFzkBz3+qSnQNEBF1GtPm0NH9WOyjBQsv4QSQl
6ATdt2+ZU9vkbWj2hXrplGMTobFVhV9PORTkT5Tazp0VLZTOTXYhk4c5+HWOAYpVdItKhyLHA6Xp
dUygba30vHkaBmSanRkTTBamhs4OTgDt9B9+sCt71dBeU7VuirHI6ewIvSSFtLbaEUnjWKKOjG2d
9K6Agj7t6kvRlVR3KH/rdCD68jm49CnnW7ox6pSPw+UJkGl+HHtPXGkFlC7oy+uExQrHCH7ZwtaO
TqDsXOcujoqsFvMZ+j1j/8IbpFeshl1jWtUcFDoyGGXt4ENtYNFh9DtlxoUPvdpR32W0GtU/kNNZ
NMZ12uxN4Me6+FQKtN4VgOeHhEdVR1eyMz8WlPs0VR12u4w94RrJKXo+LDX3crhN2HmIc/3aTRuO
6Rtc3ooJQeKtnJrerRbcwmx9tLVsvHe50Bcn7mdopES6VTp+B+c1mJPMNJ1htruzfL+DiBO62wzZ
5ikLYGbIwFPWjOk4xMeZwuGRhwqmCrg6sdq3DP0RrQNyq9jnFqURqMPqos9YWrjUC2wxSXCgP63x
8OGQk/br6l+FcsIDIWC36ah6bmXazf5NyMfM5TNiarp1I3Xb5+X4qylw6VaCnMJbEX2pj8QJ7S11
QNdvXhkHM7ZHAkJEcsB8s1muHHEed4neMPUM9bDVp+iqSoUbiOJ8FHTzYZtxG4zUZhZHYF1eHqxy
cuscepMrOatf00RE6DS1u11847uPHhblMHpFi2xif9r+9FQllAm4fUFlKC9XJptRAK80iBi2+2fi
hXp2QZMh1srvCbXw0Be83WfNHVcaRXSLbBliMND4IETxdaZdl3nDVQSRhQe+Ewbo2Fn7Xufy9Hk+
xScpShFVr0RV5Hh18cVEbljOdcrUdG9fsuKjHPXf4s8+4yG96OXd2kgAwrCpMvDYDsFZzT1adusH
a8/tspYYjTJz7RZmmAG9kWS7l3bs3srqB7E1Lc2Sn4yvOQ4uN8YpA+4xQWkILW9uMEKeFr8kcB/5
b81CrMHODvIS/L3gPbNVD9MbTDH2X5LdvH4HhUIrv9EW6hjDVCFCb1TWSNC74sEg62UZlBkDQK2f
fcbssD2wAjmtC/CEkh4Z2DoGbQ2KonieavC/3ksSpuwIrLEtdLvWBXmHPP4DeyDIRcYkA/pbMrPk
8aWmYlhaIHDj8EfYQIEjWUV4LPAvy7TudZZj66tjSqs80zvuollfn9nGKQmJ2D4F1A/4+HgmD6we
uyvFBSyo3rI/ZWA7vRyL1DZheI/pJOC9NHQYPOxwK/upDB1zjos4mnNKOTQG3WcPaa+ZpOr381ZY
wne0Lbog4ivkOa0319XAG5WxyrY9GvcPtFlCyM1Dr61biwP9VlII30PmKJm+n3HXCXySgcdtqeHo
x5MJ6ESDLg3EScSDEfA6tfJneCbs1GJM5U/6B6XQ1O+3rvV3BrheiLAdPqnWu1wmJrYVctU49539
TlHvexmKydj7PPw+VGaiOtWmsdm24O5emeJH24w17nM8Xv0OPcaMMb8AXnPAi5KcUk/o/VqoTSxa
0AsyKmcdIsagBUxU3cEv6R6zBUjCtMvyDA6xYRlYxhb/Sqq2u1tgKlKOzprKrItGs7FUbA7rvEFj
a7SQBK4cAZM2rdwNLZhG6D4z8wbxf+Jx/uK+0XxivWONinVEHSQLAYwiq0hQv0nei9Yjig4CyD9u
9Pf/zkcgoQYuoVRcOPCYpJC7MSVyCUODfQOzTvUlA8B3xY6Y9FNPo50SeqVvqnABoyPVP78zuK8z
Vbma1jRhKAGFLmgb2KUP6kuq9fR5uVWcc5C//4NOs09yZGq1chUkFUhFUlTtFsxkWDDSv0CKO0Fe
Gp3AIZt7ldlcZwuMJZ/h5+ZMQDprnDJdAmDMDskDfD07kUfZ+r+qvQ9yesf3o26uBCp8vBCUxouY
MYErisBr5K243gHWEUOK5qGCvw1MFxvd3K5QhWbkNdJFY8a4DkPpAUler6+AieQnt5wTh5mQnErq
wF/Sug3/muNd8NtB4M1lvOaJlY9kIKB+A3/Q61Apt93Rt5rtq1VvDwaXu9qhDDkZ23y2pRT7GIzD
jx4MycfbWJu/Orn6l4fxhP/3cptB1Er1NsMXXceCztfemRFLeiuY2Svjj62GV3OnwoFd50qFW4vq
KSeH9sC3dfnkGjFtgPi+ARQ8LE4jty2aVRQFHNga7HdJ7dcxSYhjVWKuiZCHi9tDOGu+shYvNwU/
2IMNNW4CRzqjM498aO6Yr9P3PRlH8EG1Qec/kyTo8e6tPXwqvamz9T5hOyxPFQChxQMVY3jWn41u
96gAxgPU3RCS+pFoQbgjwET2Lfzw+MDd96hwS5BtjM208RkHMSF5DSGcWmbshcUHGIvQAGPAB32c
xyMc0cuIxlEQDhj1S0JknYrJSNfNPik0xvU4RCcO+N0JAI1TuQcUe0jo61SN6pPbKsPR+ZR4MY+/
F+6iIASaNgiWtxpjHHUDpZvec7v9GAYhD3eDXgn4yWyRzGTQvtTrs/oDLQXoaXxWGd1BrE+pQAP9
bB1/nNCkHV+q+0aZvPj/wUyMpPlNdpuqh0ISA77fTMMkiMNEUQ9cS6ugjR+nlio/Wl6YU/30VSIs
mfy2C+40CZaS723hpXaWPk7d8p62LV7KOzVyc2e7AvYSuCJuOzyHk+URiZEHwlIclewMfXBhhrN8
j82YPFRn5IDd9xzXTQzTSLTRm7oXbj6GWeR5/5ZmyD52l9TrmoXgo+AmIWr1g7zAkfpBuvYsmHqN
LaZV3rTa6Fn6vb3m1y6aa1Eaxx/bb6sLHQl4DDxWke+bsXfizn8HoWjP3wZuXodzjbPw61+7OEHX
sjMbQgf6Bup76TrMUrwM0FLkDYqPXjAEpY/jnBORSI4zmGyGGD+UByn0n6C38F+sN6Xj8curikMk
kgt0yNYDuXcKNVni8YG5Dnbu97YHNBc/WH/P/ckKUF+H7/WrRAOQqncafBypnsobjgwumGzANFAv
OHebduDaqFR5Rx/ibVAqzAJeTNJWd34NP1gEFc2E/muxoHTBvoZYI9f3ZnQgUz3vLQSdunO9HgEn
SiPAmcrm2REG7wT377qRytGJqKRiqsZ4gy85YGyvR2CSqiLY9IHGrNRK50UZe1BkyQ1xmK4SYDrM
hSpoPmE4MeUKcoMmmY5ebIEsAeVujjkx2bcjOZDsakhvH6UfTNze2ZU2mfqAFevO+7DFyNLk6Mpp
0XOn1PuQq9uD+w076tb7xxfQJsp6D/ow+haQpgtwfCWsf7FsrSX0FE+YZkK0QaaVW15W4Tb4CTAC
TyiiI3FHwEjTFvuEcxZp13f6skIu4xaBOPV8C5f8O4PZduI8cImruX7HxCF0qYGOu5ym+JT+GwRE
QEwcDOnd6qFeGeWUacsEmX0yHvH8dEaLDmGnSoLFDaVQ0H0jI13PdLO8VFnx6Os/llt44Nu49GKM
WVQKt8chp//3e19Gp/tE66hPl9YbB9TtG0kx7Y+YTX/DTrSwxZfS4q7jGdMtrybc8cERr02qcV3A
r91KpbB4Z4kK5oItE/jTc5eH8DwHlp36BniKLyne0mDbCO0iJ7ynuGEDpAhsIN9xqrqzVyR2bDwJ
Yct3kJ/rxKzsu/iFLvpUtlFZP/IW0VKTYvhEioZR2e/ZSsClteN7Tx43O//QK/Mo+fHXFKuQ7Uea
rjxYukx4m6OQcDlYwJi40Fsa9tUKuozfBxCFpHMAEeGn53rdRJEdvY03dMfNZ9U+kyAkDAYFRBGb
jrm1mnZEeHaLvg7mTUn/M/zy2EjP56Cqydzv5v5bRdm8pGfBZQRhlTu57Uccc9B42soTlplgOyLv
tmhOaM8L7ZvieHFvyv2Vs/94bj5mzeyyDSUdBMa2k3mg9z4J5xlmKDAGrppj00c+DFb96GeY3oNE
+HhbIz7qlLQ8knORvV8Eti4qhWJyBATlba1j3jsakaCwtpUpD9lZxiwmOrSXsr3ZR3tkO/F1YqBE
XvyDQKydnBXs9IbO3l8hqRR+t7Bc8qHpmvDuV9IbOVVE+H253qPya1XRqP5qCTXsyBIiHunQ0okH
GKWX5v/UwyD+KUISL5WkWKlno47rl1w9eP9F7EsIjcOf0NkD/SfVFO47JAjOHsULMdJ37zz4nzPJ
48D0Mf+RzXZgWHG40Sg8nxBzhiSCHmfXnLTndG2HwW/evpoWN5ygrcFEn+HunUoEJYMvCIBCbPVo
8zQILeaPU3w3aV2ezxs06Lte81nAYZI6LkBX6fspblUOO1ABdH0tPvlySnj609j8GsPxWLVzsLO5
Cm8y63tfup/wvXQsIwZZSaOxd5a+WlOTMYAASl5NVmSxndMeclDOvLqCYJS8xoYyP6VO8/f9kJ59
BxNne9pmPyJ38thYrpwAgPMjSt4l+mODBEo9ShF0aO9qtxvy/xYoXjDDVVGdNvGWfBVqjBfzCLMo
7KsunUirnjzIqq3PDNBuPy/hKM6UIN+PFVHyxFHjW1r2Ys96MBgbUovDtgymJYKpBGPS9VoiUii/
7qXYHjQbmjJSPuyOGxmQJhsmtIeDwdAjbIzNjR4yacrWVR2zl/LP9OMpeTOVpONcZTgqjj/iyEs9
D9j6c3roNXXhVGo+GS6OZiCC5TtpK0ePPV0MKNxVHf+mcpr/lihQiEqYCRC6b+Q4IhmhGNzdL9MC
JagCsLKJBiDlHvf2/U0fcIGVIhAR081wbRSzirMIymwb/oY9jGuqj6fdLLn2ifM8r/HU1+c5CiWD
vaQj2UVYI6oLKVJxwvFwF4OsMq/DPk78xMV7vXcLPPa4yRjJpoVRFTD46ean3Z3GES3yhPQOmefe
vPQ0MFm3gOvXnBNPd2K/wci03NUqyR8OrgfZLdTO+Ycre8c4TjbvzSt2AUsJFW2nkDlDGEMYzOLI
lVKIq/qiaSFpBKXYEFnOeVKZ6ABgH3lNWYEwi+pELEVW+ON9dZ2AUke7cPr43TTkKONvCwNSsOXD
mpJSGsUhUjUapjKpx1oNVvURjIyVsyiCzjO3L/tlolCfO27H/hdagkXbel9Xdi+3+DWo0DbPU8C9
Qg9O2yt3AplfSTeG4gwijIRfRqBtGpo/aqIGNMcJmEVudptvx3CVrw+7f99r0GasFqAr5vhlfZMu
9lSwDLO2V+VAJTy4VGNZHTlAsro9FSmhqqGVsvJJ7FE1xuZKq2Qd1hrHF0n64DUtiNBD6J6UFQQa
Qhjc1tKyKL4map1QtXyOkjdBo8jPOWbrdUDLx/FfGY4e3xtJ1sE5qcquOFb10YtkRhmJaTE0WAux
hka5FuEoen9n38CLN4a5yiPT/lJHHM9Vp1TQUPtkKVvvWvpoOdeeaJA1DYZLFRfTFF3U8Lyjw/3c
+QRLpMnZRz/0R9sqpIyEbmSJ3Kwgj9mZc9n7xokA1f6ZdRLW4PVgg7ffKlno8wqPlbBxdtHWpCMn
b+EnOp9DfS1zzaSMS707lCSmijMwLle9+l3oUvwG8F2AxzLGhLxEKKTsgzvc/BI8pD8S58iGgvGN
2UvWD8U6v163XiR6LwZ53znUe8lK0mvBrjBDiBYAdavHkhO7eHejLU+RSH9W5WOJ6kVz0RepzwXU
SmF1LgzY6FA+GnJsEZksVjeK2azFDJR+IKQf5+18k0ppWw70mCd92PUjsseR7IQJwNlmZXOiJ5hj
vAYsiROgVEAY62rVUNFsyP3+R1tBIppQ/iGvVy3wCCKk4Cf5hesHbYaowYxCCbodqEafGB+acZE9
QyNeCaLlj6eJwHJHMyvGAu0tHIB/nsH1zPusY8HnGKIoYgcSw1Q8BWzIJGYJLwGWhofAC62SCZER
SDcMWbtnKoE5fC41dheSKeym7SRbi6ES0vtlMJQW3RlgMmxNnqji/O/MjOBgoZbDRkF2B23+ZJ5q
hRK8zslEMrDjBsXpGl+vtlVMVNNQJ/7IA1y8BpLasJeduyxrcVBqS/LbzbdewbrmZKoTfFhnuZVh
lnv8Ss75UZUlyg3aw6v2pCnhlRWpc7RJih3kjELF73lFKgJF1WyW3MrPkJc+57VJvpkMBv4u0DD9
/pceWqYDiFc7G3RoTQ/fNMByL00e2uSZRAXUgrPLmAAez5ZkGrglMIwmnLokmG3B8SixmUoR701g
0+5FkstVVLuFVQ0cvE67cBPf7pBASMCDF7v88WUAvTthkzyeM8plZssI3SuBRascvQaMF7M+wgAO
F8n4hrlURrA2o+roAHzPKdOAVllyM4z+ZU2hiKIcAahNExi6bAIz6Phk643sBdhGuSHsO+nDLGhM
/YQxEe8G5b2TsizS+ZFxsXq1DPSNlFSoBNWAy11bjCEjaw0WIpo8wLzCtb4kjTDuNTxeA3aNU0bQ
gdEUtYkmjBLc9rpOpsJzeJu71n14D2uWxPtsEx1zqlGaunLuIF/+r3xlglaSZUt5sgRGiNRiTMcY
aDAObvJl8jNjXGlQ3xNgAStVOlX5FEID14TYdYyS7W9fKtRsO32b2yF9HzizotO9tiPLkfoRp/z1
YqY+nG5ahWLxaQsGUvu3xef5+MhdksC85Ann4CF1Epd9yjcQ2QvilE3FYpiBNZcK0K9MR23JijUt
BxbaaLM31iGI8GUR7INhgDtJc0Kr0Roo3ig3j/sSbCJZKw3XBkdBexgofxrZfB9mdNwK9z2m2oJj
3Zq2N29egqH3FgF9UlelKl5vOk2xAka/tOObfDZ+SK5C++Q8n6eO0CfoanpbKvNYaLUmxq4GxUil
IcjYLoJnNks+2hekhL6lX5gmN6pNaQnLdrKuX/UVCBpEsvMK2wK9bNF6OxAa8F0oLI2VPp8ViBqj
pNCRKTffig0rk1yonsWJPzy38EUvbW83lywip4qGPVoUzB0ZDGT8aQCtb2whcttTcq88UyCoSue7
mM1Nl+GluWjqMh8KLG/gK2GBjPCj8F2yMfigIC8qLkCPAfHA8pQZoh+OlJkJ8Nsufo2f6WeofPj0
ffpAhzE9Kvm+KLyY9moEqgQYsVhpEHKwSpLk13MLT+6bOLxzXXCcGuOCDNk/Q/yfazRugdhvidcn
lakcXaDzscN4BGiN1Ybc2u7B1cQQ/1us5SC+pEpbcy2O2hx9h04m63sb98Cev6/OZmQAA/fY0f8a
zWUbhgTzGs2+8OlvpIE/GOqgGzcACAyw4G7hRN+cHEbL3UaXUCMceMX0gXJj/ziEhu9ecVpAHeIK
aw2SdUYhj8+weVo/RU97fAJK5PhU7im26USHINpiqRsv3LfDMZCTCOToF2d6ZvcfNJYanrY4mP1/
LxhL5C6+Vhntqbs3kbDxx+IoBQVxU7/0zrJqdxxTi5XxtM8vBinASSbXaDOc1TgN2lLTaTzlWLOR
7V7+5ycg6SrzyjM2aIZPoWpwrG/UECoO/j5EuQbKtgSkGzZbSDOtxRj4uCK6Hm2jGhKkTgeLpWue
OvVUY0+GyGRg4oCBaE4/juKXUp0YoweDwbOpbasOiwY42AJK5kxhAf5knMZymfw+1tzB0GbDO0PR
XoIGfUuUWlemrISr2EyZFz/baftjfNI+/v4b4b198F633RLnXlEk4jnj/AQ9nFmIIjOJJ8IGKdp0
3un94ownXgeSYnYpLu1xD8CaWJUFTNhgJ1TK/Fjzc+acyk4YKbzXD5yCSTmItao6v2rPJzPcU44U
mqVpwWrvl5Sdnc1/Fk5gBvqJhMqtMshBWLt2jCuNRV7z9AR7JUlDkaTv0GP7UcIIDMjdOBwRtJl4
YY/SyWkTBWAzI7VDSgXzIbksxltAbtmCPp5WGw35rcHXaPhm1WLbkAl6DeEigY4ju+l+NLHmWf2/
mMMydYKn7qTDp8VSa/1HA5lQ3rL/v7Rff6euUypY/M91V7V9mWLj2SMWNxDRjtuqrdeaq+1jJaDp
7ibBnoyZjB+AJsLKAR31Q0FSxIMPa9v70hl+WUlrZkij3XzKM2hhmTorK2XoQcXAQxh0abeayXls
49Rt8PVO7jRHdqnKdi775QhgUxYTGo2xo96fe4CvDkYIGgg3W5l4QTdgaNaG1Cud3E7H/NCZdVKA
jVLdRQj0V5Bb4DbDSQNUdGJJYwrCrZlxx2gVvpsLZ8UyofE7K9VPwaKHaiPNPOj3K0qsuyUxOYMg
uqMBhqPsZYPla0JAkHoo4ynT2/fwY/emwxr+Pbj2Gmopq+xgdUe2B6/eaNRolYALUrnDMNpb02VW
2D5tmJ4z+64W4gyQXLWfD8RiIgscvUtVAQG2vJGBwfYagjp3Dn0uz/o4V5DVDZy5bU1hfuM27YN8
HN1E2QDlqWTKDhZJYseHI58mLl8HwoIwgGBfgIDDNZIECLZtnDJMFcY7qFMoFS2OvozJ2SLS7eJV
BYksF6VjkF562EnHD025kvQhNvABzZxqfF+dD2QV7TFeo70sYoK/PoHWUXNT1fYmgj4/012Zf6dW
RZ0xOqnuIyn+tmqSng+/vdTpZ2s3GrzTcP4eh+6Tivy2iFm/RA1TwovGW1i35muS6xw6ttDZSBwI
PIrNP3YAvFXmEjw9UONtebpVwken0xReIT1LVrSm6zj7wV7xYHdFHjSpCYrDop6E+K31x3v5IQ/X
Jp9u1oH0liZJ+hBlhVQHvmdaD8xBlbPPwrpdzP/JbfKFsKeE4GoC2HNbFiU7cHZRTUOLivVo6wf6
KMfy+NK24MDVjoZwc/uY+ZU4QRTC5CdgIEVkOqehk320w3Vl/InK0GcLZ2RH8m4q2Por5/nDv8l7
PHl4CUEpxZUlz3PM4OzZKLsTPp4bBnxGDlxpAj/2vTW/0iGHRLJnX8uen33d7Q/vvwUnaQ8hF65r
YBZEFx5nOYc2hL1A2KJJIlWkfvxiXrLfMcDLst8QwMi970Mn5WFN7seHRkcpxZSWqHAphcgsu+pj
+rIh7Xbho1Dkip4AiFDC0B1Mu2ZqHVSU/vd1XlW1TwNeWPipnb1hHTB4QhY77CTNq1ckjopXbK55
QJpKn5xGqisVKCyD8+h/Dre55Qc68/NdhIojiz0dQdTMOzAwBcCSqChTh2q4LW5QJ4sv6rY3358K
898KigahpafsFXlHp8nTKxypFskq4AtL3grZGAaRRweoqA8xuyxD4o3SdKI0lWH6e3oWEg0vGc8G
EbtpcQj8upkJz9ewmurhsLnlf9u0ixF760oYeQdce3jEB2mloguhG2Qhj9wxkzNNfnW9DN2RkhJ+
npnq2RNNH99JieHahBeX+Pm2vvzIaFvSvda7ECCuk+hjRL3Zpeih5NqIro8rBf1ewa7qZ0Q6EUzL
3NdGr9OQEaHj4B9lAl41A1pl9jyIU62XIYm1vSgD9XjKle9jmwDSgrnk7rpmTibb18K35NiGgk3+
LSrbgMvJQGvAGTFd6RkgXqbsLU/wDJQ6FDdjDbOWDYX05QV3Q1zzc9y/ksLTHE6/hM4zZgJW/j7q
p6K9ENjJoRmWYxg3+P41SrWo5br5QnLZbehV/jMZdROo0mqw57Ba8ga8RO9+eGjzQO1a5MNTyld5
7gHnyDyMBKZplylcv+1fDkPjKrsB2Ujl5Tbi9w89CKqDesxVPxOuBEQMGj/Oik+gRxL0s/GHTiKy
XRZS5j5enfHSRMKmp4zc1Sw6DQG6gsxps8mmFVK7oR8pPtaEU9GGx5a1j8tBGFw8gAFj1gVPF8bp
Xui4rrAzqI0TI9ZEc8aYvs0vgmLX7E+111wnkJwc1Oo/SDPOifgPTbB3iWH03o+u7sJVgYlucXVM
U9dlf9xbnEYCmBNPdAsSd9HJ+jvdAJhdacMPqWxJdzoKrQijyNaIEEpnCK94Q63LF09c/l/bWXHX
oyt838veCQ2i4c+ME5C0V5KsC6ot8RV8hE3OTpBj/7wi27RKNlxsIhdwTApNSVAl/o6wtCRBAEec
IXm+E/l/NP2IgFqsCNiPcJTF+OfbwruwTEJ4TFtWt70eE1cSpxPy1E+mHbv97A89HqGGmYFpyZ38
/fBxZI3FAG1jP2qkvYQoL3AJoZWvgr3j6rLC0agShrce05mOt7wLuhy8QDQnjyUAuOrl18xvxBUd
JEAolRwTJ4BLxd/v5FO0TQbRopA9rTUjYpPA9FVaRcUnLI6Ty+eqc8Bk6q7/Vz+zO36rXDhT+j4g
9h9dN7JIbp0GOdf/gfJZqiuI5OYZjMYyi+UVl3m5usCf0hAHmS+juMK4667lXo++xYG1H6+/yEem
txCWSYmhj+vB76oSgMwxjtBKKVy8WkmSj0EwT+XTLUuZtYhvh8KBBWMBruIVIZWnswB1xe7F+JPt
fxdhxVa+iZQGhung5jUjPAHfguX0ZpTEAj+sNVfKnJ9PZy+eGRpDdLh8Du6XBDRxDL2VxGlRbaqE
d53AYRAI0E++ktvmYYDjk5iTsz0kUkdOeUchpR+nbAxtwNNr9dQVzG9qpLzdLAlJPygcxzvAbcEr
43jL+8TO75kcx1boQvI0OIIMnOPtdsWW7Whes1OzviCybrzwjIltbGmaM3glppOx9Yg4pVfDBpm8
MXTY81dZAiuBJKue6QVGYTlNMNZhdM58uHN5frZ7FZXR1KMuDhfcH3bWSX4GFF7I/BMYFEcfzwtB
8AmS8UpBRQi5haviLKkRaewRY1V4iO5HbG41LBb32tqVune5tnuRku17WY0YMqNG+YVg+P8uL6e2
1ZZSxVYXUVM1KTtaDqGX6YjMH25Wi+Dn7LyOniporn98twPCL4CVALeczDc8PfA94QeahN6IUiSW
t/rxwa72bXd6PCbI4XLcMTXhZVywNwU1IDGRmRhd6yNhPyvB1z/6l7xFJkhW5hdAzkX5WJrHRyMX
B1YaE6qnG9VXtW8IEY0cynq16r1uZGO0K+0a1Z5R9OlUGCdRS++f06xhJ9B4XoX/SQroF0jJHz6j
qqmieuOBWtDqcx94DvwHgnX3BnXXPHiLnmcwKBGcNv2BFJ5NYrq9+xUqfRXAxLIgnFoM5ML/3vPF
gAJGebHXevGdhEBZpHWYBWJqrtPlsu3nBFGj70yM0aEqi4zbuhC+9wMkNF4n0sIdnCNTwm+fujCd
L+gX4cGPvQpU13yxEBCmzYT5vD0hlSDJdBKp6zcpJEhkJ8Us/qpa6vg3QkKK0qWRorhM1QOjcQTI
vK2TGaAF4ONAUljGpVXNNBoEmG7NJjkxH3FXL60Q8hivrYHzF5sHydk0sG5N/q+ualywByhOmrvj
xepaONEaq9SjFat5H4GRh+jqPEiLOaRcpxGx8goncAvxgkI/pYwDBA5Gd2U2OLAG/V5iMXeRxZQY
HbHVxjWGMj21tsRJ5msZhw+oEtbam/eckMtMnDETRQk3JAJsLR151lKeUu/d4AdNV/DPD28hJrDg
lG2TFeY6oT5G9neUr6j+S4yuQ8XhOQjar1FlWF01iXUfWdeuS4Hd6Seh/oa6L/nnnw1hUCSoX2e2
deoFvTWDIjMFm3WIoqO3naCl43YtOErOB1YnsGmDTAk/OLG21qk5wr6KcyooDbSH/oRrm/GHlnbI
h19yPx/F3xjvQrZL6+0lySRAqS66Ia8j9FFxzaacmSDbtADw7OybDWLFO5J5wz3sw3JIXkvQo2C3
K9ydBS4S3yzNJbmFZ1aR7amw0DequXIgIUT0Xzh0e40wf7jU5xJO6J38y9NttAmPEvq104qsdF0h
jD22KlPuBV18gDTyTuy11GpJOJMwA8x0A+YVK+VghNDyqe+4sRUOHml9lxeZO1ErYmZR2DzjTr0n
m7nNBoscsK6DIzf4KMB5VOh2VCC+JZZTX7csTfBOU7VBRXnem6+vvVybup3tFXiXvFH0F2KDgepD
qtOyl53IbqedHtBgK9zsF+BrZyOC0mIZc64rBDyKY1m4FfJF2nSF5CASyHuinly7J33ghlaMkcy9
XKfdn5sO5hAnoFANahPWw3xDQKt6kF7yORcOKk45Asfv9g1bnSfxXQ8aQLSW83y/S1ZyTBb38AXq
MVi1lHMEZzW8R6ZXKxS1gPCwWEXRIfgX18yafC1NnguvEtRz5B1vPMNFjUGOkDrGzIlV5HVAODax
VmECnjtATAsLs5VSp2YCkQ8wTTqIjcOHVx3kn/ZPn/rHngwaACRXFM/QnlgHidCVk4/91vUJXAIC
nXDjxrGJHlJ8Qd9xYPz0F/p6u6VfMHgXhUQGvO07NAD5rp8NYClDq5N2IOfZXPj4llLE3zpTHwAh
5aosota7o8+Tf/CeyU1l4t9+mPojiCqBdFP70wwRYlhftBJODzaiA4/clj87jBH77kaV4F0MtLvy
/HIhVCqPeCZzDpGVOuDeBDl4GN8C0PGO3jajQv4h3NdOFS6rM7tfm0Gvve/Akr3RlkZZf0J/tu0F
0uMh2NnWOPWnbRLL95/NLSEaO1FbF5N+T6xMtyMfuVN0z3UwZdjGiARQw80O3AXTPGA5QtR15GgE
EyCcdj0g/DXwNgO0ECaN7lkhUT3sRv9MtTSOxVMoaWGmMgogA5ohbciFirq2Pz2K2sfGoqTQVD3a
wBTTtj3ApFrdWjExFbhr5w03dPrCNJjJYn9kkqLsrEM01h+DyfHQMJfltlQTvEqyilHacW+FdwUZ
x7OnhfH8UF9s4Odk6dr4sjbODmHYZqy8bEsw3lXQ4owoDNtv73nhR5VCROSw5lbgFhhq88h9SuP/
b5hBWboa0rpMX8RX5bQ9sG2zyQwLH4S4j0ADv8DOtNVSINltLsNzPO6pxP9/9kWnUZYXpkOfk9Dr
nrmf++HFBqod4oqb7xMT0RzcUx1X77WQG37EN6hafUZ8M2GtwpJth7GJLzRQVjZy3rt46D7JuZ2Q
94fAIDa5DziIrMUrJcO4XxAF/E2U0iiCgHSZBnB4Mwrvy/NpQOPZznWSyyYaNvgn0A3sRsrtmBaL
KVrVjRqpf9yKCR38rQtirHttPIhzIIiKaWwTkVRFn5uyH+mIgPIGsMHY/XbbWn0fMUqFsKgRcSeD
ba4HtpeQTgAXhiBkdraN+8AyMyYvvsLhVW2fTl3poo2E/25GOkeVNW6FmBwM5raZ7jpb8HBjFpjL
5OIYJJtZCinzWncuKCp0Rtgx2livY74T4XMqKeeLt2A5EbKwVT2tnqhpEoMaOpcbL0v79CaLNYEj
EFHoB2Nign+W2nOgweoeJOqjHKs2UG39x2d185m+1VU9Vpfo8COJt6nC9mUj7vs5qMo6sc5moqdt
awpUvCc2kCKgWIKWZ+E7UWx9PM7+B6uACwVfZ8pqB2kNAE24ZpRlbvEAMoil9f24XBZXCS10GgQO
sEPkVjZTbG8fWvamEKbyuH8acalkx9SeESnSdjHrzKPghoNonK1jcx1nArzCxIjrtKVW4J0BAs5/
w95MNHHxL/X373U955UL4SywsmWQZKb+5BZk5dkV8iKUftq+B4aJuZ7lfQ0jetbCwTQYihnqf1Fw
X2aUAHQ3XITnC0B71G81cqNWuqzg+EGfkDcLDfnl8Ms1Lw8ehZATeIKtGFC1uvQHXVsUdVX1YitD
0P6Ac7R5GdrX0El+cCPWafuWfl+Q5wfi15mMS02BbuLEnJ4nSDWOXrxbEB9NChSeW9AuTaomB3Q6
JEj7xrtrzosWyNOwIC22jJ/wIQv9Mrb/8DWg9m2ugloKAcevIqb35Q93Rr19UkvT4YJTnuRAE3f5
GAQp0Y1+0LjyaV3uBaIK6GYwBIO0SQcoLCHEiPk7Kj8XlJkOhqoMSnva+2u04/p1I36BfVjaX2QI
J38mmPnRf5m3VN2KWwT80UGj6CD9BJCb3MT5TAWw0D26w+5Qi0/5ChM8OjoEDa4oyjgVZ9bNY0+Q
3sW879LFk/RHgD+aAC0uBevQW47KIcF/ofrFBzQbAbHMPkefNubEfnjPl6hAUFZhtC48YmXZliKS
pYo3g6lVYgCQtpgBgcN+eu9dtIH76HErD37aJnemR3QvkLZtucX+EjVBoUZ26Bp94tlJ3JwA1sgr
i3mcU/8s2jDCV9mWzNPngeDmZ7FKpXOmxJVbnFMEX8CwFpHlyGSjkQhiK8cINXIIjNOJzurPxFzy
+o2lrKpH+OQAGy/h1FKwd1yfTCFtqjSBpQc6gVLn8NG+FN/l9foPUDlvJO1o6dso8gqlAr4u8KiD
+TuqlAP+9K0BsGPfgRnX4XhT3ur4nUtILA3MkMo/FPnTTHUYubXyCF3wgyMv7MypReUfUkkGwpqH
EmMGsa6WcRJvf4wgxg5O1Ew/J6AvcE/jykvJfV1A39W0qQ+kLCDprgJrFOAyxWg/g7aXvRqhH+ps
zJNSh9bz4zZ89H1x3MLVNLA3ni4FjEkUmKVZzKTpm/KQUcDxpMmKNaoTtWJXOXoLynT+jLyjxETx
c1BUfc29ea+BlYgnFa8+k/Xi2PGgjRRCmMAad6FCenq+nr5U76LKWMZ8AJHfdA8QB+1Wfliw44mH
O+xBG6UuRD6vAEogq48bj7obxFJryYHFzrWHHjmbeL8TnfkVOpji65ei1hpGDY0E5chb5ZqDjYdW
zHR/vqGtkosX1XCVCjbT47FVzdUHPq3mb5aJcKes8eis7152cm7UTRQvqxEIbCq3AwQUvTjoEQdQ
U1tUuDN++EKVA9LPyN/voF09U2Mamw1FwqB75g9oLsHLe3TQ4fizsKiFIq+qmNg6WcQEn9xbQb7K
y5l+s4ZIv0sUrKbKeCOnNH5I4a8q7OZO6KES611z/0UWyZcPBVxbV9j9DrybUN+mEh/qpevqC3C1
Wo4vX/JR8oBF9i4iT4Umtq/jCl4fZsZwn+DopHo3zbqZOE665a/O/hGAy18q1Ilc1Pnxi1GV2W5a
h1OSgILhSS43dBGftqsN+lB5fX7+bhyD9irBxf8BLXC9/0ELsZm1u+8a7gyQ5ocwhx4DqyECJDZ/
HH5TV66lLfnQpgaNKuksBU38Z8YVOkVgF+KCplTVgZ3vtF1o/UU4fMZ23FZDE4QJhiNwVE5wYJ0f
npz+dI8i4CUTjFT/9jeGKsA5SuzZUs/1WeV3wnOoqrApSmpoLLAPR24Rlqb87ZS/N7K7s0xTasfK
vRvHvLtm5oZ9VslixkAVvlrH4dxqtxTpLHu93qAqvKkIBbON256phydRBM8cQNHLanS3RI1beVXw
mWDX4lIIZEXvMtVv2Ym1R0Tb0ccRdImaiMzC1bPwJ5hNPuoXxVEyfvoAvTTfbJky/Na1G3iaUGlD
wfq0on+1+rgLs5mu0ZN0EQ2eKKow5eBO++enSQsCdsrrGIiqxtFwpfmjTeLp6N1exwM88RPH00Jc
nKQvR+I1zNOo7mzwNSerqBX99Ze/QjrC9C75wM9JHJ5Pl5lsuI+IFyT5NL3T5DaPp2Yox9jKRyHR
ZqoroZyaROcfj7AGI3Zl+qxRt++ckzQNOOQrMFmb6Br3NhqCruaDYVJy6k7YP4o/IySSUMxqE4tE
X353FdMm+qhCAzZN7WU2MdTntaHoXNwHIGEkv8Sb3e6Mc5JujZfcjj8tgpNJ3w2LX+EVldX2Gkof
oeYJqfv1dX14l8vEJw+voSh/K0wwCl/tYusSBbozvVECLn2Eehv4PTP7eq9t58Br7f4T0UG9yngI
wmVlhTrEDHXy2fZhSLLJR5xQS3WBOdX+VjbceMJMVo/7FLhF9XbEqTmwzqs5fe9MtTBU8Z7uyLtc
cjF0wJ785XFDkeWrpicqcmH10imt/NSyAF+2BER72f/ziwuwTRuP2LKytpYmgYz1M6ktUQRvGUoA
5rXZg16KRGZA6N1/oK1Vjr4ZUYcWioLbe6/whqmI4K93wXjWHMNkdC2ifM+XeRKGiAa4au0op+nt
3T0Kc5Tb2HUztnN2CaZAAYxiEiHU3aeGdWlFGKmKZ/Zj/xqwz2S1FY0z3+CFzzqpaEGL3RCD47D6
CcfsEiRY/DwB5RJbJHcRj64dj+GeKsk3x9Wa+vVuyPIZUKVP4Ml5Ji2HBKOGcv1rT37gkUTFZCLM
zaizFPoG5Z8NXEKnpwHC5la7RaQ2GtSvF4kvxTGiqM9Lol7tSoMeRsr6UUeY3OVx1JjGqFGm4ye9
D9sfW59G896SuKPtEIy4rs+FSReTnLod2cx7mhuEB9zy/hVRKyr5BQt2+WsN3/dBy8++GEIAzuX9
HtSPGVjSRlo3Qqu7FmE0mUD1InSCpQoGBBH57k52e+MqlEPUnhV78ZfsdEqAK7cRCNC0ZZVqXTOq
LaQwgixr09DZ3ZxspxwWp4mAkS4YmZ2FXCPMI5q7wm6d0ADa4qjT/5wMkzSp8kt0g3YY20XjfMbR
PWaNsLsKo0wSGeL6cgM4gR8sWBYIG+ybsy1ymTWyH2qNcaTloWtiLJN/nTKPXybs6GxBSN8/99wM
WMvWKQAmyTlWtZ43KxMVqyK1YtEsJYKV9l2cssOx/2QpqHQ0VIJqia3Q5/8Bt3CgpltDcNOSZu6y
8vWRbvvtQVKTrdg445KRpH2FzsBbBZISXAZ6x6SQcBDDizUtSC7+slPcVt1Pc05tPTTqXG2RK0iV
YQpvruZd4PgzICH/2sJoG1zq1F9RCfHBc6ntBNpDkjpOmqG4RKdf3qmRTdPA6urq2hKqin73g+fG
4Uldy+U8iW4UeGK8EPntOoOyZtbf4xqATXZo96S8usinexpgoc2IWiDFiDYIvo1pHpl0YISsQzMl
ZfTeiOpqRCx7kUWE9aR1xhN3kj4yqH7T4DZOioMtZOLhUZ5cdU8Mu/CVgQWP+U5kOoa1z/YZR5th
gt4GEO2f6GGpmZQ+zKOa7adQawUBwHA+ikEl1BQKWYDC01+ofWGVM4xFHJ/SnHMQ/2ElY2dbhewY
hi7nb3Sp2zCJgKDzSu28mcMwyydz2gI7VvPxJmbqFG++SOLZyybafDFTcrgSusEMFnNiTZbCaAs1
PO1dv3hBTi+vIpxANU3Sfg4JOghGhao/vFxe+4XvK4ezWX8oe8uFiioTpyGYqpXFUxQUM4nvZGi4
OorKtLwC11EA/vxpUPdTdMvmNXI0s+RE/UqHOpWWs12rvjad+BTbNjLjAGV41bM80d1DGlgzQzz7
SyR8ttMSPUFRGV6i+3ms95l/CDHrsNDypo0ky4CV/5H8bWNhVi3ZM5+K7cqLfzkdLN+/7tzgiesO
PyMZnBEDLNJq26SGNzKtHic7C4MuR6lK217d1onecMjspiyjmgn23iCWi75wuJVSfLAFCfF+HT1Q
DSlkH75CLC15YnDNRopeUOn+VuhfMwBlMfVIqCHUuSwHdZIcIc/rC4fqkvbK72V9AYCjTfQeq/+k
eDqY3SPWGftsiRzg+o4KlincHiNh3SMosOFGmbjQlhE1CqvRvIcrWMZ9lOTzApKoCjagmICzvZzJ
OKQy3fFUV/DdB5GbYobfIKjmbtKW18WVOBbvda/1mdt8esk30ZM1pffYyAC7Syc5D48hG+FryaLZ
4W9eC5gW7IZFBzuPdw1o6KLEr81ko9x1Og1tUyYiy6fkt8FD0SHdgJE700yFsrdo6tffTE325wju
jMRR0aja8Y0VljGe0bcfIwNusuYntnf7VEseWpE7tdQQxIWk9UDsOIE6SJX+lh4mksB7E0I/L7l7
4rxoVkBtOP5zQ25kgA3Vum5AAe+XyPfZ6GFWJioOId72GK7JRnl1Y+6GJ7uD0+hwELhMJvvSGDwI
pDazPFeXHXQwOUmuYd+D4705O4fGYQKB4Wlb0dKpF0EyrqwlzqwSYaBg/XqwRq6jZPLzc4Us5vIN
wXkXvLb2F9etOoINhs0UKKax7Qp5dSQB/Bj4h6uZ6wUEF77RfR5H2zEv6kGHmh9xPFkq4dbdHu+J
RMX7AfIpJGOBCzMHkrDXMfFGsUma8/T7se06cZxjSo0XwmvNbvUOg1sJudjitqgN8Rmi2l0UY9IJ
8qQyLGKcWQ0+MZPfrjgHqOgjEQ3ryHc6tXHxN8t/sH6DM3nvKWOKTQ/5KUOScoGQmnEOOwkgi500
JowuFw5ZeAfoy0etF/tXqyYfIeUA1GHCHRPrFLtlAvaWtuQvlNp246+SRP1FNO8xOH55wevry8of
dl+ZHMxGyupRJPKFRCXuZ72qQtj6HEk3b+6mvN7HjGcYEgjpWy6wDG2BzuVEbDSzr2lV4UEI8gtQ
ih8Ew+pcS4KWcHA6rB1GGPV/4P6o3CeKfvmAqJW1ETLbWXre9/2CnGybCb69Dyeam/aIX+7E+SfI
wmsgPsnPjkhbzc6kN0zVkJjmpuDlxmw4SLOJ2Fhi6GpN+55S53nMVt6YFNYeOAj1vS2XIXqJG2yr
QM/pZOZxphaQv5x5iJjLPWPJr8a29WFfFeyGsyhshjTmolIeW88RKcfoGP6+t0ka5OtbAF7NWFtN
Tng1nnWZxzmyaUOGKRVR5w2ZXljs5nwjcguF0KfDRpZRyJrq8tmUVw408MD58f/87MSBmbsr9wHp
dU8EiOVpGI3Dd+zPAuMienTx+YptupL9Lp1qQql65UZrxw5izhH2n4xkT9/GyRTnqBwZFDJamP10
loGQgQeDBKoz4hMyD8oM4uk5z/LjKxhibECm+X3RmaVWRHQwAYpyz0beXy7HvLjclhhiJV90Li9T
FH4xNGyWMB0LZUB/Rrmfu/7xwSXEHppx9Yt3//LtXyIB/Tp/RO6vnPlHCYwEqocmUnYPtBPrnPCo
bPk9Vey1Nteu/hNRwRZ/j88qaXa1SpXXmrsL16mYKYNw2uR9PiENOHQj2gW03oohPAIVVm9UUrBm
or3jnG9Sbd1T8FA2hiJ0YofKS4bY5kuybZ+8K2bhoSUFM2iUM/gtEe9WX+BgkskpET/fwHGUiaVY
dLxhD4MSxpAwNtLm2JTx8dHXE7EWG1WydzqwlWCfTD5Y/LiT2P/T51o0s240x5VI2EcjaD7LKDx1
j7B+OTHuhTFPdmuHMK6Nowj1qTmR8kCcYQDyYfrvcVmi0TNpquiz5AoXTShCavqIxnEXGudpasVg
cm11PTL+6iJCKtFpkDYRAEJZr9q9uKWKw0Z/QEsChO0EjZy+RlRq5w5rLcALOVpViSg01JF4jVY7
7rtIeL/Doz+MjOO5UxXsF4dGafP5mcv26GVn/7FOoa2bUauZGf1akJa5lNREiBTZx9MysEVSy2NU
VEZ8UKh3B8Zui5O+HYAUg53NoRoNjVPJ3tLnTgOnpyfnDM7Lm+309O8Y+FB0W+2cF8w8pl7PL0wO
35rrBRsts3Y+U9JX0y4/U50Bhh2TOrtnzbgmnQ/RSL0MF/UZ7wjkEJjxSLT7KXRi6bKhktsH0aka
/3iE5NNc5AzmJeFYdXB1W4UKlFl3WVEqQjWV4YUHCfvd88L7FMl6r0ZDnruDA2LVK5ink3E6V1eL
iTrE7QhKaAYbtrG/7I+J663lGqjOODM6PC0LEXLUy2gjMtm3HrwRuqU2qdYSGTNxq8DOvIgFlm1c
VSpgM/hL6pfoxN6MPWVSgEwiGW3zbmRVvAWmIvp6Gs35CXYqGWMujZYreTgRHLwxN3efatWj0Az7
7JM3r4EGLgJd7mW884E3y5bYQSP8w+ULRjFmVCMiJWQ8CGOpVRMZhXl+Ha/j7hpJzHbclq/CRCs6
ImphrJ3QTHJLBhhcIqbx/nFuRkdVhu88mRZaaiC/2XiRGCVZTTNS00n0xecHuBRzMjSTnD2sbFoT
xVzoMGImljJjp/NWZpmVBWaRkNW/zb8Nh3Rb22YPKATWBmujCx22Y073Xk7g++bx/cDgnrYSZFUm
duNajSdlo89rFiSaJ+2IDiPmsQGGWVgIkpYQNFhjunfSAWaU4zFHAES49Ijb8P4V+Zy4zMpPELDD
lnKNuMBjgR0CUAV3a0yF9m5ziYSjZADh/Edy1gMLMik8jw1OOmXU6ftgHEBmOWx0alcl2YQuadwi
Aeu6usfIT16tnQErTjRSnmlOlKxKL7MGLhooJzPr6yoEWCLASXzNGEfY0jANjeLjbNUUMdPQJp+j
BWQ69587Qy3C0Q5bEi+T3uLpesqUUSP3F7wxB2C62+WbExI+X1Ia9NpwzM1qmJPvQvpjdqUAHtAV
iTThOVh7k9LZmxVGpbz3C7EuhgATqYaznui7ejbO00+0oAGvWmRrLtrHoTvIp8Nng8GFAF6Is+rl
W7z6AscRGITg62HHlNipP+b+7GyghFC9yd2gxjoBpd/YdFMiXvKAFXmkFYZdoegD9ZsT4Q5/1uuH
kRXaa29ohcaV6cXBqbJum27688LCz5DnEIbgC8pdvKTfQbmmpiNdMw7tYbPQL3BOhm2m6PT3CxaU
mOOkzamd1JH0/DrhzumuVZSaEFackySK/tghxEm9IzGhbBA9TPbte72rNvyxJ86yD+7x6Fe3qtbv
6qyxjHdOQs47JGkbSxqWipxKhS+brpT0YjKxDkk5NUPrEN6SSCNYKoU24YiLBlPzFQtmrTZYX9s3
71ZTATu4ZAN3f/XkT8PEOFMTu1lbhAr3iMOsWsjLK0qqUbDuRoHVC1Z59pCACOv/qS17WCPSO5KF
Dpbo+CSJNLUHgL9fm6SwLAnJ8E+yJBDUF1WGbufjqGNgNn+hg4asYufrfksUIPtnT5d4lUz+8rME
Zi4K90p0wyKRswxqn8jS5O8Usoi3g5+/4l7VHuY79O8T0Lfeo8zf3KeHZ/6WTbrzbMkBZiBuDIpF
8uJmdZbw4qx7fEvNRCEvuzb3U64xrIPiVP8yA9W6LKJCougQUtwcHNxp0jLH89nQSpw2fVbREwBG
yfdLq7rfCWRiLw3h0G/c+YacFqnWKZz0/0ZLyw8uBlngKlOeOP2VZwdd1U1y7Ihb1b9aASKX8J8x
h4zWl4c40kz+kxIxt61upmg/yAozfGU3b2GqDerHSB4z4W3KaJCZprWp2p501tZtt+KlwVykClbj
4AzzxxwjPX6TuGGi/kt3YtH+RFUVJpRKthLayDFkvkZ/iHdWrJeD7yTlXUDwgQUiksMCioY+xFbk
NM9gRQsJNHVX1dcbKO8fWr6QnkPz9m5EvVdm547LUYObnUMgDFnmmDzlJ8ow02+R5o0ceH/P0ioB
JzOk5sHGfLq1K4Xqrz2i/XApl7EbApW4gGwkzeWv01XxG8tYam0aq8Y0NgGTIAnrZfPlfBsVJYXA
Dv+4RlccXrVM90sqSVaiI95yxV7Y9PownuF2iRMp67jjyiaNql9EqYD50DVWvIEuhbvFK6U/BJmr
0D6cm9qmFtCTuWkeaENAfDH8vCzDvSdhONjTfBhzt5cr2G/kLTHtIyzf/qAyDgfKr8Z2iMt1atg2
ghg1KE5m2IlAM3OBuh9fs142WldAbFCECdo5yGWjT0c19aV4NWvupdqZPVYqPrtzgCijPpKSHE5H
2ZsCvBbt1vPAM7FR87b4e3CJK27YdnmqhjI/Avx6LsYdsVGzNFRGwqsUSVMFgGsKmqCh4jqSZj0z
ZdmXuqf9O3OGxqTWKSYSaY8nW9nF9oe9q/mea0QdBYYFHQblpvcVWPlyqe1WTc4M45Gw3QkhJpTx
fIedu3kJMFNmqiPaJ3pzo93u4obJfec4OVhuO5wZXTmVOK304QZVqWU8qj4l3/qEI8BwteeGi17K
kT2cCQAkgtMYwA5WJNtc3VJZ3x0ToEX3T6zqGsEG1CVZZELs8PXIGOveBH9lEqynxjYiC2dhm+nz
qBnuTR12ghVTTN/WqbiU4bsjAnPVux8Vd5njVTWl0k4pvGD8t0DZrLO8PNr/rwkN5GkxWIfYeSXA
1amGrhuu5vHZfQ8vSbcVJ1iLV1rkMhRcwKBQe5biANasjNkahtMA6q6O5AfJz8bdce95rl999xC8
Fl5bJcjEfADrBafijwar2BR0PekwaIyb4yS0iboLrRA+QwRkN2mhIUze8nWdzfqFTTUlPiewhU8R
Yq6npUHV7SwnEL8I2H1H8dTkYQtXFV7zoYYN3wUS05WU24pENJVzdRdDgkXUn4hgmQaTvGlBdko9
0XGgLc4I/3U8l6TmfYFq9YJfO7c6xbowKdvAZ7D0TaMj4xpaM5DxTbrMnVKDY5IYVhEqwuqPwlCj
NxfcGubiC9iLF+s5lCsD9gYRK0q7jEAs985DPY1k5ejFp0kbks0KLzjy7g77wuyWWjfnY2hg8abk
WO+lTtiGQpdAWeF3nlCvIpZa4LjDKJHzM/bcP/vqoRviQ6/4RS1NhD5ymsuvet21+NJk6SffgEid
0IEb4DF+VJB4LFKjFttw8iMUVoP8xga7qLWJBn71A8+zecKzpAl2qadqLpgMl1enNTb8T8G6iZ03
EO5MbjxnKX0eozbuGfs3xWQAqUh4qnkN3kgPR+VFrs5sBrW0HdNK5cY4O6b79kt8qICluruBw5mX
/OLQS6ndXRrIH5dokbwVRsNSGE32RKJh5u8YQFU/5MS4YUWZqg/Dl5E3gvyH8V1dmWDjwdIdSlMt
7VBKB/S0bfIw5ZyOxy4k8FNo7mac4dionSEb10MiW8nHNN5PrUWrnIIzU0/8f1uahXBatWlIe6CM
w9ar6l8HKER5SnZpZlpT0Wt8ZzyyKtqCgf/5Sob1DkgaWG6xLm8jqGWMOPc0SaRrK9wqAqpoZqd6
qsG+KltYozg8GBHnLLhg5YMzuZB8mx94bAEpddq6EbpjSrORrbw3M1PMKwqtSTc/6Ri6eSQgJ/Lr
8Osv30zdXZsONrCWOt+/08BmdRd9pk2rWyjTW/ht0evox9aUSFgR2YddLdvOOfpt6mngXQjCxGFq
+OYOCT8P2y7ODB1OM9CL0jGXMeUAs7vfE/wxI/ZPpz8cQnYBnynvEqgQcAXBCGjdf9sIQdAsAvIb
5I2ASF2XTGmFClBEGRpYssLMV6FtBacbTy2Lz5n+Og1qXVrNNu+s24ESTVvkD0VXaEAyNZUaMkWv
OkH0A4dfSfKP9xDpFGusfs0ITsaRPJxY4KfOYiY/D6sfmHpFB4Iyw+aAN4PY9HR6QRiJHvo6tWc4
VXHvC8nYAXZI2ZgjqUvATZ6QfdBO6EQV0vAiWuhOHEpu6NcvBqTg7bqIudZMypPu1gjBRDrENyX8
lTcG1LL6Nszgd47Ax8eGoNHI+G7JinGrePbRtw8uh2y+mGr8lNkhjj4CoMAIu+wF/3/4xR74UsJH
lJd6c1cTAmRPkRvyZ8BqCxkJ1OjqEjGTS3TZe+OYe8ATkS+WasOdr4E1BAFkc1LW9LzYVar3QRuw
3wyx9E4gd9hfpPqYH6fZJ0PKtb3beCQsXGAUgAk6xbIuANwfUPiBYVLuJYeK5oOKcr/7TlRLqpye
aPHNiCEfJwMCXNE4f/X/AQuaqLu6Ui1i/dPxguGLn4HKoFTv5eJPzm+cDRMMQ1inhlDPSPLi77rG
E7R5U4/UpuwAw/IDPqMiJLzlCQ/CaAyuXgecVLW2zbWiSVNZBXWPSorKhY9owEHmrdFHFd6gwBVi
f/vdgq8K1qCcffa+32Mk8IzOptLJE68jvTXpCKKiSTtzuIT5McJHP/ZDCHXDTWmvEP7TTb4fUQv4
qulyO/alMKXIxSQBdj31YWu1ETf/nR4dWlwb7wrn1u57ySYkj682WU7IMKVScL/n4BDYgmUF/u+A
zQyPddzfcl5ubpul6eadwYninMTEM/eJ2meZBRjDteoNYVl1vKbe0+qZm0VDegPWrDyKvMR117x8
CpxJQmi5n2VF5Es0sn9odzUAm51vuKmA4OCP4kAQN9RGohbXRq2VYFpqPkf4ZxZpiyX2raRvtYTs
lmnkQIbDQAV6hKe2HEURr1j3K3lFYDUFALnz59Znfjj6IKA8N+K+dmq9ldAjdDnH7InLPV3gPZO2
HNNnV64xe7HGCfPQ8jfeIWrmisDULHzcl9dnoUs5Nwjr3T+sT5Jcdy7LCTMAglOEK2Ow1VfuUaR+
s/rjTMNbBxIQZsk8LH5u3qIfC5pwuCz7qx5x4u2P0FTaaULK53Gm3vcL0ftK+1RERkAAykGKGvxt
1AiI6vjTEqf8dhP3zLcS8Uhfv84edHb4DPHkDkG6OAsQ3d4hMAZmZVVG4MKWgD/uOjY8m2iEfzzP
1H9/3RTye0z3+zGP10rseZI3xr2zdVIRMlUVXYncDQuvuQb1coMm8WUt8z8O7I4ppoJ01jST08/m
yq2mCEKWmQwNoSwHHnnlOJa8utKVEV4vI7gAtAtd7MFWGJNp1e5ogMSutdkVK/dCUrdpjabXMQPQ
KxpZCiQtDLqFVtv4DK0w2Ei/RDm3Hdn9Y5Z+3f0eOsIRm80lhcrW/Vaz3jR8aCtMpaFsldPuu3gv
3Tb9Gb1SIwbDZBPbLdp6o6T6Z8bJNMW14+M35pjnARv6/J/cr3bQZa6TdqgSxc2xIowa1MEPHTFQ
8lWtOqGf5h7suDMEF9+cORmrX0NjMICNQntB+LQ4G3o/2fil7y2ajqyYZ3y83UhRjdE4ZLgduDzR
1xtaPnmUt7uay7Knlney5JySLLuctCknN0MHM7202ch1wghjDLDHsBkE82JkplekJoVEZfmcrNqD
2S1e3L8nOV/RiU+QWsKMj0VlNBP65J/glVKbOFM+S6jn1dV8bxFORHrvw1++vkFzM5yg832Jpvbv
xquzw4KzCu9UCpAyvioO9VF9Hw5CBztoHpy4NDpBxk65VRofg8DHsfw63d56WVMsIt0q4hlW2i4m
PXfjHPrNY+EYyQrhaa3inAcgiSh1YrLrz/BFVhjoIBsIsenockyl49forrzpUwKn2/NV7mxfd4SH
LfRv7IG991fEji+BGMh34zCLCGCOnD7GtVY3HgVOTYrkJP6Tw8SsvNPCt48AS4v916yjEleEo0bA
j9o55XzLuyTXnnaDZ7LENGP4Es2DxXidiZD74rlrYtAReR5tq8WKb/a+Z8K9UB0L7jpoBpvj8w4X
7x76VH8ZLmBMrQwBh8HWTgB/NQFozPJfue0HnSsbMY7xyFkaPKq4MyTpGWSdWTWxG+Pi7z9hp1cU
aQ0D+2UxPvEUbYivwHyOAyB1k+rnTdVjA0BEBCDZF+g8oGAnnfpzV8qlRnJjBvU8N2jK8fN749O8
+basSUAjEt70HmzLsW0BZdT5ZOmDPl0YlL/JvnRVvoxQA2VD2u8jq7ny28ArO37l3UTvb2G67ds6
MBfTtP5tOEkgx2JLodtbVfDfSt4uloh8HlVthTSFPkCrrSyMh3c7koJMzVFuBdR08ykkVRSRulsB
4mYm3TalewQs2Nci7trs6MOIuP9t3tKZbtU0gxAGYBz9vpfhp6Cw+2Sp41ow8cbNgfiXuZl/yoJM
1hfSGiyT40IAkX7KkYzRR0U8KovUTA+EkXf0LDkUSk7cajhFwb6auq3IcNI76zL0JrcFnTanuGHF
MBNJ7vZxuxrr5Rt3di0ZD3PalVgg5nR3rtQX7Er7CRuPvPB7ytxgGsHWEHOgW0A9y7R01I3cPRuo
3TQ93TEHCnxUyrHkphPi9ej/8rtLdR2mY0wDFNEOhmtMJ+SWCK1sIXH+QByAY5gQSpE9AXa/UaEG
1kA+OTWGAzGac7rGQbFXbEltvVwKypLXW0iISse7bTc5xr1M0gciIDX12/imewxZDf0cn6iCq5+Q
BqVHfbWhW2an2g7ZtekKOPaQpozeRKNJg7kZlVEwgNu2b7X7qeqjfm6WBquJdqfCWpBGy02NMsP0
a4612ni3W2crVTF6qtuRAlup4GbIZVg1DaSAfJSRfdW4pFhOk6V4Hcn0atAImFosqO6ZgMyfW74q
LSlZ/ka7TL2i0qvbLQqQaky60IkUfEKuQTDMGekbIWkY8rkrijqxqF51LLwIS0aSWRAZ6T/4QZST
GvXCCU84pcxIJgsgzqL15fH+ZaDDIkTf6rW0ISuBaxWZTn9PIqU9AzfSEDIfX0rT6AWrvuone1RL
t6JNTdy2xgk5nv2ZZyM57vstTE22RE2PjhBiEs/K5tzOOFgpcVzcf/Mu+zMMp7qLkFG7nLqJ1l2l
LIbeXtKw/cQAIQm4hedbFpxSzgPT7h6DyK3ANb+FxqXWHBidSM5Zd/ZRuaPCFUjREpWTL+L+UDTl
cCl1oP+cW9aiKhXSezmWMpT0W+9Jp1+umS+aBnZ/Eoymwq+vPukjr0q9/k9N9CFZHC8SwrOvnmpD
7HrnHkqGjSkAxJlRfYOrNolxkEippYVLjmN08ETfgqCc2Dwur9gdHK+KoORabLWCF23Ise38nfjC
+upZW4ezcKBlAvZlBDuVxdx5r0kqE21Q7xt8t0NzOXlI5N9GuDq2lAYF7NZmcIUfkjSYoQV2kT6T
4w91oSfyFPR7+Y7lj0dVKAUJ8yaJy4/A9i1Jw8gn14eeQlFdH2H3a4ZFjJ1CI/Qus3brFVrU3NYe
QKhnXQhUnke+qntqqhgfUMWx26WRsLGwDNYVKJjETpyEqt7MzkhZUNBrN4+EuZ6cTd1KzcpK7rW3
+FxBbJX+3P4V9QMRucIfHhsQbaxJCvrOPn/jyKak1ZBNKvTKyLL3c4KK+ZTbeVMgZA1XNf91FN4p
+97O2+9p+Da4gbl7aUjsyat7Iji+ppaJpRDnRf6WhzsDxIE0PtgjOrqTACOrvLqlFoKTwTARg8uz
XrDuE7LNTciadSkJa8Ynlwry6MUOqYrPMaJs//HKFwreu/iIRzqHsyNurDg6gCvr/zVfO3w3D8Ge
4yzmx3FFvK0q/96lDrQQ/WWnEUwFdkBSZBdGx6s5A9Jr4E+eOfEelQTWSSuoqNTxANHgwFQ5xv5o
gG3ZUdBNGWftquIeu3E1hrVhikKKp+/s76euTTbH7b+tEUKOpCI6VJAoU0Y9b3GyJGDdW3i4dbDq
LUjH8yLbeaqzlB7/WbR3g0sBvjHVNsWG2YbnmvL2e3xIHjdzYKsMt6Ch6Se5kAtiLvph/a7Zx08C
zRuJ7uYfZEy2Rlyu+XRf5noQWr7k4j9Jv1o73b6qf6F28IU6dSeBqy2n3+1OcLiL8BLM0p+Zj2Kp
hpUZZB/Sf3k2prB17T3FMKou7Ably6a/yu6KpEKLsFFM+xZSM07It3Iym4RlAW0U2dlOcDE/kLkj
tMdgCdFpJ3hY5z+gk/BNZ83LdmpZBUlLSVOCFs158EvTImU2DqTwcklqLh+NnAv8dUaTEdsMDncf
q2MSv7TmDfMD0ZdKgcrwt5Mtx+IN0pbMshV3+UMfefhxZqu0PUicO0oaA68ONPOPXwS7Fpl+wTeW
w9zHoIxwsjzeqNEzYvNUVq+/XOSaxO0nfA4NFzMsN0ZVln4Xn6MkdPVh3jPLvyrXxRvm7mYFFsNk
sVqvSBmlCldV61tnJoPJIRRkgrwey6q3Clj8FNpkNtUUjriMyjRly/itoiMRed1OPfD9WLaw8jo/
mllr+aw4pociX3K9NUyzYevciojmvm6/yPe17UfgBt8C0UtUI6AWK124LWNXrV+RL/GpAGktkctR
+Y7PuHz7SFmsvHRnhYZzd09DEnbCqD0JgsUldXOEZ5/U0BLYwFOWxGuw/g3dfitC4mtcqvoZdzvL
dQLz8yZKhsrkYmrucn1sE/GLGreRjohw2oI8cqNl2EdyxhUizWhXP1r0pkOWUESZVbanyU7CDZR8
QLemWB++OlZ772Q/KPhxdmFvF8VG0c/p3sPuY5ZrgHzfZsdQcSt3Bj+q/0Nw1h2HJu/7yDNALTZh
pwWmrDG3ZJGmjaRJmVHr1B7fOX7gBrV+HCz6awGuN/KBDMba3ohX5epKvZtmlptW5MvBorF7UJyi
BDHCHKoxdvVfeA9dUcUdYGESqQB2E8n5pFVFKr45xX1DiuSouXzv8k+Gra/CYRjjBHwclHkwH7U5
390fP0g3eoP0xLrTSmQ0VeSlt7SgOcCkdvqp7EZZAoSAnZmoLCHabNmBs38j3Ze8x/81Ocv8ToX5
Ya6RjMYN99bL9UO+AARKN4XDqP/SqzWKobYSHULLqd4WrnkTPJ3fXkvzgVGqyvbtrmH7iXFbRshm
3Zj6d87Foosvkf6LkU4XFfeb9RKb2+94XhibN3YmxMlcjBgxjPKlEujn5IlM1qLRLvSKV4iBA2wj
ofwaH7UeSMrWw9q6IgY+vm95krAXfjC3iyGWAz7+GeIzomb9611/QYBEJInjFOl8Zkd/b2zMs/pk
FxOtC574CaDXuZQfakLYytCH+Ap6MupYVhNpOrW6NHeWcu2zjfwZVjthy8A550aGfbaUhcNnPk82
VYd4rbu+i713mfURJa9z6CDVRT7QwJcj0e9ugbbwTRLpXnS39ij8sKYasI/lC7S0h8Vq3m7Dk53F
TLoS47cjBLQ4yP8DRefauxTAkJnwWLQB6WRcQt7IExlFaANYDjcoB3CzDCg1pkm2s+W718FYYSkc
faJmjjHHxtx5WhOmEhMwNYlp0Rb4pmcM2Aqi94EJATTiX8+WGbrvqQHzvApCLeMM2ylrzA1ew6kD
x4kOo/RaLr1XCZeMkcjk8tn3tubcSEU3GNgpbNyUDZbA46jk/oWrvGhLLmAEOwrOQ76+e7hRPvDg
PLrHikX2gnd9xjQ5g0tlAgPpVbcUb782dw7Yw88w6DDkKxYWNugvHPz/7Mbq1Y6sD46gKYCahtw5
JVr6sCQnkdeZsqwDvfxzuoWTOmUJXSXd6s+DpTqSWeP87rJhTE8oPMEtgUh2p1ZzHZ7GxC5jg2uB
FAvKl4aHvtKX3AFwamUFK4lSggqZavyoQF33R5MVYF9snyMPES7eN/Ji38JQ/VSX42IGRQc03mHX
XhXbzo/wc+bm0ZZL13uE/fl0nP385LImyzVz4zNkjTXFpYuvQ3ngH/rR9YImPy7dZKqnNJXkqfuS
HAAljJqYA78Vg/TKnyEnYpQ4Ka4B4aJHBNsf06uEZXZpHKALPCMmbzyv7XBtKibbFbf42WyI7e6E
7th/zrEgPHA3p0unDDW++BJv1S+o/QiFS/W0Kp0Lu1YgKuvY0Kg48a007DeLVgJ0suSmLIE9imiu
JdQuSvVctFvm1qiuDdoGdOPO1oku6H47D26NI2ZQPyIxqmxAcvSe6EKQRW3ZawKoSUOt9IH2Vi7P
BB4uSifZ+UI5CKWNOpzul31x5+kcnJwJGH/ACDFMAMJDS5A6tYeOKHpWAvsU0x8IaPyb9viCpzNZ
PH3GtHcCm+/8C8c48MA2oeSQ9XXRDCsMkOYUP6W3KE2ALxueyNc6DZjcrE5d0vXk/ncn5zYWG95E
YxI4P3EHlpq4gNhgmeUGOKpRCQyVfsAhmcz5PzUfh8i5szbjccmNekqAoA2wAOu7yQGPjULHQNJf
ZtnFdoYUwS1gaKTwge5W8fgVKvOXwwYUW900NWt/Q4I6tOWrInkVtGLrDb9VSbQ1symXKj5b931X
GnaUXY6OOO+R/GbeNXiI2powRP/8Tt5Wi8xhWV1FMnTuBzGdZFfuqyeKuuxa9Ht6LDiPZZHpchg9
rJBhgz7NZaxjhXdqnmrhRit6FhG/iYph9TqBOk5pa5PUNRU45MpzikHBBKG+Pq/BekPcnI5p2+51
Vw7deXHm851c9D2u1DHXRTBvlDSsblNu3amLdbBwzjVplrb+aItpqp2gKzyOiwiSWWWT9Gxq3wQ1
tY1TlkFBs3upRfpUg2+RzuMI1hMh515qdQFHCH46UO4rC3Uurxq3pc829P6teXu3/IngyBKeVmNv
l0Wd08fSmDE10ATNLqYMFUUHo4nLtdS4VloC5H22VBRs6T8ahyhZNHcaOSCJouDnC1Sydmt9Nm2Q
XQhxk6AXSFiR5KWiJywOzdwJjQuiGu3vZ0aIOyQ/aidjuiAMW+6U67vM/JKqNqSFJIvSH3ZUZq4J
t9Wkl54bYX6n0O8q6iZUBpdFD8yUYoFlUThZ+GqwDkMvMzJPRLcuatX4QTz/UFT5UW5lJdzKaSQt
RbeP+M7Ead6NegczYxypzBvnleBNIDg/ZsnmIMCS1WsUmt9/+x9WgXvsqnvtEfI7hPzun3jkmEKd
OuZbiTIhcjpu5ZRrZnl/K/zjNI4hg16NQr3B8u89qdgx/KMLgjKGGEm35mOL+4NL9C2hLYAr+Prk
Pd4GvtIGENvK1euc8LQGAgchy0GqXPXGcaP37ccQRIOgMUI66HuKJfoTaP4db/A1QMrwb5aEG81l
KiS6RZ4nuxEfA+dkVpDS/dUUO+6kA5RX6iEG7OVGPxFZ4DBqXZIRDJhKtYzK5weU5/TIgACQWF/k
6F94fWSofYnMCNIdWO+/HnZVqxEP6qw03VKcoDHO9CkVohCwwtRjecEJHyKBhRSgx5qIMshFCW5j
C+64DEDoSFULywyOUukFdiYLtUOuTBY4LuFv9AgQSbOmtcTCOIpwH8JpWNxl/Yq7fFaZTG04R+JK
D4+74AFTo0OKttkHGD8s1GO0Z5VSzB6iuTPk9luwSBjn7Uwgeu8Z6V2vnOAgu3RPjZq69VFf/BDv
GxfuaRSTMwRef9SQrW2OeFWflfq1fgzSHDsX572CWOraRkuf70UKX1VYTL8LQjwPRG2Z9yVc1Z2u
9Qrq+Rfcq812UqXOhG0LtR7++4d1Ih9y1OqXgLS+IXuQWW16huf1R8a2E5+luI9ZzIv3wo9jrydx
BdXGegFgITEUikHbI+UtIuSV6pq5bqwvKhwHmgHFmO7TYimu70xwnl9zeyG+kZ7OhIo/P4x7lFQy
5Jk2F6zK12euHR4XfOuDfISq1nt/CXkohiFRhLhwftzG9hCMOMRH3hY+M2BhkzNhJjuJfbSObuXl
4Am/VeyBG4dNE1yngGKzBJzRcz0A+i+p6L0oy9b34MT5wfjUWKHh7Aq/kIm4HJ7MusEehtLZqobV
bFAyur/plmXp9jw1NlU/XX9CedSu6eqKHJg3hUL9TPTLs2PPbPy+CnhF9daULoCFf6FLKh8ylTDI
FrtnyVax0Tnn0NLU6A48Fo1Xa6KEUMbvSu35djS+2isx15YzQ61PRi+qKjibf0219xnKpsdrtE8/
YqlsK7i9sifO0Dbra11U7Z7ALboXtK+h1ZcQVg0xhdIyZM8ybf39h0bbiqi0mTd3a65vqzLPNwqm
eJ5r5i79iJZ7e4QXKWzfnw8hO9Oy++n4YEJutuoNvDLS2gLEOW8tpcZH/dnWySkvNo9kZA3uIipX
EiffnUTO1MS+Q0Mf8SggXxZ0bHsMczwFAVogXUv7HeVarTEPKUNFz/ogQ0Bzm0f6JqmeEiI0f4qy
z6H0utB4xoevb6NYeoZyYU/6MTQBcJOVoaafjLAzNVQ8DMX9oG2I5Q+iQQTp1o42iPkKjxjOX5iL
nm2Jbe6jW5i8HxxU1yXEETkfkc2AIq9qAUy4mSgbXDkuvlg7SU3ogHBkBPWh3S77+DM55++9D13Y
IuEHLP9kLXW+Fx2lPajAXWyN6Q7u2xUSJc9WH50YW1JgmZKwn3LR6kg+apzJ0lKitFQ0iluV574s
Ukw8mEMWnUMu2ia9wF8/YRGz7er+R1rTsSK2uMozgwOll0XNy0kQ/spmUeIJUuoB4gCZ6NQ7ecWU
Fw/nRBndQmQ1B+7yxgvFc+CRYtEIKSJGW7J/SUWoOXn2CCZiu9o4lhiJV1VO/LdtQfyi7E5HqhTe
hA29ME/6t7kXNzfuC4n8q1V6/XE8Z9Y0wdJ91h/TZ/JpUwYdXaOKAcmDATGxFOs/khFs00HVO+jm
otHb0yrgUgC1SSTk5G9zzW3q42VoENa6EX3Z9j3+8xajGj4SwJKKosf1cbrwLQs4ZQWsyH5es4Mf
+nfy4b6InFcLL1BV4h1zRHHKaevvgf/VEnSro1dBUiqN1TICLWDstcNJkOWJ6Cyj7grp/XY57RN4
TiDVtjunQWoMZ0K64p6gqfd6Ox/HuBQEOU1ekIzpEQR2xUL+zyCbkxxBlT1p/bzFQupYHDmIn/i1
NoLyAjnQr08qmEnlr4nEBfevnBJ7DXmMinIlV8RxmIbMQpmgRvjWzAVQZsjSe7Vn2oOyfHnEfxFa
cwJIIr2S6Crt9yasiWV6D0jxDLNNHnJJEotHIIUXwxaSLnc+CQ4JofN6yTuK3YmDIn7Ls5JQfE71
ntxhVhLkTFfSHNE+7uZAtoHjigut9K2sJ5iCyQ3kqDKzngrtzBb5Lx4hMA66bgYtC/dotptSDiBA
qjUwPBVOwZgVg2ddkowTaFuOVNjt2BcglolBAo+yK29S4iZFIXKntV8RmhsXbC/qsHDx7u53s1Qt
QMugxZ6/ncALbxUFcpFu0vdvbd0cC6kWOTECJp9GHdisxJMY0w+hjCZ90d1mD++DiNRCjS3isr8F
mLIMvf8tHRl/jxMF8ovJCUkxR69y3i2b8yHnCDpOpQb6JLzTZPhfUBCatnkK0U7ARS0SwfQKp2tD
cIB7P+YOf5IOOm64hPOLlSWCAjGyhCdhy2aomRRxTRgHcJvdDax4Rlu8tLVYDeRoL6FW69E/2QAt
1VCX1bLDbdOkj9g7Z2lpGEK0f21jsdKTe0oQ1+Ltn5jdLibOTOVm3Ephwg7WJSSAtbTGgHDc0DOG
4I+DzfKRRkLJzbMJ0rHTK8DGnCaVfmaE5MAFQ3AEGw0FqHacyfoD+3CrT93xlifnXtvPDDNsDbJn
qPSx9AyBpqYR0thNQOltEo8oLCOBdtKysDKKZI1Kfd6mSMuhAyxqYnOeAFSiXHh59mTDRFBk6guA
hsjrhpHnsY6i2aauUMAtlg5017Xh1YOzGPLT3983gk0Hgb7OT0ffXHemaHAqdgH9g6Q7brAjKrtI
NpZYGvGU312ttrAWxOqYQ7/+evpCXM3APYin51HE2ffEf3T5lEywkyShQXnDaFYZhVWA0jfh0YS+
S1BFsrs1H8oBkl1SqgNNCMXGqSmoeEfqaGJL2H64OKyqtt3/KcFKka8LwnlYxXHzpOAms/q8QQVe
Bj5rK0EpnN9kRNncs99Zup6fhHOR5tmngGb7FNaadE1ReuY6FoTPlkbci8lIiwSXSYEXXv0TU5rl
r0mqJesZTwZnAi+0apTRPSX0eWQX4e20v2Cbg0DE1rAiQM0mE1xzGWAJBWXM7vwHN4P/6f5QSdHL
SM2DKLGvXM7thVFixk33CQJBHm1uPOoKKbZAgBNIm+qqGapea116sTUA50pGTzcnacLC3+ZZctSL
Q5yZJ7vDeCrMeLQrpPCwjmApSr3GvmMKc+BxeYAbpGBW0hh4O+ePjKFAJGUjUJNZ9hQ0ayKtY47n
L0bh0cKs2nNpJwizyLiUBE0MEXdhQFzUBH49XoQlT4fbw6wPkLegHaqbGmq8y6CkMeXomzRPdCyf
rbiGdo9/WiFAn+Q8Drl/4yTSeSWw8anafRcCBsfYUXwhp/3+AWFoJmmyAmSYQUzS1qtZqeiU64fm
8yXbbVk4xfFbDnXmXNu099zEdrRa+hiSPnykl7lSipyznhQMCmZhrzi+ICeiBm6eqhj7G/mNNSoz
eiwOcSSH5z5kjMoNwgSzw9boeOPZpSfItiFvvekfYqzbxmyTbS8nTQSMDPdHw2reKoj7rkbIHjsr
WOacvNylSgfa+L+AYtJuS8QsbvwVI5/Ajt4SOdVYxTn41xZXuwDBi/l/LM8Z+qyQfRAJKXBs+sHL
r2/qPAyCldCHVPmfM+JRdC07hSiazG44YZcPBCpWAbfQem6M4NKxZxDvgwccthULsK1X1t6ExUc1
rHoIFIydh2HZU6v1K8E9MORHL7JLBIMDfOyjzvHKTdVy5/8+zQJWgcBIGtoArHGzV9HvMzbVc0/a
n/SmrwzLSScCqdXJUp3F4+LujZIQyjt4+A2DYUt+wlCUY0j2yR3MB/YqI6HGuCalVv7140RSVhMD
fDxNkiIbOXv6DjP7Hx0h67bLLbclxLqVohE3J+WliflbRpnAS0Z8z078jgBDf1rirR9HvrK5n06c
bJxyEmTaNfIOfpCoMpRcHbQIxksZlFbILM5TNOcT3jsF642Txtobdp7xaCFGSTTWV6CXXJUo+xjp
hZaUB6tiP7uZ+cPxGoy2nIMYVAgqwNOB/OiRgM8H8+VUIDFlMGjz5xnjwhAxbDL0V4TqD7i0evfc
1h7GmP+WxNK6YE/WBEhG30TFJ0KNaBEvLVO2YLvE2Fsiicuqc/bKzkeT1qhPxQ702QvH3WVO/YyZ
XZ23Au0dSOsocnktq8rLfjurQGHse+CZcF1FUpVMJRs16QRsA1WJhf9J8mcR6vA/eItpmxW/VDfe
2l3f3svlwnF8whyA0v0iyXsWLMlf1XZKKj/UIzC6/Z/mMklfAi/oRIHxmk6m8vWIc9W/oKJ5HmJv
uLcZtuDmU5AbybMO7EsC9XzReARKsdF75cooma59LyLXCSV3HrJwQsNHCPj7WkSYHusj3pJQGPBf
e8wdQLFRQQFWRf4sIDvLNeB/lr+BKy7NGc9/ulmShHH/9ATLTzgi4WgwkaM9GSMmqac7haltjcx7
AOZwbl/wS+xt9Ut4UfPQI79YtqAql1DLWp1Ncs8o+uzrqha0iyFyBpR+lW1/HZNJbhmnsjoxx0+S
xszsXUJF5ggamsFy1L/WZKdaWB4RnpjdsDOGkoGCjIOAEeP71dfASCX4WTryjnJnvWOJ3RmCmVOq
5EBRxB3EzRvck/Px+sOA3p4WdeeqWbygyyOai7PlxrzyOqPfC0g74nD+O9NIdMVbyR7laWf7Xd5B
uuTXSYKCo5sGyeSDdJrppJehk+7JhT7caFSzAYpHjEs4FhDMjYtScizvuzJfBg4+IrPhIOpF1knl
/kRFhM0bNrigQ63zUshyUdQcB+zueyqYahleoua8xfw/XPFjF1tcQF/u0cWgzxP2pkmV/oAn2Tr6
VYzCi/TTjJkuTGrilfkaEVmtxCjuJiqOkq2nwhsITxy1+u3mTDsF2WCmiU9Plm9S+hY2RZBubTo6
D7z0QPDIULN+Cfjy8Wo5Mqu3583TawfQm85ATK9pmCcUk2EjDi1SXxJ1HIVqucFlw/y+tpaFQpqM
RlPtx38crQg13NyIjQ9iIn9ED4yQYgji7o6dg5xtv8rJHo9iazPzEkD0tRELNauyacG4g15XnjZl
rzQ0xFPdSeBinJUuZ112wqpVi9ZOg3DF8QMplfVbtGaI223ZL9n5gtr7/E19gq/hCPAfOCMmdU3e
eBsZVjcliP3IRMGGFMFv7R9Jb/oP1vu8MJTTZOVC/oa1ygzPFChH2pSD+jkvfGRgQqIiW8z7mImB
aqQxnZGmw/zJnXy01SvcZTsQf1yDusS36kCozD7PuOCwumMuVQ7DSWvt6p8JrSHpYr//d39EomYX
R+57AeZPb5mVXfRUb7UZVzcxa86b16Bk8ZKF/YIZLZ+o5LXnXxRgx4lNqxv7rdd7e8JOeleFuKzl
91WEqYmEsyIlM9WFanbzw52vyQ8Mh7jatrQH+L66zTOwJwFNGXBcKrxwH2lBfNsHFy3hdYv7pl6S
HDWuNTPvOE8CkyUXrEwHx1S2+lvHSbEqO9pa1d4d4gTJxD4LdPVkFA/7PZXHnWqcLpwXivDvQ+d1
cE5QG+M6KlJrclyqENyuiUAaemHTeyPUtCpZOIBDAc+QpILRmHLT4t3tqHM5idkjzfr0EoBGh7CD
370Rd0CUvnFdSOuR8pfG/1cim8jU8hzaZM/XP2hOLu83AQIX+47nl0mYzj6HTCarRUW/2SMLudVE
+hz00ec1lEdOHQj6bsbyvgONh9s7XJO6T2hCYR7HQ994waN+AF0bFfBncnYz6Ma5Nazzt8zOFQo0
8n6h14kSXn4mAMrDZzKU7QG6avCaDHQe5V20QROrntbZO/ogS3MxqnIrnw3aNa5+/irmAmbr69I7
8cySkuqIKLRF7c2QfqzpHFZnLiWR5RS9XB8pjHXwd3NTX/m6a/CdDXOEqIdv2ZQ3tI+Iq4y2xD8V
/InniwJYfaSCqA5X/uaWKFOWPH4JiFLCqYHVnG8N6sL/xcfXQ7350lZ0CXPkFxtLX6YFldeXkrI4
eQtG1gpRDVN76auh6dNSBE4gXdQ3FAJydujVE0RcP86TW4mUaNLBhJb/t5KY4LTQlD/vsR3C3AeS
XGQ09Jg7nOqTypAJgrdNCOb+Fh3YoA+I84dn+zmjpVNgWCWhvlHLbNHxX/IRH6JYPcJ1gooUA1Sm
5W+4qGGcjTv18KyVWfy5WIM8Mb9VC0FpCL44JaCdQlvIHdnkVpjajOFUOxw5s1C5Pnpr9jyocaWG
hW/s9ySAdfqGV2nVaPjCFG+mRu+TNBM9OUwxSfnM2uBcyoU60l7fI1NiyequKvDADKYu/D06H/PP
vxlvGQtyhHZOwsUDEbXQjj1RFiKEtuFGa9ge8kOP69zrUTN7zXqqwbiadDdJWmAG8lLQ6+aZcyrM
FIcW9N2G60WvyHpVYktn19P/ERroizr00AH22AzhmhH9Ud4bDwMoWAA/qbQEbmznqA/M70rPvKSF
0rX9m+668YCwAf044UlCblG+74i8k5CSVKM6YzO8ATFwNuyyqOjZCkyB87Oap8ic6QVdCFkiOXYC
h4ZK7UGyHTI9KmDKOiP58GXhUPKgBgUX5rHYvwt5jvS6fIkeE9Q5ASHsPT9dA/4/Xo+RyRL3GKg2
Q3iizFJ/SD+yFNicl0+LPRN/XE4krnfPnmzzTZN9jX70MWdG7xfA95i3enPOoKEVNkfXoHuFSRKA
aa0x1ikMt99kvTNvdPuAF+mX/afLas/lpAkSCCbpYMkKr4OomfRcEjDveua994b0bjnQ49sR8oVK
WwQCEoZcn3TCPx3EkUxa7LzMJEBCM+8JBX8+PkEtwksPtQzjt0oEHkkKjHZVqaB974vuQbcyx4vF
x9iO3fJbiMK5NPR8J8BH2v2OsrorwNZTs8vPKQNC4V4K4moAoxzDjo60bcKhGV5+fRK2m21BpBFe
lqb9w8Psbeu/Q2Y+DoG2eGbdQaTJwVOXaQk6roMqlq85SJjEViF5kjlIeuvDo8gnSu5gika59DUM
GpBjZMih0b45LLC3HgH9XJ5h9vf14YAcbUy3ZBEDj7ZIsAMJBTzSD/2m+3VSScNMnu0WqKq4diH3
LfMcjXBVnskOeutxd0Cir/KvEdok3q5QaMmR+WFubIwTIFFiz6OaKxAE4o5aEG4uSu1673L2tQ0m
5QOm92QZiXk38SkUdBm3rQ0ZMeuOtVoG1uvFyMtlhX1bLKvnlLbzSZVYfGK3pCcG9iZ3U0sq+nKp
9VFRxvy9YDsPg67gAeojNI9RZ/bff95ZflcNi5fu/dhuWgoaSw5h/zXBsSrkd41tGSQefLPSOmiB
v0LTgEyMKsfsae0xzt1JkgtD/uFPbJGmigmU1Q/7gObfLXPvr/8UfmTJ++4ypwgpaYdm1lgq5bDg
kCAmlD8lBBCYLVHksfE9ZWvZbY8hWY4UrWzVRTTn/ZEeGHJoHSZgWIslfg0u99M88mqh1TICFuS9
/VRsquudMb0CWjkktCEr0F4Jdayt++b1wtYW07AyAEaltRqI0DZYfw7HA7vZxvwncXxua0Twl6k1
x/iJN3UjpwbJYeYBI4mFnmteerAHSVUynhBLFUaDkDy6vIR8meGhlMkBv/bYmL92BCxwjzraYvCn
pzdp8y2F6V9xfvOp0hz0MFa6m/cWe6iORlvdLQ/9pUiFkEEnty9xPqosvvBJ9Skg6rkR7JOnG404
PN+GOsOht49JYYfO1Eo3HeFIN8kQ+t6fEQCd0awL14EhbUcbFW720iCBhzyFz3tKFh9a7FCoGaD0
OghPWMdAsA+gRtnIOlpRPUTrWuDfYT7XL7Mxp8anM3pTKHymyD2Xp1EWSbsR4ro8I5UzzE6ZR1/O
4b4ZpWnYtPjMtjZalQf1sHTRhrh7TJmkUc5PQTyHs+TEgnFrEWJnBa1f2P7L64NZfPVRkuACY2sb
Y/T4VcyiT9MoV/1G0AAvq6atV4AttmV7Ptn8AVwGIPxSIGpGAjXCYxRn3Vd99vrkYSOz5U/lOkdC
U9OIQ1Cb6wxfrQTlZTTbtSXFOECQPndD01XlYHANTLoem4QmFfxbUfhr7UA86xAzyXak912PQDhw
ChvojiZ3TuMWF3qn+lQBfhVdXP80+lP7iYY3yaBekRXZ75ZzKXce3mbzcbNT3ZuCQZbgZji80hQO
54NU3GUCrT/PdG4FD+m2zSy3y4SewhKzA+4i6sP1WNeY5deba/gxapGIOFC0UKuLVHIi7Szr2sW1
ul2OyWehWioDKQTznR0GVBapJKGJNv0WdUxAMsZJkqMX2LBeqyQF1HRGlGqObSmNEz9jiAxgwwEP
eKwC6Ur+QpVjqgtVaP3fH99rQ2cJT9tTkV4eXi0zY4rWyEoeAdMjm+DFD4NHB3sGnvgVdwPbK/wU
fEIEdBd40fCJ3uJK9LPwimKnDHCEKJvwJIQ7Aj69hNEIkjF6LkT6aQnAF6+oLot3PkkToG8Z6Jgf
vuToEMgHsvm0K1KisXKu0MP5We0gjizbh9IRFVFhBmUJ/P6y7BLIlURL7zTKM2YQTPfYnt3CiqdM
29RAxM7OR4fhunCe27YFGVFFuS2xcj6NMP8Em4aKmbwkADBfJ4lCLB8rb55EXofwdgyycd4A/TW/
KAaVIWFZsJQ1Uy/JthREHa2cKHoZmBFxjI+BtBHGLDfDsMNPNP28xHIZAHfguN09PxEJGoq8uXiR
XBZvFwb3yOsmF1q9RosWLOxWaMR+GWtf2zsXdO+M+gftKIBKYr7iCx4CTnUiDqxFAh6iQimAlgwX
t9SpTcKvfT0lx/2A0tyH/PQZWCFDyqKTwcr1aINmI7oDCXZNzNI2bYoVlSRCxsF/o+jszrZIXu1C
OHHTRJBJRjCPclQieex8YdTW9lawVfdxhk8tR69Teeg2alDyFFKPwNXDZvEcTToy36qksxWnEXI5
JsBxm2ueOEdhrkb0JdZ4xAq42FB7pRUSkBpyfpugQ5kpP2I2rAJZzhP4MHu82Ycuc6VWr+n9SyW9
pBxsnyTrFGbwu6gCnfVTLwNL8SjHVoJjeD1gH+va2nTOgVZvCAoqI44/qwSMcpRoYfm9jIYcqfAy
I3nRmSHRmDWPGLlVVLTmXPAItQ9XeSKUvPF9APNDmUGD7gtxsQ6d6btQFvfmop4Remunj+HMWiGQ
FiiGTGqacZEhJ+EiM/BYYAHvPuAAtZf+8es6U0PuqLnpafLI5rB1Cp0LBVNWcxXRogJ9viZaHR0B
ui5hvCPFib2otNFmp/iw4Dq2V2odPTXURmssT1MGetrUoRZc6iySzH/DjSbcB3s0GbKGVZUbtVd0
lD2ElfGeFE/NP0iKL90na7+Cnmyli2cm3h6TkAV3rBrAkgFZ/tCIktlqFA6yWC0i0/03NFMUhRUW
/osZA/08yFjm6oanh4m6/xfgK3KYKKnyc1k2000KlB8q3vwZTe3w0RUoOLdsNA6y8DS5zD0Ynutv
2mHpRkmPENG17L3Mvl+Oc2RmygeP1JfllwqYydtpxjM8bdhYCBOhwjB8nDfIBncXmReJrWZXA7KV
v0Zt+PX7r1oMy5srDcc4JM0Dw8k1AmunqQdwX7vSC68oZlKDgP8VJ5gquAYn9btv9562RaXf4wMf
7joHlw4FSUIRG07a4InQDhz4ikTRvuGQErW1EDO5tnYQCJoJi8xvU9pBMcHkDGjH6ZFL/7+8Y5rn
A1Gd+qi0Pg6fYkdDvxQT07Whox2eUzurJ/SKMwnz0j0lgrjOkwGdC4oYt+sjaxFSyBDgbNIQH6mI
1/foXt3ycUnAoDDS6x07rYIQAK0t+0uMEUfNkH/RdNd9Dq2mv8VwXkxBZtkq8BR0pl+zHZP/gFRK
GFjvFvGScrtg1P9REViFVhdY09wRLSFDRUQEPruxHwMV3CvACxMDmxPyJhoylAIF73CgPyUBZQFv
ur/D5uMTvOeA0m14ukzq/Y99JktxKSg02nV2zMgoloFnSa/G5hWb6AhsKTxXLq+nBTmccBCgkT2S
hyDSc1H4ulyZNBPNG5zC3Q/3l/HVivAAmx9ziNYUOoUoXnanfP9RWpUXYV8e0zpA0Eu6tC6FqRli
0KqIQhJUqQNZuc7Gj4xOJdADa/9B6smd4L64eITg9W2WQvccWyoG7FLyFcwpaJ4uWD75f4Mi1aWK
1KvyrsNlbXjSPEFUWR7Vbi9/yxY+3PX8VPoM4kWP/LY1VoYTygF7iRRbsUVjmQcXKKp79Y41UfXU
SXxrdlis2qKJg2Ty/ml0V5aBQ1gIdOUYUdq7d0xAsV/EhEqMBFZkJPc7PzNocNcZIwetQDIZfdp3
z/j4Lheqzztq3CtzHyuY1DxJP+mnKuV4KAPFFjh3UXqc3xH5ChcllfbvFBcTqSx8SCtE8MLpdJrC
faXii6e9xbZRVdJqLF3OgSTB4pty4K297xw/OFThpSqP5qtkZvu1wkCfbi9m53YwbX+Wd5kDkD0l
w5ED5ADVxIQUgZbpclMlNwbeG4Um3fMljKxWq4QEvppyb85Xtyhp6Bb9uowkW1YLW28EYXBrN6By
teoN3e0uSMPgKEuGif6Vag7Mv4IfXnjCrsz+/RmWBudH6askLGilusEsAo+3kzmwza4q1/btZzyp
VQ5PEUrKe1sgdsBh0GmMNraVjNUPzE7IW+PjJzLLDTvJkPTgSEwz33O+EPt9TUC0OZ5gJeCT2C7z
PzKojJ/vBRR31CKm0Lz6RdYWXx1QEbJAkEkYT+gg2ICiKxuvZTx9vCQMMnpa6ziNujlXDM47wbWe
rl95AcZe4vabuz9geU7P5xS7i7yXUlPDpIzlsCByJ9lKQ/vivBLbuFPAxL68AIp+r+JmiGEFZxd7
MhbCn7qgHA0+dsVIufZIyRYRP3A3WkEl3a1En6YsVeg/Ap4RN8ql2k/oq4msXDQbOyiuYkTGS4WA
677fXbMkFlcRcP1u+BiMzIYEY4DkNzL662fTyUpQxioF0qKelqm2r0h5ZkzUdRu2L4I2qCjG9Fmg
etWZg/FQiFAYyvXkGNUgB4fJBKTbUyi8Gpz9Phb3aN44YcwI54BzHieKTKmyy1EBnWwJ++Qw5MA9
tjAGtgXkU2K5ntdMcKphypDZO1KSILbcRQcBGbSXNaNr34x9KxZbYn/ZLgOmAHoR4PgjDlWZ64Yd
0lR7wM8doyF6cfyIYx3mMQ9F7I1NS2fGH4dlaxClRlCBCGBEXyz3GuKi4l37Ya/N7Tpasf/Otn8P
XEadt+IIG/YYUWfz8qEvGRdNWntH3KuAHoqoYiIH58tBWJEg4TVDluRhzYvmalojLX/Bvu7FWFpP
KzBRmuvsqhvYAVcMzEGrIz3j7hZ44V6uihEeAUHRHKlx7iZRKZMK+trjRQhZJWtjhZnlJ8FiiE6I
8+jtI40jCbbXHrN+fRwJVp/Xl+4rvvEupFNmWs/Vvae5vsNyisNT9A7k9TQZKRNv28U7yA9j1MsG
btfR8rvesBgQNlSBDNjdFw7StEm4aWMrOPDIb+IB9hqoVASqZC45CfXhFXAozjHmOnbUBdZ4crgb
PQKq2S8iAOoX6oeK8PAWQHXS4UdUblHvHI9BHLCkwUcK58LO/CRIWyoeF/mXGdZxmxeFgl6U7qp6
a+ilOLp7NdBTElKzJvrEwV5KTz7zvhW8K98iizdrZbgqXcL80FaMhs1OTgLoP5TTYb3bp2KbRhhm
8sOGDbL7LHdGiYgNpl1djMCWuGRhlb+Emw1pUUtT+02GVCIC/oJuTetj9MEUv66ASZFEH75VzuPM
W8Q8L5F/KdzVyktZIO7sgdILQEWr+QvBdlQWeND9A1zbCrkEyxJATSF8P5A3Tvm0DJxfz46dHqDI
E2qiyZJZa3IJk+cnkkpPG64VvzFVGAfkIQuXy6tS+umvCH/2iQZcaW5PJ2JrwVXlhda3gpDujeE1
xowk+S6KATrUtynyfWUQw3G+DHIjlSYZ56J3H+gmmhxllqOAec1GaOVy7BbfgUyfQ4Dgn0IZihfA
PWT5Ow6QaRX+zwHNDlm0SP3N6ALeHheUAPAl3110aNdk+f0zTZ1nHxNP/nv9WxJsIDP45F8DXy5x
iV7LMkGCJrnpeOHEUUr5s2ev7p0R5q6g36UUJDqXSx0VWb3jUEywBv7T7BwmcMpLPx0UckYdUINP
Hq6+EaPxt+OKQNnYk5eldNerENDaYGjwGl1yKd5ZNOFWobZKzi3zRBGp7RGyA66mD9pn8DfA+cdL
qp7gidSkQ5Pnq5haTCRoHy3we7pKn3NbBQJBqNurdIdjEXyqtDmnG/JFtyAgs+EJZEHKq6bSffJn
m8b3lSaLI5bPKZ9u/tj75mVPpFMYWAnIyZ8nunYf6XV5yX605KQdZPwqO+eqsmqGWUh/2x9BNQDY
w5wt0xAQ3eSo+aeSpplkrkdCR5vH/ibmeoErcuD/juiELUSq3CDlMXfju1FIewvxpW0qTBm5v3QC
MvAPjjNTTMJ5o/RUUjSEL09XOz61wMowktv3Ihv8XAH0uV4MN1xU+C2nYiU8Y+LVIcREA5dulHgg
VQqlf7lWOZQD8h+a3Fp6w8cHfuutmvwQwTboi1a6z06dRQ+Z6yrncEe0jAMtXaQDdAmnoAmrjIHc
X7Rs6GOLyifHqZYOQSP2Df1wSngzOZVGyehWxiuysJYbV8ASAxzWek9RbEVU9rSM1qCLJgYlO0gl
vufBi3W8dtaF7wOvfFEwLdzzFxEvTtX3qxN3JZ6wO2tS4QWoxA1Q127gIBuz2ub/8YdRElTXUjKT
CuowbVdAhKVYkJ2PT29FxjFTCAFSghoIGyHN0Jf/rtPh6xdQOQwgJH3IsMetL/OIuiv9eficBwQY
iO/fvork1jfNj/rS3S67XdhwvTrNA4YlFzwuH7zhRiml74pC+4oNZ1CY9TQ2PaSD7acw7n8riH0/
KLXN3WJ3wa4/XRroNYZ78m+yzkazFFQ5tk6dKr6lGhmUSKjPScqf1lWrq3vAoxwiofhwGaJ2oG2u
x9rOLvDxSm0t0vyJSeSJh5jK3pm8vZC9UroAiuxorHSIlDJqux2uQhsqx6/beT1wsg0KwMRmbkCo
mH9MRH5Z+rUAjoiE31uPL6oufuVBHJArT3HO0fDynDIdT+X7ao1fqX7b4aUbaOq5wQSSW5hLWu2u
NDhc/X6ihKzTI5J8iNSJxXKFFu3fkrtKaFTSy+bOUW0uiHELlp44tnGTaYOGlIlG0zdSXu7wWUMY
CW2b0iivZDaabmFK1SkfAXxoMeT5+Ja/9lJcR/3HzR6G25sf8Vk27KDcT4kdbdy5oGfYGhedp5+h
IUkrugCoU0NGFX4r/RIMLycvHH4uT+QTcoFduhOHTldddeVC7jxDNsALHuld3WX3b3tESKRvroiR
Xtdbyal4EohRJMHAGIHe2UKWe2eM1UvhKctpyvH32JWknv09f9Z96NHLUwWpxvwiaX/6XbBWAPpj
Pxk4lkPndBf8C97TqT/QtKbmv4HwUA193xAudk41GSMxHEmUpgUcuPNO7EWPnkwFCOBUjm/VbJC7
7Yy+uUVp8PEWOmm4YScmxB7hw0Kdl2BU6gBugmRLLi+z9JrnEdUvnROmhFGO/maGAHl2Asi9TbKi
0wr+Oo9RRmUSM4XJX55tDgt0JvfxKUaYZn81OKDiE7guxUo3eGFC/+V27nydHAghLSMVlrg86xa8
uTLcth1W85coKdsHz52TkgaJ/ghkpsy6OOSYXmCdb+Q3eOqPXchs8K5whi5XF8HW9HTcXZOl+UtV
1RbFhJGKtbYxtwkQ13ZoNjDKIKkyxTxLjYf2FAF0lVV87wJReeV9kfsIfvhlp3BKoWIw8LOE8ho+
lv8rCo1EzOWiny+XoGEig72nTkqiijTgpCLuYAkoYyni+tqptfyzM9lIaGkysXHTt0VSNBuPZeRP
cZDxML0rW2oV2TmyyKAi1wCpI7bVUeFVV+/bl1LBVJZ3RY4vDhJ6jdny78lmjau0ufopQPGRMeln
1TclIbQSAM7wcg9ODvqrudGmTD73i+eVNCa7LnB/wgKb4nF8YqtMzHrZbYPzQV4Xbtp3tIHh/gYF
bFoGA2/GW+6rEgZLpY65in1CcQiBI6rFM8m9rt++t7qpXFqoS/Xuyr3moUIaC5S2945YYZc7sdAl
qsDeLUx/3n0sIqyFhLCRBbgcjgbkxuQJX1kr0C8nf71RDU5GVLUxzqlgn764psP0dq74yJgwSE3Y
FoBlUPfK5iHG7jmVhfQAAvJs7Lhp7945jQD/0JWMJcymEW7FnN7pbgJrINlXtVtARGNQBLgCDkzL
L4RuD94fKlITYfsl7Z6WLipePjqrYpmcyg6QliqB9LI4AHBsb1Ed1VrLrhH52btVNpBKTIudwLoB
lRIgLGMBUSQCBGBAM3/mo/1BZ+qpw0BCIWgUax0+pqXrt5qS4B0f6083sDQct55UYuRV+Qlh6GaO
WKH5tnNsOjfhbsj3xcCnpip5R5SRNg4fEjx1xWznjHowAsE/N8RRDvZ7AB957t3y39NsHbaPUrvK
bg2v8eFaDcOd25wpv6ZQWhP/hlJWTeEX9N0H6JuiPs/L9Xzmm0C1gmsG/z4s/bqAx2UsMxGk6w7i
5PsJtZ196WwCUdeABeTui5Exk8G3EPdL36XtnyNd50fy9Pf+dYpGuFEfXI1x6ybxU6Wmr4WixBDX
DNYaOYhjcdT7JBUWFj7RX+mLdk+HL+gDq2FEyR95AYdBsbsJFTbhMLGx5N3vvIh0Ip7X+/9pzPXJ
Pp9sAXn90XLOrb/4yn4C
`protect end_protected
