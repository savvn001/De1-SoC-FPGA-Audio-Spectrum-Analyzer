��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��Ìg����yO��ǿ]�ج�/i�il��{�{�.�蛔�Ԯ��>�02&��Eqp�`�F/��]�_<*�2���#�O����2���q�����Oy�M��ߨ|�`S�5�����H]1=��L�ό�#�����&�#�:X\�7��w��Y��o
�[si^�W=c������wIs�Ubڬ�+��w7 ��6�7�4��w9,���9A=��-�֪S�6����W�S7�O�[9�k�T&=��}�aϬ���kio�K֤���C��~4���<�q�{Y��='>����m��&����dtzM�}a��[3]@�^���4�#bY�.0��Ͻ��]8(���Z��̛�a��Bf�	ך<�+lH}���>�$�]&d*�NFy����,�.*]�k�/b��!;NH	q<��!�q���P@����$�k��ܱYz�`�����f�1�]"O��m���d��e��8Y��ԁ�v،����yz���~@c��>���+�P|�Lو ��zN;N⺾A�-lc)WY����NyE�b���T��k�˕��&{½�k�!pU��J�.Vk���V&�b��uLp	Q�/��G�\����\��x�k~5�s[�4�m)���O��luh�m�?�0�4���Fi��zk`Z�L��s�B�Gl3�͋�I��������6O����my�G��C /�J��蚜�'V��1�#a�A�/m�_�!
 �lTO�ͦ	�"��]��r��;�;|�CM%�χ2�-8#��}�o->��v�V��Q��f*/FT��j�#`�&��A���m-˸=�@
W3�;L3��O��3���y<�LBp��*�V�����'	�:����u[��`�E>[��l#r����ˈf�<�CuuU��~��뫰�a�}� �3E�ƨ[�(����M�:��ꪯ�
@r�
��h����*8��V����1���<� \V��a�dD ��m�b5Q
}"�Sn���Tg�x:4���c}#��V0U����<˕0�Q *G<ɚ_��jLn����;� �ݡm,���q�e���EUB��$�~�)
����N����C���a�
�S���Bғ�x�Ìw�<F�GEs<�<y���V��ӨD�d����G�똎m�2���D��V8�	G&7~�?2[a W�'�����Tm���b�) .�L�ⵠ�2��Z*�[��O��H	!MR&�P��|K�����r���k�IĀϐD&~}�IM�=�ZI���1v���M��KS'O9nw�e	���%�a���)�!T퍿�[�j��8�e�{��G� 
6�Nd:�K�Bƌs
tn��3���ϑ�ss�����
bm��AD�x�Q�|�4�y�@P��p��JR@���1�m��}�MDJ��4х���M�!y�P	���o�]�.J�䙫��h84�#aA͞�˯��W#W��-֟��c��B�p&-�#u��QF_/��{�n��M5CSm��	V�5=x�����/,�{	��t�!�g������-�F}'�)�	���uo�����W���J�[ɕ�*֏���60R��e�u#�)g�<@��-K�j_��c�6�	���p����c�R��uT��������Z�$?%��k�m�&�9j�M�`W(��RG���X���D�szx��r_���ޜ�9�$�����`���*��p,��~*�?ؖE\P9�q.�0;���ʢH���f$1m7����q�j����;ĚM����ٹC���k����N'�� `�0ж���*�X��$$!�ٸ�lG_�q<��@�&[�R�ۂr2ɟ���༼������k��r>��I�(ᲀ	��+ۋ@@#�;��s>�W@��m��i!"�*#�Nʨ��>�[����ͮp�Z���V�(T�����k�mx�X��=�Amu��[������7�V]�774�a�d"aM	W,R���" )�כ�$�`L2|�v[�ꍓ��)�!��~�w|hg
�uxj\�$�2S!�{�]ji
�Z
_��3���@,�qn��g@������z��d��b��H'�X�(O��\��4��d/��2��;�nۻ��� s��aN8� ����=k ��~6Z��0H[�,V�H�0�����6�V@C�tkϣz&����"$�jY�;��RO��L5Xܡ��y#�z��n�f{zGR��9O��bp�e����ѯ	�1y��Q�ze��39���舢���6H0W�\�M��	��l*!�7kOl��>�m�Bu!�	��jy����ټ�'�׸�u�c�T��}k�4]�b{�DFYƟ ��Zz������Y������>�蒉�~7�&�f%Y�G��,�>Ű�UK#�C��FB�X։��h��	������)ۑ���Ri�8Je8����\Y�mU¾4���7o�\"V�0#��fO�t��ٖG�2ut!�F�|��,z�D)�i��C����n��_�wQ�4��Y��BP=Xo9$ �G�.{e�N��������s2��ub����L��%H|�zYS�=����$�"Bɝ.�+�����"�����:�W9�E�&A��}3fb��?��V ��Rp[�ޏo��'�0?�,���ǅ��c�)��&.B9��;4=YuPm�����.�F�=*+�d]��^����aoc���DrЬ��7�i�g��}˾�Lr�G���⨍�PP�]!�2Kg�c�� �N>C >䁵|v<R@�|��� n�n}S����	�K�g3ڏ���>7m:+��%q�r�m'ש_�
�#ptvM��s�|iգ�+��V�]=q�QH8�����
������O_oˉ�@-��7�-Q��&?*�ى���6%J����Y�m
c������Rl"��#Vb��>�ҁ�j�u�h)���?C���lN"F�{wa]�J�uQ"0����ņ���g<Y���0'��@E���5;�@߆�	��^��!M"N��s��=�g��1.u� N��r�T�T����CV-� /�@	V��nɥn�g6]1jB�$��8J��=�Aj�����Q*�Pc���<����xY:��T�����}��Yf �G��c6���y�l]#�MO��}�KN�C��{r�/`%_В���n�����0��sl� ��'�Jt!����|H�ίSY�&Vf��l�O4^_��@qM���(cl�e1I_A4��2�����M/X�&Zks9��К`�%ܶ^:+2}y�G:���X!ni�P9��:F:�]�_f��p(�����鋦%����$#&���9���϶:nxxN�"�fT\�0�� ���Nl9g9��P+��À�K����:��:=�ve����˓�P^B]ul�Xi��x Bq m��|y폽��U���S��*g����/UB��YK��[ϔ_�֍!t����ez;	�p�9�G6:g��M� ��_i�u�e`�)bY�ꗬ�9;�
_E�^��?0,24Sh��#K�K@�oȷq�D@�ޔh�L�U�rH)V�T���#��u��,�||���p����o�>�^�|(�o�G�3D���x�FEA��f�Uр���3��.*Y��G�^�����<ļ\�ш�"�.0�xH��C2�P�X+�ZBt�F�=���缮y�Fc��11Q\�/����u-����ĪR*����
(��ɨ� �B*:}x�#��l���#X4i��L"���E��~<r{Z����sy�\ܫ��;��9	d������j�1!˿��$�u謿��>R��CtJ��U� M&�Mk���Z�(]�}o�޼�bZj,��O�+@i}p�H4�3V@I�8p
����Z�ׄ����v;��:�
܃~�l,,0�ז֖ծkN�2� j!ҍ�cك?�,�����"z�Ջ��h�8���p8E�������O�o��<d�+�7^��%u"lb�I̤��H:k�=�/G�s�Wd)3�K=�1�q]wB�_Q�����z�Y)J%��mI�ؑ6���R�qz F�Xv3��z�Hө���A��\�A�k>V|N��U���n��ZFj+�S��� �"��ǭ(B
�Zz~j=x�F	��{���^05�	͜��B�r\?��t�U>��Jf�DGU=�0�V!1�[Ӽ�y��:���������X^W`0���*��̔���<�Ʌ�J�'�xǀ���M��*�V���ՏTo��s���.��ڌb/��ϕ�5}���6.74Mؾ��������6˚x0#)U�RRۍ����Ɖ��L��uj��F�oz4)��]@�وZXNd�c�|3��Gin�?�u�kn����!�-1�xJ{��U�� -�A��4����ߠ�w2c�_p��[
� dq=�q�|���u�u/�������"@�
Rzڣ��S���JyB����;���z�t]�F�b�������*��K� �NO��b8�Tw�۰���3�d�ק�p :l@���iYw �tr(���hU�!�"Ϝ�@6�8���1��2u`q��H��,r��s�o]��R}S�(Qc������g�jk�ٓ�2�J.�z9�7(��J��T��3������|��P�V?����Ա��'�1��j9����"�@��e�8�����2Y8;\�d�RȦ�V#�%,�p�a�s��8�����NW�s����p �
q��T�G��[��[_�~�cX����Z�S1:�1"mP6��p`�t�信%�(��A���0R�G�Ŧ},���g�uJ͌�Cn<������s�\��U,𺁾TI
�-"��̈́.��їih�C��V��(�Mխ~SB^�Kk��2'�a����0�%��*����k��_يe�!L߈���PȔ~�8��[��2\)��5hrs��\��o���הa>b����u�⧘*���Gp61Ud�G����Bퟷ��[�]�Ih�ϞN8YT!|���"}���Ӡ�������"�Y��q��H=�/�EJ�BS��,�7���р���h��<S��{����8/��k��m�� ���p{��O�����IeS����!b�@Y�~�F� ,V"����,f�<��Q��re���2�F�κ7����n��q'x�J4�5��c��N����yTT��X����j���N�G�ˈ�]u��Kނ(�:�i^��)nLA9�#%�?fg�@�	�&Ɛו��Nf�@}�Z[���M����v���7�GM�{~6��JFs�EH�lPՃ��߬C����w
J:*Qeʄ�[JD�}K��ySȸT��1�el������l?��ݬo�����t��ߗ����Q�����ƿ0vzzqwU�kc�e�^�ct���G��t���������*$F勸�T��,|n�!��L���`�� Cˎ��/n���؝�)�Y}B������U� m��oJ��
�~��]k+�H.��+���p��/Z���P�mty�5f��wU�ɓJu�n�>%���t��f�3��X����ZfN����{�q0�1VjBH�f�_S�[�u'�z>k,�=�S��ն�����,2�C�s���^0Ί�
�^��� �\h��N)ؖ�8G%6�?y���}��s�$�$��Z5w7�d�$��	b6o໽ۏ(�m�q��uvX���sj1�7��%|�*1�l�_����ɚ�.��/O|�A���X��'K�h$����*Ȱ����e�����̡\�R�{g���6d�j���c��;�_r;c���D&{tY՗]KK���ң�������`q��sBTh���b�dQ��� ��|�����~����Q���V$��f��EY�e��`��
	���4$�s�]�$�[rr����ɗl�vݴ���jͥx���C�@i89�\�mB���c�H���h|��~�7jr��8���M����� ���ϫ��4������%��Կ�~�YHF������B?��8&�Z��T1ʈ�  �h^�VJP+�&��,>,�*%�i8���3��\�ۛE���4�.��  �H%��a$����X���8���3BC��;���UH����i��&+�,B�ڰ�A�����N�Hh�^����y���0�V�n�n$���P��r6o�K<D急��ؑ_Ք(��PS�AY�ٳ����W����
t锭�g���E�;Lh*h^_�´}�a1��|x��}}>�������Xo��}	��ѦǍ�=z��m�a���Q��1n�� ~ʪ1�yr����%4W�.�@���`V_��R8�S_5ЗGf�:;4=rCb��H��-x(��=�j���M{�L
6*!��e�;�W����B��;�<q�'p�6�Db��{%5�Xd'���K�J�xO¨
�o�DlZ�cib��`!����pp��<_��Y�YdN�o\_L�[x��Q�g*��F�q�cf�@o���ԆG�nX��� ��sn�����{q���|�3�b�4�'{��mAS ��%7�d�s���ӃQS�L�/����2��d�}�f�C6��ZBڌA�=��?�_}(<���������z��Yt�N �à�E�!�N	�#T��ͮG�G*o��,���T/:�FX��Aٵ�kTn�C�/#6�ާ�=����T:챂�^�����C�ño�=�}ah���n૑}.{�YiH�LG;Ů�<mZ�Hh:�Y��.i7�m�7뜻^�e��΂��!h;J��	r�K��jI	T�����U"��e����9_��%}��v��\3m�n&��0�i��k2�K�e�� >ogH���8Jb�R� |�D�k���l�rƟ�3Wu����,��V�-�F�5���GN�v������75�C�-iY�7��tqN@�{�ʨ�G4^dX�Z�;W�u�g�e[����t'��ѓ8ځ����$�@L~�T�*�����rIQ���]��$|�Y6��{�Ga6�*�sY�e�#H�/(����8l
h��i��G�Y�6�E�hgH $�fV@�\_rBbJȳL���F���&�>����'ZX[�L$�����k�`r{�ߪ�^~��s�E�?l�h�hI@?��$���>RE�d��}Op����,S��`�������*���-b�`~�9M��T��a��ud�!T���8�3j��Ţ�HK� ���NV\�qڋ.\�e��݌�WY!>�-�@5yQ�:z-�̎T��KPo�YGW�<_Gwo`L�=X��'��5��U�X�s���7j��e1Jrs�r���f�78C��x��6����T�P�#�F�l&�����TT��X*���8Gv�k��_;����
�vЕ���K�%�1{�5d4�>[��O�=���οm�66m��J�d�9$�'�Ѽ���e���=ǷR���^�ΓHTAf�zTF�(��O��*���+w}ѭ���r`�&�"����lxJ(2��+��E��wk���J���H�nb)|k���ɩ/p��9T9V�=� �oC����d=� �tuU֨ ]_��P�⊺h��D��_$�ܒ�&#��n�M�S��6ѐ��&�u
o�w���6�1�����Ƣ��c�A�b�:*o�|JEE�����]܁f�L��M�@*W)⤥a�Fϰ�è؞���%w�\����W�,v�`�)RxwO�|���m�-��w��'}�/�B����=�+U�*��C�d�d8Ύ�MG�?��CD�8	Є�]��=��M�Ս . /��,�8���p
7��<����oC�qB��+	[��W�2�ߋW|��%���bSޤd�o��]E��S�K��+49�Lz�L|(C�(�4��o.��-�/� ���f�G�[�4d|Y�(_�nF~�/��W��_���m�[,�*ryos�'nz�A��߀�+��
�盧�YKԚT�v�4�������Ѵ��f�=Y�Y�>�dQ�GgH#|m΀Dz!�h��F-Hm��H��Dj���W(��m�������-��7��~x竪[��V���'R���b��cZ�u��<��S����N"R��@W�RZo�Nx��E���02��4sR"'̋W|T��w\ߘz~<�A�ɐ�0��ȭZw�r�ե/3{B�zJ� 	; k|�_WW=�1m�m�,� �)\��Zu��:ȸ�Z£��R�(�#�	/�h�������{��ϑP�={��Sp9Ō�}�-\�~|���0{?"�e
�"�@z�`�.$^��a&��}�ܺ*�V����i�)h��af��R�䑅p#\�$ہh��r|)Y�I��{ZPD奔����Db�t /0�p�K�?G�ɟ���F��[u����"M�J�VS!i9̿쾚�J���cmK��g��*��V�Xжqn���^�A)խ#���c��m�2�$h�&M�Щ�ܱ�R��ũ�k��-�����X�ˆM/r���V'�����.#�+V0A��2X��y	��tϥ�1j��k�P"0mv(��x��W����+*�Ndi�a�,wϕ��Z{�,?���������q����o��*�ŽbӶ F4��v7B��;7���uv�WU��*8h�(��޺#p����7<�I��¿�z]n'�*W/=.��@s;{ѓ�P(� �`{8z�z9���K�1��@�.�K>���v�3��X�d�1a�h��	��3������˚U�v�
O�l$�Gve`|Ĝ1��ݼ��#p}W���hw�|��8ԲU�E���0�&����%�5Q�O��U����|��.�U�c?�A�����^�>����3D�(B��,㣓�+��م"}e�0C�}�Q�Js=� �V������ZxIK�R�j�=hD�4���0:�_N$bC+��=`�&�;X�����mV5�a��8��K����=�_F1ۭX��4	>�e��Z������Ȳ:r��a�ގZT���R����{Uz<��ׄ�?g�ݺ=soi��C�Zj��B��nD^Բy=�f�����~b��'�2zuv&�=��b'5Z�yH{����1�4�)Z�D~24��49�P{^���S��v����_D_Ջ�S|jR�g���P]�H�x(�{E�ʳ�B?[睶�
���
�I�+61���ŰԄUqiJL1d��0�~g�9�	�h��c��3�QgycaBʀ�cBũ换%^�7TYv<m(Zd}����I#|��ps�#�xͱ�
OF���Z�Q�Q��g������>�0#1gr�\i>ُ�|h��Nɰ4�2`Ҕk�Sh�b�;@�h~*�6����S��2����7C�o���(���j.��	ƍ�}�n��|�a}R�?J W�u