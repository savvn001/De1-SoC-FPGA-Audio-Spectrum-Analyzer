-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uBGQLfcxvpHfZrsy9rUENu7p7oGLo2/XrwO0K8ThNNE23PTp+v/TNexHVmWUSq2STAyP41d2s1Yg
1W3HmvEfEKE6SfOgYIizmkQoQ0cLUGW0noktf8etDhftf72wwk3UbSLhaNL2mdUXzAVIe5PMCYer
ZCBhpIZ/oVwqE4oIPdoaWGhVjodF0pDrng2mGJR77cS72eOse3RnpMDGXYoik4b7Tn0zThyNXIN+
voL6YsbR7KhHescVyAOyhl7yQiQymqMT/ErSfAwHq6jrJEYWjuu3NVi5BheVFO0v9uHcj4JvZAyn
IYHscWQE7DGoWaX2livykSzLhcBWtrWIHy1saQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
18Rp9u4N3igcTF6CxBxwlm93uRwUnKLUQKG4XPVeqbMo+0MfK6pmbYa0wOSjX5hDUyWw/lkNL5Uo
jgvoSqvwk7AN9NFb65GZFfWC+6WhvR3KNcV55/iCvt5LiGkbQZ6+mgoH3LP6sa1FdhafPZsXJOuM
ERHOf9LoZ6CJcOVlO8mUI8Z52qpQvvcp5kg+a05hCJ+uzBc53HwTIhLvcksQINQ2AyEtYhwuJjrw
5CRlPf+5jB8HgdMu4JsA2tps3oD5w/Jy/o/N/D233JCDHUnkI8AyiUnNAhArrQYiv1rEowIGRI3N
byTnSWkDiFmaiGGm4n1ONYOs6MLiNyWFBI7MlLHlH85S9V1dhbHcIjP7mptCgqerF8MYUb9QOSHL
ydaM4O5c0An8naPj336mwFVJ1jhRIYsH1OWbDWxB9OUVDgpQP2gy0dVIVf5zsNxIfkt2KvieFeB2
GrKwDu++RvyFM085nJlzpQqd7LHml8O7Gb7fLI2hPjGXZ83Won3PVEq9uN4jR6tjI1C9SS/BjcMU
J+NKeNQRH3JjHzUQwk4h/ELbRodVzu4fVxW+I5XF2y0nuaUrecrnAQ7f6/egzd7GlcImffVjSRAJ
ZYs5uoCyCXp2RknqXjfYug+A3zJrFTduhxQ37cHP7iDi2EZqM70xDhOoFPwh1MBBM+nlzOHeq0iZ
YbjfwcVe1sW+ry1xWIHT5d/xwIpXxVo9fdwOTj3I/z3LbnyHzqQXROixAWukQeun0niiid4bCief
Cv8ysc894A8ELZycuIpXVcQsKGWzD4vqcWceW5CoWpxKO7tfaOeyxnClhUq4onqL6Ewi6sOL5Qcy
Qk/RxXNc7xTcq88+mopotfJBmvZO1aRk9j2J1gDn3IeWpv+8D33ch6uGqzI9ZzlEfFaj5I0QsLVu
ELk7qU2jKFIm+/wZ0aAEvmp80f/oEBm8rt5moEtrtx7xS/5ff+854ln1NqhCBU32yWmQ1K6XmObX
nIr3Ba3iuHcut1ZYHvgEgO9gJGFfkV9zqQM8+Bl1YWh3NLAUmMpv9ojRV2i7pS1i+kWNfowlHw1U
5p1miICOPHo5mHG/q8VlH8daET3LxvDZ6e7YDSGzpes4XzYzJ6b3rnXABWm9APnpBkVrZ4ctguLf
0bWLHwKpb1BW5W4pGv3n0i4o+Sn8IuokBcuXX8m3Qr5NjPzlxdC0In/RWPBLzHc9GM1n7D8SSiXj
zpQcUiXbO2Xtc+02jOH33GnZDw9rwLoBWYzKZ3ArgZUJFUbusiySs70yIwId/AygI8Il0bKY1c9W
13s+EamaL94cRJD/nXaxDSwrGI6wDCJZKDxg48NObK6UxGIaSQDeMlGYvOZlx8VYXbXXsa4lynhv
cuL/KDRvNpBkK8rob1C9Qak7x2PxBZoS/T2ZRHb2+s5e7SFYZXQNMB4vhRyO/2ePPxO+baiKOn0E
aqXg3HPjoVIJ5+Q1fr6jg9BOgjXSf8clIajb+eqeTSENtIpaAaKn3ld31HiLbXTg1KWq7LLlcOqF
S7nNDAhWx2PcwavChsgb79QXBkN6RR9CV9NdmBTlGjJB2xMuhfxbwgtsyuykOfJKnLVeur0ThaCP
atdF4I3wPyv19MgI6VkCbPrMNgVBHW8XSe6leOLOFk/2IwyxCmxSXeO1hE9OKyh0lrKAZHEp4bsz
QMPaUm9eVd/aNT2TorkNdVAqRO+2njWxeakz2VBClcD+pQ4LpZDGZq2t6AbjN+AYt6ClTKcg3lsw
JsAvtiy+MSO4I2cnjzCj9c5FMEYyXT37fdnEZARzQO7c/dOLEJY0pn2Ey/1BZJ/R9quOBvpcoV6D
wjDD+DRLaHuLORnuMpTc+Pii48yrLGc7KdXW5DlNUsW3qvd5r3fSWcy1ZzdxjXKQtCQnG7immp7I
MPh2kDFwyA7Rc+QhkJqlOWg1CLgkimJREDj1avw7TheoEhc46CAVU5NUDuwZw9vx/Vk37vrmnK1O
MnRvvok7K2ajwj18LgOOkcrX6lTx8fpKfUcB9TfjNKXHmTlzdq9WYZoG0mYENhef8SRDpHdVdnze
nhg1RL8q5Dk7vqTsoWjOBV6XA0X9RqkNKWZO/aD/KHfKhTH1XwhWn1bZ1corRaZGhh7d3u8SUY+j
xq+iIgso22Dotn+ixENuiF8Ehpb1MPK2w68x0W1yaIdXIJYAkCTM8o9A8dOX1u8NQT1d6sDNz3NX
aH/t71RBcc4nAfhs11GBGiwj44OQ+rFyOd+e2GuRxfBta/T4iqX/V31IgaPeRLzdB2+I/JLxPK1H
DZfuc6qW8WdpKZNMym54Yx4THUHczjlrkpamInit4oVzWC6xSUajOZw4wEY2WEzh7cPV2mEqP/Ep
/p7u2BfvrAD3yLHbhEJrirFQn6W7pJM92y4fo025ELiiaTzsJzPxzrmr3mvpRMlkma4ivgCMhFjy
RIuDLBsJP3h4w7iPEiNsy8Q+lpItPNnFhcL7YIK86rNdU+fJqjFkTzqSeXTOimEPR2wTG+QEWtgk
NUQ1mBhUpQkS1AAN1/H3Nf9n9TZYDjem1z5cmRRk5Lpv8WkNODbRkekl17R/A4AT/65jfSGLXBmo
W3Cb1AY5CsjdvI9rw5vKh4spCdneyB5EFv8gkdfdtOZGclE2Gn+7Uenqt6ui9U2rpffNHAk5dWjA
M7cxpU+3K8xcnd4gjeAS/WSeVhFlnR/0H/kAyYHfG//RHPIDdmB4Wt0VJ9kI7L+n2dJHVwL57ANP
Jsg4hJtQm3dUhcLwj06rA6JiUfkVRHsuC9vv7eLtSPMwwuQ8d7ob2a+m9AijoXsoGybBGHcI9/3C
sZDSLGDa8kZOFGPDBv1mJ//1yQTtULer0z0S84BidulEjFkQ07oM1prIQYn2yVtCJAdx/mQVKMvd
GfVsb92qJiTKxSQUEO5Z5W0p8u6Dg2I9T+2sqe8Hy+R1krVco8dLszZcz5PvmvBFlGfiu3I8EPzB
cct/pP8CYOSckAnNYyBt7DYjGnRsckyfl+92svC6LD2Ot3/c3Nxipb+/qU3GDod6jR2ajCoaLSsz
ttQo+ArFO6C9BSNSKALJeVOFtH//afUhWL8NbI6mLuzBE+s+9d8yRs0V5d3zCylBuKDGJ4d2JyNI
mL98mnPEAsKm8FbUX2IMGNBGpmTFwChV5mtzIlPHKCe8vThzfmgpFy+UnsusLytT8lZrHNjgkP8D
Cu6WNbbnJs7JmRa+lugNI1mSiHQ4EXvPHqneI0qoGjEwqGE+bOiF5P5wVGymLpAmWKSxp24GkqnY
NF8Vm1u0ymEBvXLJzMHuMHrFUSskjU+tMEb/fksJzclgvUXg1LtrXXbfbpzroopP6pDROZz5Su+r
EVfefeL32dF5jars8UrPreJYlMHf3L4a5MkVJfZ771Lshud/j3MKXmkby6MRd/fzhnOU55txYqUM
ZzAMU7XykAhSfBaJDgZJZ60D2Ivf1w9iKt/sOHiJRRT17B4yx7jLw/qOlLdYc1Ab51bo5F6fcBBt
1/j/D/gAAmXYpytTExVPqYPP1J98z3gM17Asnfozl8G0nlzy1B9dwQtACAHKj0ZVJ7wJFsQ+sMpE
8PMdnqDbQgwTNbrtXenCoEwr0Hd+VOMPSpMyET9m7qFZ1aD7qMJsPFPfFz+TNto4z5zPyvwh6nUk
gEaud29JK6JcVdl13made29o07dQCQKxZ7E0LqG/8ZEV/JUdjW2C7MFyuQ9QbsRyULRsNcv2pixx
Tvzz5CGhqfQhIlYJxjfQwAW6/VH3oZXxIzFMyO/KhYy/EdJu/DMB8Q+6wLApbX4y7QwHYO5J2FDn
VTV02+ftAhYxp4G2JGfpvXmxWi1pF3IeTeN6joe4To0f8JL6couwUUrH8xWRB3LcCmspC1KyXIv5
CnPKIlN1tTNS9sxo2JB5hClQZOHwZO+2mn+V9yeA/MPFEbnQvO65XMHq5l4fBatzGC62rxTGONF+
Aq0WrA/Soe7Zf/6dWOMD6ZcLsDtQaSK1egEmUl6G6stmtVT+uzVrjzc/uxkaYhyYfzJHzSA0BpA5
BMJn2SEMmDA9Y7RUeZR63zQmpD6RnxVmX623ct/5Z76U7YVoSInAmhmOtLq5jymVv2P/8tNCecJj
hoI/6TBJA1TPGa7lEr9/TkwjR0WYGBMzyDp+Nk7RNm0TMXIbGRH5FYKo/C6MFTMA0bWGSOtmGCfk
VMQOUfsc3HFxcH86L1AKgSuwyr3qKF8qytnmrPLN58Ry4bL1yj252GjIb/0bHSmFeIUnj20L0vMQ
e9/5kn8f6ErVnj2GPtp1+MrAM7NXGshW2Lqlx3TjeP23z2Oy/aHmXBP0RjPncLANFykSOOLjZHlK
Q6Q1UnXW0rPWbtOIFxKzCf89mzvs/qFLs4TgMZIj1cBLxXTCjib4SaWxehOQYc19HpGVkfnxDVCm
a1CGFjGZ4WYqmf/q+sAqV1phGpyZiAVP5ZL0CPruDsTPwZXpCY9Bs/Z4aymuukNi3KEw7EcwE3/g
YhQCFUEs7EhEt3z2eHu2mSg0r48lB9cqBfFFuS8bJrnB/q9XfGaCBQMB+sYGDxMcld/jAUhuDdAW
pxEAOSZ0z8Jstk1GlnBPfXEl5QmVNnpUM/9jw8/HtHDNdPsT0QMtbdvyjdb6HQlBGNA4KTAJSonc
QoLz6iKG/L8kS+Xw8iCF5ReqwLnSXjIYfNo9cYb1+z/yjjrmZrtsVsE+K+SNR0q3GljvsyK6aOTK
f2XtKK0wL6kID8ZZB8R25XThgF5DqQNjCR1pbWc3v2koP5MfRAsgRnxqT7qbudrPZ0JMKUab38DC
VWQtIEjsz2viOXxBrNWoC/hojPBaKtYi4Epb4T9/A6HbnxdWHOZNhTLKn9RcRf5UGNIFuUdZs8Va
7f/1bV6y9/+kon3l2djvMXHYXbBYkFPY6yo8sFduu+w26wlP+J61JOP8wHmRy6An7h1jU0icnjzN
tk+mEOYQdB/+GU5cv2bQGdKyI/Lz7JJxoK/MWGXlG/dkwwSauM3rX17X/qZFyKQHca9T3knN555q
8euVKB3X9nx2UqHSXNKEXKRTxBx4MPejT0oilqs6FQGT6HdphgjjVXjbgO8lWFkxtT/AjWLHK+SX
GP0z2xp10/EQN/GrduYW1YCsg0m8wVSq+DHpK5A2tn9uPWcr+jRfjv+ygobCfol9/C3CCGJCSjHL
GloYyte2/8ilyTf8ThakBfPK5f3AMvxzPtB8k3ccJIbhSDaSYIUaKIrsgDiavcI1NoGXMkSZdTR2
jbTLUUQyAfr70CkclbcxhKhIz93h9QEnR/ZUuuJJ2qPVpllNZfztjObD3rmosRQ6CyP+uoXDzT1x
nXHimYpoQHDyxNjDD3k6HEYNx0+AS4GhpgpPR1xaqbYC3cWmQE1VGbBSFiKWXwEbCVENscif5lIC
T1kHYNJxUKrgOQmO3mCVeSiGNl/+fBvHkFiB9O68FVrkhMbuuimIw6kTNrTxmxmaAU/BmazSMifX
TFH9zSW3QoVlTZiWaHBFMgMiBjcA8gfNcoPqsWecFZTLOnkVG4wiO+teV14mvyBiG8aaPruh/YyR
NZku0z8STI4QLEe06M3HuDCFV4I/VYuUIDGuWVUK+pS+2qGUcd8NrtJr9tRDf0gbgKW4PVWGFpyB
1UewMnGcL5iZwQppsz8hggD+kQ/h+ig2PXlBEvgYlvIdFk6V+Bs7xQm1B8nSO8rBQFRFXaqkRIta
RObKx//VZJ6qZ2Rm+OkASfberxyUwVADWxCdHALcgyYMRt3Ymecmsdb7kEVlJm8SfrZi3+sWMfHq
CCpdFVFwiYoDbnPzrekTC/jJUqsH+E3kAeitqXkFw1guFudqRVIRwItGHd42vrBghzkooTceVwTq
vxfDEEFbl9KCfcrf84TphErd/8z1MPk/XVPJRh7qB1z4ZB0v3/wqQE9mz2rVq5CF0xnogUmc+NWi
KXtj7MdohLxI+PlOVQGplSKXrPQxkZxIP6WwwZ8LwhprbELlriZvgPZfXJNWv6sE2HXu+Qhl+Fpy
5Pc9UfUqf+6ayMpJLnLiQfQI5MmeMATrm/AGp0hN5k2JkJ6n7fpSaYxbbL9QrSkqyJnEUHi0LXBB
c5y+Q+BiuiVtoTlxCkuHDie9EJ0tyqn5Hy1FuBIP+m0FHsxtyIK0zlkGVp3QNI4NAyAIU7pSfMuD
drhuY/Lj3FriObBaxBJnwKTLUrAOoUM2BkHTeUHOfOFyb5mdeszS3YF8HQD20/IcrB/2kWencW55
8KMB2E3Jgijn3u8o3wK704nO8HNn/Ns/hO8faH1g4C6QcBI0xGyKSQMJc/0xm2DRYEhIpYmAoRyp
vPXpkuEtO6ob8e+vObbypQnU81GzptKhAhQ3+4+0S27Q9O+6zAnrGZxArZZw8aexAP9MzvqRFlcS
M5/4o1yp40z/JYiMqs8m9nWLOFGamK0lKfucqecaEy8MBasa+3Pk27igvSH3C0iJ2tCXhSI3nVXU
zv81xutHDQ0NwTx/H3bE+rl63v6ayKs9ix3teQqwQuEP2XlsiiNvhwbcaMbybYHaZYe8biKLGi92
lOzcMCCgNQjLlww6hcDUw0zOF186eTNXfK472fV2+xZ7aajVJbrrCzh3deOPhwjsT0kaHGg+Fjqm
RE+nDHNIut448AYXaZhIigeXxsrpY7qIJd+1d4M08exTpLw2a47pX/BW7S//WdZS3HtaPqjhzsaD
leyGT/WdOFkDgCipeUJ8ZrX5+BcrgN1OeNFGz/+XbgkvHfx9oBTzUp6ds3X37ly8L9D5pf4utMgb
JGjumovdY5mKitsqzUQ1m+/owFpKIzRv1iwYB5+mFTHzOwk/P169/zeAY3ewFmVdk7bUoTh033kk
EV3tZ7R/ugz+U2BiMN/EWDBg3iN1e3RtLE7WtmayU83Wb0zd8J6lu0b++nGsYYr5jGF2uyco+qzP
n6T2j+wxP3Jbh7XizDyvEVEtuRdIYbQCYc3LxkwzptODTpDMp/TBxQONmgz7x5VgR7pb8ywghMQc
TqQdoo3zByECbxdBXdVQui1guHfIhXobyyRZ4XUMJkOj+YP6gl8XzzgCwBFspz734NMkOAPb0PSj
XcJ+o8EvaDTR8hZazYPiNm5AGkx4NJ/wz10sRXH5IWQDI7NHhmsqWl4d5wzkBjm8VKJK8ZlQv+eh
hygrwa339QrXRGGstl+1UIVpUCLO5KpfmvbYv1ZnB2e0NXgv8M/qH7shJDOIVSrOIkfBQvswqtjg
tg7h+LvEE5IhVGDLD71wD/n+ujKz9PWxoIpMbOXM9UznflLYaG2f6K16m+ep6PwVsubapkHUp6qX
M60Kyw0b21s96G8ft7sgiAolI9WcJNZexxiIJz1NX3PV6L5IF9fzDaPpTPRPxrMfffC1IXVwtLOm
4WMW8ZELvpTLoiQ6y472t6J8strTVu1JC2Ze5Guv2SXxHnJEHeRK+9j3JsjBZQfVuKZqLfzuTmqX
X/yMxh93SD5esg6d0Gxmn7QGwwbQkXTfJCklmLLNhavVz++xgvZ78as1EQLKqOJNunS0gmoBabes
vLbpRbXCydQxWhseHFiZwUEjxbWbXpfhQ938efEyU2Y3vBS/roCmeu75rvc/CGbdVX3c41FpM9Oo
xi7IK4R0wh23q5PfIwpn/6ddbGoz+6OgnbB4JcTaVt5f8cy/ec1ubrnA7A1RhoVct+xVu1vWoQMi
q7nXYHQR/40NVJhxF7qbqY75NUsw/WpjoDF6xOz8IiScT5UzuOMNi/E0lQqZsR8zf4LDY+GiF6Uv
cfihnZIalZXFdoqHhKvFWOjmjRsaL3vAcWMVXr2zb6mECXEuHMVCPUAEG+2kZJHMN3JUxxI3G+v3
7hpsty9j0EiLA6J5j1h3slM9CB5m/cuHzjabRi1TtoCrDitbgANjrl3zR5SyNoYoru6RZJkr7BKO
LpCGc5iBvERfLjv+voVwUknD2vUkeBsgoSUyqY6o6N2JjxusOIM1qT+N70I0+SH/fgUQigCQdx/f
8MoXlB7dw3OZ3aVlNJW7RRAUUM/D6oClAZgXTzIOEe8/w1VQ9kBgNtmPiKC9o2IDm3EWhROtjZsN
rIkoFICg3F6aKUO68Bcu/Eo9cHfDxW7g+h/m9tQ8wa3w3oMMHCVSS1JmZG0pGcKeqJIZ4uCILCcR
h/i40V2pfaylFsrGyJTyLeIxb6cbrsQcYhhohXxL3XQROGknAka/zUVtaQYojhx+X270XfE5vSfu
FaSKgE4ztz+HpW5wROrSwxIfETeHfcCbTBOkM0chVVCwRzIRG/9UhjghQxM8dvK/vXQSfxr/XeOx
7sTUy5fzRCRdgqeWtiK4svKbHrTwtp5YZk8tzC9/XxSk1TLSbAFywvzzHuLMbXpX51CjeBCubFKV
lAJuyqJy1IgVPNND9+qC8U+vPu2QStGiXwadOKBBvoBoercWu9kASlniqS44ZpKqU5tkAwFIqdup
+wweEret3ktTt8jVZJw5cglkRPW6hY1rKKrUsImRcbUtcCOSUuoCljawJavEg3r2zC2SsDVFjRJs
j1HmjFpnx9liwEwH0MLFuqGFt+rGQhS36l2NNpalej9mRhBi4X69YCh14HCZ+O+XO1fM5lbCOki1
aNPCzww34rWP39q9FhLifzO/hc7fD15A3v/9bgnHqsyEocHz7WlbBoKo3waO+O/ZhUZi9y79qkCa
CQKvinDc1OCF4o0+MTu+UpIItQ6XaVedkpD8bpgZVqPeMoIBxRhLHOiVa1h1Jd7DP6PDxdsA1Uby
az0xhSE5ztWjDCTWgd/lsN1TsZ1twpE/l+RcN3lcUzm1okzO4J21SxEeWD1kPG5LBL7nlP+ga4YO
cyhXKlb0wrWlMZxFzkR0q0Md78B55og8XTamKyulxZro5OmCqxkFkK5jmKg=
`protect end_protected
