-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Bp8ZKT2HZ9ufUomsHWHfMHdwj9+kgQqoxR4a+EjqG4DlOc7Pt0aZsB2IR3MrmTXIRxwF0lUF2hxT
6ioDxK3ShOftU0cr21NHkwyL+ZKWfB4ddLUmy5Rbt1/DPXS+lrux4U74ZBXqIHR5aX1Jr3k6R8+C
5lG6J3HCgSAbwFmnIV70Irvf0fm7sF6I3UlRANIFscwE86GWKZMWLSvWmdSifrC1Ri4Pt+Vctqos
DlTUdiJbt0b4gXWgYbRdf5lFS36mJu9HUEqK936VbMZH1Tp6u759PhMGm4ndJ+qkzkSIV2OEafqu
2G3XKA/L93D4r7Vj97e+iP1jttAWOQWg3zy1eQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
uo1vWw/Cb+/o1d/aBx7Kip4RaV2X6qpHrCGsZdndS1nveSOoeeZsYRkUgijEVZWDZnwoeUxXY2fl
w787doN6os5eoQdE6XseI3vAQstEmj8pbd6jw1FQEiXfrw/a+k+TJoZE+/BhsR/WELCyz+2+mjv3
3ULXJewdsgoKgG4IekeUYD47ohIEhyTFsBP1743s7QPr6jAkeKuShog5HZ+dywi8AgAhk6pUMCJh
G6M2FXzd87RrOG27AETaEZha2Fk5vOWUBme/X7xG/QsPl6FPSrttaei/gcNLxYtb6PaYFtdLOpLU
tuN0dkr8XLuzyhh2sEqZWPl1ei9zCKjUbBLgzlz1CZnSLIzQ/t3oSqhAEXOCpChvzfxuvFD+P92R
ZJ4FqOpqiWQ3g6Lu/Z3GQ5OKzmJ7N7o23o13XplJg7MyCXf5HQmuOhc6PSWvVb1x1om0k8uNLpFO
hE9ut9HGhIMZfmTmjic19r4/9OFGC0hTh3kLyL5AdlZtWJzcU8HTxkqqSeoJrBvCyeVGwxFCYt+p
JoRAf/7JRdJGsAKt5nhIA6+Y+l56XmfVbBqHraida9j+5ijMXM8b04lhm378GgSUoYZaTOylwtCv
GKJGI/nw5wPF/9C2qbBWpd0aaN06To7oBdh2dG0IbJX5tVx2/SCsQRxClHYE7QuTrQI+BtnqxFL7
qrJUOp4qCXNSIQ08asqnFGSjuOobcexeJ8o26FLIdSjt0Av1fTnGyB0TuzI+gzMV83dFU3E8rAQf
pmiiVZAk7p81w+7F1wh/14Qy7klOHHxQAf5chbe7VKxXIpHPsBrg9dX6/oL56Kui8u39XeXlSIyV
VcauZBL6JHFeLovtx3w0eX2ztX/IYN0Wmmez5k0CvVYaSYSQWhJjSIN1giEUAnCTdBSspLgmwGb8
FeG2Ri9pyY8af+DEn8yjlwywKz5mmcM4ruN7M4MJzlwzpJo9YtRAYLazGK0VDopASWeTRRJyEUwS
a2ihK0enEliPH8cAKQzUM/ugWO1xfhx2moOjhjI+qDL1sR0w7vZg3FBczJwKs6PVRWC9/uk9CQT+
vgzMyxKIILQtx2heKkL+dmEsto1nBEYz1ZKEAsPeQbu9ak+13L0Onmy4wc3Ox7xKctozV64QAYMK
AoTCAY8Z0tF4Gqen1+NtL9eD7IpfsL7M/GnRiLm0gazbhfpBCpgk3U89b6pT052/G7k9ljJNAlCe
9ikeDak05neQa7zt9ZxVBZmJY2R1ng3xKC/qpqWHgtHVm3EbBW5agzZDu1UDH/DR8zZKSF7jSdKo
zPgtLuTDPstrFZttYQ3IAqIfB59ppTXSmyGf0C31WcU1a8FBqjuP1ldQMrAiHQVfoJNiJkiPlBlA
wkNXNnntuP3hOZK8YSrH7qSPf5uiacOTLOFuR7GMNRWvL3m8j8xv30p7djBV7jbiPr2hnB6LOBza
GSfk2G3PdfPd9VGKyanMERLh25MZXtkkIQqDO0e+qZIOTkstHGuhPwQ15Fj17uhJoRP8EXeomxfh
y0H8o3+INExsLkRNfiSVeF6LLJG5ZB5w10NxLQqZxJKYrH8aOSGKmOGmpNmCrt6gRt5ToxWVV5lR
yI2wus/eyHuBSwgupsVEObDysJzuz5fcfkKhcFEy8tMrCLhKlujiyRc0KPuldDBci7Tj9IKBYDpX
WZhhOztPTBu339Zhz846FS8dDTe7X/fnHdpECOmtgJiMJmdorLGEw5+b8gdVKcr/IzITKau1eP4f
klD8JylPVHrMmVjPfnuGjIS4CgHvwsD+dkCQX/lw+HjNCD525gEqLCrlrKVE5CJo4CEKGAo9avix
l/ZzUGTzBgBblmQQmJgk5b47f/tbpGhqC4PVvbdqJ3aADsEUQvTLeyVa0/GhrwOkp00dpjZ0Inpe
b+5HisY0j6/wASLffbtZkKXmPCSED7509v85Tw1RpDfVQPzB+ZYiQ76KDc/944YLAPvdPEyopdfV
nR0ZGZHtiqaI2KfK+xqgiQc4yZ5L78k8Hu6pZx/y3K7XD3diiiD7S1qOqbT1/ulUE/sFEo9CiGll
hZ6iOvUuamSs4MT9blpKrF6iYPD0BsAH5IpU5gJQN6MM4sYbKHxNgqBiWhZj/cPcmNtjXPABilj4
lR0PG/XiyvZk2uCNpWvVA35ay8Wi6dcMF97y2ISTr/425gMPw6gVBtiDXsPdqYics+kL+juGfrUg
JZw1VuQxGqC5ZZZpsz5Dfdm9hmQIQBgkSjRxrk9SGMJjeaRHjrOzuVouzB0huvpGjqfS5CzCx+6j
i8+9di94FnOeHTn7YPii3kn0gQLAsMB54f9nRarIf6l+jnL1IAdBjdjJqPUhpJWGbKdc9v53pazg
zW1ckfWKaHYlxSnC3U9DxEauNTvUwSvMclRkuaY4bhpf9rMzkPwE61ZZiJYqbsxCuOVhAV7T0L8l
n7gAz2vgV9nPrBpxToQE0GJB2B1LXAdMI7HI56P969Sty3dwSSUISh9BIu6a8eAulsSrhj+RXd2u
ZaT/CMnb21blifxWSzR1oQzuI51Vg2ymlqY+2pmEBOmoSPUGudwEuML14qUlPLZwiJhTmmpL2ico
XocvFx+Bow8sJp8Lg1KH0Om83LbpIRYw/1xVOYs18+cAzROTw3oX8h5D3goglVpJUceFK8VVHaAq
4/ahyK7CPnpV6RmmZ1m1B8PhhmenXXUKzQbCSwl3IfphLOtcJ/JGNWs4hcU+TR9bMkJ0TepG22Fn
q3Sks0hnMPZWHZd/EaO4lgtaoT+ZNniAR97/K6FuzgKTzFPYxok/iGn0RjM8XGKEqtwdXJvSNRCz
zDnLUni8n9VAuT6pVm5IBZQaC5jwUQRkWYoIKMqAkXgXRMspuEMdx/3608TmUFE9OB06ct7EKD62
REDkzbxmr3yuxNbxF/bUKPIfpCnrJwycgVsGLXIVhOmmO/c6/PSfMfuSaUEOtVkerOFcW6xnVb+j
XGQ05K38NbfwI7nSDmhE1ADE3qZljrbzdWFMpDXhTWAez9yhkQ11QABN79NXiLEW86RepEWJvZeg
V+nDdLROU6zJGdmiMPLFZ5JH6Lw6DKHEuH/mcU9+8S3LhiIzGY0iS9CPqHe2F0A33p+EmjvalZoP
6BWlwCGC3aspJ7AWSIihDaoXWtc3iiPtgkaxKMaJR/TT2VKPKj7RhtIW6R6S3bz6e6nBh0qc8D0K
SJHpXE2c0oUaBKLuj4VpjBs5LV+/0pqVqAiHLfYfDNxRdpjLZNjWzP+YylhOOQZIsfSRsD6pcoPd
L/H/uSxyGkOjXTbVgzcdhBRybPhoCtLFnKBigxthnCQ1/tQ2fZKhaVVzeKSj2tuk0f+AMovWY6Ez
nqU/JKJco+IPbKVjxgZEGXdMk/dvudEBp8hgk3FxzKM+VsoptMhAlBLx2oUU6KDqY8tF7TkzBIYe
YzMYRvYI3U9TxIzO8O5UqJkDrXXEAbQpZ+/fMAdPqeHR2SLUNhWUMBA1TaUOWB7hdKDKIrldFSa+
qtdTCBZGMnbgUBp3c/g56dRIIHqCAUofzn4glRbBOKlX21z5jT9k3N8nGfcR1f0AQQF55j2Or/M/
PV0GOfd1knvO5HuLiykipRLb0O9+YiXjbzoeubLO1YT7a2xsOwXjq6pc7ryvg5BX4jVUdw1SkWjA
Hx3bnou0IaOBSyNux7nh6714h2LN33BgNeSoJkknFnOgCniY0jeObj1vcM+ttRhhj0NX1mpKITPr
OaDyV6h+WJ6E9phk0wcSQL1Xd2ruVaqkPf+mO3Mjv3Xpm0aUpEbL37HL4Q7yHVkgAREaY6f7voYn
1XeZrDQkFGg0wxLSIVMSyJTS3llyt84HjwcKmxsx2GfhBv/Npks8Taoo/3jZxcBCU1QWUhH7q1wS
W6OLi2YafE1gzJ/kfhE9mjw2FkcUZBimmMpKUyluYAs9n6o6potekj7Pq6BlaqnVjaVdpQ+QrNYd
viyfJmnhU16D1O47t/6YMfl2svxRmY2i/rwlKltv1HAad8IbMZ3qw3DpzWFAUEXb2MJHSmzuC4CM
v7lvNHz3A5L2o/+WsI1a5vMPkaiKVuO0+WngkpxHAgep5ZyjUQyrtMoWqQiT6EAb9qcj0kQB2P5d
4weZ74S37l86/ofD1562HN1D8kD490ba4C7V2QdTxGGS2/tnndcps419mukg3a13AOJbI3zpWtlj
ns0N+ttiRymqvqaPsVxj4t57UEyiEw+EGe4LDLKPCWTcynqBpu8n7SXzcBg0UJZPw4VZcSjyjsDB
D/z8q3C08ElcLIw9hst+GVWlEekbqrQ8w0kOJ5fx4GTqPZGCiVr1UgzmIduK+gJi0+7lWqks8Pyz
LAXi8hvAqkriAj+KOWEmh6LrUyhZiAtrjFtZ6ba/37WInlytpRglCeREe8o07vnLp/Skwk93jLSV
8+KjKE8o9gRcAVh/t6l4jDLXeNQLUDvjh9UZNY0pbONtOzz4PdS8bxE9uzFGItdgIBe79FOEyGR6
gZt4YrhL6ZrG9vhcrR/D9Mg7JmtNPTMhzHvWG78r890h3vbPBE9ipN+wlrlajwX/5v7AgdAEdKaZ
AkxVctoI+m7rMTqw+ARevVR/Ox4CzqFIlpsJYjyzB2Gxey7b2LM+JGMdrDtJ7K97vBBSmN5Pn47+
5wc4kqwDAUXQkCUutOdzTGkHd8bEhiiP19p/Bpcw1e84HWnzrw3myCAz3yPp1s5P03mhi3jw/0Gp
hpalIyqBlKn5tnhALGrHuL2ciTCp+tXQ9ppsCZYkK1nKXXRY/1GHBeZzZ/uVaczPjAlshjTrhdhe
TUUrubAiLp7eRWGbdHGM4j6bAC9V/R3bLlQYOpriRX39qV1CY2a1Lrul9z9dgDX+osRwIBEB0L6b
QgLSD7ZQVxHsfvEuRqj9ZHVHvjAjLHmJLK6V+V8asHfoB2ddK8UVKuPuUyh4pcnFJsd6f8fiPkmT
x5uphhNoylyHbzPrICNT0FJgEY3W/qtGR1/b4Dh86VSbT4Y5fw3Du66keToMi+0hSMOJgkiDkw/e
Di/kLWclB26KHlgQOyjp5/LjJwNQjKrtmf5XyhvFMfgDBkb2elar83uG9PxVAEaSdP9OiuaRlACE
J/8CCHtdUxn5L5UtlrET/LvazpVFs6+z9/Nqe/I2yLI/WRmkYAtv6TfuuUyo4mOntW6S8yXawFtW
2YGfEBiXuUoXgQvi/iz4/mEb4FLpumaC1427c04oySCC4/w8IRKXA0wMuk2b4RhVIw2rkGgClCj4
+TSapOJk3/CVpcAj4V//pmJ/csKGG0yKLMe1rjx9gWtmeoWyK1HVMBi5FkSqUqpPKXLC0JkVdDr4
y3asY3YbVMz41yAk0/jbl/fBe6JeN6OT15hy02ARbLxADlwbRU6yRHSKV6i5VtRk1tat78MxmcUC
bATo81Qem3EORG2+TNMvcggcFLOhurlVP3OiACvVCbV4a7UxQURm4rHKye0cLgnIo9Zy6noli+Fl
ZApc3ElF2ZNK2rqGKEpCph0YTzn0AfcewiOny5Bz3J3HErmW9kwOyqkrEQbL6oj2K9iT0jSbSuRk
5JFDNdtEys16Eev4TYT8L4a7nYAsXEZl6x+C95BSP1rWdYAccgSrZhj7O+IvEiTKrDJbcHmgzTOc
cLYVn5V73T/wwUq38HmTxbr9uZwbuQ0nBjkOb/VP8Hm3ofhcWVXc1M9fOUJZxvCOJo0MxzrqooIL
g+/TwoAGKhpBYtpomU7qgQ4Y/M3UdcQDUmPRbTc+hA9KfK6zFg2MsYHXLTQhMMKJUySuf3MwFXgm
C38X1wZ42NnjnxyOQnoBIQoPseOIZgcuhQ8x9zHFhPIEXnXoeJIdX3kkBAaFu+LEaanE7UZSj9Fj
tovi7/aueADNTjLv6bYZD2wDTZOXw3sL96VtLrEXSszDTlnmnHur3mlwVr+jQGVXt7CED73u7gPw
UmxrOodIfqmeVuqda2dM1A9lkDVUMlrJYxaSoSnLP/9nXja2z/FPm8S63fAgnA6OmbbTTRmQDYZS
7qaujn1MWNeTAAkBdobO/rKbGSbqgW9j9fbm+21/kpTzGoSWsbnNqGI8qs1Ivq66e/HjgFMscGxs
araff9+Qfe16JU0iRZSvEY/0s2Csb+lrZz8ZIAdEXVr4/TPKrfQhnD9vLN8ybYKF6nJVy+DQgCkb
1P3lMRxNvqWwAH8J9X/iBxHIwZVwTdSuB3sjDD9q4Rhhr5eG32H4zZl9GPCeF/5u8Nt+lMB9LTyQ
WLGngMDJgapMUn7yLZvmG9v/np+vThY6OMjZgWJg9IlmzZ1Ag/Ggw2OIHL7Lne92+lgSVdClmJS/
rhiJndEfTE8GWUpWRpkCT4VKZ9Lbcxnp4+dOwgLlOy811jsxKydR/gt/lGXi617qW6Uw8YcYQLfL
euanvOEc43JvMmJSp8qIkqz8WPuQMlNiOQN+8ph1o4aIGXIlgUjLdvBJWBEpRJRAMCIenvy9KtPY
Ao0Y8zg7PqKRewac6BaTcn9vH4wI7JWZKKp0BJ3UPoCGgLMdAWfFiPiwArJeI7YyY/CduX1zvQ3t
YiWG+ObV2/Gu+9vXNiFZMasmyshz7u82zBtVtm2w4qUrtu39lkpFb6DMYWHrOLNl9ODheQRzuWi7
+ziYW+uh+MfmLeMz0fgXwSvT4JeyXZKq2sisJc1UkKhHxqBbTfL4K3XY1Kz4V0YRsaM3DUfdRhlh
96voT88b3J43FRQQg4KTJd3Yg37/EqiPhUpUkqqdEfMHavF1KbrkMZIYEPr56WIKrBYZjr3Z1CNr
qo4aI0BrowbJMADEuTwux+EaJ3LTkKm1ZNkNI/OXSceV+K3SHFq8/SmLsUZplBs2SE2q5/v1AVA5
dTlJ/bV9h3tDvCi8RwMCyxFYhLngVRfQBcAoJeYndsNlDR3OF85Q3J3MPocsPPEiEh2axJVU1cbo
njrhGteSjomYTSydWBjr24WcdJdWMIByfbF0I69l2lCPzVpIxr3HedZvXBrEb1jr7rMJcg9oRHE8
rQmic5JCK9TYSSNsSOKPKY4Sybh0sv1mSATgpHKUZjWo6Uwi5WLc4l940meV5JHQbwTf5PrU+xDz
VOI/Gemj6SJvhcLdA7X5Hvot9/a251JP/6c6ovmDFbYqqV5sxViLd81QtRRterQS29/p141yREIm
ouGmYcGzih55wMV7bVp/TNTEbQvUzbnsAVpoY+wv6U/CTvnBKXVDfvN+sBTIcwQBcaDx3w4RKwTS
YFnod2+/1u4n8kc8l36b/FSdhnJO698uVVYZgbHdj2fuz1xwAqjqm+HxBOIjVC1tLYoTpCRkkpzx
rqY3ygxFiiXjetplaS/VLxjQljnHTAdqAEzM1wFUZvRZWh6VrbFVdpcwvpdit6ZKinlc0Hp8NhK0
UYtAYTfp6oo8pAPd4wz7RXSYIWfy4q77paYP2pYycaOEYpb+Yvqofa56JxCD4uliGkM2RR1A6bLA
R6OfOauIV/CK9OzMU+RkFSWCyqOVK7mOzYg1mKW4mePNQYiUnNd1RWXCz1q5dPgJi85MnBpWjpSN
hH9I+fgeM0Uxd1xNI5GGopp4xPiucQsv97KVRPOLkW73f4GMkNHEpvnd9qmWYqMCygbmU48tecDb
pEtH5dFd0pfQ3+QswJjGwnNNUZobk3khfs2UBu/sPExqZ1p22tQ+j/R02vHEsk0RaKSDtwUJrQmE
uLv2TNjPfCdli2Dhr/IHLwMv085IZrVOSz8JKI69Jdh/XZW7SnFZOLKUNwBOlKX8uLd+Y+EXJOLz
gKuq3/zQC5kPCA69pFjBPN5snz4q0WJkFBqKl+Qi2R5raeaa/UOL3zsRerAUpamZBdTXGf2BxEFc
03tC7ERaCXC+7D1aXSnZETbJA3Hwm9ijyklRMwJnvUzDgqJ/rO062eJvgVrXJzDiueEG/YBQsQPR
NM9xKbJM/+bw6K/6Rag/wiajqP8Nhtp9W9lr9HvbDjPRKEKvXmIezhbNQSs/h0knOq/OCi9MriXw
mvkOaRzeWX2Ba3mctilCfVWmfkog2DBA8NIIFq4yMWfDY/8Ky5z7PecUw9jF9tRtmOu7E/yFTP04
nDZoeaiseVh0to9zj/lGBeoRu8cRaB8tq5XhduGE3fyNeawcu4Mb5pmXsdHehT73lMi47ANy5ylm
LzKc4o0ly361nBBsgMWBnNPSmthEmsRS1g8BwwUO1z7pzfEt94I4N2DFYWzwfLpcL6k1c6BtW3aE
FLbCOQwMHuf0Az6iEWkarjLYZ/5wexIefCzuTyoe34e3Mg37yaCDRPf/HeCZ/yraCGkMAHZXHqJB
V+HB4BkriPdO/wGaN+Tgf1zT43f121dySh8KtP63sLqviTN7PRzy6y7gB6TfSs1VtVMrZQK1E0xd
83Otzok25pQfVYVBxoliJIBKuj5m9AXuu6KSfO79KyOuO1B5HxzbZE4ZOE66yBFyoWZj2LUeqMW7
X8vBR56xR0B7Fi21WSTIyPqOlygt9ZHyjXjsW6e8fQrgfCgsCykeADO9HmghuFup34xGxn65iw9P
BlHXNKGFHvuuuks4EJMZ12YlQEOgR6XLyjoWa1Ki7CNQnZk6cjeYaVML6IlMe10tqGGf1KfY+fCR
Z/+qHcid8viBucLYsDsj6smOUpVvHuDL1REHT7MiXDYE3Gk+SK9mzvfauLbNy/PSmXkeKiL1hmxq
wn68s0CBC0m9RkcLLJA+1dS7CuVUb1xzDSajipQcx6ZDHZwgjk+c2XZEvsv/Zgk95RCcawUFD0WV
0M1FbvVXrdM0bN5OU1OLzQVzf2ZtMv5JdsJg6VSW7i+xPShJb7M2ehVgEvJ4AFMrVQFrENB5v/Jt
IM8DqBjHeXtPfhQJAgi8XAaQCXZIdrrf2LWQ+Q9aKca2x6oJVcUsTnjySY6d5t2Zuyqj7wkmYwS2
2GYKy7Vcte/Mk5ftD4j1ZQMB+Bfw9YAEpqKmzsfr2ZiqgPDXxc9Ah1L4yBcAX+LJ6UTtYhKjyF77
n5rDuTM144VWc01ewehQT8aaozkQmEdLuiB0+sxH90Xd8SBoCkRCIC6JnvodBUIuyTG2th0ylHmT
5F518onfqOMnXZgv4ScDSN6Z2oF1cFpOI00wWHkKcS0Ddgi0EvEl9ai/uX7zpOZkS42yrEVB/cSz
tcRh3wrwy06bvS6/VyouF2z6srACPTF7SApmXPQzpvHt1wRlp1Zo9jPN1FmXSPcQYK0/sFIX3nVm
gGFqA+v8nftLuHdnDPiknB+zkGsl2+yBL+4kR9snN+VL/pUVQM8PwEcRBWYQwDDxvc4qBTupq9l3
cu97tgJeE4swY6g/CziExQjsmvaCaAsPcOre2ECaVrC1YCpUjnBexc2+ZKQBlAgkj2lUhGX1DJXF
7CCcBuORsOP8KMhyd1G8Bmtb0axLyYdIzhfjkgsn/6PJrR9XuqZRsFOIKAA/JvWjY4j9g5aqJfWk
FLCg2c7Ize86oy4II8jMl7/l4nRSkxJ9qGoffbOTa0CItVkpL+qdiDpDNcwWWq2cMNRZRz+8lgTn
GkeTMOBK3viGjUSrOVCTrjl/WmI8PCfLPPvSKrml+6xgvazbcEHk3P7uD2VZX6I3wrfv3BTT4LXG
Wpa0EV00KHMIm3SYwWWGGyarBlmFk0isFZoioxWrHxK57IjJ/Z+ODRwakgHbvxNGSSYeQgLq/d5Q
KeVX84wyvTIz1EQq9ZcOnGSPENHkxA5gWVf4ux2gl5Z1VwHB0VFGOxOPcurDgRCiVYmZ667LNXND
omUQdFbBCPyC9n93N0dxPHhF+1WGm+MH2AFF6EmeXZgz16j/IrrqUg07968w2sjNreGxWNwNUgj6
LIQM6rlbkONX3J3i/4/R4qlPUh36xX2G4zCtsTBf6kpFE2JQTHuJMO6F5xyZl/NYi5eDQga+A9iw
MNdv7oQn0RttAnvilAjJ2gYnrZs1Md49np2YxMgatSpBNHMWO0tT5m7fE/2vPSH0Rsylw1tFe5Dv
ELl76z+D6LWY46C/VcErX81N0puE78OpuxiNq9mz8ZSr9UJLpQyzjQJIJJw9JkKNMWz+8RVi2HMp
iRpdteoGxcgU69AzQxWBUeaNNm1V7RDq7aDr5g385DeIkqTvTQTJOd6hIaDHq38Jtb2euY8hZopd
sxSy4EnVAiCqeUIJ4/WKBiOVm2lvppujJnlG34CJpUUXGJDsK03VnlM+ANHlRtrnKpGuJ4LkCO+9
g2ItbCvUdPa8PerrzIqOKNeoEQfh4v4KzHLXBLDxjOqhR66fp606Uo4IUkfUX56ZgkhzUiUM4aLb
dkXQpDMskoM9bCMVGq4XII3NjRiLXLiHk0hrg+BIUTkE3loiKJ1TT29tOO9wM4D9UdUWvnfU1Ecb
XRJHwGpwAaQpcpHuqTOBllsav4OWJshnwSgg2r6SaBwQ9bDOySeYzqBoU+dgi/TvnQm+wJTrhInp
V9CUDnnl/4SZh+m+Hs4dXosbIhqckfo2vPSOWWipstEYrWJCj+MceQvcPLk/rUUQwxlr5HhVHUvP
OfLMBL60U90J6YGA/syyKQJewlLx0/zkc59yDrC/JlmUlb5yjbMojK2sgxLnBqYXqsVBeVd21aS7
B6QrmGkdp15cose8A5Pk6wz0ozTmMO3LglZFgE/ZsTFGb2HDGRnOIICLvCpOI29PQ0FKU05NUhgI
s1TdUCceOxMNj+q+0mW0l1unGpz80A9MDupwZHY7Y+xAVZLvvw06VhVzIyh22sJHJPf9sV/y7KI6
mUKSO5ROGD9F2IMPs0uXVYVWsZxvwHivcaDvU/fIlDkQgJkWBtQeu5NVyE5btsMDMxVOk/MpfcTw
eZ3hb9KHKrlV9CtpL72jqOH/+ickYf3XcBOh0B9jKcRFbtyRIvkwNfnrM4SDAfeRazyhgSDvlesp
6b0Fz7vPn7g0Ovrg3dFKx8pu/XOgMtPdBQKgRM0//E698mC+zeDfEJZ1NhH+ch2o3/KBvVrHyvuL
SfWjMdjthnO1D64us7yGgNev8KU9hfQyXMJaZliJFob7paxJdufXK9hcQ8nD70Ec66mF84CZZbxV
UPbwA2ZJEQ6Wo1dXOyU1rHvgXK3ivqtgtXV4qNfrtL563BSQdCqoeSNfmpgV9h6STsLdeyj1p83H
Imojj/CuqO0igtvfH9zRZD59aZ17D/7fYBcGDjE0ejVoyk3MRO5oO37fEkgGT0JcVhQJ7Xiu9s7E
EM2vaFaU8vSRB9bBeDL9XSlDAX/KTGqKe4QPY3+kMRfpXwcCeApDGuDwfIFQxWdwTRep/06qFNRA
9tJcqD+sqEjkOg161ONS56i1R7JhT/8g5cvdYF/wt9Uhbv9ZC01UNIu1vjRGQVTRSaB/Ls63zgIk
QrADNJU8JODUvgJSuMPfoI7vrXvTj9QYMQyWSVyNdmiHt34pl0mXlZ6pj1qn0Lhb4o/5OsR52pWL
Vqccn5uCsszw1qu8YbknmRsj1WaQw0BKtNWGrZcPKx+TebGwS3F7Pb5wv3hyN8odjGazCmA+rk6Q
1ISLigkNOLnG/1p00lSbu0NAb7yXl0/fg/ZZ86gIkBREN9NLqlydQRd/oCtLtJ+nZEbJo0n+zHyb
yBpSlFcw6dYQxBmNvrzng+oxa6Zu3wgJgx44NjXDip8MWH3evRNPWasyXIYrOb+s7IYEgu9Oi6tH
7Zzhx+wDLYnCt4uX0A6oGTMHT4881NKos4ma7qjtr+zehhzNET5ED4CSqBCoe+1wf33KjjUvhhoD
47iFkj1jRoQFs6Q8k77wMn6BKwXB9mK5BYWLV5DnxfENATb/D7L3RvH4bEKTSrRLvIW8MYBW7ys9
vrIsNalFIdajfsd6cNR6IajIelsR4WNTzzFPx007j/Qh35OKAtqLHapIzeB07oXxBF90kv24bCRf
EoDx5UpBISE+3DRv+BT43qUEQEDGCFE1CITJZ1RMNR+ajHGxrecAVS4cSPMk05b8JFAFojSzIcV0
OBG50PTrsQw5FohTrCVRwA69xPMsgJbpt/sMAIw2y2GaskbPljLQ4GWcASr8zk1KThx7Zoyi6ECk
LYxaIWyIN8uKxW//WqfIQq38+sDH+wL42x7KXKyUeu9IvcHt2II7uY1/gMNi33A8YYCRd4K+qpcP
4k7ontnoFV9kd1AWTEsayNWpEm+fvtFQnBxZy+3FympF6f5ZPF0DozNYWJj1P1StopCpNOStFjm0
XlDcMrsCWtMtBqSSdlIfNISUFNvXlztwid/gV2XXlRjgypokYAFrz9hyRjxy3wYxqlS9DGSNFuPk
t3iztg7x5qa2Lz002qsaoZKk8IqlwZEBOnnerHl8ZYlzKy7JjNqJTfcJ+kEskcR5qmdkjkb00Q8v
tMcAtPHz4CKL7wEfgzdI05+f/brodXNmvtVV39g+GIoGhxU5grgT9OYR7/LcHVtOllndCyw2pn+O
6UEEqBmzu6HEULcJCU1LF89NZWhP0azRJwFmhJVyMK5BCi/S5peQMkM/I47qjP5hllLbPIgXptWX
GT58P48uIT+WLU6DOv+kb2gQtHKCuHXM8xSaNNkBL3tDjeXwk3OJsDaqXJ7rWw8k8UpzQzzfq2JY
TQf4qRSbtuvSRQbykbvJ6Cdo8oWh6lcK+/5NhbiTeaJe7WcI+xiZxGTF/jRQlLh4H+cOasN+gO3y
9vEckpUx7oAUl9rX5byaBQ4jsjGH5oMfq+X2hL74FwhY/sFuYCPb2n3SCKjw4UA+iacffCMgACqR
wUqtpA2wlBZLmKzDtOHKEW2HOWuPGFQxx8/PaPxF47JQbZSvBzarDqOgxfHq1VtXVfDCwvQZHmnQ
rPGIRAr4q57Ff5NM7BguzUanfOeTsHXCiYnoER/BafdEEh4z1qqDhnz7yM6cMuBPXhBe5JnKOWaA
kEjD52tW1hh4Joc45MEAAQDyt71x5Idi/TT2CGnBR+UprhOPY6LnsTcfdTl+JDNDd1nUpcps8SEH
JrsVTNQNYzJUt2U/TroBM1V4fzICFX4HzZtapkDg0TBSm8f4oMahQk/nQ43mh+ERRdCv1MCg6f4n
aXOsd2TgEQQ44sLHCfwQgVC0q+Be50wip40COvTP63ZKNzEqScOfQlWORX9FYiENPJa3EPOFN17v
wThPyXO2/g+hVi10n4Kc8b8khLsWnQjzTY6JTBdGEZJvNdbgECUl4ec3ePTCy4tmAVbDtmk9B1Uj
QQZxilFKiPDFpBRw/hCG1zxna6XRxqpzglzukpeQD4M/iPdOMgQvJgMvDm6UvamIQNoooJ3vY3bJ
ZLFfLjH9G8Y2NeqY7uLq0YGvWaJ06KurMBUCNO3jOgkQz1g8o+/zrYAhEgexWEaEF/fdI/B1IwDC
QAq8jX1vQ5/oo6Zps7CSXAv/sPPWSbQIS4wZwdpBeD1zUu1kgu9hkmq87lnNUyb8s3DlhF6V99Vy
5Vxe0duRGf5Lto5qVxG4qzLf60kXjjpxDU2F7kkSTcqh9tN1Hr0HoLDjPrG9aUr26rJt3q6y/qQ9
+tAh5G/wHJuItm8NWWLtemK+5WkLyKMWr3fGtbMyo3DQc6n4n1SwARvxCDH7hclOPzdc/oMJqPDM
62SLF+QA+rSEgcGTvksyFWOanP8XyNv/jn3cGpTf6gTegiPNGPxx3rG6cKqPRnh84PxdTtEiONJv
L9M7mwMdLZBKuRlI1VhLobfr9PBqH2YCnRNpKK3EvHFQ9IhkTfzLDRToEUkK5JJ6xOqte7tO7MHX
mqzrTt8UWL7/VxALV147h/E6X+f1QD7CmvrsQswosVqU7XnuOgHuZcur5a7IyjYF38QC/dqbejor
MHh6jmiCFRj5sJnrpbKShDQeBbD84SOWflErfVD0v0j6UPIy2EhZFAFny9btNN9Kx7sswyio2mjg
84NTVvmg0hG1WJLnyb46CrPpSLzIhcsCR0VXS31bHOKTYzGl/0A55THWybRDqXa31qXYPlyN4hcZ
XEiom45U3JWkpg0ikSXwI9ZzVhFyfMqaCSppFq4jJOeD6vhItfE4G/0hWv91wGewZ5AhqDrqoAd3
cslw3jMbFXUqSHWo1BYVJxZUI5/cbG8qBqSLnWNQoy3e0vG5yCrfravbFY0uZjdsPSvuIglihUFC
ZW83jNmgOWuR7peC4YVQ3YpahAqwtaJxtsKNzvgyAo33nW+sZU5+wbzvaXFJj+lc2a35uuUX1iI0
u2p1JOKg86X4jn8eyAwLt/zIqvIpzW4OOyQmR7hnYiNlHPj54o1/0jT6k9kzwGQVkno/RsiYhsBz
XdCrSHhfdHI0f/MMguqdvmcO5yTgU1CsGlnVKkz/sfyUL9gx/JuE56HRPB3aLUaWIekbTP7ogud6
sBZ0cxRU9si8Rc5pP3yebJmcWvSLw41Y6ez4GelokWJoCIwjKYIOWdGs3fRKoOhnhVNNklxn9W7E
wfZoKprcIyWdnsYZlmVgjjcLhban8lLq+PuE7uMcni0sn37/bbiPR7MZ5kPnsKyjdPo2HVmT6oh0
Ex4xjmcZ0Kv+AkNqFsz/rXWHMrrvcJ2zLBxDWbrtBHrV2YRbsQGt33JxvYemI+ketp+IgHE2jWnj
qFOUKLZuuHybtTMDJJ8oWyKKpEHuAsweq4P9Ng4lgbtYxeyt+Fy93FVSiz9+UMnSrESCLIQO6SSn
fe8WCqCUOCur5UmI/3v4MHkJ0M9BYRq1fdpWFgGKhgAbDZS46ymvZSj4iOKvLkJEKQspS+FzhqQs
yXcu1LCcalY8Zu9CNjnf56MfZt4fOFQiF1x8QKVS8l1RDK7oVcbssf49+KasYhEPGnoETulREfY5
u4Ia4pR32Yt+QrTXPcZh93eqSCh4y60ZK4YvAQjTwXcy0uFU8g/WGRpf86fXFY0vd3BqXUGr5yOf
bPgbM3yIwl+wS8pdi7zUGvQ+2iDNiR1WQLr90H21UeRC3+1ma7V6+3kBLxatwSz+2s47AR4Eb6nW
n72lNV3X5T6NtEAUTgXQRlNekm+cQQs+x0XQInhI3T99OnVHMl/BSb1Mjs64rxbI+ca5joOKSFp9
U0iHLyJRaooTjF7f1BtAdn2zOeE6lAMP/yj2TCi1Nvn4/iz1Y/skPBUUfeu3QHfVo/YRKvjvFxPQ
PCnc2Ur1Pz3XwnwIVZWRW1KcQVIS6eoncB1qelh3zD0fDpH+GNRbw/ISuJcvnQwkna13Z7uS25ak
BER03uiw15o0oCGOTnja4S8kW3U1Wcbw6F5jVlgHVRhI9lbZihHoXxSAg2qkFCz0DsmS54sizVqS
bxOAMlIQIZL6HK5oiMCcjlhPCwx7Vuk9QXEc6YzK6F/3hTrTHNFaUB75PDJ2U60ZUAltjILLT9jJ
0rNidu09hv36LwnR4KnfWmd49UeudfmTKTCBuCutc7XHIOElwlMRyGgkXMDy91kkshDRMkckB8xV
gIc+pTR+9u9m8z3F4FPiNWQbuQ9f/0Y6zokMuCFKNNMvt+Y5kente4mQzZr9KZ2Qt6lo3mzUL/bf
mMzRBivDH4RmyMG1AX4tG1uKuUkF1P97P7swM4M9sgRfSMpnZW4aFUOnQND4xnXFPeIvI8nJjJwE
6xzmcpmx+JPWooiiYRsp9g2jOYeKj/WXXLOSWA4pwzqik0ctaV2SMGNDdWgQBURS75bWXqggehBV
5zm76OQDg9sU7gFGtLfndatOvnG01D9hJQhrSUJMMZU21PWBxI+VFyFwIO1dcB0wF+D2O8PViJyW
bT5a800GakUqOdhsW+8YIbKtUMtCcCdpBELk12v3H2vJsT1otpOkWw8rUz4Xp7EIXvQiZ5ZXorD4
umWyb+tPLA/+yTMAfpQW0/gd8yD6y3L3SjFs7Ch3eah4ihR1P33F8VSAZeX0QpqO2K7mY40oOUMN
z+7DYNF2zvh15ZZ/OqoPOeHrmiysQzRfah+HarQ+2rrJXIBEEFZ6HFd3E8t5BLODFFQndyXhkywt
EpA6iU8dBrXMKy4a5XXzbxWmknuP99Hlad5nHuK9/gPy7/WxRYJ6Grsbu9vTNuQP67TjFFFN6hy0
rhqwLjxUvYhz3RLcnraFNbK1emklOzbiGBNo3VUnMgrcJQ9G0bBhWrfKsZYQdEpcRrsz1r8/S0Us
q3olPRGFQ7NNuJPxQ8f769QqL/lt/qy2rjfnHkKzOGVZY3zvvR0JZvBOOdsepvgwHFf5/eUQJdv9
gHMfShVqcKlSpoufOLCLeQ1sFaTjeGiSzl1wFcQRBNQG5ZNLddO7RLuTuqncVqsJ8aBnjsKDJCcq
vu1YGDS+H+3MWUBVQOhyyISq4LEBjWXvCfq3kfCnrKaqt7fQJtn45HOt88c0PmOiWX3Fpypf2K/f
GCTORn8dvpSrqycRlGDrEH3gImekce56uwrv61SgAsvg6x9sPlOXUeXCHvSYXVL8289KACCJgOii
4Tbik/7obTFW0T322bdddLYIliu4n+PnKlUqLJ+YNuWugVGh6m1UZ1hr/+YOX5YzOhGU3HxFaF60
mEi2iI0N3AHsZCgda0/qn2js3APtuqZ5SODfR77Fd6iPgHmgnWzjQOWoIHI1tUEjyJbU5OfCvF4D
UulkpbEP1ZlY66XpJ0M0KlEHDuI9N8bHiUGPgnysH2JxEC/LmujGNtIH4H9P8tbEE2mn2Me31yCc
oW0MlVMN6VZeQUc2/hqdcjCGQQtyfHZO1ARTrukKOhYV0MPv69PkEd3pgvVDCdTWLOEF7wAYM/PC
vocKFGQyPuxEc1xx4B+223s5GU977LsN2cWrqaP3fB3jp5DPXP/aOMu4NRYGGPHAhh6yvsK5CLz0
nA/hzyEtQHatt7h6B8/lXiGIxga25q03PiOPAbZXfdykz3TJFI7/MrYQD/p3wXEjs7qCdOjdpGCj
JIZhk0gC5huRTDSbvfyPEp7oie+GnfiuDCBby54b1A/q7hhZzdmPfU5MMgyKnrlQVk7JL6n3w8fR
KyvjxJEQ/69oTB6MZGqSdruuNXsauZtQrXiZc6BZtXbeKXsSs+5uRNUaAMuabKbL03x98hetC7gI
T/CqVGefAOTZv679K5Y05l92dnR3jm2fYTcSh7kvK+czx9HRB3k4ag6VVn9pq5G6xQ/CRlkshcL2
ZRfL5US8JvknndPymlJ43kPF5+3CoJ8rHbNKs3ht1ILxfzVQvXcGSqmZGTkKEwUGChVKQzGsfX5F
16hQ7lIKeH282HZDJmiLDWf5llkzmDX8+M/cvWzsSmWBCTl5Qk37cqDfEtcP5hk+9tQb8eFW2xeB
CM7kSrCgMK/j5pEFQT6AA5Calgwr6474+VxVk7lWd5vJXXf9/QM9e9+MLsGvP9TtaZdY1UYYpubR
zr9t6pwhnVxxy1CljpxPHMsx+wznSFYfG4cbzbXz6/ojdkatM/3OrqmuZa0i/KHD7oSDyJv2qKJc
EHwj3TNAIWrazWY3sWIhUz6gmDp28AFyXkA0pB4CtreGp8KyL5aryOJpcNy9ZMkbFibl2hHT89PD
cgObLeviqMXGunpFxoa14r2hmhfbLM4jA4T7P5mvIba1Dg1hkVDw6pWqiEQhcKTbqn++8lFJkyXQ
7lE4VwtjqCAbHITkur96rQQbBHWej/HijP7n8A4pAjS7KgmoXaiqVC+sd0wz875ZNBz8i57wIT80
l9Z/3oE7uLYSHzVon/3S8w7aBA44k3u4ILwqephF3rr/6EDu5GG3pOTn83N25Vk2qzBzlzK331z7
wkjWFYBT1MFroV7MrDeIjvb8LRWRR+PiN5tkl34XfiP0i9uGVrM5E17kEULxrgK5OCVZk9H8L6A+
FinI0Mjjbv1RFjv0dYuLlQMW/5paZLgAL67PSBefYWmOdASbDTXx7OgPA9j1vNB7vNlih12Hgxz2
qfae5p4mDHwf9vjjQzXrpCasnlmWd0K7yawlCT7SzcGRz8dX+gPtUmRE4Z8GFgW25Zlr74A61Xfp
U/iXfIogO6IknFnMQV8Unew2PLdLSZSmnfH23qIdcWVgM6JPT37BCGneb837r5ahRU2COOyzKrbY
RbrW28oAQt+82UBW/pHqeITLy6zMzcrXKcigPlYyWohlHADUfj617uBqTm5C3r/QU3BqxuZrurRW
kwiXfXFSGb2K8Hkxcw+Z6QYcy0HIaGhMKTZNtAKgY5js/2Eqt7d9VgLCOz4JcWHkHrneQ/b0PR21
85ORHtDHSMtetiwzAZuR/G1xb3q2j5tT5vIlLAPBUOKCUbMM6yd1jlWs0fxuOZIPiT5A/46SajAM
UK3sMpzo6Mjsmh/CA3P9L10K/dbRTvWSO9eKuezLFuYOT5xeza18kbT9WD86Y67oy7I3gmnJKWJI
ECxOyHsi36f0BxdQVWJSQ/mD7sOKRnxv5wK1CgQBiG0gtOZaU3bF30l4f//nhGrXXSXyvgvDJACQ
kBwdP0QY1QFpFEXaEk16gXCLdDU0OnlSP43s3U6waUZ0d1DmfyEL9vcnz1Xo7kGQSleGn78qRn8x
j+c8ochCLdlfjQTwSSbjcyhlzbMGFl3oUbESOR08DlY2/OFP/XqEemRK2luKZ8DwSjGIpQD527IA
iDpz9u7+JH648c9rjpHQoiY6hZ5gG4UZBtzi5tLHeDpxgNYEiJCi7KdUlKt1Arq1fctFWbzQUHdj
1erVAzJE63oYgV388KlLPlgTT4knnOiTGc7q/gSWNVmg0ZyPUC7QkEm+ibDNHyMj+iLRdWy2MoTl
pP4VzTmKTwp5KRZtn2Mv9Kwv6We/QmG1LTXAq+nnauaYP6B0u0N5htIFUNS9nLx11sDattpCrtXo
RQ4KI7nHFEf6Hp7d611cZuoguFHSg07MGCUXffBSg8Atndca65BOiTfbMXMFIq5ge2t0UgUUixvT
hhhxLIpOavBeJXME9SnCZMIs4Kvc/gvTscrWNRyh5bHquYOuAiAftwI8+OVZ7dbOnd+/N5lZbstV
Jcwr0QPsw650tG6zujrbAn6ZhFP7Fs3qbXKTZ38KR46bZGBEgtnXDc8wtbN5YgnmuBSh6fhN227D
1hbluRV+1QbymAHrJEL31L89PkV3PdteDfxEuZYbEpHtFGZz3jP3tQ6OoGhiu2gVfI79rSEBdjyN
dqkeXckGmYsDoieig1E8Vc9dkas8/SbRXnCBgHVE9Ylqa9vzTIMfOEM7+g01XnZR4WsHZiqpriUB
mj3w8seaxes4yKcyIFV7MMR7+e+DdiyrtGfU+ltGbBciCHs/i6jeiFTRtRJoFLqQ1vpr4pL05KIM
aPLXZ5fHaaZEJhqDUMBTaTxqDKanVmEXp8nWYce0xZ40YW5LzMPhsifWyk9w2xPxXC+rlc9RM2Om
uXxFjsGstz3eY/k6xf/HlQ3SFRKfLEEiRXqj6dZhwH4Iz4kK1fa9Qg3Wk6OVNak7kzZ/U8MUsETb
PFV4I8LGSFE2sGKaS56LrdZLPOYqiymXcNQW1TUeR43OVlxMdc3w1M70giFmhlf0n6fTtm4NvKws
Z8k8QTHVJQAzf8MOwnTBUVAvchmDLoJgs9zFbtB4whmCGA8i9QTB9iVvB2oujJox29eifFOZpAaN
yTJ3WeRBMHAu3g1NKSbj5AdYm9dvCKhWs7Na1DtPehHZ1K5l8FsaGyFxammfNjpuyDUE6vcr5d6Y
yr5Dq4Z11+/ld0XHnNeRN2e8qM1rHvfVJEyWu0jp6VyghBvE6FrSWwY7jjQDekTPx8QzJmocgfae
l9d435IJQc/ToIkCxgYsD77ZKxxijD933QAt8dgAO8VwPf5R8LwEjf0itjf8/oiN4ZhipRCzGz3E
flGrZrlGqtssn19Y34JsEgzJvg3jZIJ86FULSFM5jgH3zb3xZ3FKxZJzCuylij6rPuD8M3JdAjm1
f/q5ukcMvTX6KLIUjIrxMhRpRXApmMoYoBsMJ5NwOgAisyzsRaFnGG8vhv67aVyQRtO7jMTub1BS
+ZK+xWNsAH4u/XYSMLdDKJrCCVbTpk2Vg3vz0gy90qL2UAH1pmmg4hXF8LpV5u7mFtAKtDaysgtU
djvkfKmgfzjwSCnFlnTgnaD9AUyYcq70xmN7yMplBI2PRaQPPys5IXN9fc3gsTW6owyIgXD+nUDz
k6rI7F5HHlRrz/8LLEsNI20uZTuP3/ZKJW970Flwi8kOMLnPzc9sgWzYzOJ8YBEBBEfthAk+UC7i
+1JXMdItL+BrQ5OA9ADMxFnd5ooWOqiZOS9SnEkPUnJBclTFUWatnZp99g1vQWTsV1PM7q70DTML
wULx5O+1D0eZj0TEQ/Ml+WQx7VOJAslSL5/lpa3DVjetL60xvuttbhNifVadnPHu8xUeftvpEqjP
LL/MSqWjY53HRzSkMjUV9C0jjG/HL2H0QhcZod82R2IrVcmQbTiZQPD9M/Hu34+XSoL+xAUh5m0J
uNnN/xmrdr8Mhaof7KqXzfb1T2pQH7PjWL+4vd60zBq2Cnyj5sETQ4b1tKg+U5YKluCG8BtvQX+L
IHTcqzYjWJ+SIn4l2fX2jBcHk+CV9PcDPPeotnyXYSUifQwwlY+ii9KinxCn6Fvdo463yC7JooW1
xdDW7mUb4dddQU2aA+F1sxoZjE2ABMDdRijSSzRQc+Yvqvmewz3T74D8ml5zNK2HhmcA9hfIXfZb
N3/8yUhGt4PcmT4pQuR9o64bTRkcTlOkYR28m0aXFsmP+fjQSwak5cbKcNWwOqc6bwDa/wiAMc13
w3k/FaFmuOnSW6azVvQ+Pw+k1I0eB84clGQMRzUlydrbtjYXU9JYXLvt5UCoAJuWhJeWOt9xNX+H
5FzvL6vYiPSJ7Xha7sq+vAYoifzvPwsrZTWvVteJcpk5VbxL3w0ik+Bnp+w4OdE3KXVP5dv5FIn6
caIyIB5DWjR7L97tplQtlAyVlHkKdVvZQqNxDp26e+6f9OpKPejtmAbB9hwAd3ycC+VT9Vohj36G
kn/nqcL+W3Uh6F7aMKyCPw8hV2uGvrArlMCwkzKlFBYt+bbxbbnNu6ZjfifRvRTqt+QzTWw7TGKC
2ZYVHONKb9qQHZAjQb545/m7F9qLGlLLusc/K1LuuRBG6lbman/BF6w5mRw03StN4+x+ux2rmhVJ
3KqRseJuJbdVsiFM0ymr5QSjL6srq/3EDENvmypswczjXJtmd44pPOXcITnAbaCwmU23YdtGSuXz
zhypFcYZHq9Xsiw4A7N7O3OJKiFQXshbnKj21AxT8P3ar7Qf7eHJg3j9oxfCQheNJKut5HxKpu5U
w1ChyDGV1HEVXcQ+3phY38/qpnAH3oL6hKfd1UwFFEH2z/eu2Oot3CulNB0mihRAId0dXgFpMwoD
n9s2HcHj0OXSOsdp0rjEICIGKlYgs/s1rAd/+s6BovQ3Z69G3w4jvG4hR4gy3EDR8R2oeKZDZut0
NsELQi1yday+K8DMBDggAJuvhGuch2pObXJDHq4a49/evs00OFZLIzqc6p5rjVoD/mG/FK1h7hLd
OjQ2+Ti/yVhEops+8b0Jsl0/Qu+/ngVJ5aNTGrobwi3WP8Khu0yZLZTxqDp0L+0C0MBFH+F0sRLQ
3ecxnDUa84M0zftjGRtirCVJgc5nWvsH4GSIf1To2JDXNJhoQvoqt27oRrcp7r3zedBMHPnS+1HA
zGokUfVqdvXmR4pWOC9Y/bdX1YsFbfQBDvj5utflZ7yYYyCo1ZCA8YNs3B0b+JQVcvp/tjSL5JBV
ouXCrVwUz4f+fQRwk/XpuqBWedyDovvoI+prOI01xdYsreVtdeFuhD4XIhSGu44zUMo2tu1bnW36
QTBTVYYfItXVz6gBxE4f8PDk/8l44W4pVxymz2IYHMcDKQYz2ec8gXqk2gKaMtbhYiZKNtrYU7xH
+rzFkPUlKj9aYZzavtx8j8ZyzxEHmYX/mrWXHV7sEWER90L1baThMmAfNuPJso0ykTfz0MwqiqPZ
/EIHWXJH5pasLc2Ofv5TtnaX1SOdWh8PRA7JSGko3qeIpqg+VxUR8Wi6aGC1OuUbny2liFO5wVgq
iTwKkvO9JCd88AvkulgQz835LAyifQgzArB2iytPnwVPUzYDo9G/iMLPXfLFpvX7p6u1M2UMk4+g
D1wW6cruLj6D6YvLCsmH8pT3NDN4hoqveZ41gtiKs38V/4jj0/yalxZTaWJidlG0oMdPI/TXg19x
Il4/CWE0w+NjzbASUL6M8WF6AwjwkMrc5kEzqRT9EqGdaH/utwIcNp78KQF2trEQRAeFmnd7ywUX
HsXmapqhxi2GD404zMzw1J/bSnka/2zPBAvlA2fh52qWOPbXjtT3y53Mr21/7IARc1aJPl4Xcjab
CFdpfzQKpSvDFuZeroN2cVYuyOTx7m+V4aD5IiqEMpmKmbBiafkz6djO4lFlH5j8K7hHbSO4nyvI
TikbBzjRjA7tyWCSqMGlqeBZAcYm8aHO6IJ5eKKSSaMjSgfj+wzHWSJom08HM5MTvOvO+EjiTR2g
NotPC8tpQtKyTFChDrYsWXPzwnUwsRuuTbF9mkDBMnt69I5dTdf4GBRY258YBj0lVAYNY8QZAbUz
8BreDMcpLUyg2kuGaGtKcFml/ExJWzoKUDzxYM3zj3MOENIx0nQzarHzSkfiFDxyqOEJOKZVxbvh
iSrd4IjOKxDf8AEwjaj83MHEszUvn///FyuHFbwMrdoYy/LkgfKQNAF9fn31yXwvUlkbBZknt05U
89ZQPmOs7b3pzgBFMzKkHyIqoZbyi5YdgDraSXpQg2pq0EB/W/B5McxQQQdeRuODot26pJ72Xlun
E461wK/dVQKmd3W6BbM/sr3O2BasBQ2Ojmo5KXz4DlMntW07xxeycRnlt5V8hnaMp6+S9CFWP1IS
ramNovIa/rXVoodpBiWWYqkTRY29cX7JtLCIHhNuNqjMo1SfQ6nBqxC4LAMhuJVlE+4sj16GPsXA
V0UbkmbjW7p8QiTLfKfA6sewWHyM0Xlns+bpqcV8XVvUdw+e87PFHokC1qRCL8PpaGVzxKbMSQrf
pRZ1fYnuYLiTAgx5rFCB1qcTgk/6tHqpDVc3IaREH+iDuzPrcefoIMf2fWv5Teh4eLgi3go6I0ko
/atFj6RET/4Imp5N0JORu2jTip/TobdenhcW2f6eLaMLAY1mOhzY4nFVL8XVh3e1k8COVRrOYS3H
S8QQhU+CJ/d1q4nSiyYhoFAKNDSXw1nyBvRAEyynsZtgE7JcY77XhBclB/0oTiidSUxDa+zfKrlo
mQ8A/iGjpPvldogaYgUH7c/C2RkesHiLU6b8BNGPlWanN00PiLpD/nXnHPN0Dj+LdrV77vDK7XEX
pY+DaXfMOR605d4/Qxk0lLrp3n4noPl0rrGqtPFGHDdExABjh8rsYDhDaspkddSSf42o6jBFx4bg
woXFJUbGafFqHKklIax+Tn1CkV+kt0g3yiAvmNvkCylq1I1wsxkJhO9VixY9vgwLDSa3rtuGCoFp
RxvA1N2kAkMFFcoeWeFcrUYcBndKADGHJRHEkM/WHTIKYnynRgnkQ5F5ItsnhTIxZgay5MDIOfBU
cigtmOmEyQaGNRgkTkFBG+3vTZC/WkBxguwMCWJ4dFSXgV9/CUZk5ZhCJ2+7mUrZEc07po1ubXV6
xCJyNc8RoS52nhaAfS45gbiaLTaMX21eHh1fStBJhKu0h2bLAuxuSb+Gx166Ubz9zFcopW7Lg0zO
rNuCWfGp9swoZ+ixrV2X7i48Hljh5kNlMUEQMJPLsUBrWT437e+uI5I3KeTr70B5A5AzvzOM0prZ
Tsee2lcdXH6GA25UytvxwTp+fHQV2R6PHJzKthvQk5KasnR7fb8bKT3tiRrsN9Mh/aH8LI4sDZSt
D6XMYXKnPXdz8+p3o1JnUNlRRpGYbirHa/veumZ2DqYZwr0d06VHe5Mku27bayERovFv/93Iha2O
9tzCLzKXNOQ2JGvnmdYIXZ6QvjYvU2wW1gaHGbCiNgnsNmYdDXUnBTlHwazlU+3LNTGDApYcqvWs
FqqBrR5V7WhB3ciCe1FhOqY+C74W457dQqvrFcsPdS9ZlKlCEvAtCt4f9RaiNKHclkk2o3AGYaQp
2bFEV6xdAOe3tt8WG8x2H53kd1AjxSjsx3e08neGvocwzRG+pbz1pR5bDX7EJuj308s94RrEGg/B
BaMu2GsR9H6bs9CWiw9QrzLPwP6VFjZZQeYQHW5Ol08CrvcL7b9BOeLxE7QmUnah/NJ3v7wm4XIN
bewuCe3LQbPUjhDHaPlNHeKdbykeCkIX7Cd3kNaJ9Vl6MYAVRusEIVqBskJvvEXgJ1+QCfLC9Jwr
0/kOQ4Tqtg8hWJKVMzpMxlgevpKdC/ySvkMQptQcZOnr0St/3nQp6PF/J5iuCX9mAh8/OgEN5sFL
3kUoVhwqK8iK3yte9kpQilCO55BnBgWJt28GsAaYe0yFosQQ5bmrij8v+CVlUc6F5aCnQBF4PE3X
uMSYIhoKUAv/Ur3C3qoWk1Do2pcJBJ1D/yKswOXDa7TicwDu6v8B/v4NdS+9XltxYeTqK6OvoBwc
sZYWp0WTjB1ECSPKDiQk4r6Jymo9qh/OR/MoRnq5hoofJy7+qJv7MNO7XzpIrP+KETckxXrEZXTv
Hg3mv5lvMBfCk0uS0QJjYJARqtxYQc/q+pj8urh1tMelPpI5NN6QEF8HElUZijj/3QwEaYrT4oi7
PG4vkc/Gg658cIwM7LSQfUAlh+xpioQXpb6m/lvsl4G/9RvV5N5KVjFN/rrsV6ki9ToBl9mrus4L
NawEtnFuVpMrxic3OSVNJmAsOJ3DUksW27tQkO2XT5RAh1lvDvl5PbaDIi8kkNdnLoUGnPyAR6Et
j01jbWxEgaAKs8QAtB13ox6pl5EvT4ZNaSguF0Aye51v9W+Ln9GsDrRmXILYx8HIQWgorojauKHG
QjFx0UdVPu8B4j8ixdhs8CITLyopO1ECCJhwoQfBwIUm/7o5i42fQU/HeXHBVRp212hUHAc7voef
HF/4Kaq5ymTKzLj3hpAHHBUJEJxzFMI8qHzw0qczuC1jLDArITH/65sf4+z31v5JmeuiaWkvazZC
Qn3F9rldyfz2RLqDXRTRBSGBVXTGyMlqxWr4LAPnTEuci+mLzjJvHZvgCv39MNBA0wIkWtjHN4yY
Nfum7l1bLoFz4X+7cXOPFxDTaS1RVtiipmB994PKknd33uA2C/I27z2iuZhUMcE7HW4O3b+2DDr/
9f99rtHt5Or+qAsW757vSbnO8UjjeDPZoco+Oxlf6lRicU/R4sVHN+AXsMVnhiStkgElgnym/Z+9
ov+FnacnDrrl/ge635eaOGvWB01BwzTOi0JTwlLRdJYY5hmDS4skVWicTuDSVRONBakfcwWjUPR8
0EjppzaIcUTPa4qFBQpN9Wm6Nv0yocczxDM60r8QFG+TbKShGo2d9Z/RmoNFJdpUq80/KAZ0dKGM
ha8Q1tGra8/pWMODFL7/iX94HGthlw2bJwLLVBtsJr7EqeBvo1jMfz1S5W68brlC4zhIOFR1NR50
saAxWZ5sL9X1DmQ7crYFhYgVeQd6tE78lSgsNxFbhcUr6P2OddpJLXIwaZKC8fAIkgtJBHSxAkrG
SNpVIg03Gdtj7fPTJvg08+QrXhtHUUMuCDJgomQI+DT/02mR0uQwJoLDURPuWpCJy02O5WarDRfZ
9Q7iK2SonK6EqrYsKIcWpKXA9u6BGBdk9l241LpOSatUB2fcyWyVqLY9rI/VqpOi18KDIuIqL2oy
fUPJvhNwYrdG8y7sol9WbJ9VIObxHGllb3+QFpPwg2GV4ZVU0942lfrZcF9BCm9qB7uMcdx9OCKf
jBVtdECVSAEKzMGicZH/blTSlNG4eJ2kjXKZVXwwFRuQ1yx5EnWceMdzwP5K2uqjpR04ENbAxLiD
ptjUqTD6yz7xlykvL99PJPW/DYfb9y2eafgLxE24co9E9KCP+F/VJ7wNc54y13fIgNZ61xcVt7IR
xpjTX9JAILa/aoKe6wu7CQRLfGCcJkyEwGIjShT4tbW7rFTCIj4g9qVXc4SfMfJ9D+/j9JLPuDBq
pDXtXtKN5sLUbBI4MbMxIEshY/WM2mi1dPYz39IL1zpNKR/3ZLjbdGUAKChag1XX48iHCBeWbunw
sSs1xArJM39vjhw2WqP78DIKUU0DMX3zq3VBsdJZ5E85sU6/KAWwzoBGaayEVws8c1OsondjEl7T
1S1vih227BFiASzVXEcDTvBL6xpscHY4IPTKiiDXU8htw5eP0INmZhAULEw4rasaWb0etrhkUzIx
k7KkZFbsDRzs5rSKLSQGMy7hWHi72w10D8z9Phi0SRvvBD3QRZCfXbyVr/tMDd16APYQ+8rt2DqS
ZStT9hJowy8Pwp8Q2yyqLRrg/+yxCHoP6IzRtFG0lMwXjioMbZloxS4Oqo8d45waOo7DFiQR6HxB
+sRJ234mDCffThkTwTuvmOyBl9eBKFRXMZXT1waWWt15RJoVoRBSL0jc31vqr0IsxfXCeUwYAMJe
EUEVDu3qasvEhE04FFKTEWG6Av/Sn5ZjuC1PP5cigWa02auLAkjjFagPErM87QV3mG2zCKBB+wRZ
pf9z8h2OXllgy1ZjCujmbH9XNijKJL21TMFCfJKrTHugMTXDgjIKa4L495Zp6ooe0l9feaujB+ij
Y249R4g5e6CpjX9+XuzISX9v3n+IbphJvzQxXnTnAbyQ4BCepUyX7vw/hc75VOpPOxKgZvDQvoo7
IkNDNHE47l8O20d8GbC+eUChj3LbCPZvbw6Gk1ELs6Y1xWZW1nbAxsHlP8p5UH8l3IOHMfw6jP+M
4s52W29e5uWwbGVh6ze1ruB/TDVyMtLpiE/1SE1/YtA7v34xlN8L74PvAN4xmCG6/IOwmAjwD8xm
+n0azPi5tC7/MjRTV1EkVINweivUFytWyBhpPGVKBPtdNtu4VFTr0xxbXnWGgZVi/XTZJa8Xa97F
No5MMUjWAxYZsmGZxpN3jbUcn/O3YAAbDiX9PMgIZsDP21LZx1Tl59rfxXFEewq3FjNaDtQUziZy
HdcPNf2l9arK5i0JKxowUpXpLttz5wK3RDYmU7qmvmoUPyy6o2Wk7btCfo3SYTU2dwAgbD6pykNH
mybEi9Z3NLzVAxVL/UoA7ecQSlqTLDSMBRPB2Br4yrh7vrMupzpYrKrctIJTLyX8PqIsKIaiux3y
YlNrRa4PSVqXi0yti6GHYAk1q6g7cqT4RKxs94BlgWuKceCbIyrAeiBW4WOPrEpUgNC+zfnGPG1E
m8A15QtdfTYQcWljW/TyNaghFobPZu8rVVYgBMtR/+IUANxg1Ly2aEjswMAgOly5upNTQT7SaLVP
ch2SSJocFJeDP40G+tepI3/Mg86z5aIFJiIx/K6Fd2h3FmwvVaqsTEyl4YWcqkhGOC/BZE5mmWvJ
nc+mDfBg5qXP1+2JwNXwB9/QCysKsgrXoB/Onuok/F/2SO1m6EoLKE3sJmuvtUQTckWVZ8WXbY/O
X2yF577N4L50ajLprjUehkWo5VfHNXHFTEx27r1HQbOxwINZ2BaRahOB6ECYZ3XXKNvOfggrOwy1
hoRetbBd4tjtSZzboJyB5xWFcbCbolYoz5tYk02kOnIXlRRutBl1Q1jRByjiRaIICQu9WUqeOIvi
hCo2cIIHjGbwjb/QzR5dhMc7bOqd0tkm69DctsOaUflvYoa9AlpvSj9+c7IQbgjdesCg3TaE9sCH
kMyRe2sKd+SfVSdWQqEKCQ02XkPdyHx62fBZKdHPl1wkR+HmObHg2YkOb1aBuZtD1Hq1FuYlhLgB
qx6+NeqsiQNwTKaAfHcLqae4E8I+TjDsdFbOae4arZXoN8E2LDhztXVTr4C04ML1V/HeyVnDysn2
9tWkbIb29Jr89zFELP1fkm8KNunfb1RUNNBwJYgQqRtHY/iFWNK46K3Hzb07RRuZr9QtyWiKXumG
MBh4qt+Gg4aedplFxduYI/aDl6pOdbYwsG9b5lefXXBt6fiG9v3qdcMJhY1ItTCE8qeo4avthDzw
CEbXOea/w4briuN1puHoDOPhF5qYLrFJPgKb4LiOAe0RV4jiuCu3dZPyLn3i2dErU5xfw2y2tkLt
g2idZttY7KzK67C9AE+0ZC+LRZ37S8rgDRwckK22ubrsrwaPhh7pNs3m0nwfwiMwISglaUBjL+bs
/UQASIAhI3JuPxXHcprR+0W45IO4NBRDXxMe/Np/XQtKrQt0627WymIIYtTShdQgPuVzg5LR0DSf
wTJWtyevPuylXBeFS4/VLkv5As1f6IOdXtieB1mN69B9qE0n0TYCGwKefaA4GTRue4i3SckubfL6
h+meFCv7w/Szt8ZU+jXS7uyajAYDU8sVClvnNkXAzXNFiJzxjkTxsNIjswCmeaaDDYYkByeTrvKF
jqlX0Bpn+lUNRyTkjXV9kRPjeq6lt2B8Bsw7wQrtjOtVmVNu/W5YwzHZEM5XZPjl8n97mkCRGk8F
nmy2oterXSoiMG1mhP9r3ojc4cnsb4uIzYLFr6DXD7uuFMG0ygf4nJOgOZmpv/dohpMYgnYxQsrT
96QytJ18nJTIBZFc4N0N10mq+Ht6S8kY/Ol7bRLDviJw30FHLcSxfc2EXAwGPsZlzvsngHKJzBgR
iavuTnmxRTIPsFGt38xq1Eywr367zG7btJKeo2qHKyVhJ2TDNHwmLOtf1x7LvXTragPFOmZczYFh
z5czdOQTfDOcWIpqo95jHO4D7wZyF+gAlwYGOeojdrEv98muFnM1vZ4ngwBNlJIFeF1Uzg3PMcqf
NJqdBrtp19D9UA4wQ1QpE4f/25xa+FxEWfOsIrdZxgehyZnt/AVKd7irTXLgqgZ7l3PK6v4B3By1
yd21mRMeH34jD5zqjPHOyvMeIlp52/B7jG/420DNvRsx5X4ggoWciB5Ns8OajnZJJjpspiKRyrtS
0BI5BVzSyMHtPYdX2FhNL8iOq1162GPuCysJzmHdSpuKCP/3qmU0dFKq8Xkfl6VGHWgxZXAEm4q4
x3PcDdMdtOv/Eq2NEs9OLd8yHJEEsQTzOFq5rdT8YD4IFncQdHHYwvxstmCsdB90Ul5flYWxnrf6
jXH+GPeErmbSILXzJDkj2JxoMgCSooq5pkmWYhyHW9iUHEtCyG55sA/pAh8KP5KUMyeqDZUhpxNl
nloqMWXG0egS4B8YX7ju9qR6cqQu2fgvWeWvAacHoZKKQ/ulHTF8RBCH1Sz3qkUO8SvYhv5TS2E2
yAdkMOmzq8Zh20id5XAj3gU208L0QJDUEWCGNGtYID4a1JDPXXjDqw9HBAVts+Fg8Y6ldd6LC6yd
CAS7bqmNpe/rTyUaeujznpIxRI050Ks5G7oYBAgtSsM/vyRvQC5zPEQlV8T38pq5bm3AKYLvdHD6
GYoMu43zjkRltwMkyUOmjJl+NP/MfA5r25/zJnnABPhIJskbQMmPnO+LaKlmTEhDcSZqEOkU/Nrv
WSKYXYdtbAJNbN3xwYhKf2oTAue44n/yASiI4VscJNZfIvW87i2er8AUSSa9QOAb3N9bSR+0EBa+
/EyBl4AyQRz099IBv/UujUYH9aw3hmlUctDG/sDlSbrwTai5qB9+Z+ufRLR0YkmHdtM0KtINt6cU
8OqjQS0vrLGjMNAfidK2Nix/zUomC5oiUxnKbZrhHEE/YoNAohMyxEurbxRfxTd1nZnDl88mDd9o
/wIZaRUXl/FEE/SJKNkKcrT68wBFbdL8F5aSwB77waIKQoe+IxjU0c/vYmdbGkipi7bDwty7y6Fr
AcFwf6wSybQkQvp23LvQu0SEAfy8NUekN6ahu5sbxReiliryiUYIrT6G47G0aVZ8xSx6RV//hP2X
Dm+Nen1cQO8kATQaRM8JZV8MUWhkzd9TC5Zc+i6zNRr/etdAfP+m+dwJIs6+B+3pThO8TwzcsRpd
+B5ZNd/ViDSQUuwOYnka9Rc308gv8ZL+nJwPLn9P1+JC4dj5+BQ8WH3ID7/TW2Yikycwhcd7ymXK
r86D76b3jIUJ89eJe89/regQ4a9nodNX3JlycuKPlhc5rOWYM3o/hzpa0X49DSylc0DThDYphKiL
IcbHi5ctlIuOMxFoQSPr/+7cYyMaH/yQho+BAo5QyhA33qIrcHOqt1lOsoH75sl6q6XWLks4+jPa
mR+scf2b7xlrRaLkNfAQHK9TEeGoc5zKzixXWcJbXTxcWiWC0ddW1tbpPkI64F7WqwEcb0ASj8/H
MHhpDkv+5XVMa4Or57zjYOIvulgRX7e44Ae7XZRCi3JoWWd70lMPZNYNyMNpnPJGNcakFc4iU7Kp
qAEZdsDhsIYlntHiI5v3iFD0kr8pOr+Tj/riVegpivglqPNXTqSOMJDCYals3dnMow11pRYmElkm
7QCPkJh9QGY5sGeSotD9ZpT22GLkg8OsBhi3r/46MuCDMdbxE0wV8wKH2WGiamPKxWG6TL9xV16p
UbBuUekUpuRpAsC5omOnAp4hP66m0tgOq/h7O/C9MEdMp+NIBncj8YZqV8LsvTc7gusJNxhQAN0V
BOQIldEixKY77X7A3nohDt77t+ZMjhwEBKUapKveW5MD0ZvAtQ4h7N3AiPy0YUqqlQTIQRMHiyxj
1aDD9TAkX8M1lWAr3R4QrtJWAlKsGxa2X1fUPkBByhfGZt7QU2dwEhMKOxIkziKBD9bOrIUuP+rN
rjytjM+sriw6Yt/J26IRvAsxLgcCRVvClaPPEf5jo4BbGUrdYlZ9+kJYiefKlmes85JGykSvrVNj
iagaATs0Cn6LL8WiL/dsSQnoqvJ/EOT+6HCaQ66sNA9ED2JYTwNBvXSX3LwXW3binMmRSQiqUOIU
urUb0pPmWl9S1DdeWcBqGG6ozB+3ybqiEEALinr0NlWttbBblHyqo224cStd8lvQUpyslrhiSuPt
48uRzrRj1OKKGcBB346SB+GqvrHNLv43FD7xnl+AHNJmanx7g2TZ+ZBg1tAqvFZqVF1DyKd8sC0k
pL0QMhQL+PFSiNv7K4gh1lK4chwepuuUM8jpAeozyE3NDqUND7P8aUY04Y1suNEPx1s+9tvkEPNr
qYU3Tbl4omu3mzVy8i079qvsBi0Wq8/E6L9bo1Wow4O1X8Cn///l/KU5Cw7cfy52E0eWL5lpXruZ
h1c/uZAXwgdBQXpR8C4+S0F8MPKSMRfsOzWAKjDd0aXSvq+tsyCEuVB8H51gt6dWwKIaMbT6+2Tf
w9ObKjTdEqYWTPcc7Xv15ogdsm6+pSBfMCFlQDnBPRQmzEfMT/LUvKURnehvKOtuKOqo12rVqrYC
/busOxN2ROVGP1hbGmUPuvXPHApirX+WGAaiUV5lmK0JUhST2zlXaXNrga6d99gP9yEHZR2u2IsQ
7blp6FORu0hzAofMQrtF/DRV0DYyh5Q8TBBl55Fp4gt598ucKDTFdq60hOUxqOac7ibq5Z3h3wV9
q1eO28ImBqSXbPki8m3pYmCfJRnBAVvCFhYFkxjLd5BYSyf19BqcW0hv2pOHgn2DqMZ2mBDbwacf
St753vgZ9jLzDIvEfQgeO/tgsw94w5k6c9ezZtcdWVK16vrD6qw43i8c6QlOIjSaejI5JL9t+gUP
iCctpuD5Jqhc8Jq4BD8pk/kYYRZk1hajKePcCx0re+DaOwCdEhgOMZAvQrU8CkO7AFxz8d6mfBUh
+V16f/GRhAGwZYMjUp9P2nUg36knHNbgQ4YjbenK28TlcLI/G0hRkjbsdzh4B9R6LWv/2JoRXBF6
xvyuJqArGxpf/jpJy6arsyZoEFwWvwtoaFnL8r58bNxPHi0Gzz8amhGwyXqqTMl978WrJaixAOkQ
Q4q5b1BvpTZ1pkyvFgLyWNThvLzt1/OlmGBcPnuFCp5aoIjxl/Oe5NYPt3kSoXMa+QTfE5g+g8wO
pGSGKkz106znD7UL0Uk2y0Tp9jg5zYTTzX03ZojTc2httF63Xc3qCva2IpRIyVOP0/+ShbpA/g9q
2EA6nPk6qhJYnqxUI6jku85bais8XZyVHYvGQ1h74xtmHtALy9bztQ8xRpwJnRb7Bx+lwatrfZJc
SZd4pzjIUq90iiGf76C211IZ0/QVeQHWSGWvYFF2slTfR/sZKYGm91HUQAIl1iEyHlIJdJM7qk4F
uaejDPBi5F/kPv5xxeQ0BfNxamRi3AAw0NQfU8N0IMfzhQ1LsUDOF6gFnH25GHUOqL8sox83d3Tx
fHzyr3AcPLeoBKadUOmNf0THT9hj56tAnhL71By8xyMhtG6srEWLIyrPbz7HSshfJ4oNEOEJ0Dix
ZwWJrDylssgLt6JZw9F25Hc2SAZbKvhuc0ShKc4vtgx5GiAkh3iXZjTUA0Y18klCYSMUnj90jRzD
t0B9Gk4OQPDpOsjVNGQYOgLsRgUhAX3UbfMw/Vgk6NAFvh7oLhIdXd4SApKg+txd6ucgwSduPV5v
nIiSWnBrg4JLDaU0MLuqsYYp+KZCPOlTBPy+Jl56aiIBZhIMmn7eSJNZZzkFfnmlLvi1UM284TJf
R8hQ6GuAlUKL77Cz8cTeia3V2GQ+7EXTbBMrpx/88SuHHwHyRE09fkmMiXXd55JQgjQx5lehT1VX
sStlY73pJwlwsQr0z+aLSVzuwGgjzOMw1yc9fVLDs2zeQscscDV8XB5PVzgAuvvuJgd8jPJBOFHL
kX16MKT5q3zvCZ925Zut5Xwk7O5ByZMMaJ5oNTJX3hbglFS+FF5dApN2d+0yoX8YwFdJ5Ak+muWe
sXoP8kPE+qPlXBv6UBWI683KAl8f1QgS1ksfESV8jp1n6SBuIhckERHEj0mFc73ZvTN2LIC5iIDi
ROa89P0yAC1GSE8rWg2MPcV7DoRb1aHnfG0ha1PZlqwLb+NebN08uBBDDbWnXnUnxrQEpz+ggGaU
gBZ7Xr9AxtIxOAorFRjiGIW/X2x9AqDnB7OyRKvBPhOkT8X+YbYytf3zyqjShveYAOLjLP67/qOs
4wwSSiGs4woDPuIb3P2n71u8h2XK5B5Ok8ht0q+OcTraXOD38a9LscyrdwGyE2KHucNZsLl/ddCh
AUZm8FSM3Es+aDuFHI3d16grqLm6s3kwaB95uHtMs+WPg2q6821whSnFD5RNe9XFbEwvnfc3s1hu
2boPj8GO0kPaPhnG6yB7TCsBrTCMLsKEywkE5H2cdAC500wZcEbIpzVY7asmMTunL59eINEmpi/g
+idSZHAeULlOxL9A1+AdSafxOmPm5GJfakSQhFTpvfiUavMWZg6XzHyhTxhIy6CaFZf7K1V5UyHy
MOgrEQlJpkRuvetcgPjwj9CpeWediqFJMv5Es5wfqxY8yj7ZApxU5BW0Y7UbnyrgulWQczMvENSv
PZk8aBY+Q6tl5SVK67h9Q4kmI+OuDhH9hwFwIYbq0NzJngtGGEjenomaczDiT7emwt9zv8z5MqsX
gbMnJIlznM4uOA5oUN509g/1EK9TGIPivoJB0b+fDrc/ek7WvJ8SVjGgyu5oQPP9hXUWzHA4PJbd
0q5FFFh9N9a8jLjpDz+sBw5uZZf2Cv4gD8IUu58ZASQO+UhaQQwUcW0yFpB5w+MtCDYWz68aP97T
E2oW6TXKPSw+IYpbjkvnN4IRd2jXugMo0GWj3zl+9b6FCd+CTSLsZhF8r9jLvW4+8WOMrwRjUoCV
fERJYeNQAPgPI3CUzy5aVhLK+pPr6fex4mlXWX8rf/Gt2VqsyIg4ExSm5tja3UaLnCCpFQsyR+7e
fxzin9LnJy5oVYaqddNd7mE3PmXtYIcqE4mKJmraHk+LXs2wYnRD3LuaJg22ioYKTbmocquhXc+m
S8opYgpRVDI4AqDM6/492WUsWmQqaVTIWhPonl2TdwPZyA0/DDWidLxbNuOxsSRgp000UYu9h3X6
wX+HoCHtU2Xy+r/JibqSlTu1n5V/DN1xsocJFlj9kA+63hVf1JqEuA3u3X7XLJzPz/75ltScsSos
orJvwP14qWyJfWXoRRy5y+Qv6HRRYReZhrW/R9KysWDfX5xHSaPIY6an1Rj6xu0HhOCKK0auCvnR
h5ZictlbxBhRxI4QWwv/ZN2dA/kWnPWtDjbTsuA8QBMQ1mAQ6bbAFFR5yyJrtooU2MxPPE8PwEeI
U+r4FPhGUR93dmnm90rRLTMoQD8dOgA7fyvqMNyu2cp7On6DX0rpw4eGqR/f+hlt7oxZYU5JRVYr
zyzjT8FG9TOa/q5Ft2GbEcJlMsm7VJoWR4ARrnKUjXdoTMXjdiJV2lLn4ecxi5eBpRJcjMArFOf4
8i8BuXTIb1fohRZ2+tmjsQS6giXus6nAJTuL5rB2vccYBn/WoL75AzgIjwH4YMivD4FNLzdnm9Ow
ZeVV5NsoL7H2WoW9sVaFFdb29PLWpvB+aBWEDtH1P78J5LPi0cP+mzoJnec8zySN96FWTanMmhwZ
AtFzwDb38VEmbzs5gaAk9BpRhPHDGhUHvOaREPo1DHMic4ZSEXZpftRZX/FOl6Wzlfr1ItVJy7A1
eIqXuf2O2Ah0Tm3+QM9BMJgdwaHRQdxLWwlYaduXDosBdR6IPNcf0mQzoRZKIf3UyYZqEY5WCzt/
e4gl/oKzsiy+IHko3WjTOZ0w+rnft3LuqwlQBisqiGdx9cjTvzUpQG0HgDIPzhFK2cCohdjcbJMB
17CIJksnW5nP3iu/5fuW9Em310vJ3sEHifHRRLjcQLwM9aY1u+MyuYgMgia0RodkZmFe+DkLm5JM
h63XnYQvpYOe/rOmhw3o4XMJVX3Lea3Wwf1Vje8r4L6E7H4MlrmYn6+BfD+wu/pSleUF85m4c28S
ruCfwazt2VcOfxZTMzb70OZCUqdNSFFAFkBJiWMPaMPxQVVQLtm5gFPRt0FoOnaRXqz0jzrS4jMG
bTzzkI43/xCeA29vUVLdmKEIdlQQ/b0Y7jDNf9wvIAWZxo1TcYbLpZy59Wcg6UACp1hd3VME0K4Q
IJRCLNHYq1TvTYYywSNc0qgc8ZunoIx5nitlZm0/V5GO1oipsA7pMdIlNAbmKjmHrPK6lnTK2bPB
mKSfa/TUZ12xN9YaodW1K9j6v7DIxE099ucHE3qLKgTGq/0pUThGaX4oBqx51hu808zEf4KzOPOU
bkzaYznRcLngBiv5Ec/oOnfeg/Mj70VhxiDqWdc7oVbuFIjwCuT86ueIPIoJuMFL7mEAc/IAqgS9
kcC137AC0bqT2BQGMzzFRVMGvqmc+YqFrXJVqq6fxchBt3/qWq5tArfMsRsqOoMkhpBikyfwWjL4
0gabjeKBe5UQIEBOM+2GtiN//c6XjzLk1lAvKYrHnkIygKbBJmY+hiVkjeyaE82v//xiG27uiL6N
fi3gM+/rGUWyiP6rPvE5LczO2cv/oMismqGELTMYT9qT3ZgdkJYoumFOTBX5r92slI2Y9eQ1xkC4
HCv8AilqjI9tk8oYlvpErbEKEYpYrTw1uZDSrX3fjlCBa+b1SxlzxVjyXGBnV+h9AJ3rSdKSseQb
sEsd0N0oRIS63BhCQVEmmtxn6Kq6yS4xLWsPO6XsDjTxySi0iWfIZQLfLPxbdFSl0lnwc9aIp7m0
4iglcwVenfTuTRzKKakF83DrAA4x7LSlXoW+yEuCe6MDpyCtkCMZgrfHUrPBH4NBgWhjAGUSG1S6
n3zTqV3lxzI/0ZCqT34FUontiu7FZbUlLE+8xjDBQbB04NNOiQOkf3MycAwaTgsgPfIegnlbUaAV
8NAgMIippQNTkQWwXqjB3nODOhKy4HnP27V25xZUscKEcZIiLHPiiSUBgHsM5Bt64DH5T4Zw7LGK
pnIupF+Wq7KgVqcDBnwl68UtIROcUgwd/Uq23zsofH5JDDDqHYysndIjNvYWCo6nwZbNyAz6TlH8
vPBq5Vm9tcUiH7vOI3wpE4exh0CtglrUhL6eVEWIYqdFfAAx/itlAy2TCfYE/i8U4jIvK37A2dek
DIqvIp02n7qdEq9Dfcz0YNqIOXDS9KJNVlnUxHyDwUMz6Gw+GO08Z97jjVBvvmqkJjjkgmVxJDGe
34+1K/bg+nJTldG3uzLDRJwydzn+4D/YqN2jy3Et+i8E9S9wIB1arMq2MVaGCZkuAHdZJLdguX0R
MeGrG/2TZRns91B+/FccBnXP6rXD0LAYYkXbZMlFboBNJxqLd9ihS0iCJa/tZO3parWAFVdAOSgj
MvvPErHZ7aFEL2Z5Bn47eSh4AfxBEEViwcrQ6lGjT0OyE/yzQ7D39CuP+kCJphIcl2U/yp76BBtx
eHTuOK1odcIcaSXlBaYxssa0MB2J3Y/Y3a8nLD++L4GIqj0f/qZRQrqbtngqD8KKLpTk3m5VwDuJ
GTH0fA1hhsPkItYhZqqknXjLEIYLoLujh4obChg6Y7OHxBsWUdOlInkOBTu4yzGo6l+/N9yiRX7J
VdB6oxhuU44tC+p3brtvdEx44Y8XkAjhsfXLgT6jfcvecV+mmljG+H8x08S08reHZH/aJX5E2atN
3b9L55BuR+8pRjky867cl+AP+el+3z1WTyDr8xmmSKLEJ9flQY4O9RVMfl7ZBlvumbB750gvv6uK
hTEBxTH35kbdeHdeUhveBdKBJcDuz6Uy7tWhbTn6WeZC9krqmOX3a84tqHDWuxG9rNy+a+WZmmEb
u5SLbeSTl6cJ3nPZWlJu7XIbJ66t5mXXIcq8c87m4kQPr88b4hPoOYmKAmgM+PhHlVFhgTYBFQFN
otubmBgJCVic9uWcelcHS3BEEKeWc7MYRefINr9chyCJTsE5ktEFg8RPe1Zn/J2TC4Cv8hnN8BEd
+AjI/9bYbM05zhW081Jv6CJB0IvYsSfLZ6CxuHE3p7RQi4ovg5cYVYOMQFuk5hJdJozMElTirwAo
4G8uCfNF+RRZFkXY2vriseIyyTQUq8w178ouB/IXasep1hiTNOknQ8IHdzSZa8GBHQR/MuKj81JE
TN6a9IoZ8uk1mFk9onoJufd+qparrEQSiwxflNAclC6yAfh+UfxkBO4PIsx3NqwLWi/fwg9vkIQ4
qINlLOJ3NX9GkDINkGZRMAim36uIVNAM0wrrDt/sIKdJp06i/ro6aslCJsWnXHyK+Q94eaCgDH6v
StG3RlZ3OyzosJs6CaLgJlADJCV6T6i2YCDocGTaN1XiwUJRKeXr8K2Z+D++vpaSD7WEtXSOx/K4
47Ptt5QIXjOUoj4CQBIt/n7GCzIN5KzesTTuXmcSafe9eT2d9ZN3sbbzsyjA0uOsGPLOPzJO3pk7
Uzufjp61jb2zbMa9uSkr/oUuqVL13Dg3hrW7Qnpsac7bsTNhMjbII9kJNPt7D4bl1N7hyFA6b/mo
Ki/4PqwoTINbmPNL127smTbZ0QhOm+eSF0VaOVRej4CvsD7AaM5sL8GyyHWa94oQV4FxbObhQclT
vp7x3lAhdhlxfYCNLVux99JHTdNO+7+IPnHcEwy6q8SAaUiTAunlPaIlbH5f8IUacqZ8hxRH/Fpv
lxXxC8iBdGLbyHNc0na4EbfqPyYv2i+PPB6NVBFFVoATFmYqn3bgNE43MkXna4Lojc+V205Lx/Tp
eaM1jgbG1odSCSBRCgROvveXfjBKylb9aLvFeDevYQgGN8+klx9VZ8XpjV6+UccbZ/zS5i7ICfHi
RtsQVtwY/R0D5fUd2n52xPAqOICstVSGTjcCc+ahdQ1eXXgiG/Kx952hQ+MS8ZtUfL2xiXkFMTlq
JOMHT3NmeguzEgyFelffOrv/doavcXhdH1nBOSicBXbMAfK4t7SkluQneh/eddlCiTRBCmp1Rkbt
5IBL8ulkwQSTt+OqS8k1+wxkyndbzdz8WMBhIR3510Jsf8s527cP0Im4ovMLahEOciruk7EOK+Rn
omdimfogcSAE9AYBIQQo7g9GweuQqM9rhC3Xv7rlNG5hPFY/tZmqE9l+YEOyUBuW0Kw6EaQQrJVD
jFhJxMdl/N5AmXBuz+a2DUYz0aehZfPoGgt1wDQQRp8GFtdE/ZdmC16BWRBdgSp5hN5FVdcy3RDj
c5zh7LCwwGl0cQoZOBmClUUSuESAaD95CjThA80o98R8CoOUdlm9FfAxTcLTnhGjzah1m/Kv7+9j
SfyT9GAZr1GwJ6oIbkMwGzq4shPsekI73N8mTHq2gVmuKGVh0xYFzzWcijYxRgtR2m3r1SonqYDu
bCLCSdyKA8ox46d1EUI3/prlcjdlq2jkFdVnsqWn96fHAiAEY4C39KRneyRLTJ+/59ON5MIk6WPj
LCCQ+dnfbKreXRCuXbP1ZrazafIMhUtfgZ0+M/zlQq2iT0pMmzzlHdLydLj6eUpCrue1a4qI/y9n
TDBSvC0wlNrZf5vKfBwktWAX6nhUYr8+YvIi8nDdQ04DFV7dxmCyFVFowaNLq1pUuk4TOCESDVnc
RFHaYi/nKIJGkWfckpPE1WPCfaY5b3rhlUlJ9VRSUoLOUQCTn8YIdUz8keot/DgQ3/kpOuh8isUC
5fajWQxaezKjSnH9IURWSGL6A2Z+0M7/kBZV3IxFDp3U4osJlUg5pJBEhQ1mVW1l2Ckp2K3Pwf9e
p50RtviFRETIvmO0l0bdNaAB0j/h1JqnnNxrsonCsdntcJIFMm58jH7QGk3PgRSjDVo6c/zWz670
vb7Ayzg26P1bbmRmvK92gx/WO04o33ggxXejIjKD0L9q/bPyYzdjxLniMYcbhbNszOdt6SMDSpZQ
US67/HQ0iK83VDqFS41PBgTT3+3ROr2LoSIOeCujMB3dEj6ZxCXyqQc0Mnd2s3eEwiprdxaaqHeL
SuFt1Y4Hg1C0GQLbHCXiKWIL/dKF3X1K/fyWJyq6h5itaEJPIM5I+Ifs0DqVM+b3hx7QFCV427wB
zCiMrpCCkjk+ATeTb0YUWh8UyBQyOrY6zJjVUX54grZjmCQslVW/H4oH+O7aLrmnneuLa3YJ8YaL
0NYohqPWttXGd6h0yJdjx+aWsXy8FE6itRzSf2YKkCxhVfhNcq1w+fdbu9TsqH0fHMioIfyAgAuH
hyABhyjIdOBNXJRXv76qtzdAQbDE7q5bsxjS4if5Gtdbq243rXlF4yq5PAOiIvA1WtS0DWiqxZFq
1DMOsaCYGRyqdOcfqo7xIXTjy5Y3pDTj3rmvzU40KwF1pPc6FPufWjFMe5QFXvvKMLdUHE4SAZlJ
CEHMxMqDUKwy5kpDz5Ra0v5N7hGTEPWLeWFHH6SnfohrJM4SC0BvUmkrwzcszPGj3jh3rCNeXDDE
X+DiOg/jDDV1fmu8PUzMMiKFu0FvenuKAdDxXqwGQ2zJtFzfo1USnj/O4yhQZ9uOcODh9JvbllKh
2IcrDZyRctrQ0bBijTQw+n5IOy4y3skKkxBDhvZm3xYn/3WwX2zPoGzw8vl0aNLFhRqdeoAdOoI1
dSmOoIOiSfpj7BJ0BWVIhOhCRnGPrVKgBw8XSrDYrGz54Mf440UUB//7zhl28SrQ88/OEh1iR+w7
xZu8wIBprjnrtK4lQuEx7txr8JQ2U+QCG06kDjDkpNIpN1JNh8wun8whRsAsFenCO1Q4aRLGe/WY
AoWziqbcULgUh5cDilQSPvE43XDlw09IPN9SLb9lBBUOFQvZnJuIMSXhPecqP+z14P/jhid/jbyx
HiR476B7n4oOLIjWRPCwulbfEuiDqXC1Z7vQUpnSpG89Fhnp0glau5Npxqb2ZH981qPrTFF0N8wX
W9xPjLpKvliNTbM4dcOkhHMW+t6Fn6FyUXCRQB+JO51+WyHDQDZlhEY0RaQReZEkC3Pz/Fz/9S7Z
QiFGL3Us9N/Z+mHwQ0bLPPbDaoLeEEck8k0zmfapkB2JqUDaZEUToyCcBopx1vudJ719n14W/l24
i7Bc2WGS7F+0LKipGhZQMJFkaOCNtW8qofS2q7YC/HFhs2KBeI9d62RwurodemRdQKSYvsFNS7FO
ciWGIpTJnxNGfpqdoGSz258A/y+dEmylZ1m5dsHWoN8nG61fFl9PA7WGFasKBTvAjQPCmg56Xals
JUEAfoRnAbw/s+jn6hmqSJkby2e3dGI9+VPw7vw2kIa+NO0SLepV10j2yvncfD7JWDgrqjfDZOeJ
vLlmj2+0m8/9EkhyJJmqwTr+IAD/7Yns5cQvmZO9dLhJxikpevyB6jkh4EmFtz09wBr4Nj2JUtYI
iBRadojGAroS1/0z8c/NzIQh//DNZQQa9Gi8CLp1BWsUhbcqXXRqr21fDh/nCkRcGrsdakvYhjTq
Ph95yBDq+cGHM8Kfrg54vIvSArJ2cFy0k4USuUR9Z8jD3qe6hsXTxv5lgR4sDvD4ADwiECYd/Ok7
q5KAsnXZRkfnPA/DVUXFfaS8LVBH4qfPBU/vAs2MZvhuoJJswo2L7iuAy5xKsjOqzgpYPNgeTm65
jgJm0U25csjn7UH0qGLKLdycGUyoqxCrLYo/nC6I0ZQzzJdtzW3xoMJImB51EUMURLC61cIinm+Y
aNTuA6h58/h2PoAQeMdanEpX12q3GL/Tda1tZCgKVg7smbS2TsKeYnoyO3p2Kqt2K+UeRbBT0SGK
/2oeJJnnabpe+DXu5r2Al4nkIAqcklt4zrr/7N4ED1Mkh399xo1R7+t2Dcu44mfFLPr0pGLOMstM
aRYQ1hQA2o7d0PPm6jF3JYPKPQ/BBI8lLTx+bJYMIPbulIymusN1jAfXeI6qjx3IuYmoxghDuQDz
Im9gTGz3z2w0ThyyCTJgjFvhXrjfiuTfhnAPjoTS4BFjUZiukO1ccmQhdwYcZWZDuqtPuJmv4y9h
3j689Ui+AYBdEQab/cF9SADB75gFuTT4QFPRLnVd4jZnzyA4j5glJR9j2kfpw0wHSkiKQYykid9m
zo5fxoB2B2/BHh2bUob4Ysy8XGoVcUuQCF8vP+epsKWy2JykbBidVvM+U8OhlxW9dU2u/BNhI5h1
DwmozdeJYp7CCFVrtGB6ZtNYuXhvKzkVH8OtU/XbkN+FbNCQccBZb7rYsuvpwzRslSFnqq5bD/nU
2FPct+XNFwWo1UPu1FpLlN0xVHZyEblhzYqdsaEeGPqIF1VPpklFH4EMImFwgdvDbPTXhEM44xe1
8NRQPgur2c8jaRhP/zoBD7tdDys+rSG+g4IzvgKAdbdTHLp0b48itvjS3mvhrXw5tXNoFjmGfmkp
IPV6PmTosmQ/ik5Yfsbv4EvesgNKHFkt2S6qFR7WFGK8RCmLnMsij+149LgGZF+RH6Qf/RjDfPtw
hGlX3HiYBvbFEkfEEMsu+q6DiFd9MIs9BzgDoXndAjZgxBCNuICH0qXBz35enZSZH+23hKReqntD
AMjoDtfdaP+YU344IU5QJPSbhNhkXqsUn9WCYaCwP4j2Njx1u5GiAYv7i7F9QX/dk1O8m4IdOQXS
lSANCXvybMiY0dS6a48moyCkd9qxDiAT2IICcAIfGjhzdy4eSwfCmmC20eGEle6KolNWaBdAdFbM
Li4yn9fxzAjs/NveJ2YAW58+1+Tu2UMnEQF4OTrUiCXuJ2/DT3vuKSw0q4s/89fdROXjmnsMnXbM
9P2GHVnotOsi0Qiu2LmMYEDRXy0JHUukaMQfjRkJe2g8lfkta8rbcJ3In6JmnSANM1XRsfbdS6vk
zLwxljSQGpXsR+/3QFoYb45Lrv3d5lx0Bnya3saYoSky8e9/6Zes3O3Lsyw0fk473I4YjVqpZBuz
YdC125bs88hl/x6MrYjsQytY8in1VV7Pqt+kVlmUoDIzzZk0gr7Izw2Ssq9FnpWocnhWLy3HXSEz
UuQIeu5OcvQZx7Xm+MpjOTNVnJJxZ/3pF6/GkmUFDEl7KvINPQgt8jNLZfEdRumQxKivzxpfmore
8UhThd/yAR8LZ7+BhCrWR0bBroFUqQNHce8fu5quafTJsSE4RUQloDucVtVyPDe7dYeDjjq+Wqza
EFneEvUBmRGUkrUgXb2h+H3vgUPsCxDv9ExbyUiDaRgry10VwUOvLAofTH476zV8CmrXVQndLA7q
/DbHXSJO6jod2SEHxiy2wZROuigvpTtUwfLzUHcjgYSTEaX/hqIEmzZ0JZUYB4VTV8CMXgReLXYs
nHuuRZ4LPGPYHQRffCGFkZGYREMhRt5cot9MDtjFT2Y/rHLV+YaJLAxsXujmlXsIzyJB20v8tlQb
wVkkLaIIDB7VwPjeBsH8QQJ47CaFGLiGwh49N56uyoO6PEsMGCYM99KiuiIVAv0sZRBXlL5EoG4l
/sJppyYM8Bd9fnt+o1GIYRzBHzal/PAYTlxYX0JqlqdNZ8UrrwvEhkdrIFL9KsOibC0X70MmTFdE
ADkp6t1r4CULfMY/9GwT8QBtHddDJ7T3HA4QN4gbtUO/zNjvaemoIVuyPy8717YUzrvkSX3yztC8
wXzk1BNG6tLrtU4QF1NhjZA8Fk/bJyARsMPCRFHRrMTwAJGVrGfDHxfSaG4KmiVYOqdoJU9TBCks
eKB3PkPWdxOLKtb0G3zJnTsvw7tlECD19RDy9bv+lazZRnj3sN0skr4tFBMvtD1ju+QkAYLuoqBS
py1eCS1AqmZVL6IUoLTxAZXyXMdqSWN4xJYVkeMsELSB0bn/XU+7cO/88qgkfl9iUhjw5zOnjcSd
yNe+OiHLoC5RHg0UBiPaaz6dpZHQOq79q6Dyj9q5hh051Hs8qTP5ea1OxHnYI6aqAZuQvjvDGzta
KaGKCLMZe+HelFa3MaGns1/ldH/7WpYSss5opXrIFX8BEEIwlIDrLgpAoh1ZPuixnZTUBJIdNVTq
hwKvToIU4RfCfbhs1z2PySZfoDtLaWSdemyMtjf9U/L7XQq/fPNi5fCWKEppYTmLsTYTiWdaqVUu
oJcTTTkzVnYDN/5h4Vt2KoZV5C7wK5rrlOqdJ341GFPC/VBKE08n/CTV1H513cndNZQh6s2WkHkS
xqbSEaEiIVGdj7r75/LS6nWyPVRql96Yl+VwTUSALOTA7/UAZqg3wFQ13XzlmUESbDkRJrkFF0oA
0ipPqiPcSmzxAa9NWztKMtmmIn4BDlEZSmNf9PuSWIxc27YnPihAcGFLSL0TTtm+ni4qL+7kRjkj
13EbJyqAmrnNNYfBJIk4WGpTaec190x+TmdHGjSyorTQNhxvQ/9T9aQWkRqQmJxJpNQxNJXFOB8j
2VCwpVbqP/ryyhlIyIFNbPCsAdejXkRNRuEi6/fJrwUIbUTApKuqiCSHq7Wc0poplzLr9VVbPHde
8TCVMu40otY+TRyxxT0aIF+4QKVpvvVVQkLJEXToEmQW67iYAgbYdvpcn3yXC6bv1L6XBy3fWaok
gBYD/BdBdzOQxz9+wf400MW306O/UkeRodw+5xrneY1WMalLqD2vwey6DcyawH7loKqd7w9P6irh
Mb2IH+IZJT9bcPWnJpuF/0dZKbrD0VQwXXdOJq3AnZ7gGuyXwquqzZBOf+kcdd/Jeov1fO2LKrFJ
7JPxHepLS5vjusl+6yXnyZkBHuLhSLgbN3U6qzco85Lu+JJx0eWBKfSUg4dGn+pZ4WbY1L2ZUyNK
wfW5DhPnVScarw3h3Xjv004xQzdoIuMQ+MrTPF/U/TuM32C4eyvSnLR2ZmmY0vvpTkx3PX4wqCPi
P08/Y0zWlm9KxEoffVWkdOwTkD6US25aOzeo6POZdAuDnWckbDoSYRo6/RJr9QBhQ5H00iEoiERc
jeIj3F4UmVibEvTex5sW1OddY6ApDun2sOARalWyDNQhWtV3rJc9Lazgp9ZGLTLdyo/JJ2Q31LXS
9GB72THkjBFqK6oF7skUglKvTroUI+1paS9xJdT5qGQUvex7PBKeK5F8COS2WbNOYpT3IQGt1StN
16Az8a4L/0CwZix2yGRyn40YQeTLg0yUpDQhnzaPxK+xTrg5kXIht0LYnuu2t0g+34FsIMcemLYf
a1gYwbQswRHsH3Z8mJAk6wr6W9bwEFGKEbveeGNWyAJmbQ8cBBaN0qVlPTwfCB6zDSUsWUqAUJ5K
eADdk6iWdR68AIF67kThkdlFfu1JGGP+58n8GzPxcGGNCJtJSHLCu76nzEyUoiltJVCZ/GzXodBk
9fhCBxMAaPgiwyKzLyQIQ3M8kbEGiVffzIf/8OaWy/0xqI7TubuID9K8md3g7a2Ibe/gYgekBgUZ
K+sqhjnli/U23jg6iosdX6gMr+1IQy5l1d9cn5wJ25uQlsgnmyCnfJD3FWFwg9To1jRD/WTvgwwm
gfervAKj76gKekjod+uKHl4WrrtGV5fnIKnc3lDtL5Bmvj5Mg4u0ZDUewnLwmFbqcqUuVV8pCMva
nNc2Ff+e5i1acXrzo4Krt1x0bZOxMkKvbiRBQdpfmgNR81x60siuHwDjn54y8WuveSsAmXwIQYUD
F037jAk+IipcIvhEmnBqP6fOWBQwu/WiGm0i27vUSa2Yv6NotzjoPAzBYmxARFRh/LHF19G3UfgB
2gC6onzrzDkBhVTAqbf5pi4y15YW7QWg/mY2dz7PNp6Ru/QM//TtUMXTte90VQ/k+rx8bDPX7R2z
fFyFDFJFLzKkEEj/ehSMP9szEmC/0/qosDLeiaJP6RPKOvF1fiBQZuvuoihu+YIqpFL5wG2AdGja
YxdTb/NV9E9Q4aWkrvpDWa5BtAJDyW/k/GcLDy/wRkUcxvoHpw8YEJO2i/vM4IYZoYHMeJCnG6vu
7JU09kmoTlgRFiam5gtb8sCWao5Bbc/X3Lmj16JYfdzbUNGKkHYww9QtWYO15NeujQ9LSPkmbaYD
7llpB2xBxF70hBKu+pgOHWCteIG95pSE7S2arewq5bdVE/eLMjn2i+YMvDazuSoX36gXSfjg5NAk
mN++ghRmSZVsClwekULR77uS+Ql5G1/ZOZT5x3Gx0enXn7c4l3Ae/08DhXf5Cnzvwz/oBwZm/lS7
4mIOqoX6Fz5TS9BLY40h/nIKP9lewWgP/xrLxRi33QV2I8xoPo8xTpZqGPluH5yhpeEtn/wqzMz/
BISiKF8c/IIULXHNtYQvQilJPEfY6hzBu09AJHj0COTt5QpIHcjVIyYRvwMPDqiD7W4zpNNtx1W5
clL9PS52558sbJYEqjPthNZMimE0NIZZbnhkgPPmgLookeAQeDVDBeG8JnLim8vpo7khGv/t24lx
aCnjtsivwGyA/wlqwcJ45I+WlfHXwRzks9a4lVYNLpU0WkV+v/nE4f0QDb0HpqgswC1NO91dSCRD
qyXpVj7nWKslg/aA/PpqR1HRjzyb4uq5kQi2xSow+knD4S6DH/nDyxC9gytOGq7K0wFmmts7YHM5
TMmDR0ecxcXhOSST0mzIjjusOZYGziLQMfTWuaH5iYv9AS0rAZBFjCix/YybIw7/7o5vsZyqC1JS
VBc86FUo4egTutPhhltZJkIcE2QW+Q1UR+tFIghrUZRaTwrL5A8AmUGe0ciM4yBsGfsa8O+o8MZi
Gzid53MYF8v1eMEpWGHiZy4Co7j479JOlKsB5EncVdVTBgsTy9J3No7xbd/MeM35OizGgDGfuE6L
KK4p3m67Xn70qCtfcOX+UsmxlnPdxt4MHybosJc4uk5C/HcliUBq++DQGnrV7YR6me2XYfsixWpM
b7pXYIpppQL8xbOCj0oi54NvLp8aP6aqv8hUyb9V7/RwsSL0h16tqaHDeHBZa1Fx6fVjPADdeB9e
LND+HIjSn3A+SEClkDsU2OU8LWIA68AlZem/Tlzv4mQJO/80nT7SoZuBOvNxumhWIo6WseX2lJ73
n9hdUKM4DPuM7omog1XEmoPFkFZLR9BHa94ak/8/Oe1IqT5Eg74gyzeWpGQhC5OG7mOVbq55+SSg
R/rwowAWEYIyUyAwd+4Cl2LFhPj8IPH52SIjQVqX9BEUVqsISnSF1QpcHHbK/t2QzxGyxM/X5cO5
DirFe+1OXlj9he0TtnZAxbF4XI4fviLlChAaq9KFbGzdYIV53Plo7nFPTIi2vFGwq3dYKEJjjCJP
X3zWoJGLs+IdzfYVgPEHhR9NAfllLuKuA2vkcgB+JidrkcBpJLvNRp/8NT3EsSUovBlF+m/1C9KV
Q3Nj1i593RaJFLBezese7dDtXw0fjFnESoZJl6dU1q54MWJzDPKhREkLmNPwY5fidOnHf/fMDrO3
E8IxgFE46TPFV/hSvHhxJZ1IRHugLU89D3Gwe/cqJZLyeikpjym+R1ibBMjwa/u+sqeEjIelowWB
KJvVMQCvqvEmUHGJvU4FpqoI2zkESDNYAwjYpVC5I50hPCrVn2G7vgzXT4Qdj5paC6lCOEb7i0SC
PlIDXUSQrcvZDlxx2kCSBJKHVRcPuQmygoqmY1sPxX+6Tzt2+wEPgT2sW8r5nsSgO6b7i07VQwr6
iXyDLupERTJsTYUxO3edAqJIGf1qJW1NDWqbc1sDenrlND6980b2n/pEFHfPvtmz0wTyHYXnYKtS
DX9Knr3nDK085p9w7IytNNe3frh4bfh5kQeEXamr57GxV6N0RASAbu0X3qTZKClSumKITVDsJtq2
AlnZNGDN7zwqt2mSOt1fTiAO1fD3iP0Kpo69TW6DoW8cKbdRLhJTeMIbOCshqhcBCTOFUlFZRh/T
yvKV0IVWoI2Ye5vMxHUZmX2CM6gOjjf8hBFWEzyRPkQcDq/5kBMmCb3M+x0D2k5uPs+E5MK61c8k
DaJxMi6aGWEUJMnPu+g3/QwN+SLfFDE77pOj7HvxBFEVkQQZqoKtC6Vq0Q601xtZ5wtHaO6TXZ+0
zRz5fdZNCzcOm/oSD1Bht9DR/6y1hMHI6+1YPhEJEfSopu3RxBTkoFIMExD+J/cZwYFfhOiujnsz
sEtiXE1MsImXVEEnTDu9VZ/xI1FUIM4VO/crrzXftwr5RNdJwWUDUAxpfCqRzPyPNuVAv/NBCANQ
rrx+O0PBrzGzInsWI2ESK2G3IjaCGfP0k4dzXcTJWcwlWmMZ7CEWhRqbSXjRAx53afVJ3rQ5wKAT
kY/S5ftAiZ3nA05/yO1LCjrC9q7Crw7xFaa4LIBUjnAp0JO1lNCNov4O/9H73QpQTM0a1XgRvZMw
teIlok1H7RzPx4X5UFaKaJxcHofP53ifN61Hz1WDgz5Z7uBT/f7AUIhUkjnBiWt1o14PhXpAqqLF
iHtlbNm1VINL9nx1sabuKoAepwgpPBSKVBF97FOEEQgOv7QXbgJ5iKUtIxtzCLOLw8KHRBuzMnt6
Ra8PHfMW5e9ZHlf6ZqyfPxIGKPnCqWiYuLovvcsJyN6CIey3Fknaunef7D7zKnOfYG/xgcfq8rdd
+HvLzF0EyLFTMW/Kn72EYdCQIJUufGFmtsdnYG+bD6N/X0t+s0h3tvwGEZ9pl52mytjWmVq0WLZW
2bl7dTz7Qw6277hh9ZSzCr4c8LJyO2tc0jyxlfpjZW03fgoaDuRuoXMv77fsCluogKkYIxwuebYD
BxUlRqBTHiAUhQ1y2/xp2hUQ+2uNvioratgtr+lkLwkDKSs5glbcbQwIOPE8/56RxUHG4uOSHqyU
GwWxz4l9bVHB3uMZCtN5Cavqs9NhoCbBTbIuhcHgdeUd1dQO7xGZOVx2IoD+4T9dOv2b2lDrmZ1S
xMEVlMkjXsLCJ/wTWPa0+BCO3ryX8TCU3iwpVttPzQFKI5Jp+Bq0/anlad/YZjs168T/LaZH4YLh
zeXgkOaSk9ukX/JfJbveP5dMexxKppcf78IQJqUIKb4dixpLeMp+lDCVhXgi1izy70gTMMGwH4wi
xEP9MesY/jOg/xV+aDO02ifAthaBzXkyXn5+vIVEGE6V2CBup9msLQyj1D67ASDgy3DgSN0sjGKl
xMnIsQiYgCsSCfqk3qaOOlb17sugCVzTT1Gt9Zf9D/2GUYRPPqXeMLOjz44r/7iipDksJkEdEzPs
Yw1Otl1HBOTM+V9JqDC8KibXK8PNX9HIeJIXL5i1wHtdJj4rhXQBB8eM+LhA9o5RaMNXICrWJCCO
8/Eiaz9CPd4HR3UdEqwmz5ep6EOvOFKZKR0qGwBg8sWiKN0vjxlRYmeyTvu2CIn3eGicAYKF8ZZq
BqKtd34HmHTEgTRjsXHjUDO3r3vkUcHOfUvoFTKNV5yF+loV7ks9CtlRIKbjwoXF3zj3qfi24HLa
rIDNui9vs6u8YI9wLJ8C0iDYMnuBLQrG0NBGlW6qS0g8SJYt73k8d2IVN0aAysCMBTW4OGn2AfNd
9bPLjCNKSu414L47y1QyE3//u6qpnp3WbK/RcpXjwgwK+nj2PsStgYi6dE92+dN0YGwA+suYN/1g
7Tw0XTQEYE+QGm2rdbXJFKEz6go+yPxK6CyVt0o5TwGVkIjNmpkzgahrN33F0BqKV4YADJXx8waz
RV3x+NCznFAMhto75MPTOyew5PvXXw1E3bEFq4Eye5qTJU95wgZTSEH2fKSS1JhD8DTQbva0jMOy
cKoNvmXprTA0xuMKObHIrkO4ca6/rjS/zjEr2Oi6o6EOEpmRX2M99QHxL+U+6Lvgf5iUPSi2i6Zr
sq9Cpb9u+zXfX0LAd2n3OZ6xbf+51v+g6kFv3+qtaYJ1xxjin+51YCovgY/2/YP5RXosn+wGC/ta
TXUB7aNM9QO5eGXesAb/94Q+jSZ7Nltm4oqHq2th7xnq6LjPtQRrbDOi12wSYFIdiCyE1YVX7WlX
jgsvNNbs/kr9Sms82v0C/VQX12WVYQmncX8mvKAMNN39nGXpbWJDA5Mri9HDrYeCzh2saqU2+zsg
HXg02tCAX3pZCLLPoObSDAcVsLGUB5bMfcFcKzahUOp/+EUAmgJzReSuXdAeXZMQvlmsikK/kq0g
Nyrf5QW0FYncoapWy4gkBRVXv5yIUuE0KoprojbXMf0SOoruUO2+PSzbebwYNncKW02usocSAMMp
misvie/6bF6Ioht3UlY0ngN94FaZneelKq/7NsxrO61jK/f1quUJyCesW1Z//X/r+KRo6fjATv/0
vbybifeLWPSG6mCqUwJ6zJ4EkEeMN2G3gvx8d3yJuJd2me74Y4FrxNlH4Ytx/2e0xHhOgeqgMUjh
v9M2BnmM8crOlEiqal/p4PFBl1Cr2GD8KmAJN9OD70vqwihHFi+uZ0i6nWP3+jwEf5eEDpy3z9gV
2Om8D2NLqWUugg6vR5YR/Ic+sP3pONAa3iCao5DOxxZHVZrmsK5EEdtVdiNYtuRyOkSL0a+hJAQ7
tIbe/YLNYUS690elDFoJbgmGHfeDlsbdq87FLFcu3Fle+IvRvjvas29dDvoCxqc9LZv5JGM7yDVW
R0acst1Ig/4vjo/z5FMdy116r37XqUfUK11go3zFmp5Ij4d99kd3PH8UWE9q6UUuFweG44m3n1Tm
SW+zJFx/TJNEiQJVxykvQH8YdFu09U9CSKa0q0AD0V02CVjgK1mCKiTIgxJopLILni8qPER9+/dw
PL9xfSB9rKLEbZM/SeeDATBDXt4D+iJ2bRPDIpr9DTDS6knZBVNHdL6nNqyjCVWVDfTUDm1BMxsP
IXvc7DF7z5hzrqKhDdximzFqHdlWXr4HpOQ3HRJEUvsEH6KO7MnQUd3LpZGwlC1leDOokDbnvQkg
3mKR2kyVdet/VHfwnBVKb0tuVouLXP0WPlKGtIiiTIAMLhKjq1pwejPiyZJlzYsDoB4yJLZ05d8c
K6fn3gCxobAnPwQO0jMiQfR5bZRiGaxez2HT3dgULis4bAlmNksjikGEjwlAkPPD0AijQ29koDl3
iTqECs3O1gcgSoJbFDlcoTZ93qB2fFtzmPVDjfvMrVzjG4D+Vsu3sEW4MCh1Maspur1YEeif+Eih
ELkesAwW/C+h3GlDk2EuUjjOcUzRyg6GhhSYFKhGz049IkSiQTxZ5HFcT+vJsB7p9dqb1QSu4Igm
NIRwtivoM5eJXTiyw0ovka83/8DIBEqUNClJO9gzLTvmYdYdoynAzFFW0xqC7sb8RV0S6AdgWFkI
KAC8Kq5aKGKKnoDICqMlJ877SNNJXNFLjNCkQDXdHgK2kQRViIzKQ4Pi/uTrhf9p080CmF0dGDNo
aXo3vfCMEQ0ajaFMu4u/I09B/G+YIMK4pbilcS2keFd0B3SyBSKcbibzFQNUsZaE1Z0cmUKaZ866
jIuLbJer1YEPJYPbCD+XArjbf84FKEYJKx3f+ytSekkLh1c81GD+TjrprmOdWYhK5X7rp8r/WEtu
ra7M5VW50UfWPO7h3+aibZP+UhAsEEtrETkjaLQ/M/WHi9DJFvqf45FDDHBgSjDhxvzMy1+AarQv
gmE5FnXWEeATJBWK0hgeDs+4idV2RwMqLXjVvQVZAwkHgz18A2whlJOUyrcZw/wwJNavN73a6tmE
FTqhBroretMPAUf4nyT76/rlttcMXIlPDkn7rm+LTbdbHcHp7Xb1ASw3yPeeMah4BnnCZw1KiEGi
KSW2MucvK0qj25PISa3I0oHvscuc8muaFSFFti7VLLUwrgiqz3Br300NyPY8mei9yBw9kmTtqsPP
FGTlqFpBMI67g5e6+etX+kghyakultNWupuV3zjAWAQXlA1q8MJLIj9pNHUSbpYj6wrCVB6XXOOt
KQ8kaW1DqfZ1toBw2pczzr9nMSG32xc8Ofn+BSgCqN6FQtoH+3fZxUpUA3voU3PU5lJIqn4VYeDX
+cQ+1cFPrhaPIITR0hlS28l7H38/o7VfAoY0rNss0YTh4dZketH/y3bgAGSthQtojGhc/7pftaJU
Ar9PRrWGM4fSto51x81w+w6KtdowVpL/R/XR41tUfm1Ow5eDGjztGCc+M3/aXwXrIpCTMDQxWvl9
dGaXcgV2n107rQN67AaOU0XvC8rYtSClmt7Cd+fwMg/IK5xeJX6PBeOBq7zHrgWYIx8xwjZ9ec4O
loo93ofmFvkyksPCPHQo20645ywiQiTOBVDjdhyw9pfDaH/a6MvgywYq2+qDi9baBuNlpH5QTion
qIMKueKadQVXLkXwxAb8amLu/x8xuHSxFCY1bLlrrqGtFdkbB06a337XwEGQm7brcmbtLGoXANaM
aIeydjD6MMgTrxoVA4mWIRtR5OZSIMybFO2p5lCfKIu4/GtB/oumumQTcgXZlgeq8sy/qjtDVzVO
cTg5/RwjoVERrV857ExeJ+BZ0glyG2KHIxnC/llryz+JQlcCuRiSsYQg0oLlYOwdJcTicdYP5PY5
MbhSRHsmg+9ZX7zUBqisUHdc9gesx8E7g2FT6lEDXkNf4+vfozQGnOsWm4iFPbXQDXqV5Xnj6psT
0bbSHVi7mv7aT0mxtBkZMg8bojbeVnlUFeokTLwjPuwLn00ZjM0+aBiQMFU0u8p/9E9kSOW7HZBS
7kl5SwX7rJCU2n5cDYXXd007L5+g/Rc/sqrl92jIBloZh4RCIHB/8qwtkCJ7zAF7he0DxyH1ikBA
OqbXPsEhTqycC8QL/YX7pBawPz/cia13bekc6YwrU27AODMr79gLLpwPjp5xAHXIMavqFRl+QG+6
fi8LVF4YEIjbMMulWOOV6dA0GnOltXNduED1HFK/wooroTdK9mvwyrKuzq+RNid0MO9sPKR0kziI
X6naMdHM39MDZdNorPv3PXYkg3W1v80t5dLHoWIpf0BDITMFXXgLyGa/eT+1i95cNGXCMCD6avA+
Z483fNYcj/87PjPs7f60uMHn/Nx6BFHSAP8XInDn3+RW18pIExwa3TzIzNODcfBszton06QlMogH
yoDhp5WvzpkiMjQRlv3jm4UPfjs5lCH+LbRvAKLsgpiGtIRmLrhdgZ0vOJU5U1Kb3X/ZWcHl+MDL
Q/MJC0xdXK358PxKoeJOHl23yq44lUFC5o33X9ARWSpLYRGVDJRoCP/2YxQrpS/lUbRJZk5xI1eg
U5mVZVJO3dBFrCFMzI37COrHJ2Xc6F+BSteCgh9SvmnCcd2V/tAcz4ZQaL8y/YVZ74oF8bD4BzpK
GH9C9XVrBqLV06jbY6QQhxGqgJwGnX9Rx5Fmcdwwe/ZDrKI3AHcJgWCWO/Pev03C65w6kIYjo4u6
R58pEHBzx9vF3i7LptMo4YLPX1boPnD47fFhG3WtP9/0RYIpcqdOIyIcVwLeu9gsBLDO0ajhxqox
YXnTEWFcM/6pIhGFeavjLSEX1wjmXk2HQfOBQlf5uxR/qiB/S7ZqG6z7DFzTf34VY1I0xSdFyBP3
p2wMXtN4aNz1yFFtvKmP8E3/QKxT9OHYSuwruIYbN+cAq3uyPCO7PY8A2BDSAyqdRRJFFM8N0Cfx
G6VCw56MeOQXOiiDEGzntKRG90jZeWQtcQw7ecC442jtHNbgWFNDzwXfZmjjdlEEUOwRATPZSTOj
CAfklzTflJo1NC0J4FmV1oJB4Eud0n91WWWNlCPL/HGKX6fvCemXMeGwRB4Dl7ygDOH5joYX9IFf
qUnszXMa3bAK1owfbONb6tzOZOWQs60BHz7E78pEOFLq+X1KA/iQ2dnJ2hz6Y9J3ibfUIUsEQ45K
88voQ6NY3ND1bBdYqgxSGIgCmD6zAKunuQ0wmfuIbBnM4HTctUrIqDql7r7Bj8ZcXgMTVzobdFm6
J/GIMDZ+7yU84QrfanSLZmgFO+A7oKC9dGKUxqxw+muB6t4yzlbsEbZdrXqdzQWsKwSApS4e4/iu
/l6f62xhb9XCcrm11VaV8LLyCd1FnIiJeuU0GDoTvgXoRsx0ica+3XpH88pV99RhhIAhN1HrSp+U
R8VnIIuQSBVCbe9D5bYKz9AKpjDPVBKOB/yi+cCTDLU1KhHZP2afnmzNxwQDVrB+Ge9wHVYgJzi7
eV3EIhqt2fIxpcDvZTxITGosiNBqg4n5QV8Y4FatVHGsr+aoeEZKJTUyUw99rREpjB/MsOB1nwhe
AolBNE3pWe7BUjo8Y9F4WKN67rg7RNQ4UmfFDWg8xhdsk1Uc7Zny6cY2xZRuQFdjZBUE2vvgrNYu
1UuDUpD9rJRC2CMGbqXaNaUhmoS3b/pdQqD9XEuPCZgBeh+Xk00A8oJ880IO732L9o/wU87hWjx/
LurMXf4UO9V9R5zPfOMT6hPDs2kzaMIu6q8mDLeyWYT4wm3kqy0zYWsNmsOzM0sb8Nptc68mDutm
n4bbDOCOG+ANXduoctDauOIOluBQ5hhn0MM6X6duq9qHdUrQ1a3mI6KdvkUQaLqrKWKNv58UJDM5
McBMedR+XcHLdDrfHu47Npqlzwk702QdSml9MQA6eqT0CKlgbwIAcixPnv78qxE/cboJuIMEEmk8
juIe7Y9/DMmBmwrx+8npjy6zJJMNGwlixtH85m7ao2biNSGPE40or+TwbObW3WmImZgQ8ObpwyFp
55m70Nm+B+hBCkaRK7jrf4DM/yEEblxRgZywxTNmHM7h7rBAmcRgdq1JCx5ZVxZJvFpgRYaHKFWm
R8eVgA5I61BzWuFOo+yfwUDAnds450Ui4odBKMVCTZx2Vifnny49/bX4q3D0vXBarz5LWZw2YBPc
NTCSCAgRGRgY8UOXDJqNmMOL71fVvQrVfDFrwQiniTtNidOq5+NlEQ4OhzWZjk0NNoIIxL82hsiu
h59qJyO79LXZrGH685PGhg70c8GgQ7MoF93iNohLO8ZhpzTK9ABxRQHGgYLlDcTlstb47ImqJHAK
u6wvgAzbqUF3+ZWCVUQ2wIn3ZJyZP5PmSQhmP5nAR2MJQu5g6c1GLhFxbIOksANlQ4EuCxkroInP
EGKruQBToJmBFkZ/Jy4FwcxA8ZoEN/5NlKaB8hnoIG7gRxDF54nOfcqIEWI7Ux5gI+fm0X6aXChn
lgNi7s13sTHwUbTwgA/ddg3lZtojGZtr1I0EwK2tN7qlM5qSnQI/8e33jbp13h2yv30Tm6AorLSl
24/np5QR61A9wMa+RdzX5A3ROXBxkiAtd3uf5zk/cjK6+0u0D4U71wXBN896nxL5Wm0I0xWI9U90
pleHwPXnx3WGI3q+wF9hGlH3Y302+bsAEvYQ+2AfAHlx2fs69bs+6X3NRHi7p6yTZ5XFNPfZO/lb
cP4nElX0RQVeiVMhQWegnc/QIlXyyEQxHg0Nzz9loxX/aBv85jxAseK9TINBtn8TDyGWh0oAjzGY
4zhz6MjpxAuwD+2bhz3jlYuAHlLqKZQiC5dea6icP50+7VWF99M834hwj9I8AsRBiONf2vu9XKLY
G2R1iFz5T5eLRgVDtOElUYPmrvg1uD1eoulMx1XT1+zuhPQ/YDLWlN+0RnFAPMy8qlba4i/EEm0Q
mGcq3kV1mD9KFiUxRqR27qL75KTr1wq3yhOE2kuzfFjvo4jxOO6wZ/LNl5kw9iGqAyjU0GjWp7g+
ZjPfmXBHxayxRx1KkbBeA5cJ5t/gmOp6XGghC8BH+UkBPglfDtAm1KsBlhSn/YzwG9VYhuEeYuy7
qTALG00sS8rure3cPowJoQP7cAAH7olSHczE/PQBEwQcwkQfucIAOHLYCfz2N1qrERkotb3/0A+3
cSgpjjTUfrtaEYrjAFcWoPkX+d6UjApZXtHFDPLcmPqx9QeWheQMwV5OKZmMPpTiMqDwAKdQFXIk
IRzJgwDn354iFY+UF/XuQ7tXnmKRt1rLPoiBgwzH9NxC4FSe4Ftm29+fG7mDOWp//EUFbWSZk/wJ
91+e6/Pdd5rmi+J+UEyJhdGnuJAR7v+1kn7XFKe2hq2qJpcKoxP9W7tMhHWx6r1eW7jkLkZEcMNx
3uVdgicQtX8J5d90yh9vri4Lbst90d9sAUcQH4JHBc3plSvmjH0aApQUsnoG9mHEAiUwZgUVUiFS
CuRM/J3GlhuDJ4bkfKVzvoSOJZrt7J/dxpV5wY+m1hiKN0OGTTyG1Xqj8OMK5UVebL+hgC6c5BvC
lUAdeDC1hfo8X/rOkZDIkalXUSRebSDp0Cl8d9AAbMkRSiKGTpAcl+JW1r3viFaumRNbjYJN4rWn
R6P1epk2/apEbO2H+natplfJwSepzhdodwWN4K8G0qWbuH2bkoNFtyMxjXcL5+cF2ymQLnmXOJqS
rXCMI10IUih5cpZkIlqkez8uFTznF+F5d8ynQyT2HIrEIb71RaCXHgh6y810ptAZOkzR9pJnqjMm
WokwoqwO2zMiVQ7kKbij0QJk5rMO8VlaV/Zmv8F1FwQuo1kvzSC1vqso5heDdTkHm8CT3dd/OGld
l4mKkriXbB/nN9shsPWMdL8TYqvRgCFpd69syovbmEMFWUtoNqq3s23r0wAMnoVjkvxM0TzuSUWO
8YU0pJkaDMrCj1e7x7VD+XHfFiP2K1y6qJKKDNwqCAuqIEkgFGxjjnKwMwcRhgssjbny6K9WImnH
OvGzLLUZbaEKC2EcKZzNq7E9RTCUiS0pzL67x3oczI9AtQFOgEhB8RgI+UXl1JSmnabL4Zsn8Lph
g7i+YXpiEW5loCx/YzOXtfhm3CelJLJqKKbc8IFhZCbALk8la09aczekPQ5kDEhG6FsO0XLxnQB2
HwEdKGmYW++IK3j1wjqV+MsTmkXRq9ptzTrSdU623RxCoT7U3Xaf/rfchwTY2qvsAcjLRkFlfx/M
MkIfS2lzhYN5WGao+PlM8qKQmm23rh5dhjfbHzfeRtDaR5jlYFu9yYDFQjUYesKZ3x5/srO2va82
8ep2UFc1hvWs+I4I8JSaT2diTtTttrQU0yP5UjpuvdY/QMCOQM9iDpNX3kbtLQcxpvzLEEavR0Py
LvGBVdJmJkWzGckhrVAapgU25tJt4QviIFZpgFoa5kl7w9/sTpKOR/VnfsG6mq2hA+LJ8xR+ASE6
YxgAmJgGDWNJHZBhk/NTjDPE8Fxh8eMzJOQFUo1InBc280lukLHIb/nE3lT6AjxZZOpJkGQNxNJ+
KL+lTH6Hysa/Q3aiIzyENBDBy9pI4tu3F40qdZAMukVUjtRFUg1V8CEth8QzT1hCo7uf1fQ1XokZ
JzLCwU4556jgArPmIm9RuDylk7+wynkmq0IQJJ6ddmyPzrWSvmMiQwjrt6lVJQCXMIGH9RIvQDDp
ziofwypkuBFrZomzAX2YGw+SvnD7VRdA/88mHh79uROhA/it0DUIVav9rAZXzMngR2NDtztEPBjL
zTUeRBS9oKLj8sroFLS9t4FYtbsiBd72HDnVJ7ZRuocM/ky2/UBebRBVUW+LmBhDaOQ4duyRVVXI
N6Df6mQAiK+i0Mpct2CUrVb8haPnvp/DQPyHnxHerwP8VYd5pRSXZmezzo237eiT01niSmUx9JII
2t6FgECuBfjVA0hlO1RvcZahowOJObVqOF/O/Zckpbe5nwaTzVrh+wOguuFhQ5Z/G9aGWgvzlxOM
rpi0o27Rp1h7cEvJLcYLqshGuf7ppHyGtTVqwzuuZvF3jEnXr/3ZJMv7g0mrPmqZmUtx/krHS7RG
tAirlwEV3dLal2v1vCrrkh0aUthVvbNfqEOjcY9VH2vsuNRvnp/MirkAl/pLfuB6UtDM0JMvfewN
rX0ufwrJSYBhCuurOv2K5sjJoCKJMunQRB8vGBAWy3VaCbTsSbWgGT/aBFDhPqjZJN6HLSnYTWrE
6q4QiBRkq+cHctjSKvDYgD45/g3ajP7gSpbnbyWlfEUISP+XF4bKNTfGPf4r8jA0p1+JzqVwUXNc
JoJXdvc1f3HnALvcL1DXAJemBYEfG4ZU7RDJP8BzZtlh0akLNG6YuthLo5RiwWYBXGws4v6WatAO
4XKBxHob6XqAZeIEUyQ6iDNV9UkdwROeYcWJ2o4RqHkdgKMuKx+QkYUxhTRdQ1w8F1936PxhwIdB
U06uq07f9DHpHcs38zg06ZQnJ7TGB2Hq3dJ/WH6bRy+WlfFCZ+Kfbvfoib1PS7SwNkk/i/VTJ4AQ
T7w/nMiYfAiRnvBlwrQEkKNN7qWK4tQcIQctqjaDXlDgnnBFvnuPw+mmIXP8XPROJYsOCh+lp9Vr
JKjW/AGYa3ko7lCJQKah60jtiss9Hx7htpj1FYvfytdp/4DPHGz9rVeYx3nuxoxAFa9gWiqnUEIR
eAOJkrqS/rt31pzT0sFihxPcFHlX9kAbMDWkFy/QMedY3jv4+zHst2V8uB2m1nfB//7JIfY7a8HI
ranKXhaHtcPnJqKTiy0pjqMppszzDzhCaBFKG4wma4NxOJ95ddKFXSRXZ8sdL6C9m4jbP7aa9yJd
Zz7fABrwEe9/g2I0kljG9daOAN3J8FnQtM8q5WEI+OddVikZoo25ctvk4fBIMCDy1oB7yd4ALrZB
ShhPh4kOgEYG97UFO9la2MlW+wXJBLOI5i7J4zUC/Fc8IJ/z8KXWDRrJOoRL6tZByJ3bxYzLjMhb
z3CdeFAt3GDSMhiTIFOqWFc6AUACTfVXWoNcnynYVpzMtcTrzlQPgW/pXLz8pKiA7hEOl/OFhwmZ
TpKx37pkYsaY56pJq2+jmXYt082VOL5oZsT8v+xEnLN/xPTRFzmNJEhmm3ZsEfw+BB1x5+6Kmdxy
aYZl+shghu6UlW2qcTUDXC2UOFtYRJfpQoHqU4t5zqApDOWgsHQjrbHiGFzToSlGWj4ijXeDCcS1
W8uamIR+vHaetlvYFv0axj/h700g026mM0dCUiXtJ7J7MMQ9+62JOSejRLUXgCXJXeJiWtdrlzkx
CSLRiBgJ6FBLOcZZgsYaJQOlczMnyXmzX/seD0LchOLNH3h4UfJSeEqChVE0ID5WcYXtHDSycQVh
WTwPDjw6jX2OQviLZ6IPSopKScZ93Z/s7bpoDo9G19ioPbyqe5gxlDaBdhfXNIE4ni44gLcy2g55
F9L95a5hNgiAKrzs3g1GvN/amQamakEZPQaUj+cUDTtX8ZieHz8wkaHjcCxFRj+yZbN0to4iRhWf
rX0k7ok2IqTr6AxhYjv7IsLhdKSvYH16j7Pu2U0Jt4INv34ZN5WWTvi5Cd/NnmjWrO5NEvT7O3fC
pMXrpJPahk4/KGkNK1q3HBTPp7ED/6iywoM6RRwa19WlHYpaXsn24S3PaUZkFdWDjZ17SjWwjMiJ
HsPCUfd5toy8+2hPDtGPuV1DTvxq2JhUm9LrsuOVDhdVxgQh2N6DkPpjzUVTGg6v6RD+FPAg3ipO
BpF6wQ2AbOI9/4HDxma0X83aXeLrGotnfq9j/aI4avR/ekl3/4ewNvbl6yHBxuUVXmue4zkc+1dj
5tElNGgWPxf7TF4YPpF+uVLC0LoVOmQ/hKsSCj60vkJVp6cJkwsOOXojuNPWThCfOkcLi6LYxgDR
ZGy2+UQUU3CqFWboVbFJn50HokRiE3LIVC2FG6ZIq86mUZjVl8kq89nUiwiYX37eTgoOypPH4ZtQ
VQwG0Bh/MTyjzuIgwxRbCPpgkcaYLDhuG3vqHlI/fMiBLkXW8ijf3bfH1NXOA760ZmYVodBItf9M
+s9Fzsnn7mvlRuUz//I1ZGL400/xuklSp27vdZvvhGMa9xGDUdKoc00r0f7zekiLrkJnJPX4iHI1
dXwYfAzIEzItZnjqQ1kz3VNsVsZwD3JjcJ+RbJ+472f4b80u9OH2yHyKJWIq0nDIoJFsLyVkj7UG
Ti2ibiFhdVO73evAF0TCwqn7YDWSAbKrf6TIblMHOYxTq65aRjtKu5x7z6gx7e6D410BHbu7+/TN
dsJCIl0T/RumtebunXVFNN0JyiRennYgIYB46/UDU3mRO96+oCM+XgiNt/lsS6cGXqqxbF+ttG4q
7hWQrGsnQxkeQOheYV7GeSWHqHFmIHuVjUdkYpSxh+grFpJSV2RNRILw5qRd3iWfBmEebK9dr5bJ
9rm/q+dgsQsBgyaOwFA5PwlGqipOglbvaV8CxaR3A2IcBsadEqfhkka7V3kVYywQuD9u9sZ02nAR
h6VkYTZrmhe8NqmF20Idzn9Hh6BZ2mULVMCYjLRqAlbyFoqLU7BgAHwDrki3iYFCaxWcebIwpyIe
a+XTiR2WfktMPWdBQm0x4N5n0beklUr99EtbFOGWcvCh0iG/fy4460VdNe6bLcDbUR0rv6FfcRii
ZDumGQhr0HZ3zwPr0Z5pZWWzBY1wiha5FkleQ0kTIw9Cp4ICwcWy5nFw5EvlKHMerL9dOxnQkrM/
wsXTldr6NQiNCZbOQDt82iHwGMRZZym4ByIbsbAQGYI069sWQMCrkKPeP9vchA/BCQN21CfDbEVx
YC/OCt7HRLlI5cEVb7dibLvjGGcjavVXl/RPw4gcNg7qzIS+rf7Z4p79o3GI5M5vjlhQh6mujHUp
/jbnhN9eNJgMgh21gnxas+3Gi3K+DOxV+rZtyW1LYJZYeFfOheQqeTaaWMttCY9cba67vOXkD2fj
PKFIMY7C5AHooC5mkRW9R3eM7hDdWT+HykCjRCaaz36aAtBFlYJ0EmX0NYlbv15KOFs7x0PrNdc+
2T4uB9txpI27agcuYbbhgZSv3PYecEcNHQSLAbSrvweRyFDKw74w1j6uVsHENcyN94irbgJVO8K7
jaPd/KwmfX8h4lW9Q/csPY0y0TVOkm2Wbk6piSBNQzjwb3v93oKX4jfNjaYUPEL+z8DXe35ilbUX
l17Z7juG0AJ8JlxvyG6cuPJEd9Cyps96ybqj/B9zn5DFZyQxXQCrHG+uojAIumO9BbxL66ZBd4VQ
Pf9IXRs0bgpkmt12LRHq1DB7Zyr4EIopFp0ROPW1k6/XalKjBzfCFt0woprpi1kjOQ+YVY1KaADm
tK8ULx5pz4myD35LzXzID2PYad0XUVXpgurbaOVDdkD3HgsTM27SrQD+gbP0vP2AyTSf3rOs/uBN
MwBkRBY4Dv2ZomfjKEUp4HWdklicFVBQSlp9ryigLMRMRiKY0a2dPXmukV66mJuDop9uQfnSYp4c
Eh5xbJ3YK9lgT08RMShx50NUxthxM29ATdcwx+v6T5Qqop2czRQlg51+xRXVmWrbJ2n+emnMdX3P
8PpDnkSylJk8B+GYbD79zwka7XOLTLwKU3RLfh1XYX6GlZh+0fu9uhxX20tYdhZ690uMHbrV03Ss
w+oiOg2AUXhDtdiAarsbS8rYmJRas1YbLTdlw0nrD0516FDflLqJ7dg/Q0ELEw8HjswjTxoOzuXL
ejJgwvpc5jpEpTFLV/UgaVa3AATldZJRwYj/Htsaue7RDqPgK8DHkrQhJLRVV8l7VIwozjU/LTEc
OYrLGLfLiaxZ/R0xNCYmrY30hWuk4U9FbtIUiTvjsWDuphtTqDpQgsbAeYPT+fC0IMspZfrYJRP0
T5Jyr+fjV/gwxbUhCzQgcVVp7eTfTtR1BnNPjAd4SCbXqdWzAnmOt2MukMaunEPS189u5GSSh87g
Dmgt/fWNo6BJgluPbPcwvM9WXZOkZ2qzczq+CQwwi3/D6W3G/uviFSMeOhzDKmhNB6AFwPav1EAo
EWMNtPhIRopwHyBLFzXgknIQGogVO5Vo2d3OY5J5wLT5W8bHBb3x8ewmxCi4CW1bbYmpbpr8NSQG
wWYHfZxAfc7b2e/AmzbAm5DCx3wLVIJ/NEGCCXiAl93RUmTPjLAcROfwASNNK0M0RzAupWS68vZd
PEjj1SM/7ApKc8uaBHAPd62sweGWpjnb6RWU7aI/gFQW63eWN96xHRs5MLRp3Aaf3m/FCH9qNhxB
xEeAd4RELQzAbv9gwETktV2hfJHvjanPWcn9Ch51zzQQ03XTQReYKlK3uihRQQWwLy0jqzstuLka
GJXxcjZxhkST1MQy7/9IH1aemxqgkLjMApilviXQXq3CuahtifCCkxwoteK3pCUpuZD3bk9I59D3
8tSyiPsr5PkTtTRAO8YfqTquxUYWbCnCrHLN6jSbxrRNl6ugv3I8m5/CrJCtwqbC/WatvSLC96ci
37ujMkVMP2u9OUly5LTJ84eHMjzi+M5Vol3Ktst8NJhYPBqwjTJ0hqTQjGOhhYV+ty2RKlpjtFbR
26h4Gvm3WLXtHHwqQ39ejj+GWk4cb2dCXHdLr4yYa1YRH9vomOgf0byvuhnpCwGp59mi64fbKbnY
IHqsWVvz8W8etGCeqKggwmvvABF3/f3XEExzKte3EnCcJhriau/0EXHwlwOc6RTSk7OUSKMbmtUK
bUx1clcxxm0E5ZnrszM+atnsU43ABV12AiaVT6P0TBQR8sLuXrTxqEiIcvIN3cl0SrQ00sykJVQC
knDKsFDZzdQ7JLAlgBIp/+HuJNmoqzM0cMomGeSFdJ4UyXmgUZMgztJaDvsEHnXBRBkaW1gQjSX9
ja7O4t1d4p9LS2lcAihXBi8NTeRtKcIkL2MSfU2ZTPqiIEjvqFuAZVwBN7sPtZbxouQ+7g/Bq62u
OgU5tS+RkSjJekILwvuT053k900YlEpb1mpIglgutxNTlGva/92eykKluMxbT2opHuROkW6L7W+f
J+Umecxz0azwLb8zQW5bzyTPcfbT2bt2ytckqepkaNgfVTxfp8yNOp3Pao3yF9iLAMOfVnrAZYGh
iFv7ce6YvbFAdizgcd3GnTh2kyMMJhNAiwDxjsCoFle1zELw7Ias17tZwR41bLwY8JYrFVHgkDgZ
HzfyzMS7KXmo5bnQ0JEyAcm5Ofyeo9lYKH66OUnqMuoSsxt94+ScQLf7xJSXMGxjsH9acXR3VbjE
qC88asP2NudSgZhpS8ZIjhlxeUsyUakpxKsKCqOuNF12/U/cT+XZ5670bKxQkvikebD2YMDSjm/6
K5gCq0iNrkLKyM8KPByDJJOIRJaKHgMccBAiT6NEqUXjH+sPGJH/WPt+jfoJBFiNk3VxmV+mopkt
6hHkHsTwb5tB22Z2vhnPXNghzbzAE8H/abKavxxGd5pkGOJHWxszzHjpCo0vs3ScMnGAZdeXYVkn
eHEoq23jX6e40kdyE5F/NfTNz1ujElaRoB4S0bUyoGfmjoDUoitCjqwf2u6y7mrJpzOAXbqUc5uh
LmvBTz/psjBIHV6XXule1H3VMthyuxOYa2nJmn4N2iPpbExlZmajOKn0/wJygCoZzOmE5GPc+Hj0
HkGWvuLhLhP2CbvtABS5x4r8Fd5Lfbe8RB7JLtaeCiXcJssXisi3a2mfsAVvOZwbfr2zmjg6qglp
TvWA33107SKeeJHz74+s7sE+QOimX/UGpTugaNvYuagFPT4AZUIoRyT8r1LxzE1ugHtcDZzbAr6m
P0CkkI9+kHB++qiFBEvQ2B7/mgFi2OnZOQNRXY9kGdQoO2XEFRMIGpUbs5aHpY9Pe54dqGoIdVph
oe8LwFpPIMAvfDFDBZaJWJTU/PZFdU817GEJz5u24GjkC0NRIgptUhnsVRXRSVXyrrueCbQ33iEs
t27y/XfM9D7JdMCy0XcjVmnuAj2WpSTvbiOCn2kdsgC36x8QT/gFh+Ec/xk9qtJYeZf5wSZw1gf6
ObKYCnZYD5nNGT42FljmQZddiC9ZkEkymSuW3IisfVoExE6aFc7ebxqwwBCEgdi3HCyLjbXBWpCO
pSliLeNkF6W9hh0PSM/qSqlRaeqO1oyN6fTfFP5OOcRhHnOKEh1gsHTA5OLaXX//ekzIqGumRWPG
k2W2BQoPTB6XJnSXvXnCakHlIe5HpitLIwddx+NKqTUeCR/rPfAyR9FIOl+jZ0rNrTQ8gYTMOiSr
AxGyefHyrwFs9Z8wNfUbvZ0eQMEzKcR6jC9yBXsOcXt25gWXpHqie0LiMwODlIFgfKOnR6Bj+K2c
HimfgEyjEBXai++43rxF1x/CYUGbfzM/TriUHLMpUfs1vcQX9YnoHcRjrtNnBu2NFnZWeJF/AMwH
5JLVS0Gja1EycA55cOzQKOYwk39yTFCfBQKiXK2Z3PVaSVvlptYiXeNZQunJ7FovFswbkewJkiSA
gVufYICCdOZMJa5NPfR45bVv3KErGz2dnydzzYljIDxVGePpH553qwmKRycyQSgTZSe8yh6szIjX
azwVfgV0jMX7clvrSof6bSmVticirbyQPgdEU0ikKN8RHKf2kMj7DSeO0/GPZvBsnfGCq4PZaHV0
KH7F3bErFfa7RgmtfpdY/qioQDwBBGDlnemSHVSBTr266gjsbiGRlCeyri+PV+lsbv2XvpAeMYJs
GZuS/KTGY55O74HjvWYmm3iJ2UN2YZIc13CaPYyMHMZbgrUJig2vwK1CUyLax5L77+TmTZYvITEn
Z/wq+p0QYc0UdcQhVcDJjMFMCeObgb1PaCc4f+m6jKAGP4kPXJShf1ROsEEot2OGSIkyihIgI34C
aL12xvZQrk0RYRrTmPZUKV4Kfdi+fjcwnTnPOFuCbYuj2kYjjuFb5ZOn/8GEUeZ7bXR+12BS7LDx
UPKw0lgsIHziEDxBIOkbfFw2kB6mL/2YcMuma13apC7c1dVUQ/cz6rF6mizGL6NOsz5tUM7PZ0KC
QdN/2aJ19PHUU5pw587MvrkR0HpOl8ekmSkLRiSZzFfe6/iFNpOmk/P613pXnIGJpSi4tagF/zhl
qyfgqFV4xTqid8rrFYUFzLnyR+za3vOytInTKZwhihBKN/Zlg9CQ8kGp97Dw9sUAqpm12MpfshAG
XTV+wr7qgQ8x6PKBKbp5ht4rEIDklakQ20fC5TyVe2XBZugHLIVbSE8RGUG6bGTr+xQXXqc01QWv
9cMFU8V7oRzzt5d9SCdnsbS9wmn1lW8mMPeDx+fD1c67p8Viy3Ok/9GzpHrYIj7PcLP9rvaH5fw8
G1PWaU2G++P5pgGoC39SlYCFbTwko53mvbeYEBG6XqypiNYJl4h0okN9faBlvTCOF1yhgkpCunjt
6zl/41D/NT7wjoadOKpKV1dHs+2Vx8Q4Y6+MyXS5aot4ZORUFyoDLysAF4FgNdQU51Q/TdiJkdqp
QPqonQKHul/5G6DGehr2kmX8ck25i5RqBHkZvZnPD1tPFWlqpPEeGjYxtYx+wiCs844C504QXNLt
+yTOTxxGMXgNtEK8PYbttX61mhhjzyP0idKJjMbOMg7hMPmbKMj8ya/lbgz4x4n1cCBgZbJ/Vnww
CNy90Qo1YxdpDiiOefR4tQOg++9iRw0IzaU6rIdcGG7gqR94KeVgvapYtYvBXngCk0wQqOD1lvMo
L/tKLCZ2owRCWZczJwZN7q/nA99IgdmY8CYfB72wov/zDN93HDAjlQwmSL51LuuWQvfxNySLaKbb
6xsNM93J/gLME+47ufLveku+0jNRhGbvssm9CytLIpcscd0oQ/tvKPbLsT7/vmN5KhfVEk+V1Hyj
f+StMFo3tCE3G9AL2XsZ/sXrQdwgNpxRqBw/z0cbZCYCe5ZICk5tN8EHkyIxZutbZUbND5ZoIIfO
o0y3YQ7m4tsCofNpXUt1NZoCNIg55CuSRLfP2Q06HA0A/1QghvoHlHPL9oaWQ6+FY0sdpo7OaZQR
WFD2MxCeumAUr3zCBrh62yUCZCT/9VB4yFUSJ56hgvf4Y4KqI2tMdZDyKiM3WDiF3cUojLcbUDWe
Mir8RFevQdLh/U9k0buIuHcjn1mhBzXWHANpYkx4VB3j1EdhsaItDA2N3UkclCX3utpxmqVztH20
/srY78yIFQ7jSm5rl6RJ3+J8R3vo1Gmo/Dy0CoJc/sKIPIwci71XkJKzvUZoQzfJJnDeXMp99xLM
7kxbwIZebp9nP/yx/Py+U1Cfl+3ZHn/yZh3bfHOpfCfirjREdDbimDYxlR1XGxnsNQs+A7Jcpg5n
V9t+9hIfzlKx6fO9txQ1ooxh/GA9P/cQdKcr+PZuE+HpnHUwF0msghOj+I16HU5YvXZ7PV1YQhb4
rHJQIaW5poa1FLUdFvLOtNWwqKGbnB6RESDhXSdMu2pE6wPI6fGnAIxW8EUpXIeuMphy1Iiedn0i
7w5rB45mjc6IqBxUaJYUBcVVZvorK7EGtUtyGWo7urGj2BzG4HgBuNu58O3mIAsKwRyKgqXDbnt5
akMPWWyUo1brkAGapvTZwk1plxVPpa28BgXypp24g1j+vdquMtb/4J8vDp6nehvu5BRDY/Oicpws
Z3kIXh0wjlsnjvnsiJ2VVfjmK4F6lbmhaT4ckKj+oy5eHVqYgarLwWdt/919jpe3HnU50f1Yu34B
pmicVUwrChVL8ajmkzbYC68CbW4PVtJyx5w7gB1uI/hqA2/I2NfYPrAPbTsCU8ZQ0G8u6ACzuz6P
bdq0uX/L/dcUjpbWCPyuzEpZqOY1frQz4P6t967xLrQXdVMETXqU4gEbGH9Sd3vkSeOLu4M047n0
/IokbFV8YvO0r+DWCzw45zTuWiIj6jtu9Y0WyFCTKrjUAAZwqkVGCNsXYx1ZCg7Tju3dOJRVvoUY
yJspZbxTrp2yOdjyVPHhNnaHsAQkcCgG0JPwDptAEvC87yol0TdMK10Hxb+5NhtjEF34U//JFA8x
EyvFUachrfL0Sn7dlmjfX8euGKnkWJrT4mB4SbOaPqgpBJnfZLYGhe7QhHMRWwaz9oBasjUtPoKv
lSI1GGlh7SOI0SmFpJe3TUfhTV6CvpRYqjB3mo2PE5+H9I5TbGcoRTtGKJDxb4/MUiYsUyLB2Vml
2Nr6k/kTzfFIp9AWPs5Th9GAndd0mnBqJP/9BtzwJbq+Kh3QEumnHn2t1HzFxq4elLToyQ1Gb5zJ
viNUZSJMIspnPE+Fdm1axKXMCOLoXeCGBbpnwMfSdTY0bdNnEuvLzUzxAdXAOcSfzlhfwFlzyCuJ
2Aknf4D1lQjTMtL2vjwy4xy7SnV2nxp2cmY4rzEllP5nt863pgtbtzLTVxwlLXcW+0FsCbgRmPI4
m6o1qK4YEP8EmB6DdcO9miKa0knYJnpu4HIMjSs1ADBZEbhKlam1+m0AjY7wE50S8n3d9AJHzF33
rrF3ErVrxJcO62AtaU0xaxDJzCp0HaEAqzmNCPBfShCiSvVX2JUFQFRnk2IQBC3nulM4nl28mGQx
/5NT4ObRvYfBjkw08JY6ZrAyv6sQTwd4u4OsoEakbhLVlrN0QVVjF72Go/Yl+KZw855IZZlCixv8
N0C754S7jtgwnUfERmTWjvT8uqUKCcpeDTO5auAo3EwCpmlS7qQlpCbdphwlzSMpzroo5pg+l7yx
83DJJbeWOg79PjeRwDmKg/2zdK0TnVw0CbBYxn//L1F++V4UHZ35CMbp6Du/r5hcNMtMdPDwWgfi
IO5st6UL8Vrq76ugHlwX0pdqRUk4SMxVP6+UYY4dXQkGjbkKJ+qC4JaXWTLvUtAY8zaVtXwdKhdR
Vq/ubdsyC1ZAfyFJngkPa0Bug0V4sLDzfhCDCbCDl6hlAYgFDmfIR7PCJzK2PrrYLOwFMXGSI9OB
Y9YaOia2uL5JOSqilIu5TNnYkAxyT5TO1mlvH7DvJiOaudOeJxJbHIkGZRnjxo6YDj97gN20zj7y
0nzgUK8uWhmKdptKnr9pVK5997vEPXOZvyFHkr9vlRdMwingDVem7kaJg92Vwo0R0V44iy5dTsEL
ErYo4eQapTQeOYa4lkUbgdxuZv4DWUwSx1VYvu8Y47yCVSgFdDnRC8huLOYu73reBTzpKeIHZsos
8zSc1x9X+r0EVNrGkA3AI4SHKxz6CANiK8u2NKeu8JVV/qpXV77+/kUwoF0sTcdsYLEcEt2xTDGL
uZnNK6NJPvBl6o7H5xeY6+UA7LffSCov/qK5VrB9pd3M28hqbVtV4Ybejza4Xg6JFHVpBxzConeb
zP3flRaTgVVPFNvxqppqlfSeXWWQ7NKUoy7KJAxu/rj2WifPyAs/3lkrfXQgB8lpKnT88EnnuLDw
vfiki5iyh6bux6qCMP4V9/ssevqrE/3V3ObWfPV+0VE0tHIoj+tI3oBQIX9mB+4Yp0OFIYezDUvB
SoqQ+Q4oKaNEuB+OsJ99yQ4aqibDDeOnlGDAkQQflGp1OO9EKxq9w9w6BXgHwBI0VPbfVI1pNx01
Tciq3RVjO0x+czsPl0Y9S09ivqYoLmTkIEJJruuaUKYstiJjGtgTuKIfhk3SeSo2oEgU7/FuKJyn
MRRomHU2w+voURSlcPstsjayMBkuOwr6Qz49J1cm+ZfoOdoMCs7Q8YmdAdh2eMKcvlrwHNiyyzvD
I2QgdkneLJI4HllW7bUbqtxrhDh6a3k21btbQBqSNKA7cVYXO8s4lSGeCTTiWaRB7GRgdUQcPql3
ioz5gcUGGC8RRLHKhp341ihe4dn0r+twroecdVil6NwwiqZPkl9vL0BvZVzlHUbypw+63VKDRkph
lCHSmFXHsc/CoC3VYQ3p3QSeSEWlqrp0xaTOWK+JXCGwCnEiqsg83WcFXrAAe+M+H1x0cc/DXY2g
TQ2YP8HFNDcYEbxRKHJBMY3lEFKm2k9JAj8gXLkGBYnsF9evCcrqeFmGx95QbRv09dIOe5+I6hkL
9OWbLp1cMn6UNMXFiRVPqEpKDmdfJ+n4tXHfd0ogpb1RCmQkXOeXaJicKO2Wx6JXtv2C/LQ3LcLI
Z98p4oo1rqbPk2bdtz5M38wo6YsKPAujf8WjXH5Tm899X+mwp/aPMfod6mjOo0CxcwuxlBJ8vqpp
fd0kZbWpjZNHT4Gg/g57MxJIepxhNHczaBCf6DoSLCRqW3CwVINpnzwh/QkSAgut2R/7EdhGxo1r
obXUWE9mnK2PiqB2iT8Q+8oebcb7VpL6lwXo3izKXIH2hheWCGhJK8XGYZk8yhMpYeVljQ7nhFaQ
jI8hP9RAmjAXinuF6PMCrk0EYxgjFUElGW1PBOk05Jsr+K92/NtnybyWkKpm/Xi811WTZStU0Kyp
XyhoMkWmWinQwRJnD6b5s9+AgGC15svs+IHXfbxoZQ+ZRePqjZGLoDSLP9xOaSRwRH6ta3idPp6U
JTEFubKL/3kg+BgUYLyFjigm9oYa6UWqQUYw8RAhmEXvjohBZ5chdz14tUV9W7SoSdaJyeBJ+HYC
1VtX/l+6rAeDRPvbtVOGZyz/fBauigwF2pbhwEHkYZq/+kTZSFDlSRn2sQUc2MgkZuxB7qaXR0FJ
/ci3+Hz8Offs6SDuoYMDqsl0ShnbO25ZZKZbDhnjTrR0BREoIdVZ5Bk9vPhiZOpCBHmXgXnhwS6l
7iCXngKCKPyoGX7iiWMWdN7yENRf/Ln6k1UjLBk9xmPJPjB54WsOzt5IYJJGAiLF3iFsbR2OVSHR
G+G4Mvdzz6fsKdwkegqUNtbG9qoEVKWj4zZJU5vrmaUNRahNBWli0ZHti1wPDE47aQD88hYBCmKR
DXTmL+EgXKm0mrLTWaUOG+J9/nOaUsg1erP8erJTqpULBs4y4a/vPFla1kIxc5czbeKv0I/40Z21
bCJpVEOO7B8+/x5mltxZ8d+EGFjls5nQoK63fVdrtPTT8BFCmknRnzjSUqCpGHrelFIUroi4PqNW
vi0YsUo5QM3YZg33ChPAJSQnzL+sm9AxSK6MYFJj7iDiEyxO5zf8YFEATVbZHxsOhIna88qC9Rn+
1RbqKMNlNOuFMhjADsYjpX6XpiOsYXHl9iYgTGZ8BBgJW0vCQfBncM9UhwG3bpUrAk76g2ozhPKW
OqYaVLvOqrXbmcTXDMi5v/V4DVICn7OGL+4GvTKwfDst7UOkrhmtbxrVJfaMQAEILOaFsO/mXafd
zOnZihixWB0TiVITlbdMkszAVgqWm789DxxEAqeJApLJzCZYllfGnfdUQyn9KghqaApgfTlyQ6Oj
rf7iYL04X1KupAdhUpiMabsTTE2vJemB50F28UD6BllzewiVyy145scOLpEQ+MFFi5/TCj1bM4f8
y+PMqUkoYy+0oU9I6gNF0dP5SqkskEhger3fCf7/olnjXo7d2T4n7miUDotUk99VXW72R3o0qZ5o
ahCQ+IzzJbKgrVTowocYnBOnFShurUMHLK57lw+bXPAaHqxE5oRdRd7Nu7z0E5NWePh7hD9UbJXq
3CVr9c46a7dVpD8YZ+1MBneRi1nfYx1rlhsvmCZ3r0xmTeaLsNXU3AAR7ABmKBwPuTZWg28bdueT
wWkl1d52Qqc+dbCiGqnpJXw6hY/gwFdtnjiKMk6WvM7GbMPas024IdKSLU/c/donsJFOGxtJg+UM
HPtwB9jyL+PuXiSZIuyf2OQNizqiwrhpGosjgEn5XcPu/adnam4Wwht7IOwGYvwKlGPXXWXZamvJ
aAj9cmUYc4kSQJ7bmE7BmQMVgcg9NS4gNh24YB3t3I4Kjxv0k8YvbSje8QrCerQTECP6KsN+R6Ye
N+hb+N1AXJQl8tcvoPBmCjfQX+fZnyq4hsH6OW6D4FC4i4qap4n85GzTo8K6/DMYvW1xqkxkn+wu
zC/Q8/OCGPmBoAb/S6JadAse2Eef2ZVYh3rrl5LTIEB4iPw0E25YkccJgHecOPnwXCwPro5ObsFO
an2vEj9Fdz0MCuy3odF4p+e6877+r000/6yRGfU9RAqFFP0R9+nHofnCv2v31yo399YDBIe2ZE7h
QLLtPEOgTRHYSML8L86L0MD7XBkwVwycVphG7Jvy7SCOA3O7tMdP6HRC7lKmXdLQKViNy/7fI1Hu
XHGc33+b2/KqcFjxhFGObHqN0C6iiFwOTs/XTiYEAVs7FaTD0TAkB5aGy0fPNIZ6QuK9kcDvadLU
qZnE11AZg97PCtqmiIMhDxC8KwZM+efcLcwmu+pLyJ2BhlWb5d1MQweW6av7Oe7yov4IAFMHSijf
YRmSXGtvkYF+2cwSp/kLc0PrAon6UAl9vmLlLYw+WIX0JMxXeaR2iZKkbIQr+h8rEuc7XVnggANY
3ml4RJC17hE4/OTGl+ozt5ZANCTqdkIdoRh36MZQhB9IedifIWYRu+UnjinPe3gAz1c8WhoWANTm
txl7cHRaByfrli5TUa4/tCXfcbnmt1LAjZ2RQZPSOC5kXLcZqEt+8Y9xX9BespCIKLyP8CeBB8SW
R7tlA5Lf8ZTHx3OqSuPSkzMfvu7pqLOaLduyeqdb0y9nNTDMBpu1uPZrIf0K2DbGrKzmsJwP9mUx
IncAweaQC7RxrUXT7UQFdosPgercbqeoB1GPtallO4gpPY6iNRWa7XsiU/Z2GDUBWqzPAgpoYjTJ
6TaFwxHxyiT3LOVQDrp47J1Ts547k0KqmzQmJ2JM90swGucZSor6Dz7Q2kaJy9pO+g6FgLWzkUOa
+TZQOmyqjujZOmf5nh7OPv4m8awGEJY5qEO2tVMbQE0Veub8AzrNd/H72q/6DNs3J8zjol3hX6mI
/VMwuED4DM19J7skTq40OTJLnlgxGggQvJL3dT1Hn8s1pkkLvkOpO0wktvd79Uu5gwxVc5js98Xr
BGx1CGTZk4Z7cn5YVcu2dcK0YXy5ykbhclXN1lddWeCFa2o+HgJnmQ46t9Y9zTbC+53E28mYJ+NT
i2EoK3qGdQuJhnlsQaIyqkj/RYMsCkvKIoQ3yUlxSZuOyHcCdY+Dy+9O9H6QOc7Jt2yJgIXH86rX
RDhAVNgqNX1jndSPlYpkFwiF6ZywfFHsJqunUpZt/NltOzVdbjNLdnnr/mBkFcm3I2px+glOg/hG
y0VWSZOr+7OU9hRZuONzr5k6s+Y6YjeOcfN48jRq86rDLCyT/+IH/x3rQaSvCFhEgzwfCziZmrbY
BOJylbNMNnhAjngrDrBw52rRUUmxRqD7UZNHRqymudK9xFI8kS3F29kTKPfDahm43mtebLDpUD/2
dRr+wLiClfkevNo81dJTCmsIHZ2jWOqDvGFIC6CQri/SQqFx/XFtz3YKxTCIdRs/OVaKivQDW/ct
ZS0QbQPuAUA8eRlF1KOHYWAz7Do72heXoiOjXlBFCw4uxi22MnfxWivk7k7an16SHuYcZnwbnKiK
4qlG0Moq3ZaQmMSGjtlrS1Idr/oP9Nk14G+QPGbF2sQTy+1o0yUqjJ8BpleMjDslsn998XyjQb2e
qrHk37c/nzqh5Kl0kXikpIfkoC6A+yxqyYBHEfMw5TL8oGMVpwczfFHKU4A4KVZE36/8FTysaE0Z
2EN3K99ghzAq8M/an0J7wQgM5jpuJ9l+KMQMQ28iQfHlbUhjEF8I1N1LhZUlTEJhy70Q+rhrKwyN
vyH4w2RZPGYT6ytgt5TvdbxH2ERLwg4TaH/FuVwZVNpQqeZzlGHs+GGXjgM9ItFrvutiQsuxcdcb
u5MeZ6JoGalRlJb+EyxkRAWifpG8dV5BP7wsL6ivJ5HmF+uMXhG6BihnEynMAqkvqm8urNZBkOct
GFescmyNZwhDU0cLN6sESzmQkodKOli7VDTQFyLmQuwk+SrZBfxmWMOXnJmEE8O2dJEseg66xmLm
lRAjv/Z9CD5P4JQxLedlyR9Tc3Gz65p7I45pio3+vgVA/MA+Y/PKD8i1/jgzgq6m4/bi2gH7Zzfo
eF4/s8EHHui28itz1Dm7opVbpDwb9w7jVtQB4gLwRul2Q0YDmQOcEP1y6iq5rVbOFLLIbgi1fKIg
FCBl1ndAoD4YvSdddoQsy/BLSzWEeTa9cE4aai6h5OalJbsj7Nf9b5jKHiah8EUx7HeoPmsOXFNF
vt/KlKTxy6tL/GJ8XahvLxmKWX75n+Wict3O0Y0sD9lk7onl/7OSEHH92JDRTAp5w2zoopj5T3+e
vO37kvOWnis43Y67ZCfTc2kcKXw4sLRMLbW4klUjRaruuvXlUdh773zfxNmWR/JOLtQ8ivwXbAbZ
7prHleFwO6PbnuKTR6BTC1msQpd7fXbBmkO/h6uLCvwlkq+wk0NPNyJhpAUK1C8aEF1WREnafVkW
6sTK1Oy9QGjHR+VJx8LieBZvvw2ydwAolLTIskR6H7KHOHZK1AA1B+yJivMQgU64q7FXRO2OfJIk
jq0QkDVlpWfqGgk4XMyKd++hFUuYS5Q611T5KFv0YvJBO35ALsLb4RQ3PUDQnNvlaCD5244FLM1o
Goc9fxB2RgdXKal6PqYhA2dtwmZIl/SAPB9bU8v5yk0nq9+KikXNbEbV8nAgBs2znTkSk6GvpU7w
Jg7AoGK3i9/mW6/eT/2zaw07eMj+PSeQ3Su3box7CcztCe8eYij+MHmvHJzrOAROJrjuhlQml5G1
9h8h7L/5U8SaT9qPQM0zvGdzs3zBQsI9/GvTk2v537xHkpaWpe4FCa+QA0STIPqdhRdmiCJuytEH
9u3GYT01gG3uKwAeZdqPfyX+bDpGMc+1vzbUltky/cYnaP72Hpvw7KB+n0eO5SH/qSxLaTbbKqc8
yVKVOGrPhejEVCc2IHJHMRPKes362Aex4t/r5an8WIpf0Bl2GMJI7P6CJ0FlrsHBT2ybTy6g/eCK
8sdNip9aMFhNnEj8yMgh0tXbCXQReSSO3AhuQiZZb7j6nr8lhYPMhpaH7d5IgrXQEPMvhj+t3WdU
DrkZmwTzNJHQ1MD6lr6wJ+3QFg3tob8pveDKXawgkgWIxuP6CsScIU7gVNcjAB4LTanYcrmZRmlv
x1+QoyVWJA29BrwIXojvjYDvcLcJb+xdWbK3P5Ee8sDwrBJUjgjPAAjf3YhRM+PpEvyNY6tkQfkN
X+I2kZZmpAtkkbR0Zc1o6z818JA3zmpLZVDBsLx1Og9WTDTRVfn76O/if9g1wbcDnQJG5am01fRJ
a8Jt0zQ4azTLuccW1OWbQB3fMlAKT4GZA8kV0/RYDlJZhmcBaJzqnwG4u5th+FnTuEz9H/cma6Nh
ADkmg+dH+MkEod/9jDpKATEY1/KmmvaeGwpAN5yEa+tOjetlT/Mk9qh3M6CcGzAITYnfuku7bpBc
i4OEGsXp//V7SlZbQyJ8DdNuU3LFiBovRR7K5JlYJjD3Z64yM2F0McD3d6aeGFNOAyX8klxpsh8q
t9X6yGLoK0kQzeIUraJaRapcP2WdchT6/jJrzCHH7NQoNhe30YhQ25YFSKreRBpe+Bg2e+4sJyHr
zBSZNhszujuthKft9+QQQf/OFNt9q3Iky8MLoQfPqhwRu8rmYInqJpdyiPW/XaVjkt6BK1RPNKq2
ufHWlzTZ/K4Gtpst+AdFnZWnV8xUGGPGHk1B3x/EXS1j+beXq44cjH7BLQskKXeBh3g1f1OmrUBL
JEhE2Wp2X+/4tw3CwLP6LdqeU37GIwKU/+1lKV8AZItrRh8gjTqNrMCVi2c97ZkuCddl9RQ9TcMv
SI5Ktwj9QxXc36M7pfE1Ox68CR7JrM4oVL4BCe/z4UHr0t9Hk3psXCQCHFnxVz/JBA4KEocEe8e6
ABPM9bMNnxXzxXxxk3sFDiSp9Jzx6jf959iuNcO6nJy/bV5cqtiM5PPAZY+acHkoSVYuIjP3ho+I
dk6ogq0HeKPQyQ0kzB91EOugS5r4N/ZUm+Ze44cE7cf/TA5INABFbrkQ+03b1ZqEMA5LnyYVXJMC
3CcQK+7K6m3X5lFBoHymfu+5TyGFkibxtr8DmW2zMckZYNAwZ5lLxdPO4lDvatzHQwBeiL0w+nf3
+sS9+mCd/HByNIAaDcBh7AyVXUArjq85R+iAft7B0yG3ICWo2ReQYSizK4tcNf/KV3MSg5cFZBtr
+f9ZgtX+a0zS6ifWTVVZ0YB4NnXOH12Tn5dtC7Fcbe9sbVLfMs5Gxg6psj6VUC0Jm8Fo1or7cCzQ
vE27qRI5w/gh+AYVFd8+VFAsXHzen3IkaqTypOPb5UQVmiLc/h/cNCDEM0i7n+J/QkHpaPF1styT
dyBrYEWCJ5Jfq9Dh4YAai7vSIJl0L6fuab7EqG7STsg6C4nn3KGSaNhgHJMKpUj3PvPZ0Sum3JPI
HzPdXhiqo2vNTkjYHTCv5SQ8ChPeK/kJM1HnQw3XvHWBAoeuATDhWCgDZqychsmGJHIyFQKH6dw4
BwWAyhEqb9K8raSJcap7S5AwtoP9imVLlloKLmdLW6xa3ouo90/UXk96XGJj0/SjZeWm3kAXU4z4
TPrJ/SyFuO9U6McgWnrCY6Lx5n9lfKfueC+PB0gb3VUwNPKiY8g91ryLCmbpqLHFdUkvy7nPOdVt
r558NhX08wByNBUT4is/VCjmBpp4IhzedIJjF5zr/ccnY4RfU3OP7OddEAzf/qWbiGVt3p7NgJFl
Rs0huObYzJIHwsRjuZZbM9/NzyH+EA88Nhx1q4KxJSTxaMSYY+mLXwNOTgRZHDzxBU24A10qWBlY
6yMtU7U4DC2ZOkU2KZBmc+gkXXLUHAwsDH0DMY2mDUi/iJIU2ez5XA0NcqgUhLT7LwHj6ltbD8BN
nGqRrJJWHokiOthglSAVUFh7hERtb77ZkhL0pBnUN2nbfuwfqCCCLg7TG8PuXCQjfexnZrO4Gwou
kjHL49zjF0pmz/EF7Bdhxr3IsYUUJQrskWgaMcIKvdhkrIfjHcXaL/2pHqTgTjmDH4wofMtEwa9k
DQhI6DZYag4zJybfaMmjQuJCkckj2GOMk/WqRd2stn/EERRCpQKeNNAhZtY5oyL0KWlF51wEEu04
8PHX9d/FWyiGlZDoJSMk9/BYWz4/ZZ0EJNocg65LecDup3o/7rp6UjIGwdcOkEyj1hi6ZC5tR2yB
9WAs92rNBnJZXbQmSEMIe6hpwfaqzJP30lGGd+oBm7OZrvyQxARi9SOiZnOueRdRnqy/mNED1b9h
9OSyXE9Li9U/awzz+q+3p3k/V0HqVPY/QI8XhynvnvqLYYjDgDFG+2M0YJIKHGc2rUA1lG8dbv33
R03BA/pWelKo0Dwvjl92F4mq6VrK+4BND8gtJ1709d27DsCMk+4EGEFPEj78JgFtGap6U8B49k0x
GZRXfbmR2k/jKyQnBYYrDRY5H5vPEhjqh2+YA2k5IkKQjnwGFwaWSxV80SQnMy1YFYGb/ivMKtrF
Hnbk5G7lC0K6kH8mMQbxuuxh1g5sxR0BigOwr7Y6pLz+PRKVUQ5ti5csWyLk2TyQGt0efFCZbERJ
61cDHcgo0AfULhetSAhmZ/Jm9B71EEYdsiCXim0r94uyRk5KVj+RQrS3U4i3G1+heLMfZ6EL3tLX
kVGEfa1zaud8ouVEi0VmxnjhygAbE23IgRxHOnHkygmkrqHYfm14ZF0kg4zy7oKxmzkojTAUHW7V
j+Z+m5UFfC0ruPtTKlPgtFp/7hMb9pY/JpEOJ9OEDzUhiZ6R+/zV/lM/hmCF17rouISroq6y4SFm
cdjWwi2wZabCADOt8mtog/l6wByI3Rnos0agd4oLDdKhUND0Tp+exVMGPoQXej2Ra/lG/qBApnaN
xE6ev7bAn7d65jlLyWB5HOFJMWHk9INxnk8O+gxcsWdpYByPW07DRmCg5SJGezPptw3fkLszjLag
DO/9+ulVsLqO+UwR+rq8omP0lF9tA026hv9mIbla+vEbQ4ws/8upT7sIWyGIwwrOO1L7DX94c2ix
cl0MZGdLpWP4MhHGbQPdr8n/dwbeIswLGo0AjeQTxUYnuFEqgBPjCc4XuKQ+yvADfVPRPSeMRkmX
YRpuCVhzsitKFalzuS6K4DU3CzUSWpl7m7zBRxEgh8cUtXUM/ZknqFD/BHVOjbAKXWUHu7R6tS81
2k4OirjndsLEzrJ3hVFoslQUmaMhheb6FpCq2LL28darbkF4JQyWdv5kTEtKS4X+naqor8yzOPFW
MjnwAoFFYHyeH1FEp8E7yPD5mOXThh1POhNpof7fUMhfbiKu3i//YwgEkQSizSBkvgrENJ1AKA5s
MGVJymUdr/Ofe05atunkJhcAugMaBkb6xYb/kVyp+dL48IcSmYvyG0RCgBDGq0qt2SQmNQm3NdJp
6yHwdAD35Pw+Jg/OSA3oWTald3GEcdt0XUdLjejfNQc/0ce3vH8hBmJ9FDnQ3QI6ToFloGmbNuwQ
tQlwhil6MTWuIH3gt8sKj0dulS3IXT1OqKA7xP8ktdtVLvQzm0r9OK0UH9wbKEnkHnxX5Jm9Slwg
5BAA7v/MIDUsZJXPD3QOnm+fvnuGf7FaAs/UwP3kN9KajIra+SeSN6sTsS5fDXgKcQ2SRixfSv1k
rQsCgWEytcTk+oKLeZREQjNSkPbvBhnKcU0n/YEmSNqWNtssrJxIueXPgRO1IpHn+5ATWSojIZCn
6XObGf22Z7OahSH1OsU9bpfmSseSOHL3YkkU4zyA63wUysW/eFknAPlwbYbi1Jxlsnh5GyO3sZd/
yezOMQMbQp7nsZJ+uV8Ac9Sjen3Rq84EvXzMG0mV9kQEcPpiZGOP1NfH4MtzPNE4ouRYPF/D7srG
I8ZtbORw/LBbDWeDys8D+t9GN6gbhms/WA/GQYvAT9huMUbA6PCUgQ/L13OT08czkJMGz/g/rQnG
OMPcSp1MOYFeb++hcxXN4vyNYeJYQIrJGZe+0N/YDiIpsBF69aapeKFWQLN7yUW/A+b6UKdWiZ5x
ZgFW81pHY1GZ3tju2Q91uLLt36hJU6bq/Htl8kSxG8f5tc811ojj40b0GF+k3zzlYcYuUqcATPmN
1wYfqBzDGzgTwRumSa6g7w67ZgbCe048uidQMPvBlkD3dOqVtBo3UETVenr1Zdv5OleDHHY3aZKN
ffyJiG8u0T+VEz6MA20NZZ6vVSkPT5zugO77uhm0qXYt8eqzbFRvVt2Mn4AZExnvgA0Wlgo7alxt
abTBsLUHGsxq2j4Xc92Fe3pRFrj5DUXeWRKEI6LYdc9JP4jPWkymwsHEr0FAgjDy2PSTq/L0SHJz
TngdoD9spuQyOVGOdUa7zyC8/UiPtk6Ud2mT/qYuR1JgTi7gPOSMIMOIg+gxTeh7rfraGQteKea4
Uzvxv0Fw/ID8O3d0XnlxyCLvnBOUX8u4cv6JwP+3M0fdrRg+RJ1MbPOM4HVGH9VZVQSwxy0Qzhk8
zROo8SNeOcnHQAvk6687+pOXpEMsNE4IQp1RKP8oi8cWr5aWF5UmFLPfR6jNXTHPQvCOmZ3I6TX8
CO/uVwn6/cLpWZvcdp4LeWW3BN0W0115a2r1zFTe1ddXAC+LAlzpMTv3qNcwwJ1BG98L4KN+jFuk
/ubvNveoBnjUGab6m0G2cZtY42lvRUwl4unKQrWypBJ+qOtd7QN6l5ejjjheydVXAqEEUZ7gBkXs
bySZLf9Iedt0HJQT9RNPAOSdYBcsiaZWVFmV1vajJGV6txnly+xbz91b55gOGypLENnztc0SG0X2
J8jz/P9sz6ixmN3cGLA1IDG/r+ylhSLcVzabCheL1FFAy+V8VA0oUQSwinl3IFfKgHkFhGta0r13
M/KGDxd6OOhhCKPkrjp0kvjW60bhEtN0u2YCBZtSncGHJfMyFWI49OSTLadFQUff0DoksGXEjdn8
IayZVyFNwL3BgNBWjiY8i6PMAkAuiAIj7Wp742A6qicl50VoQJpLltUCSTWOq0CDzbwIttSAUglJ
dFWeWvBs3GEHEj8JY2nDWrVrhc+UWe82ZOsok1x8TIxOo2/0CbpTAwjn95fTDaCR0nRLQVP7fpd8
hpIHGnSYGwvFdTbV7wh12z7eFqojTthxnob04i/72yVkqxvszvIWzc8xVEmpcGVu33t3356Rk4t8
sC/SE/HeKKQDZv62hfZbhe9MTbzDkLbKEf+Z0pvfQn4dJtstkz99Mt2dynnFJo4PwjTXQ6XBG3Ro
j7YovI9aVpsAVxO6uV7vKzV4x6lnF7F5ZxlUclc1SsNvvlfLUgYw77JWMccIrEaqL4dsBbinsKI6
N0HlhEkT3YCpAoGljGL1IPm0C/XrDK4Ie99lw1S8XTVj/TWVWosT7ua50R+hkA7Qbx+yJXqCTCDu
ThTkKYAo5sO5ZwZkDERMm70p3+XHchZKHVSCd83bcFETEksMVfdR17s2ByvZ8Z+GlsImKzs0tBlU
oVLmQ0iXfk5F3LQUKRyZNBfvlDWTKAoCpKEgsLd7KLkhnadmOBJUvkpcl177IqThtcFM8rT+UQmj
bIGGOb59YYs0iaapJo3QAfFz8bPDs14pAKLYSqm8oa6WLivQ95IvHSNRu5OcZcixjkdul90N+tUE
JNeEDXBtsrDBf5V1RSCtjEhcKBQKyIWCZhF860Yejnd0l4UXehR5gkRLXj3usJ09Rvc4S+3BVlYF
Y4Xzq+iAQJd6A2u8uvzipEPewaYrkSY+izHeZ2KrxRhaz8VvsEfiJMyZJt5X0lWoTJ8AajCtIYyc
PFkZS+Ykcia2xgfpykn5zwWeWMmlmGIPDiuznaLgVB1yLen9VIB5ShtLBiDEDCHS50cybwgGiBeu
f7t97XssdBheBPxxaNSDYJdQbROfbtzeLh9iYdBJZOEI35Kh1X7IR3GyEZU0YMGZYBV63unrbPnR
zgrqQPOk2ITRakFfAmUFu17eKPu8lD05zyWXbNTJ59uFQuxtlAZod/R4L60+WNGKYd4IGOlyPveo
8Fc7dP6xr4pmlRYMo65mg92RBF5DYl+E3lFV9HC6KCWTJ6ihPxxo0bxbs+F6A9UUJz2PEsfin0Oi
h8OYhLFE/SXV1loDPLh20J/aPU7fD9RffJ9dByghkEYZQuMk6Xab2qhPVfJcwNtYtmD3TqN08xIU
NPki24dQ5UVmGSJroFIlHjnv5K8GtcGCu1jT/MjrvXhNbgbE233wFV+5Mt3/ty+6sQEnFRSQX21M
iac+VlJ4rBKzIUmAtazK3oCVmo1os/jQ+3zymzEKfQKZ/2VeXRnLyGUsfeLNob8MmSjnOCUzsBNo
l93xlD3ExPCm1XTk/OSQbcYQp47eE9iY7BzC9tm2VHScuZ1k2pCiOyTD9CJZknAZIDaNs+jHhsb4
aCYg0rk4kKIe5hEBlkuJUjubDQjj5uojbDraEHdXnKwPqIGadAZ1vGFynsOWn/XWmH1/ryJDFwse
AUBg2RhPx5L0+4cXA4Dqnq9pgi+lxygacq2PDTKZ7ZQ9pnoZFW8m6N0W9+s3juG71g1ZXghivime
PVT3FWnPmbw83Je3azxnt+v2Tucv5uVNx7iE457oHk5SeU1wWej8xpPUzn35w4gY56URVBC7XcMK
QYZVnE9J1zJapSHcyr1AXAQklTx1v1LQ55P02Ne2lHkrGEF+Qlj52XkQKVRRYCifS8XRPlISVi8Q
q5Qn7bt95N0+rU2WWt5Hs9UhmpQoxQV9Y2g4hdCGbj15GgyslJ8+A+oSEIunRo4ICywSgf/k32RA
B84cWgyxzFHfahr6ITbqaXGTPLofo6I+Q5mxjqfSjyVY6KPb6kjbP7IV96KkyWothtsM/I0kZuj6
/6Kv+6KvGHZ/IxCtp0QWkopmWmMgDGZL0C2zhMmcIl90ePe8WqDrNZ/qI+edopy2B3mh8HrDA07J
Y7e2P+/x9NORO8gammpI4jSUKeLAQ7UrTMMQln5NqNe5EU8O7P3qWUQvr3kGuF1TnjqnlLMrE4ON
3CKg5VO1iVO1OpkJGsA5zN7oHuwjfQx4jVZx9ByOG4R8MWKEe/bMpJKxDItJ/j9efu7gK+2fAV8Y
SFX5CIX11MI5X5oqxSeWxYOKL98E3ah833bAqcHXyvkvArKbGkRoW/jL1F2AfSlYxGVqNLK4+qra
dL3S3v4Qdakt7W96yiqak828D7sfqY4G342rjr0c/qfHTKhqjj+cdzGv1H5bJm8SNR91K1fB8LS6
LEAovEjG4mDjkf0s76V7xFrTS30Oi2yOin0g0G53f6V2hp1didja9wlT2fVnKHM065DBR3c9XzIF
ZbvJhPBVj1VRbc8q7FUpnTi5FAK6+DW9h6M6g79/jPfzypNeKBpj+LxI0tvX5cuWKVP2+MdyP3U2
8yTl3kKOm6jiwFD3MUvfHWSRN/mPo7UhLoJlKAttnUkYzkF4Udau9R5N8YgunCbBrQMH6TJJkeZ3
kK7SlhkZEDJpydluz4WXTomcyiaKxNFgImhzJn8ucagQ4nUxXUN9X7Qm5vTMAZdKnfQaf2In2/ty
x1CHShiA9qafhIS331MgWIHmplgM9qAXYcI/XstJhf9E66cKNipTT/OMDS5O9O6cAJ4DZfQTq4Qc
Y+xk81/t+I/SsVUdFdQFydUngt4V8yUvNHPrtNeG0+CuI0/VKfDNsRj1o4sgty5+kvDFPwGSJXGF
hKOj1nxuRxs//j+4LygTd1xH6JD2ffKCd2fr2jlCjPW/npJ+SHcGwmOeLaN6c3MLDMJWytxkufsf
KDl4NCf0y/EmMHsJwWTgm+u/fdJ+ZLHm0FwPxC5Nnn1GJQkv06CGglFCGFli7avb0yv3QbOHAWJo
uXZOLe7V+s7EpnxTI5JvI0YfBI9XmhosJLB4tyhlApCRT3V2FNNZQANmZQImlGd9xD9MnJiglIzf
+97ZYci5H9icSX25QH6Lw7KXWDntLFXWPI3TQqDbN2YL/cWC1q91Q2+tnxoSEQAP0pg124tXMS5h
80otK3yeBeMoajrn7nCOx0R1fwxBcRl8dd4tODgbUJNYd7xKhiTrDOhW+4+9SvySrKv1gbWfW0QA
xNF1Oa538eW4dn1Y73CTZL2PX8/jpAJabskoxXX65Ll1YbBSRry8Aqu7s4ume4INL+pDQaUnUAjX
qMjI3PuY/zUBdKYkkHMbJOvdoveewedSD9VYXYGBiDZTNyjUVFa+wCBuiM0LZi0dyOYZptcQYayu
y0BHsCSv2pl/ywQVAGpwjmQ7BbEpZEnbhFpHldrIZBTE5k/flQjnS80qMvJd4YXJCyfi9IFfgyKO
lgyParRY6fg6CGdkOusiHAJs2zdtUQ6YNrqI4BSDSZHSd1bLhulYBVp1UrvDHwv+Sufj4yCqdTLR
IRIG9JQ0JXBojAL7lQQlDs0IO2JTgzPPA+ZYzIosTDiZOv03380qmoQHMDIl8jMYfc9eK+7HLsqV
Bn4V+DCik/UxMaK/c5Io3VkX6natkz9XpM8V5rUIEn+OBXkswRT+BwiCENIKxsKGy9V38wPDIrFG
ehz5gq1K+cgtvjs8Ht7eC/KtIPWInGE9ES22JTxAK4IqcnDtDHyyvAqUdmEP+FwWJYnC7WxvMPHy
tIHrN3SEGVkfer+EcIHJ6Y++hadji8n5OOPmntCai+EGyR4pXfzCGPDzEMsjPkLhIKifsIuil5YU
mKRIao4gXjMTElm1KKwxHu1ahzPZmQcw1UD1LYGcnv7ViA/byXDZfYwSJiyfDhA8yvnVzUodGSZ4
Cie2jg2TISgmfaDTkXobmVG/VbBaxpPuWnF0fEr+OonYWFGVkdWH4f36CG+InVnEcAAn3sj8SzdW
9VrF1aXzuxVsmjQCZ3m/icv6DJAJlzn886nLwuJ3A0BZK3o5CGW6NyuhkqcerDHayuoDKDhBpRtv
t+sQ+vGDeCzs2d09Eb2gsaXtgN4YPIS/OIF8gR35dnxXss28N8sq9nay1hJaBH1aKyBiCco0xq5A
nDpwRKe0oAeY/NU5cV2Ewl1NEXxcz3T5tYFx2c2uc749JnI4V1JIce54O/OXj7nzKzEx71S/guKg
SbcTpAvp4iieFKi9rIIf6bQelfXrehgXJJMtoBO8xT38Ywi5WxbzXM30ByQgxuvTumgXiMfhfpDU
FRzOLLF+DWd2R0QLk4gFqw2GlUehhmZI2UKn5WqXBP0icxrzkQFIJraxWan2yHDR448wPrB60STs
tdp7dpFCKz/4gLyIW0uz8qJz0wfFI7257qYT0rXOkRs4PXiOLuNAX7BGE5Z/iFSsMZGn7/6WfAGf
fhKhvEYp2Kc7A8uXPcPD1a1t9jRrEshYdCLJVyHQW8L92XkOJS4owmPwobU1Ym9S68uQUQ1oRrrM
DOTFkSTfnd6//lxui2rbDlfmYIBpVT+GE7G2yo/LtyY5pEDKQug/cb4jqaPASUteiOZP7IUG2VLj
Eh6RjP0sR2c+C9//b2cJ7gah0S57wHFnio0t35AMIhamYldM0mopi5xQotok7encbQf9mL4Q/geZ
MndwzFWUbK1lluKhAboJJb63l0PoiLfB0bBVNAH+iSz9r+BStmV9lpSjK/enVgkS/dW6cOblVwVz
z547+tjyVaou7XH+jVnxpNDzWvRPocLn2aRcjx2JbWCw3rNMm7jXCMH7nYNAS31b+NkUBErHGMhc
T8xSVN2vkQMRTuKhw3znj8T9cRvOa45wTPAMhW7x3bAKMOyLEyfieOZCtutj68Hx5LMthnnQrKTm
tXnhI/BDVC5ypD23URRcakvC+a0clxrf9CZXEm4OagfZu1zx8GFOc66nK8VqnkN15b7CmDYq3kS7
e9eRNwCxWMuOrgBRUnqnFXbCGGWzkd5MZPJdRngAzSW6VCgtqusSUCvlzgyVlWwSvti8uC8wcD6v
9onFe3t7ukQfz4yw3oJyNiMXhrpKgauqIT7B0v35H2gvgXFALmf9ubqGkxP/+5je5lwUGk9OhuWq
c2dhjHIS9Fk1t4ryLbWQaDGL/RSpwW5TfVGnYUFR8SrP2L9n1uEaKWP2rCulu7TFxCU0ds30hPEy
uWL5ShWcku4WyOsD1tfwoahezXp5SZjfF46QmsVgKM6Ev4CMgnMXdfDAqei/Mf3lUhrMnb+0D4UA
qcfTGhl4e0i75uhNbwG8I7beZzIYRf0mtmq5xU7zsACXVbizkrB+qB8Zssfcv0uZCrZGCbUBgpWC
xXX7YC3Y0nGar0QdHILkxX/9CqaNBk6VHjt0VfOWZuEwcUOP+2qvtD9uzrNwOzvUfXxhHo3bJGiG
s/t4ldHiThQ8tU6oC7B27WbaTxeeQeQJVaDuz395DRqlmqFJuozF5kOKQeYRxRFIW2jp8yRzCUg+
GjBt4s1HpJot1iwkRqSKbhOrpOyk9skrrSjX/gMU78hjdei60P3Mr/7RxwjbWfRIf4yNHOtpQWkw
ot51vGtzC+K4xG5EXcQXWhqrEPYLe53XEkM41T5i90NIwbZynLQwD2L+R6d2aLni89qCQ8w29AMr
3Rm/GgbxLzcaFKnKWZRz9IrEisAoJz/EjUoJKjeHCEHGA9AMPn8dZj+ZZV4Ws3YPQlxuQXHuQ0RY
C1jdEmZd5+rRF/9bFdeia69B+iusptZKXcKTqjpXqMI2FdWd0BEHnVRSi6hbbxwhkR/FziCz10tf
Hors2V322jnr4LS/IupAGgFl4V80JG8xAicEMl/Xip+PprSIBnqw0p87MeAnPGvV7h+rSUIXUHu/
HuQQwjmhyVsfLm4BF0a1yMT2mjEZ+DxGyJlQ4XS7jNMd0MHBwli3QATPsVhql7hFvTLfwTPFooC1
GYc+if/uqhAiLCCxIUfgUE4uHVP+7liM7vjT3ToMoyzoiwl0OiDJ3nInHWhOLu3No/V85zUBa3M0
R8C/j/ME/Tzb21PMNpg6Xwdj7uCFvbEQ3HNAF8ib1Rc2k0MQsSpTJuQM6XpJZXWoKR3ijuc22Ssy
U/34Yqy/FpfF1hUY8knSmhX1/x/+RIHhhxurVKnuicBBGHhtXJuY9gbdaNrxx6Wp42bmekVKDV1Q
b4t8kcSlZmvwIqRVkx7ZZcVZ03I4x+VNSI7zUkZN/3N0Hkd85+4x5uXwocO1PSu56pgYKfqujB3I
oz3BC2nEmZdgGwdSsPIUyXpIQ86rOGUPTl0kR/GIm1KktHEjDHzY80pWF0hH6UJ/WB65RwWnBdd5
ZFx7zMPECCmHQyB8aZ0VeWN9ePnFUePsC99CvDyhFJueTaySWXaAtpyJQpyPFlxZCfEZeNuEYwLq
/mGMIJBs9+fs6wKiEsWpVq9cR1qRNz2p4r0B9IVg31PscFfqyShapjN/Xx11UryIqiimYb+WgTPz
fzRrhO0NYLRS0BMXtD6ppaM67NgvbqnHG75P/LAhdeMg7d7UShS4IHNsFN/rCxUeE7qQNR5mGYl4
FQUL+EuES2TLLBA+RDF3Q4a2ekBOBaOAXSkSW5E3SU9glOEB080Fm/SKlTPX+IA7J826HdFH2vCq
8fIVCbiFfb16ieTRBQ7uglKZ7Fxxj7jdQUJBFIol+eu4AqhQdfy79ig8+OlBzgY+qxXQUYEPwOWf
GHilwB0YwaMu5tkwyOVBA2rlwLhGrW+NaAjUqJHjfzN1VLGW9+O5aeq5WT7VnmNUyPJQHbuXfbzG
87GHmK9eWXwmp7CknkmveYGFngTjzwq1JqcVkzA1xYG+mnHBKRt3AeEOpDqDFKvX/VO8lone/3K1
bgJI3Rc6vb8HT6b0d4MQ7ky92qzkwk/BwS+XTc0VVVPO28MpY5rZTkN/XUXQowBYfq2nW2+cM2qS
sKOLRlxDUlZ7mYxUazNfgFm2Ph90D/2stuBjHSM5IgQX4o55qVH0oLqZh/lKhtRtOxKjmEQlFtDD
jMCREKfkJDdrBeeKPtONbvLAX0C4NKkVkpX6t+LW76EFSD7Na8/7KHSvDy4wbYAblRw1yLn3P8ZI
NOclkP9GTqWpprqZkbqLBo/6tehC8ymoU01YOpJv85v1tfjSDp/L4/IH6cqnMd36N5BIdad84S2K
e11n3h4FRt44ZFKRTHfUIvvNtCUwZWSDzl781VPTNeNOLYsGZNsaUFE+ogIpGHxnmDufUsl+1xwj
S9+WgwwWSO5Tn9kgQPa3e2df5OcjbaunziFKWukrBil6pyQolDNXCKWjOfFw0m+MClWyekQoKTgN
rEjuqgYxpdPwLO7/3zO8FL49VxcMiWNeNkFpSfbbu1NO//SgBdSqdKgDPRuitRlqFib2X6OyL8Vk
xwCxw6XCNGLUg7P4X5/Qsq6KAvJ7pnJ7ZC8vMjGAdvPs0pezrpBAe7GYxnFYOUvjWuHYWxUYg1V9
dnjA9FYAHvk8J93oET4barxkslC3F1VgRABgTANz7xZZxNFF0o7DGY4Emr04sb53UHFnEA6TRr17
ROL6pis4tZsi0ya8S9XacO6nci/MERrs/q/uTnCAy4M5XviCa8VCf8y3YyriXrWL/NqEUPAxNNoV
UdTp7D7MLE/tnvc892mLEqJi8c/SFbuva7k+iBNh6I1AL3bSE99isXnL0ruKZh65Mx34Pq/so20M
DyX+cUUuXmD9qt+5wzX6ZEoK5hrOB7O/f9DEg0mnVaiW5CTI4TsWu9FlNlOQaVRApo5ry2RXID3C
4ukjYPGni1Ajf0caQrv24ZuGFgvaCaBwa8IN2if2m9/Y63nfRzpP2fWGR9ZNrrhy5ZgDyewGddEw
PL0lazagBogOQ221OdfztPKyY6H6jJI0SRpOSnR1KBVOqxXJOK2NQCafET17DDq5GUTZMfPcYwd3
mv9L6HjvDaedo7kdZZki7/GxpdV/xqSdHgNbr3QOh1vf17+jMnpD/N5DfhtUI9GfHuGkeEV+O1tb
xcNocHbZo/Wcv4WeW3GBGUPUP+pUjTYQ/+7aJzr9qLBc0BgZZU4HL2pkDzLCM1CvwoW5b28IS/nj
qjgoMXZDI+FiUwK12+fsuUQUHdEoXdAfHFZjh1Mi2OAn1zgQEkCCt03AVubCdxdAXki1z6tSEaUZ
DGE4uOXyoRPtSATVf0dmRLQ1zYVpMBLdL+WsrkWI09767R+Vq1CQH8J2AhDrKSA3HvB9EgJLvRdq
f+BkNhjwb4dhQZ2lTggHBt6rmrKuuwF9Ey4zXpNEutks+ANzaNmJXSAvNs5BBbb7Bz+SS3i5BDPt
B7BIbSAQBNw5f8n46vhrcTq+InXsEkMDAnvdrn+EfXRC2cFGwBvxTti/GxYkVLddeaZ9kwE8tMpO
MRYsgjPUjTbsfBRkFE1O6Fr9lLPP+RGx3LzsL5puw5AtCWsqcknGz1ze3FVlu/DgWoaIwcGNzj9z
NMIwN1/gojru3beE3Xs4YSwqIRPT9+KoRR65o4IQL+H2UjzTcvc/jAcvu+BcsV0rRESseZ8qR0D5
CBSJuV+YyAc8RBYToeAIulDNlDHLWgfEh4FKyysWZI7gq6db80O7N7AiGrGW+53oEG4ZhAoayAHr
snggoFUhiEuJIbWpxTrI3hQukgVkJ7t6Q9MZclNAkG1QtCsZXatJUz8BYYupDZiP6lbSOnhQmQsU
SVw2P58ome82V88QUjhDxl2O+IrUrnjFyMAsyRm/lCvONvEM7z6/dNPZX4SYN7BTNUEE0C4sdJee
+BvbAZVxOe244KgCqkuqzwhkcYRiJFMo8WY+F+ZfqMVDdkh155LI+BSyzNxh6OiwO+74gP7h4+ly
e221TojhtJ7XSTHzaqz0iV+HjHLGX8FPAlzTHjafsN3W7qt5XLqROLwIaGAp5YN77MBwl7r0D21z
XzK59Sj1nNTH9rCs9oKBCP5fw9hXtpscoqVpLQzbd9xkSqi+QM6R7BDil17nUrkAY5IoxbYHsR6u
uo2XvK7/mKjWWjpvmmgsbhF+QYvWpPmFtMEVKwXVbOFr6IsF4pnsPEVULEfOGirxuJfi8JB7R6wU
FKeunmlMtwqMc6/H2zRrBEfU1AL2pi/Lzk3Fs/xJKRGDZxkQ/8mVchtX1Q+FPPZOzLuC/Bv/SpkX
XKoIz7359T3ic7kddRC8MiY5NFfAQKwPxm2/KjcsAZGendQnij5MZUd0ozflLg+F5Lh8TeBodSYh
6I8NMy+RUbN+YlAwOoPm9qJNy5E4dxJVShENY3Ld1l0TBbiKugBtIX8G/tTQ0c+fxKguoc/C+Ecn
9CfVFPYKfEf1lyUjGmPrWD+U/BLjkUmxJpOq7faDJ1WnCZoeb+7EcGFx5bbiO7ihf+4mtyji6EfX
jPwRTTErIRk9waCznruDjbmnTqkSIX/AyuO4hQU4MZ7s3He1FxVntEffc+oBYUxcCNk8XtyJDbKt
BBI/pnwx86qo1iiBQCPYCHK7So9WEo3KzZpF6EIjEk/wwvGG5jf7Wsp5MQzZJ9R1rVMgorIgm7ko
MEvdWKDwCAL5hx4fDhGUbNdvfpdEHhG46V0Zeq+fGJtQa9r51J3Yt7CEIXhtxK1wScBh0pNoGwiK
NTp/0g0zr+ZFSx+pQVabHqB85ayebAwSCQW5EFzIB8vu86HmJbIhM3EdSeEGgT2mmeyKmCTmku/A
nTd+5mBlO60bAgWzFqSSm0NY32S18OqL/LV+sozoseNyJRgJTpM8F2x4YSFzSnvlM9UKZkshkPqE
p91Zb53egLzsEu2fvAF9tnTDlww2jdDmH95MW4Gaq3ytHxTwu7Ey//3UvjE85DH7kbK2Ibyq9xZt
f/oDaCf2TPfFH7EbalKN6KBDJ/s5WFtEFko3eMrbqGc8QJQnTLkPIip8z709r0/fOQL3Z/Irn2CG
OYwihyyuHa9aZIjtb24/NeNBEXKWBxheZbTffMMCSebSfSRgvgD+WE0uTtZ5cplwozIPq4zHgPTC
cZ7i2PfVp+4X+w9D2H9zs2jBkY4ZBl7omqGn4hXlaE37xUjSDlj1u4yptzSORid2VrgtnMSdAyay
h0Gxb+3+f1E9WYuLqlzSQWgc65D4i+qAA+0NeYfo56dBb7/aCbYzCoowUrH4GSuYJjgToq14b0Xr
R6SvkYNMU3FavZqP7OjkHJ/vko9JTYsTCcgpvOKx8oIvGZvzrTwnxuU3cm9azTk+xKiBY57sep1S
vgtgfGD7qF097NE5eumfpLrscPBLpdx7bxjs+lhoSwf9gGCbs3A/u/Ax0+jbJDVmKMYuaHWCgCTA
+uqKbV+PCpbsY/ZoaYCnIn39Y6F/M5911WFkTppyS8lv21/FxI3YSTQ5LI3Awrft0zkvSUsPZtBK
CnWDkpIT3kQv6rPjTpfhRXIW8DqFH54+qDCe/ekhzpoOJjR8EVTvV3Cj/1EE71NRfG63jN8Dc6/r
AOG+tdaUObKzGgGMyTL5vOlYYbpFwrvwIbP8EsGbpuapCWIKloIlAgImXm1TDaBOpWUhZlArUreh
UVc6fqhlD3w3W4xvwFCiRAcoVE1uysIBJ5IR7gGgeYcjUEHVxSXK3/LP0EkZ96PeUHAlk8afvgYJ
uufacnnPBpM/jPGkJCYBY4x2G6qKEs6bqAG4mawn+tOZ2UcF1aBEvQGRAunBCG27i8BuuZTF6VYp
NceS1KKuxxOCAFT96GCd3raaUsNDAF0m0X0v9LMWWbzVrGaJgUyI7mQbmJ3VWtVdiR1OeagTlwi6
pmMWBCmDLneaRK7lbqdCBoGcC6vi94mtlgbr+3RshkR9rR62Pz/IJoKlEJQV3uvB66vYkep0NhnT
QLn0OESgQMtWkoE7a+knc8yLDV1nvBso7UpKKbO1kIaYeD2qbP4uuPKL/BliG0NVatjyq7hiQA9Z
uRqkJbQHos0TNqbKzNodheVlbLmK4BfYv+hXXm7fRQ3opW2RIqXU4Pm6Uir/4DxJmR2v1QCjQGcz
UQl1HxTlUonUGIEeShaNsM3IWPhqKE+C3VkYHbpS24L1WmY+ICRRCi8ZKnp5MK51qXpFAqWTG1oZ
6KRNdf6KoDvFGAY5QpaF8KUllGjBFhVncrswXWuaGIGag7/n+Dlofxjx/myRLdRilVrfOuf+NYxo
9I17jvZJf4ZPiQNqeMx4xzbZtuhUsL+09UIP/4y2kE8KQzFGEp2EEXCMOe+CnkSmNvJ/wUgB8DFp
7TAHH7gvk1IC0lv0TctjVxYRBJG8jz/Xr7PQw0bP8IcOcPfsXypFKVyTKD7bso5MOuqOCFqFJ9qJ
gPxQVaKjl+uvq4lkTLaJxdAruA5WoxtmI70Ql/AGFpey4d9pFS6sb4Cs33GFkdCel7uEi8QkdcKK
8fJda6pH9g+q51TzIYXTu6P8xS0om3zGYi597XoGlDBUR6uTBNw8pQulHAXnpnmZkHg6x0airNwJ
eCx/d0iRkU27fTcWrYi4jHMDsm6aVeQuV69L6v5BmXi5bBvTi5mV5cnwwDUqVgLXCxa9C30OZjow
fa5EW6ADSzbnISkw4fWJ21km7fvHfSrHo5dPm8aLigXwhy1cPzkN/40oCLp9Ka49uFtp6IOCd0AZ
kn5o9kyt6bHWT8AcumxMPCQTb/PobOTjhGQ63yYOBrocp89YFhXwIwtSvuN694j10TnXbuMJ7r33
TuyZEihOQ0YE+GS0q/42kj4X6B6gfJqHb3ERmNjvF7rhEVe1DSTTz2KA/xD/xWsvObUH0DmBkWv2
ikLR1MpVRaUPofDwUtr5yMnaEylt+iIUEylulyoD60+WH+qHIqlZI6jo/X1oGqH1ZNHtxEK3K0uf
1NpeTwk/0W+9JbZN7JB0Wu87eaaUlu6W+2JkNqvf4rhuNS6bUQwj8gMk9BzZv51lCZ6CLQM4L8Jw
4tNQVm8oD7+ciRN8z7k5QrqQxLHGwZ29TIWO8V5e1E7lxtbT0t897tq6jMJZMggFm83/bcKWiIk2
A8+hO7X26l7+Szy60RAX+uxUig2wY4W2GAcPyR2Z2ErvI8u+/rKlcH3JDEmT2QfgPSIdzG6SPx79
o69UgJvoyUb2yV64JWu926x9fb62uWviQd9JPfLr1K4G8VTJppiYPBUAwtDYRaZ8+OwPd8zQgDBO
ahhdAao3eHTpN2GWQdGefMfvAlo5ESUnOHqi6XMnbsBxXkV6WOZ2DSRVPZmXCtAuQotws7avaqtN
CK2gPnlw90P4Wr7NwKWG+GcDPMm0phEEknglP/tYjXQhJFo3s3LdyEvXl4MpvjA1C1fYlOv6r+qO
jwKp17HIQoEu7snRNQ2WqL1dyEFu7fQ9YUX7LL0dtR9iH6ICTpk88SX76OAw80SdEHUCbJBrewfI
H7wAey+xSBtD3akzoMhET8Qal5/pR0xtUbrAdmc54CIH9KIulC5Xx84ICt+yjaeKXzxZCB3H83HT
9qh5GSEsSh5BMf1x8B+EfBsJXm88WhJ3ouQJLSl5fr8FGRFoVvqAwe1z5DVT+KfqHwjmGT+p0x5W
dj0pb5kXitdfwvTyn3S8kXUVtCp3Uhjd5XQjSH5SlKGVmL55OElw5m42G3CrKywJipIUOwH4g9fT
rtQ9TzbDodDHeTIjdsLaOQnVblG3cWcwgTv0INDRlMRwvpM9HTHIqTNi5YmuyC2RvVRuLDoEege4
4Xvl+nlpLVHianu21y2fZifJTnBdXY5EBUNCYflh/j6XCV1CRcMpBCS9lT+bJlyXr3SLbBipQ31g
eb0BrXVrkQHDCctur2br4tOekxRezFzsd6BI61bdGuti0KfzL66ps9KoLEAj4/U1IJT3U3nf9/nO
IudHxr4m39B2L0PxAYkc7rpkjBkW9qDwhq1EGxKG7EEMSb+vCPw7kokBBMnUyjbzQZImUx8jrONS
4hVXb5tnHJrgWu0IWq1gO/q3lAkBeRFsMOzPPhuXuXIDI3Yfl9jSbL1r3HFdcotn+gzeqS0UHzd2
AkwN8+lntW9ST/sS1oJewgJVNr6FFv+vG788M0xee3u0BhTAy/xo4eInnAmbDke9LxvrPnPvP2dV
YRMLz0y9pFiK+9eNyKJc0htg8w75Uad1FdpYKAvkhfR+Q6aT5bA8qg6sAHiQKSQwj1QPFkTfMwUA
NAZc4zD1fpwYsxo3MpPv7fOv75Hq7oofIHmxOqkmaEQ4cvBiXufuja7tQp2dH1ZHPY/LG//o6WEY
6xJPNlsWvsroXpb5YfRHllBUFG1BYHrXuAKy6Rev+gj0e6scBJsLUHka7HidVbhtyf4gXWQq8G2f
EIWdGF3joXBCzNhJsL0iEqOisGtDgwcpVn/RUxPScozC+569VbDGaLQVWYK764bHeSoFijJEDU/z
hnkLEQQA6VhYGk7/hEZGT9gD+f8VTRmjyQ7INVHHz7cJDg8txTe4RJaBZfOpjV6los541Tf+xdRR
/B3/hjSfR3z0GHBhvPf3SLYY5nES5x3DJELg4VpaOkar0GnQ2xeWV80PahNzR0G0kM3MIpy4NGWc
XXYcSe2zl4uW6o50pN7u1UajNzeAADUxbNeeoLunX8q5pf+E+PiJWGWMVxg7v1In7Jjelm2hl/un
Wgsdc5dIBT+pymjf66OVNlr1v9fq8tCCEyB68JvzyuaZqW/VkTR721KCJPWRYpDf04hTY1DkSxW9
2zN/C+2ElYKw5px3Pkb5O7vt5usDQbEAdSmLyI6jznqmp2s20lFW+Wue29J45gGtDzrIfVm5YUsJ
erOP697XVRDB7021Vtu7t3gwG/wpRmiRglXuzDMwSk59UnUXyRAZYhHAs/DVOe+9O0hZQwcs5IaD
96DKE7N2QnZ7nMcfl7Iw64bJMgPfPh9IQzSTKMfMgbBIGb+sQXZ6AyC7xlmy6vNA0nBgZb9wHZNr
ZNaTH9fJG7snzJiawHjnWwH4OkZtI4P2LT3xtkseP+X+ZpziJpLuy7EVT8A3JRO9J2HzKe4SgxyX
u2wvfqXpr2MQDfqQ0kliP1aP0b5hsMXsv/bLWi3DHoJ2suPIqJUNrJtFPKTDNDUHJ5JbXzyuj0WT
47JNpVNYne7No0DvEwTf6GZxPjjVYIHmKDXjBC7r+YC7t20SwlwL4KInTzOxBUSd08GRRcApbGaY
VY9z8QQHL4FF/z/VsYrdDzkHoz2IxXsCpBARjahbxB9lNuVGa95xyF95bnPtLj40MdepoAXt9Dgn
dHqRz/b8xBmpt+XOQr9l2vzI2/RFVl4UTo6ZpRY0xxU6PTCoCmt13q5l6ckLlCP+F6fVmDTzReNw
vmODMLBJzwSWaN8LVpJa5xhZqlzwwfgcpIbNZDC0UE91LUBExOi92dQl/LYwXFjh5x+dGLzjdN7A
8O/3L9pAfjsNzykDR4b6Z14Q+nywvyX445il+8mErL85VDyOgv/vzMnSEEr8RqjhvqQ2Lh4hkhCN
20/GQvKwKSd7KmnU7TSF5hpsXN8E2dT/7VSCwmzg8TXiL6Sm4bnLfAUSoeyoOkXhyK8WWRty+Wnv
ZIHm99YlFj9OLSK2o7Qh/ivsfgHOhRk9lnmtVn4rJaUvfOXBi0KbdZd2iILChqsfSyW8Nt07dRsr
7USaE4SCk++1Fv0TqqBdBRgFN766mdq7sUsBEdMG6tMP343w5Eqx+q0+spAkE4x+ByeKNXQS/Hbl
OcqJmNZTp/HlXCr+X5k/FGM3klR2dgBDTrwwzfj9mHnWLlMzO1hy0SeiPIpZIgGKeUOjeRfIrJAA
J46ri4m1lcy76/BPVC0pUVamNtbP3aLWG2jFV29eKvfDOzQF4puBruufiKoH2sraybkqMjJq3ss4
Eblc6Hebev/FC/Jdz+7/QsRuuWlw7bUMo3qYKleGPH2Ii1q6mAmXqCzKYTsDfGzaMqZ8SfeJ/9RX
OzUUcz96AZU2I72AHKLv7MqkyQXgoo0YGmYT1X+4Yh/GinZwu4ptEpJWAzB/l+VnyGqQ5gx40MJo
oZa7TUgyj1aoWawj5W97mH/RfPRI/BFa3rcBeoWRsgSlczUt1+fGYFV47/Az4cKYdgugo1T4UTX9
v5CAkk0MIIIFnxMOSRZIfiql3GPbX8YfFz2ZTqq/EMmRh+fQijZX0JrFMx0FkJSm1z7lAOSOP9XK
SgFLO2Flo/Y1zifhy1a3Yx1XH//I7atfduPJ8nN6Szvio/KAxWK5Hsr3ZE2yAUtaGmPvqSgzjrZY
vc7KLESxPzffjojLCEzPViLnWt0W23BkP+rgBY9eJpZtn2tS9nFLkEQXvK/rKsGsyk2PKOENocbB
1XgOCy8um+Srph7N3abfzT8Ag4n2el2qpW2ZDmC2ZuszI7EtbUX8oDXtL9twW/8hmHtBEkvVP+h7
zUd7jgn2CBX2veEwIxaqtRt7btgYzNDe6WC7cu+4Q+nVfqzQ69fREVlvGb4TtuAeUE04XJNvbvKk
SBvHEzquXnUNv6Ec2AUdVcBpFkZt4vz7DQf8K4ua367K8lnzgqfzF4fG1kVbbkCPMIVEJ1/5Qb61
1LCBqSZOGs2dTvtgna28C4tgkE0PyPVbpwUKryhJZp0MlBQJNB+ssRyTkyZUw7hhMR6y0K2dUQWY
C+8+TCpuuRIbrIx9qrGhaVTvYnO18OYqmTM4UNAuyyw9/kJr3s3mcH3vazULwTFoo+ZmZPgJByEU
jRx1W2g5Kk9n1VYAx+ACGCswxbzwG1CJPfzsE0/VOWag2L+9dFHTvtGw3f/IKQRYBQyPn/P/1N05
0lcZe8nf3BANRazOkq9uily++b0wRRML5Q/sgODT4s41rxPuY0XiOI93axlyjdK6kMF5YbPf8/mT
pup5m/TCWO10Z4TfZIDpaBh7OVXlb8ywWWOSDboif4Ste8fzls58X37C4Hi+n1BhVjCvYcvM4uzo
f7mBjv4dF2383MtTDd1LqJIrBiIgHHgRW8Ez1IQ6cTF+vmDmo19RW7WV8kVsgaeWi3qAej+VGY42
k4KvsFfptRhi3eZ/wF6p0UoQ3NPFxSwTP7xlk0IsOD1pUOYN0ybR1qUUqvil6zLJ3v69dHH9roaz
l0lwR0aZXW4F51xOOmWfuYbZahePolKm1BgHkGw888daYchzHNrgYZpL7MPRMcSXMqaVbS6sxDes
G0v+G/RznL6Bxyuyfwz8scADzwAfb0rnjn8UJm3E82NPbI7BYGQlEgQZ3sr9xXIY1ooGprGO80Pf
U2nEhGxhm0qJpXh0E3JaQRqy6RkjIGcMc+v3g17krXXaaYd/iuiCB7kjJMDwq98SX+Noh8CtjrZB
atUa2pyRijpKxpQda0rLVAa8XDbTQTKnLPXEdY4gF/HtNnZ5tkvKkhBZRWtA6gTO4eJlHfdxkeKH
nvgLeKquf77IMM3QHxynTqf7ZNHe9ePJWBo6c3O81PKo6aVOvoTY7/Cg17aCncLPFFGnRx+VKgpY
vJIFzbWtk2P/QiYdiC/WeABVSCQbwSiF+KEuqnUQOR0ceAS8+PRyRuE+6mKCkxFxuH9pE7D4t6kE
HSLlxhHef9A3CpYWhVbppz3a7H7jITkte46GTBnkynGjZ2ZfUraurJnx05+p0JidThbCF18ZCoYh
fhmfOH/zANZasp0nosrH4B07j5Hm/743EhFW0GhX8hWGdikP5XUyR6ZdQRtp1J2lrx8uuSxb+l6C
RAzEyNO3T0PZwBCSo3cXCh/QXV6kmbior14wVXMLs7+zSjXA5anoNGDjnmypsv6M9tk7ddHwPbzH
HGAZlzSnpijceBm/kMI0kdcTa3DypSVKcx6KPssvPNYZ8fWbiPW1ykzFV4HkLIR+bQC0MxpwVM8E
vEZIShHDrBY9cGu5Z+ACvUe0C7c3HelthVl1hHRt79AMKZ9FxdeAU8F0xNsJMvTjAHLXbP93hZjV
Ho1ZZRIzBmHGrIUTg8P/5SUglhzXSACm8jc4fODEx3Kqz7odm0oUnVQuT0xZ+xN0x4+BuDToreC3
T+peh8ykOdv78T9J1qF8e5BRt28XAWnEJ5mhGl1b9k5q7rzzGAW/L3R4iwzmvmkUMJBV1clWrLj4
59mONfBnVcKxSIsVyYKy9z/OgrNy8dhYo8D4E6E0QQpwof+LTt9bK9L9aIK/izlgG+ur2NHVnKVA
nes7Ua3BBye47ORbvhwx1NC8FlumZISRnBpp/9K/UhMAVgVLMNqF7nUMys8GfDVKXVD5nggQyuMj
x5boLgqWBq1+ZBzkCvCXn2JtkW6t45hNcZqtRxxuXS7wB0bDkR8SA3Lhqvl+5KDlylFowNmLSn9P
Rb3EikSMxU2H1lLP1rT6szAkwV2CPCXh2ZILxyY7JmZ559CTL7M9t7QkKfFxWv7mnytsX1PzVY+c
IlgqXLizOPUSYI65le3wPsE2P70vdWDzG13RhLsXxNsyjFKmN72AU6bY7V9Oz0oyt8lFuWiTSNFI
Or2vyUxxh76KN9Y0JbbEelv/lsW8ooowdNHjE8K5zOrnS1wpGeb4M4zn6ZwzQq39kT4gNv63cHgL
ciS8wIQrRhCnOx3S+YMpUusCN2IvmQ85hctWjMODvo1H6vgm7KbMBSIb5U4pxY7umA6msADeLqi0
lTMrUx7QkYAuZscFxuWuYRt0rSb2Av9lvBUie9Bp8WW4zSMxi5WMGc9gbg2/UHiuHFjAi+2CxBxS
kA063OmVESYHAX+KjqlT0mSkUamJ6kyOgd9Zsh+yiMroJkCgw1aIAIK8gzXMwwinjiYs1xvrPtFM
MScSgA7Ah4nqy09jvH6samtL1S87k67K9Snpp80xia5ScWbnSkq5JL8yAYQvm7X9DvEP7XmgOa4u
FQ8NQpie/SkCfn00GmucyEX3w2ppZRWPM06S0NOsfgWYdIQ7YwtrlxjmzoInzupkm8f218FmnsMR
EDS04Azw30pBxBYyi7nq/DGG5LwkaZp/Kh578TnUUrnj787+a2rXF9Rhzc6KIyvXAZxR8r6D51To
5IuWhfOAbm/QMIBGMqoPM0cxVsGxD7GWjMT7XyAKsgQMYO6JSTc5F2C3QkbmTPdMNCoTjhwftyKy
qGMr7DOhg5S8EjhKlUh/9VAmdrMQ+6sNMo3c2JOuhnNNfcYaz16wVnP6heK3nqIZhyJVB+ewUpj3
JRv17iXvwQ4CZyGJJrH204H6XfhFZ1raVtVG97qe/592MqLPe0eyEgJYHsL4AWYdV2+GPDm10HjV
ThaG8Bf3pvBR1jVVUslp7iSdyhvT/hgC3i/QHiSNO38cGqfGmbX3eeSKKIAS/tdBYnvGnQQiwA9A
PI7+uBe8FxScaZ9Ny1LL9dCP17+Cwh4o4Gezi3+VFYCCoYG3UYBoGZDZuy07tGPXAnFDdN9nyEF0
CCEijzS5CI2QYbhK/ps60jCTbuuygUOIaafo0t/gkmNmjRARX2GKErahT50JYp1TK4wsR6xwNlJ3
X3mDwavcPAH3hoqT+UhnM/ggZq27QjdKshVLo81YDjxCzKTIB59nDMswf0XAT9DHrm/25qg64elk
YAGDEBJbwmWEv4LH88+N8czzBNm3om4raVbvh7/d39g2/9SscxJa9KZlA4a8jbjSyeRjyuE0c2tl
h1GFGeN83wLL2ojzrAvJwg16iuknFhzNYG1ssjIwTVRSts6q1eQ0hwaThlVj2V8Iy0khc8Vljwl9
qE//97b4orUfe7CE/VlAfK5WoMeFh8GdNkeI75r9lQgYMj88PC1JfHA8OzdxiZN4ucQsMIQOgeNq
NmeZo2D6tZGhzrii0SGh4Q1Z1FTmeRTI+ngg0c0CUMFENI5DZG2abN3Bxbfo756DbZ3+li75h0lJ
WHczT+ps8QXBpQcIEW8eEOi4q4nUobJXp2/cMUxaeh5tREpIY0/AmsIj1zvrRrAE4Yj68qQflkH/
YXmsI+7NA8n+IIImTaPn5r5oO+v6/7+4KNjjW8ll4N8DOOrUdk2xjJNejT7tuGE6jUF3Ecw3c89u
pz1jBkuIbdHAHRe6DvFdGaeP6wzaO6CFZD/6F09r/7XJUNtjghtzjbBWTb9NeBOzakqIz5VwM5IO
abpjcw8S7jsgHgHSa4gg5SR7LpYX02Vun8UYWifK8cLIqe9R2Wy+y2+g0NdIIsUwiFqZHsnHprxc
3lpuIrOofaRpm35TpAhgZx/4JzM8xLlRIZpoXrw+A2RlvMkTSGipDHihAxB3wnEiCSEHiBMgtnKs
VOy76cUMn0p69rdT1zcK9TppKsfiZ7DiHyRb4/9HfciyB4WzgH2SDdcAdYILw8Rdhu8rmU3lDrL9
kMFZhTwSvf6UJFd9dof1jhyOuHnb4MJz1ZmMyxTQMxD8kc8sXIv6x2yR4R386JwVAWO+cZKAr+Rz
DoZB91hyyBADztEEJpm8iiLGePLD27XHAsuzpTz4QaQJGoMR1pFyvToulg2pRJiajZH3SSa++pHJ
dLIsXRKrSnpNnww6lbkLVW+v4zQvDtZuxGgFDt698mfVdYGrguYa6ytJi5yB7/Rpm+FHngu54Gwj
FaHsp7thi6nsWRW/ODb70Em5O9OKozKG3GAMqxYoDf6OLB4eV1yyTemdJnW6UcjgbHPI52XEvZLE
3qK9B2Jylj+bt8aIW1X2qr0jtWJb635HhRXCLFcx5hwP9rO6C9EC2N+u0yZkvmG+8aGpnz98Vut1
esQTTGn8DApj1/mBhkU/FqEzpbirKN5KbhQPGZZCxi3EGHhqJOFVmsbFgLsv/16aibWUEZHo+quZ
FEQMFUMLTMVCO65bu4KhKGViIUu46uiRcbWQE/WJGbp33cJLBvxHpqWn9/d3aH9KdHAvnyMkOlbn
G3SS2/TLtjR81J3qFaXidPOSOCiBOp3StneBXyAgH6xsaSGzzH2XiA0sSEegNIaqDxvSC1A8KDbu
ycNNTKDwfwyPGYwIrUeiLfmBLbuaSObgRxEXhW0qPCyyxIKXU8MzQbPU10enRMtmWexua37xp5HP
BmHoy2s31IFL8L8nDhOpT7K8HHsiEivaAsYLbKgRPULFse+OchdCWtJo6Atz++vz83EkRlkN4VEC
lU0jYt7BahGE2JE/SbZEp4zsa44bTqC7d+3ytAeSuFA6+Ue83xtA72JSiKA6NjlWgomWywBcZT59
0OfYpKhZ6UQVMglacXDxLfDPM/RCX2Qa+GwPEMOMKmhtI4oaEnoJhe7kyXixxl9zxRV7rJBfMRqf
NQAgTfe311O3K+Czwk5kb/SZQwxcBsSCCn2eDwq9jZCATzeKgDn9TY1HzdyebizFhqkR9j1pxXlp
Xci3np8wWsFpoRnwjK1MEFyIEMNYr0oa1dCIIfoaikAyRg++gfxP6ybESqrX62HMPfWgcehiQ5j6
ldcGpW3MORibuCSbc6/WE8nPpBSgCpYsPrL1qzpeVKWNWga+EmgUrYjxZJSxD51gazWUAWMKU8nc
E/MU3i4RwgvW/bvKdlwSauq47HFW6kPAGEb90ET1qLHtrsexvBWG/EBKsKq0Du90TswR0+CGSFbI
fLVqriWw/pP5g+GkfWsWhIJa7juaDQHvt2iw9Y51J7c/VPXWAtisTeWbF0oSmquc4zZhEh97E76P
Ezg/N0nnHpVmthzuDDO6Q14ElFmewKlBSAkEJuJeRLg5uZukGHmlK8VgRJ/HnMpPJsMEKtDhk0O3
3erElb9Cg7j6W2RKBsZLEQWgYfFhXbrwdUMZiuFMSCdqnQhJtzsu6/c4nynPqTitxQNS7XlZyRZD
RDLu8EhI4YihG3J22Mweza36cBcAFMPWgPFDAfN6obCrHDXiOfSEfAL1+KcwLVuLGL472bHGx4d7
CXKcM+HgIE2GEbBTL1LQYISKQA12L2L19KmifuOCG4MOpX/y0Ujx1sIrRZHQi9R1WzpChJy/N838
HnHnR9yJD9llqZPJg8WZddu4GhxN+0e56XxbY3JIx7fS1GkTjZCsQzIu9y6kjsJgUwtJmpCuHq2I
Oy5vWBUw3VCQLfrupPluHVB/4wrhEeVULoRVkRLsgziZlcXv3RqqDm3zS2t8GAeE3vumxiC6JybT
yoHNb7x/ZCvFwH//33gpPeRw5DOmxY7hBsCaneNiX4wHr6GSEc7YHlN/QICMOZfZeg5cADy8q8CD
P9iVi8me+DIxmd0vQM5b/WDqR0dDtZE5xpu1YM8bfAtXMda+7JRpMFnVrqaJqofUBC6xgHwwimaO
hRAuI9FcZiCx+oTchdSzqsIbw1DXLfyrxKl80NCoKIAi/XOgLSwhSrEnVxL6vc+KBMf0t5rWxpFj
JvbwFKQrN5W7gs9+d+nNqWYcJZyBpqJykLj7dXq0sNxtuVRlhrmwYi1O69TQElITg7HyWC++9S8i
ZuNQvJHLsOlLUd+eCM0fQ4ESG7NeiVNuRs0b21jdXrsg3sXoKdyk68EzQEqQgSG8Z3JTr9dmBvu4
WfJFFjBfeYxw8elVRMBJUVVrse5HxgM7ULrTi9lKDJwuLxPrd98jUV76QPPQpuuBRnLPcegit+8C
i9LRPD4wYBt8pnH8ObmLc00BSOWtCpCbKrqkEnMD5Zt9eNTCN/bFz7vuPb80Swu/1Ci64cGVIJEj
nNUPiwrZCdWSa8CqXtIz1vIhFnOpSLEsVRczIBGKpAM/SiSe++ljXsF0MbyBNNuscottkKJXwN+z
fitoGxbLYcPYl1/Sa+j/2qFmDZMe6mbLzxfLlXi4C9g+J7E+87/j1wJMm4xF1qNrfDF54i61wFPs
PqShN+cW5nMNOnHixs7v5r3Z0AM7yb7Lhy1CwPFkg+xRJtx3lHtTaoD9NV/R2757nAfb1GVvthdT
eSiD48mC/zmhyfkVOoKSe93MFXPIqbeWpQ/pkGMaT/3cnd6botPET+bUGv6/fn1+YGzMwfjfyCs8
l99t3s2kYjUi+RqLZhSw2CoeZCOMnctEHiWZ+e2qXTgcldQtTgxAbM9cF0Ypma4sfm1KTUul60SR
C1MSMMrxgC7DqsFQdPblNraTQN26/+eMUAzoB4cYYegybYY9NbqYOpnBgzeR1qAVMPz9OBY7ZFFA
KvEENwrgHl/zPUl3Xf+wsYY94g1XFucyjOcuTF34Khzd6XQrUIbhZ3fKNTNva57JL6BlSM+eqrEp
86JgM2H90R6NMbBTukc7AtPl46zX65ix3Tye24MzMYIqy0YiAATOyvHIq1UxDl+v4HotM374pqzY
u76b4JcwRHrO7VBrtyoHx8EPbWn61JfgPHOc8Z27rTTztTvzwJHgXduLYBR4+RGmxxlfcFm/7aBS
29N5cHoY3jOMT1hKb0t+KrVNOBVwWDtBgbI+q9pHHLI84y7Oe/JJfNgsFkpID+9R2YGZVJE29F/P
JxhsOHONo+e7aFd/uDNasEFhgaW7olSkbkDboNHSzgoV7NsFM/rf+5UGvx8ETFvYhEprohFG9SP7
50FfQTLhbatD5pkbQbHp1XYkvE3zOF9rUOu+W96UDO2J3clhaxKtnWWQ4wC+Ak4sUZ6qSUqrKZp+
IrYHJIekDXGla2YyKzYgjWvQsJbfz4UHk8otiMS4PuoHS/bpT+laT9KkLUGyi9JInU/o3vjaBJQM
qjSASySPfq6PEDsbQGYVUt0LML76V1PavHn0/JolILc7kSETB4fZXlaqbVarWh+ud1WY6quudpzw
6Ou8vwEXVLMiGKWKvnVR1vCaZhYkDvnGO3pWQdYKQGGoDcuCgdO4TuT7n7VqxmWMvRT7SABIVrw8
IVMsPzhq1akyOjJB3TaFLNuE87NbMvHvsvXSX51OPwQtmPu/apD3bfyaiI+HxlKCjbI5wzGTBlzn
oE0jA4mwkKz+gHWUZCXEgiqYTqxKbHE3yGSEykqq4SCBidPZg19pAana32WMVPuFrqCLUGwOfyBV
N96hWq3YWGuCR6cYoldsbRjBrXy8ZRjSSY7C0ohdsqNtJQbNp6F5XBOa/75BfbsyAcZ3ghi0WVPE
xSTZPZAEMJQ2llRVK00QPnBDH6j1KDTi3Z5LhHi0l2Lt4OpQnp8JmaVPAdj/KRB5AJC7pNxrxbwJ
oC21TAictv5bSr9ALYuXQUiN4vwQItQeQpNtqN1wxmQj5t0nrf3a1NZ9VkJmTStiEaM3YNGxoAp2
fL4xoDq5MRcRUyBwZ73aDzvp8JaSM/g2txXYiem0U2H76ugGQwj37KTAxUjiv+NBQMr4AphkhbRK
qIbItxcC0pHA3O9NUZMPnF+cNKlTkEIyMfjv9o7c9D9Jzvhc1PGVPfBXmzvRKFdl89hzs9X1WXdB
fnRW7990vMu85GGUQcEAn9sEoG4rfm38tusnG1WS02zSegEISJGP38u2V75z6yFC1veGBSmMYy62
UxfiCMavmiiBog9kdBVh95ttRfQmGpdLIsmwJKWYR6pprsDfPleBAjH64YHX+NC3zwcQeb8MS8eb
cZDSFfKtoZH3mgZriN80xwYoDMw0Ox7wieHveufOX8kePvmZXEKZ4X2aM9iE4TR/TqQ3px0yYObL
+WnGxFHB6H9oItXVrvBmoe2O4uLn0uS0EwQRUpN5BMNSoczkLqy1glWuUYeuy6BdU7EB8OEJHBRL
yKUzDzPN1CP3YTwzGYLymaBDTpAnoNNlVeYW/eH10PXHgtKEK36+2R6U6RRcFgYExAPguM+7ffOc
8wtP/jk8Pc9WZCxet73ytJiEilDqVfkAX+i+3Kc5ra+j9JdtimerYdYur1a/7Ous6u0XEQcU13sH
mVxQQeE3B1OHkGDIUR0nztjuGras84uhiZBOFHK0tgW/XKxqbyeq9WBpBj0/ejyf23W38wpG/tdA
O5qYONj+Isru4jfaBEhFo4dql80Ww3Lv0ctX2MuD8evVhWJFbwNo1VT+c8+5x5Vjr7g8Ro9HUT4K
xBAd4Z8KAJABZ/EjCafdFnf0JMnvhtOgO0pxgUzbsRklpH3Y2WwutzonzKl8SAHI7MFsmTlh48ZG
5OFoK9EHuBkARSSyA2Uo3NyLRZxpFG/8Q6HwauILFbAOcye5mlquB8jenhGz4msnbyx4xc1kdYq4
A7FLtu92VdMw1Pyd0JY1mrnl7PfjgaxanaWieOk5JOHdB+a1F0DvfvhIHhkjioH5DMAF74rgLBxH
01VRiGWP9WxZgVyiyMMeeuMfRZ6SbQAfuekT373Rsdh2VhXqVd1/T8Vx1hvoGEClGmYuRoXlJ+DS
WzKuMxMOj0D0JxLqEzULl1rPGiVx2N2tiYICn+CcqolkwHF+dvqmoPTBOrKKIJIr/P9Ijke3ZWig
+CTkDfzfTAI6PhfZKVP0P+145kOhHOt1BdCBsmjepD4F8uMIuo9Mt4fIwhBNcD8aTxbeixSvnTjA
ZG8qm33G3u5kPpPiXQnMHpEpue6faYg8V8/xndKv7NqB4QPm4Bum0KdMUtFABsWE5Un13NNklVKa
l3pULfWJ8lDO0FT8JVAk9XcA2GbljywSoeB62C8aNvX31WMEgWVY7UOmJE1q9+rBW5wvO/GSdp/r
moz80VX/0QjjWO+msmG3UlAPUIIMd1aAifM1Iy2yjp59Xyg1AHk/+iTOl8zWqX3r7b8bVkEc0pSP
BUSB58k0IrvMjkJlMJ2tIoOuHFeQVMHi2EzPYoyeFBIvs3MkBOX/dDBLOCMO+aR6tAIxl4fLMYs6
5thgppVUIrhiTFOAwhrK2bBZqJUos/fM2CHmW+BPCjRnc5bwfyBeiRzFXpD82LfUgTWPE0vGFnZM
qkjBjsKu66yK/eSpTuFy5ujQYG51OFUCzRcms4foZLxcGs/wxVg6A4XHO7m9vo5cNU3vBKKEqslP
wPhUrv9+zNIWQCOR5V6hPS+lDgtyFW8v0payGerch/kfiQeKMM/k4I0xQhgfEMWNdNkNFIw7iqa5
dpwW0Kd9pBJ5H31sxz0iLQbS6AsWaA5gy6SoknosVY6CBStRkc1+AB6zOEAOL7pUoiJaJgeckKwx
JQlavlKsXazybqbsfPiu+MATtF5JTF1rI+CxLsR2NR9KNQrtMa1yQCG1EhRb+2Z/twYNPn0dae82
OKPNjdRCfBBavFMyaCZ0LPeqlGU9TjJ+6eA4dvq6HjgpPdp/TUTdL09zJFXmgmFSINtq5+IftVvD
1frtNy8EXQDrFhu9JjepoL+MdS9reyUVX9foXcPk6GWVqTTdVchG/vsPCvLsERG0xt1s1g9T6zSL
KFptU/0vhFvNZ7zMwUx3x5DivOK1dyI8ML9y9fB7sgpGNAFWjm3fL/HAvCcs5hFxHhqg9s0Kwpwm
2IPgvTc5LePa+t01v4CAs3AlrPovhdnokTnTkAA+poV4/tCXpKqyjzK1s3T4IyC7/nSZB7yLod11
5kefbjKwUBVz1dmjhcdFkK1PzKcqqT6lLm0crwjLZo9u9qWQ0LN7+alZiCkTX9UDwwK/nWk5CnLn
pL9DveDQ58ojmQVqZ94DKjoVR97ll1m7p0Z7erBgXPBeiYcy8Zd75hxGEqtCzQ7U0UPVj9VMRKWj
TSUADrrabpWsK/0UlvDd1Fp65wediWlbZqtqYY05DdcVGMYccU2kk0WbCWktZinru4AOt4rbWjTk
BGyJRa1S0EeFqjUobm/7ZyUhzqGmhKHoK0CA4U0ZxZh9Dk7w+3+ivFewC6W20bo0nMm4+ibRF/Eg
CgUa0lIG/oOihuYw+1LqE2KEeBZfKm6Z4M8ak3N25YUctRCOwS63ad35WUlNJzIuX4gB4UFT8Bko
ISGT0nUgBW5folkv9JSvIftWHoqRI1zDK3o+jsP+zucs0a+UIL22EUPvnc8NLWterdTWOoQ35ChU
42hvBo4fTY3Xcn51oVHmSEmuvuGVsZtxhDYoCe6e5LhRBeQgbZRirkmja3Yz6AuGYKM2LYA6apod
emMeZbslJXmLJhNtN3QfwMXWx1DTjt8k0ByZA/lYADj3UwcyHXCvNBKK79/IkCT5LkqLF7qAw+6w
R9WOe3aRpyuJnJhzYT5+oXbBSrShknEogsDeJnxziMtn1g38GR439MGEwd9UbGWtuhHF/H3xMPen
sglEbEyU3qZ4L3rep7+PM0Ei60oeB8bB/xXD/R96VS5YLMXxFv35dFZUPZdKxMGC/KdEqtAzOUcj
1AHNHemFMWjoC8R4QOCcZDKzJU45GkmCAlAqRA0Jh1QAeO+p3eKfv7Jf84X48MvVpKhHblXaQOrT
KlZO2MQnmihgdOEt9cZk1ZL5RTo46gtQsVWpdUeuxPK0oVh1b4978sHSG85i0geQSdO1GAFHW7d5
H2nOZAeRHvAv9fhz6wWoRrsQP2vn4vmzQAL8QFgwDhyBPjqyuXzStA/tTil4u25TvjDZbH4yg0kL
Wah9oeg6ghEUDJU4EYJW9O2hW4hfP/SeBXkKTBvNtKtQWRlnnVRNnYjFAsxfYa7vZd7Qu9UJyeKT
oKJ927lk2ObTHChUlcSZFhm5B8jGb/s7mySJJjocAFalNhkW56fxAuYzJko2Nt7wPgp7lhY2soW7
+I5HYUzAVEYfC/cUY3nTmVA+vKAUdo9OQFyh9DkYs2r+grD2aCkkI8S0rXgKutk16Tu/dpN/iQsn
5T2FCsmr7/2dapHO0TBT/ObtLChCbqGBuV0IkPPc/o9b/C8NpPHT1UcqrYwyTs3NnhvMI8HXYjO0
Klx/POz7grrPRcwBT+RRccWS9VCbf8OzXfPQWjdTrxifwdoFu/hjwB8ZMi3ZcMT664XoGIxMFjAj
TvCj80ivAS8Wa3MXDBYCn/DJxkfChWBp87JW+d4/fwkZNMQcSGyn/HCKuLQemKPGLJESX0d2u1U6
kqE9zrSGRqYQXGcw459SZ6EpU2QXTc+tZuEC/HdbAl6mo9WUMQvS2VttRXl4X8EE4EADH+tybRlA
jGatXJduPAoKGqOTYB7sisfkQqeIF/se3rO+/GkvQ1jQUd5aKuQAZyuYOcwutjy7axqa4HcA5GXt
Ya8Qu2UuMV3PeJy/2Nju0L8Ar45/WCrtWIBT9H3uz97vwvsHv18mFUvco6qzq8GszGpZUTwS21AY
j+EP04GsF6ri31MmDryWlq9nPK1wkQWlf+nJQKzf4/95mnKHScLgUtS5/gTTmqwx0cNbAkbI2MnB
zgYn+N+3Rw3ouJlYY+K4aUMpeunKyfvDUQBS8yAL8s4pN4h6KoS5cUFML0vT89pJi3Ki7g3zfepu
agZhazYlMzS6jrWDhvnLOphOARAmhKU7aSRASOxie0vqSXHbdwmiNz1oFe5WrGFD73+XLLBTHD9X
+XPNzLxEm/IAUaHPTgdWFvsqY2o5UX4B3EYKKCxG1/olsVRsgTEU+9fhMuusG+lEIpqmTkG6m4c8
qZ5+d2I1IJvTM0je+y8ZyV+p5hCEJATFgWJXUzmxAz3ipuMplcJn1u8AXU8r1veRs0vb18+ABPAo
pOcLG/iQ3mZmrj8gEODTkcT9wDgm+E3dEhEiYy746OwKW+/H+/nrSuKltnoTG2BaRk3PKDq0TqwJ
gPLcKxVcqh63XKkKyFZCsjrjbYf6FLny3mVR/5prZ4whcz8XvjD+hqNNU0zv3bMwJoP059Bkr73D
bgk/LpbQ/kN2MH+iDmnvSWLpn80HVl1xEQ6OuCeNE4P2QHcn0xvyabWH1ai03vJPXSXy2X3ai7pS
X3dS3HnVzzO7yNR1IJanzr6gTxb0Bv7c/HbOqAojirq8MGDwya3o84b/ZsCQ3dnuV0kFrylGoBlX
g8ESZvRH2aX5bPh9T7tfeNg5788VbdyBzffr1XgCSFTurgj9BwMjqqUzg7hEw3ES4T3aaiN/56nQ
dWc36Om3fdc5b16CnriHFM90/njgZY92sW0DFhrBBokW4nacDTUqCxUpscuNWVTwRRKUe6MUxw5k
8YBjIGDPdFmt9bH1mD84iVX2Q2tCNKuS2MP1JDs8HE4y/W2viA/4ZgedFMjckRjyqKUAgedQuW4O
j9sMWo3uODOSVBWC1k9rFsJcIw6+OddQX+GzbgQBClB8EibKPTnovStmBatdqrawmyfWtzk37h/D
g4f2/8h4BLIFtIiox60BQznRfEgL5Bnctt5jDCXZ4heyOQfCmSxiKdNeQa2kKiKsUzJEMnhjvaV2
+FU/BL9jS+W8OXpoZUDc90QpZH4GTqUa06WrrCeGtk/PKtllyzyUPqLdfFUKWrF9BZ6HsWNcoQko
LIS+/hd3Qr+uRmakhMK4H/8r9/hWH920XxQ8Z20zOIk5Crf95tG9tksdvGV7+vF2nJRfVuJVGSUK
b5J/aop7Jp/mz9JXFQlHXMzm5EjvFWa/c8u/NKmID236puLl+GuWvl82ZGThX7vYwSqKkLa1KwpL
jt3O9X/lnRbT0F2MwQuFSIw7hcZA5k+2fZzAbVHllDHF68UNc3x6sF+GIGf1cGA+nWLEpMifcRfH
DJ9KiIE2GDkV8dKMxO1oCiVEg5y+goDu2QGuLCUHEuCk5DoWfQfgoLBYhZVssgwy1WxtISsFLfxi
yHZXWzEekaJIfhcrju8Xp9wJP+JfnpYMkmpGJY0OYsN33FwS8yVT2sa8Ca7D1Xjcgv2bopIC2KP5
8cnEUi398zQzLnKSOg+C6azFHWoaaDTXDAGJCiuJNM1oAObJqT6dcJ2T5TtP/HoFgzTiFDU+WIva
9zC4FlQQxJ6KzBG5WYGUotSqLx6Hv9tYH+AZdb5xUr3Wos6qmkk05kR2NVk9ejU9st/+As+Wnl7n
R8bRd6zl8+fu/yZ2q63Hgw4mfP/9YjIKUyEO/UI1GCLw29Plqxf7K4aOfoRd30uj4+RGUKkQGv/p
A9DobWZScVR7zUbhmTlijcHHtG4UxfPBhz3Xt+Q/PqUSDzAN/Y7NpU92kYEGRdmQUEFbP3ud5LSx
BHBEZXvvTAB7/SgZZVbx7wO6uH218OLU1fyWrSU4nSVNbx/Y1p8dXFJTqcE14YOG/GF2UMp+cQfg
rPORTS0Vus71GWTYA6QA/i92DS3aqT8BVjJmoa92Is4T1YBDXxZVvD4dl0XRmUyeiH6NNiF8nJ55
HeK2H+7boYDWN+zR21YcoDo5RxQ+/mQEp6ZAiwinrpJQAiqaJFGuAFi1jVaWL14nXE/pOXTzmGd5
fJPUPZUIL3p4nZJL3fFmgSQgARhRFxw2UNkI4/PYBx5mokQPH3vqiqbut/1UHSmGI6eZF/j1QJBa
nLdq41y8uCUvrAVYHxxScbZ3sgNbDmHPm6swQf2tHcYUXk8U5g/P5+7hHlkWZfU5MrsUM3diWdes
ZlPKYlBHYcWLfuA4jTK1iSo8joqGdrpsniNkniQgWX6TvdGAbmu5DF9N3Akv2DtB2eUckUJblbQ8
RTppKKralqYuFbvyF4Rp/kI6q/HaWUQr3V1uOC5tux8CMhHJf9+Mt0UUneYVBCz1mrVFIIBQYq17
85/ZXsFUh9Qp5UnlmA7i8ptGihPybx+mPi39NUtQEtNDAmTb0leVHFR5RVK57qOPenKI8iffkPIJ
HuPKLd+FXf5DhNkHDHcFoNm5PJ+n4UjalaEmqKjE/HmOQoHxNuV7QN2T0AKWgsrkqT8Hs0Gtkhxy
HmlwLM3tdbSg1mH9N+MDFMTuGOdipSURFtWu334Y8swBLVWxoWnI186m89iW5pNroQCMiqfP9640
rRo4hEAyKli9bjk86R65HQSy5SFc2/nGgmwZl/37DYGOTYsCuNACtolp9REi6OJ+72/9bGcFWzGg
vsHN7L6SJnbKk0huwxGbv9B25nTwrjDg7pT6DwJX7YIUin1KEia4NUEsNQ58ao+1Wvp7DvUSxX5u
qCCYO5Foqf9hPZY7lk07I4OVi/UL//vAJEGpDT6bw2F5SOH9pZKym3W1gy01v6rBxOmjl54Y2O8i
QoXbGmP1b10raE6W2naaUnEwOe1vBg5ukIv56kHZ95m6hBJw7HMQJVdQeqZsqlVAfyzwxuwdQUqA
vARbHn+vpYr4Putq4UV17hw4EH8aRj+ROpfJMCpDMFE2ziA6jpeMd70Xe8EXLkZKA8t5kU0NGtXH
GNdiAEMT61CapymVlTUMl9Z9BI98k3LmjsnkSjsVTOUdI5GJTofa3eflhFN1iP6n+1lNODraCHiU
2KPHgvFIiGm/8lzLzGV35obBrpIC97v0daPG9xg9uPbIfiPq3WViRVyQAgj6fCZHQeHZv3ok/LxX
pXnUQlm2n5jg8zt8dB4Yxm3SlmKsKDK+VVUAyJLTb2f3S21LDA5FGWMUjtZV839WdAq6ErMHm96P
8ctYsab/y/Och7iFnnNsi2duux92zsD4F4qoGODG5pBbfSxIv1KCQfD8Cq/O6uMwM5kJM/WMyZFy
8v0QPvA/cpY7TYK3ZPYyGK/W2b0hW78RlS+X9+kUgwsL8x3MrFgTnCITDtKxrDa3slDgUSBOWjLY
8fRyI+g4wee8BObD75pWgcrhzac7ccICsDQM2CBJ1WfyxyY4wf8tEoarf6ZCR1fWTlzuGP+SKYEK
GPzwW/KHx0XFCQc5ms6ncWmciiuEP0p2qor+quTwdmPzQI4hMGCenVI6IYRQ2p+kn6x8GvFBNnqG
ckW99jkVJaGsJxjmjbHAUfcyB4E8e7ufK4MrJr5aVyYT0ZGiwXZnwkBl/oMSZXApFe84JJyVF6QD
GFXLs+VhpiYbWHuXe6Q8jgVGWZIYaUSMsRtTd5bXf50XYs8CWIwCy07ao1JhqQ6p2ULIJJeBk6mc
oRtm3TyDWfz7eI3GNZXrpLb2Q5/unxwVBkEttqoCcH+BY27hNwVVklgYSmR4doIBCcPedFh49ouR
K0eDOf6CeCBxYMJqt2ehgchRzSkrXiUGyZfFgsIfWI0Boo5XAmLVV3n2qlUyXL8qw5L+/eVsyfZU
QoabJ3Ytz2oBSmVMF3Uvqsh5nNcenSPdyf2YaBHEuEqZW5Cy6JcEHqtVHHMR+irMCuRI9qTiH2yj
qmiS9+ParuuSOK/rK3MT5NN8mqIpp4vc0E+Q3LsOGcAMIKlLozWgr+BzPXV1eMy/kX46NkviwzTq
IjHGQyWVB6RYb2epEE2sHqQVfxHeFmVne4GoQWMUWm3Coip2PMfYBUdocL/wCs5ZRhhI5g/RVaFX
TDmt2EbysBcWz5CInVZz/8ReSGRoogAg+rr8mBUb1b4XKuYNy0WiSS8qfi3SPz4ES5ChAts5T3eM
VANire0WPnr3MHfKOPGpX6vOmfdDawyOQ/OPedI9QLNWorYDIopXr/keFQekvugHIoTJAsKqYY6e
q6TDog+6Ljn+qXddbH+TIYEcA4leb+uRE2H7rRMDY2Bd0J+wfNDj3f6NrH2qmFcGyFZ6A1ySm0X9
P+YxMRacTdqWM81YQWeHTPuPFkrThsPDHVhKQzfAI4Ih7JAh/uZfV2M4o4CCUd2QPLf3Zhhu0Uo/
f+rHuMLf6DcOA4HsJpCBtkrWvxeDhLGY06jjTRWhf2vq+s3dh0GZU84RlrjFNfpuk+i0lItB+iBv
x9frkweKqGOC3NRjikPiU3G2NSnji2iP239tdB5MzGmjD6HV/EpUWLUwVLsA93ikWiJ1CIUZ+l4c
gqUVeU7/lZS9wu8ioQPLucYi4QA9XQAH1lDYVip7XD7G4iPoTpBxEbPRoMn/dOpLJHHTve0Hf+oI
OPxvIccDqDo0NZqPqjPf2gUu0wsEwWvIRiTv2gOIZDQiTDCPDj4LEE1CYFz985gQfRB6qpj2sAwh
BHtvBv8XPkGxCGaPZlbxOS+nnLCxxnGIRN2DM9w9sC1bnc9X/5oWOXDYO3IDx/incyobd6CZ6i57
lL5OGb5uOQ72ogMP3OVf0mc//pkBu7kcI4ZKH5XZXGmaX9tVDWL10k6yUk7+OztUe3yneD0ihg61
YH2z1sfRk50KbQcb8kiolGz+InIxEImo6FBvor+ENlIVLExIK8XhF/8Ym/IzZGAXv1HYniTlEnDI
mGCkmRL9hL5GVeGhr4BJlHDMbJ5NBq37FImSGDfQJz4W2T2hpRB9T80ry+048OQv+XBGZypy3LRK
TLXLuVkB1LK/uYChYSGkvaGuMsdqT5c98BU4KwFexuvS336pqj0Gzx6fYywix2FaK6Yj9ziC4dzI
ek52xHSFvyBGda5+Ya4AjNJOzZFo2t7n3QYTOvEpD3AChHLliwli9wP44U+k1/KPY/BdoP1vP5ft
iPh8tgiEWaE8TzbAnErgprX9isRhE170JJx2JK+O6Utas7kdUbxYOApTqJt5uYGs4aVMxCOOkaDv
5KmhUTSY3CP1pOeVD17+9wir0ZimzgCZMuY1Uld+inuXdRA4gTY5GLNTm5St52xtfjYS9LIihieu
nVTDzNtATL9kP1sSouTfGFfvYgeIUp/pwgI2Ngbl8BMbe8iduaxFtGDkcdy13yKJckYQCxUdo+24
Xwf/izY1F+kRnLI7BtM7qYpMklVoTWEeRr38hFqQ6CVOKa6FwGRXHQj391xJJpV1DVWr4+mxtUIa
kt5tgpoX3drG1DM+dEzWJgeNxn4zihcQJ/ilbsOJIaGOhMMGIHDcu642+zt02AOG0SGhq386aVEM
O0JJQzFA1l2M+EZ4J46Ipd0o5JLjE5iVAWSwpSsApyLmtiXBd0FaJ0iKY9PwnNASn5P9MD6RRZu/
DJrfoi0y3b2LXoKmLMZFKCNjYN/W2YLH/QjgbmTqS/7Gh9jZYEZpYD5HkQwFrwGdQq3aF4BcpexF
nhLzHdWdXSevd0/ioCSdm9IOGto4AmtWgz/MEt+sQmVn2REzu2mr7JTGhVVLWSEtZ5BLwf2zN0jI
/CCkOl5KtYgB3rsEMbN85N8dw4vGRAPEWyFDhowJAIrhU4OyTOTdJ+nnwyT1xiuGU6KVBgkX0O3L
CMf5nzuSdS4KXt8UqyFNM2e8HbajYvfOXOgKJaQn2RLjDDQJNqprKeEKffXSUeFqTkkECuTN1cLy
x759n1LMghE0kCtAHWDnhEj4OPGy7zB84g==
`protect end_protected
