-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zb2GeFyvUEGmB3L3p6ooCAdtZNuIg4Fox5V5pv3hf5g3KLc4Tn/NLw4VQ6Xd9OBw2xSsTbL3ym8z
Lz3j4ATKFdc2G1ml0IUTQSiDkPBZqE/E9m5xdzIHiGPngt7GyAMWLXDVRTKZj1Ph2AnkxQC60hnW
BkRQNKQw9BQMvWb+REUoiXGfy28ICBQsU8bEdUNr49yK4Q/cn7+JYc78LOP0l5O2yl37Rz/vXvqb
mDLl56WimvHWeI2vdRTKy/uo/ubYxn6rQPcSmh3S7cCYYbFxVKJ1EsihhvEVPQ6B318+CNc8kKYp
HRccSg5bIK493MDy1rjRlCyhMwWa7jjne5FB2w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
s7tPpbFulECl1LC7Vuo0pEySJUchHitV4t+Bwvlq0iBNwyYKuEguz/JMNp8bp6/yfFwctgMRmoF1
xC5Ng/J8idPKwzYO1S+F8n2REJaHs3FGTBcY01aMbWyQ5Dxa3Nf2MsPjTRn0lAL1voB9sgeJTZC2
ztxQ3RBDyNr9N8XsXutRkLpvVXcuLlY6PhMfOyQJhFYhMkT/vQsx2JpK8fKNAkN7y7Q3OxbJTKEt
DWHDfnCa2lQpM3JCkL8DSrG14JgGxisHr3In7tr1fESRnrQJas/q1pbd2u72XJgO14nYd+gksWa8
L1yDqhgr7qbDLRpXn2tBzBvNSeX1aqj1EIWMTEHO09ZdcJe6iF4JlWvQA2oVbN60Xn9EG/GWciXi
4QofCEIlM8t/6Rf0kZqVj1j4gdpHMe4Qt7awgI3UKAt6LdbRGbPh2RGWL7cZrX0UVsQ2nrcWDYTL
AWDFxtVZsSVF3wi+QREVUC2UQKzwWqlM5AM7TruoOnyXjzm6XDQqumkCpnrzLZBspHDW/GZqR5Mb
Zn3oVMa8UY57KrtC5k0ogjvUWt0qlCk3Dp8lq9LZ45vSfh0of2WvxZZX+ohDC/aPo7xAOEi+ZWVZ
QUAgntXqaVEjF+pIexdxT+QAkA3xUQ0ynzjJlYTykHN2y5E+L6POazshNfrl+KFQIzY0LnR3G3Qj
joBpeTs6pK3plwnC8UXVjUGbYkfuQ/nQHhRookPKHXfGwPaAl7deH1O0wPCq2805VOgRxEerLt9e
W5kRzW8xqPOlb6wmWsIokkiOhptuEFI16I729Phm5U/4szv0RofP6fGGotWB24ASe433WhHOEkqP
LYgWCJ2rp07FGanYHy3YYsy18zyZnEJZeOfdE0IMO4CnycURx5LgT1UZVMvFfblNuH8G1ZaPQ2y8
vl0yFTaFJAmfydhByTXIwbBpoju6iiDgy+0MfOreEGx68/XQxUHQKzgONghF0jC2tfUGNDzoyNGq
aSX2t2yAXUmIoZW2rofT/9uQ3ngV68wd/he7Aj0f2c2+Famn/54nELnO9J75pYUx+nAE+EsNwowU
hi/I07W0VYIq872jKkQYHvu/jtA9r1LHGMrPY1/Yh3R1TuVLiPmC5setYlJLNi37oow4dRwhGRoI
2V0+gWX0U9fwGvwD3Ss2WfKoJ6WOFgjyrJq4DSHQ1I/l5qtwbem744cwOVhgABQ7SlUL/NWcGlP/
IimTQ6UHXaozrSvYvwOYSDtniW0s++hUEY8tLOfHRJrbG2wiTmumopwcB7GlL4O39Bcm1QGfNOxU
HWBJtMsNu6qLsce79rAtilNrfk7UzjktMp6Jt7/q9SGqWwz57dEL7Q+0aLxpU3G8uGlDOa+pmTeS
bzyK9beZICOAgsWlp4BpEn8UJClGCCCLRyMhb7q6OQed8av4XFKRvo/TYwCiMVRSUU9mxmEnpAOU
DAYXKo0EBPGswuuwjyG/cgU/QhRISjYUJLgJzFxBLeb33CSfTlggDiklaGytCBXIKfb6/8OpoOeb
f9S+8c50DLW0J8o/AEk1UphmR450mvLnLroPj8j5h5f1t4RgkMnwY8CrWeNcTWguQ1bR1LAmc+db
/RpbEh+P8Q15PobPiZo8vGE31CbxUESWstjkPgoeYskhjNKsnGqG2mkTEw7rjSMciWF+r/gf8bL0
Y2AjHCxhGGcMSUHoamd0qxPgPPqtV/YWW7N1YQGwzuovuF1E9LN7V01IJmuU6beKIujPPQAD5COu
wku37Xxh/M6+nGLcZd7AoJtWu/PrMcjSJExUUxxAFVekowHgNQuIxurxb7Z6MTXEz6OVg8nrYe6g
sfjQHr1GEGTkSeQtZsGbaOmaUhhjF/SAORoV03UpvLX+9SyZu7F7Jikb+0m/XcFOz+kMAFl450z+
H7CLwZsa5dytDPo+24VtXEPRX5e/VnFzBTBuJ3E0WSotcvzNm8TaEDdoYVOCMT7oCyI8ezyssZ9+
36a5Q6XwQ5MmMtjnVF9tokzH+LtQbBiTisgbDLSXQPrHAZrFInoSllRg0roYC02eiMHG4JW4vKBO
RwBWor++dSunAGQDq6ny5/0W4xRdiGs1cvNTybn6jFkElXqJZk2bki0K3hk5YeuRgjdoXK9ObcEZ
TtulNkrca7kTGDAQs6mtFjtHllPS0yRyXr9vf+8xS2nZ3S5m2okffYyB9nMc8ceC14c7Z35UOha/
dwANk2eeEoCm5xxUs0MHi8ehZqtxLj5vYkDiL4k6VPxWZNmfSW1999oySBVi//tljWgAl59sej/B
QWv6skCnkTu0bHaHFYnVobbCXtjh8wBYZ/ErR0yydDLbymuzjnMOjEjc9I+H+bSJmZ+MYPbX/bpP
wK5EGDJhjon0o517iSlrq8Rv03EtBj9CL1tDehKrw7b9zmY11Wsqpq3rZs2f/aRrlAmwUDIORYpC
yRcCXQ9GFx8B77e/d8IVqNgvDAxgDU4XFeJn1+Uzj3h7q89FZCFV/XgqAzA2rENbjKB/1XaMEtPi
k7hIXpd9Vn4nStc1tbZZRQL4pLr5mB31asClolekuHD2UiLiKAlSq0XtXurg2Z23xIhhPnXfUyB6
IsnUpzwpA70ufoh3gXKexc78DUdQjCcJtD9jeKEeAuwNmI8FIoFSr4n+qX7WR2xZ1/ehNjnCIN1D
/GjGXL30z+3nTFH7MBqzdJ3ROxD4WVldSZd0LtfaAUNjN+xtCqFZCAGAfFVKmOimJlKU0TeoclQV
vl3z7m4AObC+tuFkQmZ7CldtTSRy71CHYzwWazVz18Cpxv7fNn56+WTac4NZ8d8JKyXyw6XdtQGy
zzZd9AusdCOpZGyQTNOREkGIeGtoqwx+y1n2b4pFaIuLr+bQzHU59vzvpRx3IGLkX6LUJhDy+dT6
QJwXLfOeuvIYeighT/Z0todwsqv2jTcaBEdVILL4mgRRvhdgbI2VpXFF43BsbVjUFIEDEgBhnurp
xhgzXmwuD13cwNXYSwGZJFqP4CFqWfKc9AZxvuKgSmb/9PvToNGCR/6KJNKjZJ9Iqe6n+hLe918Q
X5mUj5tcDs7Kylu8jEVdYQT5iABHl2c7QNrf2XpUkvEF+CxV0/cuyItzk95OtibQzkH07YLEOsem
9vR1/OhATRHi+YseBSMsn8AQ12ZC1QuhgKzSuWfBhdb5RKicfo94M0rJgSMfsuQfjaum34yHaaqv
EUjeRf2E6Evx4bdVdUU9F1hVOhis5XDoVzYqNd6amBFFQBvIagqovgWLMtXMhNytvQWGXFBhQ13b
f1ngAwIezevhzvXTeCc+ryfOsr50wKjpXcLZEIefeB4gMmbOpHKe+upYSxX1d2J1KhXL9RWV8cE+
Rez0kzTUUvB41okptqWwnKwH8PFaxttmJaXSSb4eyxBfv0yJ7wLgZGs6Ct7dXx0MWOawml3ghzUW
I3PwyTTSt8WNmfpP4WngHnrwwhD0c+UxcQfflmFZTtzIOjJK4xyF1XUjBMYuNVKsC2cx1PQ+zchx
zT+VhuQEqiuRp5UAShPwuNeZTKOm/ufGrLm2BuK6zrRN+34EVjgcgHU5zlJMvZq4xQ4sUiaa2sDW
THXIYH/qYC+hkhREEd7kslofMMZot+hep4Hj+39dtGlUZ/ub+rw9l2szM1qINSQ4FI4JALbo2p26
dDkvJubanbeuuMR07u+VHzHBMn1u7DWKGyCToPb/C3VnVLSATWR+wNJzPJeERoomJXmuOtonJLiz
/tcwcLAksoUtjbf5Xkjkv6nOSql//QFx45Fs12cYf77QJxWPhsTqqTsJ6Jk/q/80M7a6xFktE0R0
8DS6lnlhp5wAkzebJOewXY+Sn6Aa3wxXywYiq/lp6dx/oun9RCYvtaKjqXk/rKYH4EimBvvTldlL
aJfYhL4fg2ltcGUGCEfsqbjmPBryIqxL8XlisRzGzHfI+W7l4fAhBPhr/iK3agLzc6M6RTP8qnXz
Lxs5EwDy77XLvt1tdPOFvbOYJLuC81oaNuWYaCZ9m6c0eBQlQ6L2A5Ahg4LYpfMBTpgYSCIplL9E
z5YPpiPi+ZuzkD/GKFRKXOvZGNdXj4JIBfzWltsPz0Ljre1WgTdquWFXouvHP+qXy1OqYK4uZIdA
3TepAW/MwC8gu22A1fFpsIVpMTs9X1hVfPhkS+XNjanUrKATsDtfhwnZSfAHAZDHWoYfzBLzJGbP
8bW/lEV7xwuRP2W37Cmat5HAyuKRHx7FpctYbuEj4FysMvRjEWq44x75QdbdGkjtI+bhtoevn06b
rYUmpahUcaPRtTasfdVe3ZSsaGvYx+5gb7FdqVXQxkua62c1AOtacFATNTe4bm9VixDCzPe5Hft/
/WBU4c6b5WcHLXaBfvST/QIAsobIA+i0M+VglZnMphujN/ETnUhXxXj6yYCLLbxb+Y5FbThQVPOJ
T40+V/LbYNqLkXImZaT1TF5TyS0wLUy70URdtQBqH9UkUi+XaFcKzyzRywEK11gwle4vgrrN9yZ+
yJL09H96TEhsy6FiIXIBEMgWhQ0h3aJmx0HwVjgebdftFscz6BhkufFHnt6qwbcuIH5EI2zoLoNX
Q7JVsZAbwXnwUpNTk6y3GDH8ir+7uafTxQ1weW8UskJbfgfZVYE+dLbdfJKhMr5r7E35PV8iBOgN
qrh9YptovyxYi/KWZN6ztTJmhL2rReNXUzgS3Av2Qy055qOYgoKJZFuwztTRw2L+rC2Eoe6dms79
yYDz7ujQM8V3Xcs6TfWivWvX16WeitP0abbk+gz9EWMzBMPxFoBUXCe2Y1v0+c+dUoWlF6VJZ5dc
kPAvAR/LBEdbLUc/j/XsiPnxJ3+0l5NKtI2FNOQHVWqtERQi5hY+v34du3NhEnRMHYALBBLRyRi7
El06+G0uvFZNRNM83hp1BfeOarFiSFxXUeWp4r+qSLJN4xazTK6SnjUKBK+aJKQop+HGO2RvUiST
jvghzQZgqcUask1zxM1e3b+1na6VYTfHCiuN7KLefO0Hg/orEBh8rzDeyEajSyrAl4SB4aCtsKsh
bsZDpGVWT7CAb8ueFbcXgLDtW84aawLeFwhXfMDc5vIt+utgQ2KJ78xoMpoPMgRHfh1+ZcmeLW5G
A0l8rW8bC9x0LdjpmqJX8T51gz0C5qNOu3CTbDtqbxqS/Ju7JWQWs57Ha6uYlStqBQfT4eOf1dDf
NHRttekINg02CE1ldh4XwuCcNgRbvbNHTz3SXTxPQw8eBlyB4gvokVFJZJc1zxbLtc7r0jCPQnlj
ZHKh3bpnoYDOo3ytnHe+wRLaptG+BhwTOR7OX+ji1Q9zEALySjqTODj0qAtg23ppWwvVHAfE13ko
WlQMXPPJmP2ZBYqOWUE48WZvIRf/nydJuokBNBsbKi+owVXkO/fl9owX/RY0ZCrWUwR7id8w6OlB
MGKfgiIGAElmk0oCtYg5wgBUeRMNq3Qd3jrrjx2sMz5d4Q2c15oHfCF7iGTAI/XJae4WjILaW7E9
ABJI+SYMJs//GnLgbFicNENOGU5ChNE1va44N2wKCVztVLllR5OXYjI3+2fDlTGsjWNo9RvflKNG
UpDBFMCVHA+seclNC8wZS+jFxjLKGGGqQAi00NWK/aksDzJABmiRgb602KDLabOIZUo/OK/X4kXB
B8EiuHqLZYzN1p6yyKEosYY1OC35YoCs5eOnqEu8fd2KvdldaYe2mX6hpUQV4fFfy5LM2yQTiuET
p11NZmvKUkmGnDpKQ4NSXNRLhUUvXIPA7320e72wknVcxJrEciwsW0p8pcx1ovSDL49h5cYolhj6
QAmFIM4LevsJ2nNy4+LQesMdXxdUqxYDcb6Yw2pvhK/LUq9KQAYKk1Lbf2Shq8G7SidDunWiTBnz
pwwiLwlBV6TZqKlXMaVDO8bxi7yrIGgVDXIZGhsArc+AnwxXFQb6pAfvtIYSl8RHATj/dZlrYt5P
i9w0Bax0lZEScKVC2mdgM5+nYlTHWTIVhq9jOXbkXo2EV7xq0xfb8Tvmy4BY+4FH3Mr318gE1r2b
mbpKI2jQoZtEGM9genxLf8XP6e2I+EkDaaBQpHEeZRMelNsRsHVsFZGjF6wqhbmNgxDtPt9p2U5K
puyf4wMXnOi71amf1UefNeh+sgKzSAVuRjlkIW6MiP1ehRKoO/nosRy5N/YDzjqo41g111QYKb3y
mi6YcPsndzL0vrcadACah/mhy75gujxSgv5uBszsqAMFnJ2v5L0JtK/g/1cer52oTmhM1hqYHx9m
ohR+wqbHvAjGBxTwALm2SfTB1nUZqoit556ZdiDnuOmv0jgccsBWA8DcJfW5Q7yPzoOFDPGla9bI
hVScEIZR6BOjWeJmEmBFk0N/OV3W1xfi+sC85D4N1OfrxRBWPNTpQzL5PoZceRGLjGNC3oGJMqXB
whh3NVN7QB1TDvdW5EL64F7QTqylnDJBjt15j9tW/3En5KYRs5tbe3BBWLuExW/8jSWX3C0S2iVP
vgDtSJnySy3JalAdr3Auco3nweEHw7FDynYa1NTGgN4SEY1RkTX/mMo3+7Big8l3+XPgXgz1C3V7
f9X91KbRro1smocBbt36zogHeVnHtTd1YtRen7Si5vEjsi25ho7ITbji+jJDDvddDlvdRADS+dTb
jbRPwtFT8nQlGXPaz/VtjTh9Z9zjZZbaRxZOGXF392JUYJ4fCZxno+3L7n9FgV/fp0OQ82tjEerV
SEqte052qBJvFL81e9ch9YKejpEecq15xbwhvC7cIlRInrT1s72NjCChlCVz4Qfxb1IA+Hstc2mR
fuLX40SXbC4K4QLBnRmHPfuvsl6UMzJHbw7rNgjr1+eDtjF+wsBCGcHFuwallej1eVowwyqhlThp
ewhV91rExFy9iU7hAp0y6YBNzRkZHbY+mJunk3J5wJHJ+inzAQDOV/CF8NwmjEI1SQkwmKZfbjEK
T5EXf3sQR9x6Tsm4rZsCbma6QTKv5wfBTIFRxcskcGMibXl1UYdsop4+kVKQZK57dDhC5unYzLMa
g3JLGo++uoph2J1Z3VfthEOXKEONhWfhxqVdOOOwAtmr/aSiDL4lnF4MJA31AwX3Bt2yuJVJ9QoE
FD49cGYrPslnb2c3R6v8Tu5qoIVOMIZsXSuLXtK1kkAPzUPgpnsegqulBaxLZPXLQnr9Euj/bJLn
KuJQZODBNcZl9D7rZQdUa3zUc6EHRg0loo/nPlI79kdvndjxwHQsqilWJwZIkTuOvHHJujj48h3D
/63Bzy+WIRHyRg7G80hqoltNqkIEWi64QUylJpKqu0+5IUopNDw2XOWgmOHdRNruPQYCdi9Q93xb
NJDJUa4gWRVRIwMq0SioX3IpVh0dGiduwpnAYKsvHgi0hLE3V35l8IX5UV/R5ah0IO6d0iyk5+Bp
jtm7aZo2Bn8VzsteG15K8hNOUwoE5gAKEETs3JDZhahHclPB4EogUGAIRfVeeEvbZPl42O/zh/Qb
cvpyRe3JrP4FNGWp2nISLsIhOFpwNlYxD8AIJ7XSjrovfSt5sXd0ufHbwxVblq5IO6/UYaMQxlMy
qff3h9b5FQ/Jzwu0kTgl5/WK5JbVQDo/OolP4Uvn/iKNcWvRlQQSveCOX/r3ft2u9w3RESgYJTTv
6ebsO2cLrHS7EnOQ7npzhvkF7vhTMwTXOUkezA7NvT84q5R4WvxeY1rYZXvCyRPzjNhyTHIcxOHI
0P2jLCtwMcvnQ5Y43OvozmuYbzaA+zDkBbXbOJ/eOfe6m+pn/SKg8f24b4fGkG98AFBLKELZlF+k
AXN81pZsU+kP8Ehhu2sADQxgH+narlpHCrgn1jok+xtY27uXJ4S8MANdUswYu7dTY6I2Bh9IXnyW
wcWMhBiBAcJU9hmejiaZdk9y+voXC0ZPh/EY3Rn9pegthJS5I39m6R9KgMC5ifFnxW2P+dkwTxBq
4MwOIS97YH7OPQLlceJynRVaP9LHVABMr1YXT49vaPyRMBRaau9oKlzeTMHLq3OiWVx5JJyGaV3K
l9LX0ZTelPLsCNHaGJVLibD0XIpo2/TortgUjJJ9nWSMnYMrrr3dK5n4/gcliPlFEyzFmaz8FgpJ
RM9qp71K0hoMksBdHzXxWYxlQuVT4vt8kLn43C+pagvC4R/pGeazwPSpTILerXXt2ZpfuGJgJymb
xUOzoklBhXXTkSfplv8zU7PnBVxgWpr4q0gcF3wd3/HafF7nSqMV6qYWm/dtN/ieOw+Fu9xqsXYw
prKAxA+sJYR6B6HQ2F1fdT0FeO5jDjjFSONI5mWq2wQp5oovZ2ZSTOSicTOi1cOT4/O9tN7b7upc
hjQohYf5ZWm7mNCgMzMZQLDssCoEYMiOYDCE0RmTbu1N0ZexrNSMT1glb41Ai2I4LsYjqSeM768e
K5vRLr0oQ8UOEVV1fswKwPZKszN0E2TeuBlbIjzjPwDV5dJfXNsThZEW/DgoeRWH0WcuQHF7o8YY
98/uNXSKQpRBMKUMR1ivKAeGk0OQtKnLQxTyNGt64ZNxXRvLyuL5rhrLwCK2ttqdXLRWo189LMvp
x1yGFLIFJ4DK+EMI7SY+VxjGIHiTSr2887VHU8vWdRgJC0ga2SS4mfuZnzoq/R2U4sIQiJfx/tJD
BUMGtQxSr0QOCX6VPV/Z6UzxGbO+9ZBvbKzp56pmuegJ75+qJgAXzKGANtrCDcahhCWzb4/pXQ+W
jmH05xasnwE/wKkCyc14wKdXrnaHfBfqvMdvmIBVfnCUuUzK/glcK2vwzkACDoyPt+IpTZ5W1BUy
oMrDVX1Ew8B8Ohn2e93O+wWpIgaXfKUGzbeaEabjCVI3RRKd2WRwBgE9cnduCm2YoNqknyUm4VQE
tHgCT3/U4x9hXNGN2wLFIBGcx65FuwI5ZnDiY80kD0no5GTeFdKjNcZvFMN6DSDYo2AhYgtQUWrr
C99AdZ3NINaCQe8I7YQxrDIGAxjSYQPmeNJdQgnoesEVE9MsZGlLyd5GHpUUU59mqBfeRtxFFHn+
kTIKCu4oUKzgTG9RRbStxiw8tkRqobnHo1hVmFYMz2FvsnDGfMd1iXTG1TcT8zck06A09BbGlw6V
zyGB/X+lEZcIzZ1JVaY/6GKgSw39dWbuhgdmuPwo+foeteWmqL3KO1NMMULvem5b+6iK8Oc6gu5V
OQrlFZqHv0rkVyXSU4M3aCsg4at2GGrDtmkewZ6Y+gnq/M92khWSyu7aZozA1RCDPJmiDz+eDgNP
SK3g/1aInv/sqOKaeylWxFbgoDcLYRhmpXYuKzyiRo0UdoyfG0Ok98oqBhF7DkdaYVugTRGB+hoN
u1B+h+8NfH26x8qZBQBwH0bctpNTpf9t6NtxB4Vjrz7PkR2Lr7OGhvRR0kzEq+9AqC9fpFPu7eL2
QwaLzdH9sGtzeka+EnOB72A/MA8X5jgwvAxH3k4fArHL7sp6+tgZPyAAqg8KUq1GMT+W0Pmms5zq
n/NLpBG9jEaCa5U3b9PbIgXdO9iixzqILdbI9BQLXw/0RgZE8r49Hw/WAa2aqxpsKBjGWjfEAp4a
0d9uoG7YbTFqFoWgXZQfW7E0W/WXxidCSNLmPd8bBAp3/KBuFCFnw4OeOmz2nmxAfOKWuJJWPbfD
GjVnxa86P283V4oqhy+PQtQQpw4NPJuhALGJRFlbzHvK87qhoT0M3OfVwBHxvIg4QwqfRMfYiWPy
HI3F67Y/kVyU3eXHOWfUHj1DU6UtoKYYiq8W1jxQsNOxKcDq4C2mWqIWABswJjDUHQQq0vZdk1ks
sHdml1rS/G/TggQ6Z5uxpsqpLjbRy7PyCY3tAxRzoe6XjgCcl0UtQSt+Lvz0+H+D0oQU4wmDzJ/7
5MUyFdJ5rZzHs65GpnGU+1FltpU6+mvr52bw7pPahdgjBhgAqkQzVohn5k+iNfHoKcWxDC6/QFGN
bm95yme/7olBoU1Z+khxLPH2oa1DhjgDTdh4M3qhcluzkDvynZ0iZOIUFN8heQWjMpH4sppaWXD1
sD16gZhdmylJozSYSOSFgXkslqryVmwqZwWhUch7xtBcVwdCI4Mb6KHwtR2pJ8VQARZToLwI2jy7
B2JYaN6Urbmb/sY0CpJqWHXmq7j6lK+Qv5Lw2jj9BSiU8P2j6f2ho6w9yxOj8SAn/MWohyopKZkI
2mg/AigwpW+qPisf3s93nP7zP8X4VupcQl5QyYWHBxwkA7JxqBtArXknZxBu814xbGOv7eWEGlsj
3Cme00TOW5SKuh8WRdqIJo/l01L2yxkgUEnqjPKFpwAezaUPkTJFGTqg/d8gPsV6u2KJeGKfB5/p
hkyS03siUJkd4yOSa6+1gyZE/6M0ZpIZ2B7caJoVtWwAkc++1STFFD0Loz8pTUq3NJb/KYYSPIUD
ursM6TdRRRiyzQUbB49iuGyjwj4XZrj6FT3sFv2MkZCrtFzw18aM5d8awfdpnuZkDEbx4Hkhqoc0
8C4DKf3yhd5cHdM0WqzpWc3D+pDv+AAm8MOoDnfO8R0CqUx2icXvnfSWPuuld8iBB7vDOdt6ZAex
MAP/rd3BHty+C0QmNr3+PZPC+ouThqBzxvMq5ev0RJYUIGyCT/YNOKS5v3GuEc9ENVbej+F3IdKw
7OYrCAwr34IrSBda4AZVeogO6IHcQsOqSrPSV+cHS5VbCsGn3mblLafYDIJb0c73yjSci1ekuvqy
K87Ay3YpRHfbrlNyyZcEZfXgoM07M7dNpJ9dIgdpaf+0B7Egg7ndyRYKV9L8fWwPjZPi1zRh6yHl
W8mNkkSfz22k2rZYYuE4DpQAcKWoekUr6pFLc32ThhMc8mOooWt6USqOq6i5EufvHSlLLfIoWY4x
rgtFotETqa4ZciN+yvBarv8vin+ZZjSaVwtTWWk1WtMpJkqCr0lD5GYRMGQQXDuB5bAC4dyt+hf8
fRgGGM1RBoZ2KFp/Vf3btuLuZeQIVBSeKKxEEdsul/E+uYkEEXfsnmsO+a9ACvPl37vHkreLvF+z
th39brc/TeGsCMU1mqaPN+7X3eeWdcubRHfmlBusyOKiBwxdsmytBopkbMhHrIOJ1OClHrCZAd8E
fwLNftsIYsvT/bf5TsfWZ5aF3w/tgNeXQr+vbu4lX/AovL5AHXHTE/VD6gusPs4KbsWRcyarC44e
5p1XKqLPsRErKNlUmCG8Zz/yxve4fVaLPVTcWXA84fC5Ip132nT8ABYSNG9zWdAmbEJGDaMxM9w/
U9IUrY6+ne8iK6keX8Ck+rnKzneJGsohOAvsRDZfLkPLsLxsywarLU4F95HoZUiCsq7s4CuAHa6W
c5hQZ+vsCFMVs8rOf2vrDeSMm5Gk4mKnwpdzOpcAkmVeZJ+PS+91iTFULjcVQgRYCMfurH7EEvxU
yDqPpvhS6uLtXXo5mkM9Z6bzV4CGOLv3c3F+dEqDSDqGkzxwHN6whuT3YF2TQgrmvuV1cvrK9I1x
xqGkKeArGUxRXPpRfUu0/dtXJvW1F4E35e9ZBwxtrzY/sPRgR4wKT4Cqf9XPW3Oc27ToRk1C+ChQ
2H0B/+FQWCl4jXFCo5jNayzIpiLppSfSPgP3vr9dRj5JxYf7BNLxD308NqIJlxt8HPpT/OC/ABRu
Trru3Fj3mLtJBuzlvW2eJ4yzYZgOZEVN6tvDheRGGZK54suxz51Uia2hDBTcaHKKrkODLoLc2GRD
FokaGoAlTcQH7a6dHwRllNj8z9tREq8WVmXxS9xlviF+fCykyzwXQOGfYgxjeC7nOlVpD5KBkLCj
aYQGjGmtuIYUSHFDYyQVVD0BXDoRjVtnTW50Nu1NLVI+a4hzA2OKw+em/V7YfgtzC4FUPSbPzDFQ
SOim+/7d6bRGuW9zPUG2nqycu+ouLrM9lVhhoIQy7tfjv1eStwdi0RZYJeMccWstRsFxS7ouUlV+
j+iB3EeSrbQ5ztg2rBlp8tcSq4Qz9lfAaOrD1rjEqadGS/eb1faVRNnFRoLwJpe66se3Pj+w7W5r
oy91/m+FrNnsT0bkdHkBBl6cj561tL1/Lf0kHllgiEYtIzIyvAmUXbwvNm+Fcp+VUw3QLShAo9vb
ubRbWZlLKiLH0jAL0F5DFigsTRAgqL98L0ZnmW5TUYJgtkLwLP73zMjef89BNZ3dGa3xItlUKnNT
jRcZO8EdYEIwwV5iPCPw1ZbzKwqkYI3buEEmQBfizUVVe+b53//ttWJ5u22AcXFXt7AnU2M76Ogj
c09u4WvsxcI/FCJ2hXbZFev3QzvgEzMItZbM7gCnnnnDzwiglywED0R1G7Gn/qwqSP0ek2yc42gW
TFgDbcJ3d3kfdgyqC+UQscd2syg7TGGZjy4HboHhcWn8/mAJbw37ZPxfoVXYmO2S1ijsROS/6PAN
gsDN15Xrwwao7bvDiqOwCNYlOXm1ifu+QZNM/SJ6Qcs5wzycXZLFIAECOJ/RV+cYAJjVZbehPieK
+XJuLdcFRAKcpwFmibKLjkrVaQFj/A2TqEpGCdur47/Z5vwbQkEQjznpea/t6HYtZ9CMCEixftjz
IpGfNypGPS4AcMQ86BVhD6cwb+SLi/xpNRbDiHGUaCqWxzg9SlMxl51Bq+a3i/0LxxLToc/yObF8
T+8P7guBZQaeWVP66NNzmI0/iL8d0vfIdlvgq+/UMbXaPhfRGcvwo3m3wxf5e4pXwMtS+0I1wkep
jNOdtMs3JN5DB86DjC+/gQyRTU77rvh43OipPRf2jCjHNtRO0b/M+J611ksrfsInsM3/fNDUOPD4
u1uxODLiCYLyWTUJ+0koKb+KzWsIE0kd8hYUP+DPMayhQsVXpqOvAfYuPEZU98iRDrwnAYdIsIFf
+Apf8IZalnvWcDr1FBKK5iQngW3mrfdwgyVzkct8Vo7snWFmtrD2gzmue+ZDr/BcYC7rzNm1QuVr
wJyv5RVUZppeoZzeFiknqE7U1Fe7cz3p4eGcKkimoVqC7lLLeaC4+eP3GRTDUJzMkGSXroRihSYx
eIbPLeXf27BoR0jQ4MTW+EzqhXaHryD4WZUji8L4AHcADMIiKSH5mgBtbp5HvszKs3DsGFDOL8a7
6C4D9cN8GyL6+JEkm8+RpYRex3IUKfYBvVI6QBrGYw2ew5Qc0EGBBJdqBD/5KuUEQwn2O0t61YMc
5Xsr6Lra1yssUoidlkhRGCT9ZpCy6Pvezm5HzR99eQ+qo1Q4WcIc3n35ADhdGjYw9aBYOXXY80cO
a01zkBfKVc/ZzlK5UfZuCn/374p6HD9E6qZ3CLH5hWZSwyJofIDBm70NiDXQ//viW6sH1JFHYiMV
wPxNYC3D9F0zhR9mqH2wkGwQh/dsYxsgzANvz6bgRUw/ERAuYbaPTakDbFy4plbadeevTG64N96J
Yu+rqszSjFrEik7KVKHef/DiIHwZPrd2gzxQXFHlw6+i+Crrig65jTPK7Inx7q/CAe6WjMOPAoN4
4mauQNbt2hg5M+jOgDU0RgsjkdJ7FS5HFJveGvrnVYyPkM23+VYSiqo3lUmHyM/FDrtJhCdnexuR
9Y1eZT0Kj5YZC8vwp+s9Y3N/ax6BJyZNkjP8K48JjnpgLkBjSJI/Addl0RI3aOhpZswevTG6g7Ym
/N2pL9EwJ8NP3KmW2ShHl1IeG83xNcn/StHm2Ww04IhqQO5WdK/EWQz2/RM6cxCpnaRVs+vAvZHK
aYAmuMidc4JfqFKY9yq9HDd8FAHghjmqEfkPhfGAQTNsGTJOr8eepv0CfttQBRWk1c/+7B8pFNxI
g+d/B/FcVGiCJ6b3BuXXhHwGdi/rqU/r7xrWOtQ6rpC/I8i8wf0cnZlqHFv9ev+NyfEnhwx7gTAk
jdWZIo9K6Cmowu+F3YAqbGuKw1W43qULC8gC/X/LN/JPSzMLeCA/ejWpYRz+JJBgsT9tYOv4EbCN
mbxXgpi/aa7aRW2bJRSBjHAXkqLOn3hp480Ugmui6cGC1RTypUdMH1lnYcUPVfU9Ornp2+cD8xJ1
t1bEacz0bh2bBFOiF6fARW8C93bhPZojfcWeEnmUKqTxPSmRHdxlfDFx7nRNWBZLz+VRPgrA/9+S
B6yA1Vbe5Fa3GYGFTSrjs0fnEGt7FPczbtPC5BA0TCA4D4Yw2xMxOj8nwmDwgHSkZKMftqWwH9hC
+cLMMYhAfPgEvZgER4mNnUu516yrm9YL4UHQ2JrCqxfnFUN89qrb0xGgQoFtZfedQDf//6ZqHOZ/
f68tVg5UDncdrhOfQWKgX+aRYp0rs7d2L0olQYMCgBTnjAocwKtk2iML5M8WVV7N/Jg1Uobr6wpS
no3DB7O00dIK641Zw0RAXUZtJTA8zzn7RUu+tMOP9JI39apyWcWcPBK4SseymShMYqj3FYuiz07A
hUBIOynQpGFQkKPUPD6DfJsZelmddq1yJLrDtTR8KtppAKBlAxsJBcSUYNevQM/soRtBEkXjxjkp
qmG8dQLsvCWDPm743jyvlwril+LDfVaA2wy2EiPGl5xM4FI4vIimS67vjfq74kcG/0HH2H/5kl5A
iX6Ryly2k0IBfPbAvNLpW3vvLsS/UgwIilGzs9ZCDmuO4XJsIwoJmCkLDLwaFXE8vv1ltUQjv7M+
TqgTOGTVM7XY0fq9t7BhUNajC/VMV8y+w3Dx0XeDTohTdMXsNXF5GqKu0SCWb7bhu+eh219PDd59
EHBfoNLw2GWC+cRrurCcIvso2fTegqri5hrVPDc5FVJ9F8vnQIpwB+7iq/R/+JkJiLHFEWUgT+Gz
njKQCKjGZiBqikwnBkFQM8bebg0LJaSa+2fnVJiXaCw9TorUBfAFboDwofS6S5xyvMuYlBE6ZwLH
VrBFf5UFDUrM3pcMoIhf5nVEYV3a0GYUHP2jWdHfxXe92o9GrnDJNzb5NfZoicafjcm6DcxMM0aX
MjHa8oREtbgtbcJIOAs1BMhOXZHEKNJJvBvi23nHY8UAEeOs4XLRie3ukqsWZaNQnOz7RsO1nrug
qXADlgebm10dZKIR7HBwEUxN4GE/ZpJTR5DYPFoOx9XRbz3q/LswuJvLcqQ6vT/M8HMytEPxtxvp
QNCqtKvdUyUYv7DSn06hmC9hI3sqFUYy22tIxdMzNwG2Uv9+AfdobhEU6TULyjsk3T6JtmM46oyS
+6U1mYZPeRbEJexxpPkOdHHLIXwrN752THSTwIRf5Eg/RiDqbaJGGxvu+3kCaqG1pTqIPgnkBPUG
8nejxWJsZvI+J9uT9R0JgqQ0r7aUExFqV87hUy0M9rFyEGpLM3MZTsE/K+STh9r1uaA4N1RegErO
BKQfut/qZfiHtdsRSkXIDbMavM0yECTzL1KOSOlbxAXbu5if8lhCXxi2DOREZr1rzpE5824Fyjb6
QFg8s3huHnvlDSc0dNSPhKSE8UZPw7dPF6hvqPfxJvFmGwuMnnpvJc0UcR7lCIth/WfPx0amj3Nf
CxS7YZ5p/6/It6RVaNTmF4UkoE/kH59KHia/VKVxz44y5aG+nGyClq0nL73lp2UpSTuGrf52z+qY
/paWlwJ5fXOdEInP4Y2BquK/oPZ4pV8fuIXwKa9OU2hN9+kfseVnfb+6XmHXRm+eiWqg/8OS55Eq
yyK2Mxot4ekp3kKDKtR2jivr1HrCi68sv8A6ih4louCmF8X9BY1jeUJ3pQn/uCoW/Cgg7K+lyxZA
o3d58liPXK2u8zf7bicpy7EuhsJkXvQ0xff4Ap4yc4Ljj6FptYSY2+oBK5kQWMovGWF5M+6rTTm5
YCVXJOB3cdz1oK1FbsbJhtei8DKR8sfKZjpClbGeDjgV/xowqcXWI7g//eOQW28Nu+Laecz/KtTL
KS6MYi0TKq95YoPllNR9z/tv0LLGz8oCellPuaUAEwuzPxnXl+GIBRVgCAm9QHgYC2CFwc0C2gGz
5EKAF7fiXl42qeViP6JKikRKq8RDFHSDXKcdTMQnAfxZopsnFQ6A5DbV1jaaYxponFFw7ySUBs0M
xxzaQAWRg5DwnKSEFj7rmyTwskI3whW54X4Ud3sfj2ga+jDYFKxhMWY4kytgIJ0AgUMEt4vMpC84
nLtWfW2ecg4cvLGtDBH3RD+vHkzj6/TojZnCm/cga7T68lY48M6Wt812V6vNXLJLKxXsg38b0f11
JaIvzRX99r/5fMF+V66+eNXSYRWYI2PnszXmee+hr0cFH1FH4q/FmAe2XIkLQFguNRC0Ka1g7zwy
E7rC5fYKsmieliUMZeOe/e9ORFg+jsg/QFh/N5+xYxFur0SiaUaLvw92UKtd1uvKiUp2Zj2viPbd
dmVwZQaz1V1zo66VG7lZMF7ICHjHvEFKLlT3cm77T0L4Y0a3Gs/4p9gTrnQRd6um0GnlCO5i9CyD
wy8o2lCozzM7nrUsuS1Zy+TfKfQdiUXFlNT9ixLH3IWhsQH6jFkZH0lu0jfwJ+3bz11cehZQFcZw
MNHgv4QD7GMtzKkAk1XFQ2+USG50Udr93+CV4CsaIx4CT7W0IwxRtAMO/ZWa3UKSy9+2KcaPgYUG
v6NdADhxr2ETIqpgLYCxl/9dadvbjqjyNK6ZFLOMbZDwfxJxf4LhfJ6VpOhi02YDbpJtXdMeW46i
KdKJVaAc3BoiQOi/TtLn58MHlpM45IWP6hWwsny192hsTfrZA8wDUBeZEhF0YVvuHpfJS3InFFbp
YlH/oCGY/qGKLHWpYF1oisughVpQoE/bOGL+e+cgE57eqTXJIhxHmk6iSJwI1ZuqMRrttE9JN0yL
k34cQcj3guzw+doZrMlY0Pr9+6qXjV6dqSItMdnefHeK4Djvf9LA+LjyeFWFBGWVkLa2suQnCN8n
Ao8Oo33uc2V5bYkNoQKde6YOOeDOyrw33ZYH33uAuZJ5sHX1uS+Q26Zs45hb3FS0GlSDVoqJ1/zD
KzFabLwGZLGVVUP+22JZkDV22UTv6JxgyiSRIbPCjDpVS7cYlStLlnIW2uzdcVyZtFCwDzrI8Rjj
ynt/R0mnfk7l0F3H2Ila/w83A4vsHGFCJNwVelRPxljmYNkTMIRQUAE4ZiRxbCYCs8qn+rCpKpXd
veG54kNjsuwT4pF4K/W39wVIB6nvYcXSjt8iFRAsg4N+q6cLSyXtWzzi/xcngOO+Wfd94YbJZEhZ
Dtv+Q03fkH10A02pHeFgSFSHubGNua/sf6vss4tVrokghZVvaLto2Y1/V86SC1N5EMCfOKwDdRu4
4TE+26QsXXtV0EAeLTa3UlAAqpMluDWdP7R6iDTxX0K5ld6y8aukvIydNSutXXWCf1jLgyweNGmR
N/qbGJs1Fsg/JwsX8URhUKIO1sTug+hrZnKeKBPVBHGv/y1dK6J5QjRhTzPONuv3hRdJJfdaYYQF
yMS9zDxsVjsFBhUNTUt+ZM+fpz3/b/My/5RaV6yvkKdLlQJgH0hoMpLw2dRlGl8TBUcM7LKE2/eS
mDEEPQUl0VTKj1s7XIzCuMyoQZoDoGJaLuqvz1pQt6IJTwOvV3byA+CVfRauLLoCA/xIvdDyiwh3
alsjbOMMG67xUmIF0mrWKYTTlZx9WhKb7Edz5T/AWO0Dd8Vx0XD3OG2p55Gu6ZErTN59krRsQyCr
/KdPki07w9Ry1+n1gRowEYDa0Qa7p+6ur+odjQKqKpBd38JQ9on8tbfI1NYoc3G+DjKl3JiQNQ1j
3mZW9OE2Hu7YiPvY9O7OzWdgtFbLXFlDftCFnDMVLOjIduZl7RyKTnYptJce5aoUdo1sDlNOoGS1
2F/EJmC0SkYorTZjvGPKYRX4crY0MlHOUonh8swJT7+I/3xg5QLugXfd1dXETVZ3y472wrUs/jkB
s4TTZGN2GPhlzvEgSxBYOpDSeZsOUupruA7jdQqx+1khDAbrQFyXGrdAlSxfTdFDwxi7BtBsKNCj
dq3WyzqqGmZ/gvVcTXOlSCSNaGVx6blL8vKsASZfcMEqNrvHezvjqQGv24p1Nj+iRlPHVk3vgQxh
dPgFRmaXlBH9YFd+yTohgSeaa5KYKn+MpmzlxhNVdONaK5wjKg7gf9K/BE2d4cCQtYdwtoxVHFj/
EQOImTz1GVVkypoNpNq//MEVXuBN3WxNyJ8IqZKhdNeBpH/XUIoBkOjuf3yzJZlhQ1VUxILV+bew
eOMI1AgJCbQqb2ZmF2rO+7SgTa8uj9E412pQ425nr3zBrMrc+DNUCxgHIg896qniPhXTOY4L58j6
GPSuatFUiwZvVmJ3f2YdS2Dl/x0wNy3KN0Yw7vrE5Q1fxtcK+Dh5+iFm7gjp2ACOKpQBln+MJsHI
zSILcm6TGNvb3VYN2a25cXR8a6XC58cQw5s3FnpomgS9M2daz/TilvefYggrY2muM1csWqDrj6pe
GWgVt4PSPB7TkhRVwBKGTJLe0XzF6JFLMGQgcOXFXbmLxSGh33gFoSCGExZC+i7J/r6EcBbvni2Z
TkTotVT60RV2b/T6hlHfxWweGw5I/WfpNtOY9OYTfyPbT4wK38RGScFrsRsw3nrIsh1gqJOJHAoi
q1ZCDP8awrdPLGZkzfWeBruTWXhPVK2902KwKKV3Qkj+0NXCLB42YuOk4N173KEvKHj/C//dOi1N
FcFeRfXDxqDCz4erRsp9BCR0zYIb8F/gdMLw4tDtBRHilkSP/WExAkUpOdl1ZEXcT0GbH2+mrL4e
Zu66+BSsyuSdSZahMNraWLSwSZLhnqI1tMXQDTbRq7wsscxk7vmJ83a2tP+nsoS9zVh2DWM6SE8R
qCpbO0S2/T8b0iMV71QnfcCMSS+cqgA4ZGOXYLecUvQxCPSJUytrHQp1zjU7W/5t+3IreHS2jX+7
IaOy21gQ8iuPt8ktbyveqVNwyH2KFIabGPnmXxKButrSHrCTMZ+6LgqZZujmGUEY0A9uSW+9cQLk
xcFu+MbSnWqE+c0mN/SXvuNQMBb6oO0o4x2RP/eau8RYop1gX/Ko4VX89n2B24BxyZdSfDrt5Lfd
lcaV01AqooD/fXxhBLP+Vqw5t1IlKw4GkvpqfUgK5c2nqkTjZY11SyErfmpfNflxeYvCE5bmS7gS
8lidUtmSW+nfTQMztgDhHi7XJN8VYgoCJKKjnjO3FkQE+OY1vAL1lNpVwXHyYWghyAVo+djWSLwv
H6YU/4DqdOxUuSpE5FThU3YCc/XhWq424mmNblMOoKItjIr7S2MvTITW56EqhcRNcy/Fzkim4bec
pCMzYkRJn4HlFDq8wYqqoXNmCF59ARL2Boq9V6nSZtxhtUMtCa61WLzvy5rYDhmpByxeKaiEDUgs
4pViRKpmK54yR6O/sak5xnCx609+6BCtyK2E49T4+xQq+gqOjswiLULGPCFFsF7mxJ0/I2QlZMhg
L9WJrclFitXCI9cXOirV2/glavpkSBDU9BTMJ0q8SgBK0iwwF0+M2n8QpDRDaqM3lEbNysGGoS61
AzlOvqGIgEKrX4FY6AF79kwylba8Dc3j6+WzTSKOai86y9vwqLxogekS471Tlj2mEmM4RMNvt8Q3
pigZX38te28qFJdeXBMjwg2vl3iwwQeh9I4z+9jCvI/WbduENOzCy36JO8Mpeu0b8CawSUmOc0m7
t+al+wm+uI1NVS+GxDDU+pvSTnjDqfPplU+qQDewf/dYxzYQEd0EymrJ+j3GcWcc5NWoYtI0obdo
OEdGd8jVxot5AL/v8rfUXI1enDZ4sxHsM2TWeZh50HiRjm7oX5QCWTnl7JmpGMPU365RM04kKrTO
96kvV0aFfCBJ8miCRB2RBEuiaeobHlhFyF+/6nPlALgY5XKCGTqG0r7fmwTGONWuMR/MIk6dHc9W
MAPZnASxp2JCu0ehz9RyhOOmuuiJ0NopCL+g9fHHgS81oXGxjZx8UnAQn/cS5qqy6YAatlmi5uth
ONVbK2iZ1js5AYtYRxW1qg9xI1HWZ07QEEd45syp6ZYK7JmcKWRA300RRd8eJVV9fd1pcZiHDkk4
q0+o2srercHFiEfgSEfgtZXneaLVxHMaWtQC96wDdnO2Eq3QL5YvgyZFmEf6NeXNd/PihrfifCzb
tviQnysGRAAq78TO73IkFiDWfGdcrMAzHw04DKgFRWqLs5CoCWQOqECLI4fXHi6sAnnxdOwwPn8R
WqIgxEzzPGsr8kQTKn2pVA0iCX4fMR45dLOguHONV5/u/NgI+wgR26G3uVtc9CVXRB6o/TM/jos1
ld6/umeOK+f8rjAjQy1pppIyX7AUDSJPhGISyI5q1VgkrX5nqOWO1m2fYwIe8hmafR2bYO1xXJHl
KZQH8O02GXrenijNhYKiiDvc1SOUtQvgwLt75ZqS3sjoL11P/dti4hahfH2U5DU68qjxgGLWm0R3
/xirYJcZwnka1t2Fa1k8JHmBoOQXL+Tnica/86Ah+iksFmxOXRlBeb+rSmV6EZl2FWSsrfd7mgBC
xXzr5bU/i5hO2+4jk91KpPGALoMLiCALQeeYpEyFN98bF2rV+3HM1ms+uwA+sNR+I0sHKJysFEo/
qUs159bavKoVQRvF1QSldHhKRvNJjccsRXAGY/+s+AKIxVWxCqFHNxUK3cQa3t0kiZWGTizBJnrF
HzesY08nmmPuraNosq/SU1rNLOw9ZfagXBipzSL1z7UsskL4DIHyH5Sh10uLBIknBeMV6AJdn6T1
MxDXvSIJqIzxd5rcqPd6lpjv7sl9eDx0DSQYtj7JMLGp+97AD60MyIaAOmH5BuplYsdkhMiQHlFl
tA4WCfUw0zOtoGK9KHkiMR8gZwwM+bv0bqkxwlWUbCZ0bAykFZJcEiKAgxSqHOP80KBwITHbNsEK
KBATN/cB7a4PNoxLZ2RixyqTfx+v0x7XMOngh71goenZiA4eWnm9sSsOy17LAmBCJXfTIew7hL5e
qvW/ePhgNxgOe8sqSMkTywoEhmaN6Htzu+HE/ysM1Ny5FHmpWuHnzhJQ5WVNMhCleCqSXf1SWhOa
SH4GLJQ6aVfLBmnbsbcxxHz8uKHnraGKjkn2wE16JIvo43pc1P0KfAYw+s0nFyt9vwJBhauggvt3
W0oc7BcPM69mljvqy6ZzWEoDQ+YnGlnLmtZPpEN7EgyJLpp9JFcs2otKHVFITSazHoZHzpE+A7nU
7li4N0SoKkxz8dGyZUPcZliq6xd5qV4gAWYLikicRUn6wAHP+bBQZGjcavjQUdYHTM3EhIYAe9+P
7JbTkKuaZf7VHDRUWHvn6GSlKSWe1x3Cl065oKbgsGz4cwx5tvMS+dJCkYVwBgvm0zKPqbzqd0EQ
V/J5tOHz5M77T+18gXqsfZz4bVfTJ0tZdr57gpjhjRcsJpVMt3soEZhiTTFDBOhBg5X+Hme8bvVq
wDV3KPAIixJbgOZ7QW4qIJ/XpYlGyctRI7rR8JwgBImgl1x9uxf4stc6QYNl/V1OD0uRHY5ZDPEp
LVOKTHAsgKYTTp64PovjWheijDkRzTZyW2LFRRRyK/JjosUEwiuiBjFraadpwxRN81SFX8qxYtey
VwOWmCHwXBC20N7i0Y54ni52jxGMJI2o9MbbULXlfBgzMHjzk4IyCLRuc0wuVv23qMsGOHTdU4qS
xUtkNmr+R51KCFyPhiASx9E+V8NWs473bNagMRHya5C8DdOJ6KjoKq5mlax85gDH75eM2j2dELeE
YejN5zLMnNELP+FAaaL8ssf+bZFtV5zKYrOcNnCNAXqkkwBHf1pl6nzAhnM/KcaOXPRKV8NeszIt
ti2fAsXcD8RVG9FaKtbOwMO7vb8+zWExu+aOAO4+pNzuaUOFlbKERhrHAGKKvIxsA2299K2yEQKS
JLl9uY7DU05g/R2nH2GjRbYltF6HbksO2W3iQhEKM2h3pBQRJD3SjCfCFjtJagX3bwehCzcr6rth
qTBOy5P0TJiopXPK5K4psnK1wZMmyok0zBM6Ks1ZoSA40FlKG4BMKfYx2tcjYNwN4VIBaGvML4qa
06F3XPSCizEPTAGMjEkzEZUGmHQL6AOB4gFtgLl+MPBDVfPG8eCZdzJPp6Egdcoqu608FfO8DCYZ
ZW0JrfyFA1vKu1VmNLrhC2+TTI6tMD6EzikcUGGZ3SiJ+jhMF/tNBSld/jXgcCW3hbI0LuQ14DNM
L/xBlm/G3mBOdjtUlAQJTAVNMf4Ou+Ryv/G+NVYyRks/J2vtGCYqE3e9Wh+1LjKzIhgUPFcFA8mg
Q1I1hYeCw8Gf/mNQcysfqL1eb1fTI9PFRx0plebtDfG65UwnPUAghrCtcSsId7YNJgBJcXvkU3sc
vF1nlZs4b2vTEtKIUptHRmgrOMCQc0gWHlvE8dFvDvEk1NbY7+kRxuLnoes/PUvlDF8WnwGq7pMH
Q097vm4P9BQ41pT8OknxFBWWgAI0p5E5j8NxkhFotskZy/Mxsm2Gwe8Yz4dJaKJGuGTYfbbg7V6y
GykkEYrE8AmYf8RDQmmNoeNNFLmqbwWcAcY4U2rB2hQPh7esL9Xyh7fe6osETVw+FpF9Dri/YzBg
AOs3A/EQgUsUVvbLW3DHekFpCqxiMLnVuXJMOu7MS0C+S7meOlT4o5ZmSqzafrYSLJNCmWBOvU2S
gdKs5L+wTNyVvN3ZvXRfm+JvVDE4gJWbfSW1WJBY+pugWIaBP1hVWlQJTWeywOsOl4FOnQ6gzkpt
t7CUc3GwLbCMLkKmhkiAk/foMUpCxk3stmYMryi9j7oPIT0Tv4gFZf7rFL+wOHXyvyiINbckRcAm
yBCIO9voNtrBQJgXjmbAgzlD8Qn3eaq4YS6c5Lvc76356OOcuXmasgVN6LcD0zGxXF6KalyPactx
NtCjfJpJPljDXA/cBtcm45I8fTlsojDqFROevP+YbISijCoHtCpeCZEg88XktOdPL3NfXCqtoxqO
AuRvoO6UINCWmIdyaIgLj64TLk3+J2U9L2NOwWh/qYtdBq8Jgb2/sfe5bboJA6YrfpQIaCXdHVWn
pbSqDuSNU2nC+39/N0Kdm9Jhg9KwT5StJC82PbY+1R/AQcrs49ZQorKNQ3jifR/LP4J/4BXKZ29V
BQ/TivEyr5E8EC6B0nBoMyxJfKzdlt0Vji4WUiNQc79g0LI87EQQI1MHNdEFOO9WSTGYIOs2NxuP
PlwYlCd5PdMAPRyqemPEziC2hlQxhp/a3XKH0mZql1EIabtc++axRF/eM0wMyVbcGOwA/UZsMS1+
vlAu7EeNDkDPNnxsWySXaqz8qJXhF5zHIiWpo1xhalMaZUNI5RCF5slKP7PBvhwPeGJYzOeoilLf
kNgJ9sSp2IWIcuu40jn7z41nmJFZ6XFRDvQry2vvZVv9Ohn07TP2JQ+ha3DZsqNu2WtVbDToJODX
pW32S2xLGgZtSco9nvKW9hRN09MFjgWSqk/P/c2slVzBK+9hcXPuU0NuwLivLGoZ2QTIqRwcQOD7
L+TC7iDil3OJL6giaPFTF4sbStCCLkeVS7NA9MH9T8cMtVf7uRdBngPSmG+4bhvfLEM8+XRP6XKq
Y0qibl9CP4Td4p44/Sq58YK2Z09CBFilk1+sEXoWtoFbdVvrxBjXkCQi1xerPkwcWN/+lVr2QT8G
P21SCpEWcB9ruBmR0kXU+yWBUNOxh+NEXGXvgF14n/002cNeFqZvZtbc0IiWniOizNHEjiId+JsI
qsV7zElLC8uhFJYkmBi0vvti+dtDC4dppxJ1hNmQ6xiWGi1aYNMaNTR8us37+X1YCPRSbISqRRhy
j4DRlnhg7EjSZRPilVEKnp8gpPlfkExDgTIARPoQAYYGwW13feNu9yvMvZMKLLNLZ2xBBGOiSylh
W7CpbwMdpabDYKee6BUf+4zOVEgmFRWY4JKWkWOsusgzQ90YsKLaVdFt2LxH4yETT3g/yc7WhXXU
GizqubTWcVTEmJBd9OzoRzbJmgtA1xasqSe2wby7XDlRH44J52pZ+ctm7nDDwpVZC2BXGX6HcSIe
FHco+fAgfyfnbguLUq4pP7RAPNVhWI5T4FXTVzaHRWQHHRmuQyKG0Tkngc7/sxcvbBaOabkIIZe4
xq/mGRxUYu7s/nf0WgyRHNLS2mWhQqDwcdkyGwWojq8NkeSdNl2NeHdu9KSX2gtK/gsvfzKKeNA0
7q8hpl5395+GUTQn6szS12mxg9TFYOmi5N1Nrda9lelz92HoC+yQge5lQmgvTOKQJ2qJ7gKN4MHb
l5+oat8mXHnQWyA2G+DQfCd3flrnLn3tDgczFgSnfkybgMnzEZeVuSCN9Oq5Xs7HkadqJRatptWW
lx6fpTOF01Ui1ZOJX8zF2TlWDtVr4fGZUglynqBSsZXTEUbh0+y6EjDp5wC6rg7OL3zMEmtyl8wN
9xHQWJrl1p8+KMKKWTlfsnKnozLB/o3NKAOiYx66UfG90Ao5Zg2xy75lf5XQiKWf9oAiyzA28GaQ
NcawEUPjkrkl8P7VQqN0P4HrgYtnLqIhdncjxwztwUhFr2+0eNUni/IUV8+OZkfVc9rRR5Tf5HFA
AxMOkyeiXcN8YL7xyzj2mK4tCabBnrMI/REiF6vTD8tCOLAnR8F99tJVQcr2lPptWwPccZr6CikB
KnBwT/FTTMNr8KkSD1uj0G8l2Ewco7PFQDmAtzqlQs+dLin/QMEHIijZw1UYwK2Jg+rXsQL3PSeA
vZ96BiAWaAyYM6QB6rMoFYNf2sPVs24jReUvZKpljto++AfadfyyUtohfv+ornN2sGWXJr3/6CKE
GzfHGXPyl0FdKnEv3r7MrgvvUp/jqt54yt884INF81wUJGdHiXvteTtn3HaOijcTOMQsPxyvIAo4
w51tz5lPKMDoNsZbr0r6KIJ7lvorO49nRIKT9hwjPHD3fmKc4Ufv273FSJHoZ/zJd21R6owvw6yj
Xv/5QfW8iLhASzYT0qH2KnMZnKing88/nBNlwTyJIl4fvkn3YtkKdBtqXkREaJnknXJ0iJGrhYm6
llNAaLEmwqrDiEYIRFspic80e8zDeMguMGGPK28dBeD6TRVpJlroQ24Crer3hrkRj1g8SZowzoEl
aSb31iO27vr4XUyVJfS4YhY3It2DI5iaWy9B0W3UkbHwMmSD5945A7LPwBuEPKQFHckPqmdJ7UtQ
UMXh0HLU2Hm9jrJ7cfu461F5P7JkhXj4JdOdor61wrMOmdL35ree+EESY8SClRojji8vzRhKsMNU
/IK5Oxk2DwNQNCI9pybywZh8+ofIqmqGmOPDUcQVuVePsZTqbyFHA5tLNEEs6sHMXx+Y2KcFThE1
p8e1bb3KjLVrfUo79nSwqlYG2JSeFf2DwrVHnoz97teL3IZ3Xnhqx6JHGO9oU+/2t9Sv7ZYQQBG0
0k4cM0Y8XkYtx6rXdDwLDUTy8ThbzDpg+m+LE0rVHSZqHwpI4PTweZEjZB3OcPqAvXYZ0rI+5Cc4
JrDFgC63DnhYjkTNRCicqP1iY7Y17krxSWA+EsvE9B6Yy8Kg8DKH+4sxshDJ5OMhFQ5j7Wm/mFF+
tQUuJXe6m4TgjDZvqiGhO/rUdmh2pDffLPXnjbqOWVaFNeiiUFpAKFk+Y+Pj9THtsxu/srEXjyAd
5J9UhUT/cuPJlm3cjbEPlRMlyLpxXB72J5j5nJ15C+p+0AGmHzKLQpqOeot70ML1dsJIpalPtGhx
HX5p0OfjygokFQfXPGF9o8HR1b2xOWPz+Dron+NJU5z24a9XZyXmNK3w4WU31rJ/ssnomv3urwcX
7LuAKafjhY7n1P8aVsSPUF7MGV3iAFDZSfquup1kzItDp0ews6YijzIOdtDfkMbErbEQnBJUlKi2
uUogoQZaZI/uAujTpZsBEToeSk+wzCe3PUF21sPozrSKZBig4fFmmJgUL1JX1f3UMv5JZi8NVEj7
cZNgMXunNPFOw2TzT2XUbxVreEDsiUFwm4Rb49UYG0VAoefQQ6YVxqTHtznSoB5xZgeMYkYbiL+w
0+ErviVo1bWgEhP88uJtMKTXJ0XsOA9DsOvjqky7z4JdAsSd2CbHIlpV52alTe3CCC+TVpHRWyb+
imuA4KLmAJgqrSyOa4gaFdovpm2qDoOk730V4a7kNMYlhfEqi6aVpxwmk/5T82N6Dy+rdbr+gBOF
GBdVDA1N8WZkwWlw0PNWHcdMFrWFF95lbR++7ISDBLyAvARG5NJWJz4c1bm1u4ipbex1gd204VGn
ohSAzDqeGufas13ianEXxkFkGiFXOodineC7OIp6qkrVgI5+vBKVKuWzSPvM4v9RPjcnOL1lvh8x
xDCeP7ihujrpNBXIsQYEWzUIX10KrnuXYQ7dEhy68Cj0g+o6QSuKCPjD0K8R6twGHyXsUw5XXR+u
T73DOmbT3F8b00p+LjGwe2WV3zDxLuH/3B/j2vFPM81AQjCQvRbx6xzK8djeQSj7CUQM55BT6GlX
v2RB5R35yhS2LPTHA+5176W/b5c5oQn+G1fU5jkC+AUqfBjIfX3/J+F0E8e/5HbthwwAPx3HOKOH
21NufFfGa1fNqTt66eulTLdHUZ6fQSGCERIgKYM86r5MCPP68MPPnKsaMuWXOw4qGrVl5vWjRpE1
rXI8arx+13A5qD6SJLtzPQmK947OCW5UNL97sKl9ekjfZccRO1oKvGqhJ26FQIn/aCDZA6FNpYyj
U7PQ3cbexMq/e5zAzHO9GVFm3kYXq4/nyQMfMzkDolb29EhwmPYytvMBGkITatTa3uRDR9f1BmbG
uIaPOKGkl9jboUPixnBjEivUK+0+Dkn77Xh5h6n8Qw4MDNwwQZp0sJYWLhv/NciiHEGhHGZ7Kdkx
cskf5wYTHBAQzi4DPPZfoE+K+V0g+0OZdNT7aRWE51s9ILNw1bjSUnYLkjNvUMEgbBjqfBtBB+k5
BvskVpQ20FE1Q8ghCCirQTshd1c8iyxuvs+Sx/fu1hyT6Cjl4uUE2PzEfxhxs4T4Uv7KZFuulPvj
lkWEcmkTDOqfZesmMyTnUXOzdgETDaFRZef7t89Oi/614h4T79T714h1KEVf+gvo0NtnTEzbKOq+
UpZpFHgeJ+v/1LWJMvKM0czGPDk/e6AzHsvjORNlC9gw3QyCL7jDa0EGZMsIsa5M2PzdZGe0cVI7
RLz3BRomKSW9gOGiFQPoaPcEk1t9IH+yuufoztg/lKccv/4Cz415kCNCnLkkwy80X6eRLlVcM2Yb
OJHT2TH2zyDVXmMVB1d5ddrjgj4hsq77Z8EKOhYGSD5WMiK0HSOWVB4gE4A5exNYAVr8Ln5sBu5C
LMcH/Yn/F3fG8wvEXXACLvM4bFgloTgrKhW3wAiSeixEHoj18Kst+E4z/2ItuSWMrFfWUpQfzxaX
LZ0OPy7w0fEFIH82WwxW50wOmAKWmfVrnC39Xkmx3XHwc5zJ1ear9U7L8UvFjfLTWOVX++yvfray
+ojobkWZVOxDzVVkF44nEMxSZQY4xiLNn9/GulCzgYlmsP2tVZJUS62L12vFC5FwSOVRpVxirULM
BEBnjNjNr88VyTJHA1wa0jrfwQQ7cib3cW91fkHvGKEvR9ymZ451MdGvAnsqfZUEQoxK57cKAog8
2vG382OjraOaP8l+n9J4SoppgqeFlsqsvZLNMCpDbW7aQIZXAFffoxo+EKuLHld3Xc2B9MvbNVAl
ilpx+jf/DH1fXoo+kcEw9CT79cZkbQ+oB1NbQEJpMHUClW8EEuYGNC1sfb5szB8O1ma9dZhXx/aV
78dHuw96qJFwvSmez5fNk288qq6jQ+vwHoV1OccQFjFutbXbogEH13VcBQail8NS0Uzmcqnpc8zG
3Wdc0HV18/zF2RKiKtINhIAJT46DAo2/Q/5I5gSRwu1xTCkQso5kZPB662OqDSgmNDyiBc3hTGeV
ezmgy3pFJU5g7gVdltzihV9GssAFhlcRckocF5NlG/c4lPkTJ5jiXLN2j4/tGPv857alHGF4Baht
EZIbgnXZWUtiXpwwQvgFOdyT53s9v5xVDArT6nfGUuQtUhdo74kqS4Vqvavb98YL+l0MYy7i9f45
kiuZnsCVjaVIe7dHLWP4wxli/6/SuziWpi2zjBDjcZuYSQt/jwlG0WOzNaufCSh1zWSlOw1gjypO
3AixIJat4/flYYxwR/1gtzY5I9aR/f6DFjNhX0Z682Kn5Dr8ZXBN81AAhm4erC/wGSyQ8HZlRryX
NZqSfWqTS4xdezOSxLKrxFgaHiGoWmrdbjraS0obLlljZkWzrnLvVQNX0IHwAGqmLzHLzQvAHwdZ
KZRmsIKvjl8nc03/r4ML0NmG73AGR8cpkfK2JtL3eYCk+Qj5D4hL+84bSs4Bmh+qK6ePF9VQt3Fp
ZFrXFFpUjhnCJh3Dv1JOOD0dRIhLoTbugP9//M+s13gh/b6JdA8McOO9URjK4EGMYTvgwR68PkeJ
sI5igzOu7BVelqHPmzWZgKy3kd2nMuP1lN4s68t9sCB+VxxMg+qPoYeAzLAgEDhIhpzxdKRCmRqC
pGYjstWiUaU4xwsOkKAYNBsCKd0lNwWwvYlirPIpRVKuU/vj6TKwe4sPF87r7LZD5WSWAB+bwaNP
DMu1NpcR7izN/NWg2DfHcR7AJHNHx3sbC1uXwMJkAvrwJ27Prw+RY67vwrG9nBY9NF1rVKZoG4YE
LAZfHXLoMLF1jgK25OyvCscy851OF1ufzUle5bqqWUBKy2XJ2a4dsvsOAoVTF9c55kjdXCDJAsSx
IVvC9JvJSm4/QKAB7M7l/ptQdFMiCIxL9cLwVdJbH0DUkFfM8wtyxtnyO9QnfFYj34R4QPyV7zrn
LtR/ekwr5gQQCkNfP40xEiRyurGpf705oGopululZDv6RKCLNDfYMq8Qm640qpnKvil4ylvJccXF
emv2OWEtKmk9JaD6g8MTeve2kPoqpDrThzPwtdKT0W1Ra0kq7claB75JRcDS9WfqFnbzEZNQv5BN
mczrnFtKSVF9D/Ngv6MMTq8e07wHDa8eDWcelk3XqzIsrfUE7MPkd3/xAcNh3ALVgm8gKCfCKea4
VrhCpng75LOev0XCFr6lOK5OLqZGlaJw2W7/QGFkA1wsWCjnGTyrTtocCdPmlEmEsNrhvgJJlXdT
ql4D7qGTyHHk1MTiFEKKNpeZCRKLCgeL5Gyjd6gVRIOnUewudd0VZ52GIUfyEkCCw6k4+ypQ1RdV
GkwESHKAEg7li3V3UyXcMSUzHWnTSgVmZ3763weZNuv1Vb4+TCvVT6LdBG/JPOCV/jZYMkHun8eX
T9yB0OY0Yqo9APJB/bto+4+u392dCMO541HLWvsT3voeUP6NhiE5gQOVCd85ZDOzxVPwCQIRpqka
9Qlc8ziOeRAqkaVVDy6m5EW6KQR1ZyffN0oU0bQrM8yPTFad6W5uxYH2KyuqxBRoKRZRuNMLhGUx
Hs+r8oqRqGhL4uCOgvySKHeYf0dj2X3xrdnM3zYkyd0Igm6JGRpFmcKE+5TnbQdZozn+HW+AeQ4T
+688JXhgFyu62fP5xiCoe0arVYKUEPQc90gl+d9b3+mGRHICqdk83iF12nRtNn/CfqxrpSFkG7Ut
xuNO+oEclw7WkvUHqbX7B3fiNb2q7NFnlByLmpxTXwYoImixsbyhz2celqgRgWpsw8pptkYNcYrg
KW4XzjgLKxIJEOB2EW5lNdEpdbEY7CLYYymg/+0MvTUY26DqwUlcl9Gq0q9Enw0k4N8cv5imzlzb
ro4SLw14guw2X9egafhEPBYFoJrr8peKUKVs/R5BRLLvTd4W85NcbXzPjC2cRQjSsnOWwEPUtiEB
w4cznZz52Jtkc54NaAPD1aho52eMIHE9co+hXBMZ5FgX7xdM3X2y1yjDZFaHVAcRP2ZArF92/o62
VrRY6iG2hmpwrWpGoHlibaUg3vpGaanjqVFahEeAiOtxXhfyxJktE1CMn/3K5Hd9wenzLQjuDHGV
F2/UFwhwBX7D8FYyowvGEIRFEYDSKYtYxy4MNpS26agcfhvP762ypmgza5sePEe+zAHf7hYYOaY5
0n6355DrZ2UBKLfFLAKb4yMUfr5WCxK+MIF+nU5s8ht1p/fS6hA4puZ2izBmtP+7nebD0uFfvX+5
y8290Fvbn+tm/jiy7Wz/Lbn7GWkTSnYEYy3OA7Zq2j4rF2F8I/7d0RhrXbdyeOj8Hr5LsLDjbMHB
31pixnuJSvfx+GAd9erHVgDBeBYUNNyG2YwFXo4FuKIhkEgE6RDPkr+wAanfkDY7uIDr3ar5vCIP
CZC58vEWr/zWKgfCRA9y3al1p1uUwA/AZQDPrH0E3F0TZYbACzXf/LCqNI6gCEb/v7OrW3TaKJ2F
6MUssJtC06woa3nxAiA9LxRjjIEg0whzHjY464lfZ598koOBC4yA7xHOMte2BrAPBstmZaqEqhPK
5Di831QXQLi3KM1Fj6KsJWZtR4I8j43gaNari+27je4QV/ObRCVL7UGpANI2M70U+eLe9m6V/ony
v2S8Lc0O1gyDfMLYeh16ZYODHqoji0OJfag8a+vO/LTldvZVYsxCNEOoN7fmEulH+t/vPkeFTxi5
Cl75RyHzFE6whNDrfzNAW4EcQJC/MPB3gS7ApciCmp3xZFMc3Rig+hlyg+20J7ikcAyMuhtm64N6
O0RV/4tVlNUG+M/ezFEgjONC4tiE2GnKJ956Q40tWa2jG1G+pfe/tPI2fgjBCGX+cmjhfnbYFBYE
LDz6RsidoQCPWoO/iekc3pQTWPNLIwEn2zb663QFIU2cXMwwezTxKborx2Z153Li2vTcsfBVqHNT
6ANcEG8r0Jl+lBF3+nIHhe223fieiUAe7Q9rjowQEIgLmLWi+z9GPARbpb15ErcBHbOVmlqoMgBj
c0LRFkNKgtuUNdP7J74AVwCs6UJTM9yfUtSMlqSlRXduh9aFrwv7zOg57nf5eQ/TbomXh9VX5Rxr
GosVXvdIdiR0JU79Osu2/pTH2UpQpZ2JURLhApPe8sIJglc6V3NmwePUlat3hvYMvVvUFfqJjoeL
VLaUcMttr17dvcKUKfEFmq/RBxommU06evOHpxYVS395NvQKSITkLF/d2xiTMuyybfgJwI/rB+9p
ecLPnz4Crq540UZj3Khb4DYs0ECZmxtNDIYexO3G8CpO/YNbA+n8BRNQuTdcdaDW/X+PLpp1t3IZ
/TWb5UtjMOaG9oHUMpzXpuVVXYbTK9VhVBoX6auoT64dvTAGel66eQoUTqk5qtE2WjEHCTqqMDIC
P3HTV7sd8D0lnPa1h1KxAEP1jJH7+03T1RY2GMDZmVE7csjPLiVuvGECYF+tDkfvozdMBQQbbeX0
Vo306/VBjGEOdg4U9SC4JpJnyzimJXnoqCsULxk79xcARo6XCqdojazrjLyStH+FCFCiirK3/lvR
DsKixMlLZ5CLGhfsOgKPxdSCI0vq/zWcgN86LZ82i1K1iQrs9hpCMRTty4PZkxmmEgkv7wPeRdmd
mu88qy/OEYUcHURF5U3GCPz74hwX+/yKldPYROIK74/abqIMNVJNfs0pvzDztkFgHTLuNAzAVeKp
Va5I9yOrd8bEjS2wfXdVCcTGWKV3E2J52WBWH7vs1TQ3vUFh7+Km01VWrpflSKrR7LMfoBPFMwlV
8zl++gKGz6rPqts/0QtyzShDwV4C4fskxdTqTEtIMHuo8WihoQn5NG5omHH6gxoPJlkMEZos7Cr1
mIJXgbdlIzkiGxHkU8leVeZTFDG24QBNsH0+g5tbkGpk5cPx/oKRuMY2ZbEaOdDf48PX9g7rSZyO
GUJwaZAJvoc4/Zr3jRUhZI1Ew/6OVyPKPLr86JHnMpf+Q7AK0HI3noJxXtXAE8txPn9DWQH4bT+G
s3OIS7B2qpw90JFY35xX0zFyl5lZryqWAQO1WF7ntVZ+1nUI5Ijyp+QVueaDR2yrgQSQDzrgfXA6
/Luqfl1TW2fJo9FzRvzD6YmJcQiHvLHzFiY07fJiQKz/u07U/efgQ/HprU0p9jRgQg4oGRtJ3zJn
E2UZsukKhRPH/cmCRN4GfgUIF0BFvpL1ZO5MlsMV1Ccu2ceJrsTxsYcuiA2TfFNIefOLSC++LFBT
1T2BhWHtD5u0JoTMtbEM1cLqpb1dFhLmymmABAnvg2xnm9dWcowC11FzE6S8fuc8Gz4/y01XMxad
HrXqXcMHe6MLlTkpZV4R5t4CCwqjHf+onyaHoChfMQr81OpVvJPf5XE3AecpDDgGPLltEgxoxW49
m+HUHAUjq2+jvga+PN0I7ptX1k0Pdfo/hjhbcKC46r26476U69CcA1p/427on7sUVvKD4AfBNtsT
xiO0KIVeWkWqOZEYuM++taEcYHdwdnkI8cDy5pRXA8zzRaqzA0mu2XNai81rx75MZyEKULoR1A2G
xknA8d8Nl7ZNtygk2IaBHvPWZLBLL6Ms7p/gOpVks3EzC/i2zVM+LHmpEmFebMxzo/1RlzTH1L1s
30Ws3Xdkcyc20j+SWDxE7ebeiqUyN4x9c2lL/fld4PZ4CYPC0J/KpbCLm2kOMgTi0uQeDddGhvxs
TORXhOyydjRChcXIBNICdoDcALCpt6yUHdnMfAzQEmmYXaoItb8GbC89O50wV6lDdtvat20t46Kf
EoW9inwGjnlunaMnm5YDZPyglSSIggkmvzmZ/ddl3orM15mKwW4dy9sBRH8LtaQXzSO9g4P7EubR
0Ivq1YqxS8KjIuuZ+3BZMbVeA6f5IbSN6qQpyvfHvt6Y+ehymb9ckr/bt74IoCrTx0gxXAO0ATGH
x84gNFLhOWGmvJCyA8Gz6jLEj+6vI3wRbBtRKOzN+rkPxLdUfo4h6uxqtyY8DAtOnTUIkip4X20L
2xd+Wl710tBL1107Dgrfl5dpqzRN66ANrIL4+RNd5lXpm0dNeA5FRSmj7B/Bagky3W5CtIkiCFwt
lDJ6kvZDZYVkE7ycVKDdTkv8e1q3D7XbKGqBzz3D7AQ9nfmPJ/Nb8DIbpupu2TLqkA3PRcgGG/a9
5IztHYU0EMWNLjfVXxC02noJLUxnDVyu3wZ2yGgjeKJFIlfhiqHdGpzdCw17qEJYRf6XP8nM4wAP
TPKCvGUjM6dhS6QgZbmaQ+XWoED2UZ0+z+q+Xaq4B6sxJCCk/TOLepnLVMHoQIaakrpx7zkl1uXh
u3ATADIHxJpfk8Ty7+TeM4mG68mC/LaZ1ewppeh4LXYZ2tHIAy3zccfGJhAfcWjqn8WMf0kyXDb8
2MF5hvSsHPR7vqif+wIV3WjiYQ+Ye0qvQccYVyGwZETRlcck19udvykcnPbH2jUCNxeKaVzZvhm6
E3MUs6VZ68FJa9auDYmSiJvOD0jXVkROk6Pq4JI9ELMBP3OcaAufOy/JDohwmz+H1Elo9KV0E4Me
UKiuTL0UXnlChn3Qt1I49taf5fCgg3BvwexnyMRhZMAs/Rk2b9EKSDA+aSXZtdLy15cYTDnl589u
+uC0d/acDK82QimnNACr5oFNhZeYuRs+SAqHaRagPP5IudqFRr0BsiFypmiGTA3IOaY/2NSeA5u6
31A18vV1cA2XOoxoL6dptjf8qPgaYnmC0BycusMsMXzIsd4xhWM345pExiBld7sSPuDKvhY1x1rU
AKNjD/yBbMEk7fJTCmQ204JN5dgFtuPQNzAyUAFK1k93g2FzBE27BcZ3FmRZ31SYtgJTUwgtwy8h
KdK7tZWKtauErrf/bBeFr83R2PIM0HA3tCz8EtO2j396KPSdpQ0qdg3Pi8q2gIeezxKIB0KkXy44
eLk04JajjQZ8FHj+3+/M3NCQtDIQ3/Px0TQraJErIx4gYgt4ykb5BAztKULFSl2NpsiabIKIn0Io
0vNOJR/MLKXYBfqCfVcDq8scVnifCE4v8NLWhq+Ed2iNbdgZ7iABBm9ilDimoyKZdt7J5M22PfsM
V5Zq2vVhmX5auzIw0iQ4u3WhLqxyopA6EMHcACfoiXwACQy7dMyWxJAovJPHQ/VeJgvP6mOKOa3G
fQTsr3054zz+eVA/2319kVq4t0QqLfW6cS+6WV4wSosgHynz9clKJkmr8wrpzb+66XJytAO30udt
w0gyeN3l7DQX1AYVFnkiwDtisJlgQZo62QbE1KqJRhceIO3v3Cqpfyx53eiPcL9VEcw0FfV8+ka+
tAxesPGXyPJQ4vKyVoPpYZ4ttRBiML+MjsbqGT/JYRZIuqXQBoZ02SlX4yaf4s9LoH+Icnv8KE36
u/y9BfErnLA9Dabh9/hvS7gxp4wDtwMJDV55vdQPWJVURuDMoo+0YxLq7u19EXQt+sN0hc5OTOpY
zwNeHPbBPUcBXn8HUZRAZxZf994lsvFyYhcZj58Euxw8Yn2zFMeT5df3tRbVEAdynTGjEvNvPBJ/
QDfGFAW5t8g4H4bfbUD7uTtXCxVWYYjGFWg738hW8zTuKcSxXrvdeONvkw5Rw2M+k0HICqtLRPEN
MEJ2pyH/H+u6gUArwKhoyV6w4wR9twhv4AH+n8/FL1YZBY0Zv8DWbZEkWtsDnnQehrXDaMQgjeDi
tMMD2ofOgBblXQ5Q65M/wI1D4tV7B/szL/gW0E5N3T2131LatPi62mHuuZgPvKGM4AafWsMMsNbd
D6vZCtuSsFhElS6E0Wdnb+wkFnU2sSFrVHYft+8aEaa9fm5ztXuluit2vbu0wscuR5T/1wH7dSJl
o/PbswKtfR5n8DO+rvcbDJWZx1an69/V8iN+v7HffQF4OcXZkrxWWSu8J8e1Mc0WzJZVJ/ERHsHk
H0oPz5apKhi79+60PdLr6HZkNoevsJubJ475lwHX8UWgN7k15WOzWy9HpJXn87/ZaNwV3bVC/nS2
jVKesOYYA04RvUxnPK9hzJhffM6Nr1A8IaptFNJ2j8Jh5FB9o26h1H4EPqLSn2t5k6FrPMlYWX9y
T61REbbJRvyVG527p+fzJEAUo4jybFUIV5p0TzzZLg6aKr0dRCR/e+gZEpUi5DVI1Nth2/nMJBel
s9Swj7HmoyOesT6uJmL9IZ4oY/h1hrKU9GLi05LCPUIwfeJbIZrvonmE1l2ARPSBP11PQc0iTvP+
H20FjiNBa5yIcID66Qoi8WF2GMeexZi2tRRS8iEbJoHH0ny6C/11OcVrV0ajwaYZX5cEDMXmauaE
hQD1olIIfGaSMRGTNgFze6I8vM60U235GlfUmZ8RrwCEtevDEdf0dXdA08V49w3Ls+vMFN0/QFEc
Rc9DWg6FIrxrR1mBM6cydzTYSd1/iJWfdNWY44GkUcqU2hgUV1bmK3fmz1KBcoa1iiMsP4+E3sXl
0KevqfDR18TFWkt3p4ni4PqxzKutBYmua7IMTEPhJ8De9UfknyATCMau5ywdFIk2UQWhprpJAE1A
0SZc3cIeIYguLen8EMc/KmH+qGeS4R7jGYdvKEF/bvzfS+sltHIef0S8UnWcM/f/jdUaFz8nWWqt
T5uMS2LCo9T0vTq8HRvirH9QKASatfV3+jU8yN5UlmBHsXUMoxiN6DPO3jdhf8y0PZMkc6SuslOL
3SqZqqUfiN1UBzU7WJlvcZyIvyu5K+aVH+dFau0Wd82rHFYV6kSE/nVsSVmgyGQ3Kp8uM0MTl4pM
3Ki2wuWhuMBI0KLdokoaGn/9vRPbtEGPSQYCVSKxN9yhBgk6FDhA9EYZIelfaAu9M1vb80Q1hkct
gkI5Iexowmleyc++MgElZKrApd/YCCAf1EWl78xYsoEvdH6D38bs3f7p6iyFQbX9NZ9B1t/i7gfN
Kl+Kgj6YRpM9B+xh6P/pyqc+2oGs85TCv895/WvQj/eqLYG7I7oC26gGb2B/GWMOMlxWd8+Wi1wv
jx8wQ9SNJaaxLvJsLD/pt7X+Kgu/g7aS9NcmhRdSGneB3P7JebLo9uoOmqGOFW7NUo7Ip74cuEol
DcMgdXvln8YvqWOp4VQ3rkIJ6b1m72A0gWR0q0+IHwjerFdJ5jeNxnyUlQGbwwuVzD81Wf9ncR0r
yMIOv+OUGRXnOhGrGIl1076CtW4Oai2cBp5Rr4bwCf5Mh5JWelN/C1F86TZCg4ZVUBV+exssNbYD
PiF0IyTnEDm08/rmElCEWffDRvwLz2WVjPLx3jwkwMQMFPhA+qfinCwCVaH2dL9smr96Z4J263c5
4KoQ8WrnvBKP6BK2KLWairRpuojUta2TNphCZYATziLCl3663qpBiucjKK/4Tsr9mab17koyolST
k7AcNbkO6KXI9pgkUuXZQZgAVbtaUojnRfL8KY71mWzObCmsstnwxDUR+AQ1eTxEKOE4LG/iNRl0
aIO+tflkKACuFGjbjDJzr/fezwnXJVxs3HbWlO0h5WtRJYPXaKKDHUAjee1pIDJBtkPw3NjFzFwW
Ce0HRJdNtuO1mFLj0MmSDr8XkXQuQroOoN1uXVk4qutcJrtN75u4irFHN6mtxhYcskCqcyTmrnH8
Vsp6JNfD6UT3B2c4uyqk5CSFHCkr+bCJgsVAGObrXMP0a5knulchwFycWD6n8tahrywdu3Kz9klI
u5ofWCvU1xKyvlQ+2E7g5xkA+OHNUMcNySoTu30Tdj+cXumypND5vgcW3N4mhehLzpy7jVWu8mbM
yf4hbZ/x3eDXnvhhR+s0uT84hE/ABC6SsrJSbgRDw998e/FGWQSN+qd6onjCsq4mMASCGMiRcaBE
1CC8f1sbzbgd6EXJDeMdCvluNkJ2IZ4QDq34YBWARQq340G4zN3PnXp/jXAuh3t+c4C86rSF+ZYp
J1A9ixJYwBnePpn7Znwuoig6Kb5IOj/8345ME7EQccet7gLtKCgA3pYRhUkAIC7rRb19HpSRKjZX
eIMxSEnPwZi0D7GauDJ8adbCjH0rjpf+l9n6SfVDfSMjw06q//vtrbZXbloZnqaSFmKy+1O+N8fi
25/jDrhLNV67IwJbzXKjRrPxxvqsXuo21Rzv638v6qhLcg7Llqpl1BAGr0Fbf0zBbjFUc/roEXZk
9Cg0i7AMQtHrqDHw7yMBDEBL7sU9GWJ8TdgPYPjJv1JhlZvLa/oQjcLlS3nasmDdgcqXmMlm6dnv
b0swNgRrT99s2W8XLe2huf0BTnZpGUH+QK7PWFMh6ZHi4Z3NRDhDu3nvIebTK0OTOVf3F/0IinEJ
dUCJLkneu0IWSvGoxDGkR/pG2mSm2ce37spPDXDfLfxztyBPfYOMuvFfVoxIlQ67deHc3P2mLFEr
IseA8l/4DGNkD7/lSfM5T2fr2L5v95fKWPhAR0YnI3hSwru9+iiJwuBskEa27ZJwgVDI9FvjJkxx
A643ipz2AhyHNkTnEAAkzI6ySX5bLxv6Z6R2mQ+fYauLpQm15O56fimK+xvojMWL5hppFK9rbRRR
cajVag4/ohsjgvxdNGA4+IzZ0RAX+jG2hIJNhTU75ranOkLC53qXNCTulrWjwiAY0yKX9JnW1/I0
8JlfkBpSotsrUCpPYkCO1wzRdiHt35fzi6i/0MC+7MEHmKgfl+LFqCQkqL63enxs8qwQxkZfwIhI
FuBexV6a4UmYKXg+3tz1Xqke8reIFu4PsVv7EdtK/6FObb1RKdwPXd23SOhKworadI6ajMhA3+fy
q8uVqMUnsYQacjSKFvGDiaHm8qGPI/U6eBAELkkh7Vem72Q2xP3M3GugO3X+n4E9/5zpaH+CCTKD
xJYibpF6YCWR+khQMPMGgwBBmF7ZvZKJ+KViDltTdkeYxuA/OHokQ/5n37Z8NMUyEq3JZDMvs4t0
ACqUndRyXM2e/d9CEPhCX7/UhV4IWksp/7ohWXB/1vOPqqAjNYmHZ6GW++t3jPqo1wIt0gk1yxPF
QzmE4n3PXUXAluxEWx/GTA0Td6ZP6J/Tz8wGAJM2yLYMFtB/7XMBEhEwDtmnO7WX20k+Zbz03LfF
kNK4IxXhFHScBD7xOTH/eVGfM12t1WCp5VR3Ib3OdTIGTkU6LD4zfk8Akk02H+o8451LVe+C8dq8
sEnZ2fcCp4lwXeA6110hIVty607khMTzKRYI5QxknT8CbKL+dfvUhSZRL0u945yIzc1q8yxEOaCh
FuEPZS+CUyQjzp6XkFoibOgTH+G+LKbI1gCmvf7L1GQnNa3ffvzxvw/9pOfhwQpJJPKO5A2aWCyQ
CvOY5jE/PSYPgYvmk9kbCKGfkdyVY4DbKimJYY41nvDk2UDjocDy9Kyg1fqLXggFbVm+OY4yuaa4
RwHQeIz+Mce3FYS+rHn8Ga/yu8aU2qeOfqHBTBc+HgwT+JoNAVy8gD09fQjV65fsycY2HaY8GNVt
pjQZRIYdwBVZzVMIFT4EfLQIpems66r3OMhwO/QO9ru/bYRtet0/+9VZnStraIUSTm/WuqtQMCJa
dLna1y9D8O1X60u9Vl8knvlC5UHNjptJXptiN9h5c/epiWMyBdrUw+nZoXsGH8wU9DrS76fdqmmz
jEBVycJEvWOajG4JzgQdGsHQdqCKXkpvLj01y8BTyhkMu5ZKvpoAn76RZTM7h+S9q52wg2z6bYYX
DxbXcguTfnH+NiKF2MzucskMo+dxNiCfBlcgNpUrpehX1gTsfRrm7R783lGBNaXP2ZFzasQXwUl1
sYBFn3kpm0uKBfIQl6AAk/TGANcR9pJa2e6ViqJzL3kX/avlaWC6JXd51wUiwej+1OwkGLN4rQkc
3m9406BfaFGL8vzzKqRXpwPKa5IjM3sQEUPnXZ85Vbfl64rLVyBMPqdLothuJSfi5/s36XsLVGLQ
ykC31GLkkHpIE6Yn/2cltC3k+Q31oaXnV4XtSsezAJNJ+StP85ORow9tqcXVi98NuW1M7D25zWWT
rjieWB+pNMHnPxjo83RCbxoKube2FUPvghiG/tVVIOVngMmpewRRVvS/sXlfhcIer0r2IAmuxoSb
BamLkmj46lk36ZuVO3tnRgGXjjs2MlOOG+AkdCP2xg2Lq6xtjD4ZHLX64ovLny48v5+lpdp+MF8R
2nAe10bq1TiuQZBwtQFlDsjzoawarcW0v3k4u/7XlpIgpuiiZvi+yognqx8KaRQRA7ZbxmkZncdn
eBjC1M0FN6PpmVQajVO2i7q0VSebdDe+AiKZEbUjySsmc7ot8niTNHDCzxxiz1BafwQXkSnLF6wh
572VRXz2M+4kjkvcqgFUnlcwzrl/x4xKHSmj9Hkw8vyKBdxn8gWhz+dAtvLs1ktl+tOeTFzZOif/
HfEjpTUslrVm9U+1GhfByYGHmqjzpwQVqFYnl34/3UF5rwmWI9Uz3E2nM4OC6f20ZbVt25SBPJIH
QRnL2So2PGfSKF2+xa7rs5KWjDHp7TAztPjDXgh3BnCmQ04Ck3j4MnDBCLzNPuxp2epMsNATWE7z
h4JihsNzfCZQ5eVxn5DmzLdHZvojVTv/vY74/v5L7+QnzvComKn/RM5ajfjAsMyO+fuQz6GbM6Jx
gi0koa0/mqAusI+C9heP22mqrdPrgCfBZ9QxIUdLKv324aOsw6Omp2GiBG22PbWcpLfTzdyuzBoi
eOYIwtB7LFv1tEGJAn2g4woMfmDQHUHXvvU7ZI/QhWLHYq9vUY6/TRaBMX+LmWYePZLk0tz6pHB7
AkvyE403YuEvObWkjxGd//1jkSY187RmEOC2QQbowZt8lTjLjUlF2yi57F3JHEcqEnxC6sWViwsH
u0nypapE+VFyw5fCCNDPMDGwQ4mHmD0sK5FRfJFB8qedJvS9d9SS8yLeeuiRO3gJfNFNLPtUOZTm
swYO1N8DQLodwNpbulc/wKEtLeeLyJNwRGw2LxURGmd+q7/yG1ww8JsPxpxiQM7WpyaArHWdGp5T
aHTTLLFUv1yVEq4Kdkj1zuJKeyIgb+EvO6qaqwOHyaSMDG15QBbGyd/rT0y7ZH+bnJCrCGPz00JE
S8kDZtAN1IfWk7Z/fyf79yuzkTvFiio8+s68UtRRaOqu10BLe+Cyz7ZNgDUOL9VMO+Z3YP2gfnwX
sKPKyur/98HMpcKz+tH/WiurPD9mX7q2/iQwYctn/jzlzwwbosIo1M32Yp6Mz2EWCZY1gXzLj5Ae
embgVLQIsmGRsATvBTKSxwI4lxxl116dwcQP2z8u3/jHc6x/oDf8hpjAVkZaVGKTUSVwTOsSRtE9
FnKF+YYNOwI38fiVO8dSLiyknJWlKKi7niYTStMBch6W/autu7gHVj1qWqaJdoDwEz4BPyYJ+fv9
5S6JCCKH9alXEBvtchZMEYcLdjDZQRdgTFDZfNTI/Mf+GhRxnPPsM2wZhOFbwqaRR/QK7gP06cAs
LjkGThr/x5yDnh916CXmd3BPZEFMJTdlBqwrxXV5jQTgRDng9B/l1gK59BuMHg2ovYOQU4VPoAUz
T7WN5T/kBBE29Qps+RcIbqi1X41pD/NDghh0lR4r0XBJa6wOrMVgIb8dMVfnFr96tw3fw+Uj2DHX
WKZjEzrgkJpzuLLEXQApU0ibfC+iwDchPuDk157QtaB+7uTzcQ9RtfE5H+2gMUjc1w38cUDhZ0R1
spEIHzO2+0o0iEaViQoyOtptorzClX9NuyXQvBDIpp9Aiz71ZIWw377eITZj5QQbqSG6TP3YwMU7
hWi4W4obQFmfx7VCQqiaTsxM04eGztH3f8t8stprQParVTlMo9A8yNjDCJZx3WV7OOebpgx02XAS
W72kjVOoUi19GjcO1hGo3ACUFW4ZN8o7KkmT4NXbtEFv54iYhb14RxT/wRntE5HYDV5Rp5wX3LO3
z7t1r3vbPyZvI5gsCP/vSXkU10SqVYlG817piEjER9+ODW/65/WEbSXVGBSZwrQdbMN3cuJxhs4n
XJ6pzZ/yU3MIyuk3Q03E7LE80oYpy4rhHJjBXm7oOHwe5dExnedTcNeN5DrRPr9jXBMVbqxKs+cq
rsozAvT/1JT9mNROC133vLhuzK374g6aTxVkwDuE+tb/GwYqSN8RU6Z+88do6grycAdY3/54RVNo
gA70Cwm0KAnN55i7oVDUDgKmMT5Rm/zB437V3Rq9+4xJGgW+V32r24OnC7UVae3JiL2JORX5ls+C
My/0tinVFe6txTkWDthbp2VdIoiWX4tjsvbI5sZKF8kiLe5vXrmM1NugthAJZRowj4qUx/Gj7yeK
udPmnWvGHDk0h83Yjanf9AfvLPXmyhg7tGQnhvBJ+1CGnWkK+vpLx9cTgHbUlRQEbEjtfTSMhkF8
iZ2FOn2F+PKxPhvqA+74Un0WpDb5v0Yx+nDksihQfsENxFCEAZke+3oOBHy0KRMDGEpNFGKHqor8
nzbt6LMn+3d8rLBbuSFvUcmoGkUz5h8ScI2yCG46dbJ5s5Jxo1/U5v8njR3q+JKgDT3HI8PP5F4S
fN7GZHS+xZON4up6OD1rwJOv9e1lWc70uplCoY79mHqBzfIFWdke3ig784IS4det7A0vJ9kdIpHi
ioZ2xxGrT0y/wu0S188a56KD9LahhwyM5RcsLIxzobXVojgR34EXWz5rhWejD7Rj6H/H69RTwXI/
QxW1kDat1NRAOYaD1gQcCjS5gAFfn9saKp+X0umSKEDjcGs/ob7r30swM2IvEDAySrkisvofwgfE
dG/PqhVutC3KmWxbp8v0CMgL7jSrqBp1DODjbH4bEQcfj7DE1GjZe9ahKknpdfoqBs4vXzBy+LJh
AO2UFrqEZc0v61uQPGFUPeaNEA8Y88kMY07Nnwlbv1h6AE3czbkd54JtTcbZTZ6avHH629j97NZm
poIFjyFyb/8sIE3zWuAZsHDCtB3wfdnUVA4cK2Kwl7RO5TrBKwm9ulPUXkArLyhEPGSgXqtrb88Y
GT/a01b6doBej0VNrBWMFx/luFyTr0MCFv9gdrn8khqKQC/qD3Cb7EolIEkhzYzVZIFKdS8q8MLn
vwyxMbMjDhl4H4F1oQKWxUr3lND32tBzfLNkTGVtsVR8Zy/v/HeUjGIBGKuq3v9UsWBWhxPhl0Px
ZBOqLOHX5lA5V9jNB/cbN/UMiH609m+athuhTptzjZY0egwYyYQirs99aBIY6FFPhC1KyCfU+Gw6
Xq2CJzx/mhu8BSqswjLP7TtoUyuPYRuGlEqTiBiOCEHwyNwsowK3YA0CkGfczOI2FrosYfs4SxlX
SVs2CNRy0liZnzuSwHWQwOwhjd6B0hRNChcI9pU/qvLoLPUhIcrSs2qjDDwF9wyUNVKEafjePR3Q
9NLnKDqexjBBwOHxKjyU1JZkXGO15XvwJs8Uj8WP2WL2LciROVvBne8tbuC1rwOuRYBbMGBNf7W9
SolSaT0/O/KFfONgwzYLSY8+ImSQsSpQ19thMWt39idBp1kYjpS/z6Zm8T1rkXnRgJ9llJIJiZkF
1s2fM9z58gEZA4ivKAlrfAR/jBdMXbKSpcwhjIEvRNMg6A+kJFqoLb32BvJQozlFHtX0sKLit7sB
/8HGneBjcvzU7L4z76ebBpttQ9mfKolMq0W60wROX1cBJXURhEMSIOhE0Iinj4YX2+OnedCCp1nJ
LN2BxonzTLxYk5gItspUWtzKY2IQq+hsVoVDT0lQpQPJAmUHV+mxRQUSWs063sHzPEzdlCW1YuFI
0/7pXqfqeGWdeGJICDhuZOysfhxMGOOLB76rWdu9AYbHdRpAcZOjX1OT8wv7kuJm8K+wTB+WuP96
hIY+MC7ZI5v/CyGoGJO7AUWQfP4m3TECJuDZdaBDriwo1q87WCGmQyqjrE2WehMyd9FdqcKGc50k
M5zx5zmTVO+qjt7kVhXYqBxXdEj9+LhegQrt46o7ZYWy55R+kh++ktH5F19Y64yDMy1D/yd/4n7Z
viUV1Ze4YmSxeSm5DKljs4Ws17xEWvsG8pEDwQU7uEUZjvnfjVLjyCyvXeaDQLVCffg9XQA1xBHT
wa5AJ6ps0AyWHWJ7DEDqKY1IhpLeA0NlzP5jSQrGdVmPc4P6AGVv/q3t7yhvaAA0RrmWOi0DYfAY
OCAwu1+LY5x/MqJDJ2mddKWyf2QcNmCVpAmBsHDv066d5Jjxt4h1BS1WzFtNFfigtjoCD5r91kZT
yk1nfFEk9oYnfNYc+jXm9ppN42lmGzJ7xfNOx3nojRoA/9qCliv3JbwftlOqvPBOQpNs/9rFHsq4
BOLPryKAgxOdvU98HL0YQvbm5fcXk3uFSDXzEbNWI+lfsbDDQBa/V5o65ouYrqDeaKZ09f08D+cK
tAomeb2EIhGdbjIB8IVEMpeCj5M8V4evc98MX79yJ92lWXLHZjHZL/6Yqg9PYy8TYeLkNw2TJd+b
XPo6BNDSZ28auJuovzaIF54k9wtTvhfSLZdtAWuxMh9ZFqOEit/8WE0Dyr3Owt6dg5RJS7BXzcsD
mhxsaVatsK/AkTEH08I2rKdly89lWz1rqZqNAdWFBqQ1vA5SKXyXDWO+f9dq6DqzU1RrEV+zkekl
Kitv+oAj3rPvY2WvSa5Fo+UMBQP6wP9z4SlS3P9A/7I7g1touUB+ggU7F2nMQ6DpE8BJWERoJ0MU
NJgdLxECus77svWOLTqaQxvID9NUz0wjrHCsSreH63Xg+rVxj+0PZ6mTtWSBLhY396BYGbTbzfKs
0kCyjWHy39PrMbK5fhn6jcnTVMAWThzRdyNfm+218oX3Jtt43tFecF4gC0f633vqoz0QnKMYqIno
H1UB5QchmghQeQ2WKssWgpC+JkznmrCsjx+hNVwN+S4aFMq9QXdmclVHdgOH9aqUOlLgamo6nyef
PFDzMj0qZw1CNNGRzH5XLl9D3eU1OyY3uYystsR3g0LoRwSVMFfX2InTP8UJ8TvPb4fpZs0xPTPo
V5yqekOlxMIVQidXDXklaMvERaMXNyCi4IplOPJpZa3amgP7cHvSa2BRp+SeuM7zoRtz2KPuwaNc
6aVoysVjBuDuNaOlspYJydF6TmWS0S5DsXAE9c3jdw0KExvG8xciVYIYBk0Tc6FIaRzvpR4F54sY
y5fbIpj5C1YChZOTn6Oi+Rzv7grBMEKSWMhwLRGy8CBv5K336benzeXvx10ZVSVZFj3MQ1oNHI3H
rF0s3HGsnGZyVEKzIRUESfkwZVzSsKb1P9DED0K9ulqgHFWH6IgUVJeF5wczeby3pivOME/IMNak
mkZYvCGzC67nYIwLuUejRqczztVRHYx9Avi2f1e4dG+ygzaUKMwzfKpA3p6QCMUk9IvxYgSFotTc
Cb93cDLhBGFdfOf88foe61wPaY1oBYok5fGhyZDv36v72FhP9tZpFbUwHEoz9ZtVwaoG6kc2+Di3
3Os4OFHULq0jyL1f2ketwlhrAI2MpMpUxdllXkvokLoTDAZEHr17aTO14ltezFpzj+11T1Vu9qwf
Sv8uWCdhzIZrqBrwQK/ZzPcwGJWGEJ+KoCKdWU9Bzu3z3133taW88PlWVn+gUaZtD6o1V02jMrG6
pCdkwqXl2aFYYUv1MdxseJlVf502UQiA+YLfkAOjpkYedLDtlXITAZonbVWmkrPK3KuJJNkuTRGt
7IUIF1t3yZ1DZbCwVknHIQNjxZDltHsD+4uVfoQy+A8gIyfo8TGMVn30H40d264cg4NyZcHUhvHA
k7aqItyO10SMdoPPS/GiFMXWq6bsad0hB1Lt01kdvbuF5xlscORK8EOcbULsak0YiqGp+T62UKJe
Q+mcCIKiuezOEbM+WTG0nmdNqDJS8IptH1eR+oxNL6c25I9WL1QkwEbav6MdoHB1Ktpae20No8cA
8NXgSablFfP7Y/zOAOZWF3qhXhpNG8zlEsvc75qWEHBcTZ2P1XJhrRwtAmErFOtPIEpx182kSlQ7
S1tNGsfWPLC1Cqzjq+1sE4r1Ig4q8f8fYmVjOo3Y0Ge3W8tpRwXT0wIj+k3fSa5ipvt74/kIER85
bSf/sXbfnm+L7nO+qkoku26gJQiL6B7Mfg9kBKhqimI1Q9F8+Fknw7KkSS667Wfa9gE0Q76zXgG7
2Dt6WCV/8o/OwQvoBI+uOszzTX/Kjom/eAvrwfWzRovM9fra0wxkJGpvMvV+QwVnqOiUsh9C8nty
RP9QsdhgQtMzIIbRydJh/6A124CM+wiDIjNxsgIiZJ4TBdudm64Tp97hzCWvIvQcE1VZl4hQZ/Q5
YZtSyV/DbmeebuamLBoW6XmPuEZyOxsgbCve4hvN2VYVu0dHJwZJKh/Tr2sVdhBu4vLWSpfz8c6P
nbi3UQgcLgSBLglZUi3Y1Btv09Rvzg81wHzOhbUuQ9O2p2dHc+dGw2FTct+sjTzOdDIxYM3/+xNN
CIASBOAw9bzN6fG9qnAdRpRnKQKqLLJ1JNNWtM+CnVhjC9nUaGvBF7cQ3NHFt+fjUIyX35oYbKwm
rrR27YuOGoIR1khMe9UdqfjnX6ks82Jia3r9gpwNB/38PT9EXr0V29D6z2Ogbhal++6IV+fPCMdt
+MWzF5cqt+TVS1MGqJrg3nSFsGHYRhvBk8yuJYwPwu0tDxMuhJ9kxkL6u55l3QbHGU1F0waT1fed
vpv9RqXY0wo93s5ZOUNMbAeSKwMM2lIUhEl/DoyJ8TlrC9dMzia/WgsuekKYGjOqn6t+xCH158rg
KUNrJQBbOQFe3GI5QuOkiQ3rqaTnYHwgYWNLcrasbhnbL3SV3Yd1B5HCJ9obwb9mnkFzotz4Yo8i
54/CJegsUnQb5cf6lh1IXixmd1U14fJFPRddZcspR/A6rsv3+TZlJJZ62umkCq74Gc9LR1F3Lm3g
Kdi5vvrWSKE1VpgmUuKmT1WwAYvN/bjE1jJjBgMe4syqhKG3Zmfmv2Qkevc51HcjUSVRGmtxw3QE
hbObgJRkZUEFNo1rO7RUQ9SSz22TaSa5hYZbAzgZKqIQBc61VRDHxSIcz18+mij8Lns1iSnQ09O3
2itk6JXrJoOuQDUT2ZcmP1H5fXftJENmKfo7F2m90eS0tHhttfjAR7mrqcYyl1XiLdE0s2M//+b1
nhnP/1K7VbPJHSoV1ps9BB+yQ32aabNI8mVz52S9WRg0toMp7xCwBbU7h6h+8fopvlLzVTQOoUll
EL5RmjBWeXpMNBoOPku54nnPlQSrIqiOmapUWyzfgCzISimtAHhIBklCexHz92pcPoITlQif7Iln
EL8+5YiLTvDxTHHwOyFIQVrIUlGWJBvk2Iwyemc/uVFpX0cRlPIvNLyOJfCW2g3GvwnZRmt8Fgkr
XDxqYBBrq9u1iO221JuTcMV2IZ6K9GcCwxiTtJGlwLdL8DgkpBMFoY6EbYlgR2unS9acYiVPdbkQ
U36Zwf/7XTABmDEoM0O3Pi5fytn0AYXwiPKKswgCnWKvr9T8ESEl6VzuueBqyHmy5tTz+wEbkqu0
S5Tg8XdAIRyYAap3ZwSvuXA9lnyS4wr4C8mPMI2hU23ymrn4tlD150Br81nPfWd2ewjkYUQLDcNi
1HPlxSvvFleshylgO3UQXwlUKx2E0UwZTK7c/S+eI/G4hLMVdY1GztvuzPCcCnra31MIKNXzRjtH
GzPcSBKEc4xCwSUarHqJT1AvoVPSGia+E0B2SxgwOHTkqD2AUn30JG+RRJtXx1wy01dHx4NtPO8E
J79lIEP9ijcYqrPPJi8C3vFC/hBghibemiJwBk84ZlOUhOFRIrVMvqD4GVQ+4x6TtKaKqtEtXuDk
zrZR0dIzCNUs3OdUoWs0ISAfC1TNZF8G18kiZSmHfCbbScC6+LViztV0ICvh7OmUke27AZenkZKZ
6cO03rLEGWXGcEBv5zV5KrRcMbYRs831jmFJ7Jx2p1QKcz36rdBG2Repm/Iys3npFdvIPodBKO9W
tEImHTrQZHrVfb10URF8u0JVjtrhGkYG+L59dN0/YgLCaDuNtjSS5QDY03eDItWNGrwVLlyLtsh6
JHZ/Xvm6S4FgUSTu1N2ONYLxSXyEEUMXhYT3hlfMT5Vr9AZizNnSY/RT20TKoppgidgCDZYW3x3u
7qwGOl1VMhF+I8PNwAHbm3ZTbEei8xWs10GkzAb9XxQTdXBiUR3xhRAcWVBvzJbNrxGZkkeSZgHz
PW3ezDGTpS323R4F6ajV8QA6UxYkDSjIy3V/Gdtr2EH1uNn5C4h3HWGdJ8VW0fenBGZ55rc+vM9C
V//TlpCh0Ix3m0UyaMGd3PdzGORHWqfqzdS3hrfNg6AaJjC8MxOC+eam7P9i0IUwi1GlcAkI28KR
2qeHd+GpDgb1gfvV9RDe99Z9GyMksl/GHochYfD7RJUkOC/aCD3We60Eq7WTzA5+n6R6XpqPCRC0
1OJmmvEx0yV4zCy1vKoleF+5DKjul6pCquC6L+kHZjHkxJ/yLSHSLzk371i49uojDc7+t+vYGNvC
qvpDwbnWoDN7Jf+SQB7gVWJ1pzvfaMB00p7sCB9A9oIHVUy1bh1r05hH82i5AJp81DM88KA+V0E6
fpWzcblOXiIYb4IUFNJUD1MZGLoMPD/L7paTskG6KoK4KcKemCmJcDXAvF1W5cEeU67knyOfDIzU
FST/lc4U2eFp/ib5ZgzykT6SYDzv/cVREDv8x4PNU6jLqUQswuuL+0GGeA8leg8klxIblOvy2TSm
+IVZrZDh7I3WPgi1yZn2ki+cXfKrL9GfI/ZvJ3dfXggmPYaPnet5VoRQ0ajmqeYZvnCYEQyeIO6d
XPFG+QeXw9IvJ7OUV6koi4uOGQu+4w/Ls2GTpZSepeatRg5jOHtUwVDPLGadPbRowGfHReYsQmKl
sywlhIn695IXhYaB/wK92ni21niQQB0cOAeD4RIcvjfZ2Vcw9y8RnT0Woy8x3RR3TMN4qlk1o/ZE
Ea3bvUxVwswFDNM6LZ6QZ9Cx9ztEqhEkozfEkr39AU4Dqmx7mqDYtLsFJ1P5NSKqWimDhoLG1D/A
FTuBSf7SSsXTcV7pBU7vbUjr//E2OlXzm3JBbRyaEE9HepI8yFd0JL/MHj7Rhl3+TMg8HJLr8aWp
NMtPxyqrIybNxRwxnx1Een/dBTXuiNzg+E279z4gOn0N+1KyeLynYBdgYbo5TLxpubZK7mdj4iz3
LLrjDBj0S0t7inMlTmLCM0ixAyoaVOryapKO4OXHrjkTT0QzMHb6zByjXRsynQm2j+FsZc0zhCJ8
pGwziwJ2z3VpWx+ZONq5HeNiTYG/TN5m9Nc3wV8v+TDzmAgevbuuzwgrovMyqKmuX2xw+Bi13c5Y
uqJ54h95zJ7gpIGUUUb5H4cr5+0vqmARbzf6wMPdat7/zcIRuWTdz8kQ0J+nbqdyfIbU98qam4Rg
QNEZgUfd31qSBiWWwpHk19xkL3PBe130kKn70FJQ6rSfhTItAv+5sAjM+i6WBChRvh5U8BWIfjS2
eVGfv4FBfWTpMwz82CPxm6WpnSd/84PsPpZxuvPTKrLowvty3Swj0Snizensg1LQnlfjLTGnw9lF
e5bVfShOjyprccGsBlo+LekxBYSrg2AUJ/2z+tM1r+iUjda9wgMMyxkeakMo5hHCdCbpuaZrGw18
CZhLwupW2ZUvu7tn+7EUSwcziIk9oO6sYbiStxKNh6vyaXQFGylGyrnD9jNNRzI2dKt88pzqTuOp
lHcjJBu8lJOI2cWEOLnPcNg7YpSAeiQ7jmUvkKW2LwJPqy7txD6UGnHhoBUPq8s4MjTIkIQeMLzt
K8rUwI+fu+2AfUXosgXkcxzAfDp240S+x0RFfiJ9r0FbSCzEsMNkQ/r4oG9vQDAxKkIWWPXRcr9E
8PorJjx+o3iPbwilY0YtbdsEfQXCauxutd0JH/Tk78QlCpVbq9PrvtSWfQEPiHodEWRopCXWRzlB
NK8aYmEusRpHUovTqT3AioKD8mfeAOEcRUGke7rqeWz9YEWeDz8ziaJXuP6QcGHpGfqTToIspkQV
Pk9CnP8QG06Iss3sbDXycv4Zkwsa+4DrRYTSKYYg/gVRI+eyEAKm32Kkp+/4FY9wRn9HJhJcV57f
2Ps4g4jWnbzHHzhgmlIOUguedzd7DDxwxoGcXzW7z/IpQsD97TYHm9OiPQaXH27T5WP/LX6riue+
RoGxNGnlPwbVtAB/H5cWwtJCJvfqhlC0GkC8KOW2WWjUPvcrNhICytxj4R/KUUUcSUijcUaucxiO
mzihQvvL/qbaKJbA+xPH49lW1SpfX8k2uyhDJRgyGcKDH/epOtSkQuHH/IUDW/C31DR9wsmdaFCS
lWib98lwcdKUMdxPSI5CsJ2oNINOPnYKFsYx/dd8wphI5TpLZKuNz97cuFwxPFlUfDXpUTPL245g
PemQ0W1mWhlMyGb6h2KFdi+M3SwR8pqlp4gxV9bhkzQlNet+9uU6hIne6l1q9I6joizYAXF9Ywhq
7EtjVpU3vs/8IL146Gx8BEENLJx56ZpWmNA5atr/ZnqBL8wLmVOA5VvY3hANeVt2xvALkv8VgiZF
L+qkSUXMVP9bRhG12S7SSJWhNa6SbX+VKifccGWYvgdtSaE2DQ6lNWVUh4TuyXZ0iMISRy+61/dB
E5kT3KyWfpvfRpRr7ZqmmPP9UCSChHCfYVRbBJidH4cUgt4tKqAoImTrYWa9I2jODvnaXQUAzxvy
Hqwn/zK6x4zblxH0hL/BryyTRQhZxWxtzv7GDTvnXmTX35qQdx/nMYfDLNqsPhCKT26Wnby4sQsH
2c3JFvU3ImXACXZOZORTlnq0gAUMG7U0D5qJTGqxegPDYo+maWhkaAatBREsbz2y+LQei2t86QxP
rd97Kx1oDdcuxH/kyUJcwNF+UVo+sn6rBzzj8/3q9oOfFCzsq0UYUdA9xJGjmLQ2Pf0BaicfU+uc
nC+LfV05CNmUn7K1zng+FzYCYfwtMd8BHAl6rzOBiB98GjBYIbw9LwMIgfMMpRxdUzZMfCoGUya2
BxyH30L02OWa/EuEerP2KAc6L/g+IPpR7oqhU0WTMo5b+oc8f9J9Ej7N9beM8bCTgXJBfbPJf/if
TTDEjscjrrafwDAxuPXit5SfXJZams4ERVf6BjQpBicXYMAFUcfd5O/++0JSjTUqW1sDBGLbd4sk
Xjg8KoM5UCJ03+Gb4UWeHRP2YwoO8dDA5ShY0LKL2THkLFlo9c8sALyuCEv7Ite8TaoE/IHY32Nx
Hg2tKmn4hvMZmYI4Oqqm9iMXNZcxOKSlYj2eo8Pv0ml+eJYOZCby08xGG3qj0uJh9TTG6sj+Oz88
8e5Ay0zSuIPUrMUsD1JorJgTKsLwMAV6EDQ0jzursuMWnIOwAYaGKeUzLs/VDwIurZ34j/p2aEGe
GnCoonD4qHg/0SxDD2iIUw19wDJX2iAB8otGasCQapwp+SJ376Ww3mjScAUOe28xBIORog6OOUA3
RJr7RtdSGiN9uY0tlucwGIuQZIymV0M/XWd2fmz9cyjKZ+rzkoEJtXrlrBelG5j/NCma7VXpl1LB
FMPlcemlh/sy0RD4Uv5ov5Isa0LBtBOfshIaKcbDx75iWScoJixcomYAey9L6MS7NJODbDfwpAfv
I6hZ3kM69+0urzLYwnZmW96vCd3EiubdpopY40arMjkjAd4veU+yE3ZH9/fst4Z+lsZ0qNdtzK3B
AQuEPIOKQ6jwLUPKSzJmwq0Tp4SOzOcm+Hn7js2GbTgsU8fzWJMxoXeD8N3VYzMuJCDtNMDzCI7V
HxUm0ca0ctppWtBhYfUGl7vNV7OMDKW+yqhOAD/RtY9e8DuEH7P5JdT7D5AnONmblHm93tLM+qUh
pIoOQ1TZbPxRld1NT5h6pJdLFNTqtegZNm28HMdYU17c1dLQQU2kjwgyo1hmW3OM8rV+5xk0J26Q
ZGlHi6sixShbJPICQVlGlp6bQeZATh3KdN8Igc1121CGahOVRbGAtzz81q+4VEHTiS2+Eu5oLH1q
fuFAehecV7sWQL293jf5tBj1hf2QRDKimnwVHh620NkWmcmx3nBAhSipJh7AQHnQIp14et2W+Dn9
0Pa0oz4VsxxlSyusIm1nefmpgJWgqkwQLKFdHs4+vCiK6q/pdy23/cTAaabXvouUvqi3/CHP7QRv
Uv3GT4KhiuYVrcDPtxkiZy3+iZ4sQ6R8b8oQiGDXicwry2VokZbkRvnCEY+RQ1xm3RjoAsUmeY/X
5NhzheCqlOrMtmd8QAZutgYYHcHUD8ciRK2m1BtbdvHij5hWoNHIbXj8FuV1p4ZkeM50CrLwtSpD
CQsYKnj4vklr0aJC894KYER4F25Z+uBjNbKmbpgnorOqISzQa1kM6bFkD0ITjL8aHxQnQ8kk4IS+
l692dxl5cXKHy9v7tJ9o8TTsKyMBe3Gx4s9e4F9n4bs+vx7oQOEpWSsbzn/oAC8OWUdYvmHxQuNv
8NWtqfj3dEjOekBISOjdYHtX0YURaNx1GOigMT2X5VbDW+y4I0IXFSBAiSs9XbUhw8jYvbfd+Msm
ocirPGlI7+o/A+5Gvn9v3CZ91PGaGeqc2s+oIaWTN+9NKlhQiiaGRHLsB2tl9hQPHANj032tz1b4
v5vmdRuIFGc2bFKrOrpN9k/kiX5i+40kB4sUAsOyou2WjSjLZ3yyOFV0AepcjvFH4gmQgttklYaG
6biKeHmwtwFQBJ4v0I5mVj1JfGgdE6THknXCe8137gSC5+lMN/JsUwQO8jH0wYYIB3va0au4csZH
g0GbInlCen6MfSuDZu3IMB//XJ2RewSLf2aOCqv2JW150Hk4LA8vjwyUHjEYHxOSCe4VJNdpAMFd
6M4LXq4mRZtvQffYiaJClY/HHCTDUedzXYWa/+tS6NLGGEyS9gPr+qcjI/J1VjtPSbQyleUljPoT
xNav2R0feWFkgdy4ZPWgVezP20g2dH9rgArdN4VHW5MfK0TYiqMBkck6ymGzL7HsQ8MCIh4JrNsW
1oJdoUlCOP736NrmK56gSFcxdt59Xhk7NbOW/A6R5qaEvpI6Gtbqd/utqckPmHlPDP3/tSVTZ8w3
j+1wfKXYU7/kfwipFamrCpul4Y0Eqa0mTmdBMeIyqw3Rbn7w1+/4iOb+YIQsWK5szxrZfZOS+Xzp
sjqphgP8y1nynrEW5+yH630EQStxKbDe6OdMEGMaBUG7zsY8VaCcGtPZRctgRksbE6elwxH30NQn
OJW6zbIrYsi5yfIJwdTyELXcJVakKZzDzPI37bhXE8bUdwMvlJBkKcmk3gvx9NAXWQmRG6jhN0eT
AeUJvFhbh9nqthxwcXCzwAj83XFmCJU8XElddyqbdnU9jR2LE18HhzVQ0PUjHiGAo5fLmruaueIs
AnN/38N7EbVH+CKDqs+IjcMmbmVwP5fYjaBSU2AcasRvwE5J+u7pcdOgW971YZlZ4k1HBTFl3kQr
M9rpBu+KNfcfOdZunE4IR3h+2Nw6P+bPvyVKQ23c3UtWn45hX0CkQ79KKZBVSn/4FbyKOGFN9b0D
zm4JpRAcQsu+pcGYtfQnmvU4Ve/kS3FJL5bOGT2mr5Qp+Q82KKJYytilIUSuu+NzowKiDB4xMDJ3
gkM6zJompyrh2HQyY3HU4PnMdu+2oRHLKt5SiEU0GuUK17POxY+Sm1Pp40h0oakW2Q8seUz22Afs
O7qdaXmAaX1yI/iHEa5Wi4NWPsjSxxH71lZW0ywcBJxZ5tB9DDvGvTxG1D59IzROAJmUnB0wdv0d
dMcVghVQjsvDaTI/2velnP/s1313uy0ae4VE7IGtssmQ44KWZJp4W0m2I0gBTMvL2yjcEwtWDB/9
LPJaOto0Lwb00zcrXhO/M73mrTem7kLwQ6PMHvE0A4so6y/++ua5/Xmee2trDXcQAhDxUsbsuNk/
cYH8y4paqgq56VoTJ3VvRM+9XPQJD+UFD5+Z94pEncnE69y4nkQ922tMVICKbefth9qD7zKBxeG6
4+n0+FMB/hB889KPteLbmGITkm9qhkh+7kVVni17Fyyh6qZzineA3TdI9+DPWb4KcyOVJ80O0uTH
1r2aCi9nTNmS0LjIlOOvDmQc5FKHfTzqIXDPHm4jylvB3pj33ZBqblvMwKPsAafTLqtCYrCHuNqS
B5zESP8mdmmx4B+en5U44k3Tfgo/F/LPxuEeGJGKiV8xx/jE3oDmVKaDeLxXP1RTA0QXEA0HXF6n
bOsy/39MejbH8/En2YvORQuF4LVWy02pR1AcUiFjubKFnbuvG4yJeWNWsafWMxhDbqIda9EodbRR
Da/IRt3JHeRQMJhE8T6f8uhWToEbgTnjyuLvlqp7MtyZfeXKOCdxFtPon/c3r3O4thNjJPxZVZUe
/Uh1A5fHfjN1YETe+U8AeZyGCcYkTHc7nz6xTcj5DP4pHZX/GYVWIu7nlZfqk/elVEtmM02lhD2a
fLAo6kFS6Sf4Sx6SYsX16blA9uakI+D6JDV+0RAOPAaksyQTWB/Fu+oqnNrbeBix4W5djrI0dW+q
lOeAhPROIk/TSFdLq3UYgCy0E6CcuRBZGBj/2iOZ5BwlQlK++Y487f1pTPS3KNZVXwOIsa3I15R0
+g8QYv/vzvCahDuRNnW+5/m7UUIeUUdJBC50VwBq4/7l9M4EX86/JL+QSKYnX2TebRkOhyw46kFm
5fU3wcu1IWqOBqWZI2fzptdCPXHeJGHeRK6VKBtfAb+UdqRWzgkM+ZAg6gyVIuutI+8D05jn7K0o
Qer2s/TV0h6vmAcEN+0ENMXmqc7PT7lVx9mzaWBZ2EEIf7KUBhQPDYNXpg0k7k6nmktPJ1xk0YoJ
z0nOsM+IZ0tYUGXPaqtrM/OpBfbat9s8TwYG896gNahzOJEH9QQwqmUsFaE+DR3CeJ4H2AWQsmJX
QlwIF1OqLQZLY4snQJq4q1izHsRUISg9ckSg4iQH8T8muakmZBuRc9Oy/DzW1o+rYj3n1kxkKTGg
bKPkhONlJu6DTX3Lm4SDXsBm0T0nIg8ZGDhB5Z2RYpeQL2M3L04vL74dPuei9kEcNBxs6RjGARxo
fwfJUW60uihsYUY7bRUvOp+V944ksrdSZJS/pn912eNMixNNnRy3wD3RqYIIMYsCbd5Di1wIL78m
PdCxAhx9Y88YMn60K3FpWzrmtXxOanLK6ksAQK+m8raji9snKywQNnM+n8as3NcP/MJAMQ55iWCZ
1fEgS6M2N5aNEO1ELM8O6jL61lhZ5I4gCEe2/4tS90l1Amdzol68uxOIQlS6nI6ARDm6h/29JhjB
1Tnf8L1Sn6I8VSeptxOBR+k5CWMggRwIVQEkAM1spgdMXUewlsFAzisqvB0b2RqRF1itlaiM6vX6
MBQPHMfSEqMn/FuSEHco2pPY5AKDQD7BSuXy41GCICht79V+cUMbk3nrUeL2k1FqEA8nQitH//lT
23gqNg9pyz69N2d5IZzniYU61yhAtyeW8EZYN1Ogqv1pxK+fD/m5NU9l56h4KjUQY2uvzuaivq/E
r3qRcUSccUABkVoAfP3+b6DZ1iiFi5ywdLDorH1LRxDmHhb0xjQz5KCrsTTp5TgfMrviVitfhe/Q
C0zIWzv5RBbMLOqNJfPb5lf7ZqQz1unzZkkx+KyXHumFXm6yKSkLihSzSuvm6AxUrFaKCTBO9R9t
QHmL0m1NpLyzaCH5PaVj4gF+lHG/V1CntQGEHyWlYMVkaS5Mvi0Rp5/N+Exuk5/GyLGKzrtIjeqr
0iFekz2SBFYoVBOIV4lpErX+pPHhfNxi8l+vKoNf9f3mXXAHKY0T9qeAI1mvwkvq0v0ty6Yda/Zy
je8629Va8Llx/c5m5h+NITgbJmt9bLWUU6rIwk5HTjC92C1usZN6ue0vKSMkgfmoEdHNronLWlEV
NlequoPHI56ombaVyAPiH2angIRGC0ezgF43jH2WkyWAHEcOzh+P58aw6w92D+sbdoNorRUNJ1wz
s+9/oleRAU94Yn6W9euV6QI9GBFdWcRFdQvZNNB2aRXPONwos4LqATQx4sjOgg8kR8iAP18fxRVz
14/b0jGinRUVPhqLxKyODpLLu+v2KRlgjfaSZE8hwC1hZfFk61VoFOtcl6kBvWA4Gz4uJwbbh+So
k01i3kGlorJGLPCYnSTzNxNMuq7313oxGfKWA9wSTZGr9nYNCyJTtLqWE6G1TECrZDYBGlcrfLYD
AFeZMk3k2FO/YCJiK3vksnML2t/AOZjEf9MMRm4bLLpzavMKGiy88f29cIPWpHEaS0iURJzW5VuF
1dWWF7VSbvaDtBeZjF/zDu4ilO8BwbtOVNv3R+t8c/CcrKRkCWlmehxlTdb3/JYdrB5OCp4wCto8
WI8alUu1nCLgGPaKDneeMTtB7OQYuRQYoTrm5yBVtlmeSr/53sJsnBpVydbOv/DxKyLmUCaO3PAU
8aunPc8TiZbVCcysMbAYl06H2qouYOZdzoCltGs7+80++nZLCgALgzuUg43eVmChA2dUboWicyAK
UQXgh2mP4L4uBt5WvWJzHZY3Qbbxa3bxT/QkEEhzOwSnIsC8sW38MWd6CEP5xU4OKrkzu4GhhScl
3tKOEEbLvdjCcq2rK//fR7NxVDb3Jlhc9mYfLxfck3xhflIO0YDLMxaa2PEbkcz6kP0gbA1Xje+k
lKCVzdy3H61dZYOc+qat6KP/cjv3ByRJv+0EdKMwL8nqIP4EyuMwJ2urnMXi1TQdYNOWM6N75fYX
jMLvTVN0bTk0roILVMXCcBLE7WN8EdZFKu1eb6oLQZ8KNHL2AzQbw4/osDNrrjen6sxGtocFK5VA
0H79s812IdUUN2H9ohXb+gM+SFWOxLsuRFvU2CYcIxIAuf1xuoRKJGKUt9g0dygtJ6G9whZv/qnl
fucCkWSTEs6EpcBj1RMSBsCvtylpAtTc5C2K7vtJbJeqLlO3p0UVAf5yOl/Q7iMFXZmAPRzWLnE1
YwQO+1zluAdN+TiJwMDT7XP8EwWD5OHUycrWnqR8B+puZe+GNRAm5DGB5YzyMkl0B5NgitvIWVlK
uDZwspFWtothE/1DuO/iVkLKrMbCmLnpZbd8jwe8/sBZAwnds7j6gqVv0pkdghXkFpYrJtE5pO8u
0jFQo2QmDHcPe/+3ck6aDUyvyTk4ivSvp9zqVkochLBJWxVMS2sa9CdvH1MVfcxP4SnDf1iWOYrT
jMM0XKachOzHyy1DksHN5O82ov3g3X+Lh1juLGZcaIriBrRW1wA8vObvnFgd0kk/4oeEc0h0C5zJ
/haYU0radz4ghgqSHk3szLIflUvXow1ANU33DxdA1xSjJ8VEtwVKVdtBBYaRpFOoF/TS9ebZvnE3
2QkJLDlQ6WIUUlnxcS7dv8yO/AfnTUa0lI1D6A/cA/pF/Abx2D1winMl9CN0sbaRJssk94yOcMKf
eWbdZnWw+6wJWWSOYjai4zxylHjB9n/jNspIoEgvBzkIwAKa9xbWyy2DZX8gdlQjVR1Hxs7LbHL/
9razq+H1zVfP2PWX5+v2XJDnLyhYXtnneYb3sIkiOtOzYsjdJIetFKCdVHqjGIfdI+iF0mJbrwfm
OZ8wfD+BAZoRoUudzqq4fhLBQlyr2vVMGEu4CSUtf0W2cWteuiV3aFNSnh6AY6j1ieVcXySTUPmq
YlsH8AZU5hVFGU2G3iuoFzDqjW7RgGE5GETt545JD6HjfJXN35PYS4WLgBS9egy2JvD2fNZEUhsG
lXhE1blzRTF7QaWvg2JpXRgvs7EeRWwWt54SBanw1+TmYPL27aMAGg7QK0H/ywZ9x6Psta/2p2v+
mCPEurQYDpeG7s9FTEoPOAk8hww8kv8qsRLJX9vUOOK0ayuaK0VPzTHs1sF9t55FkueOd41DyfiK
qe5MQtZ1FWCQsDrT1QHzzI3qSkjCz8P+lPhe0u7bJHJFKF7dSBEGyPkdtH6RCX7hnuuFzR1jODAj
XZ7e11KDCAduR4ufwTD+UF1Izuwj1LHlqxylkX5SWwpWf+wXLN59G7ez3oBJBYO1pynMWdLR1yeq
dkI+E36GmiP3Pc000/AfDIeBL083D9uGJtARsruu55v3J7XMFXjUBTZXBFDWtbNkpSYBlmS0eHvo
itrOaiPkL6JPLmGlT5MBVGbXRbK/nhSsf1WMVFfl8eYhD6JWkaB6xkWjUZZB1LSD4x9S55OXJz+n
PJEiDecX5kmgZ2x3udsLYkz5INTJptH1w+iFPsF2lkq75ewDMQG2ZDS/YuaPcw83vdMVAD7oSPIQ
Wet0dLdyTwolCdwAm6ZEpUkgp9jVQv2DOwGAgARMLYY5aycih9BwzhWdvSVjeT/2HKUNakEHzckA
AWNMpREyzu9B8PQJtXq0X1+Z1RbY/Au135Mfo7Z/rN7w0y4OeLDKC0QP9n1iDnRVBrIW7cTSXDwP
8hPNIAOuv8af7sDuNFzNg7zmtAL5F66cSDCnrq+BE9WZAnhVZ9kBmhmgwKlegVYRbOJg2Yc0qXvv
nw9U+n41/pSIWYN1M4bEmaFNU2PbTXwQdjdVsG1kXtu8EkRR+tS9HIq/LGVZcMJcK8yKQnov8t0z
vpb6acseztbuBQZ8U3718LgUNNNx4z0h1DZv4PCUL5AnrAtWDm0reacvxR+Y2xOm3Ijtc8RKujpU
gFHZ3UcBooLlBfuhQLS4IEiSkwjraXaux57onMJ8w9qJ7OoVLbyUxzo90ZEUYJGbjJj9wdh/VbCe
A5ZS7X6VT9xcPRJTT9fMkM8La761nalbpUZPz03bXNKrq877WffWSTRdM3Kxm2xwY5yNhNCm41e5
VCtSrdl22Z2U5qhiQYAZ6ig0/8jPB8LufPnYLnXE54wK3OyaR+AFwOGrjWmFBCgff+0A6TLaHKVX
pFXwszcbDLaeHtuKlmsm4hpEgKUOjKLYJch8yG461t79+nxf5uVQ5utuUlkuvY3hnInoAOSH9dxH
+sWscckgTPz9Cphylv+CCW/NHZWyNldobNZrQsMSp1cKiMIcptoFTnU9V5rbiFjYyRtW5hPKOXlA
vseFeCRS6GDECOmevPU9H7nwYMF+8oa642i4XbJsRc20cBviuoADHd9KKhNWi/s7awLsINw/8BqK
fsn8u4MV2Ou0/QA/D4cc2IQhfPFuvl8ORPa6FiZKwdhlF+fMub8o7sq9uL8+qHkPtRelyEHLDPWG
G/11Xx7G/EJ94SAKjTfpzT7qZy5HLjWRfa72uyU0sTo95UEk6u395lsOBHska82NwsyHW50RjHQr
4uE18F7P/mdeUy7uesbF2a2TGRlGFa99rCOceEoiWhQ5CRD9o8yDofERQIHyimkGIiBIaQIgf/Fv
A7oHZ7yhMYOCPmbwIkchQcFcD1H6lb5Zkz7itZYZ13Mz1lSFTwQxUZYvFEO52G7NJjDNPYuZ6QOf
Yi9Wd8cYcjuFNMsy//ws4ZdxEHyOR2VRIjfJRoFqw8HsjC+EKat4wrB/VDY7nv4iw+JJx41VQ4k6
EcnRoagPFye3JMuOjaWyudFi0xVXZQc/qUp3iEHBRoKf8qEPpEpgsJ2XjEXrI3+yVwndz//nkGUO
tFnE5NFwSv/5cfhmLErGThGvD3CS2u0QRAaDGrHc8bBRQIy68x7FieH2yxbx78B/BuP5ViBVHCss
RVeccODqV/RVB+hDnIa6GWLNAallMPkzMcY7bpRf7xPrrOpfjkl2ipDut5KcZj/qMJxouZ2KjYjh
i6CHnuGOYuF3GnO327Z1CeecHb6s7aRczivDmbSNQF6YANbzWqsbj5CJ9MUjuKGaO02YzG0wujGo
lUko0D3/q5tNa1eIGnMPTfXW1TKr2FhqI56jdf9+VjmodfTAyUBiVb+wTEvhrQ797It/0b4koWQw
QxX0ap9V4ZXA+sSI+m0zfKcUZ9hSzJcwE+VDEdf4pehZdXnbG0Hn5Pn/EpPoPi7h9R5/juA+tagU
9LbYSfHyzJT339sEKS9zVFExqiqOFeG556hoPB6AH+7aD1oeze2ei+iad6FoaimJZiqv5bvebzFR
/ItlM3lsSrxe7oKGAjRpOaj3BN7l5d8SrUiJSbDdN1/2plznJYwRUlc09k27XxBotZpFDTNbzmoF
IBhDFNeN23nBn0JTa9xxjdc3/T0izwP0XHlDRgjAmhRfAn9xV9OjJKNXd9n3GIwKhTztQYAfKS3x
VktGPwVd098mqSgLZORxqJAZ/BDdZ2QJC3t+O0TAhLHnkub64WZ6qrUv0FQY3UZTp3duxb7rIuNf
FubZcypqsiQZ7SnaekMrhT3TWtfnbq6d1RJwQulBW0wg4JhEI0B4+6dGb7ilvuCioFKhp/+rpYO2
R6nX6oLR0Gl0OrjDbKGHgvVlMXuEuFM17H9w1t0i8y/xisvafhB6+Mg6srAzyyEd9N+kGPlIegJD
F0gNOA4pqymKrEcar0FM0k8hPcHk3dVoTqTTf9jBGus26XxCz5fjdq892C9t5fbBG5FPVDqzIb+U
FK+vOvRm/NZb1DXsEbEhFhVABXcB4FEv+7yuhruC1++xMCLj+lGpRAexBXS322XG1wUflzK3OuSq
+LywJkRVdl4mjUZZ+3ItKlug8WZ6X831eonJbAhJDGjNHYr1tWtoT4BqNjQpzezJ56jiUoobs0vg
c+yRblmqdQRVKEwRRz6jI48u9tJ3j/YrhLNw7kPgt80th5CiqNs3oHlV3Bx1rk/YEJegbdWidaFk
ZS1nNzDxCh83614CIvgUs900UuDLkjhntyJyq9FFo7IF3uIdQXStiOax8njOKCRme8OPFyXKWcWi
qRAa00XwmT1idPwXKVazCcZy3PHhrtKibIYqAZegCVhAPsJOEs4OOZhLHxFYxfKI280Xc6o0XI5g
8NsiYkv0165g91AnNyHbjOHZlzKvuUtV5BxF7/8r+SFREnWrBWMurarV/8CZgwUU33W4VA+CwAqF
LVkCkO3nDMGkZGFRDOevdQdGFcWQhysnx5J/4Qi6mW+2XljBwCIdCL8eRam07vEKep11kgMjpgnl
dw0Vnc480ylAcdcjRTHsSeS5K0RALzQ1+HH1kHeWN4o2gjhUXZffK4rJ2QQXHPY+QSnAMI9paqBh
A8kUje468b/gYlPumHyJr8wTYfffq8HVs6MF3dLQEz9yLG0tOyzkGwMt779ff5z+lXrt4gqC88SJ
1lDKeew0AHBTrjyg1NtOvFuGvjHe9EL+3KyoAdK0FwlsVOcbKT4EtFITaydobL9FcNGPjYzQToOA
QiE4sRy4APMLX1ITq0zl27b9da9PBaaosFqH7k0Be3h8qJ9LCrRW7MHsUgO0aKNi33Bg2oBryIq9
hp1F8rKQqVKvrSZ5Pn9XqRvKOaEGeFPTQaGCI/wE6afQHCGKGVis/QzhuwCk1CLgB04KbNBWD6o9
Pu8fdymfI+i3S21gANeyx60TjSKAFR+UksT7gCkH7uM9TpB/WrUgBA2ibXRzRQqbQ/iQpDIQx188
Pc0mrcp5wUpaWfOheE2zAyUyWKdahcAtLPqJdnl/1hkxQ1rCrRa6uf1Jkqo42PqMnMBxFUybqdQI
Q+NDsoQPdcrmj7hIXvV+LnGB57Y/N5Zdi7AjPqj3AFTyzQ5VJX3iv8IVtM34X0oKuvlMR1atW+Ej
JjOds6lA05x4sx/xlkkyuMINFavBScMl6qN4kFXeg3fyRsqPTw7AfeX1Gz80ISzhfJFlwxtF+Tiv
RnunF4XXbpjEox9V+TzwQZiwcaS8TYclwW+AicQtcrIKst41Zn4bonaBx0fA6oZ2DhhOjqpHbObH
lK9/BvovFboPt+ZzPgHvgnzIk+iltI/JC6fqRbStFKl33KrZikVUps58m9SkapLu5bH3IAzXjGv5
qMMHHtJpzq0WuQuU79tOhyul1pzfeSh8dqldhUFa8duTp0iQ0cG/RKIM52FoX00h8xOiSA5pmHeI
Bqit/v1zi5RUypWOXksjWAXWZjCMxjenvCFIegQlStyxsy7v9cyuSw18QHcijU+uYtzWuGA9eAOn
Tj80GPCOZJvdC3Rk3K9frIu2uA+BnBEUuzyVhhOvCO7bE+iikBCuC8egdwUtiB1eT1v6f+Bydr5i
lwni17yg4e9XeVApHU6h+O8JTdz+g19bSz7FKVZ1Rc/EIpv3EnJFJPm3y+PGR+M8f/4WsYJkbojx
UR9DxXEIJRd8RedsCSnaOyV7PqbMkQrUzKTIgWdBa4jYXDiHdxJQ+ARCQGy1NqedemTBdK9eHrU2
jKIjTe9XfhNm7zTDLQlHQE7yofG0yjmaWY03p4HMNZV0a97sicczCzwWZFhN3WVHdjql3qzWjTKU
BpIJFMi8dyw1qIFk9W+zhmPrijsMRvxZuB5Cw44KPgB1smN8N4yh8mVaFwIh5l264TbB5mR/mB0l
EBgZdGFBEIX2Dv/e8oGOoQVNtELpTSZd0wg7pUUvu93ERAGFZPsjh9LY4WqqcHNaHjfch0fDwuMc
4FOfmXaU9HFefZ+3R73hIVYnENf7Kj4huhn4pbENZnKwPoJOaD5TRAtMUUZplk5ZayQP50+tQP3l
Gd+1VQwtZX27q2h2yLIGN5ivBoScM68kq1t778jctBEb5XNXUTaaucW210RZfwuTZxrzI7nSE+Sg
4iuXd/gw/2xOSA1RdHUarkoN3EYdYBIiGMVumnURvIk6QWRLQrzZ51qaJIUziUJfA3QwidbpVY38
vNqR0YhqtIWiWPwItH8sIeBtkQIfqw9oMi6l/RDnZFEYqoavov5W6O+nj4Kd0M1Z6c8eWsDcL649
frWbFJ/FQUEyJWi4IqhRPCNDXWznNM3AZDbpW/PJa7EMGWllWyZS+4TfflQlc3vt0NdaaffIpfvO
h1G7vlBJAC1XPxFdjJYMHOaCYegKBE6nw6miF6avQfH4LqRiT+XPv/YdNYIX3UP5RVC3N5N1/Nsx
vjekLv/fl+TsgBaX8jfSbBcONxByPMEAUxepy0Sdb7m1+KMvo2nRUikGwYBgAQd0KpW+6K/FA1Rg
AUP9E4rJQIelT2jgYc8SfUUZ2WpO2E6sRx6a0aikwWD1lOiUw9AVwdta4cii84Vx7o0rXsD4Htth
Lx51oPQV9lEMfLY2kwk0ZP4G1wELTgOUbhqAoOAEIMq83hSkohb4ln7YStywd3RzlZldZlkIyayL
dp9NxlTAbuqBUmDl/gm+uvEqVx7wNpudpDOS0Db6sLRuPuD3HIjRz118bXM1+pdD8th32kTxcgTX
eeaPMGz494QZ6vDGJ7YD0DduERXvX2Syi54wrr+LWpNbVE4qQT24v8QVZ3bJ02RbjmyZveon4HfC
CIIivbp1JMtXYK4C1zCl8tkfCuapoQVRBfzhAxwC1W6o7TPAhzgM5ffxWYN7Za1aJJXsrtEdZCxz
tLmP+PmWZgqhIfiSn7uLWCbKCeZiuB3cuHgYrnAHGjeh0CpIULtquDiFwQ3EmZqm6fuMbCEK0HCv
kT1QalBujlG5PQVZKDMh0LLtMA7hZ23wwLdBTF7PWg6TpZhbJwra/tpf6ZQegCSs3dx5WhtH/14+
DHjTcIKex08Nxk9oAgTAfx79QDcXjw9QcF+kcNPd0wVdsQ85l0uvUYlrpbDvtvqwUOr2acc44ecj
i8SmqpjgL1TM83CHA0XlBt3aVKcCpM1CLSYNPduFEaU/2a1JxDe/+hJQElCk4JO60dwVms5YC0R4
arPh6mRG6hCtGZGWz9Nq4+GznAx+/iXd5JDJeE5jegcTLfvCfO/qcPtTlG2YhaRNTcE/pcW8BvOI
4Fjg5LVvQ0u69WPqTyIU36sqp76CJfUOESUaY7x8C1N2pqTLslyKFhKGXi9Lzg7f41a+A9m4uFvq
tmGS1aGyl98/DQvOWStJm3v8oI7lT4h4k3jIssTx+pCoirp3HI6VQ19h4I+0h3B5hOMWDjaPUU+O
xPBVy/Xt2Znm1v6tvVQbzYrGIOBZe1/o6xxuv8zTcINqCCET24SXV2q3WI5/2sZenWXfDY4M9ZNh
obfG8tSy4BEGhTUjBhAX7SuUw9zAuv0f0XcCI8kz8hlLqBvkD8Mys5UahiBQVl9+H1qDFCyfxkaB
7V6zHuduOt4pR6eBfKyS9q4wbtgOD2G65W668EV7NcrcLdyyor7AL8iJ0x+2R0RjfCKtc1fusZqj
jU6ZA4CAXg1kJZWF5slBwlMJycHMSWWhx6yx9ulthlIoySEBpeek2Moq3b5PFqmHhIwPOz3TEAZr
tQvdWOKBDKH1BRgvUxpFTnHf/5BPXE416u19HWh8OQLqtT1g4MuwA+YlkLr1c2A4zvwtYolNcYf3
+tD4vp1Lr79rSYXITsJqX1sa+vo8kWhOl5kiDVHO5kFmjRyCv6n4FNhrmOCQvEVRhi2sh9qIqlKi
FlW+DBqk193hZ2FbivzRyHquuv47klTe3uxkAeF8sIpaHfXjGnfUYNc7BSrkOces/R3g4vOJgAKV
XdCaTC1aSmVxagz5ylcjCWIQwHAEekIlHenZJ8PzKxFXBj/HotsZMF/eI6oQ8KvldQXXsTlDreVx
J8o0SEbNs12otgFMEzuHoWrs2FLjLCSesPFvvkuPW0FcsZiTPr6wMiqBud8evDGqjrnWNn/1FATQ
r0R+We0lCTKOhf0LLACm4aUvWprAH0kKTmBw6POZ604ub1RHRBOh4Upe6mOqzT8p1tAvzgIr86+X
1ooBfmAKSPNiZrd17ilEEVNSzKK6ug0+9elx+u/AQ7SbOVnC0OP4ogFWP5xkL3mkP4cqYeqbXhZA
P4vVStCfL1JZG6B4vyuTFIvzrA1YCZJh7f6Daawu9JCbLF8dRlc/ypXgLxbzo5k1V4m8Q0ih2ZCW
tOw2Hvx8+DdUuV/Pumh4oNtRuI57YvMicLBI3ToT5LRtltEs00OgGtsRexSfjYWJEZiEtNkQFF6m
40ADqg3CzFASP387Lq6eLLZojnPnbjTp1dh84t+4gl5KVIgtb2t54fNNcy/PooKSP/EfUtJp8Fn/
WEXCSFJCqC/jlgsmLbA3u99Sm9XyysuCiKge7xXNBAjf1LmOGJj7kFf0R25qlBtDSQj2rkoEdU+h
5bqQfcwGHhy/hHbgjIr8JLJkP9cyEhoPmSA388F6Qgo0R4Qvk6D+Tv971/2o5CwGW0r12cUMooG4
4l59n0D6AkkC1jjZW8ToGWrDq3ylPWlfBdqQEqiP69S+1sMzr2e8SulCl9rdBGA5FqKtcXb1dtfK
0Kg7lB9W7RXAbQFKfoeV6GnDsarqiU/X5kbbvep36iqjUxPjbNVPmfMZ40C1FRRt59gPOR8r0jRj
BBcN/cbmpUX/m43koHacMreJ3yTxh2vRrxCBRUqDZi0XHf3dVrb3y/rjVvkLpuN4Bqp2KYSUsMed
eLQh7KiZWA1ElQrYVFpf3vbaqVmqdeKr3gQgjKcfIF49VF1yo4a/m1IGy4okdrH6VMU3fwQPTzn0
oAJUcU5GWO/sqUg5NZ2WdhhsAZDn/Wj8ruveFH09Y65KAGeKpU87U52J/qO0/Lhz1C0LeW2kojZJ
A30/b0Upz+JhOCF7UkpXGodpSEyr3HLYsg61SIS0yPmP73Y5TjXYZLRl1g78vshrUoQVRu7JQdcp
vuE7MOM/1zaZXnh3GNGIeijJb5jQA77+pRn5CQS73urbi587c/q9NGGJLaW2BxAAU3gWtkk4R6zX
Ogh/bO21DJDVl61FM+TnFMaPMqIvEHilfnfG8RLyX2dVyaNkJyFrZbStbTUzI5rE7PJEj/r/TwN2
kC5IFRE2OuB8JL50DWeEhd0TGMr/DQCEIglGJweKxNGzkL47MmxCtg+5Z1V61MRsjOB7FEayut/V
UEyg8Dg8//kbAGvf5JqNncg0ryHgMno3sEhbwrqgOwAidbb86H8MLmt/A/FYRzEc4TM9y0NUmvxm
nMoZTs5QavfBQzZuNjOF7gHuG7ngcLX1sVR2vkP33xKM5l+X9FrcdLbSfqps0xOGVMqJdAAcREex
nNIgIt3qqFMb+bc6P9GaIGQ/ljSLVBWSg+GzuQ9yD3g8BQBYWvPKwlhVIZtuM4dzNPkd1wKH97yL
nF/EUGEHN+xYTyAmZ2lY9sG5hWFOVdBPmRqlcz0aTGABovs6gVD8xTt3kHB754opjHLWyAtFvfuf
NdCzmS5k71AGrWhNuo0heCmfh1LbH2quEIqHuHk+kJPia5G+gud0Vo69/wY+N0DTggCjfnA7ucSD
7u/706E4vb5TUf84wonN9TIDzeemCh2QC+BXszSMH5LGjMmuA4wk0jCGUdZDbxQI8pWRaDQ5q0d4
DbtJloyO2JF7NWi0LFF8cs54/klNOjCDzopgaS1hL+nZuqmdS9jIYcGWC0gt4XPu5HtyfzqsShSY
4mzNDqSNfNIi9Ic5tBCtKB4hnY1nVFrasYr6dfHlPomvmrAdL7kGEm5PbTtAU6xCCtZIs48mPQ9g
cm3qzaEW7oq5IWYxQnry8mD50Z/1eyiip7mH5tGwRa66Xkx+N5OcqjlioTwsRCNtK/EGzuGVkvFB
5Vh6khQ+kAqPo/1UW5MDWdQytBvsfN9i6wiK/mEaIOVzJFYgJhU+GjO/FYrgXHjJXpPwFqGyD+Ua
W588mu2tv6t3s24epc4h3NuTnF6MKZ9UUz2BICl/fHmxGkHLYvZQYlW9wgUFQ6XGJzn5K3Z0xPK5
UxGTlX37Wo5XLPYYeQ30jPAO83OZuNYYXQu7NC39f73TfZEna3urklhc9Cn0nZDSrFvn8gh2LEUm
Q5/nKAwSTl/gNZ5j7OTOddW65XVaQNuT49gq/toEs4C459FK7G682dMLs86EX04Zf7JBDYCyzJr9
oyMO0YSqA+Otdf2J/bjhPO54+/f/BZHn9H1anaEplGqd/T/g9//mmfWFuDtM/eHMXG/gHoTaxfNT
FvzAZwLwwlzjz+DQLmkO7UPgEEsoqCV/0kvwmbjm1fo8axr+cw4QZOVe/thC4QsjdJJxWb6umB+6
zViKr3LqyYetFwiKwRsuT3uyI413+sZj/xty+fp0c6M/1KMnKu6P47Jd8xXP423WnmIgHzmcbdTI
XYnPJeVFTcEt/Hcb9rTc5CeeIp0rgqFquuiC1m2PDW9JMe08xNLebJ7Q+dLcAD9dlU1DXPWT+Ohx
nV/pVC4T+MzJ1LbFtJCTeNkkKMO1Cmil0CrQRhFX0ykUeAzUXdzyk81zokFZ12su1sk8wxIlrndC
VNeToEsNkNPJCXlniG3i6hSKfB5lp8yS7e6JNT8wK+Wrx4tnFm3ZBE18uoOM7JEjtP0AH9SALK66
61CZEC5uWaSm4+IELH+YCxi9CB5Fim2otm9/exiFr/L4cc4fI+gloftakw+n4wr9U3KI2eULi4dM
jWNNYaBzLEKm5HuVn6MHvgg2FvOE60QDten2XacePSkTCWtRKt9Sxb6/Tp3vgaZ+ZSCgDxrErBVM
o9l7XMhg3djanP5+ckmR3uI6VWB0AjuOcLI4ckvVIe1Y4E4h6CwwTd052eJQBVBPl1Z80/VRonLK
pTYL8oAvZrsEc1FIVOcqyNzNAzGmked+EWtj3oSSGD6dTEYOcj9O5ZD/SkAi53NbGYaXxKQ019m8
ajxGtfkihTYhRGxccWXk53i8jAvnoW/bkPF6ohDvEINf743rcSWsTSas7s87mUP/Ne33ndFs3Any
WOBcXfWP7Pq2pjSx2jSGGwxhQS6xXG02ByQfvnzptGzR3yFcU1/eBfm4oX+IK7efAzQGt35t1Phj
zF/XhIs6wPdc+cCMkNeGnhlC2EwWnFfhVvwMky4dtO1Ib8AT4BhoVERknaonogZeifGqsepOsnxH
JX0OXWJ/QJ5SlgbJbww9vfIfdTzaT9HT8ufJweF1hrpNfVA+oVkCARkJ15vqbKUdCu556Pasr80D
333eS8ur4Zr9g83cbbOuOmCC4udOwfzkSVHjf/wg6USNymtYxCAdpO16+JrYV6/q4bdtsOuTBm0l
IKM7MLLEAi7AggXDGlbbjwCfF4/k0swcN60IrymCM+dllLmAKe+e8iF+p0gSM9MpTe8ixfDg6H0f
3JerntK5atQoMK1tn7lya63SES9MS11JydoxVYELUmvzw9J9eeBeXpazT9xMcdz6Bl9PrbJWjhzX
aELifYXdAIYNgiw5mQ9eXm5kMm5kbCx1Ip2Bvnbvkdzq+Ya9jiwchKTU4EQxNE35WMmO6zlWeWrp
2OfLJmzhIwe/3BXq2B1fO2E+bfxYA9wNeFwRWpyhJPOIiRRK8hclZCU1CyskT2gqrmnBGh6OULrW
ovdenFbiCln91zxJvcKiuOFGZW4pzMvHL036GmCsFOzAJ45Q3jTlAgxtG/2/ONzGE57HKTDXDU/g
bvww3C6V7mM2ZzhTf1oIoeX/kjkPe4bUuXZMo0HTCPxILOkhgZvTv+zpwoXEsyItpEUp1D0cx2U2
u351ZD6+CoyADUDm2Z0ZtlRBvhFIFBTDDRauHsAMgXpAYqvSOfdspw6uU9cR0Eqe8erm11I2K7YD
xVITzlpjGivZmycmrl34sjrF8nnQaDxU9IwjtHOmaIFSGSxhE8zXnxf1jIa3daGmr6aMvjE8AfrR
o/bYhM43nNm9BMM6LtrvNAcbDqTEH4o4JhTgst2h8W4xt9te9GfeTg62hq8QbgxVgoboZ+pK6WXo
OC2GUXDndl1qc7FMRHrKzfITsrA96FMwRua4hwmA3n62aorDfBPvH/NSSDKLziMnoXzn6kkCVcUS
Ee0PiPLK4Cl8HCnLWn/HK/2OZr6psFDD8rFL+Tunfevfh43JMVdiLB1/RujbyIsbkhX1acGaZKAE
Uwc7ssLvTVpBCDCQ5Rxavlof/jmIw+nYSVhPPDIHP1lYGe3KNroETj5rDJu20q0QlrPdHN0x0+6T
bhODlqXhkMHtna4ipxNuB+GwIGX7cQmTupUfa5GMuKYRO59Uceu9+Dni+h2JMG7L9NocgBLjynHo
g7k6gcyMOpsqumXGWXWN3gwrOeRCnNS59BmMr5c6Pn4MRSgLhN5kbh5jv2tDtCuCrcRE33iRrPKQ
y9VeGNFPGHQDFDBla6P2EQ1YO8YcGn7AnGjghWg2/HCubAd6KwM6zf0y/9HUJrdPrvi44c8VIQB0
c9Ny+CC1QMAbTLIqSrQFnoUFgVLH1AXYjWt4dMQ4O4jIg7sHgy9p32yBXoJOZyS8wRo092oWU4Ft
tCmeE6XmNpVVxWTVX12fQwKm9kXBOCix4YsoNYqULdMzHrQXefs54w3x8OeqZtwoWK/HYrjqCxXo
PNtyjkM72uhcvitR5bu3W0y2zX6RdwMLvde2/tpP+ZOx/fPOyiA1Gp7Ber0CX0FS4Wjaeo80FcJE
W1NE62l13lhYYU1fdpdqOIlHmKvaZhVPpbl4It7A7qkvMCHGeqYwg4KP9M92ACoPuIFWU+U5Du25
gkxDBXLXLGLj9A8FPPhOQgo5c1IcdAM1gA2ht2bd4NsAMDiEDY7XFirtUABiu9A/0yNCMfnKOlab
bDrcWnvOfm11skG9WM0r2mCPWsicG5YfBP5hNQvhX9hMr8+qnzZQ1uHnY3+EDJX3WP5GdeRBDtVy
sP8tTPWixDJaDtwQNEGmWlSxCuTSzYix5yMDzH72qTZlf3vfDsCJt3xVsRfDtqmhcmwTdglTbtDu
fs4Bs/qkX0PQEcSXtTIkYZLT+RDbgPkhkceyYHXf48Cp3V7FL34fqbZAXst0RC2TpMpmVqd8xNzw
OuFLBLPLHKYnq/tOfmcP8qAyVwlHtakAfLRX9btFdPsceTgayuoMF0uPbLdKKNfug5pizdZ22nIU
cd2uB5gc5IvlNnLI4F37BBMu834V3BYkGgllAXO8pY7SfpeUNWnTXiUglR2oyrNaWrX1iff+RcUA
YcNcL5Z4qCpc3ZfbdZBhqDje4mxh0/2DkffThbLpcz9ZQ44Z0xXxNSldJe17uFZD+FDcZ2uutrLG
sT4h81e24A6L3Q2RM3dpTYvaybYpdzGP2EB4W8/agCdzPD7PvnikSmp0qXFIbKVOz+s4I7MahmI9
jPQw10PHP7aapIWFcOCvQCr5rYHXXK7oS9jquxQ2tKy3D+cDiCt8OBzdFol4KqJDrGVYu2hyuNQ6
1tkO1Vhx21g2IECYStw2ybvKnGRmSu1YnpHh00kgKN08zv+jFtktpCNdCV/Ae1mBICpoBoAgtA0F
HTUfoy377Tm9sgSJIccQrRm2jJhafzvTcP1Uc76U7YCKw6zD4D6OUyH6GLxDLT7FEOuozfLbbbko
l3BpgpUvy1Nehhaz/yCt6H/wNcFQ9ERS0QOEZ0QcQp+jiIWQwNfH7AMOd5u45DkdMxrz5JWbTTg3
OUfp4RYW+hZ5X2M5f0ltKK3KxFusSeqdIg1kFMtZCz7D9GmBpEcJ6wRQvUo2bFP2yZ1n5jJ97NgP
W1M9VLMJxES6gSEQ7/1P3xX4YqRokfLpjTzqWw58PyjoIfxFLTkeibNprH3eioPJW1TE2Hw6419M
KsH4cHPd27juNruTNs3NSHcxrXuSVYiSzwZLX9z4SkFrVZDZ8CrV8FeYIF9llGOdrvPz9FwVSZC2
sB+xQhA6lOQ0fUX7pnL7UbLrD2d81PjBCYCgERnp0wIc6woI/9EEzZPke2Xx5FXYuxQYB/MD63R9
LKp8H++zx7K6bdS5oTnW84rYd9t1GuT5tk0+T7szfDl9WrTF226ewsOZjxTE3W2I5GaS6fpqvpIZ
dXgaa8AWCBNCnpRQStVzi+DN55knQfwcxwxzWC5MJZ4oi6I21Uf/NEgwLmobY4H+LY9qxBuMetTR
I4Z6Vk6MlfY8V8K8s6YK5aUuJ7XJCDugHLl12FU7QAUhNWu5TpOdeMofZ+dpYjvDEwBMpafof79z
UjaRMSmwo5o9UQsAsqwBKy5rt+xpZyULr96SRuggZ//xFhNi1lXWGmKi0DZlj29hj22q9L6THKEj
huF99VCTRKUG23a0/elZo6L9dBcL3D4RyQVzK+AiLXUsxhU2dDoOMyN/PUlROwLN5R4IlCUNUyaX
IDKdl/FXF0QCat98AvjEvrmwsBxYwoWwbBfNfRdegm+1p73LC0mvAELV6E4ZGEiaq3WRJ+0VeuXu
4EwbAimb4rDVc92TX8fijNTVyEgSjcrFXS+M5C03SYtUU4jVbLpMs+t1JASyb90eUajsH5PD8aR5
SO7LgumHB5/u9o7fg8Q0jYDT+6PYUWmRvaGkPq3tus8ANmyBl+96Z54kfvMWv1jwYypFMDSWP7Vn
LvrqH6nDoRgpI5n6AoKiGCMwo55RJHucqk0jLlS4jBbeil0OwWC6cRZcYpR/4WpdHLuV6vn3YvO/
g6JbRMpFC7bODwy+pmtEJK8BIg0UHm+QyuPd+UvRh+1R6td4d0SEooAY8U8wSpID8VxdO2xG8Tc9
mql0Q4NnxHdaUI33HtgWCTsgOGXw0Kg7T7FW53Jg2XDfxaQSr79deOEB2wzsUk7ZK7oJDSa67zEo
1HJL2NWAIL57kQm/60k7IJVjVVlBJhcL9udXxPe2BYG3vuCYRM5b71RYCvNCGsNzSbROGjA30MDt
Z/Rp9xzVDncHRUJHEa8kP/0uiRpFRrvFxpbHIHqrqQ3LQJnES13gPG2aA2dKsu7carHCOC0DTuEm
o5Wvu+Qsg5AZQ5Z0eOk0pgApGZCNuZDTUXF0G9HPuDQpkeKNSUDU2THWp1oZLMxFNgE4ZoQAtAn0
RTOsArvwQAmYmrqA07paaObME2VZw1bd9S+gabgEIbd+jKF1x2xZPml9Wbp5qgmMvThU3a1UUhLt
KteWgbrhZltS3pYvcY59udqRSyUcSA9QxaUaKm5e4zG5wjhYWSM2tL78i/QGfI6+Ri/tGxqsCa5r
zTRLGhR+9M7eP8l89UXF05THndDuKfxRuk6MKMoJgiZk6b6CWEV57JxaD8AbvTdGaHxDbkWwWcLc
5VBWwHd+bx5vkeEbkSTCRtbL8+wrgGUYI10k/w2ql6k1HDHEQAgI2W8FVKY1vNswweWs+XGF7t5z
K9mYpYp8TWZMMYfKCUP297VqZEQvIILDIFxmWY6EseHcFoCTIg1tCqs89SMaGx7yKUg/2nx/RVB/
XC9JpwwuLLt1qT0LpWMl+maobfabb6K4DjexetrGz3oECD5ZeKLHTenGGmNVSbv711AtfrbfLD4j
2xovDQy/lfdJzpsqcOPGq/foI5sDd7nIlsVcqut+QLJXT+Kt+kDSC4BCJaS0yAxTv4sBpS1FlNZx
lMgR5lWG0PG+UotHWts2Rr0lF2eJmOmBXXZYjoHR76bs2YluJwkAjV0qtUM+nMv1LZXC1T+a89pr
StVIRFf6ONWLQJHqh+CZIA965o6/PSbH57G8eDflQiqKH74Iao16dqGNsrKOoyzjBVo05h7riY/w
1SEDnFT8zY+IdwFmEOlrObRGKtWnnhqQRS36hble5J2qBB4sW0PMLKfqYnP2kLIRhAd9ekDAuWnl
UmBi2pyRRRQvzLrNAGjukxJ/OnNoiSTd/9c1PCXeIsiMKHyQIfYAWNdundPjr6Tef+nW34oYDuRL
IC8haLrYLsiVA1b5GRRUVU9yc5Ah6nuFKm4OCiiLPyLfg/TcsLDSMRnynyNese0CRj4cf8+N04R8
LjI9GEsBaXymE2xdxl2E1UBC+Rw0MHiTH6wC8Tvo/knR/aBrFU7R5HV0sE1qMv3D2Udy0fhEAZKX
7HdSxtwmSauqnATj/LrNotweSjrnyfBdVJUpfvrRpk3vprsBGDUbk8/sMCjWOkv7Ts6/RlvHclaI
f3uvx/UECQriZcDaB/rnvLbLwGbPEomsJED58fnbdcdYSe76DpF5TxSPqh2tokOvwS7TaBv91D92
NuJgbhIyn/gjP4fQNhSSG5che96pnaLZ/qzsDQHy8r+nHFToTgS84zRGoeasy+EBdnvD0jrK2vgn
1wZ5LIPKTJEstAahRJiQUizMjPK8forh2jtVwnSQszTlW6/15ATS/0SO7OFQZ2ITDXdxh0e1PiV/
1trYCRdNZ63VTjYp50hdnW0/q3GrfuzYl0X2nquM5ks3yTWC+4VJIBq8laDVq9XYPNOATLIvyd5a
5GwwlmcUWOFiyr/wDnlt7WT1dGveD1W7+sIvV3WMgk+sR1OApP7j6/tEapKQu8fM0rgThoKdiwGA
z3Xg+49M0FCpOyGPJhYZl+8Q0MRqGZqrd7X3nm/0Lv2QdGwUy/OTGbDjseWODbHdlO+I2IpGHpjA
8Pj/ktukX/vL6UzB7yGsyAYuU8hk3dKvVst1GmPQNqapXpMM790zgVKgKDtWDx1C42c5E0zDJCpy
F/qqP0lr5YjT8QWnPCRX1W1+qn4vmqwPMfwqP6lmSMl97d0PppFLMiOtpKGJHA4xnLdX7P83K8+V
KL4vd14k9j/wbMgZZanium0wOYDF5T0tCR/Dw+4skJCd0LQcgf8bratd64TEiFm2RbT5Gp8ux1GT
onUdeGuBwE+Ckkl7fi+5vpIrRN+rGhMYuZWMJrtQmaeBcbgWiNdzEl3SGhDrqiTa3PQ4ROox12Ar
khT/n9fjA8B67Lx5ze+wK1auMjUZIcMQ1iq7XDjb6O9maXSjq+jFc7mSLoM7p1yE/yPkm1HlWmMY
JDld0dwqGZNGOgmoJu2yJW6JtSlBG5mhDmTnmdkc4q6QiUGy7+tiWOXVunzXrM3u2XRlkTWftlc0
T2at4X/i34/1ShcxJdnmZw9tnqei/d9oBZI28CC2qo+ScEdf982YrcIW2Tgudw3eE/H1RQE+7nel
8aFxhOClvbKyGgwLPEuJm7OnBTBS2iI82106uABvYgMj6oIDG8lAogTnpgDVaHSldNnWTyx4jrPk
AXHkQ4xG/FnIxpn2qi6WA5+8u3bofoQgcYIxCHGSvKfgAYx0qCzCAc+38t2uo41BOcwlbkxu6/O9
8Bc2aTh5B9sj6r5rfyZIJIH/SkjEhxSnVC840rRQQ+wwPhgKkP5RuMQpW+BKOULp2fc6LVAkFrs/
od8GIFefJavXUBjQ9kx0UCvdn0gowlaTwtU/xFBfkHe5dw4fYBk02Z0iMA/IUcpjgM2fueGZo4Dr
TZ7m9jKzz9yVSOmAa4Y+LcfHvXWulIaEpcjc6Pb9Ukn7EPVlJLZsUQSAQBHPkhEYfBRLPU27Qif2
pGWDFwo2SDW7MISGgqnEWeoNVKlrtN8ogvWXIuw1W9cwX9OuRKmTDwRedQgFuAqdyY1qdJ7MmWSr
EAgj5/jlveW7I+VJYoV8RjRRJiQ3I45XFLJqa06MmiJziQXeYh0RHe+O1cFafRNnY9p7J4Hc0JGD
Z2l9PIyWyDFcR7cG+YMwbx4gzcMIQbZon7lGBU7NGTlhpyliXw8cABqaC7iTGhnJg/Z/1uCL5Z2e
MsrcOD9LYTw5rlxhdP0al/SQ46q0NZDW/HK5LRnv73bQCFysKuTXwe37v7IOTpTJ+0f4t7iYd10J
dSDRO0UavoLAttYrvgELS+aU/93ZcQrFZTfQkVBzjLXiUO9mKzYyMXK2H2eofNrbGrqSprYVDbvt
+3HhsDVvDhNa9Z7vWqnI8zv/7IHWqiCDvCu1BER3VkGkeow6Lo/Vk5aFrRDADM+1HW22OhplEGq9
xCbztAaBe5sh+T4077vLdzG9NEJUwUQrheorfZ0tF5W/DDhfw56EZmT/U9I0tgeKJc2vNsWADIbb
XxhbcvTolgOOhevm6+EjEHcoMjphRechG/TVVykvpSMtZ6mP/rGWsrtZms2kfQ8x63ocOqneHORG
pu9fqlVBSIy+a/IbDcxYZ2QpvFogmuw7lAU2LlrYAVn9Iw9RiCQFUBpIGb/wylEa0yJoUyRIIQiK
58bjvshHfacVL1aaajeGxbVVPA7iNiNpSr3DmMglGPx68bcRmKKwemfijejPuJFX2h3FntTaPN0Z
GafnAEiNoUKBukQKYeC+HOhRfX3omUdJOllLNmEjBPV5WfleL2nFx92nyOj+zcyV4rzPXtyDkJYH
o9//zUaJrjDiQiX5DVwp0M28+caEJ2fbsvLA4INOsjCkiHDyr68v/1izgNECdr85KYU/6nxfXLnQ
7qIvgIpJ7NNWfUsMpclA98TbGXzwURp4NP8in8uoDMTNhYatIAdYs794O/q4Njh0kSoYXasc3rax
adeXN0+hGYe8aUcExLQfTz79jGrR6ltbukmkW2sfq+CGV9GmD7FJfbSq+sogwN9BpfZ6nao7z80k
+kueU8eGQUzhLgjX5/5EnVVcNBe1NvJvlKBtO+bROAJiX/W11detX+cagDz2+MW9NCsVqtBLTjeA
UIakF/KF1Dx2cyfG0ADBIzZBl8HaoqINBtiIPHr9uIKxgO1XUzetSzAiWzP4DyvdChftsna+Xbz+
ce/BU+NQMfVsgD2OGOVGtklrb7mGet0+ByE7+5SVaMwR6AekRcY+VXnw2vR6Yl/A/hRw+9IKFmlI
e/YyRiONdMCSnbwEcOXnHasYrgEC3at6xfLviTM7OSFTg/2FkYM2nAbZEW66fTSMEHVy6a8jNBsR
dmkgR5pCRINT5pcrYT65Pu8Q3vbk9G8kb/vhsP9p9AvRJSM/8qdrKeTP62lU3JdLav8DdlUL2VsS
Wwo/6SKKOUmmWCdVDhFY+8rG2aZN5qvz/BlqsexlJgsYLyy4TfhHbHbXhzbnKDa03Ma4TRHGlTk2
JzczwNKLtmAqcCUUP21vZ1ld3jZbVBjV9tAg0Z0dVCwI+seKOoytcSZlQmouTzmR82smuAqymAH5
BRPP3rPYIO4iQ9kkjBn7yNHfpwrBQ1sY5UuXf5coFzoPOmuJnFSNdMtz4gkBpNQLB8MlUfunzfrl
64TkTHhUCJDBtWMwow9NMqeooC32HO4bdhw+4KEqc0HuchQ6SFTtkry9qDaN6rObImh08t2vUo/k
rLgeYKrohebQ0/dyCBrSXckCYI0Ql+sjIuj47ysS/riG1qCTfzWO13J7tpDeT2KWLAe/OIPmu6y3
rzggDyFrJvcJj8YyVwJErofCmWKgweJcHsN2dUFJ0W/7PSFXw4sRlH0VsJVDb4pxaANVz1VvytB4
sYqiVXYxTuBjBuCRThNHzS9Eh9+vfw3PHot14Fh4U+b/Bn7OXaCoTp6L5lRw0SWtcADfOA8ZumQN
tVJJHZymzb9BiEd2sbYcW6dnZTtJ/aujB1AFCdcjRJltQV4kRoj0tARObi+HtJhjjT4ZWJ3bA+2g
dk7eJz3+ObJSF9GHuTUjYmJSJ7eSkFN3FqToykbRshALD/rFt1Kzj1GX9zF3ndL+UYKvG3EpeO30
8Q1EhqHM6W7QIhuA02e6FYjQ2eFa4XDJvUEoWlnYL+lshWsmH3rvpC3tvlYnYPrJSsy+oPwJqkHY
O47Pn30rVhznEsrj66ZRZrelgGL8gdXGn2b2P6LUj3w5pB8/OImvhrAgh9ViGm9W8Vp/LCOEz7mk
aNebyi67jbO6F1+Wkh8L6ZE2MFrCUF4qEEjh+DOKsvXNYgoHJCSMePqc2o1yfRlpSbdWWxh8SDLw
viLb0NE1S/eOnnVQIJYYhXcXj7wxH9QJebitgHGOvH4esgM1frnFVNG1rnJNxCO9FuELyPT9W/XM
xv2UAtx5I4ihYJJLXLCU96LWHTltDdMftuwgjnNizjAXuIcoripFRRcXkafURXqOMm1HEgJl4euA
wOUz6RELtM8628n0qsgvILvlzJeMxVk5dMPVqHsnK1jg7S4iwHtCxuW1AJdyqpBFZTd/Uty+qk6o
dWWcMOfK++cQHZGsQsm5xnisO7pYnoxglv/ak1p1lTqxwG39viiEgEcsx9FzePOSvdDpo8nyL8u3
1AYNewFsD2r5YWV90g2HZ4IS8jD7rpETAwRBRTF6W5XfpnQ8YZeE2puDEjfGL1wih91gjgb5pipb
yHU3RKA7hj3ZZcsz48Q5s2bz1qRf0AgXyFbl3i24W9JQPPX6T8EQIk9yR1oVQUvo3ZjnN2Ti8dWy
YMCo3Mje6SvEAyF8O33bHQqJFgsfFE42TLrCHQo1ih7SxXL30rE+HoSPz+xIppv4agJZGgDpQPrK
GF8tYw5neGueeIK4hO2DD/1YlBbktCzBUpN0sjTPoXGYlHBO/pywyHMs/riMbipeu5fxSzIdNGra
+sGuJwUxHw5nupONF6uYFgS9LWZi+Q48H5mFw1g1698L5nymgbSakn0/7r/D06QF1K4tFBdAo0CF
EXOgJ4v0rQlNkn7MSmd8RaeQhJtngTslGOcXOt0Z1xUiU9fKUmBJMR36XE50W63J1RxQPYbp3aOC
2Q4optRXUOwnx0B0OD0bN28FwESJb9j8azVQgHoMNUKDpuKY6LBK/++MO7DCXhRFYbgShgf6S/11
DBl/LHmtpYxz9rXGmZ2rqFjBKDIdhMLvSpR8Z0amN5S2BNgfPWp/4VoxYeVHPMnH0GWNPae/DulD
IGLaq425JDvXMGkDNqSLHn7NxvcQYIyuPGtzii9+UBpd6QWUpDNmcnnTkHi2SWVzDSP2HgCz6HSB
9C08+8816qOS+hQnJfXabBBzoGp+pMZjXK1jO2Ls/BpqoY/VuFr7gL/vLSs/Nq/4JZ8UqJ2N+0/D
1XarBRbGR43vkmo82LUkIv2TDR9L7b9kkHXdjciPPF6eHe9qfJKacL8EQS5A3q14XQ2k4BGmpNNK
etJcUKi8JAX3d+nE6LO/KetjDGzvtGOtywhGoSYnYGoizIrH0Rz3VqayOa3j1FyfuJQQc8pUiDLf
Op+0ehcyJjMTCWiirD0DOVVxtYIL43fmcK8T3QMy67XkbkZN5Db86l4hNtDrTk7nIb5RFlhGSm6G
7nH+udk7gyj5mP67teKWgjdJWwKb9bRBgWbr4pn4400jF225VShhwdUlwy14tHgIvBw1e4YiFtGX
hpX5yY3S7qqWHOkMwqWWiHqGOxcFuv5ro2Yn36tc5uUY3Yq3sILFXFUMbjxja0frdkBjx8Uf3rYL
hk9KrYZSVyxNCjCZwmK03O3O8Ble/HZV7+Syw05EVuv2GyFxoTTyTMQw3CDFFafehu3eAX+WJvcU
LqTOMXYAcH4x4bXkUDjLPgM0+XZdV1ZyM40bPWF6yrsKUZdQvzvm9f8ituy+e5AfzjeIF/0xEyT0
rm+09W3QubuB7+x1VYXV+OkwpOqWc+bta+xHJleo/gKdNap59LNa9GzCzuPMbaGDgmsSTvWKt5Hz
MNN5b0GQ/Fcke1CkAOmNJZyKzqquE6KGHP73kipUWQ701JwEUsWTLvpwUCD420zGmuPnCYUYi8YD
8Ne/oaZM/WeL0kz8HUev0UEnhkLWqJz28lC/5xGsou0TQvWCO/ZWYEphtBQckO0t86k4bv42oHne
GBSEuRVdqeFuDNEN7hoCia5hft6UW1MSQI4Oct4TCOMa9I7fWij12kjyujw+PlOfOfPvVVLo8N9K
e1mAlVHABypOMGp0u17rdtubI+KnEMRT+LPWj5mW9PsJrzXaajvRbxkysXviK6hP0l7Ls/68lMcu
UtaNFT14tWQkR2Jg98ZVd8D+NMIB7lMVf1MaVrowtJblwdMquztR58ydVCK5HtIVVFQeanga8hdv
5btVe7q/iAL737EVKKpCmdggrS2YsNWytfl6UmandNH1/w+tDovqmDVpoF3RHW4p3EldumH3PNZy
Eahob+6XodAMT+vbLJc5f5zel4vrY1oxfYWJsiu0ceOorLXboKO28vjIAeRnGKQgLjK7VZZr0jwv
hNRa6SRD8iHFk1CsAsGB1YwjW4tAIYnBkg1ezH39LezIUJXP6Asl1+eWTxWP2DW4YIE1KnBHsaUb
CSvoSDdfLC+gzrs1U+DpEEhumQ+jLA8G97XbFTh2vd2YcgzlwBzqUY6EniO/3yAelr2AXv/ZFRT3
xATNYSBFD4xjBJOD6KMV56rADE4nXDLkczG3CetlX/b0fkzxFouggfpdHyr46fIGCNNECFV9BVM/
krTC4JzasfxyHxbuBrXUCltp7PNVx5ZfmMMxg7IjPWXxDuPa7VUR2MhCGIgw64rS2DJepBf8rJ3U
xop4WSpYz5OdHz5a5Dct8knKPR0Fy8Da/ATnTyTnzDpQilDYbtEGaoALlQtyIJLAWHKEDgy+o6+8
5dN9M59pOTPBz/e4tU+CRHFlEMhiK5U8PlRm4ao+VyxCYRyS8OeMPqMA9WNPynr7ohnTGWKkmt+e
idT93E7zlzYIwir3+jHeR0rt0GBqrRz2Z2Upf6fpjGArbxvPk8ciDOIjk8fJOJ1b5Jl9TMP4mdn1
K12F+ap1Q75gNG6L9itZ7Ugm+wzM308uvUwOFs+aWbm6mT8bNpOAUPotfVqIDG2uqztk5Nb3Ckvy
0+IW4l+VvqG5J9UMcp/tPze63bCX2YWtiPd7gGsJh1nCdXQxZooxFs9t5qHRieTVeHRvnsIaHNxJ
tq8d8OD6HyvHCI8Cv+fdXc/nCMKyPwQZR6v5ropd0FReiAarUgKUUZMotvPT10XPlDtPEPMGgLn5
5qmX5QWcl+vVW4UMjvFVU+91x4vbtux63axzj1YKUUIP73D3zQGw8gBU8Z4JlVsfk7ZcIyPeqWV+
ghCAgs9uylVOcNBefDCD0axu4SSvGozZ+H0bCXe7S1LX6RVabDPAWWd+94Szj4Dm0g7TDCfPkEtE
dTQADqijTtEi0Wa9nVtdrCWH3Ng2jWcZpEwMPpMId35w0t/0rOjq2IrAqhJKCPidRk0aVdk0dXvH
RYWFifRtnlfQZsctKCH+4vzgXp64PqvICzy6fcGkbXvAXxbpfd/PlF3tpydIWhJKgiPZm2WQd1Rs
Fd42yyP3HUX9JG/JEMpFXebkt/a8fgmF4VU2M0nj0HdEYrDxiygigl1PJ63PFhxQDIkXemYbZV9Z
gWmM5eRvrkldQruHZH0yYZaKOzMwk0fXzNDJ/aLrIs+vVpCCkmgjhD0IjZdztIOg/Pxnbnq77qxX
RoxrOFLysRBgYxaOheatcblZkLkiXPd5Gt92JMEa+iQArIqQgnhE4fda67NJlOcwJUuIuYafbExC
bLmV5jjDwcBJttIxZkPvsahDl8YlvzKoM56LQ22Lggwk3/WzIn9JLLb3v9V65uZ8PZUxrUY1WRbV
mlD9JUzpRJaDoRS5z7llRpbUyfVK6ermA4Yw79jesoBuWvOUzD7axBX0InovC1tct0Nnl3mh6XKm
L1spl3WFhM0RU6tY9Pu/khH/FeOodHJewcTI6uaDarM45ZT76nJQ7pTYPRSz4cgWudLbXG8tgXyj
UaybcgfTyriJ0acW4+P0RToQR5PeI2DIvzNkldKAFIiFDux8HtwG6Mw+qEXMuYgKj97DdobyQ2Q/
YF3bgBYUxrw3j5ZeZf8Hblf4pDYefUXgO5nHwQPtza89E78J/ShXzo7vlS6br4phdXMe3wqt8bhH
y+oh8oYxZ4bGTMiQbnHYJuMIpb6xYz52A0ZIBYNSlFvJR/9CjRwUTW0k9fa52T3aq+B1WPGR4g0w
8Qls4y55mXsUNnhwqrGxTuUu/zWfCBFridwYv66QfrgdhQucs+G5xkzstPsPLTDDxwjR+ge+ZkUp
zjvVfXNNCnFt9HDDmiHyT2T8QiCPvhYaLMY2VFhJWXLwetXMMz9R/5XlhG7pZYOnY+bdMUbYdP+u
q+X1KuIjbnNEpsopWLhaqR42TPDEbYwbd3yP7KNYQqfFqCc6nVsukzfma4QF5Sz4w8w2Quj5TulJ
a8GWD9lnfioSM98g8e6d/jfmv6qQWJsIWeoX2rOi6bgOYisEnGXww7RPjzq7e8p0N4yI3pqcR/XX
23scnVkgTxsbZXOh5jmR0vGe3y/th2iFTEj2+c5VK/8sHZ4bEpxutMXOb6UEbbZzrlchuIVG6Ctf
cWubsd5H+FDOO6nHkFXHD+HijKrkdRANYaBo1R2k0tAKLPt8gyYs/ylu4CWXRY1wn7cO5l8MEeiI
G6L5tybGQYF3+Hohpy0+kvUQmcCbfjgAT/VBxS5bU6ubxgHJPX89qhyV49KZ2RuPa2WaB80VHJrb
41S91+qUiTCSHiCRaQVpazmdHT/3cZbAdx7btnZQL44owzIBMIUmKKv9iE58uiPz+IcUTb0+HQ5y
JyLuV+5ik1TDAuOoYW2IFf7Hvn6RWFwO5tf/x7Z+JBvHDhBY20Vv3w/n6ShdNJ5wKX/iid/l53Q6
6/96YtVc6wv2SOjTcb/KJIpVRBpiOhuN2vH6fm7RpPWGgh6LwNJo1mJ9xrFS4ExrCXmnxzgr4WaG
oINJ9Z7RLU2dnzY+ijQCxIQEkL3GpxdrP/LjoSCa2vfpujqV5rFZ+p79JLRL3NxbUPcCsApezSpn
22SBs7orvTSrNtATgrkJuWpL0Ya+/WpV7Ks8zjtT4i36Q5NgArhRLVfrqZ9DUwmCYtXp0EzGgwi/
cqxM5u2j2Dm3bMW+d3zTR4IoF9/zzf3Clvf9puK9Ryh2wJTa3tT/ArC87cWX/lZUTobMl0q4dloE
+58af4kN45qQnbrquRJZcoBrX3wUHbuxbpgy44n9+gk6TqnVaW8LQUU2oICmpeqiItnfGY6fvU5w
LFZpdl/Kr/9VbRX+Gxftem0N+/+u8hdqbpEyx1muLI3vURmw0F+w0jFHGkd/CW8GEfLU32BY6xkt
GGwyC/RsnizjvE+SaTMF5ieHWVNjbsNb8wk7N965xQzPEwseI78TipGVyKqvQT5LkUyXuZRXSDsT
2FrulXfy73Bl9JVRkh6B2ECxuQ4NTKTXnhv5YypCC2BqLUn3wrCBy9mEysdZPJvPpXmEt/qTiXl0
A8EhFiMwdXGLUO5uqVrYvMptUo61VW3FtoFqk24L3MG8IMEsSShH0it5UiotEo9GFzSieMUGn4Ym
zoDJZsfqf4Se4XDWlkrs/hJ/SUdHdTjHAaWII8cqPgoxDVqCWIGqfF+kcfxnq4PU0g2sV72nVSVS
IYndxcy0yIHxNS9yeJB8CG6r6RG58m1Up2yXhxs/5sIHrdFkFOpd4lWsStnpn8wzHrAqkXFF5yf3
raMoa1iXG2W5PSo+XduWw+06C9gCubRyRpsVvKr/xlC0lqgFRM0f443PNLJnzbG7S93mXtwjpjU+
4KRfC87n9lRuJCyTQJ8vDL30Zty2Hh1S6eQ2gG6gkkbszjC1aIFhDCqzD4oh2GRp2d4v0acEZ3ki
7q0GsBXllbz4iRsr6pkzEGtHnnzlo26jdIG5C6aVj6dGxgnJ5GrQjlRKZjVTCiVDu38L3IYdaFXZ
Hxtk8S5vzO5gAxwjA/FbdfYy+kvEXj2S9Pqct/WIW8SiOLBOFA9OVt0w41L6uvRpBvXoeINibqFL
LW+Gqg9UTAN8kisc09KICHs6M8KPXzWQJS7/0Fg6lah1fUjS9lzsHRyjpRJu0xkFsgEsMldpp0E4
5V75j0W4kU4d5RMNWrECQngoyiF3TD+F9sAp3h0nFBK9Kmy7911WZ7dhGKJxVW3O2T1lZx7UvlMW
V0GA5aWElolkoHkMrC+WyLD7QvoXl06A6Ijc3uJVN40GQKpJs/mZKOy48/IDI1WvlO69z27V66+q
YlFZs8cfBKnT8CeS/VQGRtS5v9jyXMXr01mKB4V2WcmduvktixbWBBI5B7qm0SCOC7gc9s4c2TPL
U0jEQpAJ5GaK18QGBse1wzx9X9kK4lwIdQedb8j47TiBL77MPoN8lwFe3MvQmNs7f93vtq2AMTTt
zLr4jpuIjX4+JuDw/ymZsp9ijrBS/McJBZ5xkapF15eaQPUDAGOEXUA5V1VrFYS9zBQ+mcP2CV66
ncNtXig7AWh7toGUUdO+0eYJwiB7KHKvyrOPqyrmT3vx+d1kuRWG3ga/h/0YNUTt1yW6wankWGCs
mAllcnCUwCkW45hU1WHbGu7h7UFUMXvUuZhN7rkZWq/v42rZH/HCDxZgsWkEzVCcwMyxPYrDVFXl
itdmt8sogSS5EC+52QZSWWw5T7OdwEAH0ks8wzjYHBQTBXSlYQTdUPrOTZCxg1ot7Mf4J4j2MgYh
p4+cxpudEBJ8su/LeVrXyat/aRT0fC5rjj/dDNFrh8QSL8KyWqQ+F+4mNTX3rnu7KB7/ibWuLQMr
3FVbc7f8kdxcpe6SPc6rl5TfW7GPFYnvCC1im6pA70JLfSXLxAwp0Q5N98iI44kIdTi2mjGKhhon
4vujmOhKRaURRW1d6vZOMbWlFf+NURlMBoVpcXT/s6If9xdFzWy06+q6fLtcpPv6TZvmZU8OoRKV
d4J7ISoQPPOdZhblob7ZK3REse/01qabME2q8sFu7ICEMNWLxQG9UtnHXmE/UGWcdhMdX+gF1b+F
2jQH4PNmChHGUC0tQsBrukXt7wp0kU2IiGiqjrmesWR8NwFyWnluxMDIK09AcdqJGoz26IsKLK2y
4hQ1lhpXK+BCqk8MNPwbYHYvwHn7qZwRuTQw5oPw4zwUBYfGaKTuBi3Z7TMgbg579aXcXREeJAMi
JSrb4MlpZclDkr3w3YTy4IolrJUbUycS8Zfx+5R+qvU4+8UupmqklxRJvPPHyy+4S4rdpdshwoCz
rSnYrmMQPKjN4ySkq03BmNSXyuEPc3ZFqBRo43tzMJP1/AmFwmhvQlmtGsR8RRrUP42P6VPGRyud
1FAaVMqFbJb+52Mfeo4aZ+3cCWLv/imt95QHeG1STFvbyagCE+LKKeKi9PRyIsrnI23p7mPyMpOl
I7buAH44/G5kxf7usB3IvNnNUC0iR1O+NGMTFT4wUKkgHIrIZkFb+Sspzj2Uhn8hvnbfggyG6Hxf
UnvemBmKJCdd9wuQdsdLVP/hIPTWrYS3o901FiOFF6uNJGKLNJxmfyk88GavRiO0e2Wr1t/wCRTe
mpvnmvGqPWq6yJZ4kkUrfi4aGr3sMmtEGAl728ADWx+T1qACjGMJ40GEQVQkBJKwqtpMKHQTX2Z4
WZRsEUZ87zGM1Hx6MfrHiyGP/BSeglOyWdVGYTmx0CjtEBlQ3Kmgg466zLGkLsdhgk4dWE8wXyDT
yO1xGxSWoeDDNLTE2eo+7iM3ARmvgI3aZJpV0hmrVMH5gRdM1KoEFt1rRz3nh4pZodMlWxVqSfsA
Hap3C33cyMd6YJS1N2zDLWNa5uetDik6IuXhr9U4RCXgd40NrxNcjnOap9N+NTi4PbwUlSbMhfsD
j6rcNb/UVI/Lgh5OxduKZ8AtngjbTZSX1z4aEZiRLmc309rNBNB4xqgbN2hQcEGMV5/vvrt5MDmG
rENgBX2jCKHYPv9OiwfXo8AhtC12ie9nQNIe/+7nHFGHst1plAZrCYlU1wONGvncc9rQCSMUghJv
v1JAo1ah3JtXEAABry6L2BJym/h2l24DOJA/DFWNGV8cY7LZTZs2kdEYAaRu2zSIKjVZWKJ5NXoV
D0e7F8eZbaJZ2vfkcx4GJ2xOLeg3+L3RdHFdEOZlsh9Vt0hRu22tHSaB4V24e7eikt1MX2+u1Kz4
wcrLXwqXBV7cPuFFVHixDv6QjpeYBN74CrU/N+fjwbjJUskRMHyX9xKLqkpnc0nHeifsokq/AQpO
npvt9dspdXIfQaz69gP8X+MmwetbVAHjoO1dD5rqBvhubGA9MBSXdtvis2Ijv29ouf917ZzvVZb4
ZHSxgvBPdlSAWwTdQK9SYXtnH69iMwppT9binw9CK/59GqR9r06cHbL84gil1Dq6fAPqbWLk2G1U
sPI7KNZJzEAY0J+zgcH1eAOyIcRNZCT4Qz6gzE4jGaAkS/DV8lx2gUjqC6Ab6f+Svj8w3O8YQdaY
iLTmwxXMJOe2xEbPJxSkKIoG3TLqRuZJh7EyIhd004LZn1nNw4O66m814pUj6zFL1hVtycOvDse0
kxFNCHXEGy86wRJI/5V5SFxC2aA9+pKXleyzdM4ZYV0guTOz3f+ebZmj+K+ip8ZZRxJxi6PNTqN+
nuyzuDIZ75tTqe3W7AEwXKXBZtIdQHQPkHoO1KsZzUVlhj8yfKrAQYCv6/yf6QKwgadT/3nP5Ugu
On6J5Gzt4nCaqYvjo1uRPZfC4830MSMWxZz9xFcUlHCZ/EHPSlKAwPNA0l4D3nPQ90DjRgQ34zdJ
AgfcwD4fg+hBNgUDoitQZiVxLaB8ZgbBDc1D80tVzaIz5QwBRi13sj7AVT/U26A/1qob5H/onrAO
mLywujHBgSvfdTzo1msJcMxuHp+Z7/32U5FxbUiuaJgOpKqfSIiVXVOTlTtBNPQhxluCLyYx3wYs
ytqmuf3A4C7xsyZ4D3vOgTL/GxSGNU2dWOmBEJIBA1x7ZTvfK36DKHv5pfpEgC62QykdwR0ybiHb
OluBqbMnU5smOMgDZN3hXDmC4uswTmyq4V4apCpyTx1Hg7vsabrcEihn32AGMmDWFJJetO+Kmi/0
z2UAv0pAIHjUOluzekdcUo/kea/Ogv43bFyjpC0ZJl/0suLFfT6OjasJRPKFqrXcfUT6mpiQoEBJ
RVOUwN1tlCG/17R3hAwifZ4HzfFOLAzMVQxDziivBOkhk/+UrCTSz5lV7AEnBGZoHf6LSGYiB6cQ
V+85Tt1zD1g+Rm+oYiSA2ZHxVQjonRuhMZFrPrNvmRNsxEK3U9A1GwxKBzNaPLzOf65qCr4CfHgp
SzWuKwnXPVCkhhdgnixXHJfm7ICj1U4gqxEQjPFuF/I1+DVO82jt/VVVS9sML9h3jWfCSiGUOdXi
GKJ8VqyS14r/gwBV0abAtDph0/p7kIF6QBth5ieYaNeGIJInmzzOEJXaYdtgB7Tk9/9vf2aL7vxd
ARgtnSeO2ATq0p4//diGytf9/yvRYRgg7YuIzAP5ev+QTUgr58MKseBd/+7G6qZ+4FaZjszBZSKC
GIhT4a/NdGhnT3/CETwrnv4lsOE5DbiSGwjTt3HzlYL/9XECzgWDDftSvhgJ5ts1J6d5qXfzqi84
B+h1D0vSPxPsNpEOR+ctpeMut6kmW7/gnsYFCqf9co1SwWuTWeHzfSXPa9jIhOFyi9NLuaTVM1I7
emgh9Afj1JXTLp9a3E6qeuU45AKUd3yPtljbsXq0OiQ1ap4DCiNwYw/O7fI1MGR4qY1H3NH8eDYW
jg3DpsCuzAF68hZVPAzOEPfKIDc0aYx7fHzR6D5AOsKgYlg2PIjb+5GrPVOh1lxYWCXk9DHaIXqQ
EN0yhZmYGax1nF+4RubdYfWHdOsFBYDZLYwbysSPcnurppHQvJ8JhcSPmXlWTZtoTWK4aSWC1M3u
01yQAyfsBaR7wPwrncKLT+rxl/eCZzd/TB8j+sImSU7iggx3Foollw/FnGDw8G/n1J0XJVuY+8eM
+Wr/idm8dSNqpbwQ3oqwAAneWbgPYlZnb7NkToB8HRp64RizhPrNQZiWzmxDL4+HDz6Nli5g34Yo
I8mb+d6DV0FfhJ6DduKXUfPsXGCuDR6tGr7JyeYhFBLyzgU/Fvp3L5oemW38OJvnNcIVplk0mvW7
b+4eAJZfZCKRmCcyrtDgcm25l788u1HjzVhRuNnvpmrNcbpoYTywqBgZs4n0tQdsDbbLEqaGaJvv
3fLMQ0BMu78ucSG1CPdJYMAYgAG6fZOA00z+OvJ6uvRFTB2QtOrwLoMakT5HlDDlH/w85d2W90ah
VgcxfKAic8ld0aNhHm5BK3tmHw8x/1ZaNCd0iLVta4No00Kh9TdPpJPiS118cHMMzfxdwP3j38hY
eek/KgM4exzZCf2LGcvxCVWTC7eo2zZ98lyQ02bunuyfFG/keYjzdTWTo/ZwRPPBxH+idv35aO0h
FQuN6qKTYKvz17+n3K+SmqelysUYFFCvXw8DagIInxJUR2+vVhx7EqC9gs5lf5xxsrAGkNL15n1N
7nITjsfLQXgVhQw6IbZ+cRO1ruuiAnnjJL/49moP7PsN4knPnGfGlu6t+Cs3ZCsLx/Rg81WZhNpK
58CTU2hmv0vP1NiNMYYL29XuSacj/YJTE5Yp1sHTiuJ5AfFSj4Y8/iNXkrkKpZzvIYl3BDA4qsWF
Y0CLKmN+v4OrC6vgVXfemsIYUXWdhP49eyL+76kXmugGEEhsOgzcJpd1IkH6mmDu9Efr1YjuTpHs
FgWGrEqAkbAESHYqfkkG7I9T0Y9GkIT5mEWISSW7XNyzV30205T+0lXbAeVdKQzVR+Rz0RwO6TPw
BKbVFx9j1Y5WGJAewZ5Y+r4rQRzBMcSBW54uJ/gONvYvgXbgvIWgmSZ9Cm2CIn2reB0kwszLd8eJ
N4RuOjT5EAVkbiu4kWJPMfj9LmxkDTjEaptGhePpXbnUcn/vfoFdIIzJKGhDFb1AhsXcKig20HTw
d5ZkWhAVDKi0QekKkrIKHY7bYhX4nhKy2eCAjmzJdHx/jNOi8b/UW3nEWhVDkB+JxzyhKutmQG6s
8n+gdUkzcETacoNrh1B4xo2p6pHqogYpGVAWBkVwY+OjQyeyCAhg3TCHoanQ7JNg0OfBg5Lh9I0n
UsGsHflK/WDoNXwBn/HzrNnChh4CB56DbCnrCKER+Y9WZHxQ9l0ih2B3srXVVk1kGeZ11OjpWDwZ
UrvnsJZ40cPzKfXFTDVhLQMpPbBpYS7umkKgTllCpp6kJgbkP6IiIzyJ6BAXNPd+b5Fu2o3vJxBf
h+ouIVKsqAtGMo3eEHZU7bXTFyrASolgMqNnhn8Du5/+2Bl795U1sO+L+okdkEfBL+H5txvtLmUX
TLdR6yLAGJ+cVWAHjq2xrZAd1nzxrXzEd4sOeh4anfm6yE9W1/+iJJAwV7jRkZW6WGoJYBXw7e+E
oIgJ7adTHmAPJECOa548TjLNhYR15+oDi7Oarw89WwcSOdU7pXGPs1xUQnFcC+xUps0joGvPrLRd
KZCdXDBvaNGjzXXGQV/pYJwAKiTjZeOqs1lbjmhdr5PRjt8b3LTcMNKeioBIAIJ9XaLEHnOsxVVE
DgRYLU50ET4yv7e1FjmkLtDgFvEvhzcYundsp+aLI34/08MmxWFZs5+Fq/CX11hu1vh2s0oGKOcf
9hnFxU41i3ERX8T82Wn53HYV1nUwWYzDOsM5bzdQP+z/HCN7YjkefLrk0VvljqAwx4Zp7yry3bxY
GTL3fEkox/JVnwGs46ZOu6u1l/MWdu1lj361f3ojEJOnkRmUoJpqKPEzgtJ6Ji1YrHqgVGt8bJzA
dcMCFDcBZuBkCfcEQBrYyuf/5Ni8wfvCCqCKNMYloH0aIh8+BJlVCI+N6vZkerGy6zA1Kl5WA1xd
NCguyHyZ7kOBMl4/mUhGcerIQIoX40mWAUxjE0lOZePF525KyVnGXsHkVZv0iRkApflD7sy5e8+r
b8BhXvjKBWFzjoWx9rjv88QXhwyydpm+tdiUgBiyuoAMpmasY5BU8zB8CRnt3AEt1/NReoZ6JFyW
nKLsRBto7H9Ope23WdfBi14HiVkzIPZHYa226kN5I9ERtqkiDYM4FZPmB+gQO5vzhPXgP4TBzO8w
iMbRdj9qH4QcluuFCsc1Ijejhq4Htgig7sigWGBYgocCzq/3dpHqBqogigZJEK9i876RCqp/j6cd
BRVwFLJm0jONSJdi4w7scB+Y63cTzwGPYRBob9souF/ZmBqt7DAWR2fv2F5qqSHR1n+7zTBPOYZc
DxbFohu+4Txm1UNvxBg8GV2ZpBWdjyw0d4FcKZXxtNuDBMc/elOXttAZD/kleOdq4/qme1vjJVhb
CpLHIPXgXB1/+sEDL4in9cP+SIw/C36fmo14RFoNTkBB8/bkwkbUvsW+4B3bnpAvlUkZYxWwy9MJ
1AWICkrAHcnhn9IhXsF3TD3L7V4AEcjcM+f2n3n+CqzYge1a5YDt6ERB2+L/GFWnUYLn8LHMEIqM
+IxYfAPkFI2GttQfISK2Ux7YYTIOADx+GPML2YEh3uN4nT0YvPg5rQLAvfGVbCnT/9ExZi0dCVEv
8f/jCs8xEhjsjIWvZv/ZLotsGmqg415zSr87uWaS683fY8yu5gXY2QYUbraW0UitRq8oaMZPhkae
Nikb0CUByqIg40nCOoPhNQFOxfVo6V3dIyzQMm0+7F7SExAzdqNHecT3kMPQAkedM1rlFqGYluTM
PAjxp3jYB/Noq8SlbDKsbYi3z2SLCL2O2dMnIL/V+zck4AuSn6SHoX7APfxevOBmiaMzXZFy7Gvr
Hg9ASzZaHuQXWA/siNb6XB4dLqq8omCgV6bNpSBKoctNLLzEOcZx8zHqMEVw4d+7XJwNAGR+HfwW
TCPTU4ELOHZjnX9gaXdZuqWcGu/yT7QwJ3X/iPncuXHxwgLw35Lme+vq4udYghrfFkzyOKFcFGVE
giV9ohF1EuL9lgM6fjMIgoHCXCiXW9AbvYgrfDvjW0t2NqnmEBsKPfhjrLRsE7b3Mdl4GlYrdwe+
VCSBvSWGeX5mw+v+0dJX8w48v623Pb381HgdpS/2eByGDI3WMoWLsCDuwSuIZBDguDMQHNzVSp8t
Ch9gwf5CGz+028AzBZnFU4m77TtmuCzdA+edYg8xDM+u963oXxXgRJhwe/d2TX+2byAdzErxb3PB
LDWkZ/JC7E/SXdmnKlNkhJulKkcKj42QDgpzdx2VyPpcMzcq9iHKca7r9ol7ub965VCb/qoGCmIX
+BSBhj4jLrST/1tYzYlb1f35GRxgsh9qidgcnAixdtrWRld+/adJ1712BDGXpR8w0TUD7zsf5SHA
RgR2i1UT4u8q+3dr9ujg1vPCZDMR4TnWrxRisuOAjcx3wVW4cqwS2EmQedkNGWm048x8sYQ5T/jd
W49k16YEv8voQIT4eqe8oOeBRUp0JM0ielb4C+qSNcoHhv1ctcSta9UI5BvKhInFmDKgAq9XsFck
cxO5FU/W8zH+Sm+K9z/qUAeuBuSO2GQsTHDJiQwm6TFaVgyaMhLvkCIaJ9cvBgqivYh84MMrb2BU
o9KdpyVBwe8pQewfT921YjID1NbIKp7ZWOuJ5dW0E5N9h0pdMWHY7igUd9f+kV5z/oSLbrA3MQy4
eDk9f21nZjgenLEngvxHaKUxE6dNQOLZ6DXWjm4pTYbeL6dZKM9QeD+YSrmnkwBWsp97nmV7ruEm
QV5XkIOao81luaI0J3jBXzhqFpgIvxPwovtSP7fQ3+UBx9hx08HGPcN05TZG1srjipRHGZzMr6zj
eMTLYy0/BV3cxntQsXVSP+P9sVbocmBXcDQDjbD99D9RDdmTYhiSm7Y9wCNf8dr13l3z6XQ6AqHH
dQeHu3aoexPK3zjgWYIAceM4s8JlNh2aCFxzpkZUMNBs9pGe10v5in5DylJ1PSn0sLKN4/Iy3AxF
cf3CT0DsKsX9AosFx1fbqk3pKfFyVBQ8wxbYOnpYcdvqc9tVEBm1Gnz8d1RdMt7akQ79T62POQNE
Pb3osEQUlzD76AZBPXy4tpHSC4Ijfp+rGEsHTu+1Pyb+xb7cDpxCxe7PqEzTJkKmuwjLs6RD0BRa
UYM8o0Bs/r8HZrpiXa+JX6xraXrJ3XaqgbP7wDN74wvodwt3hs7grfTEG0h10WFkajE05FSvSgFw
2eyxkE16Mf8i4ABiRMV8sur2zP2da2KhDJ5/6W1GyKZ2/prL04FP8m5EthsgcdgAynrUwau5KclW
+zMIHQf5/VGcqTXId0oJoaj8NPvnzCthozl+eU7zhAAIi3359B+gpRGsJFuIWMIxfC36ayP998Sp
wkc7fhpjM4J64xan3cSUsDYZEQt9n6Lsf/7sbZddc/6UdId2ymvyg/Howj6avSn4ga48w2sO7Vuv
vBQeP/X277V45aLezls/V89F7A4x0bkbHeGSmIQKL+CnjAO74o58xxrJufG+9fR2ayr7liZMgYrj
y3yP3+e2RkyEo6y13VbSWZ1mHp/u623TR/vtOopdvYEkZyNrBPH+k9vGECJiJ58p2SQMNyRvZrvX
YsUj87Gl+Cw/s8x7q+Q3XrBfgP00tOfzuH/tGfwTi6nfmP0r5noycTU111KGlCm70vjenJGPshxc
wkP5et5wafSPSTMBVzarMGteOMtX7+wY8HGtq+0OcpC3JO3BLZjPmxWBFk7A4H4VnMsVKT8XQidn
yHIpUJfARgfmxqmLaprwKzTpWi9PMhNokMfkqcbRlMr9veu+zOvjk6jOwki/F0Yvgk2eLGfqcMND
qu67TRMFulW8dy0EjKA7X35189nEpOql8rCNw/w4SDSKRP+IvQduRY5TQUH+dOKJuXQiW+pwH5TF
y0OEL9aGUdOS2+aFI7TraxSCrHBF+UBzZp24YcWl9MxDssUdsypLirGcyDoB3wnrJceRq/Alif/T
1nAdPIhpO/HsGiXccUOPctce1lcmZW2ukM/SwNsVvLbM20tqOJwMVFepIkq7ubS2Q4t2ljIIPYyH
GY4PdEUSmYWNCUxaWP5q6Y0gIlecV4C6drdNthd2J+siPV+GION3/ajeOoy4xOytOYr5M0I5CfgO
M39hTZac6Ie96U4d5Hx0hb0nxyx9+qFevbi5lk5IAOQirOPhodMUpR9Jsfu6jLWL/t7sYqBtkA9v
O1ukuHobF5cRnz2bBR/LmDhKItg4vYmoCCxlhKXbnbQaBeG41koFVsoy/ixkjN9QK39/6t3+4Lj3
JR/C13NhCw4+Z7mpLSE2dTTpsQMuhspxISj8RRq7oph6a9taK4lDuU0KoVn7/5extnCJgtm+UwA5
AaeO2GmiMFoid4m5nPf5DXDH0ycA2wOJN/+SWF7ugcvmnlI7LqSjNHcrp741dqMdkqpP7xWLDpa7
NJEVoVuGME4mFm+QOrQN4uhiezwCbvC55NMbAJ2/j7jU3o36SByiYCMbTxVcUsbV+233luj0zNHn
wwK4pDn1F5PPIP3KYUDmzijeYX+wp1QqzQlKlXrscwCtTyjjw1o8B6252HNGyrWLfUMEQqXo9sGO
kJdps6fCAkFgCAfBtlAI3lBxsRH4FbG4o7re3LOaHpqkza5xDoHIxDJ+dyJsXVXU2viIAETW/Lnz
fOqeUsnLo33johYkS3lu+wTnWr1lh01RXdlMjJdgc99Pma5Zi2uZWg2oqQHFtNNswoXQ7+KXVPs1
ZbYtMMOegl+UCSaJ7vz/3MULYu7bxduAWYj5iSofPdDFRGXds9I6j+bDWGzN57WVfPIbMTqSefpT
swdQnD1B4I4ePuQq7J3PV7bRK/pK8Jh7+FbheTjjvXtcZ3wcGFTgn5LnbaiEzyBAMf+QQfLL61u7
lRKEDl/5zt/hSz+jhRNemDdkEt1KNatL5NC5tN5lGPAV4yBmbfu++dbcpoYfUzXHO+e6dW3dItrJ
3DMa/IvE2tE3EMbJ746kFHW4pjT3sj9bCXRgLcgjSc7kpuy5e/uH1vvTefZSw/5+j7A+JGp+yOGJ
/9o0XeUftOR9V3TwE4geAItGuHutcpgbGff+jaPTYv25bg2EycClSrAurrHTl27mfBiSutY9ajKe
CAeEknrSCmAzoHmVvMYKDkG31GULJADekzmXOJjbUeEai54euDdFRcZzpAp75/OwOmZSbPcF2qzy
8lUTwEoJPp/U6Y+RL3tqk/xN4iIm4v/Rt06o175NbRd6TciPovAtoj6jjF04GiXnuhTO1XmQp2wV
rgurvj2phiJSmWFNRknEQ+iKgoBEzu2ogbUM+zll7aTVWFYwnFHrMXShv9blRI2GTcaTkSANS5AK
SX2LyHEpI9skwwpiS/CDA3KnfwO5wyS5YOVx6g0ISTVkVDWm1hVfVdqutmB3ey/bKrDuJKfd8fao
c4hS6prr1rnx1tlx1zqEzjboKOfp3AQjTkRN3Klgv1x0eJNiqM6dTsJ4Gk2wUdm/hqn9BTXUg5hE
ro6l6YVfZj3b7QK/qOO1OdRhGOi7IERr6W+6441s0POqDuJMNcGOtnxvAG14506oeoMVVhvQC/vd
mxUEHpQt6W0vUEUelzLlNgV1kzl26sbQNSKsZVasC9jUgMZtyD6rZH+XhEY3QF56S1Y9nyWiNkto
EYbXT4cnoG4dVGJRwbI7+8ChKpQWTT6W76dlrr3CrmLuzZd9AgLmiMqxD8snQlxZHdG6kayK8XhO
R/WQZId8mUUfIXVo6ESNwpZOte51tkKijMLgZRO3vXicSu4X9/yzilwGW2ZogPwhqpO94un5zxD0
f9mkAGvIOwNNcSSYdLZ1rFKZz91diLjUAPHRq8ukXWQ0c+ME8yhihuENoaneg67bam6v9wvpZRlk
QMQHfk2ySy63s89SABWiGXJIkYK2K55UjkpTnIwHdftFM9ENVX3W5rFWQ/M56U5phfDLW6D05FCh
f6hw7er+0rLp8kzSg4FLHMkVdX6CQvfEeMR4maT/J5iJMY1IoA8e4QQDJVGtQkGzit53fXlvuNTS
L4Fm0DrZ6hTFkC1zhH7/mpigviKbuJl678sKO3vR0j0nVOfpPBK9BDpcgES0ZWoKJNgl0yDuw+Jb
6uQ+Ns3IFnyjkGTEc0mxVOyyhxS0ETMrjCLsJgUycKeb84wnMpGMvrGVWmfbzaysDunW9z6/CZzW
qxCzmP/exJqTq9XhO15EGvOB2kKXWh8vEdFbgPpdLe7R++XaHYoeWlCxBPIg7dKFHhHiR1lpLuJ5
pgr0y3lVCPr7PJqzS6NF9SaoP1zRIVsq1U3z3+9XGbmvbGJZjCHBiYzFBcsuVtXTkX3z43ZlFLAD
4tKzm9jQ4xWMpLxKffXIEkwmK75OI4AO8W/pFMnTlMQ/Byl2RNX0JkFs6mwjSsZ1aNnmHgJKWdSU
Rhw1PQdDwoVc/f1Jm664K6Hqp/rZOtVw6hwhG/nU6PyB3xZG2AAHLkgePA9VFwEb4mrTJTpg410N
Mrsfyhwysvft8Som/gbk6PZzwl+HkAYUyOTF6AuZcfp8Tusnp1ICTVArBMvD5Ocrgi46hybWAPxK
3FkJojFTByDuaCi+s9J0jsD3+O8cTYCulbkoa5EBiO1gTDZx8pfztooGgOuRrcyC4iYYcrUeAZC6
7083BsZTxDhDCZWdKH7rn5/vdkWLWjYYfwpzmgXFoFyWj5zDom1EuPOqwgZG7gHNWeGeAlGeAXQO
iqJ5bl9/74LDUeXZcL1GWBgwU9ik2sCnVTT2RXQURaCMZiUtORxfzDZWXr66oDNqASb+WVOkxZw1
LIdJhMwKBXVp2Ive1q90/ce3aa5lhMTopj+uUxP1fmQHQirVzOpzJcUMs+AhkWUW/WQF0NA8wX3/
cRM83idESG1mA6jz6ACAU+HtUEjg89Mm0fhxBS2Xe20d4hm8wOxhrQaBfvFwclkxOxMT3s8+HP5D
Q3MR+ddgIBtSbgSOWGnQQ6cbKRf+v5HAKu5RMoI8Zf7Uokc2VqWdcfy+iUeKN4wb0SjAFadKVKNW
14ZaxzlSbZqnh+oSOyRVRJks47Q+m/AhQTtUTw1qmXjcMBTmJGLMO7Eqjg61D3LonAZ86B9m7PSo
PTddNVYz90OuoBE85ShNI8U4LARedCZOWVdpPjY+YjvRXJX+r0Jewc1qckEfxIZDe7qvjVMVgyP0
F/Gr/CIpEXaExpb7D8xuebBdtfi37Qx6GwYQvv5hxe+qipNnRo13WNKC3LPvEBGfkCyVjR4FU+Wc
Aoex+nRJ7PI0tMXqhvd2fEZ1HyMhQB1oRxCrjWftkZk6VU/VvDcyUPCG5+gcK220y6TW3r4A1ERx
UhTyNNG/HCr4/oJArMrt4D3qWWcK9BqeEZmYm5Nt3tyTbfp1a3fmUJgAoEy8i2laPN1m3tWsN0iL
xMzr0kessACnOtHjR3R7t/2h3ko7YDMSiKJIXp2lyLB6KoJiTTM70OkWAK8Opn1iq3vjrE37AbEl
DIVOINkXcwsLZ+wEKrvm3AERTrmNA1IeqLOitYbfb5HIq3L5t6jblw+SbC56cckbLtALsKTp14XS
LQa1KANCcWPFIOHafTLW957+LIO4YwT/Iu0eTiX8cRssCTZe5k0W++W3wTbDtdjSggh4Um9Ha1Dt
KtKckB82PdKJnD/tgT/wE151TzNexZ5I5GTb96ii1QlBC7RWSbNiMItnjTW4rkaGZvlqJmtvVMCV
mU3FBAF2MY+HrawY/WQKrJPYaK5HDdjUEisQPF4lilNsWYfqnaCH7wKkMIIn5thr1lffpCRn4MUf
5kRUgnTZ8OBqI2EV36HVUCHHHtx3xBDTJeBv7IJhIVJ7VPdnSB18JnZnwchmNG0fxBgGj88I/ObB
sQiipnDavDnTCrPGrhThosVe5JNZ4mFkvLkQmt3ekAEiHzYzHKofr/sfE0yze3n4vPs2dlR1VNaY
0f1QxkG45uFJ8MCnyZr3L5R15Tp/9y/pkAjdPVfCihm6ro/BJjIqcs1nPp9T/PJMEIX0eSu7kTmT
tV5G2B8Jdfzvc7YLsqwiyjOeOGh8PGEcZAcS1cQj1SSuRA/CJDoF9ksIpQG7Y0e/86UgQnzi2vV5
2XAQwhGXp5JU6LT7D44OFaUjZ2/b8B2hSX9CW8644blFyeoca6bMp9XcC7q1Z66CTM5hrg3WTmjt
ls/4oR6zNGxtzdLC2Xd2k5ERuinpXUfwr1goaoDu3gR52rP9H9c+xde61rbOCexTAb42eG9ThVJr
+5RssBTv/m599+MuG6qEt+ZlDqhaxXgt8Cin60DnfDLC++Ud1/+8E1KziCOpOIVJc6htqeL4VEv0
9Yp8tJ+WA12kFyo7jm9oY5iijzgbU+wLaim3dGFwJDw21neVA/nECVwQ7SKHQR3jQjAzGVqQQftU
uSPyD2m4H/dCH1sbskgn/9ddkNyRwGZ4zbMXeMtS/LQS51SaK+dr+hQfLPTfbNTfldvUfxlfLBg5
Z3GZUj4FJYYROVIGdzRu+0i7PyLMiDKVhe/hCrrTZxdjkwkvEtswLT0l9WJgBPLluR5lSHv33/le
AK5agHv5aCFSrk/zodHqD9/Yy9CJKlyMwvnT1U/k2BeUSA8SrxoCbERlBjzXlG/lRYMLlT8nfwxk
OCvBeQCyEraDuTksry4J+Fez8BQhrAs11y7qdP0PkDwY0b4flgeD2ApBqIqx1KX3Lr9iKWalpUMB
cR06JOl7lXjTLO0+u0sRU7gu8ZUwVPLhKrEhgTgah/gP53HeN9VuLH7hKzF5eYDYXznx+9RDhYr6
2JcgZzIN1FlD8+vs3c7996GUUkbE9x9qCtmeG9Y+u5ZSUS1Ak93JIuaK4VYuBXeXOS3D8Gi/1d4e
bGB01CHicVVSu0+fQoDepPGHSYm/cH+53J0bMSx8FtIMGUFea/QWZNWetHZzXFrfLi/0rNh/NeFW
JnqfoH3TlAByL55K93AsybD8atb+ZGS0eMXPH2wXDKpdODWRqxEd385QvPxjzRNm/QZMQQVC+rbx
Lo6a9lP9acDNYDTw6OVSfYyJxXm1tjvdOLHv1fnXJWMZ+6zG/VNp727qiBkNo71SkWCKcvvfnnrq
O20RBk3ctyf4Dn+VhWFDTYQF3xu2e4n1Thq2bj2lDlOqEw7AT2BfYYRo8uKx5g/mhOGh4Y3FpV0E
ha1xhKMWGX0svU9DP+R7mg/WWHWPI3uflkGqSYOBxLm8W16gfg46eRHRH+zZUPjkr//YTF6tGzLG
VNi4ouuu8QmYvOxCq4grgDAKINIFZ++Crmc2xsEVk4ZYvb4uPaIFfE891FahkroWfCGboXzZu98E
p3GToAn+CxKzNF8PGrpTBJrgvUf3mlJhjd9QEQNbxfJ+L0UTV4Cw1k+KIc6kD9QOzPLBt8+sqagj
xT2L4iKWM8qSuTAE2xYV7b+tVN86D2j+nNTxAqxaKN8zcKe3aNo1JGYCReNQ5PB2VhdyfT5jp0Gr
5sEoCihm3okoZ6FFkvYfiCgVJKNWrgaeEQFA3pmwpvLdnHYaLahsMKY2wSSR6T1hEEJ7P5NGhPMw
VnkuozleWrUtueM8T+6JINY0m9pKVl1Iy24MfRli8+RgzGMfKa63t+VPih2cmnqnJbtQb2dc4Gjp
I9lLUoNEiYgpW4n9BOUY155pmoXBao7obfI78lLiSdmxScwimUZicBk7HcGQXEpjskxFfscEhL1B
B8AOEAtzdMgJzoE3nQw6N/s28MF27HjbR7cF5Tl1irVk3pcYjhvARa8rUmAu+s1bUzxbWyB5Njap
y8b91voZvVToYla3qoOsOsbMV467+DzzmEpcoDE1hj7fLZOJwElSVr/nyWtSDtlAyNsDd6yDomCT
wZULWgiUoxhpWNwPsRcuRnHbPuBWBy466cahK/lRTrXzNwlacrl+ZdZt1TdjB8HLjYZUuMq7601I
duR8lrahz//vKsIVCIq5nCSb5E5AlXZ/HsWUxXPQEQcWndSpDg0DtNLrs0CKGoyWL5ylKb/oG68R
oKWXjP/rX2JfTNogKrokdbABKdt/vKN53s7gjqkm3PaJduSWYrdRHHBUyCy58qIoYTXBhGS+UNVr
j9GOyOnF5si31Qr4v8RabZMt6PadChS/x5MdDamU28ZtUduNiVZCim6tl5zTaHZxiXDmtAGd/0kY
255C9QF4KsPll3Vxc/QTgU/SIuwXKjZgSB5SIE89nl/tSX7/gI6mJpSGOsNg7iRYjtbONJzQ38Zo
l7u0zcHR042Xo64pJCv4gT1NROFe15nrPttVBIVgzKJMMr0v2pGd/a0ryQ9POT5F9knDTUxVchZh
LKNsdLB2tquT18zysJbK6u5vxdi6J52gN2il0tPKHxtF5jhOOrRTPPjT2+Pugtjij6OSntQaN2XT
Ay5U0gGoPbDApQqf9YbHZlMaeYzCRWcsvuDeivtnEapJJ81jAH0CB8gULQ3ITEjTs0bAnDlzlRb9
k1/9u5UalsngMmY9JuQQCgv0hfaXjr+cXGJFX4BjSNRhsztBTltR8G1KhsPVfcJQdEOfKVRLsm9l
KtTPDiu+ycDZD2mTw5xGvNG6LcEH9hmlRzZmTtivE2PFVk40LgMM4R558RLzVpHkNucF6YONtq5w
GDH/xzGK82UQybrw+TAUK+nHzzavomMIgDz9hgakukYy/6QS9+GmTuQiFVgJflgmPv3UtNDTFpjr
66HhbINOzz5K2M9Votexo5+dgU2JNzol3jXdS0V31AsGaWLYGMNYKwxuhkqeMTXCbKo3TZEtijbg
viwJK92QMeCOu0QLVgaw8qeORt5N18hZU3Z76xrM7wSTKR0iLYGGV2t00yEVW23bUMtjjCX36fHI
dV0QDO6N7zH+Gsbg8fWVrsbiWUY30RaNL2YGqxv8FXhiBkLe1voN2YssDa2ctbPefEQPoFSqTi7c
UIZW5z441I/xS3WGHVywUCM3SObM4FEL7v9kFUidm1goiEEeEEIU0VAWnU/88AF3ZFtyVknn/pv5
mJC3EysU2p3g9GHtWL0k/b5m4B/Odl5xKqyUzXJ1Rx0elksyX3agP7MsSZQUT0kPCRe+61RIrtJp
kOyhCnZbVOhz2xsaFNgFUoeYjnPiEFTwFbrzqn9WdXa/EXTyv6n7cVJubawFvdtTG9yxcaUVubbD
kYgkuif6ao+IsheadH8k5qgnEJGaMOJ5cezFTB2EVh2/97t/qJXoXKtIjm5WNhA7ripzHnttjHHD
qu++VzH7ydpPJJhP/dIYdG6iRTRmprzsePLGxasd0qzslU94H9jQ3BTHiFspjUhdbUaAA2khTOAx
YJEkyGNzMYaU7J7LbEIxkyYsHfRUN67oeYCyjkttiD0/u7LPbgQ4b/wRizzaZXACRKKx9N6DuCG/
kqys4EEwtxLPQgWk/RUaKnNQ2S2ZPduNHQl1s8nGIiX80kNF4fW+zVGhO/kOWvjDm0bJ1J5//ALz
XIfHI215nYRHZnk8s9JhyKH3PxzNyv9ebBeZBpC+WBT5qOKM8HCV1+fy4S8ecSc2UKWKrmoplTqT
EmIFvhueQiZL8huZukd60ZUAxFs/6Is1+t1voD/eYUFxnnTEYuAI1glrZIvifiXSvnA6pd8FHLc+
l7JriQ8Ag29xxCHcnDn+2gIgWTlXiN+3K1tqA6Ec8kma7nsVjHQhXmEMy1IKLDk6fPDLp0qCh1YV
LfByqdRtEE5noUcR6d7uzp5nDm4fR6Qib+lnT/tdbVV35+6zW7631eIWyaWIk5liaO7NH4IHjaMT
FG1qtcWmyMTXpJTmq+vquE35v1ridmyERZPmFccumOjjt0bvol44cKF2MfceT9g3adFPIuRRlF7P
lNejWZW4O+TT87UnGRBALnrdU894QsNvN40/47Ah6j6hhFd8DNHkL9XUU6LgmRGyXHlPXTj6VbWp
HSaq0rQ2Ro6VVN2bwta98QPKOApEDmPvoUTF2A8wr3x4AkocjVR08x4MOPgVhB+d0DCjRHf/INTT
fPVYlyVdTbgmselsImw9s3g9VKs5Dya/xLiQmQvgMrbSe+IV3hlrXUa63002qyDqTDlBxLUgpG5w
r7d8jNecpV9KmdaJQBo/GPOIHVIgHNCQeXEhy/EshWk6uWvhLoNEFaXVYKjM+mclCWtOS6RdbIkd
X3J6g3+ioGlTfjQxXltj1Txm3KyCPFHLv+umDTt0/JhvWI0bVefrR5wxnhZyVjcUVBr8qa2z1U0J
GdYcWLG9WxLuQEuLdco8fqG0j4/gD8VDJqvmii1+RTGKtuZxXQQ7sNQ7CW+tKHqUVYmgPt5lkoVu
pWOq1Q0fOmnG28eneb2pnJqEho8MUDZKwWPJKArSUe6R+VTQY7H5FUFZrKZ8iB4PMHbPWwCAGzwA
kG6acL+ub6REe+uIWl5ii/sfhhj4+3VOHM2y3/YejkEmYyI47wppaGEp9CDo7F2Tebgu7r7w6Kbn
qF2/OzzBTd/IX7H5qgmUSjw5pX+6Uob3Dy+s8FCnnEZic1nQ07/oZ4rKk861zdRiuJsUas62juSx
Xs1/NAqI0s/jem8WUiYc6ak0bWRQEyt/dVvRwQB4tk76LMf3WvxeDOquK5x9PPg9jE8BZz1A+nmr
rDYGbs9THAPPUPTRsn0tZK4ocCERD7rA1UzR2837iaDRUxB/TPDPA/Xi3N0MrKgwxiU2RQ/7V62X
Fgkpz8J2xlg4p3LTkmhLJWIbnpiF+LKG7i1ufAvsHm2EPqXAtal6T3WK2EFjE7tkcPmM7A+/75/H
f73pM5HWJ+9ZQ5TkbG64q5RxTBbEJsNtluEvIobxvmTI4tRPnwdQeqa8PH/EwuAFjX4W/vZiIEYl
p3u9H5s6XGDW33V50HE3YEC/lUuqcM1/qpS5MI8aiug4nKkacFR4nsLwwHJpgZXnG7iD6BIjDjpu
ujxHzZ2emPszZD7+L7apjzGXDA5VFjNcNEwXD2tK+Np/lD2uT/G+b31G/wkWi5euHJdCg2YiIx62
3y0eQrB57sVclQSg4LtvoP0kKmiaOc4+1+rmgH68nsYcnkfJjDPW9cV9fuiL5QA95GFS2AfpZ1sn
vcXfrnZu+2lEyyf4SepBv0xrQINQkNjvFa7NRLNO2rl8rpIj64EzB/mmrzIFxNxjFNWcUcoyXs9T
JA347rNsxvIKojduGbBMBlSZVPOHaqbTSMIFJ3ZxsYuS3R6rEk+G/O285a/6XFZRp5a3HWrLqajD
CYfd4hna+AlM/ApIUSmtE/Jt2Yn7Px68sAjDbupb6Wv6pJv5OhofKOyOb/CGoftc6z4M3gmAqudR
5V9LnyCGujwq3XAlZTAjXUP2oTx8icwDh6s5stcOccRKsKpnZqTkE0fTazI2hynx/NGBku6lZiz3
7oGRoYGs1z6wW7Td2pAykWFcFfqBaVi5TANxkyLTCVqmwz6g8eUOOA/bCgD2rXC+llSTs2AQRLl7
A4FVcm7D2Cm/+Q1tjAhlqp+Sq99ozvgiCvoraxW49avRPukjSEbY+l06l4M27aHJ8faCQBGCur+6
RU567yVKHb5MjQ3uw3kjBah8TFQH7yJznLOBWTN9c7Ireb372NE0WyCfRrFlMlNVrTk49P+Vi98A
AhgFZ4xsbssa/hr9tCLI0Q2lkX1T0g6ZdtBIO7LJwFv6zRoLKmI8uPWf6YL8g9NeVpVPiachkcIr
hAxzEV5lzfmB0m5s629Q73KItQaReU9d25YUjoREZnqj60MNE1i/GBc+TcvOPquo645SmCn9BmSt
dzL8XXOW3A/O47cTH3Rg5xbkpIUQzmktg8EWIOuWpihMrwP3PX4fRz9+nwHpN6vxXwCY7MUgJMZ6
YaAK3OnEv0STyqb04bmF68VF5JnnSq7x2ax0v2S+hKqew6FIpkDw776DDdJSPfg64YBWUm67W7zX
Vj3D8yYfrg3IsgonjdxzH9QoEhVPJCgaKb7kqFgVVG0D7aOIDO9pbzNKSmLi9PaoXes8LndxKIge
qRUIGLDPNYI1LyiCAJc1Z2USbalaBGTwDyzunFWaOJkdg6ZatCdKdQY9FjodcXtLlfJ4KX1nUXjf
LyyqQEXS6g7UBr8nXAwzXs7HfWgdKi+hBgMGPtkGTG74OObYBc5aD1tY4iqoM8Xa4amxeY34dRwp
Uc257KRxa4j9q4K9PJCxBketW/ZxlT8G8uvgmVamUVXzOKNQVtkTmxewWBArmJFCyhMYrTfeiXYl
4Zj8uECNv0iEkXoHZCAqnlYuDuSsXECC279YeoJEj1ONjrTw4WIPfVBeW+RC3MdRJDzMZhshG6Ns
sOo9rz0p/7HjP/094drGTQllPU3xxCojkjxexXYBP7gY+vu3DRml2a5lX5shjRiAd+bV/73g0UWe
JpZEh5NRBP8Q1HblS16SpCZdiKOP71zH0AiwAI6FOVtsXqxhEoAkjRVsmpt7PN8V8obtJgOVrCRJ
fF2FZBsh3gx4GYg0UCwluVSyQ9+VoZoegPQJGYHqOfrap1zJYTOlQSGINFOfgOmBHCBEVakteaWQ
XmzeUmC/7pXwXlQn6HZkyDQyhDyOLSIhZXd0sylBaAE17w7NNI1ev6+MLqgOSz26PzN+/n+pL6Y9
tYN3ueggY8CtlEndXF0IVhpVrkaoLtrf3DpCJE2lpox7wY1oQo5iPzPnJg1HftF677nWVyV35IDT
iqBtdX/DxYBLInPxAjPHGlZdvj/nn7O97cf8vpbVy6qcuVtZTsyrrUxqA2us6cd0vkOEvwUtRsQp
3K5VXT4Aok2qrEu4l1jxRgKyR5BwU2AQYLAHUsmij0stYBhAs4ap+Y5nMTTPMsibN1YF3/C/egsh
vXcDQD3dUV7Eo7+W2QbFuAIP8/5jE6uYiOZ6XSAQnGFD2exFqZNWGbfcEMK9v7LnbPadaivye598
aqaMRU1IOqu1wk8UUL63ZkUmp9FZ+BtQ4Mo43Ci/e6SqS2MJ7Fc8FW0dY/yPVfE9ba5Xmfx+6UYY
U+AwAjkcBTUeXsKZwj7aHlBo7oA2z74mClYwkcktTOQ+IzOGeMVmcQNYoO61ZEUJS06QsmmMDnEh
XH6kAGebTy0qauN384/C7+xHBhRtNjRl6NDfVEcfxHzoGEv3521Dhv9F1zzoTsYPwo0kEw30EwQW
/2CHP9uAajcsVJALaB7rxLvfMLCwV+VPIyWLHcG4BSEDVi4RV0/KbZh/J43hisBrl4UAanILgRpG
zGq6GRWOsT2kSXetwUBWqVYIxhEUXqO26PhFLeKSXgP1ReaLvGjTqOn1eVHfkjZtzsTgbHzACO89
hQne4bc3Eiffad5ktBlNxnCG+zTUFcqGJ70Y8rHKdkzUMelmQAnCevGQJ9S+AGkafB2ZBImld2jI
dcKCKX+YZpgajqcnAvq2RNxWl8719S3wD7iMZGc1IWsX+b+IYT4mMhIM1UzHvehATBtXOA0wDGs7
D3v6GtPnLX+KrfflQahshaRcWmb1Jn4fOcLFBg0jgzIiFCvVkYwr6L0bG88bC4yEGJndfMuyNTKI
3OiT5MldnL06naRXPkvHI2KFkXontfAPBpH+1TZv5lFTO2PKvVJy44TXDuKWFbgcp4GjgJ3Sk9kO
9fsItvzPsvLcMqiNEncprKFxxjB4syWkVKqcCwConiywZBYODwm64VQD54tLQJMtz0/7DU0Tx2hQ
/bvvGghKXhvjo5sXIWU/LlcoyipoQcqCdWlJ+WZ/aU9TO+eRb234kHZ+G5BwrWAv3i0quAENpw77
j+9q8cFz+d+12yITTwLaubtxgRqQoBrc/+2hIG4wYCB/kARuQvXdkwe5fHa1Sbhn+2AImFQfZL01
p5ayPzk7bIH1DyRgEcz4kHdWliFid30Hkj1fYxpf4YPnCB8t69ZWTfZbJzsKQspOI38wj5moLCRI
9pKWFpE0fl8GC0M6quT2A2Lc0FDv+H5iiJawGQkE+QT6RBYX1nQLk9iXR0Qlk5TivW0bWUO4Qu3O
MeNhVQviOYKTov1sJqWAmzM6sXEZldX79lZjm39bCf0P81UcH42p/JKvRwM/K+4uvn4bTRJU2Eco
ZEMzYrT5EoFoxlTIz9KAFj+IEtc1GRinx+P05CNqfv4IMMxfd3PGkuVIR1Sw7qu2KMB6ph2EOF+A
KLM0cwHrKNvoBSDxglXsewdxI6G9qY7mVO44il4Cq6KZ/n4XYPzXrumF/QmqTxQ9IO9jmwap0OL8
VoOgkP5xqGY7p1U33MVEzd2/nSVE46gguA8N/dYDPU8Q3QL9FE4QoURA4b5YoKXbvs0WvB64bkj9
zci5njlnqdxn/as2b1sIsYEtC+4ltIyR/tJa1lCTl1eAekErIo9t9fP8PW8C6Y10rT5OUu3195IX
dFMX+5r9q02D+qaVoTo0fOkpJ1ObkQuaKtHbJQ1JQvHvtYrERomN2aRfAsfdFoKR8HnkDisAkYT1
Gz7+gpPpbXhC6ySE9cB7dCPffcnZfY17faTmF+UTgqNSDOCZsfSLdCLq49xF8ZxY5tkYD0kIn12f
zh4SMeHzpoG57NG0s2/k3NQdyf8qwjv9eN5CvGxob7iQgPZxXPTlkQm08NuPqBEVMXaTrSkDwvda
3UAaWL8tRbl0rvrin9ndcImSILzK/S8cs7kMbqZPnC+KpNX3QfUIA3vA2e46rFXFl3PFfC47K5Yf
Jxvjiky1bHyCTxbuEELoYs18NcvNojmrZ+0X7xJNJYRkwBL7i/LaN3tEqZXiRcmyxBEkxSTIjcL1
XmYnXB+I80++vFnR0aVQSHj+4B58JCM8MiM1oii4fFPIuHWqfdCB48ok9wqa+KAKM7GSYaXtOgv/
p/v/jhBpgupJ7fElyA2esKRYid9Dqu25KLZ7dY/BMO0BvdiZWUGT4sZTMsxyXJ6fZSs00J1OB95h
JcFqjESLABLMDIzi9xX2WMpA4Me6YnKFlZ1fA0dlm1+OSjXqEBR82ubEsBTzIwhnXPVrAi3kn5cP
uACWDnauRtgO98mJFV7EbxtoaE+zrPyZLxM0rKHn0ke+ycFba7nwm0tnvEcPJH2w8g1MlfWmmZu+
qW7RZxK3KhfqYWcLt1K/BqqqyhqrV0+vjYEE6hbuxFI4FOTBKFbi7PnudETOqMeejtlLKeDmWEUu
djplo7bW440nUz5btRy2DGProl3+79Adu9bZzyQiNtcsyA0RY8eXw7BnswuVPs0Cuv6AtPZyg7QP
bBImJOUjQeveRGheJA9P3d9UG6mp9wT9FgTvGb/pzjyPqrP/6Ky+8d+fjrRm3KIPh6NRChpGq3J0
MtIrqX4ZV8UjlGZ2DCGUtaYp2Y/G3mYRTfrMcLs1KHMUTzpxcDvbk1Bd7aRMutKkGxRJoqoPhaeK
aulAsbuUaKn1ickXaH4m0455773dG9n5v5KvOIuMv+L8RxhG7n2xJSxuEWrgLDaRGAocJXokfW1x
ca7XexkzrZSRxy7pTB08+WZYztiC8ySD/xUh453jxRjehgAToZOVjvq3I3OkgPoC1P+zsOkParwO
w1kGrcje3E5C6BUBcXE8CkJZXgMgNDlV9lu779heEx148uwHlwTqTCHySk73thqttMbcBWrv9ZRj
yLyEBYM+fDlmXh0D0dumJSKbXKFhhlfmFJWVZoGOqY46Q8sDuosY9o28e5GNzGT2g0KSbGcEWRD1
2MU2DjJPed4WmfdgC0MaWE1aCrSBHodkPnY5uFruPXGG9FngQkflrVQWBxWyn+II7IMEUPm55+cZ
qbUTNIr28SqpS51D/wBX4TekI1GXJrujlHxwiSCX9AYkzbJglejWIHCYS0hMI8FZXWFPQG+tcKuJ
4dEchpGVywm0fX/JBBRBarivHpyn3pttS488P+YxHJ+WxMdQUvbZzLv70d1hLyjVMbZqj7vA8u+5
VqZUqp1GAAqjLKDyO8MJ0qZ6rR61SVsNff5GPMpeHUPk727xSp/HwFvy2yRlcPebFh+gzgqhT1Ir
SWZW4xMO+XtAAdK11bgx8dwyPINDyn4MFZfNLTqu4x/O+BTpLb1Ni1h+KjXaHgwUKti8HYJur+BO
43TPsldwmwJw3mby3yFbAhTaAuW+gozYjLsgWTImxzrsu+fjS4phfic+SE32M5xSRjf91LOIU8Mu
lHJLSY7aonKbalsD7WWzeigvoVTN+KMnK9jzMYbkicAyafs4d+j1C7ODZW8z2xmXcugODmTdQOqK
yMfLR+NNRI6HqzvjPOc0Z7k/vvMqe6+6V11wIlZQYGgR3/wM/q0e429G1OCuJCkSLjodMr/cKia1
SYCvjS5xHT+N+EW//f2eQyp7pcOoG7/XuWoAQBXVmLVW+278T+8fb2OT3oqU65P/2EyEw5gHZx4M
YYMB2RdOqYy8umYqu4m0BHTUPdkKX+wY600HYxxe/I4q/qrJg+Jx3e0aFs4HdgdHUA5Al3UQFG7+
Ll5K6i3S37H3dXo6yaokas4tXq22bUpfQqNU3BkXk60xXr2yqsTbOziSm1M420tm16icaAiYtf0U
Lv+3PVYe63RdZ1hHoDJNYoCz4AvvhiT64sGEOTyWPwGwd7TL1Ug/xT1XsTAQD9M4Ss9PNmffPEDF
xvOd9nwsrSOKfkt6GbiW8+F5PtYmXOisatCLotXEG/u0RIruNPT3wCgcSwQAyVx0gzuh5fXIjqgn
iMdTeLtVEkyGBgnY3HOj2nP2Mv91J9x0EkPAZwH7BVl0joRa/2RGAAyMbV9A8lAO+T2ZpLiDHK2H
c9QZm2owCnzaybXhFD2a+bSchLvGpaIFhvIwmzhNPvifs21/uaIA8AS3uNxxWQSefEEJI9weQAl/
+gGWA7maYD4GyELXkLVxQ3T2T24IKQ2EAn+S7Eis0SJfarKU75PxxcebfGygwUXzqDGtkJOo2CF1
c2ae2uJGarJzgohjKz9U/bmmmGEtW4JUsaKJTuhkKdPfMmu81tYK+KpPikkw8u8JEBOuytGQPpg6
1JcNcvTTH5goR6XsU1fbt6D81Bz0HKibI0VxuiNw9/Nt1O2X+8I6PVrWYZr2udNESpIG1nZqTGNS
ADTmyRCVhg01Cebe2Vp6VJxXds/4rwpsa7cf3OTGdxb14fR5J7x3uSDBOoMhQsjzy7m0svo2vX4O
mXjtnpA9Z3fb4RfLOA6LTv2qyumcDeWeQb1vBRed7toeeGSzvQ6KadYSw8LqLnlqwtWe7S404guA
iihnUEn2+K6v7NIS9d0Dq1zXkKxmvWeTwzkm/XmounvDhRxKg4ABYzN0GQMbpIRX8zzmP1cfZdZG
t4da2lMT4c2/CiBX6vFZTldqJwUXRczBArJzNO0exm62Fqe+eG486wDtT9L+qIvi8O1usqbM4o1k
i8h5sPutp/oRpYde0zlrv/uNE7raisl//XCo2r1MgcCpML7SvU5W7ld2/n9D57hN3HrwdaNh0wCP
MOrSU2A9mNSeJNokOH/ubXOtD0EsMlJyx8f7D5NQimP20g69TZS41Pk3BIvCfcqtNnt7rWxGMq53
ZvokAPX+tWn1rjr3SXB4xMO5jJqMB/+CPSDGqJbKcL2VmNXNnqQJwa8W4/EaPGPkbZpT6TYFFWAX
/YKQY/UEAgCgwCEs9f9AaOx8hsgakvjJ3h79h1OwbLhYdBGNFn0XuPcYxVl9eU811ssLl1N4bfvI
XkqctCNhbslHba8yePnDabthoFhHt/r87PJeEDkENZq6N6Emx6Kj7fs8PDZ9nVsatVtiE+nNnWY+
eKM9KnFK++wXWwYK66Eg51fbIC0B1EJj8BcSciSW4Cf8HfjlFVT28PHYMgmhgV4hQXeNb+M9B2rI
4sf070BRkhyoSiD+7yD2mVEZjcfkMTymhnCDzA4oj75yECYwnTzccecHiBqWqqfmlALi+XQQlRvj
Z98zFeZGkaIViiKh2AJ0SoeCDqloAL7IAp+2YiMWYXO4cwedmoWVvJYbliuGyzjb3ZOKmtn+01I7
ar8jkCqzv1x9igMavt6aCAjRpjeqZ79jh+AxdoGyID5bcDC/Wq7B/tS73Mto4iEeRG4hXdWacr8P
jwYN4HWARC0GjShg2nnfbGj9gc5owWQrh9ztoDK+SkJfNmlK2xAlJpSAJSqDQEgMoo6qzCmTZHwe
5P+rmqSKNm8kUbErrhYNlu1c/DFOAXyrRR3k/2q2AANe64vAQV8f4YT5jzrli3KV7jJq+VxtaTpc
+5PX8nc8P5axaA4/nntSVkgzi+SsrvHp6B1IDr3bA84qJ3lIauRlESf2NwwNitbi8zjrtgohUDR1
It2iYIPVxksDJHAUZKPHm8EtzMNZgIcDV3y9Ky7/iNd2zpvaEeLUZPahRCMMW9fSRRyzvU4TQf5Z
1hLt9NWtE7qhDtO+OU5nrr1s0Dcoz68aYtibYK1fElmD9XPP2FsbqbyBfGMtyvmUeWyZX6LOYKTk
ab/OKC8r/kAQO1dBLmM08HreZNW+g/Ldvf85n2Uo3GyoNKmwZVM3y6A2COlBamqxwzvjeBH5I6Yc
UNbsirhJnJCcu1Clz/yY57w1N406X58rLQEbKCwDnvISak7j3OL8NVu9Z25Qvp2RaHVox7dZlQqY
15mKPude9nLBaNj25xo0VpqgSFYQq2CkYQb9oa2exhPMO5vOi9CKZhg/sHNYTOvP0lFXcXMbIHnJ
AxdCwrS4UX/NIJ9t6i2fcnKX2q8Knl23XjcPRsnWExJbMu6710RUF8CfIUdmbVvu6gi/CmKog6dw
3jE5RRqGjsijnm7KZNAZxI0tejgp7Rl62g4ilDp9EYvQD68gpiimBpviYyfW0tdMMxGVP66YYTTE
/C3jR5OPg3yqv9jMT6611xQpJxg6OM+K1cojeAIJ88Ey75vRThG7hpC7F7eZqRdzlmj6n08Pt71t
yoZFV7vA/sbxnxBsTEXiCNr/ZCpGArNkYuGxQuQnZSlz5jIyD8UGnVwwcn/8PdZHk33ukvXMpQY/
MObFgtWyRs4rsNQ0q96esISX3ljyv1n465oxwgjlktNx5Iba+mP4OOT8CWGFp+kJ+GSiB+Q8UWDA
6HMCvF+o+ChDB87tOHc74v7qywkemgmW8QGibfVjv+1Ngl5Jk2h4oqL/2//m/U37gpJ5KXVFE1Pl
7X/YViaI8eqi2CtrVBYri0WuGDGtHt0Uu7oBBkeEVtTGS2QLJVqNtRQKD/vbU8PsvQnNqWqxFYmG
45cVjdJpPOxwapCnGY3OY4ZmKUZWSnXybe7u23YfhQbf+H8ntUF0Uh+y348u8wPWoLMpqjDWfnGY
7I48tiV4CeKQHRPFrOQfgmLCXrQq2EaE4akRzGaUZw47dEEuP7cP3yPJ5HFO7Mrsio8w3VwMiZEJ
BeG7P5wJAsX2YuNFdri6wS4hqHHUdltHgYRgiLcJdoDtk+YBHQczqTIn21Rwk5oEZAoq9nMzi524
HHOMisdrv9hoJXLa5tM1XAgWgy5FJ9rqDAbNydRMKGSC+EuXMGoNu1MMHgtSYYjFmoy2UxFT98n4
khU4AGX5L3RRIHaZZcaXx1al6MYiJKCa+Kfq9pu5jgiBt6FnDxCXg/8WNcZU2o2a4JoC8N7uB/Qi
TO+Qo9Nd68PLafyMnMFuxLQFv+KQH/aQXguy/q4PjqcNEWwRgcfwOmElL4FWLPqf4qLRcDGG8E7K
6iBDQcgXMyUozfOdgunCJuIw4QWvJhaFIqEKE5VLAgdPHuQGKq3MQv99/5pABlfIYx+eJsgMH5Zv
xSGog4DD9FDMpZhpjazPQxKNAnU+xWyoW/IREMixDePBHobZ2n3YireUqDvW+YMvZriGiXsxiEMY
NNwnzL+MkJfN7aiNImOtyvLGPMm+uFGa6zBss3RiiPh7t3ihrlTr8rbIyeLtrlQZrTeKgvbwl/ol
meBBd91G3uLlCSmvMAYOa8qmMQN0SAP23kK2uFLy3cW4h0PBxKixMs0kP8u6y/aYNGbUpCFbchu+
IpnxhlN0356hG0obdfamMkUT5D4om+2wQx0yrWsCfc9KLmwp0eCal7vt+ZilklaKT7I35c3PMAR/
33J3P7QRRbI8/BNYJW+lC66vegb0EBIhkH8/rUD8HLQLms3h2bJQxP/GP8YzEQHUStW0/H2Bgvfg
EzZyTIZpjqlc0QUMFpaRyHE0Ndqt9qI6g6f7c64QCaXC7HwFSrP8m7jEWSbQqyUJxgHOmxkGExiF
+EJo6VOuBvt34awOiuTy6hZTWPWpMSzupAdhemrNHRmZVOTNgwXBDLRuNjHAJrdgiPrexUQ3yCnF
gu6VYk+fZVYwvwDWxQv3q9USYJrdsxyDDBF+loa+Csw+HOgxmRg5JVF07mRzpXiRtrXPFXBHy7td
q7o6VJYykbBDk+65VPVKHzPB/WAp3ahnLdu/qsOp/l0kmiYLOEe8gi7P01Q6IyrbC5F2y3d/H1nq
FLYC2BbZubmjeM0w/p4kEi9q5BenlMRQ+2cjC4FBVAIPpGh9FSV1WrLc91N71Yu0It0sjtBBTQMC
RRYmi5G0sXqUqY4DwFqBDXUn3dpDPt9qYN4D2Em5rcNYkB5c2TIoWcNMN22lxA0PTZvDvpFpc8Gp
kWK/HZDcQIOJ+dz1tRp5awdQFVHADdKWriajt8ifl2zXOyq11mAxUR/jouyOXsA9Fn9WF4GPlbTm
YdOkmnBgSZaBuQSibQM2Uyff/QNAyNpxX0wV1ZpMpivKrQcmWMvLMbA8FD09sSHx3w/1mBoD4IWl
lo6jeLpFZQDiEuLjqMljL0Cg/qkeYnyMl17wj87rhdq4jC7WGzuvZPvoUZkTNyaFL3i4tdwIpEvP
FV7OWuRlwbecFcbeQk8c4IA59QxSb0NiiRr64gl4ejYgeMHzaaQecgqkV2LWXLqBaPKq/IJeO2Xb
KqlyJNNBW3uFC1shIjR4BJg+hj84A770Yde7JfRrgAXCT/iew5qLSf//13pzhLjJ8P/boGgxH6Cj
3s3O68RPXTOYWMbJRZY5IMO0xtGOm1rwf44geOD6ys1h7IOJTf3Z4hSbpf05l5MrR1Qjitj5uX3e
BJIk/ODBXddB9b41RxV4Dm0dLXyIUiocICI6WQnrZda5n5VptMwMGE4OgGlEWpb6LvxLACscGyTb
dUsG7IrIUv7vw5jJCgmcu7gq57VZkuK9ueY34nVc5LjZtO5zd1ei3gKj9ZaYGXMIsN45A0cTZxXq
QpLzRtS50CeJCIlcuJrB6WF9jPHKPbhs0CnyyQ0vOSeeusk2ceB+B8qaXWtciG4Tunw0CuvbNI4s
dFR+NfnQq6IbMl8DjdrCW2WZAHSumL4zrHDD/qMxksYVWRuyUSFr9SAQtCmsjKU3qfoV51/IhThz
2mOClq6o44iHG5kPsAlePpgNP0z3AHFQWH5pSQL9F0RP4xGLFGm/nUG8JrYZtWNshivrDb8+Lamg
mS7eTdlbckO2mHGMkK44N8Y8fWUqm+Tpye7mNCyNcfhhq4H7BiKSCrEahaB0EBY6k99kHPEaP7PW
kiFbOuja/0W40YeaEMFYfGdV2MJ7qUrHo0EFcblcVyzYnMkp5Lq0RqaUmUOB1BoeyYUdl4MJb1Tx
XjFsduNeOk4JOLtIFxBUOIzylkhFrjfkCVlvwDVv1BL8+9mu4ZHTDZF3/odbc0MNNCCiE65BjFlV
IPORpHDGJPYMOYqxx1YFsA8soqAlaRLiQpEBt4Ya2BYDeqaalAJ4APgdKL21fa5KJWOOaB9H4c3v
FCxsXy/ICb4Ywy+CjPQQAFdIbnsUXhMS2JuG2zB2Zae3Ecl1KS4RYS+WgItXHPJ2jswjtw/YLS04
8IKetZZJKOhaDQRAP75o0aHWnQCCyrZ5XZ22kAbaiyKsVYfei45BYFhvslQbm7RmpjsPbPVr0TPg
Mqz7Xf3fZCIwqyqlxUvw8leWJ/ILxIwypLH65A+zLk4bH2Jp2tEApKGpb3tG+KHKw7Ig+Vy+1fpR
TBmKxupAm351wTcwj4c2iLujyQJ1nG1xQyuoA5B5Qj+u4FHmAW2z0n0rS3Y3hVVxrkPIdBF/sUBh
1wGQ0cPxXbVNigrEk5QOpVyt3XXjSXy6/5QqZrbiASCN2GVMvjm85qFR9AvcjJSowGoEHp4s1vba
qgEyW9OUTqxuxIzKAXRs56fF+/zHChEcs8IAKPdPf1EMg/pC7S8fxLHcZMc0xFPqSca/1OSiUeeD
Y1QSdfFNqUh1TOcLNEUOpuw1ylpOKD0I8xF5rWrFXth4fReMBq00u9SgU82ZzAGQA52F3XgHwV/g
eDwZFqwe8TUgSYsC1rVhPJH6MgW7+WMhBz/ioN4rcKCqbHMs45OgM148AnJLb4xrJ6SHo4iFWHzn
1xdPiy/EjWM9CrAYD8e8Uz7QkFmCHeOTyqyitpPFWOYy9VOrKLeE6h8dG1rCxlMXMofnNzzh1lNJ
1F84IYgPdtEFDiJyRoAjD+aQAJoRJNN1MsOwL/YeL2fDRVavcirPRYVSb9PTekjcLCv3GIqAsT9p
ro1Ng09zGD5m5oYi39Jf/RlZUAyEGh0LgBhkAj/n+FA8TpFA/ebhJqLu5OONOXZNhwKXri6ZjZeF
J52t7tGakfofYaSezymV+7Kf8Hm0zI41PXX4ndAMwNajuqUiq7xXr3OyZqTCHL85jb45zAaDTmZ/
6e+/tDEN5v7Httrf8ZT+BMDNTCUxUWtOgqMwrLMGBx1cF9NRvgEgfdSBe6DtbcjzazswuMgGHTbS
F3J3C8Eei9UaCGjlD4u9l9jv2rE7UVV9KLO6DYUNqYSGiw8/kEjJMB3Mgsy6ahN/eAMj0+E/6+R5
/yooCSb9DhQtRby72Cmf/id88cBKI/USZA7HOPXyjIkNZZ5Auy7IhF5KcI44qiueLjoarUdfZQlr
/lnECnLqPGN75QpvVE/PtKRo7Mi5e5RekFOdY+zZFqnX2wo+sN68MW+rEd/G2R2nM+XHhEQyxGnd
eIRJhF69Hnf5SYOEsdYkXHMLHXjpcmptUzZCf7hEzi/0YgGGJFIQfikGgGDhmUE/1zUum8pxHBZG
qBmjvsCkTje9xrjLQAwUX5sdFgUyVFYNJPBkhyZ5OaH1zAzs7glohk1El2pySdRZIo1LFntRchHG
TbYzBdn/WMxwrhnTx61UzKHhHxwzdd3ywEvzHwcuSF4uYz69v1maq0/OaCLAjRRhFQG/qLrWkPkc
TXyD8xt+J5BJ/Vb79g2ODlD2CIcqTpt6Hsyr0eoSBOo/KbgK5t73OuRWmCwkr5Hb5S6y/1hzS7SY
NKfUe1SFL5VicGkdmGQBIgiFmN3jFtUTQrWk7w8E6WqPl0avs0/DegmWkwc8K4tn88hDxHXvsKH1
Min0q5lq6WkrVTDyV3CeDzcRDrTHqPfFzx9UQY28z1gmJFiN/TFQjzHSTdusG3UTFM1fBDoVIK0q
ESdbpxSNqhlDRKde46z5MteoBxGkC1rzVwX70A5Uyb/gh4qNusVJx+HjNFn/SXrjmxIsAOTow5NO
CIeHStquZPOWd2Qd3Ll5Iz+QVAqiBjFgfilK1NBl9WR6DcU1c4w2TPPu+T4ZDr0GX4d5lDidjIR6
lSXCBy/N229mN2dNgGb/e39xoph7oxr4Ktsj/QRa38BQK7TiQfCXemTx0p1KXtm6bgUpbUH4JFhs
h7YTjN4Z7/pFmBpxCmjmjEC6PdCubmYaqu5NEF3l7h1Ta6PowgajpHc+X5AeNQK/IA4v9sJdkCuH
Fodf83S2+31rthPPD9JR7g3KkFYejtw68LrseiE+/MZcY5ccd81lIlPnbHVC73VC+d31x2er3kbK
JQBlUphB6ZTIPr5Ic5HC4JNlVjjgocvVTxjkaV2LlGE8sUy+6lSF26xCdOO/X/VM1FcYp1AQsrdc
CzUjI1EoNJh7CSYbYotIvDIp7FPwroxhKE0TY55H+9yiuS/zm6hXjuuv63Q/IhKawewfm36zAvo8
/Tuc/osGUxTQfggwfe3y5W+klWd7xYT4aSihBBtyg0PGGSOjrh1G8I8iZiEREsgiqxZETTIfPtUz
HaJfSsVFoEdAw7Tb5KE4g2Qx6cpTh7rtdavdRCXnXSmfeElkCV0U4/kEou53oh+nNAGkMGr0psuf
/IRuZqrIeVadpmB41KNo4sUx/+b9dux+n3acHc1CPx0ZwRM0Z9tPsSWIMHAKmMe6LHvXzz+LCWw6
+c/NixScBS5Eq67Ut8bpcRXhHGp0syFCOBsFMVTPMHgIyE8K67g/0gRRztCTt0gWJ5Rmbw7w/50d
RgCcohNSQh44ecWWmoyEOfq3hA77kQotOpKHvHsvjWaJh9p7zvtaeR2w+p9Vo8rknOSRsr8m4pYD
FC1fKtVOQwINZekUFOStM7Kgg5LkyVQCUDGFQb17CL3Wr1jSxg07MOOdIXDQriJ3XGrQ0OJB6H74
ZdOjYygXXsXvKTnak+TwFScIAX83M6oqf9528as2zTYWbwW5l2bquaevCfR2OQohfRxxXDnsNuxy
4ok2hd8VI0FMyFWqv1NpkEor6AMaSrCGbrBffyIy4h6eBzHplw/0tZj7JioKBE8MmV+k89y1g3Oe
thG8g4GkBT7XeTSKqk8qK8tpCmomopdVNELRBYd5bFYJCEWiu70DKugyXnr9nCyDfZp9vpR5TtM2
scLfOWKp2jAqJ7M7zQwr2yRn/ntlJn+kcO8iixMO4XW5Fm8XBw6gC47vYs0KgWaRTWwDNWhAKxz/
1RqXfYG0Hws3jYQSbD64JohP5YPVzDSdERrgUVLy7ePi1r6OMuLcmwaNl7ixW6wXZ4hHhALAQqUv
DKT0oE7mAGlqBofvJi1Q+8Ku1Zh5NqcPHYvKSb6Y9eJoBdgpE/1Ne9tl3o0ppuiCHWzUIq2/diHQ
vgOxr+PNyDZTZGlCUHNobHdfDkioXk+EGyMn01ImNjJyYu18qqR/pCn9H6FzdDGKU32tXtuVmyBg
hbZiq2WXSJ7nI+qExDGveGyL5eBuuUf1VYBD0YojY32aDQB2NZs5EgXXoPsDHbG3A2xiGPUnmxAy
NmmSbB5HqTxaS/ZnEK29CSSBRPkOP9zPDS/B7VmeXHEowLwSVM/HK9affZimbDJWBy1VhdxncXLV
qTohKm8Y5BC9w7tVqy8blD/raZFxHglUkVtvE3Eb7TD8WQYxdG8+bRJ45OKx1Odkovq0g9veIJRq
+jxK1wePqol9igatl9Wm8LU0TrTnD6GMbmkgZ7TVdF87NNlt5gJXumsnvvEWJJH0lrZ1vEFUZpNP
R7Y6wKlqP53PW4n7KFOX74vkGBKqpFws2Xd5B9OjGKD7Vs48k0E2/7Uy/NAAzTa6z6sG+YkSpebJ
LEQKFNImFa1dPmWKwwKrRRwHk3uiHKHN0sVBxFjuGa1El4B4D0dsvoO4n93dgHqw1XoDt/2GWJBy
zRMnzwomwsR2h2UiRiNlYoeVjWnohyjgEQ/wRWHr8biVzyk73gAwZc1A1DQ7LwXbFnHnoOlTHKh0
nEuK3hBSFY/cONB5nOv/9I+WVjfgZbU6CGSOvxXu64MJyMi8vThu7mjeVraOOzPRA1Yyv8DKxN9n
PmVQTQFhbESKINAIKGRVjgCDVQG4fkBdYumcf232Y8V9AWuXlkfTJZ2iGpgcqiZsB9eIfDIlb2o5
qVxKENjf8+oQkAlrZLKIAaDpVJtUSKX3IXDQrfn5V+JTcGLRx2OPJlc701J7AMM2mMMWKBc5Z4pe
/Td47f24yOKkSAS1NIe2lsUo5/OqTAiqes2HV0/Qau4l4gUm7RydXY9AJB8rvlgnh9sgSGx317+S
tNKLE4DYUdzVROF/b1B0RnPeqWm4W059Zr+QIURh2uCNiDv40dyEmbr9vap1xamDzq9OXVgqmYrW
vnG4p1ysN6wLSSXOdW1SMJ68yFZW+v8Wxr2VQE5TS4c21L6LKb1PfKZ15+2PrnQV76VTVmwA9Jfj
Ae3mepnkYGzklv2sdwc6VU/GNh8YIJYQ5zXuNqAnMV8RDtI7i9pGSC8VHDsXByEw9DdTZxiMpnBY
6O1Rcz9RL2FSbEDOHwS8zugjfLl5dbM9ewcVA2VJexqWj6UqP8eKwCL9Riq6sE3V/7RZK7KwaAo9
pb2ozNz/JZCKmQlV2CnPBVaTYdR3jAd+5dZYj0/ucBXgLI6dAYbK4hXe/IMU/n9bcNHPXjimy/Tv
Zm62xKGhpxfqY8K6N1WeRnagh19o7KiE4vpaSNIeSWp/NvKv1OkmypyTen9Oj5K+HmTY9bp66iB0
L2/dj5P5YcHp/td4c8AtqK1wmNgydCBD3ZPX1td/pZGGqVbFpOyHX5xLzMLQgZ2gFD7hPYrI9kss
Svm75SWN2Rk/uYq0XnzzZnIqRoYYZVb7kWXDpmCJKgisB/ETsQ7NVNqnTB9/ZaEORC8cXTkoFqit
bspb0bQVgJcqxq+sBe365L+ftMFg3yzT4th2EjTeVRvTye6FxvPkjPT9AtsQYkxbpnuTL1/Syx0E
5ZLmUG6p61brIkruny5XBWRWNgkxPj1i9zWlGhjok/0TfoyPbp+NwUr1w32+izRP1JpGA47Xc6H2
7uCHFjqebMRGRooNuTLV8BrAUthL2hNvZHDLmpsJNJDrXiKND6wHTLylDGrO5qmMLNJcLJGHD1Yu
1jjI6n2gWYdnU9d3CqurocHFcmTmilJ30prdoCy7ldIGvENelRIk/g6cCMfqkmI/P62GCZUbp+Tm
iN797ZnT1D8vtinTFNlYyAcbFo4u3wOmEVK9CV2G8PrpkSyV0cYFeKD0RJH2UjQ/N60TkUx3sHf+
h1NnBEhKiT3DELhq9BKa0e9L2b0m/5mpiLsDg5zcnmxb5GNxkB7QclvtBKnvlOW4/DbzRlul6A5N
ptruyyeESWmurFvutPaBiz2ifEWZt7W1DTJUChOPi94dIQrM/5Wm1mMmqiTK7f3YZO4vtJy+ed99
UCncLDmmwP5S6edMLqX0fIYU/gXaYP1IRLjeYTfkZTShh282/E82k4hM/kGfCm/JCvZKWDsr7BD5
2xgyDh9dRFeQaB0s2yNbcENa3HSGdt3cWAAaFK1TkF8ZTqNayFtv04AqlZPHW2klOC3a5T5dZfu9
im1qWZ9Vy6Qm3fgk1L0IhPvLOeMkDNiqsAxe0Vp2k+jgtAfqXLgX8hd2KFyt4iRekSaf+8WoQeQ4
g/mj+gZXmVADFgp3GJtjWLfWOb5TJog5jaubASEjuuKdMq+59VBmPktfpIv63lCJ8AUYmt5UMSEq
HFGM2heraTeLrUlYabScTNAO/DJOdm6ugENNZp45l9Ps6iIkFcuJIQklMm5xl9kf/s6nGMerXpEu
6/8RQhxUzmDnx+m9iobHiFRlgdzHEAxv+Ku9yxAktjqUmxILkua9eXyxMDA0FH4gZwQu4tBxIA92
NahKp0kB9cMDqPd6pBCGz5OvHI1boY24Gt059s1MGgFNveAAWxfhC/l73tQJmubz21Qb01ZxKZjY
b9KVknpVIxIiWftogHvRG6uaS/wbq12b6GRn6eVHH1oZYUQznpM/dIlpkTC56clzSix50XMCBdY3
h1jpmaWSjg7k8022T9LfV84wg+BXT+MULkA4zYKJ4uOLOyO2b02HKCN09FbecXZSTbHovcxsCPzs
waCS6y3WoQB/tsqZGVwEn3leHQSTQP7DmLhUvdVcyE9z4W3chGl9E/fyA+650TC2ATFizRNMu9xa
Hry6XbaxmTo83/fVv/BvCY6Bcv5lneSm5l9PZFlD7jeMpE8wa1AbXLlFC7xc01sdDsy1bWYkKllJ
Y0/SRvZiXSyT0sdHb899HnVESdTvP0YceV9+4dFWJHALinQrsn5tyJ2rss6SZMwsgBpATmosH5wo
1BzFeMgF3vp3uq2/dsaRNJ/P3BhU7oa4FEBcBkPjoOUpbOdYXEErucIG5XsoSDfnWRsP+kIzqBNK
GsY+QBegYECL8mPLjA+nkWqI/fQmP3HoAQM577+QYV5n44okYEylss/89kPiBS6YcYjuLkGNez+2
RNYGJmSfJa1QwewiPDVtqhUkL4f73L8tF4w8cSilsqnhouP2V3jHFUtk+KqD7Z/MYfov7QRdr6Yk
zpz12xKPKz4CL2zlPwUTgAuwTYUUnoYTG7qIngtXAkbylNjIrtou0NiLigXhwodhRMnw2Y7gZxok
xmhrj4tcHDp3EHsd+k0gV1ggYZoRv3LjKVQiE/NzOyurmoZpcJyufZW7YM+dLIINbih+6rQ6H9PM
KHvPI5hwvTIq6grt8piplx5zLeVhn85p+wmVLQADz4KtZb01Zhx7KpZkVRoSVjYN5mvt0vkbBuOp
gKsujFhwMWU9JENXtSTxrEJyHqYxqxjO9XO7fAbsRajxKrX4UeUnBa+nhkneiRP9KlhAcQpB4VwP
nZ6a/hOfFGn9ucHe2oEX9ezS+j6lbt0o9fwyKJfp8T2XGQPbBs2lmp060Z09UWGvCEUOIxsyKOyz
2rvvbCeV2jidO6+kksfBbKoGcYlDzjcqx5rzSrDeIUMG3+LXPRho/tMNayz6KNcpIKQlkROmO/Ei
wDbirtArDKzxDqkweDRLWq5xy7xg8HQ5BCNFPpgzxmzXz8+FRF9n9fTemNW3v/BTyD/KwTIQubaT
5BZB2+hEtHTTAZ1OfavoBjAZhMwwcU0MKsypGqFASfoIiFXPMLQ9kh7Hxzx3GxYV/JOnaAWyJkmb
b+WUrSQxFXTBRLs8MpYScZWlGGhWTKi4cqEWNG3ZtnQG5xW8iPs2SU2X1O7KVb2H75+5LCjeWlzJ
VEzV66oitkXB+drJ3MuxAjgfYMVGGnwh9kNiPtJGFM2ROx19PNQVl6jU9s1DwDBASkcqna6R62he
P8OZ0/uXDezxNJfy06Kr8ExWH2LhxjQFOV6jtz+3xPOjXp0NzqJMZF2YzNKL0tqt3Xp9YlkCrUA/
swxyQBugFUKKy4R3kD0y3lK7qyPVitxtJJn6MZ19kheWQ8I54rsTUYkC8ShmNk/Qn1w+BtoMaQNe
NIImOvDC11+dx5IC3520BFcFlne4rJuaXYr5Wi+gRaU1bqedNqUFydnf2p5LDczr993bgJhpnQ8B
dTsc2NNsrUrTJkHpsFvf6kLhbYfLxFuNSpyA1uH5tBGdimmShw1XWZDrEM2cS6hXUbtSa6gzoF8M
tgkUORtjXkezpBzFO5C/71GCPwMu/OTh7YxB7s1cKVxQ3FBVzU5c/p+aTlyOwJgv2VBiEW5VgM4o
ifk0bFz7YISzL/TfNkoCl2z0jEX9M0vti2+e1GrTpNfFg9FydWP0bjtTGPPTtLWRN1bI1QP0uGtl
d8VKH4FsdGi6PDWC8ZAnSz0aXdPupP8I353MmASB9wxuLFp1bzPdQ4Gj1uNBSfyGH6rU9t9DvIg5
4mkw/dGiIqGoHF/qSEw/X9LiIciz5VhocGU6w4UsWI71/a7zRUmPvTEJEPhh0hozP1oikvauCxZU
flsbzCojAh9fC86HAeZvtRUntUYmUlC9UEoOROeNuNjWjfPQhzRDOhl5CIVvZQD86S+RK5lMEg8l
KiJh+L9mkiv5d1E1cplRwCMd5EAcxym8ZPnkNsXqz6mcww12glIhy2vi7aCtRIbfvBot6/dVM3lK
cMp7/WkLuTLtBEW8eqMahacqB2q53VcPzLuufJgnqksjeqU/rrhz8sJsTuDPikA4x7kFJeL1RLPA
q9mjT01ZC+vJsywjAP10RTiva+vA3VoS/EgESYZnidznX3NcNRPsg6yh/uS6le5Gd4KNs8EbX58t
Tn3yXsprTeuacKVgGh2/MeVkBdL+f42hLLFmXi23o4JlY7vfakwDgwnRrZTY/001NaeB+lJeQw5R
uWZry3G5SixcJZT7Ax0HIOn5Nv88DUtth7mFMMv6RMyuj/LZR/lX6b1ZhVblp+UJlmWu3X2q0JEE
JjxqZ5+XLqQLb5JzeXTvDdQEIFU/nQYfmaoAAPUpeimRdHDcDcGkhThk5w6XVb7OYhO3tWB8Daf+
yefdRk+mCrPG5V3/hxBwoFa8J1MXycyLLn8urBjgSHoC51NKbgMB8GSI+KczbX89NLsgkUpLBMCT
HaDIElbflXfY1WMid68vgDAHnqUdCGbcke4C1xR4pIEUWoAaHmeeQdGC7EyUyqooH45Rz83ZDiX9
5BdTeS+uPi2bTRYnXK1EYhnrQWS5JWiNA/QaliPwfxR40aui/qOhtm2ZALiV81ch7t9O92f9RC1f
cXty8eTgCp/MrY4LDmcokaVkmaHLP1if/PWznNa38oIvnEhSSivKUn9cT6g2vmmHPufjgAM+8bWi
mtl1VC2hCOb4sXPMcQJqqs4tChgNktuno10lc+sSSFDPCvrzkYVPW54MCpE9BGSbKweZPLJRLdAC
pq1Wec1N9c1008e606JeoZANKR/HcZrVsP3lpiOVPr9XLXWZJ9VkoW9g6kKgZiqOED0h0/cB2Dqp
q/S3b1963o/8/Eq7+HP5Y4Shd4nZ5tG7/ssy3Ih1L3MLTfj+Zdosqqf8Ryq+BBnKnsdytPKrgsUR
s7jZ7YvGvKSRWNOabQJzsRKI71FMf4ZoKK2e3IpMsSf8SH0Ncu09/Fa/Jf6GyMw0ozouMhKWugX1
aExDzQXY8Sr3frhnldZ9RIvKJyvdvLeNewE7uHi1jL/GItkMBNzOagfxrV9f8RpHf3SuPcpJaWp9
XBtKzCGbQwInwXU3Kkj81oZL3cCXPh8tWWzmvfW9U1ecI+aN8Awz5aihFmqcXwktG+O/lD0VtiIH
dM2PED+ZW0TDBF/UqiWMuKVmlGDthRVlZZlkmWev5kwx3ABMWUEbHCi6ehKx7EcHl7C07NFM52XT
7q62nnMedgv/d6WWz4yuo109RyxdgJw4rpmY/frqKhQBUNJ4yZa8Zyy2pME26US+frKUFXfOh50J
n91LzIpPlqOG7UpQzhIr7gCEB58m8JplGck9yOLMh/is+VBf54YsjhXqUASVgYq/QJMA6uASNDwR
Wcu4lQrsFN0e3V08wQuKc1PE8xk4seKj6oai3Rddq8wME6y+IQDtQLlEHpK1DJaj1VlifF4olVLx
ngblJpAY+R9Fk2kJ3AAXpwJKBHxEUrVHDcipFtv2GZZPiWXTob8FR9OEQIfeQ6nuYpWWi1A/+8OH
n9fQfCMuep2JTZ95N3vv7xES18a8KztHggV8G16chUqaHqRBvz1dV6lR1plRMq7W6ZbNIJENYtQL
k3kp6ko/Xs+CMmNd64K5K35xWI9RbJqNFI5T/TgKD6nKVLaqlqJ9QKvnMFCzULMOl/6GEP8z+s/p
u5uDqbJMMXZk/6OTvCZSIS9kfb1xZLC/HOv4PDP8Pz9fUnWUIJHPwVqX33DnnfYkHvoBHCsSV8w4
CMIAG+8IkpqOoyyCjLU5UQtnJ4VWvMAuLGRfcfFvzsLZ/bfdJa/TOFXTonkDzm/hePGAjlzVbi1n
3vcax4+NtSnwCNDyMCl0OjIkZjD9yAL2ORB7Zxv94B/Vvvu9sCJ1cj9wpiSXpQIkQGkKAyT9Nd0K
OiGeqM5utTRJGNuyKqqOL03LnSRbStvRSG6Wkg/XazP3VoVT56ZO/C9My5rPEFHJUlM2hytb/HmS
Ljd4g9O20V4ZZXvKGEdlUf+PTe/GTFrqMFhku10tOEVECDD5MGjXJSTFeWS7+qJcBe+l9jBElu0c
/CntuV/NwSvHy3yd2Ts/pbrDvEbAVEbk8VSL2q5g5XECqOY/TeVqoW8fbi79Z8TgYPGDIj0HJcW3
MpRTkEqQkYaGocBWFR3fKW6OyFwAvz43cChe0a8wQIh1zTaKkB9lkFLDqB3gmBIpG/tB4Tf0BRHO
krOZgp+qPJ90prsQpYOW1mmYp7OFsutuygFZ4epoHXApfK5BwBtZp1BBSMi3brdZGJ8kFDqR99Am
LUn8QwblZUIn6Njp1Qp8RgcS58x9dIuEL10zWtRvT4IdMH9vYkvbN4Tb/PAl+BFOBOSJ+7luM9Xp
PK1mIN3M4VoBplgZOESa6sMtrs8Y5gPF6VchX/lkqovsrxXT70ny20U1C/aWcWYQepDnWCKCWvHc
sZFGFlaf7wTojX4ZxSjV7kk+zTN/tdXK3BT4XAbu2Ah/bpDgmxOxmDPU38E9rxpKFOfWEmHX4ILn
+Z0C3riBDDQ7tpttOxFuQBkM2F3XBZkso4x9Xz8Zimftec7Un3WOfc7/jafysVDT95BaH/wQPUoB
a2y61cpPdqCCH0rRBggaK1eGX/ci1w26Ag3ueGf6yA1TIuz0alofKuoC6o3cBlI0z0Jrt/KDy6JE
R2+PNVwUwWruHl7PZUXMITfTvUc56ORGBm239sMtcVXpihcHh61rTsbVMgT8baskJNoNkeWTAFGL
13CNvXRVY9ba8+srLGSYga3ZPzKTSc6p8acVFUh8Qem0vHKxzCPHLSbQPf3UZ6z7ri/sFgWqDWXK
v3disSDOA36i2THuP7JcFlLgkGwL+ozz6OuOSGldtUfbAoMkFJrXZKKGeNGtYl7/pRnymt4lVYg9
X6cWEpmXiA2kqy+KkZK0JW2IboPRzHYnWFES7ihnm8mPVrGy9M6TTkbkcc4vHIaRU+iaPVDzZUTq
tUM71zkcOxvF3Dj9zIAt1g+aq6qcXQ1mkmroQVjQSl2idH/3IJCDMjviQ+Fq4pAYj/LUsl+kHvTU
4AGu9huJADRzDcnuxEs6O0hGgWe509UuJF4bZkBtUBe4w5VXJDjBLGL05l7PYj+nqm2sacEzyZrI
snjBoHvCZQzhqc2NedUR+dnf/XRfYtIspXhsm/hfhlgxJ3ebpBqeD1pl62NSoFxZ98Mhtno34X1b
UNch0PSFjiSJFIyz6JezrJYiduuizvS8d3zYNbypTEL0VzA/NUFDIT0fq/MSxoT69ZX6Tmrwy2B/
+YtMGunmTZbVpgyf3LLHP8UU+MzAOdOxql/TFBtu2Rz48xgAe4FSq1BT0uvdOMj7ZFB41llojkvb
nuaQcvN1rS8qBSJycUs8tLVsR7mWENjDegJ19zD3tdUyIkVl5GBGxtRVGQbIB8mvUze+eKKlYBeU
KCt9fdTm2nnEfUmBHHRL5O6NX4ivY7qCXytNM0iiPMqRCiehWrL/qTxzMf0Z9rAnNxDpW3Rx37n3
VRi7qZyKIXBrhv3CAcXAz8vPakd2JOUDZWgb0mR8iG4ihNJVaLp252Hyy6SHqGLhoF95fnLDLOJX
J4qjPa7vyovEu1FsRXeIjepbj8EyhKjsFSdDpoLgXmAWn/EHMkox3tRn54kf/XUivzs+R5jCJLxq
WqCLaV6czD0CDND1jn5jB+925s9OdOGUKH3pXcHjbErgZAPdxVfsPT46SMJtf+u+AYXvr8jYW3KH
Whttz13eaouA9nggofxuRAN/fO3qH9+73QGv7UNGPtX4kgOQJDXb6Yuna7BxW3i0Fpr7BeAJ/Ktp
nB5ayVTIBPa7H88uUlaCqKtbtbYbIJTR25sAOkHSyZDCt8Bg6eSJSiXHnB4VXOqgE52a
`protect end_protected
