-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pq3iBwBn0Xcu3jN17fmPqipyQWrqBciILH5HPGbHp9GbNgxw3l1J2Rr+v/bQkyFqAejiyQS+9Qc2
tzSvJ5/bSdeXUhcfrpSXOE+dRsjLfDgjUKa0wOQe2ova7iy2elv28WpNyw8l6iJWErmhaKZ60Q18
aLP3nAuAG5hoO4zLWJdHfAf5dF6TMxJdisDROyzP0D9OAp+BNx0nU3Joc53XErcv35XH2vKpalRi
RQF8HAqUB2qgCvL62ab0Ckmi8aEocv5tmzOmQzvWm7XGTu8zHDDyzfrxBqGESEeoqGBBTInbERKv
QeCWggPCTMEIETgr7CI5FM1h+SQG9mvn7axsaA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10736)
`protect data_block
eQzEjsxWnPW/aJG6rCc2/qzcg/5AfjHn9EwR/7xY5yIxOGj2gmzFBnarnjtD9aEYzFCSGTMAiFcV
auVAfO+BZsdiW89ZFTgNoR7APTBX1bTV+p1ksoV/H3eY4PBzOjS1ns+POgKVQ7C2nbOr0lsei4tJ
NvTbuguK2Tjuq8lNJQLamE20ts80g62NvLkdNL4joi6lgdW1AVMjFDG+JcxF5bIJQujxbcbriKGh
9hsOK2DImec0Zqq7wCPXUA3CZGQX2U1spZPR0QUleH/KPY9SXKFeeXJ+bXBC6EwG/S891MZwqdzy
o5d2gUJ1SnkGhksg5U6zDBuHcefJJ+N+IYtDPsqTRkSgBllTimBd/qC5sakkdUcqDNLsw/f+tNlH
q3Fd4fGcnxr5h3J7Qg9+ruWp0Xba1odZnNMmaKOvdvHkOOn0tIK1xnSrsfF0ClTs4n+qmjedcK6T
0LVAWBYYchmtvjFOh/PReGTeoT/+x2332qnXStkb0st6Ay1uOpUHcCdWbPFHyWkPb+i8PrYExtYz
tqBOvbkChJjiCnoddTjh2tJx7XPzzTiKd0lGgcm20GGWUAfNZ9MnyRJG3NwyMl7XkGGLe20ZViPj
i6JhHfLYYfhPxQtKzW2wqPpU5NfUE9gk9TyTBd/MVrqZC8heCZ4vp4QSPTa6SDz1PrJQ5AMriDY3
a9NOW9nASixFqbphmP1/Z8yiOQQ9JPD/jo+BTy2J5bqKx3G7Hyi1+CmRuJ4fs7VXsfF7fo0p2S/+
4Pr4UOyfG4DAPHCzfmONjbuZxwFD/ZFslB74zlCERTac4NhSGT1q3xvRYuzJBHJPdlLBlOWJbYu3
1V6GsrFFO4iyfHo5Mp4r7vF4+FDzHSWMexoICKT496XblqrHKYyKaD0+ihlwt5Pz3iTnQ1YuZPb+
sCYKRv3C2y3h2pjs0KORyqg9PtBX9cZA8iHh86N241V93KHryreyiprdVEj4ZeYKlFq+wZOiq1W4
9F7TrBCXNKLYScD4mXaBVwPexY1zdpBPYcGBymlpftRp/Cd8P8I1kaSorU4Ue5GLnlprwFaidQFk
YEuDK+O7/Da69rq2Y7TfMqINGE7TnPK6YY09xBDieN/XNsZqjq1S+qIENRRWCeaxQUBMb+7iWMbu
UMUnBQXjsFIlFcAhF4qv9qmLOJpywqHGYOKHPgTrtlvDHvsdThunMdh+gaxz87yvqr9FX+F8Max6
N9hAf1nYx0cZxPCa90ls3Fwn7nD4HNHOW3xddYv5kdP/5fVmjOzYUBARD0QAppB2shxroFaIBO3I
rLqyLho9mZ8+ObXTCUYkDTsvTMwNJ7j1tRWZ35bUoW2PhmdAu1OTMnDR5sTgpm1SsfAIamhMX4np
CVKcqJ+5RoTMEDHax1Pi6+QUddh9htLJsYBeCRQU9tgN6kOBw2+0sLU7sA0U0yC3TxD/ZyvY+B5c
IeKu7KmcghqzFAL1PhPG/iBsvXWLWfmKGGSPf+hAMUy5dvzzx3Bybtpiywt81NYoZkZkJse3JTb6
v0OmOW7KnWHjyDNE3t343rRrNgS4xTEEKV7x0w/lLiZIiyV7u5lGAiEepyiQMl0hG2vwV9uBAaPK
gfmQilQp7LuFJF0beIYrFVqo2lmYP5s6za9wid0eIalWPAfoF0K7tUOgnOaUOmnAlPs+Ym3wMpRP
MXLVLUO84KOG08s4qv+IBnpvEjWUA8S/lN3/DEVomdssp4mA8zkqHo0astal5Z8QRjjG4y+PlweA
VixXnBYtsIP6kaeXt9fDvYk8JmZ1DCy76IWQVh325gbJIHnPGkP9LjvXnQwGZwIAf0p8sgZAdx4W
RBZJj5wY+Pq7cQlk13vyIGlt4TLcBmiG0+cMCZOov2Ih1BJ4Hectv5M2xXIO+zN2feiBD7XaOkjw
pkbIET0L2i5B/Xekg1V7ASe+YEKI/y1yGzg0LaGPNB1OPviBypzelHqbMvC9s1kmqvX8bG5UwU1+
Dr12rZ592dmR/VqzHQCnZDWAerPd+ULNW8TKe1f8JZtgh0TaIozvXbCp3mJQjxghJ2+Y14uzzTlk
VmYrPxCP0cY67fAaMNEPM8CgIFLOE6jaKTsHaIptTEv4QDPN/syruxrKfCx9xfInayquGoQxQWn5
gUPhi52Bwoxd5DbtxMUW+RhesOE5xULpyeAzofR/HN0Vc5ZF5A39SAb7qCAsjxD8s62knthjGT3B
+Nd3RT9mHsrgqgEawcfWx3F5lLkSNbiAep6+bsGrI4EpHbRNmJgZFg2Rj0F2KzpgWM5yeYGfAL0x
a5MFpeuFXsUxxWuD6pdEwQGnnu012LuYRITAjIA8XcKIuR/vMJNEzgcd40Xyn8pJBBIpVz713mda
05KLlNG2ItJSbMueq2NDrHvYWNj2g+ImujdBEVUzSGfahf5nhaKt1byfBTwjI9PdTCNKUowP8PJ5
Thop1p6NDiUlT5HB3L/lNo6PDaKV4KPxbaDGJN5B+rcC8k2DFF4rs0FaHGZypB11ZbiYUpomLebB
kH5+ZeWkLXEwugu0Int6Lz2IrrJ/s88JDAaHXtckf6+uAkcPLBy3ZxSN6E4jtaM1EzGxkFot9ioB
sYdCUrc2PYJmcS1yMhkOa4A/uGHZVegoSXiC1EduRvminPVdE6IVw1wo314L769uzBrPI1+DfYZL
Y53btTA2j5yBOwozu1bbNRX4MYcJc8bjfzP9lq+ilLMb54gymQeRapQXzdRyKltqOJMA9EJ+rIIG
CC5sH0BkRUYaaX8tKRlL2VtmZ2aTAfUu5/z9GNIUZ//0h7tZNmYx+ZpYkO0cMv8/allSqeCkyR4A
yKR9cNBlqeH0XjYGC9rqLPPAwsU9PGyVm0Ewb0GwoDUMhoGDXtpdbZXKXoMb7wivNvSsUlnd8Vu5
80IkVW4DpytOxGQ3WAuy3MwtarrxosHzwld+QPHcrhCDx42wiBtrAleA+C/6SR+o3M4vqurQMhYA
NeS1ShyPRNU7bAn50DCMtnP9crbJJb6haXnbZytPbXvBZn7qw4WthScRWpq8CySXiuNyNX110HDg
muqfL0wxw1nwqoOaPKEf4zulEqa4k6AsaHNytCY9QtKQqy8fxDyMyxTWWFRYimCTkPAdi+EUXrlW
105JrjN4z/NmK3RsYeXJvJgT1tZPhCI5jwM+19xcNeYDEvGDF6K97pE4LXQ2YSv2iPLAtvaI4L9U
P/QT1VwP6NADCekAQZBXqX8kVdED4/FOKK7z4CeJMk9PFVPCKwyGu8ErhgU0V1RDChREpCzHj/EQ
yLml1U5yGaKKHbRtr6trgaiK0E/J6S98bR+92kwNJuthgMIKog9jPJIRV32r7wC63FHnyEBkjl6r
r8kBJZ/mpKAeKRUXMj3JNSk3aSQOevb6Y11z8M0PntpdDiRVrM1ask+/BQALHI8V4e5p1nrb+z2P
NrSGJqNFfN6CD2d5WkQkeXi/f9YGtG1YdoyEOCf0P0AFXsbG+bot3Zh8hNVuvgP6rrEsQcMBHmpM
5vepf/YUSRDoXAXbjPj2C+KpGHgHb4IBU1WKHXvIjM9b+6JC2eOnLRw7RU6RPIcoLL9CEcaBfbOE
sz4kfZ/3K3xVmry8AB9SSj8Sfo8N0bbShrUBLwl+CtLKQ1BllC7gk6CPbo+9I9NYlRIYafkJE/hj
jxCgVks72JJhDj+XbywFtCuKm/6l5nCQjExrijnLDmtArGEBCh/ne1xi+Vki9JJe9LyUlmKtrZOw
/mozV/1IY3B6EBNeAK+s/rYVkc1UyXU1wcoc9nmG5BdwUJXKvi3RdKP3clybuY5+RWD5boewpwrh
bFf98cKIzTyeGiqVShIMRD4yQ0fpJavkZ1OpClNzcJM40DL4ADDPxZWsovZ7agHj1t/DKDSXfAJS
I11MD1RG7Jf3t70bTb+CQZ8dC8rduEX6kEVcotiRER0PsTkg4SRZEWRsA6FObF6taA6CAp+xaHSB
qvqWRZ3xwi82Z/fztsUJ2o/klzmCIPnTwgXPAnzFRsLjhUHYbE5DqssFB3psKtF0msNb7ud3o1tm
ZM1J8hwHtTYJ3QNFHMJpynpczS1+shVYbbwdVy9Rp3iQ63NIpnoMNBFAajP3s77a8ncToU0ESUDF
ZQ3wo6yN5O1xaG1ZChM+TyGpovvhk4KflsUFpbEomgs9T92T4J0FHeMSDBExxb8MTNOM9UX3I+FZ
duvK5ESOuEUrB+IezuEkQYcfCdc7HtdcceEjf7qzX96wHbUXxDJPWTdz4ndn5izxlSQI9B7f0H+6
WQ3pAhYQWtHDzLQDdVjGMqMfWTxZHIkzx/MItkMvLhdLf5q3B4mICHa9rpQfjp94OSFdNDSLNCvo
Pe0LJzt5etuP5G/CYusoQpj0gtK/yaosWbsInaVDatxyRDbSF+6uAOQMxy0I8t4AHNVR9BFNkfXg
PgJ3dZcvO5Zg4lLSdl2coNEtlA7ZDajeGrgQvS313XtToildXV461FNXtDsl1MkZcs5NzqCIRsre
O8vHB+odYWjYIa9GB94LdKWVrLY0Zgh1ONbd9ks053/DptvdTle7NyuAArov1B2UKYN6X/9qI0yk
Nwshc3r77eityieWLjJcnVALkMNBd35YIJohAA3w4s3ZQKLD7JViXv5xB66S3r77pueEKU1B5c9c
i5QwNWmO7KsH3PDeWjAMp1RFyOPJCIjXG5Xd/uTMN1W8vD+nr3FdfxK4RifZkitYqAbu26ZAvb3t
9pf6Ls6Z+QPJAnZaTFYUURINpJgarUTg/lOobHkKWMcODUXnZxzwbW4u1P2PQ820Ez2KUekPFlVL
nOuHhxvSf/71HGbPUNrEvClEMPCXt1FbQhYNuQI+w5Z/G1mE9CDuLlSf7/y8AudbcWcwyw3qBWzx
r+WfYy8xmnPr12c4/53cV0VAU3gdAlz33pbaL5JHx/+qvlv7MX7+6JZBbH+pnnQ+01n8RRXiVece
qKNV9VNKF7SsMs8OlzZU4QYyYPd1XfDCw2wACovv7K82OcqRCfh8VxzH2AiCY+eNnHpaRyntjcBM
knJJWxqFdLcmvpc2ZburkVO/UNdd84+5gBp+XBK1bVPLp1N04YT8WSxhvfh3omTtoLf9h7YrBN54
n67owebT5aeOt1R8AwxhaO6ag8TjsTTjM6qY16XHTJ37/jHbWRfQg5vjIK2eiAIT0NJa39E69hjk
bkKk93N1dbXXQ5voYGaxZb8A5SQrZHXKbtr77RNe8JBIO1Dzaz7sJ4+09RoSPknPltbhx3+8gqdw
PEd4ODU4YuwhJXp5ZCjxq3CfAi5lNrt10/qUiOZCqo+ho09NSpqUEa0zd1eVkN37CBTVwJ88bkLD
0h2XP7e4FcsLn8SLms5f7yMC8sAcbJ9eN4Wy0L64cjtSG3qEKT9ALjUeHh6FsHb7TV3s9EprUvv9
S27AMBDkza0KfuRg9fHCg9rOTWkJ1KN5HeFh4e5RLoskfKm1QgA7bIzcLtIP/S+mv+2hyA370YaV
LS392ED93zPoKrTgQqCPDeWtvmcOWoV0nsWBSKC98L6XyuwshIJimPt2gWdntTl/05XW9B2CUmjY
4bop32fFu3YHRhYWB9va/HhwvrQmAR2OpOVIHF3r+6S3r4YfoS5KBZWYQab74IgZLiNL5mFJN1Oj
EngE2OivvhPNLqnLs32zp7EGcMUuYC8XIZrDDQTK90ftGd+B6amlxN4q9h90OkUlcydm09H4Vdmp
wB7DUtcx+8aNWcENVnn0wgWe0dNwk5FV1l4JSN7ll0v0QzdCmIbVhrt1Pq/q4TPVuL9PAMAOR5kp
zVCgCY1sSarm8hSrwf/7TIuo/6n7Ym/4eci0pFHjvArefgE5AzsLRKftp3MKa+togpUD0jdwq4u2
EJIGXm6fRhfwXn+PMtdKtOKiDo2/glgLXQNPxnBN2k1nJQ758cW4iF/xyqBUK+ADlK3cvQfcM3vn
rx65jvpQIHCTc+BtpJEVDV2I33RPwYMpBmJIVC8AEQPgCsq8OXqu0c/hWVG+ZSzbdUaDbowQ9gun
rcA7F34ot7/GamwYMx0bdTbj3hImDckb4Vw3rCDHhHym0g/p8p7W8QmmoYWBEZqRK5ZjfgFvEq49
frqHT7jMmu7/sC0l86ccm1fvv4Ur78OtgxRCXIFh/4inBCys9n1iP4W9q10q5ZbziaXUqFG6UWDb
9A/OzfWi7Iv1HTuKYxrjnr5cMGI6DkqDA2x+PtbpH1G7pzdIHniHfWAmJknfkKyiQdMl95v4NW0q
Yf1qqduEgVJj4+rbb7VCNAnwQxcqiS6cWnzrEeNIC8rsbSj3nvKl0Egn3EJ1Sa8kOwrO3iM4j2T0
qHd8nyC+MjjE3c7B1OuEgomtNziLj4m/hNJ8+NiR+V7K8eA/XrFvlJh87JWCFXrJrvGaNiNI2Rdq
PB++35SB4dWwmDB6Spll7gpGyVrk5W0U2y3KL2/4WiLSwnv7SdllNE06tnwXxMH0Pi45R3EMVVv5
jqaxzz5RUIS9b8N0euZVIuWDrdGSzqC6IYburs9XW84E/Oenk8LIVevYg4naoeqWw1ua+rsaFpe+
krQ9N1wZ/T1HxH35GVYHOEeqhnTLpkqOJ2hyRhRjFm3tuDHgQmxJtZBy0yk7g8FXKq/svm4DQypc
XDkInzUIP/AM7HYmfDtMP8Dy7VpxIHR5u3aw0ntJ8z/YQYz+UKiug5Itd2lnLzeucXj8g+KXo5qn
5nRQmA1ry8nIu+AioNFf9wbMOSM+fRntT1v8OeRA0AooBF0/aqrRvnVAriIHrOD3dvwEziD0hR/S
WCxca1PT0dH4vJx7i1jZFrizBrPMeeReD9IOLfYywDPqixUEPy/YdURqddezee7R6D/9ToDGMLWq
ZPoMHES6BqcO3eS7IF19fuuIC0HoCUcvF3jhBWtPLUguIkVmxSxz8G5OqWUN5IOABBQ/sN26bXzr
26XJlPFNiXhPDa0UcV5zxAEXFpWHEWR4+C1r7oD6IUyD6Yzxwt6rVhd5/2YzMdal4QfoYfXGXMTi
5PzLzFTGxbUJR3R8U0TF4ENS6l/Z5VrlgBVBM+6Sx27phwSVy/crAlI4NZOvu3dySYyYSwXORsGt
vScsK6oRIYFwPgWcbUmp9k7PstZPNe9Qf74dBjJKWg+BaUtfqYDHN3m6PecnPYwmUkZV7doNlYCV
VjLajrX/rLI257pNUZQM+wvNYfNcGb2WXGn3R7iEKLKsqYmyLQMaXpPxlzBVOv4Zg0AjDL1F0Z++
qu9tVfOoJqRsNo8SSiV5x9H/mjbPQBM6XMJ5LrAapBZIKwkZi9TpUU5sFOMwCKR9rjNnZAudBrEZ
KtPKz6IA/JbMGGxXT9bo8+SMtDiXhrhweU13AUmfHo/zL5Z6aFP9AKaY8Nq4/IfQalFpCOK7/o/w
Fu8ipKUdVl6ynqVJrAcvqbIlrG1qAcweFo64FCL/n4L5rjXZgy59oKoyvoaWCq9/8vHTcd/8tfYz
JY0CbfjOoPBSBBcG50HqXIwZVkDJD6hkcHRUOk+sqMQVI014rlxiw8lG1VxNP7t2hp20GeJABTrN
EUMnkNOINdydzn9eUlyVZb4FSG//ellhFZv746vMK14ei6SZ2zOYgOrHLQVNcm7w/QW+TW6ARmvW
BH/sGOns4RGKYqlzHgFnDZzNobbplbUldojBeuPRHlGrkKSOS6YOs2p2a02fHWdxbyYBPx+qcamY
I/BaTDfRxsbbeTKnv8RYfCAbiEJWO3ywYmyuWQheMlr6on8Jg/jAaPLS/6cLnqnh678T9MRdiMFw
Inp/a/j2B1TbIuGJV3XsWxFIMkRQOEynYpv2xUtyECLshiUiezD7ADZyv5/hRd6tHJCQVRqvMOtM
rQYXJUmjj5b5bnotTwrGsWi+c4Qov78lNfgRw6X+a5Kf+1CNgrPaXrRwsy0mCMSoYHl4uGOoQbt+
DXZ2zNG7pqN4O7Qn980ce0h2eKnBQsOqf2CMW2EHEjhFMH+/A57KSYZbqRelMKAPJ6ORUa5MqzO+
UgGLYWXvMNiFkEtwhfD2spc4VCt5Q8UrdE2jLJbSkgvxgFgO9brAoSh3zQ9gBQ0F0pA/5arRqw/k
NIph06hSGmTko+3eOeISvEuREZFkxQ/ayGegdnF729Z/F8kvV5WKzwXBtEJ0WpOdeyTufQdMVbxq
gDELe6rOuVfHu8qCdq8iArwP/W2QYekS2+T/pwF0Ziq1IW+4bhJrFDcJbCEyx3pR4v/++jNw/Rij
P4FFRO9a9jAo0WSvoEQDDN5cfHezmC4tMFu7hMCQ/uXcH2u23JoluWAlS3Wp6rexHsttzy69WBnU
dKIvxB+QgsEXSldAHduf8vZ8aX3J8EIZpH+s/X5/YirYyMvb3biEUAYF9crv1d7Yva8ls+SK71Vy
7HUg1EiJ9jmDWy/d0nelaickGFh8dD/iRTXNms6cs0TB1RBO6ROFaA1y7GAJqlCYYIf0W+xSAnDl
oAYwO9jZxaOt3kkfZJdsxIL//8MKtBe2/71bI2600UgxSMsBpsydoo6xMmu3jej9gyPN3OXSLK00
5ejmHvq+gn9tGRvSV9NLFy69DeSGPW+Xl+Ns8u26UKm+40O3okfvwHBUECnUdSdaMeVuT7IGv3IA
jaSjMneGU+rCeyiXxpbTwQU2lq4QjAivFp10KlblV57Wom1XCVCdvNQC4bD/f+1b3Ai8Y2rClokD
S6+aSLhuiZ1WLkidzd4//7rD/jOFKvujsXRtbiUogX0M6uI0R5nzQgVwF57D18Ly2tNMwaZosvYm
CobKr5bR2KbCElqMedulJe9kBsa9DgTM7LHwNGZR/4l8RenjhBgmZu5pvNmgAz89w6IdpEsw9tdl
wkc1byOs/DyGlHWdmYSvwxCbO1C9uAs2gbf/tKbMesKKZZktAPvSZrbM/B7JxmTfKDpqu9hcLiQA
t3gIlb29EqVbYJoQB0DaIPQNJTN7w1iRrBi8v5TuO0IWymmxjuQTpdQfUnM5u8+2JTjrstI9BcjK
haVbnBmJ0+ycmqoVzQR+kvg62PgHvjWiK9Azz/6IMKgyqa0QJn3pO0oTUxQnMQ2rkq45Tc5kCDsW
jCVf+amoTFdnfXyhW74p9bJbww+xmveGT160aToEJG3k8Q1I+bLkZ7XZp15pzhoIIRjxOFe1ssd9
PpfQcIJuG9ru/iuAFZRVQIoejUh7tw99zB4iwpOwPZOSTyzhU1fkkdRENVMv+e0CC3JAl5Ze4k1P
DNjZ5ZLC1cEpM13FAQ0sdLJHsKjWsHS2lEJpNboGd3TlfrYZLpJxvNZuibpOgFrgDGeFkQY1EOjd
kA0sMHJyjkfthWkwgfXgPxfx+s9KMgQCYTCsLxBKDgt+qrzEpqCKUYuaOoKy+nBrn+iFKO/rT0bj
82g0u6tyddsMezSbJZ0WebBIl9SVYsVudhtQr3FD93+vn1RrRLfSA509DgNuH0Kh0XnprYjEiY+q
UJsX/J5cuiOxSzd46+2+rJHE8vOscZiJn5l3Zc4GgaHiVENgUz9vyaxcvfhQ5XOOUb7mF9HHYSQw
F8dya+r+UnNmfJslYUZVPyuacAEzL5mSIKeMOA35YFpi85VbAk4n+KP0C5PA7+5HYHaRNm/9PgJG
E6DpbqvVbASPRowtvHlaRo6pB2gsFqODz+HTMXMX4J8Dd+ocshWcbIzK3Lxjntg3dUbp4nALwBDE
4bHVZHYCFOjLt58FPjdJeUBoGcCqHA7MH7dMUZ13MriLE54D2BMkLHvu/ZIQSPXFhtMYsU9nISpV
TBurPlDBsPwh/SK/QRfVY7Y7/eHbvewQ1PudThT6NuzuvuD9K+y44cPQHHSKurbYgnTD/F//8GDy
WaQLdT3+oELcQ9WnACsShJ9SXS8dR50sFbfOYhvj8/1NuiJaIdXqDjyapoJ8NGACyREFUXGFqy29
PmXxvCwP9LJXj32KmSY10yPogLjX4BOZO5euihYoKXUKJy+2cceye+vmgWc7961696L2Smc0VqHx
Gz/pUvBgcn/1oaRksHf81LcpPwP0fwJHCChyT547YmfVOB1Oz4xKRUp9awYeVI4vyLQ+hYmcvNrE
lad9iSxpfxrW2kUaIr8lqj/clSBiUIh7Gdcpji2z4lPiFf3NnYfiAba1STZKifwh+m5lrIDNsg3d
pk24JFCHSScNOowL8/oIxr4LAimkVOOI49B54CLC05WbB+O/4iUhkYKIW83JzX0TSrloLo+juEel
ZH70GSEGx+qrXiaOWkQp5HLCQzTu517acSSth6jYxPuCLZq19YxImJGqiy6rJrtG+oNWitnw3jZA
TGHAOSEJpUIp4IxZBZkUPNekOlqdaX5+q/t7PBxKxXARJG5udodI8UNQNUDDuridygEtg6kwZ0yX
0qECfns59I6UoOa0Dt9W9igrNB2IClrYQouqkfTaq3P1mMPTq78zBhfXRD7pKTmzmlz9r6HHUcnI
IqvZJ9DumjtIjjtDj6QMf1dykEb5LNc9I+aGFU8pHTwXXofWS8TeL7G9FRvUJfRMcQa7rcvGyp5h
iWP7fF9C2xSnuwmPk0Jk69PH60Dew6cRmKWRlNBtexEMazxJmWgNARWJrjvxUiAF3iSLp0CP6/JW
Eze3s72VE4egNGJpGqhQpwnvJpFD+cDjvueBdjkqnSLdK59V2/IxLcUoShqUeTKuyuYIywFevm1l
fNBGaz7ToISPTl9d5D4B6uaiMzm7TLY3mVbrIQUvQtNb8E0iXA2EKqT8OryrWM9I8q0zXcn+v6Rn
oSG2zTH3xxFvGDBIluazCkxyvwtNl3TVGQJOK5koPShva0TWVZVZoZYMgO7tfsbw6Rt3dYfHzkTQ
zuMZPnuywlMMD6t6+rkBEB1au56sCSFN8DPpxEeKqGOL9Z7citgL5KWGXrAld0hN+22k363jiKeO
Yxx+MYUmixAwP6DzPLtdhc8QExsH3+VPq9DJM29TN+4At1e50y5v7nZa2gIrGVr/lvQ3jfCPRgKr
+C6DuMtWEnA+oAVfyYjUhU0+J+pdleJKC16xfng2LjuRkcgEMT5WX8DGXf4/E7Tdgqp+jZyRuFRw
18c3ULemZAkYw4am0mpHTnwgrY/CDA8Fna8+hEu9OU6UggWy0paAc14v/1gFgA2Rux/oE2YbMZ04
PiyY2HHtHIwdW+a7kczs87SzxgCuvBP21VyuG/IhQ4lyMTNcJXW3pTMvZyu1nYy/hY78E6c45Q1P
UYu2ulzmODs9z/pF1s78Rm9r4M0rbhnlGAMe/Ie/yycdWbzFroK4kR6KVOVPIXeLJ/AWnqkACBQV
PzousM+96CkGfDhBzWgXDR6y3IeD70ZFSSuDb8u1aRIiqblL4E2EEh/YRm1vhQ8fVtI+dyzMPF0W
8RS0val17Spai5mzAKKd2H5zOE4ENUiYSiUfUa0LJihbNtGPcC3CRrLutdmdMuKzO5fgZag7HVsj
enTW0zdD7g3shyBFM7QKilwaV9IxJHa9ECDg3dtYdmlj8xWHQ9j1MU1Elwrb5dlwr+2uAqRygTob
xw5dIFl708UBaeMlvZNx/ZldgF05HfmyvgQyng78KmkFJPNGEBni4ut4aVkzdY0sUzzjcufZaDC0
ZeruHnORb3V5ICIjtJFtq4+fmJjO1uA5ykebM4h4ul6uoCx0h3pQvWzR/4ru06kkMWBXcGEjT6yv
bwFWSOUb/ZnQLaYItm/ne6QRY4M6R81eFKjhDORIfRfD2QqYAYpabCr0tY7sHhG4wnXArE11Rs7l
7UYcmccqhAI0XJd1gxhtg7Bex5dQ+4ReS8PiHJ8nUzYaF6obuQxgtQY0ftMxPZq3jEGiEbMj6wo9
ggVXhQ3EjhudTDBUcdVWiIMWBGbGlD0V3mhLQfLRIS09xoCsoBWJ4etA6/DxpXCLm9uz8lOrbryg
2iceqiDxSnbgZYQhwItabtDESjrRfa48kbW98a689hYYf1dGEi8L7o0Yjr3OxmVC1xmFGCyQ3Qkx
NkY8mmKNshh5Sc1OS5AhK4hHf3ODbJoyqUbmMomzp+5lJFHGUKQ5GQUpraCHvx2YJBYWGbLSGYZO
y9oRvwxw9bxZgDDrhgpYn4IrqwY8CjXHpOHn2676sbc0jhI9SiWk3zpX4egYz9AqXzbv1Ic/91Pa
h/VLWYdfKAn/dYWUZXdYMhNqbOBZbDuAME7rQy+wiuuewO+FHyUtzrKkoqB0uW2OfZDkuIKiWVjp
LSTP5usAt6V0GWIKokpcxD5IbxxQ8NEOcq04jndLdC9ud1RotB9zk+cStkWNRQ/jjHZwI0maYMmO
vn3ZiiUw7UB82TWjfHi+rmEtf+IzKqY+5MWiqfSxSz8YyYLCgnOf+5wtY/2gghZJ/6iCvkAT21zf
7OSzu0yQyt8WHbKg7HA1U/w0ykwqhLCRL6IY6ALLIkNOfbPrhr8jUMPeLkqC6FKCSkRJbpSkgXmf
gDFdXGh+t4PUxdXGq8yctvGw5eaZdH1afbRkWAip4U33WvIv4gYx7H0ry43Yjuw/VV6Mu6qFidEV
HsaiQT0yhyPic5Vx3m3p1TPOfuqLEXgJvbWEX3lsqmBoJDe919DSbER0RGPLzEob8JR1vHStGeO7
4oKCN9XjdiCvaL7lppS8+90kkHYf7aqKiW9EfUCem2ikV7VYCYWQNyiMRZ9vygXSGA+cw+gsJ1Hn
n/vLZjyac4SB0J2W82IjVh/EU2jSn+sTOriD77Xo/oe1L+2ZiyTN89pynTt1FVhVuFAfIqxyb3so
rAHrxkoIx5aAl/M0iKS9zXt9v6E8VwKnxriXR4JgESzxIwrSlqSSuveCwPj+B4Yb5//iYrz9tl/6
O5ZgqSE9L71AQLD3llIBgfLgTSHD4w5y7yqkWmL99AWVC47w0KrzIBe8CRivseBeWzY0Rpox0JYZ
A2sZhngLfkToT5eBFtqmzCV6J2URPg3dPXoir6CydknKgGtIS9tU5VxKI+sdJ2OvVUdsdoR+HpwS
7ByvucSnOjZsj5RoUnlNdM/0vLCvfaNRQarn4foqKp/1zpfuJi2tgKIVKqZ8VhP3N2TWDqjPlXPG
JbeXyhPvj+fkG9LV8ttwkw7cmWy6C6sL2P1KDFcTNFwo60rg2dVk5dTDbL2fh50tw521uS2zcO1Q
tOACcUzwixNTvW/j67usM6CJXmDfHA6moNTAm1iaYWrZ12879QwaHbq/LEwNy2VYFEwGS58Jlhyt
37NQbYvKmoSoXCJYpwjnAaYsUxKVtmMuScC5TM/T75Rp7NTFpzJfJvb0Q8gNefF3gDjVDjhdmQz5
CJau48BR/ECTc/o9hLGQyMDt6ghAD+i302eBj3+MCSvVSn3/1/u3fm1fM8LjgtQySspMQ4U1n5lp
OiSHQGZrsI/hPt5KxiTAElTeJShW9DPev2tiHwLiJsrpO4Prw9oJJElxRJZbnfJFuaizvy+xmm1i
VdnFt46+mdYzuclBxQfHQRPb+AJTKYXB9oxFXYTvRm8/Xy/Y0xT+QAJf0MurmfJmoUBQTpSEWjWt
8RFR4m5KKuOQL7S/H2FzJjvwmJPcIi8y2n6hfIcLw1Z82BSbldTrtwl7+xlAZO6hE662dhWCmUxY
UJbvV5HwJMpjWESiNlY5W86riW24W0sA2NaqA8GEO2hpOKOXfz10E6KrN3xKzUNBQ50zp5UtBETK
7ilytHgzTjrx1/8PE1cW89j2by1GdhaphqztofxsyqiXzSLuE7NaYoHjhxFYXa/4UEf4eVbRkGHq
EVUA8mKhBhEk9nzDTC49O9pzydfj2hh7EQrLWIlO51h+7JBym8pSpDLJoC+cjOF+JpPUhG3dDBLv
bKJniUjxZA2xXt2wvAQiDJjB02jEwU1HWtebYDEkJw9xB2SGUoG0nlqX4NNDdDd0Fpqx/D9rMGoL
YI98n3z+dS+gaGIvOJcjTGEwed/OtjVc3XKGI0xdBH7lrwn9uoJkLavheBgi/qf5I3iBcbCXfIFn
bpXYZUfAh+Z/vnklz340ZAbDHDNYxMu22i8qpVRK+C1ExmpjH34a6/KZUWqQBKWkfhcHoMpKdXqJ
kPhGPn/JL9dI4RziNZjAYwpcBbhQgFUipAsdLMDC5U464rRMGT7t9xjEixJ4tm0UoE9O+GtsG2mF
a2S/Q4ycYL9piDbIH7EHo8zVi9Fju95IhSNpBA4aYO0xqbGVpM1lfBEPAXsIFMbadSHMzflqEev1
A3zedhKmRJSwRM3jn1qKC7OQNmOUV0YdnzstXU9yHqwOaEtRPOu6O2ISmEFAKyMLzKqY9q0CExya
m6gZm0R+3Xkk0Nwf0u0ubiHOJiymnxGznTq4YO+r/WqJo+8ZIrZ/AZyt/+kzrE4m2ecAJ6E2XLr8
/aw4GLWfcVLj7AfqvhMuCrEG2Cc=
`protect end_protected
